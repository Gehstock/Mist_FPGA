library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
entity rominfr is
  port (
        clk  : in std_logic;
        en   : in std_logic;
        addr : in std_logic_vector(10 downto 0);
        data : out std_logic_vector(47 downto 0)
        );
end rominfr;
architecture syn of rominfr is
  type rom_type is array (1136 downto 0) of std_logic_vector (47 downto 0);
  constant ROM : rom_type :=
(
    X"000000000000",         -- len=       0 r=$00 v=$00
    X"000000000100",         -- len=       0 r=$01 v=$00
    X"000000000200",         -- len=       0 r=$02 v=$00
    X"000000000300",         -- len=       0 r=$03 v=$00
    X"000000000400",         -- len=       0 r=$04 v=$00
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000000600",         -- len=       0 r=$06 v=$00
    X"000000000700",         -- len=       0 r=$07 v=$00
    X"000000000800",         -- len=       0 r=$08 v=$00
    X"000000000900",         -- len=       0 r=$09 v=$00
    X"000000000A00",         -- len=       0 r=$0A v=$00
    X"000000000B00",         -- len=       0 r=$0B v=$00
    X"000000000C00",         -- len=       0 r=$0C v=$00
    X"000000000D00",         -- len=       0 r=$0D v=$00
    X"00000390073F",         -- len=     912 r=$07 v=$3F
    X"000000000800",         -- len=       0 r=$08 v=$00
    X"000000000900",         -- len=       0 r=$09 v=$00
    X"000000000A00",         -- len=       0 r=$0A v=$00
    X"00000000073F",         -- len=       0 r=$07 v=$3F
    X"00000000073F",         -- len=       0 r=$07 v=$3F
    X"000000000800",         -- len=       0 r=$08 v=$00
    X"00000000073F",         -- len=       0 r=$07 v=$3F
    X"000000000900",         -- len=       0 r=$09 v=$00
    X"00000000073F",         -- len=       0 r=$07 v=$3F
    X"000000000A00",         -- len=       0 r=$0A v=$00
    X"00011704073F",         -- len=   71428 r=$07 v=$3F
    X"000002D8073F",         -- len=     728 r=$07 v=$3F
    X"000000000800",         -- len=       0 r=$08 v=$00
    X"000000000900",         -- len=       0 r=$09 v=$00
    X"000000000A00",         -- len=       0 r=$0A v=$00
    X"00000000073F",         -- len=       0 r=$07 v=$3F
    X"00000000073F",         -- len=       0 r=$07 v=$3F
    X"000000000800",         -- len=       0 r=$08 v=$00
    X"00000000073F",         -- len=       0 r=$07 v=$3F
    X"000000000900",         -- len=       0 r=$09 v=$00
    X"00000000073F",         -- len=       0 r=$07 v=$3F
    X"000000000A00",         -- len=       0 r=$0A v=$00
    X"000038D40020",         -- len=   14548 r=$00 v=$20
    X"000000000100",         -- len=       0 r=$01 v=$00
    X"00000004073E",         -- len=       4 r=$07 v=$3E
    X"000000030809",         -- len=       3 r=$08 v=$09
    X"000007D70808",         -- len=    2007 r=$08 v=$08
    X"000007E30807",         -- len=    2019 r=$08 v=$07
    X"000007E30806",         -- len=    2019 r=$08 v=$06
    X"000007E30805",         -- len=    2019 r=$08 v=$05
    X"000007E10804",         -- len=    2017 r=$08 v=$04
    X"000007E40803",         -- len=    2020 r=$08 v=$03
    X"000007E30802",         -- len=    2019 r=$08 v=$02
    X"000007E30801",         -- len=    2019 r=$08 v=$01
    X"000007E20800",         -- len=    2018 r=$08 v=$00
    X"0000002F0000",         -- len=      47 r=$00 v=$00
    X"000000010103",         -- len=       1 r=$01 v=$03
    X"000000020808",         -- len=       2 r=$08 v=$08
    X"000000CB00F8",         -- len=     203 r=$00 v=$F8
    X"000000010102",         -- len=       1 r=$01 v=$02
    X"000000AF00F0",         -- len=     175 r=$00 v=$F0
    X"000000000102",         -- len=       0 r=$01 v=$02
    X"000000CB00E8",         -- len=     203 r=$00 v=$E8
    X"000000000102",         -- len=       0 r=$01 v=$02
    X"000000B000E0",         -- len=     176 r=$00 v=$E0
    X"000000000102",         -- len=       0 r=$01 v=$02
    X"000000CA00D8",         -- len=     202 r=$00 v=$D8
    X"000000000102",         -- len=       0 r=$01 v=$02
    X"000000B100D0",         -- len=     177 r=$00 v=$D0
    X"000000000102",         -- len=       0 r=$01 v=$02
    X"000000CA00C8",         -- len=     202 r=$00 v=$C8
    X"000000000102",         -- len=       0 r=$01 v=$02
    X"000000AF00C0",         -- len=     175 r=$00 v=$C0
    X"000000000102",         -- len=       0 r=$01 v=$02
    X"000000CC00B8",         -- len=     204 r=$00 v=$B8
    X"000000000102",         -- len=       0 r=$01 v=$02
    X"000000B000B0",         -- len=     176 r=$00 v=$B0
    X"000000000102",         -- len=       0 r=$01 v=$02
    X"000000C900A8",         -- len=     201 r=$00 v=$A8
    X"000000000102",         -- len=       0 r=$01 v=$02
    X"000000B000A0",         -- len=     176 r=$00 v=$A0
    X"000000000102",         -- len=       0 r=$01 v=$02
    X"000000CC0098",         -- len=     204 r=$00 v=$98
    X"000000000102",         -- len=       0 r=$01 v=$02
    X"000000B00090",         -- len=     176 r=$00 v=$90
    X"000000000102",         -- len=       0 r=$01 v=$02
    X"000000C90088",         -- len=     201 r=$00 v=$88
    X"000000000102",         -- len=       0 r=$01 v=$02
    X"0000003D073F",         -- len=      61 r=$07 v=$3F
    X"00000000073F",         -- len=       0 r=$07 v=$3F
    X"0000003F0800",         -- len=      63 r=$08 v=$00
    X"00000000073F",         -- len=       0 r=$07 v=$3F
    X"000000000900",         -- len=       0 r=$09 v=$00
    X"00000000073F",         -- len=       0 r=$07 v=$3F
    X"000000000A00",         -- len=       0 r=$0A v=$00
    X"000002AD073E",         -- len=     685 r=$07 v=$3E
    X"0000007300F0",         -- len=     115 r=$00 v=$F0
    X"000000010100",         -- len=       1 r=$01 v=$00
    X"000000030807",         -- len=       3 r=$08 v=$07
    X"00000263073C",         -- len=     611 r=$07 v=$3C
    X"00000040025D",         -- len=      64 r=$02 v=$5D
    X"000000010302",         -- len=       1 r=$03 v=$02
    X"000000030907",         -- len=       3 r=$09 v=$07
    X"0000024D0806",         -- len=     589 r=$08 v=$06
    X"0000005E0738",         -- len=      94 r=$07 v=$38
    X"000000000A00",         -- len=       0 r=$0A v=$00
    X"000002210906",         -- len=     545 r=$09 v=$06
    X"000002FD0A06",         -- len=     765 r=$0A v=$06
    X"0000045E0805",         -- len=    1118 r=$08 v=$05
    X"0000027F0905",         -- len=     639 r=$09 v=$05
    X"000002FF0A05",         -- len=     767 r=$0A v=$05
    X"0000045E0804",         -- len=    1118 r=$08 v=$04
    X"0000027E0904",         -- len=     638 r=$09 v=$04
    X"000002FF0A04",         -- len=     767 r=$0A v=$04
    X"0000045E0803",         -- len=    1118 r=$08 v=$03
    X"0000027F0903",         -- len=     639 r=$09 v=$03
    X"00000277002E",         -- len=     631 r=$00 v=$2E
    X"000000010101",         -- len=       1 r=$01 v=$01
    X"000000040807",         -- len=       4 r=$08 v=$07
    X"000000810A03",         -- len=     129 r=$0A v=$03
    X"000001FA02E0",         -- len=     506 r=$02 v=$E0
    X"000000010301",         -- len=       1 r=$03 v=$01
    X"000000030907",         -- len=       3 r=$09 v=$07
    X"000002620806",         -- len=     610 r=$08 v=$06
    X"00000096045D",         -- len=     150 r=$04 v=$5D
    X"000000010502",         -- len=       1 r=$05 v=$02
    X"000000040A07",         -- len=       4 r=$0A v=$07
    X"000001E40906",         -- len=     484 r=$09 v=$06
    X"000002FD0A06",         -- len=     765 r=$0A v=$06
    X"0000045E0805",         -- len=    1118 r=$08 v=$05
    X"000002800905",         -- len=     640 r=$09 v=$05
    X"000002FD0A05",         -- len=     765 r=$0A v=$05
    X"0000045E0804",         -- len=    1118 r=$08 v=$04
    X"0000027F0904",         -- len=     639 r=$09 v=$04
    X"000002FF0A04",         -- len=     767 r=$0A v=$04
    X"0000045E0803",         -- len=    1118 r=$08 v=$03
    X"0000027E0903",         -- len=     638 r=$09 v=$03
    X"00000000002E",         -- len=       0 r=$00 v=$2E
    X"000000000101",         -- len=       0 r=$01 v=$01
    X"0000027D0807",         -- len=     637 r=$08 v=$07
    X"000000810A03",         -- len=     129 r=$0A v=$03
    X"000001FA0227",         -- len=     506 r=$02 v=$27
    X"000000010303",         -- len=       1 r=$03 v=$03
    X"000000030907",         -- len=       3 r=$09 v=$07
    X"000002610806",         -- len=     609 r=$08 v=$06
    X"000000930A00",         -- len=     147 r=$0A v=$00
    X"000001ED0906",         -- len=     493 r=$09 v=$06
    X"000002FD0A02",         -- len=     765 r=$0A v=$02
    X"0000045E0805",         -- len=    1118 r=$08 v=$05
    X"0000027E0905",         -- len=     638 r=$09 v=$05
    X"000002FF0A01",         -- len=     767 r=$0A v=$01
    X"0000045E0804",         -- len=    1118 r=$08 v=$04
    X"0000027E0904",         -- len=     638 r=$09 v=$04
    X"000002FE0A00",         -- len=     766 r=$0A v=$00
    X"0000045F0803",         -- len=    1119 r=$08 v=$03
    X"0000027F0903",         -- len=     639 r=$09 v=$03
    X"0000000D002E",         -- len=      13 r=$00 v=$2E
    X"000000000101",         -- len=       0 r=$01 v=$01
    X"000002700807",         -- len=     624 r=$08 v=$07
    X"0000027902E0",         -- len=     633 r=$02 v=$E0
    X"000000020301",         -- len=       2 r=$03 v=$01
    X"000000030907",         -- len=       3 r=$09 v=$07
    X"000002610806",         -- len=     609 r=$08 v=$06
    X"00000000045D",         -- len=       0 r=$04 v=$5D
    X"000000000502",         -- len=       0 r=$05 v=$02
    X"0000009D0A07",         -- len=     157 r=$0A v=$07
    X"000001E30906",         -- len=     483 r=$09 v=$06
    X"000002FC0A06",         -- len=     764 r=$0A v=$06
    X"000004600805",         -- len=    1120 r=$08 v=$05
    X"0000027F0905",         -- len=     639 r=$09 v=$05
    X"000002FC0A05",         -- len=     764 r=$0A v=$05
    X"0000045F0804",         -- len=    1119 r=$08 v=$04
    X"000002800904",         -- len=     640 r=$09 v=$04
    X"000002FD0A04",         -- len=     765 r=$0A v=$04
    X"0000045E0803",         -- len=    1118 r=$08 v=$03
    X"000002800903",         -- len=     640 r=$09 v=$03
    X"0000027700F0",         -- len=     631 r=$00 v=$F0
    X"000000010100",         -- len=       1 r=$01 v=$00
    X"000000030807",         -- len=       3 r=$08 v=$07
    X"000000820A03",         -- len=     130 r=$0A v=$03
    X"000001F9025D",         -- len=     505 r=$02 v=$5D
    X"000000010302",         -- len=       1 r=$03 v=$02
    X"000000030907",         -- len=       3 r=$09 v=$07
    X"000002610806",         -- len=     609 r=$08 v=$06
    X"000000950A00",         -- len=     149 r=$0A v=$00
    X"000001EB0906",         -- len=     491 r=$09 v=$06
    X"000002FD0A02",         -- len=     765 r=$0A v=$02
    X"0000045E0805",         -- len=    1118 r=$08 v=$05
    X"000002810905",         -- len=     641 r=$09 v=$05
    X"000002FC0A01",         -- len=     764 r=$0A v=$01
    X"0000045F0804",         -- len=    1119 r=$08 v=$04
    X"000002800904",         -- len=     640 r=$09 v=$04
    X"000002FD0A00",         -- len=     765 r=$0A v=$00
    X"0000045E0803",         -- len=    1118 r=$08 v=$03
    X"000002800903",         -- len=     640 r=$09 v=$03
    X"00000277002E",         -- len=     631 r=$00 v=$2E
    X"000000010101",         -- len=       1 r=$01 v=$01
    X"000000030807",         -- len=       3 r=$08 v=$07
    X"0000027C02E0",         -- len=     636 r=$02 v=$E0
    X"000000010301",         -- len=       1 r=$03 v=$01
    X"000000040907",         -- len=       4 r=$09 v=$07
    X"000002610806",         -- len=     609 r=$08 v=$06
    X"00000000045D",         -- len=       0 r=$04 v=$5D
    X"000000000502",         -- len=       0 r=$05 v=$02
    X"0000009A0A07",         -- len=     154 r=$0A v=$07
    X"000001E50906",         -- len=     485 r=$09 v=$06
    X"000002FD0A06",         -- len=     765 r=$0A v=$06
    X"0000045E0805",         -- len=    1118 r=$08 v=$05
    X"0000027E0905",         -- len=     638 r=$09 v=$05
    X"000002FF0A05",         -- len=     767 r=$0A v=$05
    X"0000045E0804",         -- len=    1118 r=$08 v=$04
    X"0000027F0904",         -- len=     639 r=$09 v=$04
    X"000002FC0A04",         -- len=     764 r=$0A v=$04
    X"000004610803",         -- len=    1121 r=$08 v=$03
    X"0000027E0903",         -- len=     638 r=$09 v=$03
    X"000001280738",         -- len=     296 r=$07 v=$38
    X"000000DE04BE",         -- len=     222 r=$04 v=$BE
    X"000000010500",         -- len=       1 r=$05 v=$00
    X"000000050A09",         -- len=       5 r=$0A v=$09
    X"00000000002E",         -- len=       0 r=$00 v=$2E
    X"000000000101",         -- len=       0 r=$01 v=$01
    X"000000EE0807",         -- len=     238 r=$08 v=$07
    X"000000560A08",         -- len=      86 r=$0A v=$08
    X"000002250227",         -- len=     549 r=$02 v=$27
    X"000000010303",         -- len=       1 r=$03 v=$03
    X"000000040907",         -- len=       4 r=$09 v=$07
    X"0000004D0A07",         -- len=      77 r=$0A v=$07
    X"000001370497",         -- len=     311 r=$04 v=$97
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000050A09",         -- len=       5 r=$0A v=$09
    X"000000D70806",         -- len=     215 r=$08 v=$06
    X"000000620A08",         -- len=      98 r=$0A v=$08
    X"0000021E0906",         -- len=     542 r=$09 v=$06
    X"0000005A0A07",         -- len=      90 r=$0A v=$07
    X"00000137047F",         -- len=     311 r=$04 v=$7F
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000050A09",         -- len=       5 r=$0A v=$09
    X"0000013C0A08",         -- len=     316 r=$0A v=$08
    X"000002760A07",         -- len=     630 r=$0A v=$07
    X"00000136045F",         -- len=     310 r=$04 v=$5F
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000050A09",         -- len=       5 r=$0A v=$09
    X"000000D90805",         -- len=     217 r=$08 v=$05
    X"000000620A08",         -- len=      98 r=$0A v=$08
    X"0000021D0905",         -- len=     541 r=$09 v=$05
    X"0000005A0A07",         -- len=      90 r=$0A v=$07
    X"0000013A0471",         -- len=     314 r=$04 v=$71
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000050A09",         -- len=       5 r=$0A v=$09
    X"000001380A08",         -- len=     312 r=$0A v=$08
    X"000002760A07",         -- len=     630 r=$0A v=$07
    X"000002150804",         -- len=     533 r=$08 v=$04
    X"000000630A06",         -- len=      99 r=$0A v=$06
    X"0000021C0904",         -- len=     540 r=$09 v=$04
    X"0000005A0A05",         -- len=      90 r=$0A v=$05
    X"000002770A04",         -- len=     631 r=$0A v=$04
    X"000002760A03",         -- len=     630 r=$0A v=$03
    X"000002140803",         -- len=     532 r=$08 v=$03
    X"000000630A02",         -- len=      99 r=$0A v=$02
    X"0000021D0903",         -- len=     541 r=$09 v=$03
    X"0000005A0A01",         -- len=      90 r=$0A v=$01
    X"000000AE002E",         -- len=     174 r=$00 v=$2E
    X"000000000101",         -- len=       0 r=$01 v=$01
    X"000001730807",         -- len=     371 r=$08 v=$07
    X"000000560A00",         -- len=      86 r=$0A v=$00
    X"0000022502E0",         -- len=     549 r=$02 v=$E0
    X"000000010301",         -- len=       1 r=$03 v=$01
    X"000000040907",         -- len=       4 r=$09 v=$07
    X"000002620806",         -- len=     610 r=$08 v=$06
    X"000002320738",         -- len=     562 r=$07 v=$38
    X"000000980906",         -- len=     152 r=$09 v=$06
    X"0000004604BE",         -- len=      70 r=$04 v=$BE
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000050A09",         -- len=       5 r=$0A v=$09
    X"0000013D0A08",         -- len=     317 r=$0A v=$08
    X"000002780A07",         -- len=     632 r=$0A v=$07
    X"000001390497",         -- len=     313 r=$04 v=$97
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000050A09",         -- len=       5 r=$0A v=$09
    X"000001390A08",         -- len=     313 r=$0A v=$08
    X"000001180805",         -- len=     280 r=$08 v=$05
    X"0000015E0A07",         -- len=     350 r=$0A v=$07
    X"000001200905",         -- len=     288 r=$09 v=$05
    X"0000001D047F",         -- len=      29 r=$04 v=$7F
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000050A09",         -- len=       5 r=$0A v=$09
    X"000001360A08",         -- len=     310 r=$0A v=$08
    X"000002760A07",         -- len=     630 r=$0A v=$07
    X"00000138045F",         -- len=     312 r=$04 v=$5F
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000050A09",         -- len=       5 r=$0A v=$09
    X"000001390A08",         -- len=     313 r=$0A v=$08
    X"000001180804",         -- len=     280 r=$08 v=$04
    X"0000015F0A07",         -- len=     351 r=$0A v=$07
    X"000001220904",         -- len=     290 r=$09 v=$04
    X"0000001E0471",         -- len=      30 r=$04 v=$71
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000060A09",         -- len=       6 r=$0A v=$09
    X"000001310A08",         -- len=     305 r=$0A v=$08
    X"000002780A07",         -- len=     632 r=$0A v=$07
    X"000002760A06",         -- len=     630 r=$0A v=$06
    X"000001170803",         -- len=     279 r=$08 v=$03
    X"0000015F0A05",         -- len=     351 r=$0A v=$05
    X"000001220903",         -- len=     290 r=$09 v=$03
    X"000001560A04",         -- len=     342 r=$0A v=$04
    X"0000012000E3",         -- len=     288 r=$00 v=$E3
    X"000000010100",         -- len=       1 r=$01 v=$00
    X"000000030807",         -- len=       3 r=$08 v=$07
    X"000001530A03",         -- len=     339 r=$0A v=$03
    X"00000128021B",         -- len=     296 r=$02 v=$1B
    X"000000020302",         -- len=       2 r=$03 v=$02
    X"000000030907",         -- len=       3 r=$09 v=$07
    X"0000014A0A02",         -- len=     330 r=$0A v=$02
    X"000001170806",         -- len=     279 r=$08 v=$06
    X"0000015E0A01",         -- len=     350 r=$0A v=$01
    X"000001200906",         -- len=     288 r=$09 v=$06
    X"000001580A00",         -- len=     344 r=$0A v=$00
    X"000006050805",         -- len=    1541 r=$08 v=$05
    X"000002800905",         -- len=     640 r=$09 v=$05
    X"0000075C0804",         -- len=    1884 r=$08 v=$04
    X"0000027E0904",         -- len=     638 r=$09 v=$04
    X"000000000A00",         -- len=       0 r=$0A v=$00
    X"00000058073C",         -- len=      88 r=$07 v=$3C
    X"000000000A00",         -- len=       0 r=$0A v=$00
    X"00000000073C",         -- len=       0 r=$07 v=$3C
    X"000000000A00",         -- len=       0 r=$0A v=$00
    X"000007040803",         -- len=    1796 r=$08 v=$03
    X"000002810903",         -- len=     641 r=$09 v=$03
    X"0000014600E3",         -- len=     326 r=$00 v=$E3
    X"000000000100",         -- len=       0 r=$01 v=$00
    X"000001350807",         -- len=     309 r=$08 v=$07
    X"0000027902C5",         -- len=     633 r=$02 v=$C5
    X"000000010301",         -- len=       1 r=$03 v=$01
    X"000000040907",         -- len=       4 r=$09 v=$07
    X"000002620806",         -- len=     610 r=$08 v=$06
    X"0000027F0906",         -- len=     639 r=$09 v=$06
    X"000000210738",         -- len=      33 r=$07 v=$38
    X"0000006B04BE",         -- len=     107 r=$04 v=$BE
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000050A09",         -- len=       5 r=$0A v=$09
    X"000001430A08",         -- len=     323 r=$0A v=$08
    X"000002780A07",         -- len=     632 r=$0A v=$07
    X"000001360497",         -- len=     310 r=$04 v=$97
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000060A09",         -- len=       6 r=$0A v=$09
    X"0000013B0A08",         -- len=     315 r=$0A v=$08
    X"000000E50805",         -- len=     229 r=$08 v=$05
    X"000001910A07",         -- len=     401 r=$0A v=$07
    X"000000EE0905",         -- len=     238 r=$09 v=$05
    X"00000048047F",         -- len=      72 r=$04 v=$7F
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000060A09",         -- len=       6 r=$0A v=$09
    X"0000013B0A08",         -- len=     315 r=$0A v=$08
    X"000002760A07",         -- len=     630 r=$0A v=$07
    X"00000136045F",         -- len=     310 r=$04 v=$5F
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000060A09",         -- len=       6 r=$0A v=$09
    X"0000013B0A08",         -- len=     315 r=$0A v=$08
    X"000000E50804",         -- len=     229 r=$08 v=$04
    X"000001910A07",         -- len=     401 r=$0A v=$07
    X"000000F00904",         -- len=     240 r=$09 v=$04
    X"0000004B0471",         -- len=      75 r=$04 v=$71
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000050A09",         -- len=       5 r=$0A v=$09
    X"000001370A08",         -- len=     311 r=$0A v=$08
    X"000002780A07",         -- len=     632 r=$0A v=$07
    X"000002760A06",         -- len=     630 r=$0A v=$06
    X"000000E50803",         -- len=     229 r=$08 v=$03
    X"000001910A05",         -- len=     401 r=$0A v=$05
    X"000000F00903",         -- len=     240 r=$09 v=$03
    X"000001880A04",         -- len=     392 r=$0A v=$04
    X"000000EE00F0",         -- len=     238 r=$00 v=$F0
    X"000000000100",         -- len=       0 r=$01 v=$00
    X"000000050807",         -- len=       5 r=$08 v=$07
    X"000001B60A03",         -- len=     438 r=$0A v=$03
    X"000000F70227",         -- len=     247 r=$02 v=$27
    X"000000010303",         -- len=       1 r=$03 v=$03
    X"000000030907",         -- len=       3 r=$09 v=$07
    X"0000017D0A02",         -- len=     381 r=$0A v=$02
    X"000000E50806",         -- len=     229 r=$08 v=$06
    X"000001910A01",         -- len=     401 r=$0A v=$01
    X"000000EE0906",         -- len=     238 r=$09 v=$06
    X"000001880A00",         -- len=     392 r=$0A v=$00
    X"000005D30805",         -- len=    1491 r=$08 v=$05
    X"000000FF0738",         -- len=     255 r=$07 v=$38
    X"000000C404BE",         -- len=     196 r=$04 v=$BE
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000050A09",         -- len=       5 r=$0A v=$09
    X"000001040905",         -- len=     260 r=$09 v=$05
    X"000000410A08",         -- len=      65 r=$0A v=$08
    X"000002760A07",         -- len=     630 r=$0A v=$07
    X"000001500497",         -- len=     336 r=$04 v=$97
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000050A09",         -- len=       5 r=$0A v=$09
    X"0000016E0A08",         -- len=     366 r=$0A v=$08
    X"000002140804",         -- len=     532 r=$08 v=$04
    X"000000620A07",         -- len=      98 r=$0A v=$07
    X"00000136047F",         -- len=     310 r=$04 v=$7F
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000060A09",         -- len=       6 r=$0A v=$09
    X"000000E10904",         -- len=     225 r=$09 v=$04
    X"0000005A0A08",         -- len=      90 r=$0A v=$08
    X"000002760A07",         -- len=     630 r=$0A v=$07
    X"00000139045F",         -- len=     313 r=$04 v=$5F
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000050A09",         -- len=       5 r=$0A v=$09
    X"0000013A0A08",         -- len=     314 r=$0A v=$08
    X"000002150803",         -- len=     533 r=$08 v=$03
    X"000000620A07",         -- len=      98 r=$0A v=$07
    X"000001390471",         -- len=     313 r=$04 v=$71
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000050A09",         -- len=       5 r=$0A v=$09
    X"000000DE0903",         -- len=     222 r=$09 v=$03
    X"0000005A0A08",         -- len=      90 r=$0A v=$08
    X"000000AE00F0",         -- len=     174 r=$00 v=$F0
    X"000000000100",         -- len=       0 r=$01 v=$00
    X"000001740807",         -- len=     372 r=$08 v=$07
    X"000000550A07",         -- len=      85 r=$0A v=$07
    X"0000022602C5",         -- len=     550 r=$02 v=$C5
    X"000000010301",         -- len=       1 r=$03 v=$01
    X"000000040907",         -- len=       4 r=$09 v=$07
    X"0000004B0A06",         -- len=      75 r=$0A v=$06
    X"000002160806",         -- len=     534 r=$08 v=$06
    X"000000630A05",         -- len=      99 r=$0A v=$05
    X"0000021C0906",         -- len=     540 r=$09 v=$06
    X"0000005A0A04",         -- len=      90 r=$0A v=$04
    X"000002300738",         -- len=     560 r=$07 v=$38
    X"000000AA04BE",         -- len=     170 r=$04 v=$BE
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000050A09",         -- len=       5 r=$0A v=$09
    X"000001450A08",         -- len=     325 r=$0A v=$08
    X"000002760A07",         -- len=     630 r=$0A v=$07
    X"000000B40805",         -- len=     180 r=$08 v=$05
    X"0000009C0497",         -- len=     156 r=$04 v=$97
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000060A09",         -- len=       6 r=$0A v=$09
    X"0000016D0A08",         -- len=     365 r=$0A v=$08
    X"000000A20905",         -- len=     162 r=$09 v=$05
    X"000001D40A07",         -- len=     468 r=$0A v=$07
    X"00000137047F",         -- len=     311 r=$04 v=$7F
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000050A09",         -- len=       5 r=$0A v=$09
    X"0000013B0A08",         -- len=     315 r=$0A v=$08
    X"000002770A07",         -- len=     631 r=$0A v=$07
    X"000000990804",         -- len=     153 r=$08 v=$04
    X"0000009D045F",         -- len=     157 r=$04 v=$5F
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000050A09",         -- len=       5 r=$0A v=$09
    X"0000013B0A08",         -- len=     315 r=$0A v=$08
    X"000000A30904",         -- len=     163 r=$09 v=$04
    X"000001D50A07",         -- len=     469 r=$0A v=$07
    X"000001390471",         -- len=     313 r=$04 v=$71
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000060A09",         -- len=       6 r=$0A v=$09
    X"000001370A08",         -- len=     311 r=$0A v=$08
    X"000002780A07",         -- len=     632 r=$0A v=$07
    X"0000009A0803",         -- len=     154 r=$08 v=$03
    X"000001DC0A06",         -- len=     476 r=$0A v=$06
    X"000000A20903",         -- len=     162 r=$09 v=$03
    X"000001D60A05",         -- len=     470 r=$0A v=$05
    X"000000A2000D",         -- len=     162 r=$00 v=$0D
    X"000000010101",         -- len=       1 r=$01 v=$01
    X"000000030807",         -- len=       3 r=$08 v=$07
    X"000001440738",         -- len=     324 r=$07 v=$38
    X"000000BC04BE",         -- len=     188 r=$04 v=$BE
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000050A09",         -- len=       5 r=$0A v=$09
    X"000000C2021B",         -- len=     194 r=$02 v=$1B
    X"000000010302",         -- len=       1 r=$03 v=$02
    X"000000030907",         -- len=       3 r=$09 v=$07
    X"000000B10A08",         -- len=     177 r=$0A v=$08
    X"000001E10806",         -- len=     481 r=$08 v=$06
    X"000000970A07",         -- len=     151 r=$0A v=$07
    X"000001500497",         -- len=     336 r=$04 v=$97
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000050A09",         -- len=       5 r=$0A v=$09
    X"000000E00906",         -- len=     224 r=$09 v=$06
    X"0000008C0A08",         -- len=     140 r=$0A v=$08
    X"000002780A07",         -- len=     632 r=$0A v=$07
    X"00000136047F",         -- len=     310 r=$04 v=$7F
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000050A09",         -- len=       5 r=$0A v=$09
    X"0000013C0A08",         -- len=     316 r=$0A v=$08
    X"000001E20805",         -- len=     482 r=$08 v=$05
    X"000000940A07",         -- len=     148 r=$0A v=$07
    X"00000136045F",         -- len=     310 r=$04 v=$5F
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000050A09",         -- len=       5 r=$0A v=$09
    X"000000B00905",         -- len=     176 r=$09 v=$05
    X"0000008C0A08",         -- len=     140 r=$0A v=$08
    X"000002760A07",         -- len=     630 r=$0A v=$07
    X"0000013B0471",         -- len=     315 r=$04 v=$71
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000050A09",         -- len=       5 r=$0A v=$09
    X"000001380A08",         -- len=     312 r=$0A v=$08
    X"000001E10804",         -- len=     481 r=$08 v=$04
    X"000000940A07",         -- len=     148 r=$0A v=$07
    X"000001EC0904",         -- len=     492 r=$09 v=$04
    X"0000008C0A06",         -- len=     140 r=$0A v=$06
    X"000002760A05",         -- len=     630 r=$0A v=$05
    X"000002780A04",         -- len=     632 r=$0A v=$04
    X"000001E10803",         -- len=     481 r=$08 v=$03
    X"000000240738",         -- len=      36 r=$07 v=$38
    X"000000A104BE",         -- len=     161 r=$04 v=$BE
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000050A09",         -- len=       5 r=$0A v=$09
    X"000001460A08",         -- len=     326 r=$0A v=$08
    X"000000A20903",         -- len=     162 r=$09 v=$03
    X"000001D40A07",         -- len=     468 r=$0A v=$07
    X"000001390497",         -- len=     313 r=$04 v=$97
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000050A09",         -- len=       5 r=$0A v=$09
    X"000001390A08",         -- len=     313 r=$0A v=$08
    X"000000AB02C5",         -- len=     171 r=$02 v=$C5
    X"000000010301",         -- len=       1 r=$03 v=$01
    X"000000030907",         -- len=       3 r=$09 v=$07
    X"000001C80A07",         -- len=     456 r=$0A v=$07
    X"0000009A0802",         -- len=     154 r=$08 v=$02
    X"0000009C047F",         -- len=     156 r=$04 v=$7F
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000060A09",         -- len=       6 r=$0A v=$09
    X"0000013B0A08",         -- len=     315 r=$0A v=$08
    X"000000A30906",         -- len=     163 r=$09 v=$06
    X"000001D30A07",         -- len=     467 r=$0A v=$07
    X"00000139045F",         -- len=     313 r=$04 v=$5F
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000050A09",         -- len=       5 r=$0A v=$09
    X"000001390A08",         -- len=     313 r=$0A v=$08
    X"000002780A07",         -- len=     632 r=$0A v=$07
    X"0000009A0801",         -- len=     154 r=$08 v=$01
    X"0000009F0471",         -- len=     159 r=$04 v=$71
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000050A09",         -- len=       5 r=$0A v=$09
    X"000001380A08",         -- len=     312 r=$0A v=$08
    X"000000A20905",         -- len=     162 r=$09 v=$05
    X"000001D60A07",         -- len=     470 r=$0A v=$07
    X"000002750A06",         -- len=     629 r=$0A v=$06
    X"000002790A05",         -- len=     633 r=$0A v=$05
    X"0000009A0800",         -- len=     154 r=$08 v=$00
    X"000001DC0A04",         -- len=     476 r=$0A v=$04
    X"000000A20904",         -- len=     162 r=$09 v=$04
    X"000001D30A03",         -- len=     467 r=$0A v=$03
    X"000002780A02",         -- len=     632 r=$0A v=$02
    X"000002760A01",         -- len=     630 r=$0A v=$01
    X"000002770A00",         -- len=     631 r=$0A v=$00
    X"000000A20903",         -- len=     162 r=$09 v=$03
    X"000000A90800",         -- len=     169 r=$08 v=$00
    X"0000044E0227",         -- len=    1102 r=$02 v=$27
    X"000000010303",         -- len=       1 r=$03 v=$03
    X"000000030907",         -- len=       3 r=$09 v=$07
    X"000004E10906",         -- len=    1249 r=$09 v=$06
    X"000007DB0A00",         -- len=    2011 r=$0A v=$00
    X"00000060073C",         -- len=      96 r=$07 v=$3C
    X"000000000A00",         -- len=       0 r=$0A v=$00
    X"00000000073C",         -- len=       0 r=$07 v=$3C
    X"000000000A00",         -- len=       0 r=$0A v=$00
    X"000001A00905",         -- len=     416 r=$09 v=$05
    X"000003D90738",         -- len=     985 r=$07 v=$38
    X"000000A304BE",         -- len=     163 r=$04 v=$BE
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000050A09",         -- len=       5 r=$0A v=$09
    X"000001460A08",         -- len=     326 r=$0A v=$08
    X"000002770A07",         -- len=     631 r=$0A v=$07
    X"000001360497",         -- len=     310 r=$04 v=$97
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000060A09",         -- len=       6 r=$0A v=$09
    X"000000DF0904",         -- len=     223 r=$09 v=$04
    X"0000005A0A08",         -- len=      90 r=$0A v=$08
    X"000002780A07",         -- len=     632 r=$0A v=$07
    X"00000136047F",         -- len=     310 r=$04 v=$7F
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000050A09",         -- len=       5 r=$0A v=$09
    X"0000013C0A08",         -- len=     316 r=$0A v=$08
    X"000002770A07",         -- len=     631 r=$0A v=$07
    X"00000136045F",         -- len=     310 r=$04 v=$5F
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000060A09",         -- len=       6 r=$0A v=$09
    X"000000DF0903",         -- len=     223 r=$09 v=$03
    X"0000005A0A08",         -- len=      90 r=$0A v=$08
    X"000002780A07",         -- len=     632 r=$0A v=$07
    X"000001390471",         -- len=     313 r=$04 v=$71
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000050A09",         -- len=       5 r=$0A v=$09
    X"000000E702C5",         -- len=     231 r=$02 v=$C5
    X"000000010301",         -- len=       1 r=$03 v=$01
    X"000000030907",         -- len=       3 r=$09 v=$07
    X"0000004E0A08",         -- len=      78 r=$0A v=$08
    X"000002760A07",         -- len=     630 r=$0A v=$07
    X"0000021C0906",         -- len=     540 r=$09 v=$06
    X"0000005A0A06",         -- len=      90 r=$0A v=$06
    X"000002780A05",         -- len=     632 r=$0A v=$05
    X"000002760A04",         -- len=     630 r=$0A v=$04
    X"000002770A03",         -- len=     631 r=$0A v=$03
    X"000000000738",         -- len=       0 r=$07 v=$38
    X"000000AF04BE",         -- len=     175 r=$04 v=$BE
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000050A09",         -- len=       5 r=$0A v=$09
    X"000001450A08",         -- len=     325 r=$0A v=$08
    X"000000710905",         -- len=     113 r=$09 v=$05
    X"000002050A07",         -- len=     517 r=$0A v=$07
    X"000001360497",         -- len=     310 r=$04 v=$97
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000060A09",         -- len=       6 r=$0A v=$09
    X"0000013B0A08",         -- len=     315 r=$0A v=$08
    X"000002760A07",         -- len=     630 r=$0A v=$07
    X"00000138047F",         -- len=     312 r=$04 v=$7F
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000050A09",         -- len=       5 r=$0A v=$09
    X"0000013C0A08",         -- len=     316 r=$0A v=$08
    X"000000700904",         -- len=     112 r=$09 v=$04
    X"000002050A07",         -- len=     517 r=$0A v=$07
    X"00000137045F",         -- len=     311 r=$04 v=$5F
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000050A09",         -- len=       5 r=$0A v=$09
    X"0000013C0A08",         -- len=     316 r=$0A v=$08
    X"000002760A07",         -- len=     630 r=$0A v=$07
    X"000001390471",         -- len=     313 r=$04 v=$71
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000060A09",         -- len=       6 r=$0A v=$09
    X"000001390A08",         -- len=     313 r=$0A v=$08
    X"0000006E0903",         -- len=     110 r=$09 v=$03
    X"000002080A07",         -- len=     520 r=$0A v=$07
    X"0000007000E3",         -- len=     112 r=$00 v=$E3
    X"000000020100",         -- len=       2 r=$01 v=$00
    X"000000030807",         -- len=       3 r=$08 v=$07
    X"000002350A06",         -- len=     565 r=$0A v=$06
    X"00000079021B",         -- len=     121 r=$02 v=$1B
    X"000000010302",         -- len=       1 r=$03 v=$02
    X"000000030907",         -- len=       3 r=$09 v=$07
    X"000001F90A05",         -- len=     505 r=$0A v=$05
    X"000000680806",         -- len=     104 r=$08 v=$06
    X"0000020E0A04",         -- len=     526 r=$0A v=$04
    X"000000700906",         -- len=     112 r=$09 v=$06
    X"000002080A03",         -- len=     520 r=$0A v=$03
    X"000002770A02",         -- len=     631 r=$0A v=$02
    X"000002770A01",         -- len=     631 r=$0A v=$01
    X"000000660805",         -- len=     102 r=$08 v=$05
    X"000002100A00",         -- len=     528 r=$0A v=$00
    X"000000700905",         -- len=     112 r=$09 v=$05
    X"0000075C0804",         -- len=    1884 r=$08 v=$04
    X"000002800904",         -- len=     640 r=$09 v=$04
    X"0000075A0803",         -- len=    1882 r=$08 v=$03
    X"000000700A00",         -- len=     112 r=$0A v=$00
    X"000000A3073C",         -- len=     163 r=$07 v=$3C
    X"000000000A00",         -- len=       0 r=$0A v=$00
    X"00000000073C",         -- len=       0 r=$07 v=$3C
    X"000000000A00",         -- len=       0 r=$0A v=$00
    X"0000016D0903",         -- len=     365 r=$09 v=$03
    X"000000C700E3",         -- len=     199 r=$00 v=$E3
    X"000000000100",         -- len=       0 r=$01 v=$00
    X"000001B50807",         -- len=     437 r=$08 v=$07
    X"0000027C02C5",         -- len=     636 r=$02 v=$C5
    X"000000010301",         -- len=       1 r=$03 v=$01
    X"000000030907",         -- len=       3 r=$09 v=$07
    X"000002600806",         -- len=     608 r=$08 v=$06
    X"0000027E0906",         -- len=     638 r=$09 v=$06
    X"0000075E0805",         -- len=    1886 r=$08 v=$05
    X"0000027F0905",         -- len=     639 r=$09 v=$05
    X"0000075B0804",         -- len=    1883 r=$08 v=$04
    X"0000027F0904",         -- len=     639 r=$09 v=$04
    X"0000075D0803",         -- len=    1885 r=$08 v=$03
    X"0000027F0903",         -- len=     639 r=$09 v=$03
    X"0000027700F0",         -- len=     631 r=$00 v=$F0
    X"000000000100",         -- len=       0 r=$01 v=$00
    X"000000050807",         -- len=       5 r=$08 v=$07
    X"0000027B0227",         -- len=     635 r=$02 v=$27
    X"000000010303",         -- len=       1 r=$03 v=$03
    X"000000030907",         -- len=       3 r=$09 v=$07
    X"000002600806",         -- len=     608 r=$08 v=$06
    X"0000027F0906",         -- len=     639 r=$09 v=$06
    X"000005C30738",         -- len=    1475 r=$07 v=$38
    X"0000006704BE",         -- len=     103 r=$04 v=$BE
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000050A09",         -- len=       5 r=$0A v=$09
    X"000001450A08",         -- len=     325 r=$0A v=$08
    X"000000340805",         -- len=      52 r=$08 v=$05
    X"000002420A07",         -- len=     578 r=$0A v=$07
    X"0000003E0905",         -- len=      62 r=$09 v=$05
    X"000001120497",         -- len=     274 r=$04 v=$97
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000050A09",         -- len=       5 r=$0A v=$09
    X"0000016E0A08",         -- len=     366 r=$0A v=$08
    X"000002760A07",         -- len=     630 r=$0A v=$07
    X"00000138047F",         -- len=     312 r=$04 v=$7F
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000060A09",         -- len=       6 r=$0A v=$09
    X"000001390A08",         -- len=     313 r=$0A v=$08
    X"0000001C0804",         -- len=      28 r=$08 v=$04
    X"0000025C0A07",         -- len=     604 r=$0A v=$07
    X"000000230904",         -- len=      35 r=$09 v=$04
    X"00000114045F",         -- len=     276 r=$04 v=$5F
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000050A09",         -- len=       5 r=$0A v=$09
    X"0000013A0A08",         -- len=     314 r=$0A v=$08
    X"000002770A07",         -- len=     631 r=$0A v=$07
    X"000001390471",         -- len=     313 r=$04 v=$71
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000050A09",         -- len=       5 r=$0A v=$09
    X"0000013A0A08",         -- len=     314 r=$0A v=$08
    X"0000001A0803",         -- len=      26 r=$08 v=$03
    X"0000025C0A07",         -- len=     604 r=$0A v=$07
    X"000000250903",         -- len=      37 r=$09 v=$03
    X"000002510A06",         -- len=     593 r=$0A v=$06
    X"0000000000F0",         -- len=       0 r=$00 v=$F0
    X"000000000100",         -- len=       0 r=$01 v=$00
    X"000000290807",         -- len=      41 r=$08 v=$07
    X"0000024D0A05",         -- len=     589 r=$0A v=$05
    X"0000002E02C5",         -- len=      46 r=$02 v=$C5
    X"000000010301",         -- len=       1 r=$03 v=$01
    X"000000040907",         -- len=       4 r=$09 v=$07
    X"000002450A04",         -- len=     581 r=$0A v=$04
    X"0000001C0806",         -- len=      28 r=$08 v=$06
    X"0000025C0A03",         -- len=     604 r=$0A v=$03
    X"000000230906",         -- len=      35 r=$09 v=$06
    X"000002520A02",         -- len=     594 r=$0A v=$02
    X"000002760A01",         -- len=     630 r=$0A v=$01
    X"000002790A00",         -- len=     633 r=$0A v=$00
    X"0000001C0805",         -- len=      28 r=$08 v=$05
    X"0000027D0905",         -- len=     637 r=$09 v=$05
    X"0000075C0804",         -- len=    1884 r=$08 v=$04
    X"000002800904",         -- len=     640 r=$09 v=$04
    X"000005900A00",         -- len=    1424 r=$0A v=$00
    X"000000B2073C",         -- len=     178 r=$07 v=$3C
    X"000000000A00",         -- len=       0 r=$0A v=$00
    X"00000000073C",         -- len=       0 r=$07 v=$3C
    X"000000000A00",         -- len=       0 r=$0A v=$00
    X"0000011A0803",         -- len=     282 r=$08 v=$03
    X"0000027F0903",         -- len=     639 r=$09 v=$03
    X"00000277000D",         -- len=     631 r=$00 v=$0D
    X"000000010101",         -- len=       1 r=$01 v=$01
    X"000000030807",         -- len=       3 r=$08 v=$07
    X"0000027C021B",         -- len=     636 r=$02 v=$1B
    X"000000010302",         -- len=       1 r=$03 v=$02
    X"000000030907",         -- len=       3 r=$09 v=$07
    X"000002620806",         -- len=     610 r=$08 v=$06
    X"0000027F0906",         -- len=     639 r=$09 v=$06
    X"0000075B0805",         -- len=    1883 r=$08 v=$05
    X"0000027F0905",         -- len=     639 r=$09 v=$05
    X"0000075E0804",         -- len=    1886 r=$08 v=$04
    X"0000027E0904",         -- len=     638 r=$09 v=$04
    X"0000075C0803",         -- len=    1884 r=$08 v=$03
    X"0000027E0903",         -- len=     638 r=$09 v=$03
    X"000001C4000D",         -- len=     452 r=$00 v=$0D
    X"000000000101",         -- len=       0 r=$01 v=$01
    X"000000B80807",         -- len=     184 r=$08 v=$07
    X"0000027B02C5",         -- len=     635 r=$02 v=$C5
    X"000000010301",         -- len=       1 r=$03 v=$01
    X"000000030907",         -- len=       3 r=$09 v=$07
    X"000002620806",         -- len=     610 r=$08 v=$06
    X"000002800906",         -- len=     640 r=$09 v=$06
    X"0000075B0805",         -- len=    1883 r=$08 v=$05
    X"0000027F0905",         -- len=     639 r=$09 v=$05
    X"0000075D0804",         -- len=    1885 r=$08 v=$04
    X"0000027F0904",         -- len=     639 r=$09 v=$04
    X"0000075B0803",         -- len=    1883 r=$08 v=$03
    X"0000027F0903",         -- len=     639 r=$09 v=$03
    X"0000027900B4",         -- len=     633 r=$00 v=$B4
    X"000000010100",         -- len=       1 r=$01 v=$00
    X"000000030807",         -- len=       3 r=$08 v=$07
    X"0000027A0227",         -- len=     634 r=$02 v=$27
    X"000000010303",         -- len=       1 r=$03 v=$03
    X"000000040907",         -- len=       4 r=$09 v=$07
    X"000002610806",         -- len=     609 r=$08 v=$06
    X"0000027F0906",         -- len=     639 r=$09 v=$06
    X"0000075B0805",         -- len=    1883 r=$08 v=$05
    X"000002810905",         -- len=     641 r=$09 v=$05
    X"000005530738",         -- len=    1363 r=$07 v=$38
    X"000000A304BE",         -- len=     163 r=$04 v=$BE
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000050A09",         -- len=       5 r=$0A v=$09
    X"000001450A08",         -- len=     325 r=$0A v=$08
    X"0000009A0804",         -- len=     154 r=$08 v=$04
    X"000001DC0A07",         -- len=     476 r=$0A v=$07
    X"000000A20904",         -- len=     162 r=$09 v=$04
    X"000000940497",         -- len=     148 r=$04 v=$97
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000060A09",         -- len=       6 r=$0A v=$09
    X"0000013B0A08",         -- len=     315 r=$0A v=$08
    X"000002760A07",         -- len=     630 r=$0A v=$07
    X"00000137047F",         -- len=     311 r=$04 v=$7F
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000050A09",         -- len=       5 r=$0A v=$09
    X"0000013C0A08",         -- len=     316 r=$0A v=$08
    X"000000990803",         -- len=     153 r=$08 v=$03
    X"000001DC0A07",         -- len=     476 r=$0A v=$07
    X"000000A30903",         -- len=     163 r=$09 v=$03
    X"00000096045F",         -- len=     150 r=$04 v=$5F
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000050A09",         -- len=       5 r=$0A v=$09
    X"0000013A0A08",         -- len=     314 r=$0A v=$08
    X"0000002D00B4",         -- len=      45 r=$00 v=$B4
    X"000000000100",         -- len=       0 r=$01 v=$00
    X"0000007A0807",         -- len=     122 r=$08 v=$07
    X"000001D00A07",         -- len=     464 r=$0A v=$07
    X"000000AB02C5",         -- len=     171 r=$02 v=$C5
    X"000000010301",         -- len=       1 r=$03 v=$01
    X"000000030907",         -- len=       3 r=$09 v=$07
    X"0000008A0471",         -- len=     138 r=$04 v=$71
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000060A09",         -- len=       6 r=$0A v=$09
    X"000001370A08",         -- len=     311 r=$0A v=$08
    X"0000009A0806",         -- len=     154 r=$08 v=$06
    X"000001DE0A07",         -- len=     478 r=$0A v=$07
    X"000000A20906",         -- len=     162 r=$09 v=$06
    X"000001D40A06",         -- len=     468 r=$0A v=$06
    X"000002780A05",         -- len=     632 r=$0A v=$05
    X"000002750A04",         -- len=     629 r=$0A v=$04
    X"0000009A0805",         -- len=     154 r=$08 v=$05
    X"000001DD0A03",         -- len=     477 r=$0A v=$03
    X"000000A20905",         -- len=     162 r=$09 v=$05
    X"000001D60A02",         -- len=     470 r=$0A v=$02
    X"000002750A01",         -- len=     629 r=$0A v=$01
    X"000002780A00",         -- len=     632 r=$0A v=$00
    X"0000009A0804",         -- len=     154 r=$08 v=$04
    X"000002800904",         -- len=     640 r=$09 v=$04
    X"0000075C0803",         -- len=    1884 r=$08 v=$03
    X"0000027D0903",         -- len=     637 r=$09 v=$03
    X"0000027700CA",         -- len=     631 r=$00 v=$CA
    X"000000000100",         -- len=       0 r=$01 v=$00
    X"000000050807",         -- len=       5 r=$08 v=$07
    X"0000027C021B",         -- len=     636 r=$02 v=$1B
    X"000000010302",         -- len=       1 r=$03 v=$02
    X"000000030907",         -- len=       3 r=$09 v=$07
    X"0000003D0A00",         -- len=      61 r=$0A v=$00
    X"0000008B073C",         -- len=     139 r=$07 v=$3C
    X"000000000A00",         -- len=       0 r=$0A v=$00
    X"00000000073C",         -- len=       0 r=$07 v=$3C
    X"000000000A00",         -- len=       0 r=$0A v=$00
    X"000001990806",         -- len=     409 r=$08 v=$06
    X"0000027F0906",         -- len=     639 r=$09 v=$06
    X"0000075D0805",         -- len=    1885 r=$08 v=$05
    X"0000027F0905",         -- len=     639 r=$09 v=$05
    X"0000075B0804",         -- len=    1883 r=$08 v=$04
    X"0000027F0904",         -- len=     639 r=$09 v=$04
    X"0000075D0803",         -- len=    1885 r=$08 v=$03
    X"000002800903",         -- len=     640 r=$09 v=$03
    X"0000027600E3",         -- len=     630 r=$00 v=$E3
    X"000000000100",         -- len=       0 r=$01 v=$00
    X"000000040807",         -- len=       4 r=$08 v=$07
    X"0000027C02C5",         -- len=     636 r=$02 v=$C5
    X"000000010301",         -- len=       1 r=$03 v=$01
    X"000000030907",         -- len=       3 r=$09 v=$07
    X"000002610806",         -- len=     609 r=$08 v=$06
    X"0000027E0906",         -- len=     638 r=$09 v=$06
    X"0000075D0805",         -- len=    1885 r=$08 v=$05
    X"0000027F0905",         -- len=     639 r=$09 v=$05
    X"0000075B0804",         -- len=    1883 r=$08 v=$04
    X"000002800904",         -- len=     640 r=$09 v=$04
    X"0000075D0803",         -- len=    1885 r=$08 v=$03
    X"000000290738",         -- len=      41 r=$07 v=$38
    X"0000006904BE",         -- len=     105 r=$04 v=$BE
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000050A09",         -- len=       5 r=$0A v=$09
    X"000001450A08",         -- len=     325 r=$0A v=$08
    X"000000EE0903",         -- len=     238 r=$09 v=$03
    X"0000018A0A07",         -- len=     394 r=$0A v=$07
    X"000000EE00F0",         -- len=     238 r=$00 v=$F0
    X"000000000100",         -- len=       0 r=$01 v=$00
    X"000000040807",         -- len=       4 r=$08 v=$07
    X"0000008F0497",         -- len=     143 r=$04 v=$97
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000050A09",         -- len=       5 r=$0A v=$09
    X"0000016F0A08",         -- len=     367 r=$0A v=$08
    X"000000F60227",         -- len=     246 r=$02 v=$27
    X"000000010303",         -- len=       1 r=$03 v=$03
    X"000000040907",         -- len=       4 r=$09 v=$07
    X"000001AE0A07",         -- len=     430 r=$0A v=$07
    X"000000E60806",         -- len=     230 r=$08 v=$06
    X"0000006B047F",         -- len=     107 r=$04 v=$7F
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000050A09",         -- len=       5 r=$0A v=$09
    X"0000016B0A08",         -- len=     363 r=$0A v=$08
    X"000000EE0906",         -- len=     238 r=$09 v=$06
    X"0000018A0A07",         -- len=     394 r=$0A v=$07
    X"00000137045F",         -- len=     311 r=$04 v=$5F
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000050A09",         -- len=       5 r=$0A v=$09
    X"0000013A0A08",         -- len=     314 r=$0A v=$08
    X"000002780A07",         -- len=     632 r=$0A v=$07
    X"000000E50805",         -- len=     229 r=$08 v=$05
    X"000000530471",         -- len=      83 r=$04 v=$71
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000060A09",         -- len=       6 r=$0A v=$09
    X"000001390A08",         -- len=     313 r=$0A v=$08
    X"000000ED0905",         -- len=     237 r=$09 v=$05
    X"000001890A07",         -- len=     393 r=$0A v=$07
    X"000002760A06",         -- len=     630 r=$0A v=$06
    X"000000DD0738",         -- len=     221 r=$07 v=$38
    X"000000D004BE",         -- len=     208 r=$04 v=$BE
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000050A09",         -- len=       5 r=$0A v=$09
    X"000001430A08",         -- len=     323 r=$0A v=$08
    X"000000E70804",         -- len=     231 r=$08 v=$04
    X"000001910A07",         -- len=     401 r=$0A v=$07
    X"000000EE0904",         -- len=     238 r=$09 v=$04
    X"000000480497",         -- len=      72 r=$04 v=$97
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000060A09",         -- len=       6 r=$0A v=$09
    X"0000013B0A08",         -- len=     315 r=$0A v=$08
    X"000002750A07",         -- len=     629 r=$0A v=$07
    X"00000137047F",         -- len=     311 r=$04 v=$7F
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000050A09",         -- len=       5 r=$0A v=$09
    X"0000013C0A08",         -- len=     316 r=$0A v=$08
    X"000000E50803",         -- len=     229 r=$08 v=$03
    X"000001910A07",         -- len=     401 r=$0A v=$07
    X"000000EE0903",         -- len=     238 r=$09 v=$03
    X"00000048045F",         -- len=      72 r=$04 v=$5F
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000060A09",         -- len=       6 r=$0A v=$09
    X"0000013B0A08",         -- len=     315 r=$0A v=$08
    X"000000EE000D",         -- len=     238 r=$00 v=$0D
    X"000000010101",         -- len=       1 r=$01 v=$01
    X"000000030807",         -- len=       3 r=$08 v=$07
    X"000001B70A07",         -- len=     439 r=$0A v=$07
    X"000000F702C5",         -- len=     247 r=$02 v=$C5
    X"000000010301",         -- len=       1 r=$03 v=$01
    X"000000040907",         -- len=       4 r=$09 v=$07
    X"000000580471",         -- len=      88 r=$04 v=$71
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000050A09",         -- len=       5 r=$0A v=$09
    X"0000016A0A08",         -- len=     362 r=$0A v=$08
    X"000000E50806",         -- len=     229 r=$08 v=$06
    X"000001910A07",         -- len=     401 r=$0A v=$07
    X"000000EF0906",         -- len=     239 r=$09 v=$06
    X"000001890A06",         -- len=     393 r=$0A v=$06
    X"000002760A05",         -- len=     630 r=$0A v=$05
    X"000002780A04",         -- len=     632 r=$0A v=$04
    X"000000E50805",         -- len=     229 r=$08 v=$05
    X"000001900A03",         -- len=     400 r=$0A v=$03
    X"000000EE0905",         -- len=     238 r=$09 v=$05
    X"0000018B0A02",         -- len=     395 r=$0A v=$02
    X"000002760A01",         -- len=     630 r=$0A v=$01
    X"000002750A00",         -- len=     629 r=$0A v=$00
    X"000000E80804",         -- len=     232 r=$08 v=$04
    X"0000027D0904",         -- len=     637 r=$09 v=$04
    X"0000075C0803",         -- len=    1884 r=$08 v=$03
    X"000002800903",         -- len=     640 r=$09 v=$03
    X"00000278002E",         -- len=     632 r=$00 v=$2E
    X"000000000101",         -- len=       0 r=$01 v=$01
    X"000000040807",         -- len=       4 r=$08 v=$07
    X"000002AD02E0",         -- len=     685 r=$02 v=$E0
    X"000000000301",         -- len=       0 r=$03 v=$01
    X"000000050907",         -- len=       5 r=$09 v=$07
    X"000000000A00",         -- len=       0 r=$0A v=$00
    X"0000007C073C",         -- len=     124 r=$07 v=$3C
    X"000000000A00",         -- len=       0 r=$0A v=$00
    X"00000000073C",         -- len=       0 r=$07 v=$3C
    X"000000000A00",         -- len=       0 r=$0A v=$00
    X"000001E60806",         -- len=     486 r=$08 v=$06
    X"0000027E0906",         -- len=     638 r=$09 v=$06
    X"0000075B0805",         -- len=    1883 r=$08 v=$05
    X"0000027F0905",         -- len=     639 r=$09 v=$05
    X"0000075D0804",         -- len=    1885 r=$08 v=$04
    X"000002800904",         -- len=     640 r=$09 v=$04
    X"0000075B0803",         -- len=    1883 r=$08 v=$03
    X"0000027F0903",         -- len=     639 r=$09 v=$03
    X"0000075D0802",         -- len=    1885 r=$08 v=$02
    X"0000027F0902",         -- len=     639 r=$09 v=$02
    X"0000075B0801",         -- len=    1883 r=$08 v=$01
    X"0000027F0901",         -- len=     639 r=$09 v=$01
    X"0000075D0800",         -- len=    1885 r=$08 v=$00
    X"0000027F0900",         -- len=     639 r=$09 v=$00
    X"00000BFB0800",         -- len=    3067 r=$08 v=$00
    X"000000000900",         -- len=       0 r=$09 v=$00
    X"00000B940738",         -- len=    2964 r=$07 v=$38
    X"000000A304BE",         -- len=     163 r=$04 v=$BE
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000060A09",         -- len=       6 r=$0A v=$09
    X"000001430A08",         -- len=     323 r=$0A v=$08
    X"000002770A07",         -- len=     631 r=$0A v=$07
    X"000001390497",         -- len=     313 r=$04 v=$97
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000050A09",         -- len=       5 r=$0A v=$09
    X"0000013A0A08",         -- len=     314 r=$0A v=$08
    X"000002760A07",         -- len=     630 r=$0A v=$07
    X"00000136047F",         -- len=     310 r=$04 v=$7F
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000060A09",         -- len=       6 r=$0A v=$09
    X"000000B4073F",         -- len=     180 r=$07 v=$3F
    X"00000009073C",         -- len=       9 r=$07 v=$3C
    X"000000030A00",         -- len=       3 r=$0A v=$00
    X"00000014073D",         -- len=      20 r=$07 v=$3D
    X"000000000800",         -- len=       0 r=$08 v=$00
    X"00000013073F",         -- len=      19 r=$07 v=$3F
    X"000000000900",         -- len=       0 r=$09 v=$00
    X"000002B0080D",         -- len=     688 r=$08 v=$0D
    X"000000030050",         -- len=       3 r=$00 v=$50
    X"000000010100",         -- len=       1 r=$01 v=$00
    X"00000004073E",         -- len=       4 r=$07 v=$3E
    X"00000031005A",         -- len=      49 r=$00 v=$5A
    X"000000000100",         -- len=       0 r=$01 v=$00
    X"0000004A0050",         -- len=      74 r=$00 v=$50
    X"000000000100",         -- len=       0 r=$01 v=$00
    X"00000033005A",         -- len=      51 r=$00 v=$5A
    X"000000000100",         -- len=       0 r=$01 v=$00
    X"0000004D0050",         -- len=      77 r=$00 v=$50
    X"000000000100",         -- len=       0 r=$01 v=$00
    X"00000031005A",         -- len=      49 r=$00 v=$5A
    X"000000000100",         -- len=       0 r=$01 v=$00
    X"0000004C0050",         -- len=      76 r=$00 v=$50
    X"000000000100",         -- len=       0 r=$01 v=$00
    X"00000031005A",         -- len=      49 r=$00 v=$5A
    X"000000000100",         -- len=       0 r=$01 v=$00
    X"0000004D0050",         -- len=      77 r=$00 v=$50
    X"000000000100",         -- len=       0 r=$01 v=$00
    X"00000033005A",         -- len=      51 r=$00 v=$5A
    X"000000000100",         -- len=       0 r=$01 v=$00
    X"000000060800",         -- len=       6 r=$08 v=$00
    X"000000CD073C",         -- len=     205 r=$07 v=$3C
    X"000000A50287",         -- len=     165 r=$02 v=$87
    X"000000010300",         -- len=       1 r=$03 v=$00
    X"000000030906",         -- len=       3 r=$09 v=$06
    X"000002190738",         -- len=     537 r=$07 v=$38
    X"0000005804A0",         -- len=      88 r=$04 v=$A0
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000040A06",         -- len=       4 r=$0A v=$06
    X"000001CE0905",         -- len=     462 r=$09 v=$05
    X"000002320A05",         -- len=     562 r=$0A v=$05
    X"000001B3080D",         -- len=     435 r=$08 v=$0D
    X"000000370050",         -- len=      55 r=$00 v=$50
    X"000000000100",         -- len=       0 r=$01 v=$00
    X"0000004A005A",         -- len=      74 r=$00 v=$5A
    X"000000000100",         -- len=       0 r=$01 v=$00
    X"000000330050",         -- len=      51 r=$00 v=$50
    X"000000000100",         -- len=       0 r=$01 v=$00
    X"0000004C005A",         -- len=      76 r=$00 v=$5A
    X"000000000100",         -- len=       0 r=$01 v=$00
    X"000000330050",         -- len=      51 r=$00 v=$50
    X"000000000100",         -- len=       0 r=$01 v=$00
    X"0000004C005A",         -- len=      76 r=$00 v=$5A
    X"000000000100",         -- len=       0 r=$01 v=$00
    X"000000330050",         -- len=      51 r=$00 v=$50
    X"000000000100",         -- len=       0 r=$01 v=$00
    X"0000004B005A",         -- len=      75 r=$00 v=$5A
    X"000000000100",         -- len=       0 r=$01 v=$00
    X"000000330050",         -- len=      51 r=$00 v=$50
    X"000000000100",         -- len=       0 r=$01 v=$00
    X"000000060800",         -- len=       6 r=$08 v=$00
    X"000001C70904",         -- len=     455 r=$09 v=$04
    X"000002320A04",         -- len=     562 r=$0A v=$04
    X"00000266080D",         -- len=     614 r=$08 v=$0D
    X"000000000050",         -- len=       0 r=$00 v=$50
    X"000000000100",         -- len=       0 r=$01 v=$00
    X"000000000738",         -- len=       0 r=$07 v=$38
    X"0000000E0800",         -- len=      14 r=$08 v=$00
    X"00000040005A",         -- len=      64 r=$00 v=$5A
    X"000000000100",         -- len=       0 r=$01 v=$00
    X"000000330050",         -- len=      51 r=$00 v=$50
    X"000000000100",         -- len=       0 r=$01 v=$00
    X"0000004C005A",         -- len=      76 r=$00 v=$5A
    X"000000000100",         -- len=       0 r=$01 v=$00
    X"000000330050",         -- len=      51 r=$00 v=$50
    X"000000000100",         -- len=       0 r=$01 v=$00
    X"0000004A005A",         -- len=      74 r=$00 v=$5A
    X"000000000100",         -- len=       0 r=$01 v=$00
    X"000000320050",         -- len=      50 r=$00 v=$50
    X"000000000100",         -- len=       0 r=$01 v=$00
    X"0000004C005A",         -- len=      76 r=$00 v=$5A
    X"000000000100",         -- len=       0 r=$01 v=$00
    X"000000330050",         -- len=      51 r=$00 v=$50
    X"000000000100",         -- len=       0 r=$01 v=$00
    X"0000004C005A",         -- len=      76 r=$00 v=$5A
    X"000000000100",         -- len=       0 r=$01 v=$00
    X"000000000800",         -- len=       0 r=$08 v=$00
    X"000001030903",         -- len=     259 r=$09 v=$03
    X"000002320A03",         -- len=     562 r=$0A v=$03
    X"000005A7080D",         -- len=    1447 r=$08 v=$0D
    X"0000000F0902",         -- len=      15 r=$09 v=$02
    X"000000260050",         -- len=      38 r=$00 v=$50
    X"000000000100",         -- len=       0 r=$01 v=$00
    X"0000004C005A",         -- len=      76 r=$00 v=$5A
    X"000000000100",         -- len=       0 r=$01 v=$00
    X"000000320050",         -- len=      50 r=$00 v=$50
    X"000000000100",         -- len=       0 r=$01 v=$00
    X"0000004C005A",         -- len=      76 r=$00 v=$5A
    X"000000000100",         -- len=       0 r=$01 v=$00
    X"000000330050",         -- len=      51 r=$00 v=$50
    X"000000000100",         -- len=       0 r=$01 v=$00
    X"0000004C005A",         -- len=      76 r=$00 v=$5A
    X"000000000100",         -- len=       0 r=$01 v=$00
    X"000000320050",         -- len=      50 r=$00 v=$50
    X"000000000100",         -- len=       0 r=$01 v=$00
    X"0000004A005A",         -- len=      74 r=$00 v=$5A
    X"000000000100",         -- len=       0 r=$01 v=$00
    X"000000330050",         -- len=      51 r=$00 v=$50
    X"000000000100",         -- len=       0 r=$01 v=$00
    X"000000060800",         -- len=       6 r=$08 v=$00
    X"000000170A02",         -- len=      23 r=$0A v=$02
    X"000001B50900",         -- len=     437 r=$09 v=$00
    X"000002350A00",         -- len=     565 r=$0A v=$00
    X"000001B80901",         -- len=     440 r=$09 v=$01
    X"0000002F0800",         -- len=      47 r=$08 v=$00
    X"0000007B0739",         -- len=     123 r=$07 v=$39
    X"000000000800",         -- len=       0 r=$08 v=$00
    X"000000000739",         -- len=       0 r=$07 v=$39
    X"000000000800",         -- len=       0 r=$08 v=$00
    X"000001840A01",         -- len=     388 r=$0A v=$01
    X"000005AF0900",         -- len=    1455 r=$09 v=$00
    X"000002340A00",         -- len=     564 r=$0A v=$00
    X"000001C60278",         -- len=     454 r=$02 v=$78
    X"000000000300",         -- len=       0 r=$03 v=$00
    X"000000040906",         -- len=       4 r=$09 v=$06
    X"0000023004AA",         -- len=     560 r=$04 v=$AA
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000040A06",         -- len=       4 r=$0A v=$06
    X"000001B10905",         -- len=     433 r=$09 v=$05
    X"000002340A05",         -- len=     564 r=$0A v=$05
    X"000005AE0904",         -- len=    1454 r=$09 v=$04
    X"000002340A04",         -- len=     564 r=$0A v=$04
    X"000001C80287",         -- len=     456 r=$02 v=$87
    X"000000000300",         -- len=       0 r=$03 v=$00
    X"000000040906",         -- len=       4 r=$09 v=$06
    X"0000022F04A0",         -- len=     559 r=$04 v=$A0
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000040A06",         -- len=       4 r=$0A v=$06
    X"000001B10905",         -- len=     433 r=$09 v=$05
    X"000002310A05",         -- len=     561 r=$0A v=$05
    X"000005B10904",         -- len=    1457 r=$09 v=$04
    X"000002330A04",         -- len=     563 r=$0A v=$04
    X"000005AF0903",         -- len=    1455 r=$09 v=$03
    X"000002340A03",         -- len=     564 r=$0A v=$03
    X"000005AF0902",         -- len=    1455 r=$09 v=$02
    X"000002330A02",         -- len=     563 r=$0A v=$02
    X"000005AF0901",         -- len=    1455 r=$09 v=$01
    X"000002340A01",         -- len=     564 r=$0A v=$01
    X"000005AE0900",         -- len=    1454 r=$09 v=$00
    X"000002340A00",         -- len=     564 r=$0A v=$00
    X"0000118C02C5",         -- len=    4492 r=$02 v=$C5
    X"000000010301",         -- len=       1 r=$03 v=$01
    X"000000030906",         -- len=       3 r=$09 v=$06
    X"0000022F04CA",         -- len=     559 r=$04 v=$CA
    X"000000000500",         -- len=       0 r=$05 v=$00
    X"000000040A06",         -- len=       4 r=$0A v=$06
    X"000001B10905",         -- len=     433 r=$09 v=$05
    X"000002340A05",         -- len=     564 r=$0A v=$05
    X"000005AE0904",         -- len=    1454 r=$09 v=$04
    X"000002340A04",         -- len=     564 r=$0A v=$04
    X"000005AE0903",         -- len=    1454 r=$09 v=$03
    X"000002340A03",         -- len=     564 r=$0A v=$03
    X"000005AF0902",         -- len=    1455 r=$09 v=$02
    X"000002330A02"          -- len=     563 r=$0A v=$02
);
signal raddr : std_logic_vector(10 downto 0);
begin
  process (clk)
    begin
      if (clk'event and clk = '1') then
          if (en = '1') then
              raddr <= addr;
          end if;
      end if;
  end process;
  data <= ROM(conv_integer(raddr));
end syn;
