library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity snd_rom is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of snd_rom is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"F3",X"ED",X"56",X"31",X"00",X"88",X"C3",X"7E",X"00",X"9D",X"1B",X"AA",X"1B",X"B7",X"1B",X"C4",
		X"1B",X"D1",X"1B",X"DE",X"1B",X"EB",X"1B",X"80",X"20",X"00",X"00",X"00",X"01",X"00",X"F8",X"1B",
		X"00",X"20",X"00",X"00",X"80",X"21",X"00",X"00",X"00",X"01",X"00",X"F0",X"1C",X"00",X"20",X"00",
		X"00",X"00",X"22",X"00",X"00",X"00",X"01",X"00",X"F5",X"E5",X"21",X"00",X"80",X"35",X"E1",X"F1",
		X"FB",X"C9",X"00",X"01",X"00",X"42",X"1E",X"00",X"20",X"00",X"00",X"00",X"10",X"00",X"00",X"00",
		X"01",X"00",X"E8",X"1D",X"00",X"20",X"00",X"00",X"80",X"11",X"00",X"00",X"00",X"01",X"00",X"17",
		X"1E",X"00",X"20",X"00",X"00",X"80",X"F3",X"F5",X"3A",X"00",X"E0",X"FE",X"90",X"C2",X"77",X"00",
		X"08",X"3E",X"01",X"32",X"02",X"81",X"08",X"32",X"00",X"81",X"F1",X"FB",X"ED",X"45",X"CD",X"66",
		X"04",X"21",X"00",X"80",X"11",X"01",X"80",X"01",X"FF",X"07",X"36",X"00",X"ED",X"B0",X"FB",X"CD",
		X"8B",X"04",X"21",X"00",X"80",X"7E",X"B7",X"28",X"F6",X"36",X"00",X"DD",X"21",X"00",X"82",X"06",
		X"14",X"C5",X"DD",X"CB",X"00",X"7E",X"C4",X"B4",X"00",X"11",X"20",X"00",X"DD",X"19",X"C1",X"10",
		X"F0",X"C3",X"8F",X"00",X"DD",X"CB",X"00",X"66",X"C2",X"E0",X"03",X"DD",X"5E",X"03",X"DD",X"56",
		X"04",X"13",X"DD",X"73",X"03",X"DD",X"72",X"04",X"DD",X"6E",X"05",X"DD",X"66",X"06",X"B7",X"ED",
		X"52",X"CC",X"41",X"02",X"DD",X"CB",X"03",X"46",X"C0",X"DD",X"5E",X"11",X"DD",X"56",X"12",X"7B",
		X"B2",X"20",X"07",X"DD",X"36",X"17",X"0F",X"C3",X"B6",X"01",X"DD",X"CB",X"00",X"6E",X"20",X"33",
		X"DD",X"7E",X"0B",X"B7",X"20",X"08",X"DD",X"73",X"13",X"DD",X"72",X"14",X"18",X"59",X"3D",X"21",
		X"DD",X"06",X"23",X"DD",X"4E",X"0E",X"06",X"00",X"09",X"09",X"4E",X"23",X"66",X"69",X"0E",X"04",
		X"09",X"4E",X"23",X"66",X"69",X"4F",X"06",X"00",X"09",X"09",X"7E",X"23",X"66",X"6F",X"CD",X"0E",
		X"02",X"18",X"34",X"D5",X"DD",X"6E",X"15",X"DD",X"66",X"16",X"B7",X"ED",X"52",X"F5",X"7D",X"F2",
		X"34",X"01",X"ED",X"44",X"67",X"DD",X"5E",X"03",X"CD",X"96",X"06",X"DD",X"5E",X"05",X"CD",X"A2",
		X"06",X"5F",X"16",X"00",X"F1",X"7B",X"F2",X"4F",X"01",X"ED",X"44",X"28",X"02",X"15",X"5F",X"E1",
		X"19",X"DD",X"75",X"13",X"DD",X"74",X"14",X"DD",X"7E",X"0C",X"B7",X"20",X"0B",X"DD",X"7E",X"0D",
		X"2F",X"E6",X"0F",X"DD",X"77",X"17",X"18",X"23",X"3D",X"21",X"DD",X"06",X"23",X"DD",X"4E",X"0E",
		X"06",X"00",X"09",X"09",X"4E",X"23",X"66",X"69",X"0E",X"02",X"09",X"4E",X"23",X"66",X"69",X"4F",
		X"06",X"00",X"09",X"09",X"7E",X"23",X"66",X"6F",X"CD",X"D4",X"01",X"DD",X"CB",X"00",X"76",X"20",
		X"25",X"DD",X"7E",X"01",X"E6",X"0F",X"4F",X"06",X"00",X"21",X"C9",X"01",X"09",X"4E",X"DD",X"7E",
		X"13",X"E6",X"0F",X"B1",X"CD",X"00",X"04",X"DD",X"7E",X"13",X"E6",X"F0",X"DD",X"B6",X"14",X"0F",
		X"0F",X"0F",X"0F",X"CD",X"00",X"04",X"DD",X"7E",X"01",X"E6",X"0F",X"4F",X"06",X"00",X"21",X"CD",
		X"01",X"09",X"7E",X"DD",X"B6",X"17",X"C3",X"00",X"04",X"80",X"A0",X"C0",X"C0",X"90",X"B0",X"D0",
		X"F0",X"DD",X"77",X"0F",X"E5",X"DD",X"7E",X"0F",X"CB",X"3F",X"F5",X"4F",X"06",X"00",X"09",X"F1",
		X"7E",X"E1",X"38",X"14",X"0F",X"0F",X"0F",X"0F",X"B7",X"28",X"E6",X"FE",X"10",X"20",X"05",X"DD",
		X"35",X"0F",X"18",X"E0",X"FE",X"20",X"28",X"0B",X"DD",X"34",X"0F",X"F6",X"F0",X"DD",X"86",X"0D",
		X"3C",X"38",X"01",X"AF",X"2F",X"E6",X"0F",X"DD",X"77",X"17",X"C9",X"DD",X"77",X"10",X"E5",X"DD",
		X"7E",X"10",X"CB",X"3F",X"F5",X"4F",X"06",X"00",X"09",X"F1",X"7E",X"E1",X"38",X"11",X"0F",X"0F",
		X"0F",X"0F",X"B7",X"CA",X"0B",X"02",X"FE",X"10",X"20",X"05",X"DD",X"35",X"10",X"18",X"DF",X"DD",
		X"34",X"10",X"2F",X"E6",X"0F",X"6F",X"26",X"00",X"EB",X"19",X"DD",X"75",X"13",X"DD",X"74",X"14",
		X"C9",X"DD",X"5E",X"07",X"DD",X"56",X"08",X"1A",X"13",X"B7",X"FA",X"C6",X"02",X"DD",X"CB",X"00",
		X"5E",X"20",X"59",X"B7",X"28",X"03",X"DD",X"86",X"09",X"21",X"1C",X"06",X"4F",X"06",X"00",X"09",
		X"09",X"7E",X"DD",X"77",X"11",X"23",X"7E",X"DD",X"77",X"12",X"DD",X"CB",X"00",X"6E",X"28",X"16",
		X"1A",X"13",X"DD",X"86",X"09",X"21",X"1C",X"06",X"4F",X"06",X"00",X"09",X"09",X"7E",X"DD",X"77",
		X"15",X"23",X"7E",X"DD",X"77",X"16",X"D5",X"1A",X"67",X"DD",X"5E",X"02",X"CD",X"96",X"06",X"D1",
		X"DD",X"75",X"05",X"DD",X"74",X"06",X"AF",X"DD",X"77",X"0F",X"DD",X"77",X"10",X"13",X"DD",X"73",
		X"07",X"DD",X"72",X"08",X"AF",X"DD",X"77",X"03",X"DD",X"77",X"04",X"C9",X"DD",X"77",X"12",X"1A",
		X"13",X"DD",X"77",X"11",X"DD",X"CB",X"00",X"6E",X"28",X"CC",X"1A",X"13",X"DD",X"77",X"16",X"1A",
		X"13",X"DD",X"77",X"15",X"18",X"C0",X"21",X"D9",X"02",X"E5",X"E6",X"3F",X"21",X"DD",X"02",X"4F",
		X"06",X"00",X"09",X"09",X"7E",X"23",X"66",X"6F",X"E9",X"13",X"C3",X"47",X"02",X"AA",X"03",X"03",
		X"03",X"08",X"03",X"1D",X"03",X"CF",X"03",X"31",X"03",X"48",X"03",X"4D",X"03",X"58",X"03",X"73",
		X"03",X"52",X"03",X"86",X"03",X"8E",X"03",X"A6",X"03",X"AC",X"03",X"B2",X"03",X"B8",X"03",X"BE",
		X"03",X"C6",X"03",X"1A",X"DD",X"77",X"02",X"C9",X"1A",X"DD",X"77",X"0D",X"C9",X"0F",X"0E",X"0D",
		X"0C",X"0B",X"0A",X"09",X"07",X"08",X"06",X"05",X"04",X"03",X"02",X"01",X"00",X"1A",X"D5",X"5F",
		X"DD",X"66",X"02",X"CD",X"96",X"06",X"DD",X"75",X"03",X"DD",X"74",X"04",X"D1",X"E1",X"C3",X"9D",
		X"02",X"1A",X"F6",X"E0",X"F5",X"CD",X"00",X"04",X"F1",X"F6",X"FC",X"3C",X"20",X"05",X"DD",X"CB",
		X"00",X"B6",X"C9",X"DD",X"CB",X"00",X"F6",X"C9",X"1A",X"DD",X"77",X"0C",X"C9",X"1A",X"DD",X"77",
		X"0B",X"C9",X"EB",X"5E",X"23",X"56",X"1B",X"C9",X"1A",X"4F",X"13",X"1A",X"47",X"C5",X"DD",X"E5",
		X"E1",X"DD",X"35",X"0A",X"DD",X"4E",X"0A",X"DD",X"35",X"0A",X"06",X"00",X"09",X"72",X"2B",X"73",
		X"D1",X"1B",X"C9",X"DD",X"E5",X"E1",X"DD",X"4E",X"0A",X"06",X"00",X"09",X"5E",X"23",X"56",X"DD",
		X"34",X"0A",X"DD",X"34",X"0A",X"C9",X"1A",X"DD",X"86",X"09",X"DD",X"77",X"09",X"C9",X"1A",X"13",
		X"C6",X"18",X"4F",X"06",X"00",X"DD",X"E5",X"E1",X"09",X"7E",X"B7",X"20",X"02",X"1A",X"77",X"13",
		X"35",X"C2",X"52",X"03",X"13",X"C9",X"DD",X"CB",X"00",X"EE",X"1B",X"C9",X"DD",X"CB",X"00",X"AE",
		X"1B",X"C9",X"DD",X"CB",X"00",X"DE",X"1B",X"C9",X"DD",X"CB",X"00",X"9E",X"1B",X"C9",X"1A",X"DD",
		X"B6",X"00",X"DD",X"77",X"00",X"C9",X"1A",X"2F",X"DD",X"A6",X"00",X"DD",X"77",X"00",X"C9",X"CD",
		X"F1",X"03",X"DD",X"36",X"00",X"00",X"E1",X"E1",X"CD",X"C9",X"06",X"AF",X"32",X"02",X"81",X"C9",
		X"DD",X"35",X"04",X"C0",X"DD",X"7E",X"03",X"DD",X"77",X"04",X"DD",X"6E",X"05",X"DD",X"66",X"06",
		X"E9",X"DD",X"7E",X"01",X"E6",X"0F",X"4F",X"06",X"00",X"21",X"CD",X"01",X"09",X"7E",X"F6",X"0F",
		X"DD",X"CB",X"00",X"56",X"C0",X"ED",X"47",X"DD",X"7E",X"01",X"E6",X"F0",X"FE",X"30",X"28",X"10",
		X"FE",X"10",X"28",X"06",X"ED",X"57",X"32",X"00",X"A0",X"C9",X"ED",X"57",X"32",X"00",X"C0",X"C9",
		X"ED",X"57",X"C9",X"C5",X"E5",X"ED",X"47",X"E6",X"03",X"06",X"00",X"4F",X"21",X"87",X"04",X"09",
		X"4E",X"ED",X"57",X"E6",X"30",X"FE",X"30",X"28",X"0F",X"CB",X"67",X"79",X"20",X"05",X"32",X"00",
		X"C0",X"18",X"06",X"32",X"00",X"A0",X"18",X"01",X"79",X"E1",X"C1",X"C9",X"21",X"00",X"82",X"11",
		X"01",X"82",X"01",X"7F",X"02",X"36",X"00",X"ED",X"B0",X"21",X"00",X"82",X"11",X"01",X"82",X"01",
		X"A0",X"01",X"36",X"00",X"ED",X"B0",X"21",X"87",X"04",X"11",X"00",X"A0",X"01",X"04",X"00",X"ED",
		X"B0",X"21",X"87",X"04",X"11",X"00",X"C0",X"01",X"04",X"00",X"ED",X"B0",X"C9",X"21",X"00",X"80",
		X"7E",X"B7",X"28",X"FC",X"36",X"00",X"C9",X"9F",X"BF",X"DF",X"FF",X"3A",X"00",X"81",X"CB",X"7F",
		X"CA",X"4C",X"04",X"FE",X"00",X"CA",X"4C",X"04",X"FE",X"FF",X"CA",X"4C",X"04",X"21",X"BF",X"04",
		X"01",X"10",X"00",X"ED",X"B9",X"C0",X"21",X"BF",X"04",X"09",X"09",X"7E",X"23",X"66",X"6F",X"E9",
		X"82",X"84",X"85",X"86",X"88",X"89",X"8A",X"8B",X"8C",X"8D",X"8E",X"90",X"93",X"94",X"95",X"DD",
		X"04",X"EB",X"04",X"FA",X"04",X"09",X"05",X"2D",X"05",X"3C",X"05",X"4B",X"05",X"5A",X"05",X"76",
		X"05",X"8A",X"05",X"9E",X"05",X"AD",X"05",X"BC",X"05",X"CB",X"05",X"DA",X"05",X"CD",X"4C",X"04",
		X"21",X"00",X"10",X"11",X"00",X"82",X"AF",X"08",X"C3",X"E9",X"05",X"CD",X"4C",X"04",X"21",X"7C",
		X"10",X"11",X"00",X"82",X"3E",X"01",X"08",X"C3",X"E9",X"05",X"CD",X"4C",X"04",X"21",X"A4",X"11",
		X"11",X"00",X"82",X"3E",X"02",X"08",X"C3",X"E9",X"05",X"3A",X"02",X"81",X"CB",X"47",X"C2",X"0E",
		X"06",X"21",X"01",X"81",X"36",X"FF",X"CD",X"B5",X"06",X"CD",X"66",X"04",X"21",X"02",X"81",X"CB",
		X"CE",X"21",X"CC",X"12",X"11",X"00",X"83",X"3E",X"03",X"08",X"C3",X"E9",X"05",X"CD",X"4C",X"04",
		X"21",X"3F",X"13",X"11",X"00",X"82",X"3E",X"04",X"08",X"C3",X"E9",X"05",X"CD",X"59",X"04",X"21",
		X"4D",X"14",X"11",X"00",X"82",X"3E",X"05",X"08",X"C3",X"E9",X"05",X"CD",X"59",X"04",X"21",X"CF",
		X"15",X"11",X"00",X"82",X"3E",X"06",X"08",X"C3",X"E9",X"05",X"3A",X"02",X"81",X"CB",X"47",X"C2",
		X"0E",X"06",X"3A",X"02",X"81",X"CB",X"4F",X"C2",X"0E",X"06",X"21",X"81",X"17",X"11",X"E0",X"82",
		X"3E",X"07",X"08",X"C3",X"E9",X"05",X"3A",X"02",X"81",X"CB",X"47",X"C2",X"0E",X"06",X"21",X"CE",
		X"17",X"11",X"80",X"82",X"3E",X"08",X"08",X"C3",X"E9",X"05",X"3A",X"02",X"81",X"CB",X"47",X"C2",
		X"0E",X"06",X"21",X"10",X"18",X"11",X"60",X"82",X"3E",X"09",X"08",X"C3",X"E9",X"05",X"CD",X"4C",
		X"04",X"21",X"8A",X"18",X"11",X"00",X"82",X"3E",X"0A",X"08",X"C3",X"E9",X"05",X"CD",X"4C",X"04",
		X"21",X"1D",X"19",X"11",X"E0",X"82",X"3E",X"0B",X"08",X"C3",X"E9",X"05",X"CD",X"4C",X"04",X"21",
		X"3F",X"1A",X"11",X"00",X"82",X"3E",X"0C",X"08",X"C3",X"E9",X"05",X"CD",X"4C",X"04",X"21",X"E5",
		X"1A",X"11",X"00",X"82",X"3E",X"0D",X"08",X"C3",X"E9",X"05",X"CD",X"4C",X"04",X"21",X"79",X"1B",
		X"11",X"00",X"82",X"3E",X"0E",X"08",X"C3",X"E9",X"05",X"7E",X"23",X"66",X"6F",X"46",X"23",X"C5",
		X"7E",X"23",X"E5",X"FE",X"FF",X"28",X"1D",X"66",X"6F",X"01",X"0E",X"00",X"ED",X"B0",X"08",X"12",
		X"08",X"13",X"AF",X"06",X"11",X"12",X"13",X"10",X"FC",X"E1",X"23",X"C1",X"10",X"E1",X"3E",X"80",
		X"32",X"00",X"81",X"C9",X"EB",X"01",X"20",X"00",X"09",X"EB",X"18",X"ED",X"00",X"00",X"FF",X"03",
		X"C7",X"03",X"90",X"03",X"5D",X"03",X"2D",X"03",X"FF",X"02",X"D4",X"02",X"AB",X"02",X"85",X"02",
		X"61",X"02",X"3F",X"02",X"1E",X"02",X"00",X"02",X"E3",X"01",X"C8",X"01",X"AF",X"01",X"96",X"01",
		X"80",X"01",X"6A",X"01",X"56",X"01",X"43",X"01",X"30",X"01",X"1F",X"01",X"0F",X"01",X"00",X"01",
		X"F2",X"00",X"E4",X"00",X"D7",X"00",X"CB",X"00",X"C0",X"00",X"B5",X"00",X"AB",X"00",X"A1",X"00",
		X"98",X"00",X"90",X"00",X"88",X"00",X"80",X"00",X"79",X"00",X"72",X"00",X"6C",X"00",X"66",X"00",
		X"60",X"00",X"5B",X"00",X"55",X"00",X"51",X"00",X"4C",X"00",X"48",X"00",X"44",X"00",X"40",X"00",
		X"3C",X"00",X"39",X"00",X"36",X"00",X"33",X"00",X"30",X"00",X"2D",X"00",X"2B",X"00",X"28",X"00",
		X"26",X"00",X"24",X"00",X"22",X"00",X"16",X"00",X"6A",X"06",X"08",X"29",X"30",X"01",X"19",X"10",
		X"FA",X"C9",X"06",X"08",X"ED",X"6A",X"7C",X"38",X"03",X"BB",X"38",X"03",X"93",X"67",X"B7",X"10",
		X"F3",X"7D",X"17",X"2F",X"C9",X"06",X"24",X"11",X"20",X"00",X"21",X"00",X"82",X"3A",X"01",X"81",
		X"0F",X"30",X"02",X"CB",X"D6",X"19",X"10",X"F8",X"C9",X"3A",X"01",X"81",X"06",X"08",X"21",X"00",
		X"82",X"11",X"20",X"00",X"0F",X"30",X"02",X"CB",X"96",X"19",X"10",X"F8",X"C9",X"0F",X"00",X"10",
		X"7C",X"10",X"A4",X"11",X"CC",X"12",X"3F",X"13",X"4D",X"14",X"CF",X"15",X"81",X"17",X"CE",X"17",
		X"10",X"18",X"8A",X"18",X"1D",X"19",X"3F",X"1A",X"E5",X"1A",X"79",X"1B",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"06",X"10",X"59",X"10",X"75",X"10",X"01",X"09",X"10",X"80",X"20",X"00",X"00",X"00",X"01",X"00",
		X"16",X"10",X"02",X"20",X"00",X"00",X"81",X"06",X"86",X"02",X"87",X"00",X"82",X"0E",X"1B",X"06",
		X"1B",X"03",X"22",X"03",X"27",X"03",X"2A",X"06",X"23",X"06",X"22",X"06",X"1E",X"06",X"1E",X"03",
		X"22",X"03",X"25",X"03",X"2A",X"03",X"25",X"03",X"22",X"03",X"20",X"06",X"20",X"03",X"24",X"03",
		X"27",X"03",X"2C",X"06",X"27",X"06",X"24",X"06",X"23",X"06",X"22",X"03",X"22",X"03",X"24",X"06",
		X"24",X"03",X"24",X"03",X"26",X"06",X"8A",X"1E",X"10",X"5D",X"10",X"6E",X"10",X"AB",X"BC",X"CD",
		X"DE",X"EF",X"FF",X"FE",X"ED",X"DC",X"CB",X"BA",X"A9",X"98",X"87",X"76",X"65",X"01",X"CD",X"EF",
		X"FE",X"DC",X"BA",X"98",X"01",X"77",X"10",X"AB",X"CD",X"DC",X"BA",X"00",X"82",X"10",X"91",X"11",
		X"9F",X"11",X"08",X"93",X"10",X"A0",X"10",X"AD",X"10",X"BA",X"10",X"C7",X"10",X"D4",X"10",X"E1",
		X"10",X"EE",X"10",X"80",X"20",X"00",X"00",X"00",X"01",X"00",X"FB",X"10",X"02",X"20",X"00",X"00",
		X"80",X"21",X"00",X"00",X"00",X"20",X"00",X"46",X"11",X"02",X"20",X"00",X"00",X"00",X"22",X"00",
		X"00",X"00",X"20",X"00",X"46",X"11",X"02",X"20",X"00",X"00",X"00",X"23",X"00",X"00",X"00",X"20",
		X"00",X"46",X"11",X"02",X"20",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"20",X"00",X"46",X"11",
		X"02",X"20",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"20",X"00",X"46",X"11",X"02",X"20",X"00",
		X"00",X"00",X"12",X"00",X"00",X"00",X"20",X"00",X"46",X"11",X"02",X"20",X"00",X"00",X"00",X"13",
		X"00",X"00",X"00",X"20",X"00",X"46",X"11",X"02",X"20",X"00",X"00",X"81",X"0B",X"86",X"01",X"82",
		X"0A",X"87",X"01",X"86",X"02",X"22",X"02",X"86",X"02",X"27",X"02",X"86",X"02",X"22",X"02",X"86",
		X"02",X"27",X"02",X"86",X"02",X"20",X"02",X"86",X"02",X"25",X"02",X"86",X"02",X"20",X"02",X"86",
		X"02",X"25",X"02",X"86",X"02",X"1E",X"02",X"86",X"02",X"24",X"02",X"86",X"02",X"1E",X"02",X"86",
		X"02",X"24",X"02",X"86",X"02",X"1D",X"02",X"86",X"02",X"22",X"02",X"86",X"02",X"1D",X"02",X"86",
		X"02",X"22",X"02",X"8A",X"03",X"11",X"81",X"0B",X"86",X"01",X"82",X"0A",X"87",X"01",X"86",X"02",
		X"22",X"02",X"86",X"02",X"27",X"02",X"86",X"02",X"22",X"02",X"86",X"02",X"27",X"02",X"86",X"02",
		X"20",X"02",X"86",X"02",X"25",X"02",X"86",X"02",X"20",X"02",X"86",X"02",X"25",X"02",X"86",X"02",
		X"1E",X"02",X"86",X"02",X"24",X"02",X"86",X"02",X"1E",X"02",X"86",X"02",X"24",X"02",X"86",X"02",
		X"1D",X"02",X"86",X"02",X"22",X"02",X"86",X"02",X"1D",X"02",X"86",X"02",X"22",X"02",X"8A",X"4E",
		X"11",X"95",X"11",X"9A",X"11",X"EF",X"FE",X"DC",X"BA",X"02",X"EF",X"FE",X"DC",X"BA",X"01",X"A1",
		X"11",X"CD",X"ED",X"00",X"AA",X"11",X"B9",X"12",X"C7",X"12",X"08",X"BB",X"11",X"C8",X"11",X"D5",
		X"11",X"E2",X"11",X"EF",X"11",X"FC",X"11",X"09",X"12",X"16",X"12",X"80",X"20",X"00",X"00",X"00",
		X"01",X"00",X"23",X"12",X"02",X"20",X"00",X"00",X"80",X"21",X"00",X"00",X"00",X"20",X"00",X"6E",
		X"12",X"02",X"20",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"20",X"00",X"6E",X"12",X"02",X"20",
		X"00",X"00",X"00",X"23",X"00",X"00",X"00",X"20",X"00",X"6E",X"12",X"02",X"20",X"00",X"00",X"00",
		X"10",X"00",X"00",X"00",X"20",X"00",X"6E",X"12",X"02",X"20",X"00",X"00",X"00",X"11",X"00",X"00",
		X"00",X"20",X"00",X"6E",X"12",X"02",X"20",X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"20",X"00",
		X"6E",X"12",X"02",X"20",X"00",X"00",X"00",X"13",X"00",X"00",X"00",X"20",X"00",X"6E",X"12",X"02",
		X"20",X"00",X"00",X"81",X"0B",X"86",X"01",X"82",X"0D",X"87",X"01",X"86",X"02",X"22",X"02",X"86",
		X"02",X"27",X"02",X"86",X"02",X"22",X"02",X"86",X"02",X"27",X"02",X"86",X"02",X"20",X"02",X"86",
		X"02",X"25",X"02",X"86",X"02",X"20",X"02",X"86",X"02",X"25",X"02",X"86",X"02",X"1E",X"02",X"86",
		X"02",X"24",X"02",X"86",X"02",X"1E",X"02",X"86",X"02",X"24",X"02",X"86",X"02",X"1D",X"02",X"86",
		X"02",X"22",X"02",X"86",X"02",X"1D",X"02",X"86",X"02",X"22",X"02",X"8A",X"2B",X"12",X"81",X"0B",
		X"86",X"01",X"82",X"0D",X"87",X"01",X"86",X"02",X"22",X"02",X"86",X"02",X"27",X"02",X"86",X"02",
		X"22",X"02",X"86",X"02",X"27",X"02",X"86",X"02",X"20",X"02",X"86",X"02",X"25",X"02",X"86",X"02",
		X"20",X"02",X"86",X"02",X"25",X"02",X"86",X"02",X"1E",X"02",X"86",X"02",X"24",X"02",X"86",X"02",
		X"1E",X"02",X"86",X"02",X"24",X"02",X"86",X"02",X"1D",X"02",X"86",X"02",X"22",X"02",X"86",X"02",
		X"1D",X"02",X"86",X"02",X"22",X"02",X"8A",X"76",X"12",X"BD",X"12",X"C2",X"12",X"EF",X"FE",X"DC",
		X"BA",X"02",X"EF",X"FE",X"DC",X"BA",X"01",X"C9",X"12",X"CD",X"ED",X"00",X"D2",X"12",X"FF",X"12",
		X"0F",X"13",X"01",X"D5",X"12",X"80",X"11",X"00",X"00",X"00",X"01",X"00",X"E2",X"12",X"00",X"20",
		X"00",X"00",X"82",X"0F",X"81",X"03",X"87",X"00",X"86",X"01",X"30",X"05",X"34",X"05",X"32",X"05",
		X"37",X"05",X"32",X"05",X"34",X"05",X"30",X"05",X"34",X"05",X"32",X"05",X"37",X"05",X"84",X"03",
		X"13",X"0B",X"13",X"DE",X"FF",X"FE",X"DC",X"BA",X"98",X"76",X"01",X"EF",X"FE",X"DC",X"02",X"13",
		X"13",X"29",X"13",X"FF",X"FF",X"FF",X"FF",X"EE",X"DD",X"EE",X"DD",X"EE",X"DD",X"EE",X"DD",X"EE",
		X"DD",X"EE",X"DD",X"EE",X"DD",X"EE",X"DD",X"EE",X"02",X"FF",X"FF",X"FF",X"FF",X"EE",X"EE",X"DD",
		X"DD",X"EE",X"EE",X"DD",X"DD",X"EE",X"EE",X"DD",X"DD",X"EE",X"EE",X"DD",X"DD",X"DD",X"02",X"45",
		X"13",X"24",X"14",X"3F",X"14",X"08",X"56",X"13",X"63",X"13",X"70",X"13",X"7D",X"13",X"8A",X"13",
		X"97",X"13",X"A4",X"13",X"B1",X"13",X"80",X"20",X"00",X"00",X"00",X"01",X"00",X"BE",X"13",X"02",
		X"20",X"00",X"00",X"80",X"21",X"00",X"00",X"00",X"01",X"00",X"D9",X"13",X"02",X"20",X"00",X"00",
		X"00",X"22",X"00",X"00",X"00",X"01",X"00",X"D9",X"13",X"02",X"20",X"00",X"00",X"00",X"23",X"00",
		X"00",X"00",X"01",X"00",X"D9",X"13",X"02",X"20",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"01",
		X"00",X"D9",X"13",X"02",X"20",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"01",X"00",X"D9",X"13",
		X"02",X"20",X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"01",X"00",X"D9",X"13",X"02",X"20",X"00",
		X"00",X"00",X"13",X"00",X"00",X"00",X"01",X"00",X"D9",X"13",X"02",X"20",X"00",X"00",X"81",X"0B",
		X"86",X"01",X"82",X"0D",X"87",X"00",X"1D",X"02",X"1F",X"02",X"20",X"02",X"22",X"02",X"20",X"02",
		X"1F",X"02",X"1D",X"02",X"1D",X"02",X"8A",X"C6",X"13",X"81",X"0B",X"86",X"01",X"82",X"0D",X"87",
		X"00",X"1D",X"02",X"20",X"02",X"1D",X"02",X"20",X"02",X"1D",X"02",X"20",X"02",X"1D",X"02",X"20",
		X"02",X"1B",X"02",X"1F",X"02",X"1B",X"02",X"1F",X"02",X"1B",X"02",X"1F",X"02",X"1B",X"02",X"1F",
		X"02",X"19",X"02",X"1D",X"02",X"19",X"02",X"1D",X"02",X"19",X"02",X"1D",X"02",X"19",X"02",X"1D",
		X"02",X"1B",X"02",X"1F",X"02",X"1B",X"02",X"1F",X"02",X"1B",X"02",X"1F",X"02",X"1B",X"02",X"1F",
		X"02",X"8A",X"E1",X"13",X"2A",X"14",X"31",X"14",X"38",X"14",X"EF",X"FE",X"DC",X"BA",X"A9",X"87",
		X"01",X"9A",X"AB",X"BC",X"CD",X"DE",X"EE",X"01",X"EF",X"FF",X"FF",X"FD",X"A8",X"65",X"01",X"43",
		X"14",X"47",X"14",X"DE",X"FF",X"ED",X"00",X"CD",X"ED",X"DC",X"BA",X"BC",X"00",X"53",X"14",X"4C",
		X"15",X"93",X"15",X"08",X"64",X"14",X"71",X"14",X"7E",X"14",X"8B",X"14",X"98",X"14",X"A5",X"14",
		X"B2",X"14",X"BF",X"14",X"80",X"20",X"00",X"00",X"00",X"05",X"00",X"CC",X"14",X"02",X"20",X"00",
		X"00",X"80",X"21",X"00",X"00",X"00",X"01",X"00",X"F4",X"14",X"02",X"20",X"00",X"00",X"00",X"22",
		X"00",X"00",X"00",X"01",X"00",X"F4",X"14",X"02",X"20",X"00",X"00",X"00",X"23",X"00",X"00",X"00",
		X"01",X"00",X"F4",X"14",X"02",X"20",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"01",X"00",X"F4",
		X"14",X"02",X"20",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"01",X"00",X"F4",X"14",X"02",X"20",
		X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"01",X"00",X"F4",X"14",X"02",X"20",X"00",X"00",X"00",
		X"13",X"00",X"00",X"00",X"01",X"00",X"F4",X"14",X"02",X"20",X"00",X"00",X"81",X"11",X"86",X"01",
		X"87",X"00",X"82",X"0F",X"8D",X"2A",X"0D",X"0D",X"8E",X"81",X"0B",X"86",X"02",X"82",X"0E",X"87",
		X"00",X"1D",X"02",X"1F",X"02",X"20",X"02",X"22",X"02",X"20",X"02",X"1F",X"02",X"1D",X"02",X"1D",
		X"02",X"8A",X"E1",X"14",X"81",X"11",X"86",X"01",X"87",X"00",X"82",X"0F",X"8D",X"2C",X"0D",X"0D",
		X"8E",X"81",X"0B",X"86",X"02",X"82",X"0E",X"87",X"00",X"1D",X"02",X"20",X"02",X"1D",X"02",X"20",
		X"02",X"1D",X"02",X"20",X"02",X"1D",X"02",X"20",X"02",X"1B",X"02",X"1F",X"02",X"1B",X"02",X"1F",
		X"02",X"1B",X"02",X"1F",X"02",X"1B",X"02",X"1F",X"02",X"19",X"02",X"1D",X"02",X"19",X"02",X"1D",
		X"02",X"19",X"02",X"1D",X"02",X"19",X"02",X"1D",X"02",X"1B",X"02",X"1F",X"02",X"1B",X"02",X"1F",
		X"02",X"1B",X"02",X"1F",X"02",X"1B",X"02",X"1F",X"02",X"8A",X"09",X"15",X"54",X"15",X"80",X"15",
		X"85",X"15",X"8C",X"15",X"11",X"12",X"23",X"34",X"45",X"56",X"67",X"78",X"89",X"9A",X"AB",X"BC",
		X"CD",X"DE",X"EF",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"FE",X"FE",X"FE",X"FE",X"ED",X"DC",X"CB",X"BA",X"A9",X"98",X"87",X"76",X"65",X"43",X"21",X"01",
		X"EF",X"FE",X"DC",X"BA",X"01",X"9A",X"AB",X"BC",X"CD",X"DE",X"EE",X"01",X"EF",X"FF",X"FF",X"FD",
		X"A8",X"65",X"01",X"9B",X"15",X"B0",X"15",X"C5",X"15",X"C9",X"15",X"DD",X"DD",X"EF",X"FE",X"DC",
		X"BB",X"CD",X"DE",X"EF",X"FE",X"DC",X"BB",X"CD",X"EF",X"FE",X"DC",X"BB",X"CD",X"EF",X"FE",X"00",
		X"EE",X"EE",X"DD",X"DD",X"EE",X"EE",X"DD",X"DD",X"EE",X"EE",X"DD",X"DD",X"EE",X"EE",X"DD",X"DD",
		X"EE",X"EE",X"DD",X"DD",X"00",X"DE",X"FF",X"ED",X"00",X"CD",X"ED",X"DC",X"BA",X"BC",X"00",X"D5",
		X"15",X"00",X"17",X"47",X"17",X"08",X"E6",X"15",X"F3",X"15",X"00",X"16",X"0D",X"16",X"1A",X"16",
		X"27",X"16",X"34",X"16",X"41",X"16",X"80",X"20",X"00",X"00",X"00",X"01",X"00",X"4E",X"16",X"02",
		X"20",X"00",X"00",X"80",X"21",X"00",X"00",X"00",X"05",X"00",X"A6",X"16",X"02",X"20",X"00",X"00",
		X"00",X"22",X"00",X"00",X"00",X"05",X"00",X"A6",X"16",X"02",X"20",X"00",X"00",X"00",X"23",X"00",
		X"00",X"00",X"05",X"00",X"A6",X"16",X"02",X"20",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"05",
		X"00",X"A6",X"16",X"02",X"20",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"05",X"00",X"A6",X"16",
		X"02",X"20",X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"05",X"00",X"A6",X"16",X"02",X"20",X"00",
		X"00",X"00",X"13",X"00",X"00",X"00",X"05",X"00",X"A6",X"16",X"02",X"20",X"00",X"00",X"81",X"11",
		X"86",X"01",X"87",X"00",X"82",X"0F",X"8D",X"2C",X"0D",X"0D",X"8E",X"81",X"0B",X"86",X"03",X"82",
		X"0D",X"87",X"04",X"86",X"02",X"22",X"02",X"86",X"02",X"27",X"02",X"86",X"02",X"22",X"02",X"86",
		X"02",X"27",X"02",X"86",X"02",X"20",X"02",X"86",X"02",X"25",X"02",X"86",X"02",X"20",X"02",X"86",
		X"02",X"25",X"02",X"86",X"02",X"1E",X"02",X"86",X"02",X"24",X"02",X"86",X"02",X"1E",X"02",X"86",
		X"02",X"24",X"02",X"86",X"02",X"1D",X"02",X"86",X"02",X"22",X"02",X"86",X"02",X"1D",X"02",X"86",
		X"02",X"22",X"02",X"8A",X"63",X"16",X"81",X"11",X"86",X"01",X"87",X"00",X"82",X"0F",X"00",X"03",
		X"8D",X"2C",X"0D",X"0A",X"8E",X"81",X"0B",X"86",X"04",X"82",X"0D",X"87",X"04",X"86",X"02",X"22",
		X"02",X"86",X"02",X"27",X"02",X"86",X"02",X"22",X"02",X"86",X"02",X"27",X"02",X"86",X"02",X"20",
		X"02",X"86",X"02",X"25",X"02",X"86",X"02",X"20",X"02",X"86",X"02",X"25",X"02",X"86",X"02",X"1E",
		X"02",X"86",X"02",X"24",X"02",X"86",X"02",X"1E",X"02",X"86",X"02",X"24",X"02",X"86",X"02",X"1D",
		X"02",X"86",X"02",X"22",X"02",X"86",X"02",X"1D",X"02",X"86",X"02",X"22",X"02",X"8A",X"BD",X"16",
		X"08",X"17",X"34",X"17",X"39",X"17",X"40",X"17",X"11",X"12",X"23",X"34",X"45",X"56",X"67",X"78",
		X"89",X"9A",X"AB",X"BC",X"CD",X"DE",X"EF",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"ED",X"DC",X"CB",X"BA",X"A9",X"98",X"87",X"76",
		X"65",X"43",X"21",X"01",X"EF",X"FE",X"DC",X"BA",X"01",X"9A",X"AB",X"BC",X"CD",X"DE",X"EE",X"01",
		X"EF",X"FF",X"FF",X"FD",X"A8",X"65",X"01",X"4F",X"17",X"64",X"17",X"79",X"17",X"7D",X"17",X"DD",
		X"DD",X"EF",X"FE",X"DC",X"BB",X"CD",X"DE",X"EF",X"FE",X"DC",X"BB",X"CD",X"EF",X"FE",X"DC",X"BB",
		X"CD",X"EF",X"FE",X"00",X"EE",X"EE",X"DD",X"DD",X"EE",X"EE",X"DD",X"DD",X"EE",X"EE",X"DD",X"DD",
		X"EE",X"EE",X"DD",X"DD",X"EE",X"EE",X"DD",X"DD",X"00",X"DE",X"FF",X"ED",X"00",X"CD",X"ED",X"DC",
		X"00",X"87",X"17",X"AB",X"17",X"C7",X"17",X"01",X"8A",X"17",X"80",X"13",X"00",X"00",X"00",X"01",
		X"00",X"97",X"17",X"00",X"20",X"00",X"00",X"82",X"0D",X"81",X"04",X"86",X"00",X"85",X"03",X"87",
		X"00",X"8F",X"8D",X"00",X"09",X"00",X"03",X"08",X"8E",X"90",X"84",X"AF",X"17",X"BF",X"17",X"FE",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"ED",X"DC",X"CB",X"BA",X"A9",X"98",X"86",X"01",X"FF",
		X"FF",X"DD",X"BB",X"AA",X"88",X"66",X"02",X"C9",X"17",X"CD",X"EF",X"FE",X"DC",X"00",X"D2",X"17",
		X"0B",X"18",X"01",X"D5",X"17",X"80",X"10",X"00",X"00",X"00",X"01",X"00",X"E2",X"17",X"08",X"20",
		X"00",X"00",X"82",X"0A",X"86",X"00",X"81",X"04",X"87",X"01",X"8D",X"2A",X"27",X"03",X"8E",X"8D",
		X"27",X"24",X"04",X"8E",X"8D",X"24",X"1F",X"04",X"8E",X"8D",X"21",X"1E",X"05",X"8E",X"8D",X"1E",
		X"1B",X"06",X"8E",X"8D",X"1B",X"24",X"07",X"8E",X"84",X"0B",X"18",X"CD",X"EF",X"FE",X"DC",X"00",
		X"14",X"18",X"6E",X"18",X"01",X"17",X"18",X"80",X"23",X"00",X"00",X"00",X"01",X"00",X"24",X"18",
		X"00",X"20",X"00",X"00",X"82",X"0F",X"81",X"04",X"86",X"00",X"85",X"03",X"8F",X"00",X"07",X"02",
		X"90",X"8F",X"00",X"05",X"02",X"90",X"8F",X"00",X"03",X"01",X"90",X"8F",X"00",X"01",X"02",X"90",
		X"8F",X"00",X"08",X"01",X"90",X"8F",X"00",X"06",X"01",X"90",X"8F",X"00",X"04",X"01",X"90",X"8F",
		X"00",X"02",X"01",X"90",X"8F",X"00",X"01",X"02",X"90",X"8F",X"00",X"08",X"01",X"90",X"8F",X"00",
		X"02",X"02",X"90",X"8F",X"00",X"06",X"01",X"90",X"8F",X"00",X"08",X"01",X"90",X"84",X"72",X"18",
		X"82",X"18",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"ED",X"DC",X"CB",X"BA",X"A9",X"98",
		X"86",X"01",X"FF",X"FF",X"DD",X"BB",X"AA",X"88",X"66",X"02",X"90",X"18",X"DD",X"18",X"ED",X"18",
		X"02",X"95",X"18",X"A2",X"18",X"80",X"20",X"00",X"00",X"00",X"01",X"00",X"AF",X"18",X"0E",X"20",
		X"00",X"00",X"80",X"21",X"00",X"00",X"00",X"14",X"00",X"C6",X"18",X"0E",X"20",X"00",X"00",X"82",
		X"0F",X"81",X"04",X"87",X"00",X"86",X"01",X"19",X"05",X"1C",X"05",X"1E",X"05",X"86",X"02",X"21",
		X"05",X"00",X"05",X"8A",X"B5",X"18",X"82",X"0F",X"81",X"04",X"87",X"00",X"86",X"01",X"19",X"05",
		X"1C",X"05",X"1E",X"05",X"86",X"02",X"21",X"05",X"00",X"05",X"8A",X"CC",X"18",X"E1",X"18",X"E7",
		X"18",X"DE",X"FF",X"FF",X"FF",X"ED",X"01",X"DC",X"BA",X"98",X"76",X"54",X"01",X"F1",X"18",X"07",
		X"19",X"FF",X"FF",X"FF",X"FF",X"EE",X"DD",X"EE",X"DD",X"EE",X"DD",X"EE",X"DD",X"EE",X"DD",X"EE",
		X"DD",X"EE",X"DD",X"EE",X"DD",X"EE",X"00",X"FF",X"FF",X"FF",X"FF",X"EE",X"EE",X"DD",X"DD",X"EE",
		X"EE",X"DD",X"DD",X"EE",X"EE",X"DD",X"DD",X"EE",X"EE",X"DD",X"DD",X"DD",X"00",X"23",X"19",X"90",
		X"19",X"9F",X"19",X"01",X"26",X"19",X"80",X"13",X"00",X"00",X"00",X"01",X"00",X"33",X"19",X"00",
		X"20",X"00",X"00",X"81",X"06",X"86",X"00",X"85",X"03",X"85",X"07",X"82",X"0F",X"8F",X"00",X"20",
		X"05",X"90",X"82",X"0E",X"8F",X"00",X"21",X"05",X"90",X"82",X"0D",X"8F",X"00",X"1F",X"05",X"90",
		X"82",X"0C",X"8F",X"00",X"21",X"05",X"90",X"82",X"0B",X"8F",X"00",X"1F",X"05",X"90",X"82",X"0A",
		X"8F",X"00",X"21",X"04",X"90",X"82",X"09",X"8F",X"00",X"1F",X"04",X"90",X"82",X"08",X"8F",X"00",
		X"21",X"04",X"90",X"82",X"07",X"8F",X"00",X"1F",X"04",X"90",X"82",X"06",X"8F",X"00",X"21",X"04",
		X"90",X"82",X"05",X"8F",X"00",X"1F",X"03",X"90",X"82",X"04",X"8F",X"00",X"21",X"03",X"90",X"84",
		X"92",X"19",X"FE",X"FE",X"DE",X"DE",X"CD",X"CD",X"BC",X"BC",X"AB",X"AB",X"89",X"89",X"02",X"A1",
		X"19",X"FF",X"DD",X"FF",X"DD",X"00",X"AA",X"19",X"2C",X"1A",X"01",X"AD",X"19",X"80",X"11",X"00",
		X"00",X"00",X"01",X"00",X"BA",X"19",X"00",X"20",X"00",X"00",X"82",X"0F",X"81",X"04",X"86",X"00",
		X"87",X"00",X"82",X"0F",X"8D",X"33",X"3B",X"06",X"8E",X"82",X"0E",X"8D",X"33",X"3B",X"06",X"8E",
		X"82",X"0D",X"8D",X"33",X"3B",X"06",X"8E",X"82",X"0C",X"8D",X"33",X"3B",X"06",X"8E",X"82",X"0B",
		X"8D",X"33",X"3B",X"06",X"8E",X"82",X"0A",X"8D",X"33",X"3B",X"06",X"8E",X"82",X"09",X"8D",X"33",
		X"3B",X"06",X"8E",X"82",X"08",X"8D",X"33",X"3B",X"06",X"8E",X"82",X"07",X"8D",X"33",X"3B",X"06",
		X"8E",X"82",X"06",X"8D",X"33",X"3B",X"06",X"8E",X"82",X"05",X"8D",X"33",X"3B",X"06",X"8E",X"82",
		X"04",X"8D",X"33",X"3B",X"06",X"8E",X"82",X"03",X"8D",X"33",X"3B",X"06",X"8E",X"82",X"02",X"8D",
		X"33",X"3B",X"06",X"8E",X"82",X"01",X"8D",X"33",X"3B",X"06",X"8E",X"84",X"30",X"1A",X"37",X"1A",
		X"FE",X"DC",X"BA",X"98",X"87",X"65",X"01",X"FF",X"FF",X"DD",X"BB",X"AA",X"88",X"66",X"02",X"45",
		X"1A",X"CC",X"1A",X"DE",X"1A",X"02",X"4A",X"1A",X"57",X"1A",X"80",X"20",X"00",X"00",X"00",X"01",
		X"00",X"64",X"1A",X"03",X"20",X"00",X"00",X"80",X"21",X"00",X"00",X"00",X"01",X"00",X"98",X"1A",
		X"03",X"20",X"00",X"00",X"81",X"0B",X"86",X"02",X"87",X"00",X"82",X"0F",X"19",X"04",X"00",X"02",
		X"86",X"02",X"18",X"02",X"18",X"02",X"18",X"02",X"86",X"01",X"19",X"04",X"00",X"02",X"1B",X"02",
		X"1B",X"02",X"1B",X"02",X"8C",X"00",X"02",X"6C",X"1A",X"86",X"02",X"19",X"02",X"00",X"02",X"1B",
		X"02",X"00",X"02",X"86",X"01",X"1D",X"0C",X"84",X"81",X"0B",X"86",X"02",X"87",X"00",X"82",X"0F",
		X"20",X"04",X"00",X"02",X"86",X"02",X"1F",X"02",X"1F",X"02",X"1F",X"02",X"86",X"01",X"20",X"04",
		X"00",X"02",X"22",X"02",X"22",X"02",X"22",X"02",X"8C",X"01",X"02",X"A0",X"1A",X"86",X"02",X"20",
		X"02",X"00",X"02",X"22",X"02",X"00",X"02",X"86",X"01",X"24",X"0C",X"84",X"D0",X"1A",X"D9",X"1A",
		X"EF",X"FF",X"FE",X"ED",X"DC",X"CB",X"BA",X"98",X"01",X"EF",X"FE",X"DC",X"BA",X"01",X"E0",X"1A",
		X"AB",X"CD",X"DC",X"BA",X"00",X"EB",X"1A",X"5E",X"1B",X"70",X"1B",X"02",X"F0",X"1A",X"FD",X"1A",
		X"80",X"20",X"00",X"00",X"00",X"01",X"00",X"0A",X"1B",X"FC",X"20",X"00",X"00",X"80",X"21",X"00",
		X"00",X"00",X"05",X"00",X"34",X"1B",X"08",X"20",X"00",X"00",X"81",X"04",X"86",X"02",X"87",X"00",
		X"82",X"0F",X"1E",X"06",X"22",X"06",X"24",X"06",X"2A",X"06",X"29",X"06",X"27",X"06",X"25",X"06",
		X"24",X"06",X"22",X"06",X"21",X"06",X"20",X"06",X"1E",X"06",X"1F",X"06",X"27",X"06",X"8C",X"00",
		X"02",X"18",X"1B",X"84",X"81",X"04",X"86",X"02",X"87",X"00",X"82",X"0F",X"1E",X"06",X"22",X"06",
		X"24",X"06",X"2A",X"06",X"29",X"06",X"27",X"06",X"25",X"06",X"24",X"06",X"22",X"06",X"21",X"06",
		X"20",X"06",X"1E",X"06",X"1F",X"06",X"27",X"06",X"8C",X"01",X"02",X"42",X"1B",X"84",X"62",X"1B",
		X"69",X"1B",X"CD",X"EF",X"FE",X"ED",X"DC",X"CB",X"01",X"CD",X"EF",X"FE",X"DC",X"BA",X"98",X"01",
		X"72",X"1B",X"AB",X"CD",X"EF",X"FE",X"DC",X"BA",X"00",X"7F",X"1B",X"6F",X"1E",X"A1",X"1E",X"08",
		X"90",X"1B",X"9D",X"1B",X"AA",X"1B",X"B7",X"1B",X"C4",X"1B",X"D1",X"1B",X"DE",X"1B",X"EB",X"1B",
		X"80",X"20",X"00",X"00",X"00",X"01",X"00",X"F8",X"1B",X"00",X"20",X"00",X"00",X"80",X"21",X"00",
		X"00",X"00",X"01",X"00",X"F0",X"1C",X"00",X"20",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"01",
		X"00",X"E8",X"1D",X"00",X"20",X"00",X"00",X"00",X"23",X"00",X"00",X"00",X"01",X"00",X"42",X"1E",
		X"00",X"20",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"01",X"00",X"E8",X"1D",X"00",X"20",X"00",
		X"00",X"80",X"11",X"00",X"00",X"00",X"01",X"00",X"17",X"1E",X"00",X"20",X"00",X"00",X"80",X"12",
		X"00",X"00",X"00",X"01",X"00",X"42",X"1E",X"00",X"20",X"00",X"00",X"00",X"13",X"00",X"00",X"00",
		X"01",X"00",X"42",X"1E",X"00",X"20",X"00",X"00",X"86",X"01",X"87",X"00",X"82",X"0F",X"81",X"0A",
		X"00",X"0A",X"8D",X"12",X"19",X"07",X"19",X"25",X"0B",X"25",X"31",X"11",X"31",X"3C",X"14",X"8E",
		X"81",X"0C",X"86",X"00",X"87",X"00",X"82",X"0F",X"8D",X"30",X"38",X"06",X"8E",X"82",X"0F",X"8D",
		X"2C",X"34",X"06",X"8E",X"82",X"0F",X"8D",X"2C",X"34",X"06",X"8E",X"82",X"0E",X"8D",X"30",X"38",
		X"06",X"8E",X"82",X"0E",X"8D",X"30",X"38",X"06",X"8E",X"82",X"0D",X"8D",X"30",X"38",X"06",X"8E",
		X"82",X"0D",X"8D",X"30",X"38",X"06",X"8E",X"82",X"0C",X"8D",X"30",X"38",X"06",X"8E",X"82",X"0C",
		X"8D",X"30",X"38",X"06",X"8E",X"82",X"0B",X"8D",X"30",X"38",X"06",X"8E",X"82",X"0B",X"8D",X"30",
		X"38",X"06",X"8E",X"82",X"0A",X"8D",X"30",X"38",X"06",X"8E",X"82",X"0A",X"8D",X"30",X"38",X"06",
		X"8E",X"82",X"09",X"8D",X"30",X"38",X"06",X"8E",X"82",X"09",X"8D",X"30",X"38",X"06",X"8E",X"82",
		X"08",X"8D",X"30",X"38",X"06",X"8E",X"82",X"08",X"8D",X"30",X"38",X"06",X"8E",X"82",X"07",X"8D",
		X"30",X"38",X"06",X"8E",X"82",X"07",X"8D",X"30",X"38",X"06",X"8E",X"82",X"06",X"8D",X"30",X"38",
		X"06",X"8E",X"82",X"06",X"8D",X"30",X"38",X"06",X"8E",X"82",X"05",X"8D",X"30",X"38",X"06",X"8E",
		X"82",X"05",X"8D",X"30",X"38",X"06",X"8E",X"82",X"04",X"8D",X"30",X"38",X"06",X"8E",X"82",X"04",
		X"8D",X"30",X"38",X"06",X"8E",X"82",X"03",X"8D",X"30",X"38",X"06",X"8E",X"82",X"03",X"8D",X"30",
		X"38",X"06",X"8E",X"82",X"02",X"8D",X"30",X"38",X"06",X"8E",X"82",X"02",X"8D",X"30",X"38",X"06",
		X"8E",X"82",X"01",X"8D",X"30",X"38",X"06",X"8E",X"82",X"01",X"8D",X"30",X"38",X"06",X"8E",X"84",
		X"86",X"01",X"87",X"00",X"82",X"0F",X"81",X"0A",X"00",X"0F",X"8D",X"12",X"1B",X"05",X"1B",X"27",
		X"0A",X"27",X"33",X"0F",X"31",X"3C",X"14",X"8E",X"81",X"0C",X"86",X"00",X"87",X"00",X"82",X"0F",
		X"8D",X"2C",X"34",X"06",X"8E",X"82",X"0F",X"8D",X"2C",X"34",X"06",X"8E",X"82",X"0F",X"8D",X"2C",
		X"34",X"06",X"8E",X"82",X"0E",X"8D",X"2C",X"34",X"06",X"8E",X"82",X"0E",X"8D",X"2C",X"34",X"06",
		X"8E",X"82",X"0D",X"8D",X"2C",X"34",X"06",X"8E",X"82",X"0D",X"8D",X"2C",X"34",X"06",X"8E",X"82",
		X"0C",X"8D",X"2C",X"34",X"06",X"8E",X"82",X"0C",X"8D",X"2C",X"34",X"06",X"8E",X"82",X"0B",X"8D",
		X"2C",X"34",X"06",X"8E",X"82",X"0B",X"8D",X"2C",X"34",X"06",X"8E",X"82",X"0A",X"8D",X"2C",X"34",
		X"06",X"8E",X"82",X"0A",X"8D",X"2C",X"34",X"06",X"8E",X"82",X"09",X"8D",X"2C",X"34",X"06",X"8E",
		X"82",X"09",X"8D",X"2C",X"34",X"06",X"8E",X"82",X"08",X"8D",X"2C",X"34",X"06",X"8E",X"82",X"08",
		X"8D",X"2C",X"34",X"06",X"8E",X"82",X"07",X"8D",X"2C",X"34",X"06",X"8E",X"82",X"07",X"8D",X"2C",
		X"34",X"06",X"8E",X"82",X"06",X"8D",X"2C",X"34",X"06",X"8E",X"82",X"06",X"8D",X"2C",X"34",X"06",
		X"8E",X"82",X"05",X"8D",X"2C",X"34",X"06",X"8E",X"82",X"05",X"8D",X"2C",X"34",X"06",X"8E",X"82",
		X"04",X"8D",X"2C",X"34",X"06",X"8E",X"82",X"04",X"8D",X"2C",X"34",X"06",X"8E",X"82",X"03",X"8D",
		X"2C",X"34",X"06",X"8E",X"82",X"03",X"8D",X"2C",X"34",X"06",X"8E",X"82",X"02",X"8D",X"2C",X"34",
		X"06",X"8E",X"82",X"02",X"8D",X"2C",X"34",X"06",X"8E",X"82",X"01",X"8D",X"2C",X"34",X"06",X"8E",
		X"82",X"01",X"8D",X"2C",X"34",X"06",X"8E",X"84",X"81",X"05",X"86",X"00",X"87",X"00",X"82",X"0F",
		X"81",X"05",X"82",X"0F",X"8F",X"00",X"14",X"02",X"00",X"10",X"02",X"00",X"0C",X"02",X"00",X"10",
		X"02",X"90",X"81",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",
		X"00",X"0C",X"00",X"0C",X"00",X"06",X"84",X"86",X"01",X"87",X"00",X"82",X"0F",X"81",X"0A",X"8D",
		X"12",X"19",X"0A",X"19",X"25",X"0F",X"25",X"31",X"14",X"31",X"3C",X"14",X"8E",X"81",X"0C",X"00",
		X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",
		X"06",X"84",X"86",X"01",X"87",X"00",X"82",X"0F",X"81",X"0A",X"00",X"05",X"8D",X"0D",X"1E",X"0A",
		X"1E",X"25",X"0F",X"25",X"31",X"0F",X"31",X"3C",X"14",X"8E",X"81",X"0C",X"00",X"0C",X"00",X"0C",
		X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"06",X"84",X"73",
		X"1E",X"75",X"1E",X"F9",X"00",X"11",X"12",X"23",X"34",X"45",X"56",X"67",X"78",X"89",X"9A",X"AB",
		X"BC",X"CD",X"DE",X"EF",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"ED",X"DC",X"CB",X"BA",X"A9",X"98",X"87",X"76",X"65",X"43",X"21",
		X"01",X"A3",X"1E",X"DE",X"FE",X"DC",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
