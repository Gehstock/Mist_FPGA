library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity GALAXIAN_1K is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of GALAXIAN_1K is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
    x"38",x"7C",x"C2",x"82",x"86",x"7C",x"38",x"00", -- 0x0000
    x"02",x"02",x"FE",x"FE",x"42",x"02",x"00",x"00", -- 0x0008
    x"62",x"F2",x"BA",x"9A",x"9E",x"CE",x"46",x"00", -- 0x0010
    x"8C",x"DE",x"F2",x"B2",x"92",x"86",x"04",x"00", -- 0x0018
    x"08",x"FE",x"FE",x"C8",x"68",x"38",x"18",x"00", -- 0x0020
    x"1C",x"BE",x"A2",x"A2",x"A2",x"E6",x"E4",x"00", -- 0x0028
    x"0C",x"9E",x"92",x"92",x"D2",x"7E",x"3C",x"00", -- 0x0030
    x"C0",x"E0",x"B0",x"9E",x"8E",x"C0",x"C0",x"00", -- 0x0038
    x"0C",x"6E",x"9A",x"9A",x"B2",x"F2",x"6C",x"00", -- 0x0040
    x"78",x"FC",x"96",x"92",x"92",x"F2",x"60",x"00", -- 0x0048
    x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00", -- 0x0050
    x"00",x"00",x"00",x"00",x"08",x"FE",x"F0",x"F0", -- 0x0058
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0060
    x"00",x"00",x"00",x"04",x"06",x"00",x"00",x"02", -- 0x0068
    x"08",x"08",x"0C",x"08",x"08",x"00",x"00",x"00", -- 0x0070
    x"00",x"27",x"62",x"C0",x"90",x"62",x"27",x"00", -- 0x0078
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0080
    x"3E",x"7E",x"C8",x"88",x"C8",x"7E",x"3E",x"00", -- 0x0088
    x"6C",x"FE",x"92",x"92",x"92",x"FE",x"FE",x"00", -- 0x0090
    x"44",x"C6",x"82",x"82",x"C6",x"7C",x"38",x"00", -- 0x0098
    x"38",x"7C",x"C6",x"82",x"82",x"FE",x"FE",x"00", -- 0x00A0
    x"82",x"92",x"92",x"92",x"FE",x"FE",x"00",x"00", -- 0x00A8
    x"80",x"90",x"90",x"90",x"90",x"FE",x"FE",x"00", -- 0x00B0
    x"9E",x"9E",x"92",x"82",x"C6",x"7C",x"38",x"00", -- 0x00B8
    x"FE",x"FE",x"10",x"10",x"10",x"FE",x"FE",x"00", -- 0x00C0
    x"82",x"82",x"FE",x"FE",x"82",x"82",x"00",x"00", -- 0x00C8
    x"FC",x"FE",x"02",x"02",x"02",x"06",x"04",x"00", -- 0x00D0
    x"82",x"C6",x"6E",x"3C",x"18",x"FE",x"FE",x"00", -- 0x00D8
    x"02",x"02",x"02",x"02",x"FE",x"FE",x"00",x"00", -- 0x00E0
    x"FE",x"FE",x"70",x"38",x"70",x"FE",x"FE",x"00", -- 0x00E8
    x"FE",x"FE",x"1C",x"38",x"70",x"FE",x"FE",x"00", -- 0x00F0
    x"7C",x"FE",x"82",x"82",x"82",x"FE",x"7C",x"00", -- 0x00F8
    x"70",x"F8",x"88",x"88",x"88",x"FE",x"FE",x"00", -- 0x0100
    x"7A",x"FC",x"8E",x"8A",x"82",x"FE",x"7C",x"00", -- 0x0108
    x"72",x"F6",x"9E",x"8C",x"88",x"FE",x"FE",x"00", -- 0x0110
    x"0C",x"5E",x"D2",x"92",x"92",x"F6",x"64",x"00", -- 0x0118
    x"80",x"80",x"FE",x"FE",x"80",x"80",x"00",x"00", -- 0x0120
    x"FC",x"FE",x"02",x"02",x"02",x"FE",x"FC",x"00", -- 0x0128
    x"F0",x"F8",x"1C",x"0E",x"1C",x"F8",x"F0",x"00", -- 0x0130
    x"F8",x"FE",x"1C",x"38",x"1C",x"FE",x"F8",x"00", -- 0x0138
    x"C6",x"EE",x"7C",x"38",x"7C",x"EE",x"C6",x"00", -- 0x0140
    x"C0",x"F0",x"1E",x"1E",x"F0",x"C0",x"00",x"00", -- 0x0148
    x"C2",x"E2",x"F2",x"BA",x"9E",x"8E",x"86",x"00", -- 0x0150
    x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00", -- 0x0158
    x"00",x"02",x"07",x"02",x"00",x"00",x"00",x"00", -- 0x0160
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0168
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0170
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0178
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0180
    x"0F",x"1F",x"3F",x"3F",x"1F",x"1F",x"1F",x"03", -- 0x0188
    x"0F",x"07",x"03",x"01",x"00",x"01",x"01",x"03", -- 0x0190
    x"7F",x"7F",x"7F",x"7F",x"7F",x"3F",x"3F",x"1F", -- 0x0198
    x"1C",x"1C",x"3E",x"3E",x"3E",x"3E",x"7E",x"7F", -- 0x01A0
    x"00",x"00",x"00",x"00",x"00",x"0C",x"0C",x"1C", -- 0x01A8
    x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01B0
    x"07",x"01",x"00",x"03",x"03",x"03",x"01",x"01", -- 0x01B8
    x"FF",x"7F",x"3F",x"1F",x"1F",x"1F",x"0F",x"0F", -- 0x01C0
    x"00",x"80",x"E0",x"F0",x"6C",x"07",x"0F",x"A7", -- 0x01C8
    x"FF",x"FE",x"FE",x"3C",x"0C",x"00",x"00",x"00", -- 0x01D0
    x"03",x"0F",x"07",x"07",x"07",x"03",x"82",x"E3", -- 0x01D8
    x"00",x"00",x"00",x"00",x"00",x"04",x"0E",x"07", -- 0x01E0
    x"00",x"00",x"01",x"03",x"01",x"01",x"00",x"00", -- 0x01E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01F0
    x"FF",x"FF",x"FF",x"FF",x"F7",x"C3",x"81",x"00", -- 0x01F8
    x"00",x"00",x"00",x"00",x"00",x"03",x"0F",x"03", -- 0x0200
    x"3C",x"18",x"18",x"38",x"78",x"F8",x"F8",x"F8", -- 0x0208
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0210
    x"78",x"38",x"18",x"18",x"3C",x"00",x"00",x"00", -- 0x0218
    x"00",x"01",x"01",x"03",x"03",x"03",x"03",x"03", -- 0x0220
    x"00",x"00",x"00",x"80",x"80",x"80",x"80",x"80", -- 0x0228
    x"07",x"07",x"2F",x"3F",x"3F",x"3F",x"20",x"00", -- 0x0230
    x"C0",x"C0",x"E8",x"F8",x"F8",x"F8",x"08",x"00", -- 0x0238
    x"00",x"40",x"70",x"30",x"38",x"3C",x"1F",x"1F", -- 0x0240
    x"00",x"00",x"00",x"40",x"60",x"70",x"C0",x"80", -- 0x0248
    x"0F",x"0E",x"0E",x"0C",x"38",x"30",x"10",x"00", -- 0x0250
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0258
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0260
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0268
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0270
    x"18",x"18",x"78",x"9C",x"9C",x"78",x"18",x"18", -- 0x0278
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0280
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0288
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0290
    x"3F",x"0F",x"1E",x"44",x"44",x"1E",x"0F",x"3F", -- 0x0298
    x"01",x"02",x"04",x"09",x"11",x"23",x"47",x"8E", -- 0x02A0
    x"80",x"40",x"20",x"90",x"88",x"C4",x"E2",x"71", -- 0x02A8
    x"8E",x"47",x"23",x"11",x"09",x"04",x"02",x"01", -- 0x02B0
    x"71",x"E2",x"C4",x"88",x"90",x"20",x"40",x"80", -- 0x02B8
    x"00",x"00",x"07",x"1C",x"1B",x"32",x"2E",x"2C", -- 0x02C0
    x"00",x"00",x"E0",x"38",x"D8",x"4C",x"34",x"34", -- 0x02C8
    x"2C",x"2E",x"32",x"1B",x"1C",x"07",x"00",x"00", -- 0x02D0
    x"34",x"34",x"4C",x"D8",x"38",x"E0",x"00",x"00", -- 0x02D8
    x"FF",x"FF",x"FF",x"80",x"AF",x"A5",x"DB",x"81", -- 0x02E0
    x"80",x"60",x"B0",x"58",x"EC",x"76",x"3B",x"5D", -- 0x02E8
    x"9D",x"87",x"FF",x"FB",x"DB",x"C3",x"DE",x"F6", -- 0x02F0
    x"69",x"76",x"47",x"D6",x"A9",x"9F",x"B7",x"F7", -- 0x02F8
    x"03",x"06",x"0C",x"FC",x"CE",x"E7",x"71",x"3C", -- 0x0300
    x"C0",x"60",x"30",x"3F",x"73",x"E7",x"8E",x"3C", -- 0x0308
    x"3C",x"71",x"E7",x"CE",x"FC",x"0C",x"06",x"03", -- 0x0310
    x"3C",x"8E",x"E7",x"73",x"3E",x"30",x"60",x"C0", -- 0x0318
    x"0E",x"0E",x"07",x"07",x"03",x"03",x"07",x"01", -- 0x0320
    x"01",x"01",x"03",x"03",x"07",x"07",x"0E",x"0E", -- 0x0328
    x"FF",x"FF",x"70",x"7E",x"3A",x"3E",x"1C",x"1C", -- 0x0330
    x"1C",x"1C",x"3E",x"3A",x"7E",x"70",x"FF",x"FF", -- 0x0338
    x"E0",x"FC",x"FF",x"3F",x"07",x"00",x"00",x"00", -- 0x0340
    x"00",x"00",x"00",x"07",x"3F",x"FF",x"FC",x"E0", -- 0x0348
    x"03",x"1F",x"FF",x"FE",x"F0",x"E0",x"E0",x"E0", -- 0x0350
    x"E0",x"E0",x"E0",x"F0",x"FE",x"FF",x"1F",x"03", -- 0x0358
    x"E3",x"E1",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0", -- 0x0360
    x"E0",x"F0",x"F8",x"FC",x"FE",x"FF",x"EF",x"E7", -- 0x0368
    x"07",x"07",x"07",x"07",x"07",x"07",x"87",x"C7", -- 0x0370
    x"E7",x"F7",x"FF",x"7F",x"3F",x"1F",x"0F",x"07", -- 0x0378
    x"00",x"01",x"03",x"07",x"03",x"07",x"0F",x"3F", -- 0x0380
    x"80",x"80",x"D8",x"F8",x"F8",x"F0",x"F0",x"F0", -- 0x0388
    x"1F",x"1F",x"1F",x"0F",x"03",x"07",x"07",x"01", -- 0x0390
    x"F8",x"F8",x"F0",x"E0",x"F8",x"FC",x"78",x"00", -- 0x0398
    x"00",x"00",x"00",x"00",x"00",x"04",x"01",x"03", -- 0x03A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"40",x"90", -- 0x03A8
    x"07",x"02",x"02",x"08",x"00",x"00",x"00",x"00", -- 0x03B0
    x"C0",x"80",x"A0",x"10",x"00",x"00",x"00",x"00", -- 0x03B8
    x"00",x"00",x"00",x"04",x"24",x"04",x"4E",x"27", -- 0x03C0
    x"00",x"00",x"20",x"40",x"11",x"80",x"A4",x"C8", -- 0x03C8
    x"07",x"03",x"25",x"00",x"08",x"00",x"00",x"00", -- 0x03D0
    x"C0",x"20",x"90",x"A0",x"20",x"50",x"00",x"00", -- 0x03D8
    x"00",x"00",x"42",x"20",x"04",x"0F",x"E7",x"3F", -- 0x03E0
    x"00",x"20",x"44",x"C8",x"80",x"80",x"D0",x"EC", -- 0x03E8
    x"07",x"07",x"0D",x"1D",x"29",x"42",x"01",x"00", -- 0x03F0
    x"C0",x"A0",x"B0",x"88",x"44",x"20",x"10",x"08", -- 0x03F8
    x"00",x"00",x"00",x"00",x"80",x"80",x"C0",x"E1", -- 0x0400
    x"70",x"30",x"60",x"40",x"C0",x"00",x"00",x"00", -- 0x0408
    x"1F",x"07",x"01",x"00",x"00",x"00",x"00",x"00", -- 0x0410
    x"1F",x"1F",x"3F",x"3F",x"7F",x"7F",x"FF",x"FF", -- 0x0418
    x"00",x"00",x"00",x"00",x"00",x"00",x"03",x"0F", -- 0x0420
    x"FF",x"7F",x"07",x"00",x"00",x"00",x"00",x"00", -- 0x0428
    x"FF",x"FF",x"FF",x"F8",x"00",x"00",x"00",x"00", -- 0x0430
    x"03",x"07",x"07",x"0F",x"1F",x"FF",x"FF",x"FF", -- 0x0438
    x"FF",x"FF",x"FF",x"7F",x"1F",x"0F",x"07",x"03", -- 0x0440
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0448
    x"00",x"00",x"00",x"00",x"00",x"02",x"03",x"01", -- 0x0450
    x"C0",x"60",x"60",x"30",x"30",x"30",x"18",x"18", -- 0x0458
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"80", -- 0x0460
    x"03",x"03",x"01",x"01",x"01",x"00",x"00",x"00", -- 0x0468
    x"00",x"C0",x"50",x"34",x"1A",x"0D",x"06",x"06", -- 0x0470
    x"40",x"40",x"A0",x"A0",x"A0",x"D0",x"D0",x"D0", -- 0x0478
    x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"80", -- 0x0480
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0488
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0490
    x"FF",x"FF",x"FE",x"FE",x"FE",x"FC",x"FC",x"FC", -- 0x0498
    x"F8",x"F8",x"F8",x"F8",x"F0",x"F0",x"F0",x"F0", -- 0x04A0
    x"E0",x"E0",x"C0",x"C0",x"C0",x"80",x"80",x"80", -- 0x04A8
    x"FF",x"FF",x"FF",x"FE",x"FE",x"FC",x"FC",x"F8", -- 0x04B0
    x"F8",x"F8",x"F0",x"F0",x"E0",x"E0",x"C0",x"C0", -- 0x04B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x04C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"FE",x"FC", -- 0x04C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"FE",x"FC", -- 0x04D0
    x"FC",x"F8",x"F8",x"F0",x"E0",x"C0",x"C0",x"80", -- 0x04D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x04E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x04E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x04F0
    x"C0",x"80",x"80",x"00",x"00",x"00",x"00",x"00", -- 0x04F8
    x"FC",x"F8",x"F8",x"F0",x"F0",x"E0",x"E0",x"E0", -- 0x0500
    x"80",x"80",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0508
    x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"00", -- 0x0510
    x"33",x"3F",x"1F",x"00",x"00",x"00",x"00",x"00", -- 0x0518
    x"C0",x"80",x"80",x"00",x"00",x"00",x"00",x"00", -- 0x0520
    x"C0",x"40",x"40",x"40",x"60",x"60",x"40",x"C0", -- 0x0528
    x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"C0", -- 0x0530
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0538
    x"0F",x"38",x"E0",x"C0",x"80",x"00",x"00",x"00", -- 0x0540
    x"00",x"00",x"00",x"00",x"00",x"00",x"06",x"07", -- 0x0548
    x"C0",x"C0",x"C0",x"C0",x"C0",x"80",x"80",x"00", -- 0x0550
    x"E0",x"E0",x"40",x"00",x"00",x"00",x"00",x"00", -- 0x0558
    x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF", -- 0x0560
    x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00", -- 0x0568
    x"F0",x"F8",x"FC",x"FE",x"1F",x"0F",x"07",x"07", -- 0x0570
    x"07",x"07",x"0F",x"1F",x"FE",x"FC",x"F8",x"F0", -- 0x0578
    x"E1",x"E1",x"E1",x"E1",x"FF",x"FF",x"FF",x"FF", -- 0x0580
    x"1E",x"3F",x"7F",x"FF",x"F3",x"E1",x"E1",x"E1", -- 0x0588
    x"07",x"0F",x"9F",x"FF",x"FC",x"F8",x"F0",x"E0", -- 0x0590
    x"C0",x"C0",x"C0",x"C0",x"FF",x"FF",x"FF",x"FF", -- 0x0598
    x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF", -- 0x05A0
    x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05A8
    x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"01",x"07", -- 0x05B0
    x"1F",x"7F",x"FE",x"F8",x"FF",x"FF",x"FF",x"FF", -- 0x05B8
    x"FF",x"FF",x"FF",x"FF",x"1F",x"7F",x"FE",x"F8", -- 0x05C0
    x"E0",x"80",x"00",x"00",x"FF",x"FF",x"FF",x"FF", -- 0x05C8
    x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"FF", -- 0x05D0
    x"FF",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0", -- 0x05D8
    x"38",x"78",x"F8",x"F8",x"F0",x"E0",x"E0",x"E0", -- 0x05E0
    x"E0",x"E0",x"E0",x"F0",x"FF",x"FF",x"7F",x"3F", -- 0x05E8
    x"1C",x"1E",x"1F",x"1F",x"0F",x"07",x"07",x"07", -- 0x05F0
    x"07",x"07",x"07",x"0F",x"FF",x"FF",x"FE",x"FC", -- 0x05F8
    x"80",x"C0",x"E0",x"F0",x"F8",x"7C",x"3E",x"1F", -- 0x0600
    x"0F",x"07",x"03",x"03",x"FF",x"FF",x"FF",x"FF", -- 0x0608
    x"01",x"03",x"07",x"0F",x"1F",x"3E",x"7C",x"F8", -- 0x0610
    x"F0",x"E0",x"C0",x"C0",x"FF",x"FF",x"FF",x"FF", -- 0x0618
    x"00",x"00",x"C3",x"2C",x"10",x"11",x"00",x"00", -- 0x0620
    x"00",x"00",x"00",x"80",x"40",x"20",x"10",x"10", -- 0x0628
    x"00",x"FE",x"FF",x"FE",x"70",x"E0",x"FC",x"F0", -- 0x0630
    x"08",x"08",x"14",x"14",x"28",x"48",x"10",x"20", -- 0x0638
    x"00",x"00",x"00",x"04",x"06",x"0F",x"0C",x"08", -- 0x0640
    x"00",x"00",x"00",x"00",x"67",x"06",x"06",x"01", -- 0x0648
    x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00", -- 0x0650
    x"20",x"20",x"60",x"58",x"B8",x"50",x"00",x"00", -- 0x0658
    x"F0",x"E7",x"FF",x"DE",x"D0",x"C6",x"FD",x"F7", -- 0x0660
    x"C7",x"D7",x"7F",x"00",x"DC",x"70",x"C0",x"00", -- 0x0668
    x"DF",x"FF",x"FD",x"F9",x"F5",x"ED",x"C7",x"A7", -- 0x0670
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0678
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0680
    x"00",x"00",x"00",x"00",x"18",x"0D",x"02",x"04", -- 0x0688
    x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"02", -- 0x0690
    x"62",x"27",x"10",x"E6",x"92",x"0C",x"68",x"20", -- 0x0698
    x"00",x"00",x"00",x"00",x"00",x"C0",x"61",x"13", -- 0x06A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x06A8
    x"12",x"04",x"F1",x"52",x"31",x"36",x"05",x"04", -- 0x06B0
    x"C0",x"20",x"A0",x"20",x"20",x"40",x"40",x"80", -- 0x06B8
    x"05",x"04",x"02",x"01",x"00",x"01",x"01",x"01", -- 0x06C0
    x"C0",x"40",x"40",x"40",x"C0",x"C0",x"FC",x"8A", -- 0x06C8
    x"01",x"06",x"08",x"00",x"00",x"00",x"00",x"00", -- 0x06D0
    x"72",x"01",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x06D8
    x"00",x"00",x"00",x"00",x"00",x"08",x"0C",x"02", -- 0x06E0
    x"00",x"78",x"20",x"20",x"10",x"10",x"20",x"20", -- 0x06E8
    x"13",x"0F",x"E3",x"00",x"00",x"00",x"00",x"00", -- 0x06F0
    x"70",x"D0",x"10",x"0C",x"04",x"00",x"00",x"00", -- 0x06F8
    x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"03", -- 0x0700
    x"00",x"00",x"00",x"10",x"7C",x"FF",x"FF",x"DF", -- 0x0708
    x"03",x"07",x"07",x"09",x"0F",x"0F",x"05",x"0D", -- 0x0710
    x"37",x"8F",x"C7",x"82",x"01",x"87",x"E1",x"F9", -- 0x0718
    x"00",x"00",x"00",x"00",x"00",x"0F",x"9F",x"FF", -- 0x0720
    x"00",x"00",x"00",x"00",x"00",x"40",x"B8",x"78", -- 0x0728
    x"9C",x"2F",x"74",x"F8",x"F1",x"A7",x"0F",x"CF", -- 0x0730
    x"70",x"60",x"F0",x"E0",x"E0",x"C0",x"C0",x"E0", -- 0x0738
    x"0E",x"07",x"07",x"0B",x"07",x"03",x"01",x"01", -- 0x0740
    x"FF",x"7F",x"EF",x"F6",x"74",x"8F",x"8B",x"8E", -- 0x0748
    x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0750
    x"DF",x"77",x"23",x"03",x"03",x"03",x"00",x"00", -- 0x0758
    x"EF",x"EF",x"7F",x"2F",x"8F",x"9F",x"3F",x"7E", -- 0x0760
    x"E0",x"D0",x"F0",x"F0",x"E0",x"E0",x"80",x"10", -- 0x0768
    x"6E",x"3E",x"DC",x"F8",x"F8",x"30",x"00",x"00", -- 0x0770
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0778
    x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00", -- 0x0780
    x"00",x"00",x"00",x"00",x"00",x"94",x"F7",x"33", -- 0x0788
    x"00",x"01",x"00",x"00",x"00",x"03",x"02",x"00", -- 0x0790
    x"1A",x"8E",x"C8",x"FA",x"D6",x"33",x"7D",x"FF", -- 0x0798
    x"00",x"00",x"00",x"00",x"00",x"02",x"14",x"35", -- 0x07A0
    x"00",x"00",x"00",x"00",x"00",x"40",x"80",x"00", -- 0x07A8
    x"24",x"28",x"49",x"DF",x"D7",x"77",x"CE",x"F8", -- 0x07B0
    x"00",x"00",x"00",x"00",x"80",x"80",x"20",x"00", -- 0x07B8
    x"01",x"00",x"00",x"01",x"00",x"01",x"00",x"00", -- 0x07C0
    x"87",x"FB",x"8E",x"19",x"F7",x"63",x"42",x"9C", -- 0x07C8
    x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07D0
    x"66",x"82",x"01",x"01",x"00",x"00",x"00",x"00", -- 0x07D8
    x"FF",x"FF",x"F8",x"EA",x"AE",x"79",x"DC",x"4A", -- 0x07E0
    x"C0",x"80",x"40",x"00",x"00",x"00",x"80",x"00", -- 0x07E8
    x"40",x"70",x"58",x"08",x"00",x"00",x"00",x"00", -- 0x07F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"  -- 0x07F8
  );

begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
