library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity journey_bg_bits_1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of journey_bg_bits_1 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"15",X"BC",X"15",X"AC",X"15",X"AC",X"15",X"AB",X"15",X"FF",X"D5",X"FF",X"D5",X"55",X"D5",
		X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"15",X"C0",X"15",X"C0",X"15",X"F0",X"15",
		X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"15",
		X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"15",X"00",X"15",
		X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"5F",X"FF",X"57",X"FF",X"7F",X"FD",
		X"FD",X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",X"FF",
		X"D7",X"DF",X"DF",X"DF",X"DF",X"FF",X"FF",X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",X"FF",
		X"FA",X"AA",X"FA",X"AA",X"FA",X"AA",X"FA",X"AA",X"FA",X"AB",X"FA",X"BF",X"FA",X"FF",X"FF",X"D5",
		X"FA",X"B0",X"FA",X"BC",X"FA",X"BC",X"FA",X"AF",X"FA",X"AF",X"FA",X"AB",X"FA",X"AB",X"FA",X"AA",
		X"B0",X"00",X"BC",X"00",X"BC",X"00",X"BF",X"00",X"BF",X"00",X"BF",X"C0",X"FA",X"C0",X"FA",X"F0",
		X"F0",X"00",X"C0",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"B0",X"00",
		X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",
		X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",
		X"F1",X"D5",X"F1",X"50",X"F1",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",
		X"F1",X"DD",X"F1",X"DD",X"F1",X"DD",X"F1",X"DD",X"F1",X"DD",X"F1",X"DD",X"F1",X"D5",X"F1",X"D5",
		X"AA",X"FF",X"A7",X"FF",X"BF",X"FF",X"FD",X"FF",X"7F",X"FF",X"FF",X"DF",X"FF",X"57",X"F5",X"55",
		X"FE",X"AA",X"FA",X"AA",X"EA",X"AB",X"6A",X"AB",X"AA",X"AF",X"AA",X"AF",X"AA",X"BF",X"AA",X"BF",
		X"55",X"AA",X"75",X"AA",X"F5",X"AA",X"F5",X"AA",X"F5",X"AA",X"D5",X"AA",X"56",X"AA",X"56",X"AA",
		X"F7",X"FF",X"55",X"FF",X"55",X"AA",X"01",X"AA",X"01",X"AA",X"01",X"AA",X"05",X"AA",X"15",X"AA",
		X"F5",X"57",X"FD",X"55",X"FD",X"55",X"FD",X"55",X"FD",X"57",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"5F",X"FF",X"57",X"FF",X"57",X"FF",X"55",X"FF",X"D5",X"7F",X"D5",X"7F",X"F5",X"5F",X"F5",X"5F",
		X"FF",X"FD",X"FF",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"7F",X"FF",X"5F",X"FF",
		X"DF",X"7D",X"DF",X"7D",X"FF",X"7D",X"FF",X"7D",X"FF",X"7D",X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",
		X"DF",X"7D",X"DF",X"7D",X"DF",X"7D",X"DF",X"7D",X"DF",X"7D",X"DF",X"7D",X"DF",X"7D",X"DF",X"7D",
		X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"55",X"4F",X"55",X"0D",X"00",X"0D",X"00",X"3D",X"C0",X"7D",
		X"FD",X"DA",X"7F",X"FA",X"7F",X"FE",X"7F",X"DF",X"5F",X"FD",X"D7",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F5",X"FF",X"D7",X"FF",X"1F",X"FF",X"0F",X"55",X"0D",X"55",X"05",X"7E",X"F5",X"FA",X"F5",X"DA",
		X"00",X"00",X"00",X"01",X"00",X"05",X"01",X"55",X"55",X"55",X"FF",X"FF",X"FF",X"55",X"FD",X"55",
		X"FF",X"FF",X"FF",X"FF",X"5F",X"F5",X"55",X"55",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"FF",X"AB",X"FF",X"AF",X"FF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FD",X"FF",X"A9",X"FF",X"A9",X"FE",X"AF",X"FA",X"AF",X"EA",X"BF",X"AA",X"BF",
		X"FD",X"5F",X"FD",X"57",X"FF",X"57",X"FF",X"D5",X"FF",X"D5",X"FF",X"F5",X"FF",X"F5",X"FF",X"F5",
		X"57",X"FF",X"57",X"FF",X"D7",X"FF",X"15",X"FF",X"15",X"FF",X"D5",X"7F",X"F5",X"7F",X"FD",X"5F",
		X"FF",X"F7",X"FF",X"F7",X"FF",X"F7",X"FF",X"F7",X"7F",X"F7",X"7F",X"FF",X"5F",X"FF",X"5F",X"FF",
		X"7D",X"47",X"FD",X"05",X"FD",X"05",X"FD",X"01",X"FD",X"C0",X"FD",X"F0",X"FD",X"F4",X"FD",X"F7",
		X"FF",X"FF",X"FF",X"FD",X"FF",X"F5",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AF",X"55",X"AF",X"55",X"AF",X"55",X"A5",X"55",X"57",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"03",X"00",X"00",X"00",X"00",X"2F",X"00",X"AF",X"C0",X"AF",X"FC",X"AF",X"FF",X"AF",X"D5",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"FF",X"FF",X"C0",X"3F",X"00",X"0F",
		X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"D5",X"FD",X"55",X"55",X"50",X"50",X"00",X"00",X"00",
		X"FF",X"FA",X"FF",X"EA",X"FF",X"AA",X"FA",X"AA",X"EA",X"AA",X"AA",X"AA",X"AA",X"BF",X"AB",X"FF",
		X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"0F",
		X"00",X"D7",X"00",X"17",X"00",X"15",X"00",X"15",X"00",X"05",X"00",X"0D",X"00",X"01",X"00",X"01",
		X"01",X"FF",X"01",X"FF",X"01",X"7F",X"01",X"7F",X"01",X"7F",X"03",X"5F",X"00",X"5F",X"00",X"5F",
		X"FF",X"FF",X"0F",X"FF",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"0A",X"AA",X"28",X"02",X"20",X"02",X"20",X"02",X"20",X"02",X"22",X"AA",X"22",X"AA",X"00",X"00",
		X"00",X"00",X"00",X"02",X"2A",X"AA",X"2A",X"AA",X"20",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"22",X"82",X"22",X"82",X"20",X"82",X"20",X"82",X"20",X"82",X"20",X"AA",X"20",X"AA",X"00",X"00",
		X"22",X"AA",X"20",X"82",X"20",X"82",X"20",X"82",X"20",X"02",X"20",X"0A",X"20",X"0A",X"00",X"00",
		X"00",X"80",X"2A",X"AA",X"00",X"80",X"00",X"80",X"00",X"80",X"0A",X"80",X"0A",X"80",X"00",X"00",
		X"20",X"AA",X"20",X"82",X"20",X"82",X"20",X"82",X"20",X"82",X"22",X"8A",X"22",X"8A",X"00",X"00",
		X"20",X"AA",X"20",X"82",X"20",X"82",X"20",X"82",X"20",X"82",X"22",X"AA",X"22",X"AA",X"00",X"00",
		X"28",X"00",X"22",X"00",X"22",X"80",X"20",X"AA",X"20",X"2A",X"20",X"00",X"20",X"00",X"00",X"00",
		X"2A",X"AA",X"20",X"82",X"20",X"82",X"20",X"82",X"20",X"82",X"22",X"AA",X"22",X"AA",X"00",X"00",
		X"2A",X"AA",X"2A",X"AA",X"20",X"80",X"20",X"80",X"20",X"80",X"20",X"80",X"22",X"80",X"00",X"00",
		X"FF",X"F5",X"FF",X"F5",X"FF",X"F5",X"FF",X"F5",X"FF",X"F5",X"FF",X"F5",X"FF",X"F7",X"FF",X"CF",
		X"F5",X"40",X"F4",X"00",X"F0",X"00",X"C0",X"00",X"00",X"01",X"00",X"15",X"03",X"D5",X"0F",X"D5",
		X"55",X"44",X"55",X"50",X"D5",X"40",X"D5",X"40",X"D5",X"55",X"F5",X"5F",X"F5",X"5F",X"F5",X"5C",
		X"AA",X"AA",X"AA",X"AB",X"AA",X"BF",X"AF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"D5",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FE",X"AA",X"EA",X"AA",
		X"00",X"3F",X"0F",X"FF",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"57",X"FF",X"55",X"7F",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"2A",X"AA",X"2A",X"AA",X"20",X"80",X"20",X"80",X"20",X"80",X"22",X"AA",X"22",X"AA",X"00",X"00",
		X"2A",X"2A",X"22",X"A2",X"20",X"82",X"20",X"82",X"20",X"82",X"22",X"AA",X"22",X"AA",X"00",X"00",
		X"20",X"0A",X"20",X"0A",X"20",X"0A",X"20",X"0A",X"20",X"0A",X"22",X"AA",X"22",X"A8",X"00",X"00",
		X"0A",X"A8",X"28",X"0A",X"20",X"02",X"20",X"02",X"20",X"02",X"22",X"AA",X"22",X"AA",X"00",X"00",
		X"20",X"02",X"20",X"02",X"20",X"82",X"20",X"82",X"20",X"82",X"22",X"AA",X"22",X"AA",X"00",X"00",
		X"20",X"00",X"20",X"00",X"20",X"80",X"20",X"80",X"20",X"80",X"22",X"AA",X"22",X"AA",X"00",X"00",
		X"20",X"AA",X"20",X"82",X"20",X"82",X"20",X"02",X"20",X"02",X"22",X"AA",X"22",X"A8",X"00",X"00",
		X"2A",X"AA",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"0A",X"AA",X"0A",X"AA",X"00",X"00",
		X"00",X"00",X"00",X"00",X"20",X"02",X"2A",X"AA",X"2A",X"AA",X"20",X"02",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0A",X"AA",X"0A",X"AA",X"00",X"02",X"00",X"02",X"00",X"0A",X"00",X"0A",X"00",X"00",
		X"28",X"02",X"0A",X"0A",X"02",X"A8",X"00",X"A0",X"00",X"20",X"0A",X"AA",X"0A",X"AA",X"00",X"00",
		X"00",X"0A",X"00",X"0A",X"00",X"02",X"00",X"02",X"00",X"02",X"0A",X"AA",X"0A",X"AA",X"00",X"00",
		X"2A",X"AA",X"0A",X"00",X"02",X"A0",X"02",X"A0",X"0A",X"00",X"2A",X"AA",X"2A",X"AA",X"00",X"00",
		X"2A",X"AA",X"00",X"2A",X"02",X"A0",X"2A",X"00",X"20",X"00",X"22",X"AA",X"22",X"AA",X"00",X"00",
		X"2A",X"AA",X"20",X"02",X"20",X"02",X"20",X"02",X"20",X"02",X"22",X"AA",X"22",X"AA",X"00",X"00",
		X"2A",X"80",X"20",X"80",X"20",X"80",X"20",X"80",X"20",X"80",X"22",X"AA",X"22",X"AA",X"00",X"00",
		X"2A",X"AA",X"20",X"28",X"20",X"2A",X"20",X"02",X"20",X"02",X"22",X"AA",X"22",X"AA",X"00",X"00",
		X"2A",X"8A",X"20",X"AA",X"20",X"A0",X"20",X"80",X"20",X"80",X"22",X"AA",X"22",X"AA",X"00",X"00",
		X"20",X"AA",X"20",X"AA",X"20",X"82",X"20",X"82",X"20",X"82",X"22",X"8A",X"22",X"8A",X"00",X"00",
		X"00",X"00",X"20",X"00",X"20",X"00",X"2A",X"AA",X"2A",X"AA",X"20",X"00",X"20",X"00",X"00",X"00",
		X"2A",X"AA",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"0A",X"AA",X"0A",X"AA",X"00",X"00",
		X"2A",X"A0",X"00",X"28",X"00",X"0A",X"00",X"2A",X"00",X"A8",X"0A",X"A0",X"0A",X"80",X"00",X"00",
		X"2A",X"AA",X"00",X"28",X"02",X"A0",X"02",X"A0",X"00",X"28",X"0A",X"AA",X"0A",X"AA",X"00",X"00",
		X"28",X"0A",X"0A",X"28",X"02",X"A0",X"00",X"80",X"02",X"A0",X"0A",X"28",X"00",X"0A",X"00",X"00",
		X"28",X"00",X"0A",X"00",X"02",X"80",X"00",X"AA",X"02",X"AA",X"0A",X"80",X"0A",X"00",X"00",X"00",
		X"20",X"02",X"22",X"02",X"22",X"82",X"20",X"82",X"20",X"A2",X"20",X"2A",X"20",X"0A",X"00",X"00",
		X"FC",X"00",X"F0",X"0F",X"C0",X"3F",X"00",X"FF",X"0F",X"FF",X"1F",X"FF",X"5F",X"FF",X"5F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"FF",X"C0",X"FF",X"00",
		X"FF",X"55",X"55",X"55",X"55",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"EA",X"FA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"BF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"54",X"00",X"50",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"50",X"55",X"50",X"55",X"50",X"55",X"50",X"55",X"50",X"55",X"40",X"55",X"40",X"55",X"00",
		X"00",X"00",X"00",X"00",X"55",X"00",X"55",X"40",X"55",X"40",X"55",X"50",X"55",X"50",X"55",X"50",
		X"FF",X"F0",X"FF",X"F0",X"FF",X"F0",X"FF",X"F0",X"FF",X"F0",X"FF",X"C0",X"3F",X"C0",X"03",X"C0",
		X"FF",X"01",X"FF",X"D5",X"FF",X"D5",X"FD",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FF",X"F0",X"FF",X"C0",X"FF",X"C1",
		X"FF",X"FF",X"FF",X"FD",X"FD",X"55",X"55",X"57",X"57",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AB",X"FF",
		X"FE",X"00",X"FA",X"00",X"F8",X"00",X"E8",X"00",X"A0",X"00",X"80",X"00",X"00",X"0F",X"FF",X"FF",
		X"BF",X"F9",X"BF",X"F9",X"BF",X"E9",X"EF",X"E5",X"FF",X"E4",X"FF",X"A0",X"FF",X"80",X"FE",X"80",
		X"FE",X"95",X"FF",X"95",X"FF",X"95",X"BF",X"A5",X"BF",X"E5",X"BF",X"E5",X"BF",X"E5",X"BF",X"E9",
		X"00",X"00",X"00",X"00",X"95",X"55",X"A5",X"55",X"E9",X"55",X"F9",X"55",X"FA",X"55",X"FE",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",X"00",X"00",
		X"55",X"FF",X"55",X"7F",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"5F",X"FF",X"57",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"D5",X"55",X"55",X"55",X"55",X"5F",X"5F",X"FF",X"5F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FE",X"FF",X"FF",
		X"FE",X"FE",X"BF",X"FA",X"BF",X"EA",X"AA",X"AA",X"AA",X"AB",X"FA",X"AF",X"BF",X"FF",X"BF",X"FF",
		X"EA",X"AF",X"AA",X"AB",X"AF",X"EA",X"BF",X"FA",X"BF",X"FE",X"BE",X"FE",X"FB",X"BE",X"FB",X"BE",
		X"FF",X"FA",X"FF",X"FE",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",
		X"FD",X"55",X"D5",X"55",X"55",X"7F",X"55",X"FF",X"57",X"FF",X"57",X"FF",X"57",X"FF",X"55",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"AA",
		X"3F",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"03",X"FF",X"03",X"FF",X"03",X"FF",X"0F",X"FF",X"0F",X"FE",X"0F",X"FE",X"3F",X"FE",X"3F",X"FE",
		X"00",X"0F",X"00",X"0F",X"00",X"3F",X"00",X"3F",X"00",X"3F",X"00",X"3F",X"00",X"FF",X"00",X"FF",
		X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"D5",X"F5",X"55",X"D5",X"55",X"55",X"7F",X"FF",X"F5",
		X"BF",X"FF",X"BF",X"FF",X"AB",X"FF",X"AA",X"FF",X"AA",X"BF",X"AA",X"AF",X"AA",X"AA",X"AA",X"AA",
		X"00",X"3F",X"00",X"FF",X"03",X"FF",X"0F",X"FF",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"03",X"00",X"0F",X"00",X"0F",X"00",X"3F",
		X"15",X"40",X"55",X"40",X"55",X"40",X"55",X"00",X"55",X"00",X"54",X"00",X"54",X"00",X"54",X"00",
		X"00",X"54",X"01",X"54",X"01",X"50",X"01",X"50",X"01",X"50",X"01",X"50",X"05",X"50",X"15",X"50",
		X"FF",X"FF",X"55",X"5F",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"F5",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"FF",X"03",X"FF",X"2B",X"FF",X"2A",X"FF",X"AA",X"BF",X"AA",X"AF",X"AA",X"AB",X"AA",X"AA",
		X"55",X"40",X"55",X"00",X"54",X"00",X"50",X"00",X"40",X"00",X"00",X"00",X"00",X"03",X"00",X"0F",
		X"40",X"00",X"50",X"00",X"50",X"00",X"55",X"00",X"55",X"00",X"55",X"40",X"55",X"50",X"55",X"54",
		X"01",X"55",X"00",X"55",X"00",X"55",X"00",X"15",X"00",X"15",X"00",X"05",X"00",X"01",X"00",X"00",
		X"15",X"40",X"15",X"40",X"15",X"50",X"05",X"50",X"05",X"50",X"05",X"54",X"05",X"54",X"01",X"55",
		X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"15",X"00",
		X"FF",X"FF",X"FF",X"FF",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FA",X"AA",X"AA",
		X"15",X"55",X"05",X"55",X"00",X"55",X"00",X"15",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"01",X"40",X"00",X"50",X"00",X"54",X"00",X"55",X"00",X"55",X"40",X"55",X"50",X"55",X"55",
		X"15",X"56",X"05",X"55",X"05",X"55",X"01",X"55",X"01",X"55",X"00",X"55",X"00",X"15",X"00",X"05",
		X"55",X"6A",X"55",X"6A",X"55",X"6A",X"55",X"6A",X"55",X"6A",X"15",X"6A",X"15",X"5A",X"15",X"5A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"05",X"55",X"00",X"00",X"00",X"00",
		X"55",X"55",X"15",X"55",X"01",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"FF",X"AA",X"AA",X"6A",X"AA",X"5A",X"AA",X"55",X"AA",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FA",X"FF",X"FA",X"FF",X"FE",X"BF",X"FE",X"BF",X"BF",X"AF",X"BF",X"AA",X"AF",X"EA",X"AB",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"57",X"FF",X"55",X"7F",
		X"FA",X"AA",X"FF",X"AA",X"FF",X"FA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"55",X"55",X"55",X"05",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"5F",X"FF",X"55",X"FF",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"EA",X"AA",X"FE",X"AA",X"FF",X"AA",X"FF",X"EA",X"FF",X"FA",X"FF",X"FF",
		X"01",X"55",X"00",X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"AA",X"00",X"AA",X"A0",
		X"40",X"00",X"50",X"00",X"55",X"00",X"55",X"54",X"55",X"55",X"55",X"55",X"55",X"55",X"15",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"57",X"FF",X"55",X"FF",X"55",X"7F",
		X"FF",X"FA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"A8",X"00",X"AA",X"00",X"AA",X"A0",X"EA",X"A8",X"FA",X"AA",X"FE",X"AA",X"FF",X"AA",X"FF",X"EA",
		X"55",X"55",X"15",X"55",X"05",X"55",X"01",X"55",X"00",X"55",X"00",X"15",X"00",X"01",X"A0",X"00",
		X"55",X"7F",X"55",X"5F",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"7F",X"FF",X"5F",X"FF",X"5F",X"FF",X"55",X"FF",X"55",X"7F",
		X"E8",X"00",X"EA",X"00",X"FA",X"80",X"FA",X"A0",X"FE",X"A0",X"FF",X"A8",X"FF",X"AA",X"FF",X"EA",
		X"01",X"55",X"01",X"55",X"00",X"55",X"00",X"55",X"80",X"15",X"80",X"05",X"A0",X"05",X"A0",X"01",
		X"55",X"40",X"55",X"40",X"55",X"50",X"55",X"50",X"55",X"54",X"15",X"54",X"15",X"55",X"05",X"55",
		X"50",X"00",X"50",X"00",X"54",X"00",X"54",X"00",X"54",X"00",X"55",X"00",X"55",X"00",X"55",X"40",
		X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"00",
		X"57",X"FF",X"57",X"FF",X"55",X"FF",X"55",X"FF",X"55",X"7F",X"55",X"7F",X"55",X"5F",X"55",X"5F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"7F",X"FF",X"7F",X"FF",X"5F",X"FF",
		X"FF",X"F8",X"FF",X"F8",X"FF",X"FA",X"FF",X"FA",X"FF",X"FE",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"81",X"FF",X"81",X"FF",X"E1",X"FF",X"E0",X"FF",X"E0",X"FF",X"E0",X"FF",X"E0",X"FF",X"E8",
		X"FC",X"15",X"FF",X"15",X"FF",X"15",X"FF",X"15",X"FF",X"05",X"FF",X"85",X"FF",X"85",X"FF",X"81",
		X"F0",X"15",X"FC",X"15",X"FC",X"15",X"FC",X"15",X"FC",X"15",X"FC",X"15",X"FC",X"15",X"FC",X"15",
		X"55",X"57",X"55",X"57",X"55",X"57",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"7F",X"55",X"7F",X"55",X"7F",X"55",X"7F",X"55",X"5F",X"55",X"5F",X"55",X"5F",X"55",X"5F",
		X"55",X"FF",X"55",X"FF",X"55",X"FF",X"55",X"FF",X"55",X"FF",X"55",X"FF",X"55",X"7F",X"55",X"7F",
		X"57",X"FF",X"57",X"FF",X"57",X"FF",X"57",X"FF",X"57",X"FF",X"57",X"FF",X"57",X"FF",X"57",X"FF",
		X"5F",X"FF",X"5F",X"FF",X"5F",X"FF",X"5F",X"FF",X"5F",X"FF",X"5F",X"FF",X"5F",X"FF",X"5F",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"2A",X"A8",X"A0",X"0A",X"88",X"22",X"88",X"22",X"88",X"22",X"8A",X"A2",X"A0",X"0A",X"2A",X"A8",
		X"5A",X"AA",X"DA",X"AA",X"DA",X"AA",X"DA",X"AA",X"FA",X"AA",X"FA",X"AA",X"FA",X"EA",X"FA",X"AA",
		X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",
		X"6A",X"AA",X"6A",X"AA",X"6A",X"AA",X"6A",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",
		X"6A",X"AA",X"6A",X"AA",X"6A",X"AA",X"6A",X"AA",X"6A",X"AA",X"6A",X"AA",X"6A",X"AA",X"6A",X"AA",
		X"FF",X"F5",X"FF",X"F5",X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"55",X"FF",X"55",X"FF",X"55",X"FF",X"D5",X"FF",X"D5",X"FF",X"D5",X"FF",X"D5",X"FF",X"F5",
		X"F5",X"55",X"F5",X"55",X"F5",X"55",X"F5",X"55",X"FD",X"55",X"FD",X"55",X"FD",X"55",X"FD",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",
		X"FF",X"D5",X"FF",X"D5",X"FF",X"D5",X"FF",X"D5",X"FF",X"D5",X"FF",X"D5",X"FF",X"D5",X"FF",X"D5",
		X"FF",X"55",X"FF",X"55",X"FF",X"55",X"FF",X"55",X"FF",X"55",X"FF",X"55",X"FF",X"55",X"FF",X"55",
		X"FD",X"55",X"FD",X"55",X"FD",X"55",X"FD",X"55",X"FD",X"55",X"FD",X"55",X"FD",X"55",X"FD",X"55",
		X"FF",X"15",X"FF",X"D5",X"FF",X"D5",X"FF",X"55",X"FF",X"55",X"FF",X"55",X"FF",X"55",X"FF",X"55",
		X"FF",X"F5",X"FF",X"F5",X"FF",X"F5",X"FF",X"D5",X"FF",X"D5",X"FF",X"D5",X"FF",X"D5",X"FF",X"D5",
		X"F5",X"55",X"F5",X"55",X"F5",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",
		X"55",X"55",X"55",X"56",X"55",X"5A",X"55",X"6A",X"55",X"6A",X"55",X"AA",X"55",X"AA",X"56",X"AA",
		X"56",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"6A",X"AA",X"6A",X"AA",
		X"55",X"6A",X"55",X"6A",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"56",X"AA",X"56",X"AA",
		X"55",X"5A",X"55",X"5A",X"55",X"5A",X"55",X"6A",X"55",X"6A",X"55",X"6A",X"55",X"6A",X"55",X"6A",
		X"55",X"56",X"55",X"56",X"55",X"5A",X"55",X"5A",X"55",X"5A",X"55",X"5A",X"55",X"5A",X"55",X"5A",
		X"55",X"56",X"55",X"56",X"55",X"56",X"55",X"56",X"55",X"56",X"55",X"56",X"55",X"56",X"55",X"56",
		X"55",X"55",X"59",X"55",X"59",X"55",X"59",X"55",X"59",X"55",X"59",X"55",X"59",X"55",X"59",X"55",
		X"AA",X"55",X"AA",X"95",X"AA",X"95",X"AA",X"95",X"AA",X"95",X"AA",X"95",X"AA",X"95",X"AA",X"A6",
		X"95",X"56",X"95",X"56",X"95",X"56",X"95",X"5A",X"95",X"5A",X"94",X"5A",X"95",X"5A",X"95",X"5A",
		X"95",X"6A",X"95",X"6A",X"95",X"6A",X"95",X"6A",X"95",X"6A",X"95",X"6A",X"95",X"6A",X"95",X"6A",
		X"95",X"AA",X"95",X"AA",X"95",X"AA",X"95",X"AA",X"95",X"AA",X"95",X"AA",X"95",X"AA",X"95",X"AA",
		X"96",X"AA",X"96",X"AA",X"A6",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"C0",X"00",X"F0",X"00",X"FC",X"00",X"F0",X"00",X"FF",X"00",X"FF",X"C0",X"FF",X"FF",
		X"00",X"03",X"00",X"0F",X"00",X"3F",X"00",X"0F",X"03",X"CF",X"0F",X"FF",X"3F",X"FF",X"FF",X"FF",
		X"55",X"55",X"85",X"55",X"00",X"55",X"0C",X"95",X"00",X"05",X"00",X"C1",X"00",X"01",X"00",X"00",
		X"D5",X"F7",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"57",X"55",X"5F",X"55",X"7F",X"55",X"FF",X"55",X"7F",X"55",X"7F",X"57",X"FF",X"7F",X"FF",
		X"FF",X"FF",X"7F",X"FF",X"5F",X"FF",X"57",X"FF",X"5F",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"5F",X"FF",X"57",X"FF",X"5F",X"FF",X"7F",X"FF",X"FF",X"FF",X"7F",X"FF",X"7F",X"FF",
		X"FF",X"FF",X"7F",X"FF",X"5F",X"FF",X"5F",X"FF",X"57",X"FF",X"55",X"FF",X"55",X"5F",X"55",X"57",
		X"FF",X"FE",X"EF",X"E7",X"FF",X"BE",X"FD",X"FB",X"FA",X"EE",X"6F",X"6F",X"FE",X"FB",X"EF",X"AE",
		X"55",X"7F",X"55",X"FF",X"55",X"FF",X"57",X"FF",X"5F",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"57",X"FF",X"57",X"FF",X"57",X"FF",X"57",X"FF",X"57",X"FF",X"57",X"FF",X"57",X"FF",X"57",X"FF",
		X"55",X"FF",X"55",X"FF",X"55",X"FF",X"55",X"FF",X"57",X"FF",X"57",X"FF",X"57",X"FF",X"57",X"FF",
		X"55",X"5F",X"55",X"5F",X"55",X"5F",X"55",X"5F",X"55",X"5F",X"55",X"5F",X"55",X"7F",X"55",X"7F",
		X"55",X"57",X"55",X"57",X"55",X"57",X"55",X"57",X"55",X"57",X"55",X"57",X"55",X"57",X"55",X"57",
		X"55",X"5F",X"55",X"5F",X"55",X"57",X"55",X"57",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"5F",X"55",X"5F",X"55",X"7F",X"55",X"7F",X"55",X"7F",X"55",X"7F",X"55",X"7F",X"55",X"5F",
		X"55",X"57",X"55",X"D7",X"55",X"57",X"55",X"57",X"55",X"5F",X"55",X"5F",X"55",X"5F",X"55",X"5F",
		X"55",X"57",X"55",X"57",X"55",X"57",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"57",X"FF",X"55",X"FF",X"55",X"FF",X"55",X"7F",X"55",X"7F",X"55",X"5F",X"55",X"5F",X"55",X"57",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"5F",X"FF",
		X"55",X"7F",X"55",X"7F",X"55",X"7F",X"55",X"7F",X"55",X"7F",X"55",X"7F",X"55",X"7F",X"55",X"7F",
		X"5F",X"FF",X"5F",X"FF",X"5F",X"FF",X"57",X"FF",X"57",X"FF",X"57",X"FF",X"57",X"FF",X"57",X"FF",
		X"57",X"FF",X"5F",X"FF",X"5F",X"FF",X"7F",X"FF",X"7F",X"FF",X"5F",X"FF",X"5F",X"FF",X"5F",X"FF",
		X"55",X"7F",X"55",X"7F",X"55",X"7F",X"55",X"7F",X"55",X"7F",X"55",X"7F",X"55",X"7F",X"55",X"7F",
		X"55",X"5F",X"55",X"5F",X"55",X"5F",X"55",X"5F",X"55",X"5F",X"55",X"5F",X"55",X"5F",X"55",X"5F",
		X"5F",X"FF",X"5F",X"FF",X"5F",X"FF",X"57",X"FF",X"57",X"FF",X"57",X"FF",X"55",X"FF",X"55",X"7F",
		X"55",X"5F",X"55",X"5F",X"55",X"5F",X"55",X"5F",X"55",X"7F",X"55",X"7F",X"55",X"FF",X"55",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CF",X"FF",X"CF",X"FF",X"FF",X"FF",X"7F",X"FF",
		X"73",X"FF",X"73",X"FF",X"73",X"FF",X"7C",X"FF",X"5C",X"FF",X"5C",X"FF",X"5F",X"3F",X"57",X"3F",
		X"57",X"0F",X"57",X"0F",X"57",X"CF",X"55",X"C3",X"55",X"F0",X"55",X"70",X"55",X"7C",X"55",X"5C",
		X"55",X"5F",X"55",X"57",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"FE",X"FF",X"FF",X"FB",X"FC",X"FF",X"FF",X"BF",X"FF",X"2E",X"FF",X"FF",X"FD",X"D3",
		X"FF",X"39",X"FF",X"FF",X"FE",X"F3",X"FF",X"FE",X"FF",X"FC",X"FF",X"FF",X"FF",X"EF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"FF",X"3F",X"FF",
		X"0F",X"FF",X"CF",X"FF",X"F0",X"FF",X"70",X"3F",X"7C",X"0F",X"5F",X"03",X"57",X"C0",X"55",X"F0",
		X"7F",X"FF",X"FF",X"FE",X"3F",X"BF",X"CD",X"F3",X"FC",X"FF",X"7B",X"7F",X"E3",X"CF",X"37",X"FD",
		X"FF",X"1B",X"73",X"F1",X"FF",X"7F",X"FF",X"ED",X"FB",X"FF",X"FF",X"FB",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",
		X"ED",X"DC",X"FC",X"7F",X"DF",X"CF",X"3D",X"F7",X"F3",X"FF",X"DF",X"8F",X"36",X"7F",X"BF",X"3F",
		X"73",X"1F",X"2F",X"FF",X"FB",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"7C",X"55",X"5F",X"55",X"57",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"FF",X"00",X"03",X"F0",X"00",X"7C",X"00",X"5F",X"C0",X"55",X"FF",X"55",X"57",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"03",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"5F",X"FF",
		X"57",X"FF",X"5F",X"FF",X"5F",X"FF",X"5F",X"FF",X"7F",X"FF",X"7F",X"FF",X"7F",X"FF",X"7F",X"FF",
		X"55",X"5F",X"55",X"7F",X"55",X"7F",X"55",X"FF",X"55",X"FF",X"57",X"FF",X"57",X"FF",X"57",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"57",X"55",X"5F",
		X"55",X"FF",X"57",X"FF",X"5F",X"FF",X"7F",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"57",X"55",X"5F",X"55",X"7F",
		X"55",X"55",X"55",X"5F",X"55",X"FF",X"5F",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"57",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AD",X"AA",X"AB",X"AA",X"AB",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"B5",X"AA",X"B5",X"AA",X"B5",X"AA",X"B5",X"AA",X"B5",X"AA",X"AD",X"AA",X"AD",X"AA",X"AD",
		X"AA",X"D5",X"AA",X"D5",X"AA",X"D5",X"AA",X"D5",X"AA",X"D5",X"AA",X"D5",X"AA",X"D5",X"AA",X"B5",
		X"AD",X"7A",X"AD",X"7A",X"AB",X"7A",X"AB",X"EA",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",
		X"B5",X"57",X"B5",X"57",X"B5",X"D7",X"B5",X"5E",X"B7",X"5E",X"B5",X"5E",X"B5",X"5E",X"AD",X"7A",
		X"B5",X"55",X"B5",X"55",X"B5",X"D5",X"B5",X"55",X"B7",X"55",X"B5",X"55",X"B5",X"55",X"B5",X"55",
		X"AB",X"55",X"AD",X"55",X"AD",X"75",X"AD",X"55",X"AD",X"D5",X"AD",X"55",X"AD",X"55",X"B5",X"55",
		X"AA",X"D5",X"AA",X"D5",X"AA",X"D5",X"AA",X"D5",X"AB",X"75",X"AB",X"55",X"AB",X"55",X"AB",X"55",
		X"AA",X"AB",X"AA",X"AB",X"AA",X"AD",X"AA",X"AD",X"AA",X"AD",X"AA",X"B5",X"AA",X"B5",X"AA",X"B5",
		X"55",X"55",X"55",X"55",X"55",X"55",X"D5",X"55",X"B5",X"55",X"AF",X"55",X"AA",X"FF",X"AA",X"AA",
		X"B5",X"56",X"D5",X"55",X"DD",X"55",X"D5",X"55",X"75",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"D6",X"AA",X"D6",X"AB",X"56",X"AB",X"56",X"AB",X"56",X"AD",X"56",X"AD",X"56",X"AD",X"56",
		X"5E",X"AA",X"5E",X"AB",X"7A",X"AB",X"7A",X"AB",X"7A",X"AE",X"7A",X"AE",X"EA",X"B6",X"EA",X"B6",
		X"55",X"5B",X"55",X"5D",X"5D",X"79",X"55",X"79",X"75",X"E9",X"55",X"E9",X"57",X"A9",X"57",X"A9",
		X"AD",X"55",X"AD",X"55",X"B5",X"75",X"B5",X"55",X"D7",X"55",X"D5",X"55",X"D5",X"55",X"55",X"55",
		X"AA",X"AD",X"AA",X"B5",X"AA",X"B5",X"AA",X"D5",X"AA",X"D5",X"AB",X"75",X"AB",X"55",X"AD",X"55",
		X"57",X"AA",X"5E",X"AA",X"7A",X"AA",X"7A",X"AA",X"EA",X"AA",X"EA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"55",X"55",X"55",X"57",X"5D",X"57",X"55",X"5E",X"75",X"7A",X"55",X"7A",X"55",X"EA",X"55",X"EA",
		X"55",X"6A",X"55",X"6A",X"5D",X"6A",X"55",X"5A",X"75",X"5A",X"55",X"5A",X"55",X"56",X"55",X"56",
		X"55",X"AA",X"55",X"AA",X"5D",X"AA",X"55",X"AA",X"75",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",
		X"59",X"AA",X"59",X"AA",X"5D",X"AA",X"56",X"AA",X"76",X"AA",X"56",X"AA",X"56",X"AA",X"56",X"AA",
		X"A1",X"AA",X"A1",X"AA",X"AD",X"AA",X"A1",X"AA",X"B1",X"AA",X"69",X"AA",X"69",X"AA",X"59",X"AA",
		X"81",X"AA",X"81",X"AA",X"AD",X"AA",X"A1",X"AA",X"B1",X"AA",X"A1",X"AA",X"A1",X"AA",X"A1",X"AA",
		X"E0",X"6A",X"A0",X"6A",X"AC",X"6A",X"80",X"6A",X"B0",X"6A",X"81",X"AA",X"81",X"AA",X"81",X"AA",
		X"57",X"D6",X"57",X"1A",X"57",X"1A",X"5C",X"1A",X"5C",X"1A",X"5C",X"1A",X"70",X"1A",X"70",X"5A",
		X"AB",X"F5",X"AF",X"F7",X"B7",X"F5",X"B7",X"FF",X"77",X"FF",X"D7",X"FF",X"D7",X"FE",X"D7",X"F6",
		X"AA",X"A5",X"AA",X"AA",X"AE",X"AA",X"AA",X"AA",X"B8",X"AB",X"A8",X"AB",X"A8",X"2F",X"A8",X"FD",
		X"6A",X"54",X"6D",X"54",X"69",X"54",X"75",X"54",X"65",X"54",X"A9",X"54",X"AA",X"54",X"AA",X"94",
		X"56",X"A8",X"56",X"A0",X"5E",X"A0",X"5A",X"A0",X"7A",X"94",X"5A",X"94",X"5A",X"94",X"6A",X"54",
		X"AB",X"5A",X"AD",X"6A",X"AD",X"6A",X"B5",X"7A",X"B5",X"AA",X"D7",X"AA",X"D5",X"AA",X"55",X"A8",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AE",X"AA",X"BA",X"AA",X"DA",
		X"AA",X"55",X"AA",X"95",X"AA",X"95",X"AA",X"A5",X"AA",X"A9",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"D5",X"55",X"55",X"55",X"95",X"55",X"95",X"55",X"A5",X"55",X"A5",X"55",X"A9",X"55",X"AA",X"55",
		X"AA",X"D5",X"AA",X"D5",X"AB",X"55",X"AD",X"55",X"AD",X"55",X"B5",X"55",X"B5",X"55",X"D5",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AE",X"AA",X"AA",X"AB",X"BA",X"AB",X"AA",X"AD",X"AA",X"B5",X"AA",X"B5",
		X"AA",X"D5",X"AA",X"D5",X"AA",X"55",X"AA",X"95",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"7F",X"FF",X"7F",X"FF",X"7F",X"FF",X"EB",X"FF",X"AB",X"FD",X"AB",X"FD",X"AA",X"F5",X"AA",X"F5",
		X"00",X"00",X"00",X"00",X"FF",X"C0",X"FF",X"F0",X"57",X"F0",X"77",X"FC",X"57",X"FC",X"5F",X"FF",
		X"02",X"00",X"0A",X"00",X"08",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"A0",X"0A",X"A0",X"0A",X"A0",X"0A",X"80",X"0A",X"80",X"02",X"80",X"02",X"00",X"02",X"00",
		X"00",X"00",X"00",X"00",X"00",X"2A",X"02",X"AA",X"0A",X"AA",X"AA",X"AA",X"0A",X"A8",X"0A",X"A8",
		X"AA",X"00",X"AA",X"00",X"A8",X"00",X"A8",X"00",X"A0",X"00",X"A0",X"00",X"80",X"00",X"80",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"AA",X"A0",X"AA",X"A0",X"AA",X"80",X"AA",X"80",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"54",X"55",X"50",X"15",X"42",X"05",X"0A",
		X"75",X"55",X"D5",X"55",X"D5",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AE",X"AB",X"AA",X"AD",X"BA",X"B5",X"AA",X"D5",X"AB",X"55",X"AD",X"55",
		X"AA",X"95",X"AA",X"95",X"AE",X"95",X"AA",X"A5",X"BA",X"A5",X"AA",X"A5",X"AA",X"A9",X"AA",X"AA",
		X"55",X"40",X"55",X"50",X"55",X"54",X"A5",X"54",X"A9",X"55",X"A9",X"55",X"AA",X"55",X"AA",X"55",
		X"00",X"00",X"C0",X"00",X"C0",X"00",X"50",X"00",X"54",X"00",X"54",X"00",X"55",X"00",X"55",X"40",
		X"00",X"00",X"00",X"00",X"A0",X"00",X"80",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A8",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"AA",X"A0",X"AA",X"80",X"AA",X"00",
		X"43",X"AA",X"43",X"AA",X"03",X"AA",X"0E",X"AA",X"3A",X"AA",X"EA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"50",X"3A",X"50",X"3A",X"50",X"3A",X"50",X"3A",X"50",X"3A",X"50",X"3A",X"40",X"EA",X"40",X"EA",
		X"54",X"0E",X"54",X"0E",X"54",X"0E",X"50",X"0E",X"50",X"0E",X"50",X"3E",X"50",X"3A",X"50",X"3A",
		X"55",X"03",X"55",X"03",X"55",X"03",X"54",X"0F",X"54",X"0E",X"54",X"0E",X"54",X"0E",X"54",X"0E",
		X"D5",X"50",X"D5",X"40",X"55",X"40",X"55",X"40",X"55",X"40",X"55",X"40",X"55",X"40",X"55",X"03",
		X"AA",X"AA",X"AA",X"AB",X"AE",X"AD",X"AA",X"B4",X"BA",X"D4",X"AB",X"50",X"AD",X"50",X"B5",X"50",
		X"AB",X"EB",X"AA",X"AF",X"AE",X"AA",X"AA",X"AA",X"BA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"5E",X"AE",X"5E",X"BE",X"5E",X"BE",X"5E",X"BA",X"5E",X"FA",X"5E",X"FA",X"7E",X"FA",X"7A",X"EB",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"54",X"00",X"57",X"80",
		X"AA",X"00",X"A8",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AF",X"AA",X"80",
		X"02",X"AA",X"06",X"AA",X"0A",X"AA",X"1A",X"AA",X"2A",X"AA",X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"05",X"AA",X"15",X"A8",X"15",X"A8",X"17",X"A0",X"67",X"A0",X"AB",X"81",X"AA",X"82",X"AA",
		X"AA",X"80",X"AA",X"80",X"AA",X"80",X"AA",X"01",X"AA",X"01",X"AA",X"01",X"AA",X"05",X"AA",X"05",
		X"3E",X"A8",X"3A",X"A8",X"3A",X"A0",X"FA",X"A0",X"EA",X"A0",X"EA",X"A0",X"EA",X"80",X"EA",X"80",
		X"C0",X"3E",X"00",X"3E",X"00",X"FA",X"00",X"FA",X"03",X"EA",X"03",X"AA",X"0F",X"AA",X"0E",X"A8",
		X"AF",X"BF",X"BE",X"BE",X"AA",X"D5",X"AB",X"54",X"AD",X"43",X"AD",X"0F",X"B4",X"3F",X"C0",X"3F",
		X"AA",X"BA",X"BA",X"FF",X"BA",X"FB",X"FA",X"EB",X"FB",X"EB",X"EB",X"EB",X"EB",X"AF",X"EB",X"AF",
		X"00",X"EA",X"00",X"EA",X"00",X"EA",X"00",X"EA",X"00",X"EA",X"00",X"FA",X"00",X"3A",X"00",X"3A",
		X"00",X"EA",X"00",X"EA",X"00",X"EA",X"00",X"EA",X"00",X"EA",X"00",X"EA",X"00",X"EA",X"00",X"EA",
		X"00",X"0C",X"00",X"0D",X"00",X"0A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"FA",X"00",X"EA",
		X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"0F",
		X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"03",X"C0",X"03",X"00",X"0F",X"FC",X"3F",X"0C",
		X"0F",X"00",X"03",X"00",X"03",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"FE",X"C0",X"32",X"3C",X"02",
		X"AF",X"EA",X"AB",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"5D",X"A9",X"7F",X"A5",X"FF",X"A5",X"FF",X"E5",X"FF",X"E5",X"FF",X"FC",X"FF",X"FF",X"BF",X"EA",
		X"2A",X"6A",X"2A",X"6A",X"E9",X"6A",X"E9",X"AA",X"F9",X"A9",X"79",X"A9",X"7D",X"A9",X"5D",X"A9",
		X"05",X"6A",X"05",X"6A",X"15",X"6A",X"16",X"6A",X"1A",X"6A",X"1A",X"6A",X"2A",X"6A",X"2A",X"6A",
		X"81",X"55",X"81",X"55",X"81",X"55",X"01",X"55",X"01",X"55",X"05",X"56",X"05",X"5A",X"05",X"6A",
		X"BF",X"EF",X"BF",X"AF",X"FE",X"BF",X"FA",X"17",X"E8",X"17",X"A8",X"57",X"A0",X"55",X"A0",X"55",
		X"83",X"AF",X"F3",X"FF",X"F3",X"FF",X"EF",X"FF",X"EF",X"FF",X"EF",X"FF",X"AF",X"FF",X"BF",X"FB",
		X"0E",X"AF",X"0E",X"AF",X"0E",X"AF",X"0E",X"AF",X"0E",X"AF",X"0E",X"AF",X"0E",X"AF",X"0E",X"AF",
		X"02",X"AA",X"42",X"A5",X"56",X"57",X"81",X"6B",X"83",X"AB",X"83",X"AB",X"03",X"AF",X"0E",X"AF",
		X"00",X"FE",X"02",X"FE",X"02",X"EA",X"02",X"AA",X"02",X"AA",X"02",X"AA",X"0A",X"AA",X"0A",X"AA",
		X"C0",X"FE",X"C0",X"FE",X"C0",X"FE",X"C0",X"FE",X"C0",X"FE",X"00",X"FE",X"00",X"FE",X"00",X"FE",
		X"F0",X"FE",X"F0",X"FE",X"C0",X"FE",X"C0",X"FE",X"C0",X"FE",X"C0",X"FE",X"C0",X"FE",X"C0",X"FE",
		X"30",X"0A",X"30",X"0A",X"30",X"0A",X"30",X"0A",X"30",X"2A",X"30",X"FE",X"30",X"FE",X"30",X"FE",
		X"03",X"FA",X"03",X"FA",X"00",X"FA",X"C0",X"2A",X"C0",X"0A",X"F0",X"0A",X"30",X"0A",X"30",X"0A",
		X"3F",X"EA",X"3F",X"FA",X"3F",X"FA",X"3F",X"FA",X"0F",X"FA",X"0F",X"FA",X"0F",X"FA",X"03",X"FA",
		X"AA",X"A0",X"AA",X"A8",X"2A",X"AA",X"3E",X"AA",X"3F",X"AA",X"3F",X"AA",X"3F",X"EA",X"3F",X"EA",
		X"AA",X"AA",X"AA",X"BE",X"AA",X"FE",X"AB",X"F2",X"AF",X"E0",X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"40",X"AA",X"02",X"AA",X"02",X"AA",X"02",X"AA",X"0E",X"AA",X"3E",X"AA",X"FA",X"AA",X"AA",X"AA",
		X"40",X"AA",X"40",X"AA",X"40",X"AA",X"40",X"AA",X"40",X"AA",X"40",X"AA",X"40",X"AA",X"40",X"AA",
		X"40",X"AA",X"50",X"AA",X"90",X"AA",X"90",X"AA",X"90",X"AA",X"90",X"AA",X"90",X"AA",X"50",X"AA",
		X"FE",X"AA",X"FE",X"AA",X"7E",X"AA",X"7E",X"AA",X"7E",X"AA",X"4F",X"AA",X"43",X"AA",X"40",X"AA",
		X"FF",X"FF",X"EA",X"FF",X"EA",X"AF",X"FA",X"AB",X"FA",X"AB",X"FE",X"AA",X"FE",X"AA",X"FE",X"AA",
		X"55",X"EA",X"55",X"F9",X"57",X"F9",X"5F",X"FE",X"5F",X"FE",X"7F",X"FF",X"7F",X"FF",X"FF",X"FF",
		X"4E",X"9A",X"4F",X"9A",X"57",X"5A",X"57",X"5A",X"57",X"6A",X"57",X"6A",X"57",X"6A",X"57",X"EA",
		X"E1",X"55",X"E1",X"55",X"E1",X"55",X"E2",X"55",X"8A",X"95",X"8A",X"99",X"8A",X"9A",X"4A",X"9A",
		X"5A",X"15",X"78",X"15",X"F8",X"15",X"F8",X"55",X"E8",X"55",X"E8",X"55",X"E8",X"55",X"E1",X"55",
		X"AA",X"A0",X"AA",X"A0",X"AA",X"83",X"AA",X"83",X"AA",X"8F",X"AA",X"87",X"AA",X"05",X"AA",X"05",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"AA",X"A8",X"AA",X"A8",X"AA",X"A0",X"AA",X"A0",
		X"AA",X"AF",X"AA",X"AF",X"AA",X"AF",X"AA",X"AF",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AA",
		X"AA",X"A0",X"AA",X"82",X"AA",X"82",X"AA",X"82",X"AA",X"82",X"AA",X"8F",X"AA",X"BF",X"AA",X"BF",
		X"AB",X"F2",X"AA",X"FF",X"AA",X"FF",X"AA",X"BF",X"AA",X"BC",X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",
		X"80",X"EA",X"83",X"FC",X"83",X"F2",X"8E",X"B2",X"AE",X"82",X"AF",X"82",X"AF",X"82",X"AB",X"C2",
		X"00",X"AA",X"02",X"2A",X"08",X"2A",X"28",X"2A",X"A0",X"AA",X"A0",X"AA",X"80",X"AA",X"80",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"2A",X"AA",X"0A",X"AA",
		X"FE",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"68",X"02",X"68",X"02",X"A8",X"0A",X"A0",X"2A",X"A0",X"2A",X"80",X"AA",X"C0",X"AA",X"C2",X"AA",
		X"9A",X"02",X"9A",X"02",X"9A",X"02",X"9A",X"02",X"58",X"02",X"68",X"02",X"68",X"02",X"68",X"02",
		X"55",X"FE",X"55",X"FE",X"55",X"FE",X"55",X"FE",X"55",X"FE",X"55",X"FE",X"55",X"FE",X"99",X"3E",
		X"5F",X"EA",X"5F",X"FA",X"5F",X"FA",X"57",X"FA",X"57",X"FA",X"57",X"FA",X"57",X"FE",X"55",X"FE",
		X"AA",X"AA",X"AA",X"AA",X"FA",X"AA",X"FF",X"AA",X"FF",X"AA",X"FF",X"AA",X"FF",X"EA",X"7F",X"EA",
		X"C2",X"AA",X"02",X"AA",X"0A",X"AA",X"0A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"AA",X"AA",
		X"FF",X"CA",X"FF",X"2A",X"FF",X"2A",X"FC",X"2A",X"FC",X"AA",X"F0",X"AA",X"F0",X"AA",X"C2",X"AA",
		X"FC",X"AA",X"F2",X"AA",X"A2",X"AA",X"A2",X"AA",X"A2",X"AA",X"A2",X"AA",X"A2",X"8A",X"EF",X"CA",
		X"AA",X"AA",X"CA",X"AA",X"CA",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"AA",X"AA",X"EB",X"AA",
		X"55",X"55",X"55",X"55",X"5D",X"55",X"55",X"55",X"75",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AE",X"AA",X"AA",X"AA",X"BA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"6A",X"55",X"6A",X"55",X"AA",X"55",X"AA",X"56",X"AA",X"5A",X"AA",X"6A",X"AA",X"AA",X"AA",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"56",X"55",X"5A",
		X"AA",X"BF",X"AA",X"BF",X"AA",X"FF",X"AA",X"FF",X"AB",X"FF",X"AF",X"FF",X"BF",X"FF",X"FF",X"FF",
		X"6A",X"AA",X"6A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AB",X"AA",X"AB",X"AA",X"AF",
		X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"6A",X"AA",
		X"AA",X"AA",X"6A",X"AA",X"6A",X"AA",X"6A",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",
		X"BF",X"FF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AF",X"FF",X"AF",X"FF",X"AF",X"FF",X"AF",X"FF",X"AF",X"FF",X"AF",X"FF",X"BF",X"FF",X"BF",X"FF",
		X"FF",X"FF",X"BF",X"FF",X"BF",X"FF",X"BF",X"FF",X"AF",X"FF",X"AF",X"FF",X"AF",X"FF",X"AF",X"FF",
		X"FA",X"AA",X"FA",X"AA",X"FA",X"AA",X"FA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"AA",X"AA",
		X"FE",X"AA",X"FE",X"AA",X"FE",X"AA",X"FE",X"AA",X"FE",X"AA",X"FE",X"AA",X"FE",X"AA",X"FE",X"AA",
		X"55",X"AA",X"55",X"6A",X"55",X"5A",X"55",X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"6A",X"FF",X"5A",X"FF",X"5A",X"FF",X"5A",X"BF",X"56",X"BF",X"56",X"AF",X"56",X"AF",X"55",X"AB",
		X"AF",X"FF",X"AB",X"FF",X"6B",X"FF",X"6B",X"FF",X"6B",X"FF",X"6B",X"FF",X"6B",X"FF",X"6B",X"FF",
		X"AF",X"FF",X"AF",X"FF",X"AF",X"FF",X"AF",X"FF",X"AF",X"FF",X"AF",X"FF",X"AF",X"FF",X"AF",X"FF",
		X"55",X"55",X"55",X"55",X"6D",X"55",X"AF",X"55",X"AF",X"D5",X"AF",X"F5",X"AF",X"FD",X"AF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"BF",X"FF",X"AF",X"FF",X"AB",X"FF",X"6A",X"FF",X"5A",X"BF",X"56",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"A9",X"55",X"A9",X"55",X"A9",X"55",X"A9",X"55",X"A9",X"55",X"A9",X"55",X"A9",X"55",X"A9",X"55",
		X"56",X"A5",X"56",X"A5",X"56",X"A5",X"DA",X"A5",X"5A",X"A5",X"6A",X"95",X"6A",X"95",X"AA",X"55",
		X"55",X"6A",X"55",X"6A",X"55",X"AA",X"55",X"A9",X"55",X"A9",X"55",X"A9",X"55",X"A9",X"55",X"A9",
		X"55",X"AB",X"55",X"AB",X"55",X"AB",X"56",X"AB",X"56",X"AB",X"56",X"AF",X"5A",X"AF",X"5A",X"AF",
		X"55",X"6A",X"55",X"6A",X"55",X"6A",X"55",X"6A",X"55",X"6A",X"55",X"6A",X"55",X"AB",X"55",X"AB",
		X"FF",X"FD",X"FF",X"F5",X"FF",X"D5",X"FF",X"55",X"FD",X"55",X"F5",X"55",X"D5",X"55",X"55",X"55",
		X"FF",X"FD",X"FF",X"F5",X"FF",X"D5",X"FF",X"55",X"FD",X"55",X"F5",X"55",X"D5",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"AA",X"FF",X"AA",X"FF",X"AA",X"FF",X"AA",X"FF",X"AA",X"FF",X"AA",X"FF",X"AA",X"FF",X"AA",
		X"AA",X"AA",X"AA",X"A9",X"AA",X"A5",X"AA",X"95",X"AA",X"55",X"A9",X"55",X"A5",X"55",X"95",X"55",
		X"FF",X"AA",X"FF",X"AA",X"FE",X"AA",X"FE",X"AA",X"FA",X"AA",X"FA",X"AA",X"EA",X"AA",X"AA",X"AA",
		X"FF",X"EA",X"FF",X"EA",X"FF",X"EA",X"FF",X"EA",X"FF",X"EA",X"FF",X"AA",X"FF",X"AA",X"FF",X"AA",
		X"FF",X"FA",X"FF",X"FA",X"FF",X"FA",X"FF",X"FA",X"FF",X"FA",X"FF",X"FA",X"FF",X"FA",X"FF",X"FA",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"51",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"75",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"54",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"FF",X"AB",X"FF",X"AB",X"FF",X"AB",X"FF",X"AF",X"FF",X"AF",X"FF",X"BF",X"FF",X"FF",X"FF",
		X"AA",X"BF",X"AA",X"BF",X"AA",X"BF",X"AA",X"BF",X"AA",X"BF",X"AA",X"FF",X"AA",X"FF",X"AA",X"FF",
		X"AA",X"AF",X"AA",X"AF",X"AA",X"AF",X"AA",X"AF",X"AA",X"AF",X"AA",X"AF",X"AA",X"AF",X"AA",X"AF",
		X"FF",X"AA",X"FE",X"AA",X"FE",X"AA",X"FE",X"AA",X"FA",X"AA",X"FA",X"AA",X"EA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"FF",X"EA",X"FF",X"EA",X"FF",X"EA",X"FF",X"AA",X"FF",X"AA",X"FF",X"AA",
		X"55",X"5A",X"55",X"5A",X"55",X"5A",X"55",X"5A",X"55",X"5A",X"55",X"5A",X"55",X"5A",X"55",X"5A",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"AA",X"AA",X"AA",X"AA",
		X"55",X"5A",X"55",X"5A",X"55",X"5A",X"55",X"5A",X"55",X"5A",X"55",X"5A",X"55",X"5A",X"55",X"5A",
		X"FF",X"FA",X"FF",X"FA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"A5",X"FF",X"A5",X"FF",X"A5",X"FF",X"A5",X"FF",X"A5",X"FF",X"A5",X"FF",X"A5",X"FF",X"A5",
		X"AA",X"AA",X"AA",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"0A",X"AA",
		X"BF",X"77",X"AB",X"DF",X"AF",X"FF",X"83",X"FF",X"A0",X"00",X"00",X"00",X"A8",X"00",X"AA",X"FF",
		X"EA",X"AA",X"FE",X"AA",X"AA",X"AA",X"2A",X"AA",X"02",X"AA",X"2A",X"AA",X"AA",X"A8",X"FA",X"A8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"50",X"00",X"50",X"00",X"54",X"00",X"55",X"00",
		X"02",X"AA",X"00",X"AA",X"00",X"2A",X"00",X"0A",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AF",X"FF",X"BF",X"FF",X"AF",X"FF",X"A8",X"00",X"AA",X"00",X"2A",X"82",X"02",X"A2",X"00",X"00",
		X"FE",X"A8",X"FA",X"A0",X"EA",X"A0",X"AA",X"80",X"AA",X"80",X"A8",X"00",X"80",X"00",X"00",X"00",
		X"55",X"50",X"55",X"54",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"54",X"00",X"55",X"40",X"55",X"50",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"05",
		X"55",X"55",X"55",X"55",X"55",X"55",X"15",X"55",X"05",X"55",X"05",X"55",X"01",X"55",X"00",X"55",
		X"00",X"05",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"15",X"55",X"01",X"55",X"00",X"15",X"00",X"05",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"05",X"50",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"65",X"55",X"59",X"55",X"56",X"55",X"56",X"55",X"56",X"55",X"56",X"55",X"56",X"55",X"56",
		X"59",X"55",X"59",X"55",X"59",X"55",X"59",X"55",X"59",X"55",X"59",X"55",X"59",X"55",X"59",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"59",X"55",X"59",X"55",X"59",X"55",X"59",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"59",X"55",X"59",X"55",X"59",X"55",X"59",X"55",X"59",X"55",X"59",X"55",X"59",X"55",X"59",X"55",
		X"55",X"65",X"55",X"65",X"55",X"65",X"55",X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"56",X"55",X"56",X"55",X"56",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"59",X"55",X"65",X"55",X"65",X"55",X"65",
		X"55",X"55",X"55",X"65",X"59",X"55",X"59",X"55",X"59",X"55",X"59",X"55",X"59",X"55",X"59",X"55",
		X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"59",X"56",X"55",
		X"55",X"56",X"55",X"56",X"55",X"56",X"55",X"56",X"55",X"95",X"65",X"55",X"55",X"55",X"55",X"55",
		X"59",X"55",X"59",X"55",X"59",X"55",X"59",X"55",X"59",X"55",X"59",X"55",X"59",X"55",X"59",X"55",
		X"55",X"95",X"55",X"95",X"55",X"95",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"95",X"55",X"95",X"55",X"95",X"55",X"95",X"55",X"95",X"55",X"95",X"55",X"95",
		X"55",X"56",X"55",X"56",X"55",X"56",X"55",X"56",X"55",X"56",X"55",X"56",X"55",X"56",X"55",X"56",
		X"03",X"0C",X"21",X"2C",X"89",X"A0",X"AD",X"80",X"89",X"A0",X"21",X"2C",X"03",X"0C",X"00",X"00",
		X"FF",X"FF",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",
		X"55",X"D5",X"55",X"F5",X"55",X"75",X"55",X"7D",X"55",X"5D",X"55",X"5F",X"55",X"55",X"55",X"55",
		X"5D",X"55",X"5D",X"55",X"5D",X"55",X"5D",X"55",X"5F",X"55",X"57",X"55",X"57",X"55",X"57",X"D5",
		X"55",X"F5",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"D7",X"D5",X"FF",X"55",X"55",X"55",
		X"55",X"75",X"55",X"75",X"55",X"75",X"55",X"75",X"55",X"75",X"55",X"75",X"55",X"75",X"55",X"75",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"C0",X"00",X"F0",X"00",X"30",X"00",X"30",X"00",X"FF",X"FF",X"F5",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"F3",X"FC",X"7B",X"FE",X"CC",X"FF",X"FF",X"FF",X"FC",X"FF",X"F7",X"FF",X"CF",X"FF",X"FF",
		X"CF",X"FF",X"FD",X"F7",X"CC",X"DF",X"FF",X"BD",X"FF",X"FF",X"F7",X"7B",X"FC",X"CF",X"FF",X"FF",
		X"CF",X"FF",X"DF",X"FF",X"3C",X"CF",X"F7",X"BF",X"EF",X"DF",X"73",X"FF",X"FE",X"CF",X"5F",X"FF",
		X"FF",X"FF",X"CF",X"FF",X"FF",X"FF",X"B7",X"FF",X"CF",X"FF",X"BC",X"FF",X"DF",X"7F",X"FF",X"3F",
		X"3F",X"FF",X"FF",X"FF",X"BF",X"F3",X"DF",X"FF",X"FF",X"FF",X"FF",X"FE",X"B3",X"F3",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F3",X"FF",X"FF",X"FF",X"FF",X"FF",X"F3",
		X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FD",X"DF",X"FF",X"F3",X"FF",X"DF",X"FF",X"FF",X"FF",X"FB",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"FD",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"04",X"55",X"C0",X"55",X"F0",X"45",X"FC",X"01",X"F0",X"01",X"FF",X"00",X"FF",X"C0",X"FF",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"51",X"55",X"40",X"55",X"41",X"55",X"15",X"55",
		X"51",X"43",X"51",X"0F",X"40",X"3F",X"00",X"0F",X"03",X"CF",X"0F",X"FF",X"3F",X"FF",X"FF",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"45",X"55",X"41",X"55",X"11",X"55",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"59",X"55",X"59",X"55",X"59",X"55",X"59",X"55",
		X"55",X"55",X"55",X"55",X"56",X"55",X"56",X"55",X"56",X"55",X"56",X"55",X"56",X"55",X"59",X"55",
		X"55",X"56",X"55",X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
