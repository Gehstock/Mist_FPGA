library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_PGM is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_PGM is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"F3",X"C3",X"69",X"00",X"FF",X"FF",X"FF",X"C3",X"DE",X"06",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C3",X"12",X"1C",X"FF",X"FF",X"FF",X"FF",X"FF",X"C3",X"1E",X"1C",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C3",X"31",X"1C",X"FF",X"FF",X"FF",X"FF",X"FF",X"C3",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C3",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"C3",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C3",X"DB",X"07",X"AF",X"21",X"00",X"A8",X"06",X"08",X"77",
		X"23",X"10",X"FC",X"3E",X"9B",X"32",X"03",X"98",X"3A",X"01",X"98",X"CB",X"57",X"CA",X"9B",X"3B",
		X"21",X"00",X"88",X"11",X"00",X"8C",X"FD",X"21",X"8D",X"00",X"C3",X"3B",X"01",X"FD",X"21",X"94",
		X"00",X"C3",X"18",X"02",X"21",X"9A",X"00",X"C3",X"4B",X"02",X"52",X"41",X"4D",X"20",X"31",X"47",
		X"48",X"4A",X"4B",X"00",X"21",X"00",X"80",X"11",X"00",X"88",X"FD",X"21",X"B1",X"00",X"C3",X"3B",
		X"01",X"21",X"B7",X"00",X"C3",X"4B",X"02",X"32",X"43",X"20",X"52",X"4F",X"4D",X"20",X"20",X"20",
		X"00",X"21",X"00",X"00",X"DD",X"21",X"CB",X"00",X"C3",X"14",X"01",X"21",X"D1",X"00",X"C3",X"4B",
		X"02",X"32",X"45",X"00",X"21",X"00",X"10",X"DD",X"21",X"DE",X"00",X"C3",X"14",X"01",X"21",X"E4",
		X"00",X"C3",X"4B",X"02",X"32",X"46",X"00",X"21",X"00",X"20",X"DD",X"21",X"F1",X"00",X"C3",X"14",
		X"01",X"21",X"F7",X"00",X"C3",X"4B",X"02",X"32",X"48",X"00",X"21",X"00",X"30",X"DD",X"21",X"04",
		X"01",X"C3",X"14",X"01",X"21",X"0A",X"01",X"C3",X"4B",X"02",X"20",X"20",X"20",X"20",X"20",X"20",
		X"00",X"C3",X"D0",X"04",X"01",X"00",X"10",X"AF",X"16",X"FF",X"86",X"5F",X"7A",X"A6",X"57",X"7B",
		X"23",X"0D",X"C2",X"1A",X"01",X"08",X"3A",X"00",X"70",X"08",X"10",X"EE",X"FE",X"FF",X"C2",X"33",
		X"01",X"DD",X"E9",X"7A",X"FE",X"FF",X"C2",X"6C",X"02",X"DD",X"E9",X"DD",X"21",X"42",X"01",X"C3",
		X"82",X"01",X"44",X"4D",X"36",X"00",X"23",X"7D",X"BB",X"C2",X"44",X"01",X"08",X"3A",X"00",X"B0",
		X"08",X"7C",X"BA",X"C2",X"44",X"01",X"69",X"60",X"01",X"55",X"00",X"DD",X"21",X"62",X"01",X"C3",
		X"93",X"01",X"01",X"AA",X"55",X"DD",X"21",X"6C",X"01",X"C3",X"D5",X"01",X"01",X"FF",X"AA",X"DD",
		X"21",X"76",X"01",X"C3",X"93",X"01",X"01",X"00",X"FF",X"DD",X"21",X"80",X"01",X"C3",X"D5",X"01",
		X"FD",X"E9",X"06",X"00",X"70",X"7E",X"B8",X"C2",X"72",X"02",X"08",X"3A",X"00",X"B0",X"08",X"10",
		X"F3",X"DD",X"E9",X"08",X"3A",X"00",X"B0",X"08",X"7C",X"D9",X"67",X"D9",X"7D",X"D9",X"6F",X"D9",
		X"7B",X"D9",X"5F",X"D9",X"7A",X"D9",X"57",X"D9",X"7E",X"A8",X"C2",X"72",X"02",X"71",X"7E",X"A9",
		X"C2",X"72",X"02",X"23",X"7D",X"BB",X"C2",X"A8",X"01",X"08",X"3A",X"00",X"B0",X"08",X"7C",X"BA",
		X"C2",X"A8",X"01",X"D9",X"7C",X"D9",X"67",X"D9",X"7D",X"D9",X"6F",X"D9",X"7B",X"D9",X"5F",X"D9",
		X"7A",X"D9",X"57",X"DD",X"E9",X"08",X"3A",X"00",X"B0",X"08",X"7C",X"D9",X"67",X"D9",X"7D",X"D9",
		X"6F",X"D9",X"7B",X"D9",X"5F",X"D9",X"7A",X"D9",X"57",X"D9",X"EB",X"2B",X"7E",X"A8",X"C2",X"72",
		X"02",X"71",X"7E",X"A9",X"C2",X"72",X"02",X"08",X"3A",X"00",X"B0",X"08",X"7D",X"BB",X"C2",X"EB",
		X"01",X"7C",X"BA",X"C2",X"EB",X"01",X"D9",X"7C",X"D9",X"67",X"D9",X"7D",X"D9",X"6F",X"D9",X"7B",
		X"D9",X"5F",X"D9",X"7A",X"D9",X"57",X"DD",X"E9",X"21",X"00",X"88",X"11",X"00",X"8C",X"06",X"10",
		X"DD",X"21",X"27",X"02",X"C3",X"38",X"02",X"21",X"00",X"90",X"11",X"00",X"94",X"06",X"00",X"DD",
		X"21",X"36",X"02",X"C3",X"38",X"02",X"FD",X"E9",X"70",X"23",X"7D",X"BB",X"C2",X"38",X"02",X"08",
		X"3A",X"00",X"B0",X"08",X"7C",X"BA",X"C2",X"38",X"02",X"DD",X"E9",X"EB",X"21",X"6E",X"8B",X"1A",
		X"B7",X"CA",X"69",X"02",X"D6",X"30",X"F2",X"5B",X"02",X"3E",X"10",X"77",X"08",X"3A",X"00",X"B0",
		X"08",X"01",X"E0",X"FF",X"09",X"13",X"C3",X"4F",X"02",X"EB",X"23",X"E9",X"3A",X"00",X"B0",X"C3",
		X"6C",X"02",X"3A",X"00",X"B0",X"C3",X"72",X"02",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"1A",X"CD",X"DC",X"14",X"D2",X"9E",X"15",X"CD",X"97",X"02",X"CD",X"1A",X"03",X"CD",X"6A",X"03",
		X"3E",X"01",X"CD",X"CE",X"15",X"18",X"F3",X"21",X"2B",X"86",X"01",X"18",X"01",X"36",X"00",X"23",
		X"0B",X"78",X"B1",X"20",X"F8",X"C9",X"CD",X"07",X"03",X"D0",X"DD",X"7E",X"0B",X"E6",X"07",X"FE",
		X"01",X"C0",X"CD",X"FF",X"02",X"77",X"23",X"FD",X"5E",X"03",X"FD",X"56",X"04",X"CB",X"7A",X"C4",
		X"F5",X"22",X"CB",X"23",X"CB",X"12",X"73",X"23",X"72",X"23",X"AF",X"77",X"23",X"EB",X"2A",X"5D",
		X"87",X"3A",X"1D",X"82",X"4F",X"06",X"00",X"DD",X"7E",X"08",X"CB",X"7F",X"20",X"0B",X"B7",X"ED",
		X"42",X"01",X"18",X"00",X"B7",X"ED",X"42",X"18",X"08",X"79",X"2F",X"4F",X"09",X"01",X"18",X"00",
		X"09",X"EB",X"73",X"23",X"72",X"23",X"DD",X"7E",X"0A",X"77",X"21",X"C2",X"87",X"35",X"C9",X"DD",
		X"CB",X"08",X"7E",X"C8",X"CB",X"FF",X"C9",X"21",X"2B",X"86",X"11",X"07",X"00",X"06",X"28",X"7E",
		X"B7",X"20",X"02",X"37",X"C9",X"19",X"10",X"F7",X"B7",X"C9",X"21",X"2B",X"86",X"11",X"07",X"00",
		X"06",X"28",X"7E",X"B7",X"28",X"06",X"CD",X"30",X"03",X"CD",X"4D",X"03",X"19",X"10",X"F3",X"C9",
		X"C5",X"D5",X"E5",X"23",X"4E",X"23",X"46",X"23",X"7E",X"23",X"E5",X"66",X"6F",X"09",X"EB",X"E1",
		X"23",X"7E",X"CE",X"00",X"77",X"2B",X"72",X"2B",X"73",X"E1",X"D1",X"C1",X"C9",X"D5",X"E5",X"11",
		X"04",X"00",X"19",X"5E",X"23",X"56",X"EB",X"ED",X"5B",X"8C",X"87",X"B7",X"ED",X"52",X"38",X"07",
		X"E1",X"E5",X"23",X"AF",X"77",X"23",X"77",X"E1",X"D1",X"C9",X"21",X"2B",X"86",X"11",X"07",X"00",
		X"06",X"28",X"7E",X"B7",X"28",X"0A",X"CD",X"85",X"03",X"30",X"05",X"CD",X"CA",X"03",X"37",X"C9",
		X"19",X"10",X"EF",X"B7",X"C9",X"3A",X"9F",X"87",X"B7",X"28",X"02",X"37",X"C9",X"C5",X"D5",X"E5",
		X"2A",X"5D",X"87",X"3A",X"3A",X"81",X"5F",X"16",X"00",X"B7",X"ED",X"52",X"EB",X"E1",X"E5",X"23",
		X"23",X"23",X"23",X"7E",X"23",X"66",X"6F",X"EB",X"B7",X"ED",X"52",X"30",X"19",X"2A",X"5D",X"87",
		X"3A",X"3A",X"81",X"2F",X"5F",X"16",X"00",X"19",X"EB",X"E1",X"E5",X"23",X"23",X"23",X"23",X"7E",
		X"23",X"66",X"6F",X"B7",X"ED",X"52",X"E1",X"D1",X"C1",X"C9",X"3A",X"7D",X"87",X"FE",X"05",X"D0",
		X"E5",X"11",X"96",X"87",X"01",X"07",X"00",X"ED",X"B0",X"E1",X"06",X"07",X"AF",X"77",X"23",X"10",
		X"FC",X"3A",X"96",X"87",X"E6",X"07",X"FE",X"01",X"20",X"08",X"FD",X"21",X"78",X"31",X"CD",X"62",
		X"15",X"C9",X"FE",X"02",X"20",X"08",X"FD",X"21",X"20",X"36",X"CD",X"62",X"15",X"C9",X"FE",X"03",
		X"20",X"08",X"FD",X"21",X"BC",X"1F",X"CD",X"62",X"15",X"C9",X"FE",X"04",X"C0",X"FD",X"21",X"40",
		X"34",X"CD",X"62",X"15",X"C9",X"CD",X"97",X"02",X"2A",X"5D",X"87",X"3A",X"3A",X"81",X"5F",X"16",
		X"00",X"B7",X"ED",X"52",X"25",X"22",X"92",X"87",X"21",X"2B",X"86",X"22",X"94",X"87",X"06",X"08",
		X"FD",X"21",X"57",X"87",X"78",X"32",X"C0",X"87",X"FD",X"7E",X"00",X"B7",X"28",X"0C",X"4F",X"C5",
		X"CD",X"4F",X"04",X"CD",X"78",X"04",X"C1",X"0D",X"20",X"F5",X"FD",X"2B",X"10",X"E6",X"C9",X"2A",
		X"92",X"87",X"CD",X"46",X"21",X"E6",X"3F",X"F6",X"40",X"5F",X"16",X"00",X"19",X"22",X"92",X"87",
		X"ED",X"5B",X"8C",X"87",X"B7",X"ED",X"52",X"D8",X"2A",X"5D",X"87",X"3A",X"3A",X"81",X"5F",X"16",
		X"00",X"B7",X"ED",X"52",X"22",X"92",X"87",X"C9",X"CD",X"07",X"03",X"D0",X"3A",X"C0",X"87",X"F6",
		X"80",X"77",X"23",X"CD",X"98",X"04",X"73",X"23",X"72",X"23",X"23",X"ED",X"5B",X"92",X"87",X"73",
		X"23",X"72",X"23",X"CD",X"DF",X"2A",X"77",X"C9",X"CD",X"46",X"21",X"F6",X"7F",X"5F",X"3A",X"4B",
		X"87",X"4F",X"CD",X"46",X"21",X"A1",X"57",X"C9",X"21",X"2B",X"86",X"11",X"07",X"00",X"06",X"28",
		X"0E",X"05",X"7E",X"E6",X"03",X"FE",X"01",X"20",X"05",X"CD",X"C2",X"04",X"0D",X"C8",X"19",X"10",
		X"F1",X"C9",X"E5",X"23",X"7E",X"23",X"B6",X"20",X"05",X"3E",X"01",X"CD",X"28",X"2C",X"E1",X"C9",
		X"3E",X"00",X"32",X"01",X"A8",X"32",X"02",X"A8",X"32",X"03",X"A8",X"32",X"04",X"A8",X"32",X"07",
		X"A8",X"32",X"06",X"A8",X"3E",X"93",X"32",X"03",X"98",X"3E",X"88",X"32",X"03",X"A0",X"31",X"68",
		X"80",X"21",X"68",X"80",X"0E",X"08",X"CD",X"88",X"07",X"3E",X"FF",X"32",X"EB",X"80",X"32",X"EC",
		X"80",X"21",X"0F",X"05",X"11",X"F2",X"80",X"01",X"3C",X"00",X"ED",X"B0",X"C3",X"2C",X"14",X"02",
		X"04",X"30",X"52",X"41",X"51",X"01",X"61",X"20",X"4A",X"4F",X"4E",X"01",X"39",X"90",X"41",X"52",
		X"4D",X"01",X"17",X"80",X"41",X"4A",X"4D",X"00",X"98",X"60",X"54",X"4A",X"43",X"00",X"85",X"70",
		X"45",X"4C",X"50",X"00",X"65",X"50",X"44",X"52",X"4A",X"00",X"43",X"30",X"4A",X"49",X"4D",X"00",
		X"30",X"10",X"44",X"41",X"4E",X"00",X"25",X"40",X"42",X"49",X"4C",X"3E",X"00",X"CD",X"F4",X"2B",
		X"21",X"18",X"00",X"01",X"01",X"20",X"CD",X"93",X"07",X"DF",X"1A",X"3A",X"1E",X"86",X"FE",X"02",
		X"20",X"2A",X"CF",X"38",X"18",X"50",X"4C",X"41",X"59",X"45",X"52",X"20",X"00",X"21",X"18",X"70",
		X"11",X"43",X"87",X"06",X"01",X"CD",X"06",X"07",X"CF",X"78",X"18",X"20",X"47",X"41",X"4D",X"45",
		X"20",X"4F",X"56",X"45",X"52",X"00",X"3E",X"3C",X"CD",X"CE",X"15",X"C9",X"CF",X"58",X"18",X"47",
		X"41",X"4D",X"45",X"20",X"4F",X"56",X"45",X"52",X"00",X"3E",X"3C",X"CD",X"CE",X"15",X"C9",X"CD",
		X"61",X"07",X"3E",X"FF",X"32",X"04",X"A8",X"CD",X"46",X"0B",X"CD",X"68",X"0B",X"CD",X"9E",X"0B",
		X"DF",X"2A",X"DF",X"3B",X"DF",X"4C",X"DF",X"5D",X"E7",X"07",X"0D",X"02",X"E7",X"05",X"15",X"01",
		X"CF",X"40",X"28",X"5B",X"20",X"48",X"49",X"47",X"48",X"20",X"53",X"43",X"4F",X"52",X"45",X"53",
		X"20",X"5B",X"00",X"11",X"F2",X"80",X"21",X"38",X"38",X"3E",X"01",X"08",X"D5",X"EB",X"7E",X"23",
		X"B6",X"23",X"B6",X"EB",X"D1",X"C8",X"E5",X"D5",X"08",X"32",X"00",X"80",X"08",X"06",X"02",X"11",
		X"00",X"80",X"CD",X"06",X"07",X"01",X"00",X"20",X"09",X"D1",X"06",X"06",X"CD",X"06",X"07",X"13",
		X"13",X"13",X"01",X"00",X"30",X"09",X"CD",X"B8",X"06",X"06",X"03",X"3E",X"20",X"CD",X"49",X"07",
		X"10",X"F9",X"06",X"03",X"1A",X"13",X"CD",X"49",X"07",X"10",X"F9",X"E1",X"01",X"10",X"00",X"09",
		X"08",X"C6",X"01",X"27",X"FE",X"11",X"DA",X"DB",X"05",X"C9",X"3A",X"F1",X"80",X"B7",X"C8",X"21",
		X"B8",X"00",X"01",X"05",X"20",X"CD",X"93",X"07",X"E7",X"05",X"17",X"05",X"3A",X"F1",X"80",X"FE",
		X"01",X"20",X"40",X"CF",X"18",X"B8",X"50",X"55",X"53",X"48",X"20",X"31",X"20",X"50",X"4C",X"41",
		X"59",X"45",X"52",X"20",X"53",X"54",X"41",X"52",X"54",X"20",X"42",X"55",X"54",X"54",X"4F",X"4E",
		X"00",X"CF",X"68",X"C8",X"5B",X"20",X"4F",X"52",X"20",X"5B",X"00",X"CF",X"30",X"D8",X"49",X"4E",
		X"53",X"45",X"52",X"54",X"20",X"41",X"4E",X"4F",X"54",X"48",X"45",X"52",X"20",X"43",X"4F",X"49",
		X"4E",X"00",X"C9",X"CF",X"48",X"B8",X"50",X"55",X"53",X"48",X"20",X"31",X"20",X"50",X"4C",X"41",
		X"59",X"45",X"52",X"00",X"CF",X"68",X"C8",X"5B",X"20",X"4F",X"52",X"20",X"5B",X"00",X"CF",X"28",
		X"D8",X"32",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"20",X"53",X"54",X"41",X"52",X"54",X"20",
		X"42",X"55",X"54",X"54",X"4F",X"4E",X"00",X"C9",X"F5",X"AF",X"C3",X"C1",X"06",X"F5",X"3A",X"C8",
		X"80",X"94",X"3D",X"67",X"CB",X"3C",X"CB",X"3C",X"CB",X"3C",X"CB",X"3C",X"CB",X"1D",X"CB",X"3C",
		X"CB",X"1D",X"CB",X"3C",X"CB",X"1D",X"D5",X"11",X"00",X"88",X"19",X"D1",X"F1",X"C9",X"E3",X"F5",
		X"C5",X"D5",X"56",X"23",X"5E",X"23",X"EB",X"CD",X"B8",X"06",X"1A",X"13",X"B7",X"CA",X"F6",X"06",
		X"CD",X"49",X"07",X"C3",X"EA",X"06",X"EB",X"D1",X"C1",X"F1",X"E3",X"C9",X"0E",X"03",X"C3",X"08",
		X"07",X"0E",X"00",X"C3",X"08",X"07",X"0E",X"01",X"F5",X"C5",X"D5",X"E5",X"CD",X"B8",X"06",X"78",
		X"3D",X"20",X"02",X"CB",X"81",X"1A",X"CB",X"40",X"20",X"05",X"07",X"07",X"07",X"07",X"1B",X"13",
		X"E6",X"0F",X"C2",X"34",X"07",X"CB",X"41",X"CA",X"36",X"07",X"3E",X"20",X"CB",X"49",X"C2",X"42",
		X"07",X"C3",X"3F",X"07",X"CB",X"81",X"C6",X"30",X"FE",X"3A",X"DA",X"3F",X"07",X"C6",X"07",X"CD",
		X"49",X"07",X"10",X"CB",X"E1",X"D1",X"C1",X"F1",X"C9",X"C5",X"D6",X"30",X"F2",X"51",X"07",X"3E",
		X"10",X"77",X"01",X"E0",X"FF",X"09",X"7C",X"FE",X"88",X"30",X"04",X"01",X"00",X"04",X"09",X"C1",
		X"C9",X"F5",X"C5",X"E5",X"21",X"00",X"88",X"0E",X"04",X"3E",X"10",X"CD",X"89",X"07",X"21",X"00",
		X"90",X"0E",X"01",X"CD",X"88",X"07",X"3E",X"00",X"32",X"03",X"A8",X"32",X"04",X"A8",X"32",X"07",
		X"A8",X"32",X"06",X"A8",X"E1",X"C1",X"F1",X"C9",X"AF",X"06",X"00",X"77",X"23",X"10",X"FC",X"0D",
		X"20",X"F9",X"C9",X"F5",X"C5",X"D5",X"E5",X"50",X"E5",X"CD",X"B8",X"06",X"3E",X"20",X"CD",X"49",
		X"07",X"10",X"F9",X"E1",X"7D",X"C6",X"08",X"6F",X"42",X"0D",X"20",X"EC",X"E1",X"D1",X"C1",X"F1",
		X"C9",X"E3",X"F5",X"C5",X"D5",X"56",X"23",X"5E",X"23",X"EB",X"CD",X"BD",X"06",X"1A",X"13",X"B7",
		X"CA",X"C9",X"07",X"CD",X"49",X"07",X"C3",X"BD",X"07",X"EB",X"D1",X"C1",X"F1",X"E3",X"C9",X"F5",
		X"C5",X"D5",X"E5",X"CD",X"BD",X"06",X"0E",X"01",X"C3",X"0F",X"07",X"F5",X"E5",X"C5",X"3A",X"00",
		X"B0",X"AF",X"32",X"01",X"A8",X"3C",X"32",X"01",X"A8",X"21",X"25",X"86",X"CB",X"0E",X"DA",X"98",
		X"09",X"3A",X"26",X"86",X"B7",X"C2",X"9B",X"09",X"3C",X"32",X"26",X"86",X"ED",X"73",X"BC",X"80",
		X"31",X"40",X"80",X"08",X"F5",X"D5",X"DD",X"E5",X"FD",X"E5",X"D9",X"C5",X"D5",X"E5",X"21",X"34",
		X"81",X"11",X"40",X"90",X"06",X"08",X"C5",X"CB",X"46",X"CC",X"39",X"0B",X"01",X"06",X"00",X"09",
		X"7E",X"12",X"23",X"13",X"7E",X"12",X"23",X"13",X"7E",X"12",X"09",X"13",X"7E",X"12",X"23",X"13",
		X"C1",X"10",X"E3",X"21",X"AC",X"81",X"11",X"61",X"90",X"06",X"07",X"C5",X"CB",X"46",X"CC",X"39",
		X"0B",X"01",X"06",X"00",X"09",X"3A",X"43",X"87",X"FE",X"02",X"20",X"17",X"3A",X"02",X"98",X"E6",
		X"08",X"28",X"10",X"7E",X"C6",X"08",X"12",X"01",X"08",X"00",X"09",X"13",X"13",X"7E",X"C6",X"01",
		X"C3",X"71",X"08",X"7E",X"C6",X"08",X"12",X"01",X"08",X"00",X"09",X"13",X"13",X"7E",X"2F",X"C6",
		X"F1",X"12",X"23",X"13",X"13",X"C1",X"10",X"C3",X"CD",X"6E",X"27",X"CD",X"CF",X"27",X"2A",X"C0",
		X"80",X"CB",X"7C",X"28",X"2B",X"29",X"ED",X"5B",X"C7",X"80",X"19",X"22",X"C7",X"80",X"7C",X"21",
		X"08",X"90",X"06",X"1C",X"77",X"23",X"23",X"10",X"FB",X"2A",X"C0",X"80",X"29",X"EB",X"2A",X"C4",
		X"80",X"B7",X"ED",X"52",X"22",X"C4",X"80",X"3A",X"C6",X"80",X"3F",X"CE",X"00",X"32",X"C6",X"80",
		X"3A",X"C5",X"80",X"47",X"21",X"27",X"86",X"AE",X"CB",X"5F",X"28",X"70",X"78",X"77",X"CB",X"3F",
		X"CB",X"3F",X"CB",X"3F",X"D6",X"20",X"ED",X"44",X"26",X"00",X"06",X"05",X"CB",X"27",X"CB",X"14",
		X"10",X"FA",X"6F",X"11",X"04",X"88",X"19",X"EB",X"21",X"28",X"86",X"7E",X"23",X"66",X"6F",X"23",
		X"7E",X"47",X"FE",X"01",X"28",X"1E",X"CD",X"46",X"21",X"0F",X"0F",X"E6",X"1F",X"FE",X"1B",X"30",
		X"F5",X"3C",X"32",X"2A",X"86",X"CD",X"46",X"21",X"0F",X"0F",X"0F",X"E6",X"0F",X"90",X"F2",X"FD",
		X"08",X"80",X"3C",X"47",X"23",X"10",X"FD",X"4E",X"21",X"60",X"26",X"09",X"09",X"7E",X"23",X"66",
		X"6F",X"E5",X"3A",X"2A",X"86",X"06",X"00",X"4F",X"09",X"06",X"1D",X"7E",X"B7",X"20",X"07",X"22",
		X"28",X"86",X"E1",X"10",X"01",X"04",X"7E",X"12",X"13",X"23",X"10",X"EF",X"21",X"71",X"82",X"06",
		X"0D",X"C5",X"CB",X"7E",X"C4",X"9F",X"09",X"11",X"2E",X"00",X"19",X"C1",X"10",X"F3",X"CD",X"38",
		X"0E",X"21",X"15",X"82",X"06",X"16",X"C5",X"46",X"CB",X"40",X"C4",X"C4",X"09",X"CB",X"58",X"C4",
		X"A1",X"0A",X"11",X"2E",X"00",X"19",X"C1",X"10",X"ED",X"3A",X"CB",X"80",X"4F",X"06",X"00",X"3C",
		X"FE",X"0F",X"38",X"01",X"AF",X"32",X"CB",X"80",X"21",X"CC",X"80",X"09",X"09",X"5E",X"23",X"56",
		X"ED",X"53",X"C0",X"80",X"ED",X"5B",X"37",X"81",X"7B",X"2F",X"5F",X"7A",X"2F",X"57",X"13",X"72",
		X"2B",X"73",X"CD",X"AF",X"16",X"E1",X"D1",X"C1",X"D9",X"FD",X"E1",X"DD",X"E1",X"D1",X"F1",X"08",
		X"ED",X"7B",X"BC",X"80",X"AF",X"32",X"26",X"86",X"CD",X"A6",X"19",X"C1",X"E1",X"F1",X"C9",X"CB",
		X"4E",X"C8",X"CB",X"5E",X"C0",X"E5",X"01",X"05",X"00",X"09",X"5E",X"23",X"56",X"13",X"13",X"13",
		X"23",X"23",X"46",X"23",X"23",X"7E",X"C6",X"04",X"6F",X"78",X"C6",X"04",X"67",X"1A",X"CD",X"BD",
		X"06",X"77",X"E1",X"C9",X"E5",X"CB",X"48",X"CA",X"81",X"0A",X"23",X"5E",X"23",X"56",X"D5",X"FD",
		X"E1",X"23",X"CB",X"68",X"28",X"05",X"35",X"20",X"02",X"CB",X"A8",X"23",X"CB",X"60",X"28",X"6D",
		X"35",X"20",X"6A",X"CB",X"F8",X"23",X"5E",X"23",X"56",X"13",X"13",X"13",X"13",X"13",X"1A",X"B7",
		X"C2",X"04",X"0A",X"13",X"1A",X"B7",X"C2",X"FD",X"09",X"CB",X"A0",X"CB",X"B8",X"EB",X"23",X"7E",
		X"23",X"66",X"6F",X"EB",X"72",X"2B",X"73",X"13",X"13",X"1A",X"CB",X"7F",X"28",X"3D",X"4F",X"C5",
		X"FD",X"7E",X"03",X"FD",X"AE",X"04",X"4F",X"FD",X"7E",X"04",X"B7",X"F2",X"1F",X"0A",X"2F",X"1F",
		X"CB",X"19",X"1F",X"CB",X"19",X"FD",X"7E",X"0B",X"FD",X"AE",X"0C",X"47",X"FD",X"7E",X"0C",X"B7",
		X"F2",X"34",X"0A",X"2F",X"1F",X"CB",X"18",X"1F",X"CB",X"18",X"78",X"B1",X"C1",X"CB",X"3F",X"CB",
		X"3F",X"4F",X"1A",X"CB",X"BF",X"91",X"F2",X"4A",X"0A",X"AF",X"3C",X"2B",X"77",X"CB",X"50",X"28",
		X"30",X"23",X"23",X"23",X"E5",X"5E",X"23",X"56",X"2A",X"C0",X"80",X"19",X"EB",X"E1",X"73",X"23",
		X"72",X"CB",X"88",X"7A",X"FE",X"02",X"38",X"19",X"FE",X"F8",X"30",X"15",X"CB",X"C8",X"23",X"23",
		X"7E",X"FE",X"1F",X"30",X"05",X"3E",X"E8",X"C3",X"80",X"0A",X"FE",X"E9",X"38",X"03",X"3E",X"20",
		X"77",X"E1",X"70",X"C9",X"CB",X"BE",X"21",X"1A",X"82",X"11",X"3B",X"81",X"7E",X"23",X"66",X"6F",
		X"23",X"23",X"23",X"7E",X"B7",X"28",X"01",X"12",X"23",X"13",X"7E",X"12",X"21",X"15",X"82",X"46",
		X"C9",X"CB",X"48",X"C8",X"E5",X"DD",X"E1",X"CB",X"78",X"28",X"14",X"CB",X"BE",X"DD",X"66",X"06",
		X"DD",X"6E",X"05",X"23",X"23",X"23",X"7E",X"FD",X"77",X"07",X"23",X"7E",X"FD",X"77",X"08",X"CB",
		X"50",X"28",X"72",X"DD",X"7E",X"07",X"FD",X"77",X"05",X"DD",X"7E",X"08",X"FD",X"77",X"06",X"DD",
		X"7E",X"09",X"FD",X"77",X"0D",X"DD",X"7E",X"0A",X"FD",X"77",X"0E",X"FD",X"E5",X"E1",X"CB",X"76",
		X"20",X"53",X"23",X"5E",X"23",X"56",X"23",X"4E",X"23",X"46",X"EB",X"09",X"EB",X"2B",X"73",X"23",
		X"72",X"23",X"4E",X"23",X"46",X"EB",X"09",X"EB",X"2B",X"73",X"DD",X"73",X"07",X"23",X"72",X"DD",
		X"72",X"08",X"7A",X"FD",X"CB",X"00",X"F6",X"FE",X"09",X"38",X"08",X"FE",X"F1",X"30",X"04",X"FD",
		X"CB",X"00",X"B6",X"23",X"23",X"23",X"5E",X"23",X"56",X"23",X"4E",X"23",X"46",X"EB",X"09",X"EB",
		X"2B",X"73",X"23",X"72",X"23",X"4E",X"23",X"46",X"EB",X"09",X"EB",X"2B",X"73",X"DD",X"73",X"09",
		X"23",X"72",X"DD",X"72",X"0A",X"DD",X"E5",X"E1",X"C9",X"AF",X"E5",X"DD",X"E1",X"DD",X"77",X"06",
		X"DD",X"77",X"0E",X"C9",X"00",X"00",X"DF",X"FF",X"CF",X"10",X"F8",X"3B",X"31",X"39",X"38",X"31",
		X"20",X"53",X"54",X"45",X"52",X"4E",X"20",X"45",X"4C",X"45",X"43",X"54",X"52",X"4F",X"4E",X"49",
		X"43",X"53",X"20",X"49",X"4E",X"43",X"00",X"C9",X"3A",X"F1",X"80",X"B7",X"28",X"1E",X"DF",X"F0",
		X"CD",X"B1",X"07",X"18",X"F0",X"43",X"52",X"45",X"44",X"49",X"54",X"53",X"20",X"5B",X"20",X"00",
		X"21",X"F0",X"68",X"11",X"F1",X"80",X"06",X"02",X"CD",X"CF",X"07",X"C9",X"DF",X"F3",X"CF",X"18",
		X"F0",X"49",X"4E",X"53",X"45",X"52",X"54",X"20",X"43",X"4F",X"49",X"4E",X"00",X"C9",X"AF",X"32",
		X"1A",X"86",X"DF",X"03",X"DF",X"0A",X"CF",X"20",X"00",X"31",X"53",X"54",X"00",X"21",X"08",X"10",
		X"11",X"2E",X"81",X"06",X"06",X"CD",X"06",X"07",X"CF",X"58",X"00",X"48",X"49",X"47",X"48",X"20",
		X"53",X"43",X"4F",X"52",X"45",X"00",X"21",X"08",X"68",X"11",X"F2",X"80",X"06",X"06",X"CD",X"06",
		X"07",X"3A",X"1E",X"86",X"FE",X"02",X"C0",X"CF",X"D0",X"00",X"32",X"4E",X"44",X"00",X"21",X"08",
		X"C0",X"11",X"31",X"81",X"06",X"06",X"CD",X"06",X"07",X"C9",X"DF",X"F5",X"CF",X"18",X"F0",X"53",
		X"48",X"49",X"50",X"53",X"20",X"4C",X"45",X"46",X"54",X"20",X"5B",X"20",X"00",X"21",X"F0",X"80",
		X"11",X"44",X"87",X"06",X"02",X"CD",X"06",X"07",X"C9",X"DF",X"7E",X"CF",X"40",X"78",X"50",X"4C",
		X"41",X"59",X"45",X"52",X"20",X"00",X"21",X"78",X"78",X"11",X"43",X"87",X"06",X"01",X"CD",X"06",
		X"07",X"CF",X"80",X"78",X"20",X"55",X"50",X"00",X"C9",X"CD",X"C5",X"0C",X"3E",X"00",X"32",X"B9",
		X"87",X"CD",X"F4",X"2B",X"21",X"43",X"87",X"36",X"01",X"23",X"CD",X"2A",X"0D",X"23",X"23",X"36",
		X"01",X"21",X"60",X"87",X"36",X"02",X"23",X"CD",X"2A",X"0D",X"23",X"23",X"36",X"01",X"3A",X"1E",
		X"86",X"FE",X"02",X"28",X"04",X"AF",X"32",X"61",X"87",X"CD",X"6E",X"21",X"CD",X"05",X"0E",X"FB",
		X"3E",X"99",X"32",X"5A",X"87",X"3E",X"99",X"32",X"58",X"87",X"AF",X"32",X"7D",X"87",X"32",X"7E",
		X"87",X"32",X"7F",X"87",X"32",X"1B",X"86",X"32",X"BF",X"87",X"32",X"BA",X"87",X"32",X"BB",X"87",
		X"32",X"C2",X"87",X"3C",X"32",X"C6",X"80",X"CD",X"43",X"0D",X"3E",X"3C",X"CD",X"CE",X"15",X"CD",
		X"27",X"16",X"CD",X"6E",X"21",X"3E",X"00",X"CD",X"F4",X"2B",X"21",X"44",X"87",X"7E",X"C6",X"99",
		X"27",X"77",X"B7",X"CC",X"4B",X"05",X"CD",X"EB",X"0C",X"3A",X"44",X"87",X"B7",X"C2",X"59",X"0C",
		X"3A",X"61",X"87",X"B7",X"20",X"F0",X"CD",X"EB",X"0C",X"CD",X"7D",X"12",X"CD",X"EB",X"0C",X"CD",
		X"7D",X"12",X"C3",X"32",X"14",X"21",X"00",X"00",X"22",X"2E",X"81",X"22",X"30",X"81",X"22",X"32",
		X"81",X"22",X"ED",X"80",X"22",X"EF",X"80",X"AF",X"21",X"43",X"87",X"06",X"1D",X"77",X"23",X"10",
		X"FC",X"21",X"60",X"87",X"06",X"1D",X"77",X"23",X"10",X"FC",X"C9",X"E5",X"21",X"43",X"87",X"11",
		X"60",X"87",X"06",X"1D",X"1A",X"4E",X"EB",X"12",X"71",X"EB",X"23",X"13",X"10",X"F6",X"E1",X"C9",
		X"3A",X"43",X"87",X"FE",X"02",X"20",X"15",X"3A",X"02",X"98",X"E6",X"08",X"28",X"0E",X"3E",X"00",
		X"32",X"02",X"98",X"3E",X"FF",X"32",X"07",X"A8",X"32",X"06",X"A8",X"C9",X"3E",X"10",X"32",X"02",
		X"98",X"3E",X"00",X"32",X"07",X"A8",X"32",X"06",X"A8",X"C9",X"3A",X"01",X"98",X"2F",X"E6",X"03",
		X"28",X"0E",X"FE",X"01",X"20",X"03",X"36",X"05",X"C9",X"FE",X"02",X"20",X"03",X"36",X"04",X"C9",
		X"36",X"03",X"C9",X"CD",X"61",X"07",X"CD",X"00",X"0D",X"21",X"CB",X"80",X"06",X"1F",X"AF",X"77",
		X"23",X"10",X"FC",X"3E",X"82",X"32",X"C1",X"87",X"CD",X"9E",X"0B",X"CD",X"52",X"27",X"CD",X"B6",
		X"27",X"CD",X"4F",X"3E",X"CD",X"E8",X"25",X"FD",X"21",X"B2",X"0E",X"CD",X"62",X"15",X"FD",X"21",
		X"81",X"02",X"CD",X"62",X"15",X"FD",X"21",X"67",X"28",X"CD",X"62",X"15",X"FD",X"21",X"9E",X"15",
		X"CD",X"62",X"15",X"DD",X"21",X"15",X"82",X"DD",X"7E",X"00",X"B7",X"C8",X"3A",X"B9",X"87",X"B7",
		X"28",X"06",X"CD",X"C5",X"19",X"C2",X"5D",X"14",X"CD",X"2A",X"19",X"DD",X"21",X"43",X"82",X"DD",
		X"CB",X"00",X"6E",X"C2",X"D8",X"0D",X"CD",X"DE",X"0D",X"CD",X"ED",X"1D",X"CD",X"E3",X"1D",X"CD",
		X"91",X"27",X"DD",X"36",X"03",X"03",X"DD",X"CB",X"00",X"EE",X"21",X"1F",X"86",X"34",X"7E",X"FE",
		X"09",X"20",X"15",X"AF",X"77",X"21",X"20",X"86",X"34",X"CD",X"62",X"27",X"CD",X"C3",X"27",X"3A",
		X"1A",X"86",X"B7",X"28",X"03",X"CD",X"9E",X"0B",X"CD",X"7A",X"15",X"C3",X"83",X"0D",X"3A",X"C1",
		X"87",X"3D",X"28",X"0E",X"32",X"C1",X"87",X"3A",X"1A",X"86",X"B7",X"C8",X"3E",X"82",X"32",X"C1",
		X"87",X"C9",X"3A",X"7D",X"87",X"FE",X"05",X"D0",X"3E",X"82",X"32",X"C1",X"87",X"FD",X"21",X"EE",
		X"37",X"CD",X"62",X"15",X"C9",X"CD",X"61",X"07",X"CD",X"00",X"0D",X"CD",X"EA",X"0B",X"3A",X"1E",
		X"86",X"3D",X"06",X"03",X"28",X"07",X"06",X"05",X"3E",X"04",X"CD",X"F4",X"2B",X"C5",X"CD",X"09",
		X"0C",X"3E",X"0C",X"CD",X"CE",X"15",X"21",X"70",X"38",X"01",X"03",X"0E",X"CD",X"93",X"07",X"3E",
		X"05",X"CD",X"CE",X"15",X"C1",X"10",X"E6",X"C9",X"3A",X"B9",X"87",X"B7",X"C0",X"3A",X"02",X"98",
		X"E6",X"08",X"28",X"07",X"3A",X"00",X"98",X"EE",X"10",X"18",X"03",X"3A",X"00",X"98",X"47",X"21",
		X"21",X"86",X"E6",X"0F",X"56",X"77",X"92",X"E6",X"0F",X"21",X"EA",X"80",X"CB",X"60",X"20",X"06",
		X"57",X"7E",X"92",X"C3",X"67",X"0E",X"86",X"77",X"CB",X"3F",X"E6",X"3F",X"32",X"22",X"86",X"C9",
		X"00",X"00",X"01",X"00",X"00",X"06",X"06",X"02",X"3F",X"07",X"06",X"06",X"02",X"3F",X"07",X"00",
		X"01",X"A8",X"87",X"00",X"00",X"01",X"00",X"00",X"01",X"00",X"01",X"3A",X"06",X"01",X"00",X"02",
		X"39",X"06",X"01",X"00",X"01",X"79",X"02",X"01",X"00",X"01",X"B8",X"02",X"01",X"00",X"01",X"38",
		X"03",X"01",X"00",X"01",X"77",X"03",X"01",X"00",X"01",X"B7",X"03",X"01",X"00",X"01",X"F7",X"03",
		X"00",X"00",X"CD",X"96",X"14",X"DD",X"21",X"15",X"82",X"FD",X"21",X"34",X"81",X"DD",X"36",X"08",
		X"6C",X"DD",X"36",X"0A",X"80",X"CD",X"04",X"11",X"3A",X"B9",X"87",X"B7",X"C4",X"26",X"11",X"DD",
		X"CB",X"00",X"D6",X"3E",X"06",X"32",X"23",X"86",X"3E",X"06",X"32",X"24",X"86",X"DD",X"CB",X"0C",
		X"CE",X"DD",X"CB",X"00",X"F6",X"CD",X"7A",X"15",X"01",X"FF",X"00",X"FD",X"21",X"34",X"81",X"FD",
		X"CB",X"00",X"76",X"C2",X"2B",X"11",X"3A",X"8E",X"87",X"B7",X"20",X"1B",X"DD",X"7E",X"0D",X"B7",
		X"CA",X"17",X"0F",X"CB",X"77",X"C2",X"17",X"0F",X"CB",X"6F",X"C2",X"2B",X"11",X"CB",X"67",X"C2",
		X"2B",X"11",X"CB",X"7F",X"C2",X"2B",X"11",X"DD",X"36",X"0D",X"00",X"2A",X"C5",X"80",X"22",X"5D",
		X"87",X"CD",X"54",X"10",X"E5",X"CB",X"61",X"C4",X"57",X"0F",X"CB",X"71",X"C4",X"C1",X"0F",X"CB",
		X"71",X"CC",X"63",X"0F",X"CB",X"79",X"C5",X"C4",X"AC",X"0F",X"C1",X"CB",X"69",X"CC",X"A6",X"0F",
		X"CB",X"69",X"C4",X"8E",X"0F",X"3A",X"B9",X"87",X"B7",X"28",X"05",X"3E",X"01",X"CD",X"CE",X"15",
		X"CD",X"7A",X"15",X"C1",X"C3",X"EB",X"0E",X"3A",X"EA",X"80",X"C6",X"40",X"30",X"01",X"3D",X"32",
		X"EA",X"80",X"C9",X"C5",X"CD",X"72",X"11",X"CD",X"80",X"0F",X"21",X"37",X"81",X"CD",X"1B",X"10",
		X"21",X"3F",X"81",X"CD",X"1B",X"10",X"CD",X"C0",X"10",X"3E",X"00",X"32",X"BF",X"87",X"C1",X"C9",
		X"AF",X"FD",X"77",X"01",X"FD",X"77",X"02",X"FD",X"77",X"09",X"FD",X"77",X"0A",X"C9",X"3A",X"5A",
		X"87",X"B7",X"28",X"12",X"3A",X"8E",X"87",X"B7",X"C0",X"3E",X"FF",X"32",X"8E",X"87",X"FD",X"21",
		X"4B",X"2B",X"CD",X"62",X"15",X"C9",X"3E",X"00",X"32",X"8E",X"87",X"C9",X"DD",X"7E",X"03",X"B7",
		X"C0",X"3A",X"7F",X"87",X"FE",X"03",X"D0",X"06",X"00",X"FD",X"21",X"47",X"1A",X"CD",X"62",X"15",
		X"C9",X"C5",X"CD",X"67",X"11",X"3A",X"22",X"86",X"E6",X"3F",X"CB",X"27",X"5F",X"16",X"00",X"21",
		X"12",X"1B",X"19",X"19",X"5E",X"23",X"56",X"06",X"05",X"CB",X"2A",X"CB",X"1B",X"10",X"FA",X"FD",
		X"73",X"01",X"FD",X"72",X"02",X"23",X"5E",X"23",X"56",X"06",X"05",X"CB",X"2A",X"CB",X"1B",X"10",
		X"FA",X"FD",X"73",X"09",X"FD",X"72",X"0A",X"2A",X"35",X"81",X"ED",X"5B",X"37",X"81",X"CD",X"35",
		X"10",X"22",X"35",X"81",X"2A",X"3D",X"81",X"ED",X"5B",X"3F",X"81",X"CD",X"35",X"10",X"22",X"3D",
		X"81",X"CD",X"B5",X"10",X"3E",X"FF",X"32",X"BF",X"87",X"C1",X"C9",X"5E",X"23",X"56",X"7A",X"B3",
		X"C8",X"EB",X"01",X"FE",X"FF",X"CB",X"7C",X"28",X"03",X"01",X"02",X"00",X"09",X"CD",X"49",X"10",
		X"EB",X"72",X"2B",X"73",X"C9",X"CD",X"F5",X"22",X"06",X"04",X"3A",X"58",X"87",X"B7",X"20",X"01",
		X"05",X"CB",X"2A",X"CB",X"1B",X"10",X"FA",X"19",X"C9",X"7C",X"B7",X"C0",X"7D",X"E6",X"F0",X"C0",
		X"21",X"00",X"00",X"C9",X"3A",X"B9",X"87",X"B7",X"20",X"46",X"3A",X"43",X"87",X"FE",X"02",X"20",
		X"27",X"3A",X"02",X"98",X"E6",X"08",X"28",X"20",X"06",X"00",X"3A",X"00",X"98",X"CB",X"6F",X"20",
		X"02",X"CB",X"E8",X"3A",X"01",X"98",X"CB",X"67",X"20",X"02",X"CB",X"F0",X"3A",X"02",X"98",X"CB",
		X"47",X"20",X"02",X"CB",X"F8",X"78",X"18",X"10",X"3A",X"01",X"98",X"2F",X"47",X"3A",X"02",X"98",
		X"CB",X"5F",X"78",X"28",X"03",X"47",X"E6",X"EF",X"57",X"A9",X"F6",X"E0",X"A2",X"6A",X"4F",X"C9",
		X"FD",X"7E",X"04",X"FD",X"B6",X"0C",X"20",X"03",X"0E",X"00",X"C9",X"0E",X"E0",X"06",X"00",X"3E",
		X"10",X"32",X"22",X"86",X"C9",X"21",X"7D",X"11",X"3A",X"BF",X"87",X"B7",X"28",X"16",X"18",X"09",
		X"21",X"FD",X"11",X"3A",X"BF",X"87",X"B7",X"20",X"0B",X"3A",X"B8",X"87",X"47",X"3A",X"22",X"86",
		X"E6",X"3F",X"B8",X"C8",X"3A",X"22",X"86",X"32",X"B8",X"87",X"16",X"00",X"5F",X"19",X"19",X"4E",
		X"23",X"46",X"DD",X"CB",X"00",X"A6",X"DD",X"E5",X"DD",X"21",X"A3",X"87",X"11",X"05",X"00",X"DD",
		X"19",X"DD",X"71",X"03",X"DD",X"19",X"DD",X"70",X"03",X"DD",X"E1",X"DD",X"36",X"04",X"01",X"DD",
		X"CB",X"00",X"E6",X"C9",X"21",X"70",X"0E",X"11",X"A3",X"87",X"01",X"14",X"00",X"ED",X"B0",X"21",
		X"A3",X"87",X"DD",X"75",X"05",X"DD",X"74",X"06",X"DD",X"36",X"04",X"01",X"DD",X"CB",X"00",X"E6",
		X"3E",X"20",X"32",X"EA",X"80",X"C9",X"FD",X"36",X"04",X"01",X"C9",X"3E",X"08",X"CD",X"F4",X"2B",
		X"CD",X"80",X"0F",X"CD",X"A6",X"0F",X"DD",X"CB",X"0B",X"C6",X"DD",X"CB",X"00",X"A6",X"21",X"83",
		X"0E",X"DD",X"75",X"05",X"DD",X"74",X"06",X"DD",X"36",X"04",X"01",X"DD",X"CB",X"00",X"E6",X"DD",
		X"CB",X"00",X"66",X"28",X"05",X"CD",X"7A",X"15",X"18",X"F5",X"3E",X"19",X"32",X"7D",X"87",X"CD",
		X"F4",X"15",X"CD",X"7A",X"15",X"18",X"FB",X"3A",X"00",X"A0",X"FE",X"0F",X"C8",X"3E",X"0F",X"C3",
		X"F4",X"2B",X"3A",X"00",X"A0",X"FE",X"0E",X"C8",X"3E",X"0E",X"C3",X"F4",X"2B",X"13",X"18",X"13",
		X"18",X"14",X"19",X"14",X"19",X"14",X"19",X"14",X"19",X"15",X"1A",X"15",X"1A",X"15",X"1A",X"15",
		X"1A",X"16",X"1B",X"16",X"1B",X"16",X"1B",X"16",X"1B",X"17",X"1C",X"17",X"1C",X"17",X"1C",X"17",
		X"1C",X"56",X"5B",X"56",X"5B",X"56",X"5B",X"56",X"5B",X"55",X"5A",X"55",X"5A",X"55",X"5A",X"55",
		X"5A",X"54",X"59",X"54",X"59",X"54",X"59",X"54",X"59",X"53",X"58",X"53",X"58",X"53",X"58",X"53",
		X"58",X"D4",X"D9",X"D4",X"D9",X"D4",X"D9",X"D4",X"D9",X"D5",X"DA",X"D5",X"DA",X"D5",X"DA",X"D5",
		X"DA",X"D6",X"DB",X"D6",X"DB",X"D6",X"DB",X"D6",X"DB",X"D7",X"DC",X"D7",X"DC",X"D7",X"DC",X"D7",
		X"DC",X"96",X"9B",X"96",X"9B",X"96",X"9B",X"96",X"9B",X"95",X"9A",X"95",X"9A",X"95",X"9A",X"95",
		X"9A",X"94",X"99",X"94",X"99",X"94",X"99",X"94",X"99",X"93",X"98",X"93",X"98",X"3B",X"3B",X"3B",
		X"3B",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3D",X"3D",X"3D",X"3D",X"3D",X"3D",X"3D",
		X"3D",X"3E",X"3E",X"3E",X"3E",X"3E",X"3E",X"3E",X"3E",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",
		X"7D",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",
		X"7B",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",
		X"FD",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BD",X"BD",X"BD",X"BD",X"BD",X"BD",X"BD",
		X"BD",X"BC",X"BC",X"BC",X"BC",X"BC",X"BC",X"BC",X"BC",X"3B",X"3B",X"3B",X"3B",X"CD",X"E6",X"13",
		X"0E",X"0A",X"11",X"F2",X"80",X"E5",X"D5",X"06",X"03",X"1A",X"BE",X"38",X"11",X"20",X"04",X"13",
		X"23",X"10",X"F6",X"D1",X"21",X"06",X"00",X"19",X"EB",X"E1",X"0D",X"20",X"E8",X"C9",X"D1",X"D5",
		X"CD",X"1E",X"14",X"0D",X"28",X"16",X"06",X"00",X"21",X"00",X"00",X"09",X"29",X"09",X"29",X"E5",
		X"19",X"2B",X"54",X"5D",X"01",X"06",X"00",X"09",X"EB",X"C1",X"ED",X"B8",X"D1",X"E1",X"01",X"03",
		X"00",X"ED",X"B0",X"D5",X"CD",X"61",X"07",X"CD",X"00",X"0D",X"CD",X"9E",X"0B",X"DF",X"1A",X"CF",
		X"20",X"28",X"43",X"4F",X"4E",X"47",X"52",X"41",X"54",X"55",X"4C",X"41",X"54",X"49",X"4F",X"4E",
		X"53",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"00",X"21",X"28",X"D8",X"11",X"43",X"87",X"06",
		X"01",X"CD",X"06",X"07",X"E7",X"0F",X"07",X"04",X"CF",X"28",X"38",X"59",X"4F",X"55",X"20",X"20",
		X"48",X"41",X"56",X"45",X"20",X"20",X"4A",X"4F",X"49",X"4E",X"45",X"44",X"20",X"20",X"54",X"48",
		X"45",X"00",X"CF",X"18",X"48",X"41",X"53",X"54",X"52",X"4F",X"4E",X"41",X"55",X"54",X"53",X"20",
		X"49",X"4E",X"20",X"54",X"48",X"45",X"20",X"4D",X"4F",X"4F",X"4E",X"20",X"57",X"41",X"52",X"00",
		X"CF",X"50",X"58",X"48",X"41",X"4C",X"4C",X"20",X"4F",X"46",X"20",X"46",X"41",X"4D",X"45",X"00",
		X"E7",X"03",X"0F",X"05",X"CF",X"28",X"78",X"45",X"4E",X"54",X"45",X"52",X"20",X"59",X"4F",X"55",
		X"52",X"20",X"49",X"4E",X"49",X"54",X"49",X"41",X"4C",X"53",X"20",X"5B",X"00",X"CF",X"70",X"88",
		X"5B",X"5B",X"5B",X"00",X"E7",X"03",X"16",X"07",X"CF",X"10",X"B0",X"4D",X"4F",X"56",X"45",X"20",
		X"57",X"48",X"45",X"45",X"4C",X"20",X"54",X"4F",X"20",X"43",X"48",X"41",X"4E",X"47",X"45",X"20",
		X"4C",X"45",X"54",X"54",X"45",X"52",X"00",X"CF",X"18",X"C0",X"50",X"52",X"45",X"53",X"53",X"20",
		X"53",X"48",X"49",X"45",X"4C",X"44",X"53",X"20",X"54",X"4F",X"20",X"53",X"54",X"4F",X"52",X"45",
		X"20",X"49",X"54",X"00",X"E1",X"E5",X"06",X"03",X"36",X"20",X"23",X"10",X"FB",X"21",X"88",X"70",
		X"CD",X"B8",X"06",X"D1",X"06",X"03",X"0E",X"41",X"3E",X"FF",X"32",X"44",X"87",X"CD",X"F3",X"13",
		X"20",X"FB",X"79",X"E5",X"CD",X"49",X"07",X"CD",X"0F",X"14",X"E1",X"3A",X"44",X"87",X"3D",X"32",
		X"44",X"87",X"C8",X"CD",X"F3",X"13",X"20",X"05",X"CD",X"00",X"14",X"18",X"E0",X"79",X"12",X"13",
		X"CD",X"49",X"07",X"10",X"D3",X"C9",X"3A",X"43",X"87",X"FE",X"02",X"21",X"31",X"81",X"C8",X"21",
		X"2E",X"81",X"C9",X"C5",X"D5",X"E5",X"CD",X"54",X"10",X"78",X"E6",X"20",X"E1",X"D1",X"C1",X"C9",
		X"3A",X"22",X"86",X"E6",X"1F",X"C6",X"41",X"FE",X"5B",X"38",X"02",X"3E",X"20",X"4F",X"C9",X"D5",
		X"C5",X"3E",X"03",X"F5",X"CD",X"C5",X"18",X"F1",X"3D",X"20",X"F8",X"C1",X"D1",X"C9",X"79",X"FE",
		X"0A",X"3E",X"01",X"CA",X"F4",X"2B",X"3E",X"02",X"C3",X"F4",X"2B",X"C2",X"31",X"68",X"80",X"CD",
		X"54",X"16",X"CD",X"63",X"14",X"CD",X"50",X"14",X"CD",X"9F",X"05",X"CD",X"92",X"18",X"CD",X"2A",
		X"06",X"CD",X"92",X"18",X"CD",X"5F",X"1C",X"CD",X"92",X"18",X"CD",X"40",X"18",X"C3",X"32",X"14",
		X"3A",X"01",X"98",X"2F",X"E6",X"03",X"C0",X"3E",X"99",X"32",X"F1",X"80",X"C9",X"CD",X"63",X"14",
		X"CD",X"F3",X"18",X"E1",X"22",X"0B",X"86",X"32",X"0D",X"86",X"CD",X"27",X"16",X"CD",X"80",X"14",
		X"AF",X"32",X"26",X"86",X"3E",X"FF",X"32",X"01",X"A8",X"2A",X"0B",X"86",X"3A",X"0D",X"86",X"E9",
		X"FD",X"E1",X"DD",X"21",X"43",X"82",X"DD",X"CB",X"00",X"C6",X"DD",X"CB",X"00",X"CE",X"CD",X"3E",
		X"15",X"31",X"90",X"80",X"FD",X"E9",X"FD",X"E1",X"DD",X"21",X"15",X"82",X"DD",X"CB",X"00",X"C6",
		X"DD",X"CB",X"00",X"CE",X"CD",X"3E",X"15",X"31",X"B8",X"80",X"DD",X"21",X"34",X"81",X"DD",X"CB",
		X"00",X"C6",X"CD",X"27",X"15",X"CD",X"52",X"15",X"FD",X"E9",X"D9",X"21",X"75",X"16",X"CD",X"0C",
		X"15",X"D9",X"D0",X"CD",X"27",X"15",X"CD",X"52",X"15",X"37",X"C9",X"D9",X"21",X"85",X"16",X"CD",
		X"0C",X"15",X"D9",X"D0",X"CD",X"27",X"15",X"CD",X"52",X"15",X"37",X"C9",X"E1",X"D9",X"21",X"95",
		X"16",X"CD",X"0C",X"15",X"D9",X"D2",X"F3",X"14",X"DD",X"22",X"BA",X"80",X"CD",X"3E",X"15",X"CD",
		X"E7",X"15",X"37",X"E9",X"E1",X"D9",X"21",X"69",X"16",X"C3",X"E1",X"14",X"E1",X"D9",X"21",X"5F",
		X"16",X"C3",X"E1",X"14",X"E1",X"D9",X"21",X"71",X"16",X"C3",X"E1",X"14",X"E5",X"D1",X"7E",X"23",
		X"66",X"6F",X"B4",X"C8",X"7E",X"B7",X"28",X"06",X"13",X"13",X"D5",X"E1",X"18",X"F0",X"E5",X"DD",
		X"E1",X"DD",X"CB",X"00",X"C6",X"37",X"C9",X"D9",X"DD",X"E5",X"E1",X"DD",X"2A",X"BA",X"80",X"DD",
		X"75",X"01",X"DD",X"74",X"02",X"DD",X"CB",X"00",X"DE",X"E5",X"DD",X"E1",X"D9",X"C9",X"D9",X"DD",
		X"CB",X"00",X"CE",X"DD",X"E5",X"E1",X"22",X"BA",X"80",X"AF",X"06",X"0F",X"23",X"77",X"10",X"FC",
		X"D9",X"C9",X"D9",X"DD",X"E5",X"E1",X"22",X"B8",X"80",X"AF",X"06",X"0E",X"23",X"77",X"10",X"FC",
		X"D9",X"C9",X"21",X"00",X"00",X"39",X"31",X"68",X"80",X"FD",X"E5",X"FD",X"2A",X"BA",X"80",X"FD",
		X"22",X"BE",X"80",X"FD",X"75",X"0E",X"FD",X"74",X"0F",X"C9",X"21",X"00",X"00",X"39",X"31",X"68",
		X"80",X"DD",X"2A",X"BA",X"80",X"DD",X"75",X"0E",X"DD",X"74",X"0F",X"2A",X"BE",X"80",X"7C",X"B5",
		X"28",X"0C",X"DD",X"2A",X"BE",X"80",X"21",X"00",X"00",X"22",X"BE",X"80",X"18",X"04",X"DD",X"2A",
		X"BA",X"80",X"CD",X"B7",X"15",X"DD",X"CB",X"00",X"46",X"28",X"F7",X"DD",X"22",X"BA",X"80",X"DD",
		X"66",X"0F",X"DD",X"6E",X"0E",X"F9",X"C9",X"D9",X"01",X"2E",X"00",X"DD",X"09",X"DD",X"E5",X"E1",
		X"01",X"09",X"86",X"B7",X"ED",X"42",X"38",X"04",X"DD",X"21",X"15",X"82",X"D9",X"C9",X"DD",X"2A",
		X"BA",X"80",X"DD",X"77",X"03",X"DD",X"CB",X"00",X"EE",X"CD",X"7A",X"15",X"DD",X"2A",X"BA",X"80",
		X"DD",X"CB",X"00",X"6E",X"20",X"F3",X"C9",X"D9",X"D1",X"01",X"2E",X"00",X"DD",X"E5",X"E1",X"09",
		X"F9",X"D5",X"D9",X"C9",X"CD",X"04",X"16",X"D9",X"2A",X"BA",X"80",X"06",X"10",X"AF",X"77",X"23",
		X"10",X"FC",X"D9",X"C9",X"DD",X"2A",X"BA",X"80",X"DD",X"CB",X"00",X"5E",X"C8",X"DD",X"CB",X"00",
		X"9E",X"D9",X"DD",X"6E",X"01",X"DD",X"66",X"02",X"06",X"0F",X"AF",X"77",X"23",X"10",X"FC",X"DD",
		X"77",X"01",X"DD",X"77",X"01",X"D9",X"C9",X"CD",X"43",X"3E",X"DD",X"21",X"15",X"82",X"AF",X"DD",
		X"77",X"00",X"DD",X"21",X"71",X"82",X"DD",X"77",X"00",X"CD",X"B7",X"15",X"30",X"02",X"18",X"F6",
		X"DD",X"21",X"34",X"81",X"11",X"0F",X"00",X"06",X"0F",X"DD",X"77",X"00",X"DD",X"19",X"10",X"F9",
		X"CD",X"49",X"3E",X"C9",X"D9",X"21",X"00",X"50",X"0E",X"01",X"CD",X"88",X"07",X"D9",X"C9",X"C7",
		X"84",X"F5",X"84",X"23",X"85",X"51",X"85",X"00",X"00",X"7F",X"85",X"AD",X"85",X"DB",X"85",X"00",
		X"00",X"99",X"84",X"00",X"00",X"43",X"81",X"52",X"81",X"61",X"81",X"70",X"81",X"7F",X"81",X"8E",
		X"81",X"9D",X"81",X"00",X"00",X"AC",X"81",X"BB",X"81",X"CA",X"81",X"D9",X"81",X"E8",X"81",X"F7",
		X"81",X"06",X"82",X"00",X"00",X"71",X"82",X"9F",X"82",X"CD",X"82",X"FB",X"82",X"29",X"83",X"57",
		X"83",X"85",X"83",X"B3",X"83",X"E1",X"83",X"0F",X"84",X"3D",X"84",X"6B",X"84",X"00",X"00",X"DD",
		X"21",X"15",X"82",X"FD",X"21",X"71",X"82",X"3A",X"24",X"86",X"6F",X"DD",X"4E",X"0A",X"D9",X"3A",
		X"23",X"86",X"6F",X"DD",X"4E",X"08",X"06",X"0D",X"FD",X"7E",X"00",X"E6",X"41",X"EE",X"41",X"20",
		X"37",X"FD",X"56",X"06",X"FD",X"5E",X"05",X"1A",X"67",X"13",X"1A",X"D9",X"85",X"1F",X"67",X"FD",
		X"7E",X"0A",X"91",X"30",X"02",X"ED",X"44",X"BC",X"D9",X"30",X"1D",X"7C",X"85",X"1F",X"67",X"FD",
		X"7E",X"08",X"91",X"30",X"02",X"ED",X"44",X"BC",X"30",X"0E",X"DD",X"7E",X"0D",X"FD",X"56",X"0C",
		X"B2",X"DD",X"77",X"0D",X"FD",X"CB",X"0D",X"CE",X"11",X"2E",X"00",X"FD",X"19",X"10",X"B9",X"FD",
		X"21",X"C7",X"84",X"06",X"04",X"FD",X"7E",X"00",X"E6",X"41",X"EE",X"41",X"20",X"26",X"65",X"CB",
		X"3C",X"FD",X"7E",X"08",X"91",X"30",X"02",X"ED",X"44",X"BC",X"30",X"18",X"D9",X"65",X"CB",X"3C",
		X"FD",X"7E",X"0A",X"91",X"30",X"02",X"ED",X"44",X"BC",X"D9",X"30",X"08",X"FD",X"CB",X"0D",X"CE",
		X"DD",X"CB",X"0D",X"E6",X"11",X"2E",X"00",X"FD",X"19",X"10",X"CA",X"21",X"89",X"85",X"4E",X"21",
		X"B7",X"85",X"7E",X"21",X"E5",X"85",X"6E",X"67",X"D9",X"21",X"87",X"85",X"4E",X"21",X"B5",X"85",
		X"7E",X"21",X"E3",X"85",X"6E",X"67",X"06",X"0D",X"FD",X"21",X"71",X"82",X"FD",X"7E",X"00",X"E6",
		X"41",X"EE",X"41",X"20",X"74",X"FD",X"56",X"06",X"FD",X"5E",X"05",X"1A",X"08",X"13",X"1A",X"D9",
		X"CB",X"3F",X"5F",X"FD",X"7E",X"0A",X"57",X"91",X"30",X"02",X"ED",X"44",X"BB",X"08",X"D9",X"CB",
		X"3F",X"5F",X"FD",X"7E",X"08",X"57",X"91",X"30",X"02",X"ED",X"44",X"BB",X"30",X"0A",X"08",X"30",
		X"07",X"DD",X"21",X"7F",X"85",X"C3",X"DB",X"17",X"D9",X"7A",X"94",X"30",X"02",X"ED",X"44",X"BB",
		X"D9",X"30",X"10",X"7A",X"94",X"30",X"02",X"ED",X"44",X"BB",X"30",X"07",X"DD",X"21",X"AD",X"85",
		X"C3",X"DB",X"17",X"D9",X"7A",X"95",X"30",X"02",X"ED",X"44",X"BB",X"D9",X"30",X"1B",X"7A",X"95",
		X"30",X"02",X"ED",X"44",X"BB",X"30",X"12",X"DD",X"21",X"DB",X"85",X"DD",X"7E",X"0D",X"FD",X"56",
		X"0C",X"B2",X"DD",X"77",X"0D",X"FD",X"CB",X"0D",X"D6",X"11",X"2E",X"00",X"FD",X"19",X"05",X"C2",
		X"6C",X"17",X"DD",X"21",X"99",X"84",X"FD",X"21",X"C7",X"84",X"3E",X"0E",X"6F",X"DD",X"4E",X"0A",
		X"D9",X"3E",X"0E",X"6F",X"DD",X"4E",X"08",X"06",X"04",X"FD",X"7E",X"00",X"E6",X"41",X"EE",X"41",
		X"20",X"26",X"65",X"CB",X"3C",X"FD",X"7E",X"08",X"91",X"30",X"02",X"ED",X"44",X"BC",X"30",X"18",
		X"D9",X"65",X"CB",X"3C",X"FD",X"7E",X"0A",X"91",X"30",X"02",X"ED",X"44",X"BC",X"D9",X"30",X"08",
		X"FD",X"CB",X"0D",X"F6",X"DD",X"CB",X"0D",X"E6",X"11",X"2E",X"00",X"FD",X"19",X"10",X"CA",X"C9",
		X"3E",X"FF",X"32",X"B9",X"87",X"3E",X"00",X"CD",X"F4",X"2B",X"21",X"43",X"87",X"36",X"01",X"23",
		X"36",X"01",X"23",X"23",X"36",X"01",X"3E",X"01",X"32",X"5C",X"87",X"32",X"C6",X"80",X"3E",X"09",
		X"32",X"46",X"87",X"21",X"80",X"04",X"22",X"BD",X"87",X"3E",X"99",X"32",X"5A",X"87",X"3E",X"36",
		X"32",X"58",X"87",X"AF",X"32",X"7D",X"87",X"32",X"7E",X"87",X"32",X"7F",X"87",X"32",X"1B",X"86",
		X"32",X"BF",X"87",X"CD",X"43",X"0D",X"3E",X"1E",X"CD",X"CE",X"15",X"CD",X"27",X"16",X"CD",X"6E",
		X"21",X"C9",X"0E",X"04",X"DD",X"2A",X"BA",X"80",X"DD",X"CB",X"00",X"EE",X"DD",X"36",X"03",X"1E",
		X"3A",X"F1",X"80",X"47",X"C5",X"CD",X"2A",X"19",X"C1",X"C5",X"3A",X"F1",X"80",X"B8",X"C4",X"68",
		X"0B",X"C1",X"CD",X"46",X"21",X"CD",X"C5",X"19",X"C2",X"5D",X"14",X"DD",X"CB",X"00",X"6E",X"20",
		X"DF",X"0D",X"20",X"D0",X"C9",X"DD",X"2A",X"BA",X"80",X"DD",X"CB",X"00",X"EE",X"DD",X"36",X"03",
		X"01",X"3A",X"F1",X"80",X"47",X"C5",X"CD",X"2A",X"19",X"C1",X"C5",X"3A",X"F1",X"80",X"B8",X"C4",
		X"68",X"0B",X"C1",X"CD",X"46",X"21",X"CD",X"C5",X"19",X"C2",X"5D",X"14",X"DD",X"CB",X"00",X"6E",
		X"20",X"DF",X"C9",X"47",X"CD",X"09",X"19",X"CB",X"58",X"3E",X"01",X"28",X"05",X"CD",X"09",X"19",
		X"3E",X"02",X"32",X"1E",X"86",X"E1",X"C3",X"29",X"0C",X"3A",X"F1",X"80",X"C6",X"99",X"27",X"32",
		X"F1",X"80",X"C9",X"47",X"B7",X"C8",X"3A",X"F1",X"80",X"FE",X"99",X"C8",X"80",X"27",X"30",X"02",
		X"3E",X"99",X"32",X"F1",X"80",X"3E",X"05",X"C3",X"F4",X"2B",X"11",X"ED",X"80",X"3A",X"EF",X"80",
		X"4F",X"21",X"DD",X"19",X"CD",X"53",X"19",X"CD",X"13",X"19",X"79",X"32",X"EF",X"80",X"11",X"EE",
		X"80",X"3A",X"F0",X"80",X"4F",X"21",X"0D",X"1A",X"CD",X"53",X"19",X"CD",X"13",X"19",X"79",X"32",
		X"F0",X"80",X"C9",X"3A",X"02",X"98",X"2F",X"E6",X"06",X"CB",X"3F",X"47",X"28",X"08",X"D5",X"11",
		X"0C",X"00",X"19",X"10",X"FD",X"D1",X"1A",X"B7",X"C8",X"09",X"AF",X"86",X"08",X"79",X"FE",X"0B",
		X"20",X"0B",X"D5",X"11",X"0C",X"00",X"AF",X"ED",X"52",X"4F",X"D1",X"18",X"02",X"0C",X"23",X"08",
		X"EB",X"35",X"CD",X"89",X"19",X"EB",X"20",X"E3",X"C9",X"F5",X"C5",X"D5",X"E5",X"3E",X"FF",X"32",
		X"02",X"A8",X"3E",X"03",X"CD",X"CE",X"15",X"3E",X"00",X"32",X"02",X"A8",X"3E",X"0C",X"CD",X"CE",
		X"15",X"E1",X"D1",X"C1",X"F1",X"C9",X"21",X"EB",X"80",X"7E",X"23",X"46",X"A8",X"4F",X"3A",X"00",
		X"98",X"2F",X"77",X"2B",X"70",X"A1",X"E6",X"C0",X"23",X"23",X"CB",X"7F",X"28",X"01",X"34",X"23",
		X"CB",X"77",X"C8",X"34",X"C9",X"C5",X"06",X"00",X"3A",X"F1",X"80",X"B7",X"28",X"08",X"FE",X"01",
		X"06",X"04",X"28",X"02",X"06",X"0C",X"3A",X"01",X"98",X"2F",X"A0",X"C1",X"C9",X"04",X"04",X"04",
		X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"03",X"03",X"03",X"03",X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"01",X"00",X"00",X"01",X"00",
		X"00",X"01",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"01",
		X"00",X"00",X"01",X"02",X"00",X"00",X"00",X"CD",X"F4",X"14",X"D2",X"9E",X"15",X"DD",X"E5",X"CD",
		X"CB",X"14",X"D2",X"EE",X"1A",X"FD",X"E1",X"21",X"7F",X"87",X"34",X"CD",X"0E",X"2C",X"CD",X"FA",
		X"1A",X"DD",X"E5",X"DD",X"21",X"15",X"82",X"DD",X"36",X"03",X"04",X"DD",X"CB",X"00",X"EE",X"DD",
		X"7E",X"08",X"FD",X"77",X"08",X"DD",X"7E",X"0A",X"FD",X"77",X"0A",X"DD",X"21",X"34",X"81",X"D5",
		X"DD",X"56",X"0C",X"DD",X"5E",X"0B",X"19",X"D1",X"E5",X"EB",X"DD",X"56",X"04",X"DD",X"5E",X"03",
		X"19",X"D1",X"DD",X"E1",X"DD",X"72",X"0C",X"DD",X"73",X"0B",X"DD",X"74",X"04",X"DD",X"75",X"03",
		X"FD",X"CB",X"0C",X"D6",X"3E",X"14",X"FD",X"77",X"03",X"FD",X"CB",X"00",X"EE",X"FD",X"CB",X"00",
		X"F6",X"FD",X"CB",X"00",X"D6",X"21",X"3D",X"1A",X"FD",X"75",X"05",X"FD",X"74",X"06",X"DD",X"E5",
		X"CD",X"7A",X"15",X"FD",X"E1",X"DD",X"CB",X"00",X"4E",X"CA",X"EE",X"1A",X"DD",X"7E",X"0D",X"B7",
		X"28",X"04",X"CB",X"77",X"28",X"18",X"DD",X"36",X"0D",X"00",X"DD",X"CB",X"00",X"6E",X"28",X"0E",
		X"FD",X"CB",X"00",X"76",X"C2",X"EE",X"1A",X"FD",X"E5",X"CD",X"7A",X"15",X"18",X"D5",X"21",X"7F",
		X"87",X"35",X"CD",X"F4",X"15",X"CD",X"7A",X"15",X"18",X"FB",X"3A",X"22",X"86",X"E6",X"3F",X"CB",
		X"27",X"5F",X"16",X"00",X"21",X"12",X"1B",X"19",X"19",X"5E",X"23",X"56",X"23",X"7E",X"23",X"66",
		X"6F",X"C9",X"00",X"00",X"AB",X"FA",X"85",X"00",X"B2",X"FA",X"0A",X"01",X"C5",X"FA",X"8C",X"01",
		X"E6",X"FA",X"0A",X"02",X"13",X"FB",X"83",X"02",X"4C",X"FB",X"F6",X"02",X"91",X"FB",X"62",X"03",
		X"E1",X"FB",X"C5",X"03",X"3B",X"FC",X"1F",X"04",X"9E",X"FC",X"6F",X"04",X"0A",X"FD",X"B4",X"04",
		X"7D",X"FD",X"ED",X"04",X"F6",X"FD",X"1A",X"05",X"74",X"FE",X"3B",X"05",X"F6",X"FE",X"4E",X"05",
		X"7B",X"FF",X"55",X"05",X"00",X"00",X"4E",X"05",X"85",X"00",X"3B",X"05",X"0A",X"01",X"1A",X"05",
		X"8C",X"01",X"ED",X"04",X"0A",X"02",X"B4",X"04",X"83",X"02",X"6F",X"04",X"F6",X"02",X"1F",X"04",
		X"62",X"03",X"C5",X"03",X"C5",X"03",X"62",X"03",X"1F",X"04",X"F6",X"02",X"6F",X"04",X"83",X"02",
		X"B4",X"04",X"0A",X"02",X"ED",X"04",X"8C",X"01",X"1A",X"05",X"03",X"01",X"3B",X"05",X"85",X"00",
		X"4E",X"05",X"00",X"00",X"55",X"05",X"7B",X"FF",X"4E",X"05",X"F6",X"FE",X"3B",X"05",X"74",X"FE",
		X"1A",X"05",X"F6",X"FD",X"ED",X"04",X"7D",X"FD",X"B4",X"04",X"0A",X"FD",X"6F",X"04",X"9E",X"FC",
		X"1F",X"04",X"3B",X"FC",X"C5",X"03",X"E1",X"FB",X"62",X"03",X"91",X"FB",X"F6",X"02",X"4C",X"FB",
		X"83",X"02",X"13",X"FB",X"0A",X"02",X"E6",X"FA",X"8C",X"01",X"C5",X"FA",X"0A",X"01",X"B2",X"FA",
		X"85",X"00",X"AB",X"FA",X"00",X"00",X"B2",X"FA",X"7B",X"FF",X"C5",X"FA",X"F6",X"FE",X"E6",X"FA",
		X"74",X"FE",X"13",X"FB",X"F6",X"FD",X"4C",X"FB",X"7D",X"FD",X"91",X"FB",X"0A",X"FD",X"E1",X"FB",
		X"9E",X"FC",X"3B",X"FC",X"3B",X"FC",X"9E",X"FC",X"E1",X"FB",X"0A",X"FD",X"91",X"FB",X"7D",X"FD",
		X"4C",X"FB",X"F6",X"FD",X"13",X"FB",X"74",X"FE",X"E6",X"FA",X"F6",X"FE",X"C5",X"FA",X"7B",X"FF",
		X"B2",X"FA",X"E1",X"7E",X"23",X"E5",X"11",X"00",X"00",X"06",X"20",X"C3",X"3B",X"1C",X"E1",X"7E",
		X"23",X"E5",X"47",X"0F",X"0F",X"E6",X"3E",X"4F",X"78",X"06",X"00",X"21",X"01",X"90",X"09",X"77",
		X"C9",X"E1",X"46",X"23",X"5E",X"16",X"00",X"23",X"7E",X"23",X"E5",X"21",X"01",X"90",X"19",X"19",
		X"77",X"23",X"23",X"10",X"FB",X"C9",X"21",X"01",X"90",X"19",X"19",X"77",X"23",X"23",X"10",X"FB",
		X"C9",X"77",X"3C",X"23",X"77",X"3C",X"11",X"1F",X"00",X"19",X"77",X"3C",X"23",X"77",X"C9",X"CD",
		X"61",X"07",X"3E",X"00",X"32",X"07",X"A8",X"32",X"06",X"A8",X"3E",X"FF",X"32",X"04",X"A8",X"CD",
		X"46",X"0B",X"CD",X"68",X"0B",X"CD",X"9E",X"0B",X"DF",X"1A",X"CF",X"00",X"18",X"4D",X"4F",X"4F",
		X"4E",X"57",X"41",X"52",X"00",X"0E",X"00",X"06",X"60",X"0C",X"79",X"32",X"06",X"90",X"C5",X"CD",
		X"C5",X"18",X"C1",X"10",X"F4",X"0E",X"01",X"CD",X"94",X"18",X"E7",X"10",X"06",X"02",X"21",X"66",
		X"8B",X"3E",X"D0",X"CD",X"51",X"1C",X"CF",X"28",X"30",X"20",X"20",X"5B",X"20",X"20",X"52",X"45",
		X"46",X"55",X"45",X"4C",X"49",X"4E",X"47",X"20",X"42",X"41",X"53",X"45",X"00",X"0E",X"01",X"CD",
		X"94",X"18",X"21",X"68",X"8B",X"3E",X"34",X"CD",X"51",X"1C",X"CF",X"28",X"40",X"20",X"20",X"5B",
		X"20",X"20",X"53",X"41",X"54",X"45",X"4C",X"4C",X"49",X"54",X"45",X"20",X"5B",X"20",X"31",X"30",
		X"30",X"20",X"50",X"54",X"53",X"00",X"0E",X"01",X"CD",X"94",X"18",X"21",X"6A",X"8B",X"3E",X"B0",
		X"CD",X"51",X"1C",X"CF",X"28",X"50",X"20",X"20",X"5B",X"20",X"20",X"46",X"49",X"47",X"48",X"54",
		X"45",X"52",X"20",X"20",X"20",X"5B",X"20",X"31",X"35",X"30",X"20",X"50",X"54",X"53",X"00",X"0E",
		X"01",X"CD",X"94",X"18",X"21",X"6C",X"8B",X"3E",X"B8",X"CD",X"51",X"1C",X"CF",X"28",X"60",X"20",
		X"20",X"5B",X"20",X"20",X"42",X"4F",X"4D",X"42",X"45",X"52",X"20",X"20",X"20",X"20",X"5B",X"20",
		X"32",X"30",X"30",X"20",X"50",X"54",X"53",X"00",X"0E",X"01",X"CD",X"94",X"18",X"21",X"6E",X"8B",
		X"3E",X"BC",X"CD",X"51",X"1C",X"CF",X"28",X"70",X"20",X"20",X"5B",X"20",X"20",X"53",X"54",X"52",
		X"41",X"46",X"45",X"52",X"20",X"20",X"20",X"5B",X"20",X"33",X"30",X"30",X"20",X"50",X"54",X"53",
		X"00",X"0E",X"01",X"CD",X"94",X"18",X"21",X"70",X"8B",X"3E",X"7C",X"CD",X"51",X"1C",X"CF",X"28",
		X"80",X"20",X"20",X"5B",X"20",X"20",X"54",X"52",X"41",X"43",X"45",X"52",X"20",X"20",X"20",X"20",
		X"5B",X"20",X"35",X"30",X"30",X"20",X"50",X"54",X"53",X"00",X"0E",X"01",X"CD",X"94",X"18",X"21",
		X"72",X"8B",X"3E",X"74",X"CD",X"51",X"1C",X"CF",X"28",X"90",X"20",X"20",X"5B",X"20",X"20",X"41",
		X"57",X"41",X"52",X"44",X"53",X"20",X"42",X"4F",X"4E",X"55",X"53",X"20",X"53",X"48",X"49",X"50",
		X"00",X"0E",X"01",X"CD",X"94",X"18",X"AF",X"0E",X"60",X"06",X"80",X"3C",X"E6",X"07",X"0C",X"0C",
		X"08",X"79",X"32",X"06",X"90",X"08",X"F5",X"C5",X"11",X"06",X"00",X"06",X"0E",X"CD",X"46",X"1C",
		X"CD",X"C5",X"18",X"C1",X"F1",X"10",X"E4",X"E7",X"0E",X"06",X"02",X"0E",X"01",X"CD",X"94",X"18",
		X"C3",X"2A",X"06",X"21",X"80",X"87",X"06",X"08",X"34",X"23",X"10",X"FC",X"C9",X"C9",X"3A",X"7D",
		X"87",X"FE",X"05",X"D0",X"CD",X"6A",X"03",X"D8",X"3A",X"4A",X"87",X"CB",X"3F",X"3C",X"47",X"3A",
		X"7D",X"87",X"90",X"D0",X"21",X"96",X"87",X"36",X"00",X"23",X"CD",X"98",X"04",X"73",X"23",X"72",
		X"21",X"9C",X"87",X"CD",X"DF",X"2A",X"77",X"21",X"51",X"87",X"CD",X"46",X"21",X"BE",X"30",X"08",
		X"FD",X"21",X"20",X"36",X"CD",X"62",X"15",X"C9",X"23",X"BE",X"30",X"08",X"FD",X"21",X"BC",X"1F",
		X"CD",X"62",X"15",X"C9",X"23",X"BE",X"30",X"08",X"FD",X"21",X"40",X"34",X"CD",X"62",X"15",X"C9",
		X"FD",X"21",X"78",X"31",X"CD",X"62",X"15",X"C9",X"3A",X"1B",X"86",X"B7",X"C0",X"21",X"6B",X"1E",
		X"3A",X"46",X"87",X"BE",X"28",X"0B",X"3E",X"FF",X"BE",X"C8",X"11",X"12",X"00",X"19",X"C3",X"50",
		X"1E",X"23",X"01",X"11",X"00",X"11",X"47",X"87",X"ED",X"B0",X"C9",X"01",X"40",X"60",X"00",X"01",
		X"01",X"01",X"FF",X"01",X"01",X"06",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"02",X"30",X"80",
		X"00",X"02",X"01",X"01",X"FF",X"02",X"01",X"05",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"03",
		X"20",X"A0",X"00",X"03",X"03",X"02",X"7F",X"03",X"02",X"06",X"02",X"04",X"00",X"00",X"00",X"00",
		X"00",X"04",X"20",X"B0",X"00",X"04",X"03",X"02",X"7F",X"03",X"02",X"06",X"02",X"05",X"01",X"00",
		X"00",X"00",X"00",X"06",X"10",X"D0",X"00",X"05",X"03",X"03",X"3F",X"03",X"03",X"06",X"03",X"05",
		X"02",X"00",X"00",X"00",X"00",X"08",X"10",X"E0",X"00",X"05",X"03",X"04",X"3F",X"03",X"04",X"06",
		X"04",X"06",X"03",X"00",X"00",X"00",X"00",X"09",X"10",X"F0",X"00",X"05",X"03",X"04",X"3F",X"03",
		X"05",X"06",X"05",X"06",X"04",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"01",X"05",X"03",X"04",
		X"1F",X"03",X"05",X"08",X"06",X"08",X"05",X"00",X"00",X"00",X"00",X"15",X"10",X"50",X"01",X"05",
		X"03",X"04",X"1F",X"03",X"06",X"0A",X"07",X"0A",X"06",X"00",X"00",X"00",X"00",X"20",X"10",X"A0",
		X"01",X"05",X"03",X"04",X"0F",X"03",X"07",X"0A",X"08",X"0C",X"07",X"00",X"00",X"00",X"00",X"30",
		X"10",X"F0",X"01",X"05",X"03",X"04",X"0F",X"03",X"08",X"0C",X"07",X"0F",X"06",X"00",X"00",X"00",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3A",X"4C",X"87",X"47",X"3A",X"7E",
		X"87",X"B8",X"D0",X"DD",X"7E",X"08",X"FE",X"09",X"38",X"06",X"FE",X"F1",X"30",X"02",X"37",X"C9",
		X"B7",X"C9",X"00",X"00",X"01",X"00",X"00",X"0A",X"0A",X"05",X"0D",X"06",X"0A",X"0A",X"05",X"0E",
		X"06",X"0A",X"0A",X"05",X"0F",X"06",X"0A",X"0A",X"05",X"10",X"06",X"0A",X"0A",X"05",X"0D",X"07",
		X"0A",X"0A",X"05",X"0E",X"07",X"0A",X"0A",X"05",X"0F",X"07",X"0A",X"0A",X"05",X"10",X"07",X"00",
		X"01",X"57",X"1F",X"00",X"00",X"01",X"00",X"00",X"0C",X"0A",X"03",X"6D",X"06",X"0C",X"0A",X"01",
		X"6D",X"07",X"00",X"01",X"88",X"1F",X"00",X"00",X"01",X"00",X"00",X"0C",X"0A",X"03",X"AD",X"06",
		X"0C",X"0A",X"01",X"AD",X"07",X"00",X"01",X"9B",X"1F",X"00",X"00",X"01",X"00",X"00",X"0C",X"0A",
		X"03",X"ED",X"06",X"0C",X"0A",X"01",X"ED",X"07",X"00",X"01",X"AE",X"1F",X"CD",X"DC",X"14",X"D2",
		X"9E",X"15",X"21",X"7D",X"87",X"34",X"CD",X"BA",X"14",X"D2",X"9B",X"20",X"DD",X"E5",X"FD",X"E1",
		X"DD",X"2A",X"BA",X"80",X"CD",X"A7",X"20",X"CD",X"D2",X"20",X"CD",X"BC",X"20",X"CD",X"37",X"21",
		X"DD",X"77",X"03",X"DD",X"CB",X"00",X"EE",X"DD",X"CB",X"00",X"F6",X"DD",X"CB",X"0C",X"EE",X"DD",
		X"36",X"0B",X"03",X"DD",X"CB",X"00",X"D6",X"3E",X"02",X"CD",X"3A",X"3E",X"FD",X"E5",X"CD",X"7A",
		X"15",X"FD",X"E1",X"DD",X"CB",X"00",X"4E",X"CA",X"9B",X"20",X"DD",X"7E",X"0D",X"B7",X"20",X"38",
		X"FD",X"CB",X"00",X"76",X"CA",X"1E",X"20",X"CD",X"D2",X"20",X"FD",X"CB",X"00",X"B6",X"CD",X"1B",
		X"23",X"FD",X"E5",X"DD",X"CB",X"00",X"6E",X"20",X"1A",X"CD",X"3A",X"1F",X"30",X"15",X"CD",X"37",
		X"21",X"DD",X"77",X"03",X"DD",X"CB",X"00",X"EE",X"DD",X"22",X"88",X"87",X"FD",X"21",X"D8",X"21",
		X"CD",X"62",X"15",X"CD",X"7A",X"15",X"18",X"B9",X"CD",X"16",X"2C",X"FD",X"E5",X"E1",X"E5",X"11",
		X"01",X"00",X"19",X"AF",X"06",X"04",X"77",X"23",X"10",X"FC",X"E1",X"11",X"09",X"00",X"19",X"06",
		X"05",X"77",X"23",X"10",X"FC",X"DD",X"CB",X"0C",X"AE",X"DD",X"CB",X"00",X"A6",X"21",X"83",X"0E",
		X"DD",X"75",X"05",X"DD",X"74",X"06",X"DD",X"36",X"04",X"01",X"DD",X"CB",X"00",X"E6",X"06",X"02",
		X"0E",X"01",X"CD",X"8B",X"21",X"3E",X"02",X"CD",X"31",X"3E",X"DD",X"CB",X"00",X"66",X"28",X"0B",
		X"DD",X"CB",X"00",X"4E",X"28",X"05",X"CD",X"7A",X"15",X"18",X"EF",X"21",X"7D",X"87",X"35",X"CD",
		X"F4",X"15",X"CD",X"7A",X"15",X"18",X"FB",X"CD",X"46",X"21",X"FE",X"20",X"38",X"F9",X"FE",X"E8",
		X"30",X"F5",X"47",X"3E",X"EF",X"DD",X"77",X"08",X"DD",X"70",X"0A",X"C9",X"DD",X"CB",X"00",X"A6",
		X"21",X"52",X"1F",X"DD",X"75",X"05",X"DD",X"74",X"06",X"DD",X"36",X"04",X"01",X"DD",X"CB",X"00",
		X"E6",X"C9",X"FD",X"E5",X"FD",X"21",X"34",X"81",X"26",X"00",X"FD",X"6E",X"06",X"16",X"00",X"DD",
		X"5E",X"08",X"ED",X"52",X"3A",X"4E",X"87",X"47",X"CB",X"25",X"CB",X"14",X"10",X"FA",X"CD",X"24",
		X"21",X"ED",X"4B",X"37",X"81",X"09",X"EB",X"26",X"00",X"FD",X"6E",X"0E",X"06",X"00",X"DD",X"4E",
		X"0A",X"ED",X"42",X"3A",X"4E",X"87",X"47",X"CB",X"05",X"CB",X"14",X"10",X"FA",X"CD",X"24",X"21",
		X"ED",X"4B",X"3F",X"81",X"09",X"FD",X"E1",X"FD",X"72",X"04",X"FD",X"73",X"03",X"FD",X"74",X"0C",
		X"FD",X"75",X"0B",X"C9",X"CD",X"46",X"21",X"F6",X"10",X"4F",X"06",X"00",X"CB",X"21",X"CB",X"10",
		X"CB",X"7F",X"28",X"01",X"05",X"09",X"C9",X"3A",X"4D",X"87",X"47",X"4F",X"CB",X"39",X"CB",X"39",
		X"CD",X"46",X"21",X"A0",X"B1",X"C9",X"D9",X"2A",X"09",X"86",X"AF",X"57",X"5F",X"06",X"67",X"CB",
		X"40",X"28",X"03",X"EB",X"19",X"EB",X"29",X"CB",X"08",X"3C",X"FE",X"08",X"20",X"02",X"06",X"7A",
		X"FE",X"10",X"20",X"EB",X"21",X"2E",X"6A",X"19",X"22",X"09",X"86",X"7C",X"D9",X"C9",X"21",X"00",
		X"00",X"22",X"37",X"81",X"22",X"3F",X"81",X"21",X"CB",X"80",X"06",X"1F",X"AF",X"77",X"23",X"10",
		X"FC",X"21",X"00",X"00",X"22",X"C0",X"80",X"22",X"C7",X"80",X"C9",X"3A",X"B9",X"87",X"B7",X"C0",
		X"3E",X"FF",X"32",X"1A",X"86",X"1E",X"04",X"CD",X"E6",X"13",X"23",X"23",X"23",X"CB",X"38",X"08",
		X"04",X"2B",X"1D",X"10",X"FC",X"08",X"30",X"08",X"CB",X"21",X"CB",X"21",X"CB",X"21",X"CB",X"21",
		X"79",X"86",X"27",X"77",X"D0",X"2B",X"1D",X"C8",X"0E",X"01",X"18",X"F4",X"21",X"44",X"87",X"7E",
		X"C6",X"01",X"27",X"77",X"3E",X"03",X"CD",X"F4",X"2B",X"AF",X"C9",X"06",X"0A",X"C9",X"00",X"00",
		X"01",X"00",X"00",X"01",X"02",X"00",X"00",X"00",X"CD",X"FC",X"14",X"D2",X"9E",X"15",X"DD",X"E5",
		X"21",X"7E",X"87",X"34",X"CD",X"CB",X"14",X"D2",X"5C",X"22",X"FD",X"E1",X"CD",X"12",X"2C",X"CD",
		X"68",X"22",X"CD",X"04",X"23",X"DD",X"2A",X"BA",X"80",X"21",X"CE",X"21",X"DD",X"75",X"05",X"DD",
		X"74",X"06",X"DD",X"CB",X"0C",X"E6",X"3E",X"96",X"DD",X"77",X"03",X"DD",X"CB",X"00",X"EE",X"DD",
		X"CB",X"00",X"F6",X"DD",X"CB",X"00",X"D6",X"FD",X"E5",X"CD",X"7A",X"15",X"FD",X"E1",X"DD",X"CB",
		X"00",X"4E",X"CA",X"5C",X"22",X"DD",X"7E",X"0D",X"B7",X"20",X"31",X"FD",X"CB",X"00",X"76",X"C2",
		X"5C",X"22",X"DD",X"CB",X"00",X"6E",X"28",X"24",X"CD",X"1B",X"23",X"30",X"04",X"DD",X"36",X"03",
		X"0A",X"FD",X"7E",X"04",X"CD",X"FF",X"22",X"FE",X"08",X"30",X"11",X"FD",X"7E",X"0C",X"CD",X"FF",
		X"22",X"FE",X"08",X"30",X"07",X"FD",X"E5",X"CD",X"7A",X"15",X"18",X"C0",X"21",X"7E",X"87",X"35",
		X"CD",X"F4",X"15",X"CD",X"7A",X"15",X"18",X"FB",X"FD",X"21",X"34",X"81",X"DD",X"E5",X"DD",X"2A",
		X"88",X"87",X"26",X"00",X"FD",X"6E",X"06",X"16",X"00",X"DD",X"5E",X"08",X"B7",X"ED",X"52",X"3A",
		X"4E",X"87",X"47",X"3A",X"B7",X"87",X"B7",X"28",X"02",X"06",X"03",X"CB",X"05",X"CB",X"14",X"10",
		X"FA",X"CD",X"D4",X"22",X"ED",X"4B",X"37",X"81",X"09",X"EB",X"26",X"00",X"FD",X"6E",X"0E",X"06",
		X"00",X"DD",X"4E",X"0A",X"B7",X"ED",X"42",X"3A",X"4E",X"87",X"47",X"3A",X"B7",X"87",X"B7",X"28",
		X"02",X"06",X"03",X"CB",X"05",X"CB",X"14",X"10",X"FA",X"CD",X"D4",X"22",X"ED",X"4B",X"3F",X"81",
		X"09",X"FD",X"E1",X"FD",X"72",X"04",X"FD",X"73",X"03",X"FD",X"74",X"0C",X"FD",X"75",X"0B",X"AF",
		X"32",X"B7",X"87",X"C9",X"3A",X"B7",X"87",X"B7",X"C0",X"CD",X"46",X"21",X"4F",X"3A",X"4F",X"87",
		X"B7",X"28",X"05",X"47",X"CB",X"29",X"10",X"FC",X"06",X"00",X"CB",X"79",X"28",X"01",X"05",X"CB",
		X"21",X"CB",X"10",X"09",X"C9",X"F5",X"7A",X"2F",X"57",X"7B",X"2F",X"5F",X"13",X"F1",X"C9",X"B7",
		X"F0",X"ED",X"44",X"C9",X"DD",X"2A",X"88",X"87",X"2A",X"BA",X"80",X"11",X"08",X"00",X"19",X"DD",
		X"7E",X"08",X"77",X"23",X"23",X"DD",X"7E",X"0A",X"77",X"C9",X"9F",X"DD",X"6E",X"01",X"DD",X"66",
		X"02",X"E5",X"FD",X"E1",X"DD",X"E5",X"DD",X"21",X"15",X"82",X"DD",X"7E",X"08",X"FD",X"96",X"06",
		X"D2",X"35",X"23",X"ED",X"44",X"47",X"DD",X"7E",X"0A",X"FD",X"96",X"0E",X"D2",X"41",X"23",X"ED",
		X"44",X"4F",X"16",X"00",X"3E",X"0F",X"B9",X"38",X"03",X"B8",X"30",X"07",X"CB",X"38",X"CB",X"39",
		X"14",X"18",X"F3",X"79",X"07",X"07",X"07",X"07",X"B0",X"CB",X"22",X"D5",X"5F",X"16",X"00",X"21",
		X"E8",X"23",X"19",X"19",X"7E",X"23",X"66",X"6F",X"E5",X"7B",X"0F",X"0F",X"0F",X"0F",X"5F",X"D5",
		X"D1",X"21",X"E8",X"23",X"19",X"19",X"5E",X"23",X"56",X"E1",X"06",X"02",X"CB",X"25",X"CB",X"14",
		X"CB",X"23",X"CB",X"12",X"10",X"F6",X"F1",X"F5",X"B7",X"28",X"0B",X"47",X"CB",X"2A",X"CB",X"1B",
		X"CB",X"2C",X"CB",X"1D",X"10",X"F6",X"DD",X"7E",X"08",X"FD",X"BE",X"06",X"DC",X"DE",X"23",X"DD",
		X"7E",X"0A",X"FD",X"BE",X"0E",X"EB",X"DC",X"DE",X"23",X"EB",X"F1",X"B7",X"20",X"1B",X"3A",X"8E",
		X"87",X"B7",X"28",X"15",X"3A",X"5A",X"87",X"FE",X"01",X"28",X"0E",X"CD",X"6E",X"27",X"CD",X"DE",
		X"23",X"EB",X"CD",X"DE",X"23",X"EB",X"37",X"18",X"06",X"21",X"00",X"00",X"11",X"00",X"00",X"FD",
		X"74",X"02",X"FD",X"75",X"01",X"FD",X"72",X"0A",X"FD",X"73",X"09",X"DD",X"E1",X"C9",X"F5",X"7C",
		X"2F",X"67",X"7D",X"2F",X"6F",X"23",X"F1",X"C9",X"00",X"00",X"FF",X"3F",X"00",X"10",X"1C",X"07",
		X"00",X"04",X"8F",X"02",X"C7",X"01",X"4E",X"01",X"00",X"01",X"CA",X"00",X"A4",X"00",X"87",X"00",
		X"72",X"00",X"61",X"00",X"54",X"00",X"49",X"00",X"00",X"00",X"A1",X"16",X"73",X"0B",X"12",X"06",
		X"A7",X"03",X"6A",X"02",X"B5",X"01",X"44",X"01",X"FA",X"00",X"C7",X"00",X"A1",X"00",X"86",X"00",
		X"71",X"00",X"60",X"00",X"53",X"00",X"48",X"00",X"00",X"00",X"B9",X"05",X"A8",X"05",X"19",X"04",
		X"DD",X"02",X"0D",X"02",X"85",X"01",X"29",X"01",X"EA",X"00",X"BC",X"00",X"9A",X"00",X"81",X"00",
		X"6D",X"00",X"5E",X"00",X"51",X"00",X"47",X"00",X"00",X"00",X"06",X"02",X"BB",X"02",X"84",X"02",
		X"0C",X"02",X"9D",X"01",X"46",X"01",X"04",X"01",X"D2",X"00",X"AD",X"00",X"90",X"00",X"7A",X"00",
		X"68",X"00",X"5A",X"00",X"4E",X"00",X"45",X"00",X"00",X"00",X"EA",X"00",X"6E",X"01",X"89",X"01",
		X"6A",X"01",X"D5",X"00",X"06",X"01",X"DB",X"00",X"B7",X"00",X"9A",X"00",X"83",X"00",X"70",X"00",
		X"61",X"00",X"55",X"00",X"4A",X"00",X"42",X"00",X"00",X"00",X"7C",X"00",X"D2",X"00",X"F8",X"00",
		X"FA",X"00",X"E8",X"00",X"CE",X"00",X"B4",X"00",X"9C",X"00",X"87",X"00",X"75",X"00",X"66",X"00",
		X"59",X"00",X"4F",X"00",X"46",X"00",X"3E",X"00",X"00",X"00",X"49",X"00",X"82",X"00",X"A3",X"00",
		X"AF",X"00",X"AC",X"00",X"A1",X"00",X"92",X"00",X"83",X"00",X"75",X"00",X"67",X"00",X"5C",X"00",
		X"51",X"00",X"49",X"00",X"41",X"00",X"3A",X"00",X"00",X"00",X"2E",X"00",X"55",X"00",X"6F",X"00",
		X"7D",X"00",X"81",X"00",X"7D",X"00",X"76",X"00",X"6D",X"00",X"63",X"00",X"5A",X"00",X"51",X"00",
		X"49",X"00",X"42",X"00",X"3C",X"00",X"36",X"00",X"00",X"00",X"1F",X"00",X"3A",X"00",X"4F",X"00",
		X"5C",X"00",X"62",X"00",X"62",X"00",X"5F",X"00",X"5B",X"00",X"54",X"00",X"4E",X"00",X"48",X"00",
		X"42",X"00",X"3C",X"00",X"37",X"00",X"32",X"00",X"00",X"00",X"16",X"00",X"2A",X"00",X"3A",X"00",
		X"45",X"00",X"4B",X"00",X"4E",X"00",X"4D",X"00",X"4B",X"00",X"48",X"00",X"43",X"00",X"3F",X"00",
		X"3A",X"00",X"36",X"00",X"32",X"00",X"2E",X"00",X"00",X"00",X"10",X"00",X"1F",X"00",X"2B",X"00",
		X"34",X"00",X"3B",X"00",X"3E",X"00",X"3F",X"00",X"3E",X"00",X"3D",X"00",X"3A",X"00",X"37",X"00",
		X"34",X"00",X"30",X"00",X"2D",X"00",X"2A",X"00",X"00",X"00",X"0C",X"00",X"17",X"00",X"17",X"00",
		X"29",X"00",X"2E",X"00",X"32",X"00",X"34",X"00",X"34",X"00",X"33",X"00",X"32",X"00",X"30",X"00",
		X"2E",X"00",X"2B",X"00",X"29",X"00",X"26",X"00",X"00",X"00",X"09",X"00",X"12",X"00",X"1A",X"00",
		X"20",X"00",X"25",X"00",X"29",X"00",X"2B",X"00",X"2C",X"00",X"2C",X"00",X"2B",X"00",X"2A",X"00",
		X"28",X"00",X"26",X"00",X"25",X"00",X"23",X"00",X"00",X"00",X"07",X"00",X"0E",X"00",X"15",X"00",
		X"1A",X"00",X"1E",X"00",X"21",X"00",X"24",X"00",X"25",X"00",X"25",X"00",X"25",X"00",X"24",X"00",
		X"24",X"00",X"22",X"00",X"21",X"00",X"1F",X"00",X"00",X"00",X"06",X"00",X"0C",X"00",X"11",X"00",
		X"15",X"00",X"19",X"00",X"1C",X"00",X"1E",X"00",X"1F",X"00",X"20",X"00",X"20",X"00",X"20",X"00",
		X"1F",X"00",X"1F",X"00",X"1E",X"00",X"1C",X"00",X"00",X"00",X"05",X"00",X"09",X"00",X"0E",X"00",
		X"12",X"00",X"15",X"00",X"17",X"00",X"19",X"00",X"1B",X"00",X"1C",X"00",X"1C",X"00",X"1C",X"00",
		X"1C",X"00",X"1B",X"00",X"1B",X"00",X"1A",X"00",X"E7",X"1D",X"04",X"00",X"AF",X"32",X"2A",X"86",
		X"11",X"1F",X"8C",X"06",X"20",X"21",X"6E",X"26",X"22",X"28",X"86",X"C5",X"21",X"C4",X"FF",X"19",
		X"EB",X"21",X"28",X"86",X"7E",X"23",X"66",X"6F",X"23",X"7E",X"47",X"FE",X"01",X"28",X"1E",X"CD",
		X"46",X"21",X"0F",X"0F",X"E6",X"1F",X"FE",X"1B",X"30",X"F5",X"3C",X"32",X"2A",X"86",X"CD",X"46",
		X"21",X"0F",X"0F",X"0F",X"E6",X"0F",X"90",X"F2",X"26",X"26",X"80",X"3C",X"47",X"23",X"10",X"FD",
		X"4E",X"21",X"60",X"26",X"09",X"09",X"7E",X"23",X"66",X"6F",X"E5",X"3A",X"2A",X"86",X"06",X"00",
		X"4F",X"09",X"06",X"1D",X"7E",X"B7",X"20",X"07",X"22",X"28",X"86",X"E1",X"10",X"01",X"04",X"7E",
		X"12",X"13",X"23",X"10",X"EF",X"C1",X"10",X"A3",X"AF",X"32",X"27",X"86",X"32",X"C5",X"80",X"C9",
		X"71",X"26",X"92",X"26",X"B1",X"26",X"D2",X"26",X"F1",X"26",X"12",X"27",X"31",X"27",X"00",X"01",
		X"00",X"89",X"9F",X"91",X"93",X"9F",X"98",X"99",X"9F",X"8F",X"9B",X"8B",X"8C",X"9F",X"9F",X"8E",
		X"9A",X"8A",X"8D",X"9F",X"9F",X"90",X"93",X"88",X"89",X"9F",X"9B",X"99",X"9F",X"00",X"03",X"01",
		X"03",X"05",X"82",X"83",X"9F",X"92",X"93",X"91",X"9F",X"9F",X"9E",X"8D",X"99",X"91",X"9F",X"8C",
		X"9B",X"96",X"8E",X"9F",X"91",X"9F",X"9B",X"9F",X"9A",X"89",X"9F",X"99",X"8B",X"8E",X"00",X"01",
		X"02",X"80",X"81",X"9B",X"9A",X"9F",X"8C",X"8E",X"9F",X"9D",X"8C",X"9F",X"9A",X"93",X"98",X"9F",
		X"94",X"9F",X"88",X"89",X"9F",X"9F",X"90",X"91",X"8D",X"9F",X"8C",X"9F",X"9A",X"00",X"03",X"00",
		X"03",X"05",X"86",X"87",X"99",X"9F",X"9F",X"91",X"8D",X"8A",X"9F",X"9F",X"9E",X"8C",X"9F",X"98",
		X"96",X"8E",X"99",X"9F",X"9A",X"9F",X"96",X"8E",X"9F",X"9F",X"9F",X"8B",X"9F",X"8E",X"00",X"01",
		X"04",X"84",X"85",X"8C",X"8F",X"90",X"93",X"9A",X"9F",X"8E",X"9B",X"9C",X"9F",X"8F",X"8D",X"95",
		X"9B",X"9F",X"89",X"9F",X"98",X"94",X"99",X"9B",X"91",X"93",X"98",X"8C",X"9F",X"00",X"03",X"00",
		X"01",X"05",X"9E",X"8B",X"9A",X"98",X"8D",X"88",X"89",X"9F",X"8C",X"9A",X"96",X"8D",X"8E",X"9E",
		X"9F",X"91",X"9B",X"8B",X"89",X"8C",X"98",X"97",X"9F",X"9B",X"99",X"9A",X"9F",X"9F",X"00",X"01",
		X"06",X"9C",X"9F",X"8E",X"8C",X"90",X"9B",X"8C",X"9A",X"93",X"9F",X"95",X"9F",X"9F",X"9D",X"9F",
		X"91",X"93",X"9F",X"9A",X"93",X"8F",X"95",X"8C",X"9F",X"9F",X"8A",X"98",X"91",X"00",X"03",X"00",
		X"01",X"03",X"DF",X"16",X"CF",X"10",X"10",X"53",X"48",X"49",X"45",X"4C",X"44",X"53",X"20",X"5B",
		X"20",X"00",X"21",X"10",X"60",X"11",X"5A",X"87",X"06",X"02",X"CD",X"06",X"07",X"C9",X"08",X"D9",
		X"3A",X"8E",X"87",X"B7",X"28",X"18",X"3A",X"5A",X"87",X"B7",X"28",X"12",X"3A",X"5B",X"87",X"D6",
		X"0C",X"27",X"32",X"5B",X"87",X"3A",X"5A",X"87",X"DE",X"00",X"27",X"32",X"5A",X"87",X"D9",X"08",
		X"C9",X"08",X"D9",X"3A",X"B9",X"87",X"B7",X"20",X"1A",X"3A",X"8E",X"87",X"B7",X"20",X"14",X"21",
		X"20",X"82",X"CB",X"46",X"20",X"0D",X"3A",X"5A",X"87",X"FE",X"99",X"28",X"06",X"C6",X"01",X"27",
		X"32",X"5A",X"87",X"D9",X"08",X"C9",X"DF",X"16",X"CF",X"A0",X"10",X"46",X"55",X"45",X"4C",X"20",
		X"5B",X"20",X"00",X"21",X"10",X"D8",X"11",X"58",X"87",X"06",X"02",X"CD",X"06",X"07",X"C9",X"08",
		X"D9",X"2A",X"37",X"81",X"7C",X"B5",X"20",X"07",X"2A",X"3F",X"81",X"7C",X"B5",X"28",X"21",X"3A",
		X"58",X"87",X"B7",X"28",X"1B",X"3A",X"59",X"87",X"D6",X"06",X"27",X"32",X"59",X"87",X"3A",X"58",
		X"87",X"DE",X"00",X"27",X"32",X"58",X"87",X"FE",X"10",X"20",X"05",X"3E",X"15",X"CD",X"F4",X"2B",
		X"D9",X"08",X"C9",X"08",X"D9",X"3A",X"58",X"87",X"FE",X"99",X"28",X"0A",X"C6",X"01",X"27",X"32",
		X"58",X"87",X"21",X"1A",X"86",X"35",X"D9",X"08",X"C9",X"21",X"C7",X"80",X"ED",X"5B",X"37",X"81",
		X"7A",X"B7",X"F8",X"7B",X"86",X"77",X"2B",X"7A",X"8E",X"27",X"77",X"2B",X"7E",X"CE",X"00",X"27",
		X"77",X"C9",X"00",X"00",X"01",X"00",X"00",X"0C",X"0C",X"82",X"36",X"04",X"0C",X"0C",X"82",X"35",
		X"04",X"0C",X"0C",X"82",X"B4",X"04",X"0C",X"0C",X"82",X"34",X"04",X"0C",X"0C",X"82",X"B5",X"04",
		X"00",X"01",X"37",X"28",X"00",X"00",X"01",X"00",X"00",X"0C",X"0C",X"02",X"36",X"06",X"0C",X"0C",
		X"03",X"36",X"07",X"00",X"01",X"59",X"28",X"CD",X"04",X"15",X"30",X"FB",X"CD",X"44",X"2C",X"CD",
		X"03",X"2B",X"AF",X"32",X"9F",X"87",X"32",X"A0",X"87",X"3E",X"99",X"32",X"90",X"87",X"CD",X"48",
		X"1E",X"CD",X"15",X"04",X"CD",X"7A",X"15",X"CD",X"CB",X"2A",X"38",X"1C",X"DD",X"CB",X"00",X"6E",
		X"20",X"0F",X"CD",X"A8",X"04",X"CD",X"1A",X"2C",X"3A",X"90",X"87",X"B7",X"20",X"03",X"C3",X"6F",
		X"2A",X"3E",X"1E",X"CD",X"CE",X"15",X"18",X"DF",X"CD",X"BA",X"14",X"38",X"05",X"CD",X"7A",X"15",
		X"18",X"F6",X"DD",X"E5",X"FD",X"E1",X"FD",X"22",X"A1",X"87",X"DD",X"2A",X"BA",X"80",X"3E",X"EF",
		X"DD",X"77",X"08",X"CD",X"EB",X"2A",X"DD",X"77",X"0A",X"CD",X"B5",X"2A",X"DD",X"CB",X"00",X"D6",
		X"DD",X"CB",X"00",X"F6",X"DD",X"CB",X"0C",X"F6",X"CD",X"7A",X"15",X"FD",X"2A",X"A1",X"87",X"FD",
		X"CB",X"00",X"76",X"C2",X"79",X"2A",X"3A",X"90",X"87",X"B7",X"CA",X"44",X"2A",X"DD",X"7E",X"08",
		X"32",X"9F",X"87",X"DD",X"7E",X"0A",X"32",X"A0",X"87",X"DD",X"7E",X"0D",X"CB",X"4F",X"C2",X"09",
		X"29",X"CD",X"EE",X"2A",X"CD",X"7A",X"15",X"18",X"D2",X"DD",X"CB",X"00",X"A6",X"21",X"54",X"28",
		X"DD",X"75",X"05",X"DD",X"74",X"06",X"DD",X"36",X"04",X"01",X"DD",X"CB",X"00",X"E6",X"FD",X"21",
		X"15",X"82",X"DD",X"7E",X"08",X"FD",X"77",X"08",X"DD",X"7E",X"0A",X"FD",X"77",X"0A",X"FD",X"21",
		X"34",X"81",X"AF",X"FD",X"77",X"03",X"FD",X"77",X"04",X"FD",X"77",X"0B",X"FD",X"77",X"0C",X"FD",
		X"77",X"01",X"FD",X"77",X"02",X"FD",X"77",X"09",X"FD",X"77",X"0A",X"3E",X"2D",X"32",X"8F",X"87",
		X"FD",X"2A",X"A1",X"87",X"DD",X"CB",X"0D",X"4E",X"20",X"12",X"DD",X"7E",X"08",X"32",X"9F",X"87",
		X"DD",X"7E",X"0A",X"32",X"A0",X"87",X"CD",X"B5",X"2A",X"C3",X"04",X"29",X"CD",X"EE",X"2A",X"DD",
		X"CB",X"00",X"4E",X"CA",X"79",X"2A",X"3A",X"90",X"87",X"B7",X"CA",X"44",X"2A",X"3E",X"01",X"CD",
		X"CE",X"15",X"21",X"8F",X"87",X"35",X"20",X"C8",X"3E",X"14",X"32",X"D4",X"87",X"FD",X"2A",X"A1",
		X"87",X"DD",X"CB",X"0D",X"4E",X"20",X"05",X"CD",X"B5",X"2A",X"18",X"78",X"DD",X"7E",X"08",X"32",
		X"9F",X"87",X"DD",X"7E",X"0A",X"32",X"A0",X"87",X"CD",X"EE",X"2A",X"CD",X"C3",X"27",X"3E",X"0A",
		X"CD",X"F4",X"2B",X"DD",X"CB",X"00",X"4E",X"CA",X"79",X"2A",X"3A",X"90",X"87",X"B7",X"CA",X"44",
		X"2A",X"3A",X"D4",X"87",X"FE",X"01",X"28",X"04",X"3D",X"32",X"D4",X"87",X"CD",X"CE",X"15",X"CD",
		X"03",X"28",X"CD",X"03",X"28",X"CD",X"03",X"28",X"3A",X"58",X"87",X"FE",X"99",X"C2",X"8D",X"29",
		X"3E",X"00",X"CD",X"F4",X"2B",X"CD",X"B5",X"2A",X"CD",X"74",X"3C",X"06",X"16",X"FD",X"2A",X"A1",
		X"87",X"FD",X"CB",X"00",X"76",X"C2",X"79",X"2A",X"DD",X"CB",X"00",X"4E",X"CA",X"79",X"2A",X"3E",
		X"82",X"32",X"C1",X"87",X"3A",X"90",X"87",X"B7",X"CA",X"44",X"2A",X"C5",X"3E",X"01",X"CD",X"CE",
		X"15",X"C1",X"10",X"D9",X"FD",X"2A",X"A1",X"87",X"DD",X"CB",X"00",X"D6",X"FD",X"36",X"04",X"FF",
		X"FD",X"CB",X"00",X"76",X"C2",X"79",X"2A",X"DD",X"CB",X"00",X"4E",X"CA",X"79",X"2A",X"DD",X"7E",
		X"08",X"32",X"9F",X"87",X"DD",X"7E",X"0A",X"32",X"A0",X"87",X"3E",X"82",X"32",X"C1",X"87",X"CD",
		X"7A",X"15",X"18",X"D0",X"3E",X"07",X"CD",X"F4",X"2B",X"DD",X"CB",X"00",X"A6",X"21",X"83",X"0E",
		X"DD",X"75",X"05",X"DD",X"74",X"06",X"DD",X"36",X"04",X"01",X"DD",X"CB",X"00",X"E6",X"DD",X"CB",
		X"00",X"66",X"28",X"1E",X"DD",X"CB",X"00",X"4E",X"28",X"18",X"CD",X"7A",X"15",X"18",X"EF",X"CD",
		X"01",X"2D",X"3E",X"3C",X"CD",X"CE",X"15",X"18",X"09",X"3A",X"5C",X"87",X"C6",X"01",X"27",X"32",
		X"5C",X"87",X"CD",X"04",X"16",X"DD",X"CB",X"00",X"A6",X"DD",X"CB",X"00",X"96",X"DD",X"CB",X"00",
		X"BE",X"DD",X"CB",X"00",X"B6",X"DD",X"CB",X"0C",X"B6",X"DD",X"CB",X"00",X"CE",X"DD",X"36",X"0D",
		X"00",X"DD",X"36",X"08",X"00",X"DD",X"36",X"0A",X"00",X"3A",X"46",X"87",X"C6",X"01",X"27",X"32",
		X"46",X"87",X"C3",X"6F",X"28",X"DD",X"CB",X"00",X"A6",X"21",X"32",X"28",X"DD",X"75",X"05",X"DD",
		X"74",X"06",X"DD",X"36",X"04",X"01",X"DD",X"CB",X"00",X"E6",X"C9",X"2A",X"5D",X"87",X"ED",X"5B",
		X"8C",X"87",X"3A",X"1D",X"82",X"2F",X"4F",X"06",X"00",X"09",X"EB",X"B7",X"ED",X"52",X"C9",X"CD",
		X"46",X"21",X"FE",X"20",X"38",X"F9",X"FE",X"E8",X"30",X"F5",X"C9",X"3E",X"80",X"C9",X"C5",X"DD",
		X"CB",X"0D",X"66",X"28",X"08",X"3E",X"03",X"CD",X"28",X"2C",X"CD",X"1A",X"2C",X"DD",X"36",X"0D",
		X"00",X"C1",X"C9",X"3A",X"46",X"87",X"FE",X"07",X"30",X"0F",X"21",X"25",X"2B",X"5F",X"16",X"00",
		X"19",X"19",X"5E",X"23",X"56",X"ED",X"53",X"BD",X"87",X"2A",X"5D",X"87",X"ED",X"5B",X"BD",X"87",
		X"19",X"22",X"8C",X"87",X"C9",X"30",X"02",X"80",X"03",X"30",X"05",X"80",X"07",X"00",X"09",X"30",
		X"0A",X"40",X"0B",X"00",X"00",X"01",X"00",X"00",X"01",X"00",X"05",X"3A",X"04",X"01",X"00",X"05",
		X"3A",X"03",X"01",X"00",X"05",X"3A",X"02",X"00",X"01",X"38",X"2B",X"CD",X"DC",X"14",X"D2",X"9E",
		X"15",X"CD",X"BA",X"14",X"D2",X"DB",X"2B",X"DD",X"E5",X"FD",X"E1",X"DD",X"2A",X"BA",X"80",X"CD",
		X"B1",X"2B",X"21",X"33",X"2B",X"DD",X"75",X"05",X"DD",X"74",X"06",X"DD",X"36",X"04",X"01",X"DD",
		X"CB",X"00",X"E6",X"DD",X"CB",X"00",X"D6",X"FD",X"E5",X"CD",X"7A",X"15",X"FD",X"E1",X"DD",X"CB",
		X"00",X"4E",X"CA",X"DB",X"2B",X"FD",X"CB",X"00",X"76",X"C2",X"DB",X"2B",X"3A",X"8E",X"87",X"B7",
		X"28",X"49",X"3A",X"5A",X"87",X"B7",X"28",X"43",X"DD",X"CB",X"0B",X"C6",X"3E",X"0C",X"CD",X"F4",
		X"2B",X"CD",X"B1",X"2B",X"CD",X"C6",X"2B",X"CD",X"6E",X"27",X"FD",X"E5",X"CD",X"7A",X"15",X"18",
		X"CB",X"FD",X"E5",X"FD",X"21",X"15",X"82",X"FD",X"7E",X"08",X"DD",X"77",X"08",X"FD",X"7E",X"0A",
		X"DD",X"77",X"0A",X"FD",X"E1",X"C9",X"DD",X"E5",X"DD",X"21",X"34",X"81",X"DD",X"7E",X"04",X"FD",
		X"77",X"04",X"DD",X"7E",X"0C",X"FD",X"77",X"0C",X"DD",X"E1",X"C9",X"DD",X"CB",X"0B",X"46",X"CA",
		X"E7",X"2B",X"3E",X"17",X"CD",X"F4",X"2B",X"3E",X"00",X"32",X"8E",X"87",X"CD",X"F4",X"15",X"CD",
		X"7A",X"15",X"18",X"FB",X"F3",X"32",X"00",X"A0",X"3A",X"B9",X"87",X"B7",X"C0",X"AF",X"32",X"01",
		X"A0",X"E3",X"E3",X"3E",X"08",X"32",X"01",X"A0",X"FB",X"C9",X"3E",X"08",X"18",X"E6",X"3E",X"06",
		X"18",X"E2",X"3E",X"12",X"18",X"DE",X"3E",X"14",X"18",X"DA",X"3A",X"90",X"87",X"FE",X"99",X"C8",
		X"FE",X"90",X"D2",X"72",X"2C",X"C3",X"A8",X"2C",X"D9",X"47",X"3A",X"90",X"87",X"B8",X"30",X"03",
		X"AF",X"18",X"02",X"90",X"27",X"32",X"90",X"87",X"D9",X"C9",X"21",X"18",X"00",X"01",X"01",X"20",
		X"CD",X"93",X"07",X"C9",X"CD",X"B1",X"07",X"48",X"A0",X"20",X"46",X"55",X"45",X"4C",X"20",X"42",
		X"41",X"53",X"45",X"20",X"3F",X"20",X"00",X"C9",X"21",X"18",X"00",X"01",X"01",X"20",X"CD",X"93",
		X"07",X"DF",X"19",X"CF",X"58",X"18",X"42",X"4F",X"4E",X"55",X"53",X"20",X"53",X"48",X"49",X"50",
		X"00",X"C9",X"DF",X"1C",X"21",X"18",X"00",X"01",X"01",X"20",X"CD",X"93",X"07",X"CF",X"20",X"18",
		X"46",X"55",X"45",X"4C",X"20",X"42",X"41",X"53",X"45",X"20",X"00",X"21",X"18",X"70",X"11",X"46",
		X"87",X"06",X"02",X"CD",X"06",X"07",X"CF",X"80",X"18",X"20",X"55",X"4E",X"44",X"45",X"52",X"20",
		X"41",X"54",X"54",X"41",X"43",X"4B",X"00",X"C9",X"3A",X"90",X"87",X"FE",X"20",X"30",X"04",X"DF",
		X"1C",X"18",X"42",X"FE",X"50",X"30",X"04",X"DF",X"1B",X"18",X"3A",X"FE",X"80",X"30",X"04",X"DF",
		X"1A",X"18",X"32",X"DF",X"1D",X"21",X"18",X"00",X"01",X"01",X"20",X"CD",X"93",X"07",X"CF",X"20",
		X"18",X"46",X"55",X"45",X"4C",X"20",X"42",X"41",X"53",X"45",X"20",X"20",X"20",X"20",X"53",X"48",
		X"49",X"45",X"4C",X"44",X"53",X"20",X"20",X"20",X"3E",X"00",X"21",X"18",X"70",X"11",X"46",X"87",
		X"06",X"02",X"CD",X"06",X"07",X"21",X"18",X"C8",X"11",X"90",X"87",X"06",X"02",X"CD",X"06",X"07",
		X"C9",X"DF",X"19",X"21",X"18",X"00",X"01",X"01",X"20",X"CD",X"93",X"07",X"CF",X"30",X"18",X"46",
		X"55",X"45",X"4C",X"20",X"42",X"41",X"53",X"45",X"20",X"44",X"45",X"53",X"54",X"52",X"4F",X"59",
		X"45",X"44",X"00",X"3E",X"07",X"CD",X"F4",X"2B",X"3A",X"9F",X"87",X"B7",X"C0",X"3A",X"7D",X"87",
		X"D6",X"05",X"D0",X"FD",X"21",X"10",X"38",X"CD",X"62",X"15",X"C9",X"CD",X"DC",X"14",X"D2",X"9E",
		X"15",X"21",X"7D",X"87",X"34",X"CD",X"BA",X"14",X"D2",X"A9",X"2E",X"DD",X"E5",X"FD",X"E1",X"DD",
		X"2A",X"BA",X"80",X"CD",X"D9",X"2E",X"C3",X"74",X"2D",X"CD",X"DC",X"14",X"D2",X"9E",X"15",X"21",
		X"7D",X"87",X"34",X"CD",X"BA",X"14",X"D2",X"A9",X"2E",X"DD",X"E5",X"FD",X"E1",X"DD",X"2A",X"BA",
		X"80",X"CD",X"B5",X"2E",X"CD",X"0D",X"2F",X"E5",X"DD",X"36",X"03",X"14",X"DD",X"CB",X"00",X"EE",
		X"DD",X"CB",X"00",X"F6",X"DD",X"CB",X"0C",X"EE",X"DD",X"36",X"0B",X"02",X"DD",X"CB",X"00",X"D6",
		X"3E",X"04",X"CD",X"3A",X"3E",X"CD",X"7A",X"15",X"DD",X"6E",X"01",X"DD",X"66",X"02",X"E5",X"FD",
		X"E1",X"DD",X"CB",X"00",X"4E",X"CA",X"A9",X"2E",X"DD",X"7E",X"0D",X"B7",X"C2",X"4F",X"2E",X"CD",
		X"1B",X"23",X"30",X"09",X"3E",X"05",X"DD",X"77",X"03",X"DD",X"CB",X"00",X"EE",X"FD",X"CB",X"00",
		X"76",X"C2",X"A9",X"2E",X"DD",X"CB",X"00",X"6E",X"20",X"16",X"CD",X"46",X"21",X"07",X"07",X"07",
		X"E6",X"07",X"C6",X"01",X"DD",X"77",X"03",X"DD",X"CB",X"00",X"EE",X"E1",X"CD",X"E5",X"2D",X"E5",
		X"CD",X"7A",X"15",X"18",X"B3",X"1E",X"00",X"3A",X"1D",X"82",X"DD",X"BE",X"08",X"30",X"01",X"1C",
		X"3A",X"1F",X"82",X"DD",X"BE",X"0A",X"30",X"02",X"1C",X"1C",X"7B",X"BE",X"20",X"38",X"DD",X"7E",
		X"0B",X"E6",X"38",X"0F",X"0F",X"0F",X"3C",X"FE",X"07",X"28",X"15",X"CB",X"27",X"CB",X"27",X"CB",
		X"27",X"5F",X"DD",X"7E",X"0B",X"E6",X"C7",X"B3",X"DD",X"77",X"0B",X"2B",X"2B",X"C3",X"23",X"2F",
		X"CD",X"3A",X"1F",X"30",X"11",X"FD",X"E5",X"E5",X"DD",X"22",X"88",X"87",X"FD",X"21",X"D8",X"21",
		X"CD",X"62",X"15",X"E1",X"FD",X"E1",X"DD",X"7E",X"0B",X"E6",X"C7",X"DD",X"77",X"0B",X"23",X"7E",
		X"B7",X"20",X"09",X"23",X"7E",X"2B",X"B7",X"20",X"03",X"21",X"6D",X"2F",X"C3",X"0D",X"2F",X"CD",
		X"16",X"2C",X"FD",X"E5",X"E1",X"E5",X"11",X"01",X"00",X"19",X"AF",X"06",X"04",X"77",X"23",X"10",
		X"FC",X"E1",X"11",X"09",X"00",X"19",X"06",X"05",X"77",X"23",X"10",X"FC",X"DD",X"CB",X"0C",X"AE",
		X"DD",X"CB",X"00",X"A6",X"21",X"83",X"0E",X"DD",X"75",X"05",X"DD",X"74",X"06",X"DD",X"36",X"04",
		X"01",X"DD",X"CB",X"00",X"E6",X"06",X"02",X"0E",X"01",X"CD",X"8B",X"21",X"06",X"01",X"0E",X"05",
		X"CD",X"8B",X"21",X"3E",X"04",X"CD",X"31",X"3E",X"DD",X"CB",X"00",X"66",X"28",X"0B",X"DD",X"CB",
		X"00",X"4E",X"28",X"05",X"CD",X"7A",X"15",X"18",X"EF",X"21",X"7D",X"87",X"35",X"CD",X"F4",X"15",
		X"CD",X"7A",X"15",X"18",X"FB",X"FD",X"E5",X"FD",X"2A",X"9D",X"87",X"FD",X"7E",X"08",X"DD",X"77",
		X"08",X"FD",X"7E",X"0A",X"DD",X"77",X"0A",X"CD",X"46",X"21",X"07",X"07",X"E6",X"01",X"21",X"6D",
		X"2F",X"28",X"03",X"21",X"BD",X"2F",X"FD",X"E1",X"C9",X"CD",X"46",X"21",X"07",X"07",X"E6",X"01",
		X"28",X"13",X"CD",X"46",X"21",X"FE",X"20",X"38",X"F9",X"FE",X"E8",X"30",X"F5",X"47",X"3E",X"0B",
		X"21",X"6D",X"2F",X"18",X"11",X"CD",X"46",X"21",X"FE",X"20",X"38",X"F9",X"FE",X"E8",X"30",X"F5",
		X"47",X"3E",X"EF",X"21",X"95",X"2F",X"DD",X"77",X"08",X"DD",X"70",X"0A",X"C9",X"DD",X"CB",X"00",
		X"A6",X"7E",X"DD",X"77",X"05",X"23",X"7E",X"DD",X"77",X"06",X"DD",X"36",X"04",X"01",X"DD",X"CB",
		X"00",X"E6",X"23",X"7E",X"E5",X"ED",X"5B",X"48",X"87",X"B7",X"47",X"F2",X"34",X"2F",X"ED",X"44",
		X"47",X"CD",X"F5",X"22",X"04",X"21",X"00",X"00",X"19",X"10",X"FD",X"ED",X"52",X"ED",X"4B",X"37",
		X"81",X"09",X"FD",X"74",X"04",X"FD",X"75",X"03",X"E1",X"23",X"7E",X"E5",X"ED",X"5B",X"48",X"87",
		X"B7",X"47",X"F2",X"5B",X"2F",X"ED",X"44",X"47",X"CD",X"F5",X"22",X"04",X"21",X"00",X"00",X"19",
		X"10",X"FD",X"ED",X"52",X"FD",X"74",X"0C",X"FD",X"75",X"0B",X"E1",X"23",X"C9",X"0F",X"30",X"04",
		X"00",X"02",X"22",X"30",X"03",X"FF",X"02",X"35",X"30",X"02",X"FE",X"02",X"48",X"30",X"01",X"FD",
		X"02",X"5B",X"30",X"00",X"FC",X"03",X"6E",X"30",X"FF",X"FD",X"03",X"81",X"30",X"FE",X"FE",X"03",
		X"94",X"30",X"FD",X"FF",X"03",X"A7",X"30",X"FC",X"00",X"01",X"94",X"30",X"FD",X"FF",X"03",X"81",
		X"30",X"FE",X"FE",X"03",X"6E",X"30",X"FF",X"FD",X"03",X"5B",X"30",X"00",X"FC",X"03",X"48",X"30",
		X"01",X"FD",X"02",X"35",X"30",X"02",X"FE",X"02",X"22",X"30",X"03",X"FF",X"02",X"0F",X"30",X"04",
		X"00",X"02",X"2C",X"31",X"03",X"01",X"00",X"19",X"31",X"02",X"02",X"00",X"06",X"31",X"01",X"03",
		X"00",X"F3",X"30",X"00",X"04",X"00",X"E0",X"30",X"FF",X"03",X"01",X"CD",X"30",X"FE",X"02",X"01",
		X"BA",X"30",X"FD",X"01",X"01",X"A7",X"30",X"FC",X"00",X"01",X"BA",X"30",X"FD",X"01",X"01",X"CD",
		X"30",X"FE",X"02",X"01",X"E0",X"30",X"FF",X"03",X"01",X"F3",X"30",X"00",X"04",X"00",X"06",X"31",
		X"01",X"03",X"00",X"19",X"31",X"02",X"02",X"00",X"2C",X"31",X"03",X"01",X"00",X"00",X"00",X"00",
		X"00",X"01",X"00",X"00",X"09",X"09",X"04",X"28",X"06",X"09",X"09",X"04",X"28",X"05",X"00",X"01",
		X"14",X"30",X"00",X"00",X"01",X"00",X"00",X"09",X"09",X"04",X"29",X"06",X"09",X"09",X"04",X"29",
		X"05",X"00",X"01",X"27",X"30",X"00",X"00",X"01",X"00",X"00",X"09",X"09",X"04",X"2A",X"06",X"09",
		X"09",X"04",X"2A",X"05",X"00",X"01",X"3A",X"30",X"00",X"00",X"01",X"00",X"00",X"09",X"09",X"04",
		X"2B",X"06",X"09",X"09",X"04",X"2B",X"05",X"00",X"01",X"4D",X"30",X"00",X"00",X"01",X"00",X"00",
		X"09",X"09",X"04",X"2C",X"06",X"09",X"09",X"04",X"2C",X"05",X"00",X"01",X"60",X"30",X"00",X"00",
		X"01",X"00",X"00",X"09",X"09",X"04",X"AB",X"06",X"09",X"09",X"04",X"AB",X"05",X"00",X"01",X"73",
		X"30",X"00",X"00",X"01",X"00",X"00",X"09",X"09",X"04",X"AA",X"06",X"09",X"09",X"04",X"AA",X"05",
		X"00",X"01",X"86",X"30",X"00",X"00",X"01",X"00",X"00",X"09",X"09",X"04",X"A9",X"06",X"09",X"09",
		X"04",X"A9",X"05",X"00",X"01",X"99",X"30",X"00",X"00",X"01",X"00",X"00",X"09",X"09",X"04",X"A8",
		X"06",X"09",X"09",X"04",X"A8",X"05",X"00",X"01",X"AC",X"30",X"00",X"00",X"01",X"00",X"00",X"09",
		X"09",X"04",X"E9",X"06",X"09",X"09",X"04",X"E9",X"05",X"00",X"01",X"BF",X"30",X"00",X"00",X"01",
		X"00",X"00",X"09",X"09",X"04",X"EA",X"06",X"09",X"09",X"04",X"EA",X"05",X"00",X"01",X"D2",X"30",
		X"00",X"00",X"01",X"00",X"00",X"09",X"09",X"04",X"EB",X"06",X"09",X"09",X"04",X"EB",X"05",X"00",
		X"01",X"E5",X"30",X"00",X"00",X"01",X"00",X"00",X"09",X"09",X"04",X"6C",X"06",X"09",X"09",X"04",
		X"6C",X"05",X"00",X"01",X"F8",X"30",X"00",X"00",X"01",X"00",X"00",X"09",X"09",X"04",X"6B",X"06",
		X"09",X"09",X"04",X"6B",X"05",X"00",X"01",X"0B",X"31",X"00",X"00",X"01",X"00",X"00",X"09",X"09",
		X"04",X"6A",X"06",X"09",X"09",X"04",X"6A",X"05",X"00",X"01",X"1E",X"31",X"00",X"00",X"01",X"00",
		X"00",X"09",X"09",X"04",X"69",X"06",X"09",X"09",X"04",X"69",X"05",X"00",X"01",X"31",X"31",X"00",
		X"00",X"01",X"00",X"00",X"0F",X"0A",X"09",X"2E",X"01",X"0F",X"0A",X"09",X"2E",X"04",X"00",X"01",
		X"44",X"31",X"00",X"00",X"01",X"00",X"00",X"0E",X"08",X"03",X"32",X"01",X"0E",X"08",X"03",X"32",
		X"04",X"00",X"01",X"57",X"31",X"00",X"00",X"01",X"00",X"00",X"0E",X"08",X"01",X"33",X"01",X"0E",
		X"08",X"01",X"33",X"04",X"00",X"01",X"6A",X"31",X"CD",X"DC",X"14",X"D2",X"9E",X"15",X"21",X"7D",
		X"87",X"34",X"CD",X"BA",X"14",X"D2",X"CA",X"32",X"DD",X"E5",X"FD",X"E1",X"DD",X"2A",X"BA",X"80",
		X"CD",X"D9",X"32",X"CD",X"32",X"33",X"CD",X"EF",X"32",X"CD",X"37",X"21",X"DD",X"77",X"03",X"DD",
		X"CB",X"00",X"EE",X"DD",X"CB",X"00",X"F6",X"DD",X"CB",X"0C",X"FE",X"DD",X"36",X"0B",X"01",X"DD",
		X"CB",X"00",X"D6",X"3E",X"11",X"CD",X"F4",X"2B",X"AF",X"CD",X"3A",X"3E",X"FD",X"E5",X"CD",X"7A",
		X"15",X"FD",X"E1",X"FD",X"CB",X"00",X"76",X"C2",X"CA",X"32",X"CD",X"1B",X"23",X"DD",X"7E",X"0D",
		X"B7",X"C4",X"5C",X"32",X"3A",X"9F",X"87",X"B7",X"28",X"2A",X"DD",X"96",X"08",X"DA",X"E9",X"31",
		X"FE",X"3C",X"38",X"16",X"CD",X"47",X"33",X"18",X"1B",X"ED",X"44",X"FE",X"3C",X"38",X"0B",X"21",
		X"BC",X"FE",X"FD",X"75",X"03",X"FD",X"74",X"04",X"18",X"0A",X"FD",X"36",X"04",X"00",X"FD",X"36",
		X"03",X"00",X"18",X"00",X"FD",X"E5",X"DD",X"CB",X"00",X"6E",X"20",X"4A",X"3A",X"9F",X"87",X"B7",
		X"28",X"26",X"CD",X"3A",X"1F",X"30",X"21",X"CD",X"37",X"21",X"DD",X"77",X"03",X"DD",X"CB",X"00",
		X"EE",X"3E",X"13",X"CD",X"F4",X"2B",X"DD",X"22",X"88",X"87",X"FD",X"21",X"56",X"33",X"CD",X"62",
		X"15",X"3A",X"7D",X"87",X"FE",X"02",X"38",X"1E",X"3A",X"7D",X"87",X"21",X"4A",X"87",X"BE",X"30",
		X"15",X"CD",X"37",X"21",X"DD",X"77",X"03",X"DD",X"CB",X"00",X"EE",X"DD",X"22",X"9D",X"87",X"FD",
		X"21",X"59",X"2D",X"CD",X"62",X"15",X"CD",X"7A",X"15",X"C3",X"C1",X"31",X"DD",X"CB",X"0D",X"56",
		X"20",X"00",X"3E",X"14",X"CD",X"F4",X"2B",X"CD",X"05",X"33",X"DD",X"7E",X"0B",X"C6",X"10",X"DD",
		X"77",X"0B",X"E6",X"F0",X"FE",X"30",X"DD",X"36",X"0D",X"00",X"C0",X"FD",X"E5",X"E1",X"E5",X"11",
		X"01",X"00",X"19",X"AF",X"06",X"04",X"77",X"23",X"10",X"FC",X"E1",X"11",X"09",X"00",X"19",X"06",
		X"05",X"77",X"23",X"10",X"FC",X"DD",X"CB",X"0C",X"BE",X"DD",X"CB",X"00",X"A6",X"21",X"83",X"0E",
		X"DD",X"75",X"05",X"DD",X"74",X"06",X"DD",X"36",X"04",X"01",X"DD",X"CB",X"00",X"E6",X"01",X"05",
		X"01",X"CD",X"8B",X"21",X"3E",X"00",X"CD",X"31",X"3E",X"DD",X"CB",X"00",X"66",X"28",X"0E",X"DD",
		X"CB",X"00",X"4E",X"28",X"08",X"CD",X"7A",X"15",X"18",X"EF",X"CD",X"A6",X"02",X"21",X"7D",X"87",
		X"35",X"CD",X"F4",X"15",X"CD",X"7A",X"15",X"18",X"FB",X"06",X"0B",X"21",X"96",X"87",X"CB",X"7E",
		X"28",X"02",X"06",X"EF",X"21",X"9C",X"87",X"7E",X"DD",X"70",X"08",X"DD",X"77",X"0A",X"C9",X"21",
		X"3F",X"31",X"DD",X"CB",X"00",X"A6",X"DD",X"75",X"05",X"DD",X"74",X"06",X"DD",X"36",X"04",X"01",
		X"DD",X"CB",X"00",X"E6",X"C9",X"01",X"05",X"01",X"CD",X"8B",X"21",X"DD",X"7E",X"0B",X"E6",X"F0",
		X"FE",X"00",X"20",X"05",X"21",X"52",X"31",X"18",X"06",X"FE",X"10",X"C0",X"21",X"65",X"31",X"DD",
		X"CB",X"00",X"A6",X"DD",X"75",X"05",X"DD",X"74",X"06",X"DD",X"36",X"04",X"01",X"DD",X"CB",X"00",
		X"E6",X"C9",X"21",X"96",X"87",X"01",X"00",X"00",X"CB",X"7E",X"28",X"0B",X"23",X"7E",X"23",X"B6",
		X"28",X"08",X"01",X"BC",X"FE",X"18",X"03",X"01",X"44",X"01",X"2A",X"37",X"81",X"09",X"FD",X"74",
		X"04",X"FD",X"75",X"03",X"C9",X"CC",X"CD",X"FC",X"14",X"D2",X"9E",X"15",X"21",X"7E",X"87",X"34",
		X"CD",X"CB",X"14",X"D2",X"D4",X"33",X"DD",X"E5",X"FD",X"E1",X"DD",X"2A",X"BA",X"80",X"CD",X"12",
		X"2C",X"CD",X"E0",X"33",X"CD",X"26",X"34",X"21",X"CE",X"21",X"DD",X"75",X"05",X"DD",X"74",X"06",
		X"DD",X"CB",X"0C",X"E6",X"3E",X"96",X"DD",X"77",X"03",X"DD",X"CB",X"00",X"EE",X"DD",X"CB",X"00",
		X"F6",X"DD",X"CB",X"00",X"D6",X"FD",X"E5",X"CD",X"7A",X"15",X"FD",X"E1",X"DD",X"CB",X"00",X"4E",
		X"CA",X"D4",X"33",X"DD",X"7E",X"0D",X"B7",X"20",X"2B",X"FD",X"CB",X"00",X"76",X"C2",X"D4",X"33",
		X"DD",X"CB",X"00",X"6E",X"28",X"1E",X"CD",X"1B",X"23",X"FD",X"7E",X"04",X"CD",X"FF",X"22",X"FE",
		X"08",X"30",X"11",X"FD",X"7E",X"0C",X"CD",X"FF",X"22",X"FE",X"08",X"30",X"07",X"FD",X"E5",X"CD",
		X"7A",X"15",X"18",X"C6",X"21",X"7E",X"87",X"35",X"CD",X"F4",X"15",X"CD",X"7A",X"15",X"18",X"FB",
		X"FD",X"E5",X"DD",X"2A",X"88",X"87",X"26",X"00",X"3A",X"9F",X"87",X"6F",X"16",X"00",X"DD",X"5E",
		X"08",X"B7",X"ED",X"52",X"06",X"03",X"CB",X"05",X"CB",X"14",X"10",X"FA",X"EB",X"26",X"00",X"3A",
		X"A0",X"87",X"6F",X"06",X"00",X"DD",X"4E",X"0A",X"B7",X"ED",X"42",X"06",X"03",X"CB",X"05",X"CB",
		X"14",X"10",X"FA",X"FD",X"E1",X"FD",X"72",X"04",X"FD",X"73",X"03",X"FD",X"74",X"0C",X"FD",X"75",
		X"0B",X"DD",X"2A",X"BA",X"80",X"C9",X"DD",X"2A",X"88",X"87",X"2A",X"BA",X"80",X"11",X"08",X"00",
		X"19",X"DD",X"7E",X"08",X"77",X"23",X"23",X"DD",X"7E",X"0A",X"77",X"DD",X"2A",X"BA",X"80",X"C9",
		X"CD",X"DC",X"14",X"D2",X"9E",X"15",X"21",X"7D",X"87",X"34",X"CD",X"BA",X"14",X"D2",X"61",X"35",
		X"DD",X"E5",X"FD",X"E1",X"DD",X"2A",X"BA",X"80",X"CD",X"6D",X"35",X"CD",X"85",X"35",X"E5",X"DD",
		X"36",X"03",X"05",X"DD",X"CB",X"00",X"EE",X"DD",X"CB",X"00",X"F6",X"DD",X"CB",X"0C",X"EE",X"DD",
		X"36",X"0B",X"04",X"DD",X"CB",X"00",X"D6",X"3E",X"03",X"CD",X"3A",X"3E",X"CD",X"7A",X"15",X"DD",
		X"6E",X"01",X"DD",X"66",X"02",X"E5",X"FD",X"E1",X"DD",X"CB",X"00",X"4E",X"CA",X"61",X"35",X"DD",
		X"7E",X"0D",X"B7",X"C2",X"0E",X"35",X"CD",X"1B",X"23",X"30",X"09",X"3E",X"05",X"DD",X"77",X"03",
		X"DD",X"CB",X"00",X"EE",X"FD",X"CB",X"00",X"76",X"C2",X"61",X"35",X"DD",X"CB",X"00",X"6E",X"20",
		X"0E",X"E1",X"CD",X"C4",X"34",X"E5",X"3E",X"05",X"DD",X"77",X"03",X"DD",X"CB",X"00",X"EE",X"CD",
		X"7A",X"15",X"18",X"BB",X"7E",X"B7",X"28",X"1D",X"3A",X"7E",X"87",X"FE",X"04",X"30",X"2E",X"FD",
		X"E5",X"E5",X"DD",X"22",X"88",X"87",X"FD",X"21",X"D8",X"21",X"CD",X"62",X"15",X"E1",X"FD",X"E1",
		X"2B",X"2B",X"C3",X"9B",X"35",X"CD",X"46",X"21",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"47",X"3A",
		X"1D",X"82",X"90",X"DD",X"BE",X"08",X"38",X"05",X"2B",X"2B",X"C3",X"9B",X"35",X"23",X"7E",X"B7",
		X"20",X"09",X"23",X"7E",X"2B",X"B7",X"20",X"03",X"21",X"EF",X"35",X"C3",X"85",X"35",X"CD",X"16",
		X"2C",X"FD",X"E5",X"E1",X"E5",X"11",X"01",X"00",X"19",X"AF",X"06",X"04",X"77",X"23",X"10",X"FC",
		X"E1",X"11",X"09",X"00",X"19",X"06",X"05",X"77",X"23",X"10",X"FC",X"DD",X"CB",X"0C",X"AE",X"DD",
		X"CB",X"00",X"A6",X"21",X"83",X"0E",X"DD",X"75",X"05",X"DD",X"74",X"06",X"DD",X"36",X"04",X"01",
		X"DD",X"CB",X"00",X"E6",X"06",X"02",X"0E",X"03",X"CD",X"8B",X"21",X"3E",X"03",X"CD",X"31",X"3E",
		X"DD",X"CB",X"00",X"66",X"28",X"0B",X"DD",X"CB",X"00",X"4E",X"28",X"05",X"CD",X"7A",X"15",X"18",
		X"EF",X"21",X"7D",X"87",X"35",X"CD",X"F4",X"15",X"CD",X"7A",X"15",X"18",X"FB",X"CD",X"46",X"21",
		X"FE",X"20",X"38",X"F9",X"FE",X"E8",X"30",X"F5",X"47",X"3E",X"0B",X"DD",X"77",X"08",X"DD",X"70",
		X"0A",X"21",X"E5",X"35",X"C9",X"DD",X"CB",X"00",X"A6",X"7E",X"DD",X"77",X"05",X"23",X"7E",X"DD",
		X"77",X"06",X"DD",X"36",X"04",X"01",X"DD",X"CB",X"00",X"E6",X"23",X"7E",X"E5",X"ED",X"5B",X"48",
		X"87",X"B7",X"47",X"F2",X"AC",X"35",X"ED",X"44",X"47",X"CD",X"F5",X"22",X"04",X"21",X"00",X"00",
		X"19",X"10",X"FD",X"ED",X"52",X"ED",X"4B",X"37",X"81",X"09",X"FD",X"74",X"04",X"FD",X"75",X"03",
		X"E1",X"23",X"7E",X"E5",X"ED",X"5B",X"48",X"87",X"B7",X"47",X"F2",X"D3",X"35",X"ED",X"44",X"47",
		X"CD",X"F5",X"22",X"04",X"21",X"00",X"00",X"19",X"10",X"FD",X"ED",X"52",X"FD",X"74",X"0C",X"FD",
		X"75",X"0B",X"E1",X"23",X"C9",X"04",X"36",X"03",X"03",X"00",X"F6",X"35",X"00",X"00",X"01",X"12",
		X"36",X"03",X"FD",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"09",X"09",X"04",X"2F",X"02",
		X"00",X"01",X"FB",X"35",X"00",X"00",X"01",X"00",X"00",X"09",X"09",X"04",X"30",X"02",X"00",X"01",
		X"09",X"36",X"00",X"00",X"01",X"00",X"00",X"09",X"09",X"04",X"70",X"02",X"00",X"01",X"17",X"36",
		X"CD",X"DC",X"14",X"D2",X"9E",X"15",X"21",X"7D",X"87",X"34",X"CD",X"BA",X"14",X"D2",X"42",X"37",
		X"DD",X"E5",X"FD",X"E1",X"DD",X"2A",X"BA",X"80",X"CD",X"51",X"37",X"CD",X"66",X"37",X"DD",X"CB",
		X"00",X"A6",X"21",X"95",X"37",X"DD",X"75",X"05",X"DD",X"74",X"06",X"DD",X"36",X"04",X"01",X"DD",
		X"CB",X"00",X"E6",X"DD",X"36",X"03",X"0A",X"DD",X"CB",X"00",X"EE",X"DD",X"CB",X"00",X"F6",X"DD",
		X"CB",X"0C",X"EE",X"DD",X"36",X"0B",X"04",X"DD",X"CB",X"00",X"D6",X"3E",X"01",X"CD",X"3A",X"3E",
		X"CD",X"7A",X"15",X"DD",X"6E",X"01",X"DD",X"66",X"02",X"E5",X"FD",X"E1",X"DD",X"CB",X"00",X"4E",
		X"CA",X"42",X"37",X"DD",X"7E",X"0D",X"B7",X"C2",X"EF",X"36",X"CD",X"1B",X"23",X"30",X"09",X"3E",
		X"05",X"DD",X"77",X"03",X"DD",X"CB",X"00",X"EE",X"FD",X"CB",X"00",X"76",X"C2",X"42",X"37",X"DD",
		X"CB",X"00",X"6E",X"20",X"0B",X"CD",X"85",X"37",X"DD",X"CB",X"0B",X"AE",X"DD",X"CB",X"00",X"EE",
		X"DD",X"CB",X"0B",X"6E",X"20",X"34",X"3A",X"1F",X"82",X"DD",X"96",X"0A",X"F2",X"C1",X"36",X"ED",
		X"44",X"FE",X"05",X"30",X"25",X"3A",X"7E",X"87",X"FE",X"04",X"30",X"0F",X"DD",X"22",X"88",X"87",
		X"FD",X"21",X"D8",X"21",X"CD",X"62",X"15",X"DD",X"CB",X"0B",X"EE",X"3A",X"1D",X"82",X"DD",X"96",
		X"08",X"CB",X"3F",X"DD",X"77",X"03",X"DD",X"CB",X"00",X"EE",X"CD",X"7A",X"15",X"18",X"84",X"CD",
		X"16",X"2C",X"FD",X"E5",X"E1",X"E5",X"11",X"01",X"00",X"19",X"AF",X"06",X"04",X"77",X"23",X"10",
		X"FC",X"E1",X"11",X"09",X"00",X"19",X"06",X"05",X"77",X"23",X"10",X"FC",X"DD",X"CB",X"0C",X"AE",
		X"DD",X"CB",X"00",X"A6",X"21",X"83",X"0E",X"DD",X"75",X"05",X"DD",X"74",X"06",X"DD",X"36",X"04",
		X"01",X"DD",X"CB",X"00",X"E6",X"06",X"02",X"0E",X"04",X"CD",X"8B",X"21",X"3E",X"01",X"CD",X"31",
		X"3E",X"DD",X"CB",X"00",X"66",X"28",X"0E",X"DD",X"CB",X"00",X"4E",X"28",X"08",X"CD",X"7A",X"15",
		X"18",X"EF",X"CD",X"A6",X"02",X"21",X"7D",X"87",X"35",X"CD",X"F4",X"15",X"CD",X"7A",X"15",X"18",
		X"FB",X"CD",X"46",X"21",X"FE",X"20",X"38",X"F9",X"FE",X"E8",X"30",X"F5",X"47",X"3E",X"0B",X"DD",
		X"77",X"08",X"DD",X"70",X"0A",X"C9",X"21",X"60",X"00",X"ED",X"4B",X"37",X"81",X"09",X"FD",X"74",
		X"04",X"FD",X"75",X"03",X"ED",X"5B",X"48",X"87",X"2A",X"48",X"87",X"19",X"29",X"19",X"FD",X"74",
		X"0C",X"FD",X"75",X"0B",X"C9",X"FD",X"56",X"0C",X"FD",X"5E",X"0B",X"CD",X"F5",X"22",X"FD",X"72",
		X"0C",X"FD",X"73",X"0B",X"C9",X"00",X"00",X"01",X"00",X"00",X"09",X"09",X"10",X"1F",X"02",X"09",
		X"09",X"10",X"0C",X"02",X"09",X"09",X"10",X"11",X"02",X"09",X"09",X"10",X"12",X"02",X"09",X"09",
		X"10",X"1F",X"03",X"09",X"09",X"10",X"0C",X"03",X"09",X"09",X"10",X"11",X"03",X"09",X"09",X"10",
		X"12",X"03",X"09",X"09",X"10",X"1F",X"04",X"09",X"09",X"10",X"0C",X"04",X"09",X"09",X"10",X"11",
		X"04",X"09",X"09",X"10",X"12",X"04",X"09",X"09",X"10",X"1F",X"01",X"09",X"09",X"10",X"0C",X"01",
		X"09",X"09",X"10",X"11",X"01",X"09",X"09",X"10",X"12",X"01",X"00",X"01",X"9A",X"37",X"CD",X"DC",
		X"14",X"D2",X"9E",X"15",X"21",X"7D",X"87",X"34",X"CD",X"BA",X"14",X"D2",X"93",X"39",X"DD",X"E5",
		X"FD",X"E1",X"DD",X"2A",X"BA",X"80",X"DD",X"36",X"0B",X"02",X"DD",X"CB",X"0B",X"FE",X"18",X"1C",
		X"CD",X"DC",X"14",X"D2",X"9E",X"15",X"21",X"7D",X"87",X"34",X"CD",X"BA",X"14",X"D2",X"93",X"39",
		X"DD",X"E5",X"FD",X"E1",X"DD",X"2A",X"BA",X"80",X"DD",X"36",X"0B",X"02",X"DD",X"6E",X"01",X"DD",
		X"66",X"02",X"E5",X"FD",X"E1",X"DD",X"CB",X"00",X"CE",X"FD",X"CB",X"00",X"B6",X"DD",X"CB",X"00",
		X"A6",X"21",X"47",X"3A",X"DD",X"75",X"05",X"DD",X"74",X"06",X"DD",X"36",X"04",X"01",X"DD",X"CB",
		X"00",X"E6",X"CD",X"B1",X"39",X"21",X"15",X"3A",X"CD",X"C6",X"39",X"E5",X"DD",X"36",X"03",X"10",
		X"DD",X"CB",X"00",X"EE",X"DD",X"CB",X"00",X"F6",X"DD",X"CB",X"0C",X"EE",X"DD",X"CB",X"00",X"D6",
		X"CD",X"7A",X"15",X"DD",X"6E",X"01",X"DD",X"66",X"02",X"E5",X"FD",X"E1",X"DD",X"CB",X"00",X"4E",
		X"CA",X"93",X"39",X"DD",X"7E",X"0D",X"B7",X"C2",X"42",X"39",X"3A",X"9F",X"87",X"B7",X"28",X"13",
		X"DD",X"CB",X"0B",X"F6",X"DD",X"CB",X"0B",X"7E",X"20",X"09",X"3E",X"0A",X"DD",X"77",X"03",X"DD",
		X"CB",X"00",X"EE",X"CD",X"1B",X"23",X"30",X"09",X"3E",X"05",X"DD",X"77",X"03",X"DD",X"CB",X"00",
		X"EE",X"FD",X"CB",X"00",X"76",X"C2",X"93",X"39",X"DD",X"CB",X"00",X"6E",X"20",X"0D",X"E1",X"CD",
		X"D0",X"38",X"E5",X"DD",X"36",X"03",X"05",X"DD",X"CB",X"00",X"EE",X"CD",X"7A",X"15",X"18",X"A3",
		X"DD",X"CB",X"0B",X"6E",X"20",X"0B",X"3A",X"38",X"81",X"FE",X"02",X"30",X"50",X"DD",X"CB",X"0B",
		X"EE",X"1E",X"00",X"3A",X"1D",X"82",X"DD",X"BE",X"08",X"30",X"01",X"1C",X"3A",X"1F",X"82",X"DD",
		X"BE",X"0A",X"30",X"02",X"1C",X"1C",X"7B",X"BE",X"20",X"05",X"2B",X"2B",X"C3",X"C6",X"39",X"3A",
		X"7E",X"87",X"FE",X"03",X"30",X"16",X"FD",X"E5",X"E5",X"3E",X"FF",X"32",X"B7",X"87",X"DD",X"22",
		X"88",X"87",X"FD",X"21",X"D8",X"21",X"CD",X"62",X"15",X"E1",X"FD",X"E1",X"23",X"7E",X"B7",X"20",
		X"09",X"23",X"7E",X"2B",X"B7",X"20",X"03",X"21",X"15",X"3A",X"C3",X"C6",X"39",X"ED",X"5B",X"37",
		X"81",X"FD",X"72",X"04",X"FD",X"73",X"03",X"ED",X"5B",X"3F",X"81",X"FD",X"72",X"0C",X"FD",X"73",
		X"0B",X"C9",X"CD",X"16",X"2C",X"FD",X"E5",X"E1",X"E5",X"11",X"01",X"00",X"19",X"AF",X"06",X"04",
		X"77",X"23",X"10",X"FC",X"E1",X"11",X"09",X"00",X"19",X"06",X"05",X"77",X"23",X"10",X"FC",X"DD",
		X"CB",X"0C",X"AE",X"DD",X"CB",X"00",X"A6",X"21",X"83",X"0E",X"DD",X"75",X"05",X"DD",X"74",X"06",
		X"DD",X"36",X"04",X"01",X"DD",X"CB",X"00",X"E6",X"06",X"02",X"0E",X"01",X"CD",X"8B",X"21",X"CD",
		X"31",X"3E",X"DD",X"CB",X"00",X"66",X"28",X"0B",X"DD",X"CB",X"00",X"4E",X"28",X"05",X"CD",X"7A",
		X"15",X"18",X"EF",X"DD",X"36",X"0D",X"00",X"E1",X"DD",X"CB",X"0B",X"7E",X"20",X"07",X"DD",X"CB",
		X"0B",X"76",X"CA",X"2C",X"38",X"21",X"7D",X"87",X"35",X"CD",X"F4",X"15",X"CD",X"7A",X"15",X"18",
		X"FB",X"CD",X"46",X"21",X"FE",X"20",X"38",X"F9",X"FE",X"E8",X"30",X"F5",X"47",X"3E",X"0B",X"DD",
		X"77",X"08",X"DD",X"70",X"0A",X"C9",X"7E",X"E5",X"11",X"B0",X"00",X"B7",X"47",X"F2",X"D6",X"39",
		X"ED",X"44",X"47",X"CD",X"F5",X"22",X"04",X"21",X"00",X"00",X"19",X"10",X"FD",X"ED",X"52",X"29",
		X"ED",X"4B",X"37",X"81",X"09",X"FD",X"74",X"04",X"FD",X"75",X"03",X"E1",X"23",X"7E",X"E5",X"11",
		X"B0",X"00",X"B7",X"47",X"F2",X"FD",X"39",X"ED",X"44",X"47",X"CD",X"F5",X"22",X"04",X"21",X"00",
		X"00",X"19",X"10",X"FD",X"ED",X"52",X"29",X"ED",X"4B",X"3F",X"81",X"09",X"FD",X"74",X"0C",X"FD",
		X"75",X"0B",X"E1",X"23",X"C9",X"04",X"00",X"02",X"03",X"FF",X"02",X"02",X"FE",X"02",X"01",X"FD",
		X"02",X"00",X"FC",X"03",X"FF",X"FD",X"03",X"FE",X"FE",X"03",X"FD",X"FF",X"03",X"FC",X"00",X"01",
		X"FD",X"01",X"01",X"FE",X"02",X"01",X"FF",X"03",X"01",X"00",X"04",X"00",X"01",X"03",X"00",X"02",
		X"02",X"00",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"06",X"06",X"04",X"31",
		X"07",X"00",X"01",X"4C",X"3A",X"CD",X"DC",X"14",X"D2",X"9E",X"15",X"3A",X"7D",X"87",X"FE",X"05",
		X"30",X"06",X"CD",X"BA",X"14",X"DA",X"6D",X"3A",X"CD",X"7A",X"15",X"18",X"EE",X"21",X"7D",X"87",
		X"34",X"DD",X"E5",X"FD",X"E1",X"DD",X"2A",X"BA",X"80",X"DD",X"CB",X"00",X"CE",X"DD",X"CB",X"00",
		X"A6",X"21",X"8D",X"3B",X"DD",X"75",X"05",X"DD",X"74",X"06",X"DD",X"36",X"04",X"01",X"DD",X"CB",
		X"00",X"E6",X"CD",X"4B",X"3B",X"CD",X"7E",X"3B",X"DD",X"CB",X"00",X"F6",X"DD",X"CB",X"0C",X"EE",
		X"DD",X"36",X"0B",X"02",X"DD",X"CB",X"00",X"D6",X"3E",X"0D",X"CD",X"F4",X"2B",X"CD",X"7A",X"15",
		X"DD",X"6E",X"01",X"DD",X"66",X"02",X"E5",X"FD",X"E1",X"DD",X"CB",X"00",X"4E",X"CA",X"3F",X"3B",
		X"DD",X"7E",X"0D",X"B7",X"C2",X"F2",X"3A",X"CD",X"1B",X"23",X"30",X"09",X"3E",X"05",X"DD",X"77",
		X"03",X"DD",X"CB",X"00",X"EE",X"FD",X"CB",X"00",X"76",X"C2",X"3F",X"3B",X"DD",X"CB",X"00",X"6E",
		X"20",X"0B",X"CD",X"60",X"3B",X"DD",X"36",X"03",X"05",X"DD",X"CB",X"00",X"EE",X"CD",X"7A",X"15",
		X"18",X"BE",X"CD",X"16",X"2C",X"CD",X"BC",X"21",X"FD",X"E5",X"E1",X"E5",X"11",X"01",X"00",X"19",
		X"AF",X"06",X"04",X"77",X"23",X"10",X"FC",X"E1",X"11",X"09",X"00",X"19",X"06",X"05",X"77",X"23",
		X"10",X"FC",X"DD",X"CB",X"0C",X"AE",X"DD",X"CB",X"00",X"A6",X"21",X"83",X"0E",X"DD",X"75",X"05",
		X"DD",X"74",X"06",X"DD",X"36",X"04",X"01",X"DD",X"CB",X"00",X"E6",X"CD",X"58",X"2C",X"DD",X"CB",
		X"00",X"66",X"28",X"0B",X"DD",X"CB",X"00",X"4E",X"28",X"05",X"CD",X"7A",X"15",X"18",X"EF",X"21",
		X"7D",X"87",X"35",X"CD",X"F4",X"15",X"CD",X"7A",X"15",X"18",X"FB",X"CD",X"46",X"21",X"FE",X"20",
		X"38",X"F9",X"FE",X"E8",X"30",X"F5",X"47",X"3E",X"0B",X"DD",X"77",X"08",X"DD",X"70",X"0A",X"C9",
		X"CD",X"46",X"21",X"1F",X"1F",X"1F",X"1F",X"E6",X"07",X"67",X"CD",X"46",X"21",X"CB",X"77",X"20",
		X"04",X"7C",X"ED",X"44",X"67",X"CD",X"46",X"21",X"FD",X"74",X"0C",X"FD",X"77",X"0B",X"2A",X"48",
		X"87",X"ED",X"4B",X"37",X"81",X"09",X"FD",X"74",X"04",X"FD",X"75",X"03",X"C9",X"00",X"00",X"01",
		X"00",X"00",X"0E",X"0A",X"10",X"1D",X"02",X"00",X"01",X"92",X"3B",X"31",X"80",X"80",X"F5",X"3A",
		X"00",X"B0",X"F1",X"CD",X"61",X"07",X"F5",X"3A",X"00",X"B0",X"F1",X"D7",X"00",X"E7",X"04",X"04",
		X"01",X"E7",X"04",X"08",X"02",X"E7",X"04",X"0C",X"03",X"E7",X"04",X"10",X"04",X"3E",X"93",X"32",
		X"03",X"98",X"3E",X"88",X"32",X"03",X"A0",X"F5",X"3A",X"00",X"B0",X"F1",X"3E",X"10",X"32",X"02",
		X"98",X"CF",X"60",X"20",X"50",X"4F",X"52",X"54",X"20",X"41",X"20",X"31",X"00",X"21",X"30",X"40",
		X"CD",X"B8",X"06",X"3A",X"00",X"98",X"CD",X"5C",X"3C",X"3E",X"00",X"32",X"02",X"98",X"CF",X"60",
		X"40",X"50",X"4F",X"52",X"54",X"20",X"41",X"20",X"32",X"00",X"21",X"50",X"40",X"CD",X"B8",X"06",
		X"3A",X"00",X"98",X"CD",X"5C",X"3C",X"CF",X"68",X"60",X"50",X"4F",X"52",X"54",X"20",X"42",X"00",
		X"21",X"70",X"40",X"CD",X"B8",X"06",X"3A",X"01",X"98",X"CD",X"5C",X"3C",X"CF",X"68",X"80",X"50",
		X"4F",X"52",X"54",X"20",X"43",X"00",X"21",X"90",X"40",X"CD",X"B8",X"06",X"3A",X"02",X"98",X"CD",
		X"5C",X"3C",X"CF",X"40",X"A8",X"37",X"20",X"36",X"20",X"35",X"20",X"34",X"20",X"33",X"20",X"32",
		X"20",X"31",X"20",X"30",X"00",X"CF",X"50",X"B0",X"42",X"49",X"54",X"20",X"4E",X"55",X"4D",X"42",
		X"45",X"52",X"53",X"00",X"2E",X"00",X"2D",X"20",X"FD",X"C3",X"C7",X"3B",X"06",X"08",X"07",X"F5",
		X"E6",X"01",X"F6",X"30",X"CD",X"49",X"07",X"AF",X"CD",X"49",X"07",X"F5",X"3A",X"00",X"B0",X"F1",
		X"F1",X"10",X"EB",X"C9",X"AF",X"CD",X"F4",X"2B",X"21",X"C8",X"87",X"11",X"C2",X"87",X"06",X"06",
		X"1A",X"CD",X"5A",X"3E",X"12",X"F5",X"7E",X"CD",X"5A",X"3E",X"77",X"F1",X"BE",X"30",X"02",X"7E",
		X"12",X"23",X"13",X"10",X"EB",X"CD",X"43",X"3E",X"21",X"18",X"00",X"01",X"1D",X"20",X"CD",X"93",
		X"07",X"21",X"00",X"90",X"0E",X"01",X"CD",X"88",X"07",X"F5",X"3A",X"00",X"B0",X"F1",X"CF",X"68",
		X"20",X"42",X"4F",X"4E",X"55",X"53",X"00",X"CD",X"C3",X"27",X"CD",X"62",X"27",X"CD",X"9E",X"0B",
		X"E7",X"1C",X"04",X"02",X"21",X"00",X"00",X"22",X"CE",X"87",X"3A",X"CE",X"87",X"FE",X"05",X"38",
		X"09",X"C3",X"BE",X"3D",X"21",X"CE",X"87",X"34",X"18",X"F0",X"F5",X"3A",X"00",X"B0",X"F1",X"11",
		X"C2",X"87",X"2A",X"CE",X"87",X"19",X"7E",X"B7",X"CA",X"D4",X"3C",X"11",X"60",X"3E",X"2A",X"CE",
		X"87",X"29",X"19",X"5E",X"23",X"56",X"D5",X"11",X"C7",X"3E",X"2A",X"CE",X"87",X"19",X"5E",X"7B",
		X"32",X"D3",X"87",X"16",X"10",X"E1",X"CD",X"F4",X"3D",X"3E",X"18",X"32",X"D2",X"87",X"3A",X"D3",
		X"87",X"C6",X"08",X"32",X"D3",X"87",X"21",X"01",X"00",X"22",X"D0",X"87",X"2A",X"D0",X"87",X"E5",
		X"11",X"C2",X"87",X"2A",X"CE",X"87",X"19",X"7E",X"E1",X"BD",X"D2",X"36",X"3D",X"C3",X"69",X"3D",
		X"21",X"D0",X"87",X"34",X"18",X"E6",X"3A",X"D2",X"87",X"67",X"3A",X"D3",X"87",X"6F",X"CD",X"B8",
		X"06",X"E5",X"11",X"B8",X"3E",X"2A",X"CE",X"87",X"19",X"7E",X"87",X"87",X"E1",X"CD",X"51",X"1C",
		X"3A",X"D2",X"87",X"C6",X"10",X"FE",X"EF",X"38",X"0A",X"3A",X"D3",X"87",X"C6",X"10",X"32",X"D3",
		X"87",X"3E",X"18",X"32",X"D2",X"87",X"C3",X"30",X"3D",X"01",X"00",X"20",X"CD",X"E5",X"3D",X"11",
		X"C8",X"87",X"2A",X"CE",X"87",X"19",X"7E",X"B7",X"CA",X"D4",X"3C",X"35",X"11",X"FA",X"FF",X"19",
		X"35",X"3A",X"D2",X"87",X"D6",X"10",X"FE",X"18",X"30",X"0A",X"3A",X"D3",X"87",X"D6",X"10",X"32",
		X"D3",X"87",X"3E",X"E8",X"32",X"D2",X"87",X"3A",X"D2",X"87",X"67",X"3A",X"D3",X"87",X"6F",X"CD",
		X"B8",X"06",X"3E",X"DC",X"CD",X"51",X"1C",X"11",X"BD",X"3E",X"2A",X"CE",X"87",X"29",X"19",X"4E",
		X"23",X"46",X"CD",X"8B",X"21",X"CD",X"0E",X"3E",X"CD",X"16",X"2C",X"C3",X"69",X"3D",X"CD",X"4F",
		X"3E",X"01",X"00",X"40",X"CD",X"E5",X"3D",X"21",X"00",X"00",X"22",X"C7",X"80",X"AF",X"32",X"C4",
		X"80",X"CD",X"E8",X"25",X"CD",X"49",X"3E",X"3A",X"46",X"87",X"E6",X"0F",X"C0",X"FD",X"21",X"55",
		X"3A",X"CD",X"62",X"15",X"C9",X"DD",X"E5",X"DD",X"E1",X"F5",X"3A",X"00",X"B0",X"F1",X"0D",X"20",
		X"F4",X"10",X"F2",X"C9",X"EB",X"CD",X"B8",X"06",X"1A",X"13",X"B7",X"28",X"05",X"CD",X"49",X"07",
		X"18",X"F6",X"11",X"AB",X"3E",X"1A",X"13",X"B7",X"C8",X"CD",X"49",X"07",X"18",X"F7",X"AF",X"32",
		X"1A",X"86",X"3A",X"43",X"87",X"FE",X"02",X"28",X"0C",X"21",X"08",X"10",X"11",X"2E",X"81",X"06",
		X"06",X"CD",X"06",X"07",X"C9",X"21",X"08",X"C0",X"11",X"31",X"81",X"06",X"06",X"CD",X"06",X"07",
		X"C9",X"21",X"C8",X"87",X"5F",X"16",X"00",X"19",X"34",X"C9",X"21",X"C2",X"87",X"5F",X"16",X"00",
		X"19",X"34",X"C9",X"3E",X"FF",X"32",X"25",X"86",X"C9",X"3E",X"55",X"32",X"25",X"86",X"C9",X"21",
		X"C2",X"87",X"06",X"0C",X"36",X"00",X"23",X"10",X"FB",X"C9",X"FE",X"1D",X"D8",X"3E",X"1C",X"C9",
		X"6A",X"3E",X"76",X"3E",X"82",X"3E",X"91",X"3E",X"9E",X"3E",X"42",X"4F",X"4D",X"42",X"45",X"52",
		X"20",X"5B",X"20",X"32",X"30",X"00",X"54",X"52",X"41",X"43",X"45",X"52",X"20",X"5B",X"20",X"35",
		X"30",X"00",X"53",X"41",X"54",X"45",X"4C",X"4C",X"49",X"54",X"45",X"20",X"5B",X"20",X"31",X"30",
		X"00",X"53",X"54",X"52",X"41",X"46",X"45",X"52",X"20",X"5B",X"20",X"33",X"30",X"00",X"46",X"49",
		X"47",X"48",X"54",X"45",X"52",X"20",X"5B",X"20",X"31",X"30",X"00",X"20",X"50",X"4F",X"49",X"4E",
		X"54",X"53",X"20",X"45",X"41",X"43",X"48",X"00",X"2E",X"1F",X"0D",X"30",X"28",X"02",X"01",X"05",
		X"01",X"01",X"01",X"03",X"01",X"01",X"01",X"30",X"58",X"80",X"A8",X"D0",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
