library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_SND_0 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_SND_0 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"F3",X"31",X"00",X"81",X"C3",X"5B",X"0A",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C3",X"E9",X"0D",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"7C",X"00",X"3C",X"89",X"07",X"3C",X"B6",X"07",X"3C",X"E3",X"07",X"3B",X"10",X"08",X"3D",
		X"3D",X"08",X"78",X"98",X"08",X"7D",X"B9",X"08",X"64",X"EF",X"08",X"64",X"13",X"09",X"5F",X"31",
		X"09",X"73",X"58",X"09",X"74",X"8F",X"09",X"74",X"C9",X"09",X"79",X"03",X"0A",X"7E",X"24",X"0A",
		X"64",X"7D",X"00",X"00",X"7C",X"00",X"32",X"7B",X"01",X"7E",X"D4",X"06",X"21",X"18",X"01",X"01",
		X"01",X"01",X"01",X"01",X"19",X"57",X"03",X"55",X"03",X"59",X"03",X"1F",X"2C",X"01",X"0D",X"1D",
		X"10",X"10",X"10",X"07",X"BB",X"00",X"05",X"81",X"13",X"05",X"81",X"19",X"A7",X"02",X"A5",X"02",
		X"A9",X"02",X"1F",X"2C",X"01",X"0D",X"1D",X"10",X"10",X"10",X"07",X"BB",X"00",X"05",X"81",X"13",
		X"05",X"81",X"19",X"3B",X"02",X"39",X"02",X"3D",X"02",X"1F",X"2C",X"01",X"0D",X"1D",X"10",X"10",
		X"10",X"07",X"BB",X"00",X"05",X"81",X"13",X"05",X"81",X"19",X"FC",X"01",X"FA",X"01",X"FE",X"01",
		X"1F",X"2C",X"01",X"0D",X"1D",X"10",X"10",X"10",X"07",X"BB",X"00",X"05",X"81",X"13",X"05",X"81",
		X"19",X"A7",X"02",X"A5",X"02",X"A9",X"02",X"1F",X"2C",X"01",X"0D",X"1D",X"10",X"10",X"10",X"07",
		X"5D",X"00",X"05",X"81",X"13",X"05",X"81",X"11",X"FC",X"01",X"FA",X"01",X"FE",X"01",X"1F",X"2C",
		X"01",X"0D",X"1D",X"10",X"10",X"10",X"07",X"BB",X"00",X"05",X"81",X"13",X"05",X"81",X"1F",X"40",
		X"1F",X"00",X"1D",X"10",X"10",X"10",X"07",X"1F",X"00",X"05",X"81",X"13",X"05",X"81",X"19",X"AC",
		X"01",X"AA",X"01",X"AE",X"01",X"1F",X"2C",X"01",X"0D",X"1D",X"10",X"10",X"10",X"07",X"BB",X"00",
		X"05",X"81",X"13",X"05",X"81",X"19",X"7D",X"01",X"7B",X"01",X"7F",X"01",X"1F",X"2C",X"01",X"0D",
		X"1D",X"10",X"10",X"10",X"07",X"BB",X"00",X"05",X"81",X"13",X"05",X"81",X"19",X"3B",X"02",X"39",
		X"02",X"3D",X"02",X"1F",X"2C",X"01",X"0D",X"1D",X"10",X"10",X"10",X"07",X"BB",X"00",X"05",X"81",
		X"13",X"05",X"81",X"19",X"AC",X"01",X"AA",X"01",X"AE",X"01",X"1F",X"2C",X"01",X"0D",X"1D",X"10",
		X"10",X"10",X"07",X"FA",X"00",X"05",X"81",X"13",X"05",X"81",X"10",X"18",X"01",X"01",X"01",X"01",
		X"01",X"01",X"19",X"D6",X"00",X"D4",X"00",X"D8",X"00",X"1F",X"2C",X"01",X"0D",X"1D",X"10",X"10",
		X"10",X"07",X"1F",X"00",X"05",X"81",X"13",X"05",X"81",X"19",X"E2",X"00",X"E0",X"00",X"E4",X"00",
		X"1F",X"2C",X"01",X"0D",X"1D",X"10",X"10",X"10",X"07",X"1F",X"00",X"05",X"81",X"13",X"05",X"81",
		X"19",X"D6",X"00",X"D4",X"00",X"D8",X"00",X"1F",X"2C",X"01",X"0D",X"1D",X"10",X"10",X"10",X"07",
		X"3E",X"00",X"05",X"81",X"13",X"05",X"81",X"1F",X"40",X"1F",X"00",X"1D",X"10",X"10",X"10",X"07",
		X"07",X"00",X"05",X"81",X"13",X"05",X"81",X"19",X"AC",X"01",X"AA",X"01",X"AE",X"01",X"1F",X"2C",
		X"01",X"0D",X"1D",X"10",X"10",X"10",X"07",X"3E",X"00",X"05",X"81",X"13",X"05",X"81",X"1F",X"40",
		X"1F",X"00",X"1D",X"10",X"10",X"10",X"07",X"07",X"00",X"05",X"81",X"13",X"05",X"81",X"19",X"AC",
		X"01",X"AA",X"01",X"AE",X"01",X"1F",X"2C",X"01",X"0D",X"1D",X"10",X"10",X"10",X"07",X"3E",X"00",
		X"05",X"81",X"13",X"05",X"81",X"19",X"1D",X"01",X"1B",X"01",X"1F",X"01",X"1F",X"2C",X"01",X"0D",
		X"1D",X"10",X"10",X"10",X"07",X"1F",X"00",X"05",X"81",X"13",X"05",X"81",X"19",X"40",X"01",X"3E",
		X"01",X"42",X"01",X"1F",X"2C",X"01",X"0D",X"1D",X"10",X"10",X"10",X"07",X"1F",X"00",X"05",X"81",
		X"13",X"05",X"81",X"19",X"53",X"01",X"51",X"01",X"55",X"01",X"1F",X"2C",X"01",X"0D",X"1D",X"10",
		X"10",X"10",X"07",X"1F",X"00",X"05",X"81",X"13",X"05",X"81",X"19",X"1D",X"01",X"1B",X"01",X"1F",
		X"01",X"1F",X"2C",X"01",X"0D",X"1D",X"10",X"10",X"10",X"07",X"1F",X"00",X"05",X"81",X"13",X"05",
		X"81",X"19",X"D6",X"00",X"D4",X"00",X"D8",X"00",X"1F",X"2C",X"01",X"0D",X"1D",X"10",X"10",X"10",
		X"07",X"1F",X"00",X"05",X"81",X"13",X"05",X"81",X"19",X"E2",X"00",X"E0",X"00",X"E4",X"00",X"1F",
		X"2C",X"01",X"0D",X"1D",X"10",X"10",X"10",X"07",X"1F",X"00",X"05",X"81",X"13",X"05",X"81",X"19",
		X"D6",X"00",X"D4",X"00",X"D8",X"00",X"1F",X"2C",X"01",X"0D",X"1D",X"10",X"10",X"10",X"07",X"1F",
		X"00",X"05",X"81",X"13",X"05",X"81",X"19",X"AA",X"00",X"A8",X"00",X"AC",X"00",X"1F",X"2C",X"01",
		X"0D",X"1D",X"10",X"10",X"10",X"07",X"1F",X"00",X"05",X"81",X"13",X"05",X"81",X"19",X"BE",X"00",
		X"BC",X"00",X"C0",X"00",X"1F",X"2C",X"01",X"0D",X"1D",X"10",X"10",X"10",X"07",X"1F",X"00",X"05",
		X"81",X"13",X"05",X"81",X"19",X"D6",X"00",X"D4",X"00",X"D8",X"00",X"1F",X"2C",X"01",X"0D",X"1D",
		X"10",X"10",X"10",X"07",X"1F",X"00",X"05",X"81",X"13",X"05",X"81",X"19",X"BE",X"00",X"BC",X"00",
		X"C0",X"00",X"1F",X"2C",X"01",X"0D",X"1D",X"10",X"10",X"10",X"07",X"1F",X"00",X"05",X"81",X"13",
		X"05",X"81",X"1F",X"40",X"1F",X"00",X"1D",X"10",X"10",X"10",X"07",X"07",X"00",X"05",X"81",X"13",
		X"05",X"81",X"19",X"7D",X"01",X"7B",X"01",X"7F",X"01",X"1F",X"2C",X"01",X"0D",X"1D",X"10",X"10",
		X"10",X"07",X"3E",X"00",X"05",X"81",X"13",X"05",X"81",X"1F",X"40",X"1F",X"00",X"1D",X"10",X"10",
		X"10",X"07",X"07",X"00",X"05",X"81",X"13",X"05",X"81",X"19",X"7D",X"01",X"7B",X"01",X"7F",X"01",
		X"1F",X"2C",X"01",X"0D",X"1D",X"10",X"10",X"10",X"07",X"3E",X"00",X"05",X"81",X"13",X"05",X"81",
		X"1F",X"40",X"1F",X"00",X"1D",X"10",X"10",X"10",X"07",X"07",X"00",X"05",X"81",X"13",X"05",X"81",
		X"19",X"7D",X"01",X"7B",X"01",X"7F",X"01",X"1F",X"2C",X"01",X"0D",X"1D",X"10",X"10",X"10",X"07",
		X"1F",X"00",X"05",X"81",X"13",X"05",X"81",X"19",X"AC",X"01",X"AA",X"01",X"AE",X"01",X"1F",X"2C",
		X"01",X"0D",X"1D",X"10",X"10",X"10",X"07",X"1F",X"00",X"05",X"81",X"13",X"05",X"81",X"19",X"C5",
		X"01",X"C3",X"01",X"C7",X"01",X"1F",X"2C",X"01",X"0D",X"1D",X"10",X"10",X"10",X"07",X"1F",X"00",
		X"05",X"81",X"13",X"05",X"81",X"19",X"7D",X"01",X"7B",X"01",X"7F",X"01",X"1F",X"2C",X"01",X"0D",
		X"1D",X"10",X"10",X"10",X"07",X"1F",X"00",X"05",X"81",X"13",X"05",X"81",X"19",X"1D",X"01",X"1B",
		X"01",X"1F",X"01",X"1F",X"2C",X"01",X"0D",X"1D",X"10",X"10",X"10",X"07",X"1F",X"00",X"05",X"81",
		X"13",X"05",X"81",X"19",X"2E",X"01",X"2C",X"01",X"30",X"01",X"1F",X"2C",X"01",X"0D",X"1D",X"10",
		X"10",X"10",X"07",X"1F",X"00",X"05",X"81",X"13",X"05",X"81",X"19",X"1D",X"01",X"1B",X"01",X"1F",
		X"01",X"1F",X"2C",X"01",X"0D",X"1D",X"10",X"10",X"10",X"07",X"1F",X"00",X"05",X"81",X"13",X"05",
		X"81",X"19",X"1D",X"01",X"1B",X"01",X"1F",X"01",X"1F",X"2C",X"01",X"0D",X"1D",X"10",X"10",X"10",
		X"07",X"1F",X"00",X"05",X"81",X"13",X"05",X"81",X"19",X"FE",X"00",X"FC",X"00",X"00",X"01",X"1F",
		X"2C",X"01",X"0D",X"1D",X"10",X"10",X"10",X"07",X"1F",X"00",X"05",X"81",X"13",X"05",X"81",X"19",
		X"E2",X"00",X"E0",X"00",X"E4",X"00",X"1F",X"2C",X"01",X"0D",X"1D",X"10",X"10",X"10",X"07",X"1F",
		X"00",X"05",X"81",X"13",X"05",X"81",X"19",X"D6",X"00",X"D4",X"00",X"D8",X"00",X"1F",X"2C",X"01",
		X"0D",X"1D",X"10",X"10",X"10",X"07",X"1F",X"00",X"05",X"81",X"13",X"05",X"81",X"19",X"E2",X"00",
		X"E0",X"00",X"E4",X"00",X"1F",X"2C",X"01",X"0D",X"1D",X"10",X"10",X"10",X"07",X"1F",X"00",X"05",
		X"81",X"13",X"05",X"81",X"19",X"FE",X"00",X"FC",X"00",X"00",X"01",X"1F",X"2C",X"01",X"0D",X"1D",
		X"10",X"10",X"10",X"07",X"1F",X"00",X"05",X"81",X"13",X"05",X"81",X"19",X"1D",X"01",X"1B",X"01",
		X"1F",X"01",X"1F",X"2C",X"01",X"0D",X"1D",X"10",X"10",X"10",X"07",X"1F",X"00",X"05",X"81",X"13",
		X"05",X"81",X"19",X"FE",X"00",X"FC",X"00",X"00",X"01",X"1F",X"2C",X"01",X"0D",X"1D",X"10",X"10",
		X"10",X"07",X"1F",X"00",X"05",X"81",X"13",X"05",X"81",X"19",X"1D",X"01",X"1B",X"01",X"1F",X"01",
		X"1F",X"2C",X"01",X"0D",X"1D",X"10",X"10",X"10",X"07",X"1F",X"00",X"05",X"81",X"13",X"05",X"81",
		X"19",X"40",X"01",X"3E",X"01",X"42",X"01",X"1F",X"2C",X"01",X"0D",X"1D",X"10",X"10",X"10",X"07",
		X"1F",X"00",X"05",X"81",X"13",X"05",X"81",X"19",X"53",X"01",X"51",X"01",X"55",X"01",X"1F",X"2C",
		X"01",X"0D",X"1D",X"10",X"10",X"10",X"07",X"1F",X"00",X"05",X"81",X"13",X"05",X"81",X"19",X"40",
		X"01",X"3E",X"01",X"42",X"01",X"1F",X"2C",X"01",X"0D",X"1D",X"10",X"10",X"10",X"07",X"1F",X"00",
		X"05",X"81",X"13",X"05",X"81",X"19",X"53",X"01",X"51",X"01",X"55",X"01",X"1F",X"2C",X"01",X"0D",
		X"1D",X"10",X"10",X"10",X"07",X"1F",X"00",X"05",X"81",X"13",X"05",X"81",X"19",X"7D",X"01",X"7B",
		X"01",X"7F",X"01",X"1F",X"2C",X"01",X"0D",X"1D",X"10",X"10",X"10",X"07",X"1F",X"00",X"05",X"81",
		X"13",X"05",X"81",X"19",X"AC",X"01",X"AA",X"01",X"AE",X"01",X"1F",X"2C",X"01",X"0D",X"1D",X"10",
		X"10",X"10",X"07",X"1F",X"00",X"05",X"81",X"13",X"05",X"81",X"19",X"7D",X"01",X"7B",X"01",X"7F",
		X"01",X"1F",X"2C",X"01",X"0D",X"1D",X"10",X"10",X"10",X"07",X"1F",X"00",X"05",X"81",X"13",X"05",
		X"81",X"19",X"AC",X"01",X"AA",X"01",X"AE",X"01",X"1F",X"2C",X"01",X"0D",X"1D",X"10",X"10",X"10",
		X"07",X"1F",X"00",X"05",X"81",X"13",X"05",X"81",X"19",X"C5",X"01",X"C3",X"01",X"C7",X"01",X"1F",
		X"2C",X"01",X"0D",X"1D",X"10",X"10",X"10",X"07",X"1F",X"00",X"05",X"81",X"13",X"05",X"81",X"19",
		X"FC",X"01",X"FA",X"01",X"FE",X"01",X"1F",X"2C",X"01",X"0D",X"1D",X"10",X"10",X"10",X"07",X"1F",
		X"00",X"05",X"81",X"13",X"05",X"81",X"19",X"3B",X"02",X"39",X"02",X"3D",X"02",X"1F",X"2C",X"01",
		X"0D",X"1D",X"10",X"10",X"10",X"07",X"1F",X"00",X"05",X"81",X"13",X"05",X"81",X"19",X"AC",X"01",
		X"AA",X"01",X"AE",X"01",X"1F",X"2C",X"01",X"0D",X"1D",X"10",X"10",X"10",X"07",X"1F",X"00",X"05",
		X"81",X"13",X"05",X"81",X"19",X"C5",X"01",X"C3",X"01",X"C7",X"01",X"1F",X"2C",X"01",X"0D",X"1D",
		X"10",X"10",X"10",X"07",X"1F",X"00",X"05",X"81",X"13",X"05",X"81",X"19",X"7D",X"01",X"7B",X"01",
		X"7F",X"01",X"1F",X"2C",X"01",X"0D",X"1D",X"10",X"10",X"10",X"07",X"1F",X"00",X"05",X"81",X"13",
		X"05",X"81",X"19",X"AC",X"01",X"AA",X"01",X"AE",X"01",X"1F",X"2C",X"01",X"0D",X"1D",X"10",X"10",
		X"10",X"07",X"1F",X"00",X"05",X"81",X"13",X"05",X"81",X"19",X"53",X"01",X"51",X"01",X"55",X"01",
		X"1F",X"2C",X"01",X"0D",X"1D",X"10",X"10",X"10",X"07",X"1F",X"00",X"05",X"81",X"13",X"05",X"81",
		X"19",X"7D",X"01",X"7B",X"01",X"7F",X"01",X"1F",X"2C",X"01",X"0D",X"1D",X"10",X"10",X"10",X"07",
		X"1F",X"00",X"05",X"81",X"13",X"05",X"81",X"19",X"40",X"01",X"3E",X"01",X"42",X"01",X"1F",X"2C",
		X"01",X"0D",X"1D",X"10",X"10",X"10",X"07",X"1F",X"00",X"05",X"81",X"13",X"05",X"81",X"19",X"53",
		X"01",X"51",X"01",X"55",X"01",X"1F",X"2C",X"01",X"0D",X"1D",X"10",X"10",X"10",X"07",X"1F",X"00",
		X"05",X"81",X"13",X"05",X"81",X"19",X"AC",X"01",X"AA",X"01",X"AE",X"01",X"1F",X"2C",X"01",X"0D",
		X"1D",X"10",X"10",X"10",X"07",X"3E",X"00",X"05",X"81",X"13",X"05",X"81",X"1F",X"40",X"1F",X"00",
		X"1D",X"10",X"10",X"10",X"07",X"07",X"00",X"05",X"81",X"13",X"05",X"81",X"19",X"AC",X"01",X"AA",
		X"01",X"AE",X"01",X"1F",X"2C",X"01",X"0D",X"1D",X"10",X"10",X"10",X"07",X"7D",X"00",X"05",X"81",
		X"13",X"05",X"81",X"10",X"18",X"02",X"02",X"02",X"02",X"02",X"02",X"06",X"04",X"11",X"81",X"19",
		X"9B",X"0A",X"99",X"0A",X"9D",X"0A",X"1F",X"2C",X"01",X"0D",X"1D",X"10",X"10",X"10",X"07",X"7D",
		X"00",X"05",X"81",X"13",X"05",X"81",X"1F",X"40",X"1F",X"00",X"1D",X"10",X"10",X"10",X"07",X"3E",
		X"00",X"05",X"81",X"13",X"05",X"81",X"19",X"02",X"0A",X"00",X"0A",X"04",X"0A",X"1F",X"2C",X"01",
		X"0D",X"1D",X"10",X"10",X"10",X"07",X"7D",X"00",X"05",X"81",X"13",X"05",X"81",X"1F",X"40",X"1F",
		X"00",X"1D",X"10",X"10",X"10",X"07",X"3E",X"00",X"05",X"81",X"13",X"05",X"81",X"03",X"11",X"81",
		X"AE",X"06",X"05",X"11",X"81",X"19",X"9B",X"0A",X"99",X"0A",X"9D",X"0A",X"1F",X"2C",X"01",X"0D",
		X"1D",X"10",X"10",X"10",X"07",X"3E",X"00",X"05",X"81",X"13",X"05",X"81",X"1F",X"40",X"1F",X"00",
		X"1D",X"10",X"10",X"10",X"07",X"1F",X"00",X"05",X"81",X"13",X"05",X"81",X"19",X"02",X"0A",X"00",
		X"0A",X"04",X"0A",X"1F",X"2C",X"01",X"0D",X"1D",X"10",X"10",X"10",X"07",X"3E",X"00",X"05",X"81",
		X"13",X"05",X"81",X"1F",X"40",X"1F",X"00",X"1D",X"10",X"10",X"10",X"07",X"1F",X"00",X"05",X"81",
		X"13",X"05",X"81",X"03",X"11",X"81",X"AE",X"02",X"A8",X"19",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1D",X"10",X"10",X"10",X"18",X"03",X"03",X"02",X"03",X"03",X"03",X"1F",X"00",X"20",X"01",X"1B",
		X"1F",X"04",X"06",X"FF",X"03",X"81",X"0B",X"06",X"00",X"23",X"81",X"0B",X"07",X"00",X"25",X"81",
		X"01",X"03",X"03",X"81",X"F1",X"10",X"19",X"00",X"00",X"00",X"00",X"00",X"00",X"1D",X"10",X"10",
		X"10",X"18",X"03",X"03",X"02",X"03",X"03",X"03",X"1F",X"00",X"20",X"01",X"1B",X"10",X"04",X"06",
		X"FF",X"03",X"81",X"0B",X"06",X"00",X"23",X"81",X"0B",X"07",X"00",X"25",X"81",X"01",X"03",X"03",
		X"81",X"F1",X"10",X"19",X"06",X"06",X"05",X"05",X"07",X"00",X"1D",X"10",X"10",X"10",X"18",X"02",
		X"02",X"02",X"03",X"03",X"03",X"1F",X"00",X"20",X"01",X"1B",X"1F",X"04",X"06",X"FF",X"03",X"81");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
