library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_PGM_1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_PGM_1 is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"F3",X"97",X"32",X"00",X"50",X"32",X"C0",X"50",X"DB",X"02",X"ED",X"56",X"31",X"F0",X"4F",X"06",
		X"64",X"DB",X"03",X"CD",X"65",X"03",X"3A",X"00",X"3F",X"00",X"97",X"21",X"00",X"4C",X"01",X"04",
		X"00",X"77",X"23",X"10",X"FC",X"32",X"C0",X"50",X"0D",X"20",X"F6",X"DB",X"04",X"DB",X"0A",X"CD",
		X"ED",X"06",X"C3",X"07",X"02",X"07",X"37",X"00",X"F5",X"C5",X"D5",X"E5",X"3A",X"3B",X"4C",X"A7",
		X"CA",X"32",X"01",X"DB",X"07",X"11",X"F2",X"4F",X"01",X"62",X"50",X"21",X"8C",X"4E",X"DB",X"08",
		X"DB",X"0A",X"DB",X"0B",X"3E",X"06",X"00",X"F5",X"DB",X"14",X"DB",X"15",X"F1",X"F5",X"3A",X"A8",
		X"4C",X"A7",X"28",X"26",X"3A",X"A9",X"4C",X"A7",X"28",X"20",X"7E",X"3D",X"CB",X"4E",X"20",X"02",
		X"C6",X"04",X"12",X"13",X"23",X"7E",X"12",X"13",X"23",X"3E",X"E6",X"96",X"C6",X"26",X"02",X"03",
		X"23",X"7E",X"D6",X"18",X"D6",X"F8",X"ED",X"44",X"18",X"0D",X"7E",X"12",X"13",X"23",X"7E",X"12",
		X"13",X"23",X"7E",X"02",X"03",X"23",X"7E",X"02",X"03",X"23",X"F1",X"3D",X"20",X"BF",X"3A",X"A7",
		X"4C",X"A7",X"20",X"6C",X"21",X"CA",X"4E",X"3A",X"34",X"4F",X"47",X"97",X"32",X"34",X"4F",X"78",
		X"06",X"04",X"0F",X"F5",X"30",X"53",X"E5",X"11",X"05",X"00",X"19",X"E5",X"5E",X"23",X"56",X"D5",
		X"2B",X"2B",X"7E",X"4F",X"EE",X"01",X"77",X"2B",X"2B",X"7E",X"CB",X"2F",X"CB",X"2F",X"ED",X"44",
		X"EB",X"CB",X"7F",X"16",X"00",X"5F",X"3E",X"FF",X"28",X"02",X"2F",X"15",X"A9",X"E6",X"01",X"20",
		X"03",X"11",X"00",X"00",X"D5",X"11",X"FB",X"01",X"CB",X"41",X"28",X"03",X"11",X"01",X"02",X"CD",
		X"5B",X"01",X"D1",X"E1",X"19",X"D1",X"EB",X"73",X"23",X"72",X"EB",X"11",X"FB",X"01",X"CB",X"41",
		X"20",X"03",X"11",X"01",X"02",X"CD",X"44",X"01",X"E1",X"11",X"F4",X"FF",X"19",X"F1",X"10",X"A2",
		X"21",X"09",X"4C",X"35",X"23",X"36",X"00",X"23",X"35",X"20",X"03",X"CD",X"32",X"07",X"CD",X"32",
		X"07",X"CD",X"8B",X"01",X"E1",X"D1",X"C1",X"97",X"32",X"00",X"50",X"3C",X"32",X"00",X"50",X"F1",
		X"FB",X"C9",X"3A",X"A7",X"4C",X"A7",X"20",X"D8",X"21",X"F2",X"4F",X"97",X"06",X"0C",X"77",X"23",
		X"10",X"FC",X"18",X"CC",X"C5",X"0E",X"02",X"06",X"06",X"D5",X"1A",X"86",X"77",X"13",X"2B",X"10",
		X"F9",X"11",X"E6",X"FF",X"19",X"D1",X"0D",X"20",X"EE",X"C1",X"C9",X"C5",X"0E",X"02",X"06",X"06",
		X"D5",X"1A",X"96",X"ED",X"44",X"77",X"13",X"2B",X"10",X"F7",X"11",X"E6",X"FF",X"19",X"D1",X"0D",
		X"20",X"EC",X"C1",X"C9",X"F5",X"C5",X"06",X"FF",X"3A",X"0D",X"4C",X"CB",X"77",X"20",X"02",X"06",
		X"BF",X"CD",X"81",X"02",X"A0",X"32",X"0D",X"4C",X"D1",X"F1",X"C9",X"F5",X"DB",X"1E",X"E5",X"DB",
		X"1F",X"3A",X"AC",X"4C",X"A7",X"20",X"19",X"CD",X"B3",X"01",X"3A",X"00",X"50",X"E6",X"10",X"00",
		X"00",X"00",X"3A",X"A8",X"4C",X"A7",X"20",X"08",X"3A",X"40",X"50",X"E6",X"10",X"00",X"00",X"00",
		X"E1",X"F1",X"C9",X"3A",X"0F",X"4C",X"A7",X"28",X"2C",X"3A",X"00",X"50",X"CB",X"6F",X"C0",X"97",
		X"32",X"0F",X"4C",X"3C",X"32",X"15",X"4C",X"CD",X"ED",X"06",X"3E",X"16",X"CD",X"7A",X"09",X"21",
		X"36",X"4C",X"7E",X"FE",X"99",X"C8",X"C6",X"01",X"27",X"77",X"3E",X"0F",X"32",X"0C",X"4C",X"3E",
		X"01",X"32",X"07",X"50",X"C9",X"21",X"0C",X"4C",X"35",X"C0",X"36",X"01",X"3A",X"00",X"50",X"CB",
		X"6F",X"C8",X"97",X"32",X"07",X"50",X"3C",X"32",X"0F",X"4C",X"C9",X"7C",X"02",X"02",X"02",X"80",
		X"00",X"7E",X"02",X"02",X"02",X"02",X"82",X"97",X"32",X"03",X"50",X"3C",X"32",X"93",X"4C",X"32",
		X"A3",X"4C",X"32",X"0F",X"4C",X"32",X"17",X"4C",X"21",X"48",X"4C",X"36",X"4D",X"23",X"36",X"4F",
		X"23",X"36",X"42",X"23",X"36",X"00",X"23",X"36",X"01",X"23",X"36",X"00",X"CD",X"F0",X"20",X"3A",
		X"40",X"50",X"CB",X"7F",X"3E",X"01",X"28",X"01",X"97",X"32",X"A8",X"4C",X"C3",X"00",X"12",X"FB",
		X"3E",X"0B",X"CD",X"7A",X"09",X"CD",X"A1",X"03",X"C3",X"93",X"3B",X"F5",X"E6",X"F0",X"0F",X"0F",
		X"0F",X"0F",X"47",X"F1",X"E6",X"0F",X"4F",X"C9",X"F5",X"3A",X"8A",X"4C",X"18",X"04",X"F5",X"3A",
		X"4B",X"4D",X"C5",X"47",X"3A",X"A8",X"4C",X"A7",X"28",X"0F",X"78",X"06",X"00",X"FE",X"01",X"28",
		X"01",X"04",X"78",X"32",X"03",X"50",X"32",X"A9",X"4C",X"C1",X"F1",X"C9",X"3A",X"8A",X"4C",X"18",
		X"03",X"3A",X"4B",X"4D",X"C5",X"47",X"3A",X"A8",X"4C",X"A7",X"28",X"1B",X"78",X"FE",X"01",X"28",
		X"16",X"3A",X"40",X"50",X"47",X"E6",X"0F",X"4F",X"78",X"E6",X"10",X"07",X"B1",X"4F",X"3A",X"00",
		X"50",X"E6",X"80",X"0F",X"B1",X"C1",X"C9",X"3A",X"00",X"50",X"E6",X"0F",X"4F",X"3A",X"40",X"50",
		X"E6",X"60",X"18",X"F0",X"CD",X"BD",X"02",X"06",X"1E",X"CD",X"72",X"03",X"C9",X"CD",X"D1",X"02",
		X"CD",X"E2",X"02",X"CD",X"15",X"03",X"C9",X"CD",X"F3",X"02",X"CD",X"04",X"03",X"CD",X"1A",X"03",
		X"C9",X"21",X"C2",X"43",X"01",X"01",X"1C",X"CD",X"20",X"03",X"21",X"E2",X"43",X"01",X"01",X"1C",
		X"18",X"3E",X"21",X"02",X"40",X"01",X"01",X"1C",X"CD",X"20",X"03",X"21",X"22",X"40",X"01",X"01",
		X"1C",X"18",X"2D",X"21",X"C2",X"47",X"01",X"01",X"1C",X"CD",X"20",X"03",X"21",X"E2",X"47",X"01",
		X"01",X"1C",X"18",X"1C",X"21",X"02",X"44",X"01",X"01",X"1C",X"CD",X"20",X"03",X"21",X"22",X"44",
		X"01",X"01",X"1C",X"18",X"0B",X"21",X"40",X"40",X"18",X"03",X"21",X"40",X"44",X"01",X"04",X"80",
		X"77",X"23",X"10",X"FC",X"32",X"C0",X"50",X"0D",X"20",X"F6",X"C9",X"06",X"3C",X"CD",X"49",X"03",
		X"3E",X"01",X"32",X"00",X"50",X"FB",X"3A",X"0A",X"4C",X"A7",X"20",X"F1",X"32",X"C0",X"50",X"3C",
		X"32",X"0A",X"4C",X"10",X"E8",X"0D",X"20",X"E3",X"C9",X"F5",X"3A",X"36",X"4C",X"A7",X"20",X"02",
		X"F1",X"C9",X"31",X"F0",X"4F",X"97",X"32",X"14",X"4C",X"32",X"3B",X"4C",X"3E",X"01",X"32",X"00",
		X"50",X"FB",X"C3",X"85",X"19",X"C5",X"0E",X"00",X"0D",X"20",X"FD",X"32",X"C0",X"50",X"10",X"F8",
		X"C1",X"C9",X"F5",X"C5",X"78",X"32",X"09",X"4C",X"3E",X"01",X"32",X"00",X"50",X"FB",X"32",X"C0",
		X"50",X"3A",X"09",X"4C",X"A7",X"20",X"F1",X"C1",X"F1",X"C9",X"F5",X"3E",X"01",X"32",X"0A",X"4C",
		X"3E",X"01",X"32",X"00",X"50",X"FB",X"32",X"C0",X"50",X"3A",X"0A",X"4C",X"A7",X"20",X"F1",X"F1",
		X"C9",X"06",X"02",X"CD",X"72",X"03",X"D5",X"E5",X"21",X"B1",X"4C",X"11",X"04",X"00",X"06",X"03",
		X"4E",X"B9",X"28",X"05",X"19",X"10",X"F9",X"18",X"1D",X"2B",X"3A",X"14",X"4C",X"A7",X"28",X"06",
		X"3A",X"15",X"4C",X"A7",X"28",X"10",X"3E",X"01",X"32",X"00",X"50",X"32",X"01",X"50",X"FB",X"7E",
		X"32",X"C0",X"50",X"A7",X"20",X"E4",X"E1",X"D1",X"C9",X"D5",X"3E",X"01",X"32",X"08",X"4C",X"1A",
		X"CD",X"F3",X"03",X"13",X"1A",X"CD",X"F3",X"03",X"13",X"97",X"32",X"08",X"4C",X"1A",X"CD",X"F3",
		X"03",X"D1",X"C9",X"C5",X"CD",X"4B",X"02",X"78",X"CD",X"01",X"04",X"79",X"CD",X"01",X"04",X"C1",
		X"C9",X"D5",X"5F",X"3A",X"08",X"4C",X"57",X"A7",X"28",X"09",X"7B",X"A7",X"3E",X"00",X"20",X"03",
		X"1E",X"D0",X"7A",X"32",X"08",X"4C",X"7B",X"C6",X"30",X"D1",X"D5",X"77",X"E5",X"11",X"00",X"04",
		X"19",X"3A",X"02",X"4C",X"77",X"E1",X"3A",X"A3",X"4C",X"A7",X"11",X"FF",X"FF",X"28",X"03",X"11",
		X"E0",X"FF",X"19",X"D1",X"C9",X"C5",X"D5",X"CD",X"4B",X"02",X"78",X"FE",X"0A",X"16",X"30",X"38",
		X"02",X"16",X"37",X"82",X"CD",X"1A",X"04",X"79",X"FE",X"0A",X"16",X"30",X"38",X"02",X"16",X"37",
		X"82",X"CD",X"1A",X"04",X"D1",X"C1",X"C9",X"77",X"19",X"10",X"FC",X"C9",X"F5",X"4E",X"81",X"77",
		X"F1",X"19",X"10",X"F8",X"C9",X"C5",X"01",X"01",X"00",X"18",X"04",X"C5",X"01",X"E0",X"FF",X"ED",
		X"43",X"04",X"4C",X"F5",X"22",X"06",X"4C",X"C5",X"0E",X"32",X"F3",X"ED",X"40",X"1A",X"0D",X"ED",
		X"40",X"FB",X"C1",X"FE",X"FF",X"28",X"15",X"77",X"C5",X"E5",X"01",X"00",X"04",X"09",X"3A",X"02",
		X"4C",X"77",X"E1",X"C1",X"13",X"ED",X"4B",X"04",X"4C",X"09",X"18",X"DB",X"13",X"0E",X"14",X"F3",
		X"ED",X"40",X"1A",X"0C",X"13",X"ED",X"40",X"FB",X"FE",X"FF",X"20",X"03",X"F1",X"C1",X"C9",X"FE",
		X"FE",X"20",X"09",X"2A",X"06",X"4C",X"23",X"22",X"06",X"4C",X"18",X"BB",X"32",X"02",X"4C",X"18",
		X"B6",X"D5",X"EB",X"97",X"67",X"6F",X"3C",X"32",X"01",X"50",X"32",X"00",X"50",X"00",X"D5",X"16",
		X"00",X"5F",X"19",X"D1",X"13",X"10",X"F6",X"32",X"C0",X"50",X"0D",X"20",X"F0",X"D1",X"19",X"7C",
		X"21",X"CB",X"37",X"E9",X"E5",X"11",X"04",X"05",X"21",X"9A",X"42",X"CD",X"6B",X"04",X"3A",X"03",
		X"4C",X"32",X"02",X"4C",X"3E",X"01",X"32",X"08",X"4C",X"3A",X"36",X"4C",X"21",X"BA",X"41",X"CD",
		X"F3",X"03",X"E1",X"C9",X"FF",X"05",X"43",X"52",X"45",X"44",X"49",X"54",X"FF",X"FF",X"21",X"DD",
		X"43",X"11",X"96",X"4C",X"18",X"06",X"21",X"FD",X"43",X"11",X"99",X"4C",X"32",X"02",X"4C",X"CD",
		X"D9",X"03",X"C9",X"F5",X"C5",X"D5",X"E5",X"07",X"16",X"00",X"5F",X"3A",X"14",X"4C",X"FE",X"01",
		X"CA",X"5E",X"05",X"21",X"88",X"05",X"19",X"01",X"98",X"4C",X"11",X"A0",X"4C",X"3A",X"4B",X"4D",
		X"FE",X"01",X"28",X"06",X"01",X"9B",X"4C",X"11",X"A2",X"4C",X"0A",X"86",X"27",X"02",X"2B",X"0B",
		X"0A",X"8E",X"27",X"02",X"0B",X"0A",X"CE",X"00",X"27",X"02",X"EB",X"CD",X"63",X"05",X"E1",X"D1",
		X"C1",X"F1",X"C9",X"3A",X"92",X"4C",X"57",X"0A",X"BA",X"D8",X"7E",X"A7",X"C8",X"2B",X"34",X"3A",
		X"4B",X"4D",X"FE",X"01",X"28",X"05",X"CD",X"9E",X"05",X"18",X"03",X"CD",X"95",X"05",X"3E",X"12",
		X"CD",X"7A",X"09",X"23",X"36",X"00",X"C9",X"50",X"00",X"00",X"55",X"00",X"66",X"00",X"77",X"00",
		X"88",X"00",X"99",X"01",X"00",X"E5",X"01",X"9F",X"4C",X"21",X"D6",X"43",X"18",X"07",X"E5",X"01",
		X"A1",X"4C",X"21",X"F6",X"43",X"0A",X"A7",X"28",X"19",X"FE",X"07",X"38",X"02",X"3E",X"06",X"47",
		X"36",X"01",X"2B",X"3E",X"09",X"77",X"E5",X"11",X"00",X"04",X"19",X"77",X"23",X"77",X"E1",X"2B",
		X"10",X"EE",X"E1",X"C9",X"21",X"C5",X"43",X"01",X"4D",X"4D",X"18",X"06",X"21",X"E5",X"43",X"01",
		X"50",X"4D",X"11",X"E1",X"05",X"CD",X"65",X"04",X"11",X"F9",X"FF",X"19",X"0A",X"CD",X"F3",X"03",
		X"C9",X"20",X"20",X"44",X"4C",X"49",X"42",X"FF",X"FF",X"D5",X"E5",X"11",X"00",X"06",X"21",X"CD",
		X"43",X"CD",X"65",X"04",X"11",X"0A",X"06",X"21",X"ED",X"43",X"CD",X"65",X"04",X"E1",X"D1",X"C9",
		X"FF",X"08",X"71",X"70",X"6F",X"6E",X"6D",X"6C",X"FF",X"FF",X"77",X"76",X"75",X"74",X"73",X"72",
		X"FF",X"FF",X"F5",X"C5",X"D5",X"E5",X"3E",X"01",X"32",X"3B",X"4C",X"32",X"A7",X"4C",X"06",X"18",
		X"21",X"8C",X"4E",X"11",X"31",X"06",X"1A",X"77",X"13",X"23",X"10",X"FA",X"E1",X"D1",X"C1",X"F1",
		X"C9",X"D0",X"08",X"95",X"F8",X"D4",X"08",X"85",X"F8",X"D8",X"08",X"76",X"F8",X"DC",X"08",X"96",
		X"E8",X"E0",X"08",X"86",X"E8",X"E4",X"08",X"76",X"E8",X"11",X"53",X"06",X"21",X"24",X"40",X"CD",
		X"65",X"04",X"C9",X"FF",X"07",X"20",X"20",X"52",X"4F",X"42",X"41",X"4C",X"20",X"45",X"52",X"41",
		X"57",X"54",X"46",X"4F",X"53",X"20",X"34",X"38",X"39",X"31",X"20",X"40",X"FF",X"FF",X"3E",X"A8",
		X"32",X"A6",X"4C",X"21",X"02",X"44",X"11",X"01",X"00",X"3E",X"12",X"06",X"3C",X"CD",X"57",X"04",
		X"21",X"02",X"40",X"22",X"A4",X"4C",X"11",X"01",X"00",X"3E",X"60",X"06",X"15",X"CD",X"57",X"04",
		X"21",X"22",X"40",X"06",X"15",X"CD",X"57",X"04",X"11",X"AB",X"06",X"21",X"17",X"40",X"CD",X"65",
		X"04",X"11",X"E1",X"05",X"21",X"37",X"40",X"CD",X"65",X"04",X"C9",X"FF",X"08",X"20",X"20",X"20",
		X"54",X"49",X"45",X"5A",X"FF",X"FF",X"21",X"26",X"4E",X"35",X"C0",X"32",X"26",X"4E",X"3A",X"14",
		X"4C",X"A7",X"C0",X"2A",X"A4",X"4C",X"34",X"11",X"20",X"00",X"19",X"34",X"21",X"A6",X"4C",X"35",
		X"20",X"05",X"3E",X"01",X"32",X"A5",X"4E",X"7E",X"FE",X"32",X"30",X"05",X"3E",X"03",X"CD",X"7A",
		X"09",X"7E",X"E6",X"07",X"C0",X"2A",X"A4",X"4C",X"23",X"22",X"A4",X"4C",X"C9",X"F5",X"C5",X"E5",
		X"97",X"21",X"08",X"4D",X"06",X"40",X"77",X"23",X"10",X"FC",X"21",X"08",X"4D",X"11",X"50",X"50",
		X"01",X"10",X"00",X"ED",X"B0",X"21",X"08",X"4D",X"11",X"40",X"50",X"01",X"10",X"00",X"ED",X"B0",
		X"3E",X"04",X"32",X"4A",X"50",X"3E",X"05",X"32",X"45",X"50",X"32",X"4F",X"50",X"21",X"B0",X"4C",
		X"06",X"0C",X"97",X"77",X"23",X"10",X"FC",X"32",X"01",X"50",X"3C",X"32",X"01",X"50",X"E1",X"C1",
		X"F1",X"C9",X"F5",X"C5",X"D5",X"E5",X"06",X"00",X"11",X"04",X"00",X"21",X"B0",X"4C",X"7E",X"FE",
		X"00",X"C4",X"59",X"07",X"19",X"04",X"7E",X"FE",X"00",X"C4",X"59",X"07",X"19",X"04",X"7E",X"FE",
		X"00",X"C4",X"59",X"07",X"E1",X"D1",X"C1",X"F1",X"C9",X"DB",X"64",X"C5",X"D5",X"E5",X"78",X"32",
		X"49",X"4D",X"23",X"23",X"E5",X"DB",X"6B",X"5E",X"23",X"56",X"DB",X"64",X"1A",X"D5",X"5F",X"DB",
		X"6B",X"7B",X"E6",X"E0",X"07",X"07",X"07",X"21",X"82",X"07",X"5F",X"07",X"83",X"16",X"00",X"5F",
		X"19",X"E9",X"C3",X"9E",X"07",X"C3",X"C0",X"07",X"C3",X"E3",X"07",X"C3",X"14",X"08",X"C3",X"42",
		X"08",X"C3",X"B8",X"08",X"C3",X"BC",X"08",X"C3",X"C5",X"08",X"E1",X"D1",X"C1",X"C9",X"E1",X"CD",
		X"B0",X"0C",X"E6",X"1F",X"23",X"F5",X"CD",X"B0",X"0C",X"47",X"F1",X"23",X"E5",X"CD",X"20",X"09",
		X"07",X"16",X"00",X"5F",X"21",X"08",X"4D",X"19",X"70",X"23",X"36",X"00",X"D1",X"C3",X"6A",X"07",
		X"E1",X"CD",X"B0",X"0C",X"E6",X"1F",X"23",X"F5",X"CD",X"B0",X"0C",X"4F",X"23",X"CD",X"B0",X"0C",
		X"47",X"F1",X"23",X"E5",X"07",X"16",X"00",X"5F",X"21",X"BC",X"4C",X"19",X"71",X"23",X"70",X"D1",
		X"C3",X"6A",X"07",X"E1",X"CD",X"B0",X"0C",X"E6",X"1F",X"23",X"F5",X"CD",X"B0",X"0C",X"4F",X"23",
		X"CD",X"B0",X"0C",X"47",X"F1",X"23",X"E5",X"F5",X"07",X"16",X"00",X"5F",X"21",X"08",X"4D",X"19",
		X"E5",X"7E",X"23",X"6E",X"67",X"09",X"44",X"4D",X"E1",X"70",X"23",X"71",X"F1",X"CD",X"20",X"09",
		X"D1",X"C3",X"6A",X"07",X"E1",X"CD",X"B0",X"0C",X"E6",X"1F",X"23",X"F5",X"CD",X"B0",X"0C",X"47",
		X"F1",X"23",X"E5",X"07",X"16",X"00",X"5F",X"21",X"08",X"4D",X"19",X"7E",X"B8",X"28",X"0D",X"E1",
		X"CD",X"B0",X"0C",X"5F",X"23",X"CD",X"B0",X"0C",X"57",X"C3",X"BE",X"08",X"D1",X"13",X"13",X"C3",
		X"6A",X"07",X"E1",X"CD",X"B0",X"0C",X"E6",X"1F",X"23",X"F5",X"CD",X"B0",X"0C",X"47",X"23",X"CD",
		X"B0",X"0C",X"4F",X"F1",X"23",X"E5",X"F5",X"07",X"16",X"00",X"5F",X"21",X"08",X"4D",X"19",X"97",
		X"BE",X"28",X"06",X"35",X"F1",X"D1",X"C3",X"6A",X"07",X"78",X"E6",X"E0",X"07",X"07",X"07",X"07",
		X"16",X"00",X"5F",X"21",X"BC",X"4C",X"19",X"5E",X"23",X"56",X"F1",X"E5",X"07",X"D5",X"16",X"00",
		X"5F",X"21",X"08",X"4D",X"19",X"D1",X"1A",X"77",X"13",X"78",X"E6",X"1F",X"32",X"48",X"4D",X"79",
		X"07",X"D5",X"16",X"00",X"5F",X"21",X"08",X"4D",X"19",X"D1",X"1A",X"13",X"47",X"79",X"CD",X"20",
		X"09",X"0C",X"70",X"23",X"36",X"00",X"23",X"3A",X"48",X"4D",X"3D",X"32",X"48",X"4D",X"20",X"EA",
		X"E1",X"72",X"2B",X"73",X"D1",X"C3",X"6A",X"07",X"E1",X"C3",X"9A",X"07",X"D1",X"13",X"E1",X"73",
		X"23",X"72",X"C3",X"9A",X"07",X"E1",X"E1",X"3A",X"49",X"4D",X"07",X"07",X"16",X"00",X"5F",X"21",
		X"B0",X"4C",X"19",X"46",X"23",X"4E",X"79",X"07",X"16",X"00",X"5F",X"21",X"C9",X"4C",X"19",X"7E",
		X"FE",X"00",X"28",X"10",X"57",X"2B",X"5E",X"97",X"77",X"23",X"77",X"3A",X"49",X"4D",X"CD",X"D8",
		X"09",X"C3",X"9A",X"07",X"3A",X"49",X"4D",X"F5",X"3C",X"47",X"07",X"80",X"F5",X"06",X"00",X"CD",
		X"20",X"09",X"21",X"08",X"4D",X"F1",X"07",X"5F",X"16",X"00",X"19",X"72",X"23",X"72",X"F1",X"07",
		X"07",X"5F",X"21",X"B0",X"4C",X"19",X"36",X"00",X"C3",X"9A",X"07",X"78",X"32",X"4F",X"50",X"C9",
		X"FE",X"1B",X"28",X"F7",X"FE",X"0A",X"D0",X"F5",X"C5",X"E5",X"D5",X"11",X"66",X"09",X"07",X"83",
		X"5F",X"7A",X"CE",X"00",X"57",X"1A",X"67",X"13",X"1A",X"6F",X"97",X"D1",X"E9",X"C6",X"05",X"C6",
		X"05",X"3C",X"C6",X"04",X"26",X"50",X"C6",X"50",X"6F",X"70",X"18",X"16",X"C6",X"02",X"C6",X"03",
		X"C6",X"02",X"C6",X"04",X"C6",X"02",X"26",X"50",X"C6",X"50",X"6F",X"78",X"CD",X"4B",X"02",X"71",
		X"23",X"70",X"E1",X"C1",X"F1",X"C9",X"09",X"56",X"09",X"54",X"09",X"42",X"09",X"41",X"09",X"52",
		X"09",X"50",X"09",X"3F",X"09",X"4E",X"09",X"4C",X"09",X"3D",X"F5",X"C5",X"D5",X"E5",X"F5",X"3A",
		X"14",X"4C",X"FE",X"01",X"20",X"0A",X"3A",X"15",X"4C",X"FE",X"01",X"28",X"03",X"F1",X"18",X"43",
		X"F1",X"32",X"4A",X"4D",X"4F",X"07",X"07",X"16",X"00",X"5F",X"21",X"EB",X"09",X"19",X"E5",X"23",
		X"23",X"46",X"23",X"7E",X"C5",X"E5",X"07",X"07",X"16",X"00",X"5F",X"21",X"B0",X"4C",X"19",X"7E",
		X"B8",X"38",X"07",X"20",X"09",X"23",X"7E",X"B9",X"28",X"04",X"3E",X"01",X"18",X"01",X"97",X"E1",
		X"C1",X"A7",X"E1",X"28",X"0E",X"5E",X"23",X"56",X"23",X"23",X"7E",X"CD",X"D8",X"09",X"3E",X"01",
		X"32",X"01",X"50",X"E1",X"D1",X"C1",X"F1",X"C9",X"D5",X"07",X"07",X"16",X"00",X"5F",X"21",X"B0",
		X"4C",X"19",X"70",X"23",X"71",X"23",X"D1",X"73",X"23",X"72",X"C9",X"4B",X"0A",X"02",X"00",X"5B",
		X"0A",X"02",X"00",X"6B",X"0A",X"01",X"01",X"8C",X"0A",X"03",X"01",X"9C",X"0A",X"02",X"00",X"49",
		X"10",X"01",X"00",X"78",X"0C",X"01",X"00",X"09",X"0B",X"02",X"00",X"29",X"0B",X"02",X"00",X"E9",
		X"0A",X"02",X"00",X"79",X"0A",X"02",X"00",X"49",X"0B",X"01",X"00",X"86",X"0B",X"04",X"00",X"A0",
		X"0B",X"04",X"00",X"BA",X"0B",X"03",X"01",X"12",X"0C",X"03",X"00",X"F9",X"0B",X"01",X"00",X"27",
		X"0C",X"01",X"00",X"5E",X"0C",X"04",X"01",X"D6",X"0B",X"03",X"00",X"CD",X"0A",X"03",X"00",X"94",
		X"0C",X"01",X"02",X"B5",X"0A",X"03",X"01",X"CD",X"0A",X"03",X"00",X"03",X"07",X"00",X"05",X"01",
		X"01",X"02",X"01",X"40",X"00",X"01",X"60",X"BF",X"53",X"0A",X"0A",X"03",X"07",X"00",X"BF",X"01",
		X"01",X"02",X"01",X"40",X"00",X"FF",X"60",X"05",X"63",X"0A",X"E0",X"06",X"0F",X"04",X"FF",X"05",
		X"10",X"46",X"80",X"FF",X"66",X"00",X"71",X"0A",X"E0",X"03",X"09",X"00",X"00",X"01",X"0D",X"02",
		X"0A",X"43",X"80",X"FF",X"40",X"00",X"02",X"63",X"00",X"81",X"0A",X"E0",X"06",X"0F",X"04",X"0F",
		X"05",X"07",X"11",X"06",X"51",X"00",X"FF",X"71",X"00",X"94",X"0A",X"E0",X"03",X"07",X"10",X"03",
		X"01",X"04",X"02",X"00",X"00",X"28",X"40",X"00",X"FB",X"60",X"0A",X"A6",X"0A",X"50",X"00",X"FF",
		X"70",X"00",X"A4",X"0A",X"E0",X"06",X"0F",X"11",X"03",X"04",X"08",X"05",X"02",X"04",X"28",X"44",
		X"80",X"FF",X"45",X"80",X"00",X"64",X"0A",X"BF",X"0A",X"45",X"84",X"7B",X"E0",X"03",X"07",X"10",
		X"01",X"01",X"08",X"02",X"00",X"00",X"28",X"40",X"00",X"FB",X"41",X"C0",X"FF",X"60",X"0A",X"D7",
		X"0A",X"50",X"00",X"FF",X"70",X"00",X"51",X"8E",X"E0",X"03",X"02",X"00",X"18",X"01",X"05",X"02",
		X"00",X"10",X"02",X"43",X"00",X"02",X"41",X"00",X"FF",X"63",X"0A",X"F3",X"0A",X"03",X"04",X"00",
		X"18",X"50",X"00",X"FF",X"70",X"00",X"F3",X"0A",X"E0",X"03",X"08",X"00",X"18",X"01",X"02",X"02",
		X"00",X"10",X"01",X"43",X"80",X"00",X"41",X"80",X"00",X"63",X"10",X"13",X"0B",X"03",X"08",X"00",
		X"18",X"50",X"00",X"FF",X"70",X"00",X"07",X"8F",X"E0",X"03",X"08",X"00",X"18",X"01",X"28",X"02",
		X"00",X"10",X"01",X"43",X"80",X"00",X"41",X"80",X"7B",X"63",X"10",X"33",X"0B",X"03",X"08",X"00",
		X"18",X"50",X"00",X"FF",X"70",X"00",X"27",X"8F",X"E0",X"03",X"07",X"00",X"00",X"01",X"08",X"02",
		X"00",X"04",X"04",X"05",X"00",X"06",X"07",X"07",X"0F",X"08",X"00",X"09",X"07",X"10",X"7F",X"40",
		X"00",X"08",X"44",X"00",X"04",X"47",X"00",X"FD",X"50",X"00",X"FF",X"70",X"00",X"5F",X"0B",X"40",
		X"7F",X"41",X"00",X"FC",X"45",X"00",X"F8",X"48",X"00",X"04",X"50",X"00",X"FF",X"70",X"00",X"71",
		X"0B",X"06",X"00",X"09",X"00",X"E0",X"03",X"0A",X"02",X"00",X"20",X"05",X"0F",X"16",X"15",X"13",
		X"00",X"93",X"02",X"00",X"73",X"00",X"91",X"0B",X"56",X"00",X"FF",X"76",X"00",X"91",X"0B",X"E0",
		X"03",X"0A",X"02",X"00",X"20",X"9B",X"0F",X"16",X"3A",X"13",X"00",X"93",X"02",X"00",X"73",X"00",
		X"AB",X"0B",X"56",X"00",X"FF",X"76",X"00",X"AB",X"0B",X"E0",X"06",X"0F",X"04",X"10",X"05",X"01",
		X"11",X"04",X"14",X"10",X"44",X"00",X"04",X"54",X"00",X"FE",X"74",X"00",X"C4",X"0B",X"51",X"00",
		X"FE",X"71",X"00",X"C2",X"0B",X"E0",X"01",X"00",X"02",X"00",X"10",X"05",X"03",X"0B",X"00",X"F0",
		X"40",X"00",X"E0",X"60",X"50",X"E0",X"0B",X"40",X"00",X"10",X"60",X"A0",X"E7",X"0B",X"41",X"00",
		X"01",X"50",X"00",X"FF",X"70",X"00",X"DE",X"0B",X"E0",X"00",X"7F",X"01",X"00",X"02",X"00",X"03",
		X"03",X"10",X"05",X"50",X"00",X"FF",X"70",X"00",X"03",X"0C",X"43",X"00",X"01",X"63",X"0A",X"0A",
		X"0C",X"E0",X"00",X"1C",X"01",X"00",X"02",X"00",X"03",X"0F",X"10",X"0C",X"50",X"00",X"FF",X"40",
		X"00",X"68",X"70",X"00",X"1C",X"0C",X"E0",X"03",X"08",X"00",X"18",X"01",X"0A",X"02",X"00",X"10",
		X"03",X"43",X"00",X"02",X"41",X"80",X"FF",X"63",X"10",X"31",X"0C",X"03",X"08",X"00",X"18",X"50",
		X"00",X"FF",X"70",X"00",X"31",X"0C",X"03",X"0A",X"20",X"44",X"0F",X"16",X"1D",X"13",X"00",X"93",
		X"02",X"00",X"73",X"00",X"4F",X"0C",X"56",X"00",X"FF",X"76",X"00",X"4F",X"0C",X"E0",X"06",X"0A",
		X"05",X"00",X"21",X"A5",X"0E",X"17",X"20",X"14",X"00",X"94",X"22",X"04",X"74",X"00",X"69",X"0C",
		X"57",X"00",X"FF",X"77",X"00",X"69",X"0C",X"E0",X"03",X"0A",X"10",X"04",X"01",X"00",X"02",X"00",
		X"00",X"0A",X"40",X"00",X"05",X"41",X"80",X"00",X"60",X"5A",X"82",X"0C",X"50",X"00",X"FF",X"70",
		X"00",X"80",X"0C",X"E0",X"09",X"01",X"08",X"00",X"1B",X"03",X"22",X"B9",X"0C",X"18",X"78",X"15",
		X"00",X"95",X"42",X"07",X"75",X"00",X"A1",X"0C",X"58",X"00",X"FF",X"78",X"00",X"A1",X"0C",X"E0",
		X"D5",X"DB",X"64",X"5E",X"DB",X"6B",X"7B",X"D1",X"C9",X"03",X"96",X"01",X"03",X"00",X"00",X"03",
		X"6A",X"01",X"03",X"00",X"00",X"03",X"60",X"02",X"03",X"00",X"00",X"03",X"AC",X"02",X"03",X"00",
		X"00",X"03",X"80",X"01",X"03",X"00",X"00",X"03",X"AE",X"01",X"03",X"00",X"00",X"03",X"C8",X"01",
		X"03",X"00",X"00",X"03",X"00",X"00",X"03",X"00",X"00",X"03",X"C8",X"01",X"03",X"00",X"00",X"03",
		X"E0",X"01",X"03",X"00",X"00",X"03",X"20",X"02",X"03",X"00",X"00",X"03",X"58",X"05",X"03",X"00",
		X"00",X"03",X"00",X"00",X"03",X"00",X"00",X"03",X"00",X"00",X"03",X"00",X"00",X"03",X"00",X"00",
		X"03",X"00",X"00",X"03",X"00",X"00",X"03",X"00",X"00",X"03",X"00",X"00",X"03",X"00",X"00",X"03",
		X"B5",X"00",X"03",X"00",X"00",X"03",X"B5",X"00",X"03",X"00",X"00",X"03",X"B5",X"00",X"03",X"00",
		X"00",X"03",X"C0",X"00",X"03",X"00",X"00",X"03",X"B5",X"00",X"03",X"B5",X"00",X"03",X"B5",X"00",
		X"03",X"B5",X"00",X"03",X"00",X"00",X"03",X"00",X"00",X"03",X"00",X"00",X"03",X"00",X"00",X"03",
		X"10",X"01",X"03",X"00",X"00",X"03",X"10",X"01",X"03",X"00",X"00",X"03",X"10",X"01",X"03",X"00",
		X"00",X"03",X"1E",X"01",X"03",X"00",X"00",X"03",X"10",X"01",X"03",X"10",X"01",X"03",X"10",X"01",
		X"03",X"10",X"01",X"03",X"00",X"00",X"03",X"00",X"00",X"03",X"30",X"01",X"03",X"00",X"00",X"03",
		X"56",X"01",X"03",X"00",X"00",X"03",X"C0",X"00",X"03",X"00",X"00",X"03",X"CB",X"00",X"03",X"00",
		X"00",X"03",X"30",X"01",X"03",X"00",X"00",X"03",X"56",X"01",X"03",X"00",X"00",X"03",X"C0",X"00",
		X"03",X"00",X"00",X"03",X"CB",X"00",X"03",X"00",X"00",X"03",X"2C",X"03",X"03",X"2C",X"03",X"03",
		X"2C",X"03",X"03",X"00",X"00",X"03",X"90",X"03",X"33",X"00",X"00",X"03",X"00",X"03",X"03",X"00",
		X"03",X"03",X"00",X"03",X"03",X"00",X"00",X"03",X"2C",X"03",X"03",X"00",X"00",X"03",X"D4",X"02",
		X"03",X"00",X"00",X"03",X"2C",X"03",X"03",X"00",X"00",X"03",X"D4",X"02",X"03",X"00",X"00",X"03",
		X"2C",X"03",X"03",X"00",X"00",X"03",X"D4",X"02",X"03",X"D4",X"02",X"03",X"5C",X"03",X"03",X"58",
		X"05",X"03",X"00",X"00",X"03",X"00",X"00",X"03",X"30",X"01",X"03",X"00",X"00",X"03",X"56",X"01",
		X"03",X"00",X"00",X"03",X"B5",X"00",X"03",X"00",X"00",X"03",X"B5",X"00",X"03",X"00",X"00",X"03",
		X"B5",X"00",X"03",X"00",X"00",X"03",X"56",X"01",X"03",X"00",X"00",X"03",X"30",X"01",X"03",X"00",
		X"00",X"32",X"00",X"00",X"02",X"E8",X"01",X"01",X"00",X"00",X"02",X"83",X"01",X"01",X"00",X"00",
		X"02",X"45",X"01",X"01",X"00",X"00",X"06",X"7A",X"00",X"06",X"00",X"00",X"04",X"91",X"00",X"02",
		X"00",X"00",X"0A",X"7A",X"00",X"12",X"00",X"00",X"03",X"23",X"01",X"01",X"00",X"00",X"03",X"00",
		X"01",X"01",X"00",X"00",X"05",X"3C",X"00",X"01",X"00",X"00",X"05",X"78",X"00",X"01",X"00",X"00",
		X"05",X"55",X"00",X"01",X"00",X"00",X"05",X"C8",X"00",X"01",X"00",X"00",X"03",X"4B",X"01",X"01",
		X"00",X"00",X"03",X"78",X"00",X"01",X"00",X"00",X"03",X"55",X"00",X"01",X"00",X"00",X"02",X"C3",
		X"00",X"01",X"00",X"00",X"02",X"41",X"00",X"02",X"00",X"00",X"03",X"3C",X"00",X"02",X"00",X"00",
		X"02",X"37",X"00",X"02",X"00",X"00",X"02",X"32",X"00",X"02",X"00",X"00",X"02",X"2F",X"00",X"02",
		X"00",X"00",X"03",X"2C",X"00",X"04",X"81",X"00",X"03",X"00",X"00",X"04",X"34",X"01",X"03",X"00",
		X"00",X"02",X"B0",X"02",X"02",X"0E",X"03",X"01",X"00",X"00",X"02",X"A1",X"03",X"01",X"00",X"00",
		X"04",X"A9",X"03",X"02",X"00",X"00",X"02",X"00",X"01",X"02",X"00",X"00",X"02",X"F3",X"02",X"03",
		X"00",X"00",X"02",X"CD",X"00",X"03",X"00",X"00",X"01",X"B7",X"00",X"03",X"00",X"00",X"05",X"6A",
		X"00",X"02",X"00",X"00",X"03",X"93",X"00",X"03",X"00",X"00",X"03",X"52",X"00",X"02",X"00",X"00",
		X"03",X"32",X"00",X"02",X"00",X"00",X"03",X"2B",X"00",X"02",X"00",X"00",X"03",X"32",X"00",X"02",
		X"00",X"00",X"08",X"64",X"00",X"07",X"7F",X"01",X"01",X"00",X"00",X"02",X"32",X"02",X"02",X"64",
		X"02",X"02",X"96",X"02",X"01",X"00",X"00",X"01",X"C8",X"06",X"01",X"00",X"00",X"01",X"C8",X"06",
		X"01",X"00",X"00",X"01",X"C8",X"06",X"01",X"00",X"00",X"01",X"C8",X"06",X"01",X"00",X"00",X"01",
		X"C8",X"06",X"01",X"00",X"00",X"01",X"C8",X"06",X"01",X"00",X"00",X"01",X"C8",X"06",X"01",X"00",
		X"00",X"03",X"00",X"05",X"03",X"F0",X"00",X"01",X"00",X"00",X"02",X"1E",X"01",X"01",X"00",X"00",
		X"02",X"1E",X"02",X"01",X"00",X"00",X"02",X"1E",X"03",X"01",X"00",X"00",X"02",X"1E",X"04",X"01",
		X"00",X"00",X"02",X"1E",X"05",X"01",X"00",X"00",X"02",X"1E",X"06",X"01",X"00",X"00",X"05",X"1E",
		X"07",X"01",X"00",X"00",X"02",X"1E",X"06",X"01",X"00",X"00",X"02",X"1E",X"05",X"01",X"00",X"00",
		X"02",X"1E",X"04",X"01",X"00",X"00",X"02",X"1E",X"03",X"01",X"00",X"00",X"02",X"1E",X"02",X"01",
		X"00",X"00",X"02",X"1E",X"01",X"01",X"00",X"00",X"05",X"64",X"00",X"01",X"96",X"03",X"04",X"00",
		X"00",X"01",X"C8",X"03",X"04",X"00",X"00",X"01",X"64",X"03",X"04",X"00",X"00",X"01",X"96",X"02",
		X"04",X"00",X"00",X"01",X"C8",X"02",X"04",X"00",X"00",X"01",X"64",X"02",X"04",X"00",X"00",X"01",
		X"96",X"01",X"04",X"00",X"00",X"01",X"C8",X"01",X"04",X"00",X"00",X"01",X"64",X"01",X"04",X"00",
		X"00",X"01",X"96",X"00",X"04",X"00",X"00",X"01",X"C8",X"00",X"04",X"00",X"00",X"01",X"64",X"00",
		X"04",X"00",X"00",X"01",X"78",X"01",X"03",X"00",X"00",X"01",X"A0",X"01",X"03",X"00",X"00",X"01",
		X"4B",X"01",X"03",X"00",X"00",X"01",X"78",X"00",X"03",X"00",X"00",X"01",X"A0",X"00",X"03",X"00",
		X"00",X"01",X"4B",X"00",X"01",X"5A",X"01",X"02",X"00",X"00",X"01",X"78",X"01",X"02",X"00",X"00",
		X"01",X"32",X"01",X"02",X"00",X"00",X"01",X"5A",X"00",X"02",X"00",X"00",X"01",X"78",X"00",X"02",
		X"00",X"00",X"01",X"32",X"00",X"02",X"00",X"00",X"01",X"3C",X"01",X"01",X"00",X"00",X"01",X"50",
		X"01",X"01",X"00",X"01",X"1E",X"01",X"01",X"00",X"00",X"01",X"3C",X"00",X"01",X"00",X"00",X"01",
		X"50",X"00",X"01",X"00",X"00",X"01",X"1E",X"00",X"00",X"03",X"07",X"00",X"05",X"01",X"00",X"02",
		X"00",X"40",X"80",X"00",X"60",X"BF",X"51",X"10",X"E0",X"CD",X"ED",X"06",X"3E",X"01",X"32",X"AC",
		X"4C",X"32",X"00",X"50",X"32",X"4B",X"4D",X"CD",X"5E",X"02",X"FB",X"06",X"01",X"97",X"32",X"14",
		X"4C",X"C5",X"CD",X"B4",X"02",X"CD",X"12",X"06",X"11",X"A9",X"97",X"42",X"A7",X"10",X"1E",X"F6",
		X"42",X"B6",X"10",X"27",X"D6",X"42",X"E0",X"10",X"39",X"F6",X"42",X"05",X"11",X"30",X"57",X"42",
		X"42",X"11",X"28",X"57",X"42",X"4C",X"11",X"3C",X"57",X"42",X"57",X"11",X"50",X"57",X"42",X"61",
		X"11",X"4A",X"57",X"42",X"6C",X"11",X"FF",X"20",X"20",X"53",X"55",X"50",X"45",X"52",X"20",X"20",
		X"47",X"4C",X"4F",X"42",X"FF",X"FF",X"41",X"4C",X"4C",X"45",X"20",X"46",X"52",X"55",X"45",X"43",
		X"48",X"54",X"45",X"20",X"53",X"55",X"43",X"48",X"45",X"4E",X"FF",X"FE",X"5A",X"55",X"4D",X"20",
		X"4E",X"41",X"45",X"43",X"48",X"53",X"54",X"45",X"4E",X"20",X"42",X"49",X"4C",X"44",X"FF",X"FF",
		X"54",X"41",X"53",X"54",X"45",X"20",X"52",X"55",X"46",X"54",X"20",X"4C",X"49",X"46",X"54",X"20",
		X"FF",X"FE",X"48",X"45",X"42",X"45",X"4C",X"3E",X"4F",X"42",X"45",X"4E",X"20",X"55",X"4E",X"54",
		X"45",X"4E",X"20",X"FF",X"FF",X"4D",X"49",X"54",X"20",X"44",X"45",X"52",X"20",X"54",X"41",X"53",
		X"54",X"45",X"20",X"20",X"20",X"20",X"20",X"20",X"FF",X"FE",X"41",X"55",X"46",X"20",X"44",X"49",
		X"45",X"20",X"56",X"45",X"52",X"46",X"4F",X"4C",X"47",X"45",X"52",X"20",X"20",X"FF",X"FE",X"53",
		X"50",X"52",X"49",X"4E",X"47",X"45",X"4E",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"FF",X"FF",X"2E",X"2E",X"2E",X"47",X"41",X"54",X"4F",X"52",X"FF",X"FF",X"2E",X"2E",X"2E",X"46",
		X"52",X"4F",X"47",X"47",X"59",X"FF",X"FF",X"2E",X"2E",X"2E",X"42",X"55",X"4E",X"4E",X"59",X"FF",
		X"FF",X"2E",X"2E",X"2E",X"4D",X"4F",X"4E",X"4B",X"45",X"59",X"FF",X"FF",X"2E",X"2E",X"2E",X"50",
		X"4F",X"52",X"4B",X"45",X"52",X"FF",X"FF",X"F5",X"D5",X"E5",X"21",X"D7",X"4E",X"35",X"20",X"11",
		X"36",X"05",X"2B",X"35",X"28",X"09",X"21",X"DC",X"46",X"7E",X"EE",X"0D",X"77",X"18",X"02",X"36",
		X"01",X"21",X"33",X"4C",X"97",X"BE",X"28",X"03",X"35",X"18",X"2E",X"21",X"32",X"4C",X"97",X"34",
		X"CB",X"46",X"28",X"02",X"3E",X"03",X"32",X"02",X"4C",X"2A",X"34",X"4C",X"5E",X"23",X"56",X"23",
		X"D5",X"5E",X"23",X"56",X"23",X"3A",X"02",X"4C",X"A7",X"7E",X"20",X"06",X"23",X"22",X"34",X"4C",
		X"3E",X"05",X"32",X"33",X"4C",X"E1",X"CD",X"6B",X"04",X"E1",X"D1",X"F1",X"C9",X"06",X"97",X"34",
		X"CB",X"46",X"28",X"02",X"3E",X"03",X"32",X"02",X"4C",X"2A",X"34",X"4C",X"5E",X"23",X"56",X"23",
		X"D5",X"5E",X"23",X"56",X"23",X"3A",X"02",X"4C",X"A7",X"7E",X"20",X"06",X"23",X"22",X"34",X"4C",
		X"3E",X"05",X"32",X"33",X"4C",X"E1",X"CD",X"6B",X"04",X"E1",X"D1",X"F1",X"C9",X"06",X"8B",X"B0",
		X"E5",X"D5",X"C5",X"4F",X"21",X"80",X"14",X"46",X"04",X"05",X"28",X"0E",X"23",X"5E",X"23",X"56",
		X"23",X"DD",X"1A",X"86",X"23",X"BE",X"20",X"16",X"10",X"F2",X"AF",X"ED",X"47",X"79",X"C1",X"D1",
		X"E1",X"C3",X"7F",X"3B",X"45",X"FF",X"06",X"20",X"54",X"49",X"48",X"FF",X"FF",X"F5",X"C5",X"97",
		X"CD",X"B4",X"02",X"3E",X"06",X"CD",X"1A",X"03",X"CD",X"12",X"06",X"11",X"E5",X"12",X"21",X"A6",
		X"42",X"CD",X"6B",X"04",X"11",X"13",X"12",X"21",X"07",X"40",X"CD",X"65",X"04",X"11",X"F6",X"12",
		X"21",X"90",X"43",X"CD",X"65",X"04",X"11",X"00",X"13",X"21",X"70",X"42",X"CD",X"6B",X"04",X"11",
		X"14",X"13",X"21",X"B2",X"42",X"CD",X"6B",X"04",X"11",X"3A",X"13",X"21",X"B5",X"42",X"CD",X"6B",
		X"04",X"3A",X"40",X"50",X"E6",X"80",X"21",X"CC",X"42",X"11",X"58",X"13",X"28",X"03",X"11",X"69",
		X"13",X"CD",X"6B",X"04",X"32",X"C0",X"50",X"3A",X"80",X"50",X"E6",X"3F",X"4F",X"21",X"50",X"43",
		X"06",X"06",X"0F",X"11",X"4E",X"13",X"30",X"03",X"11",X"53",X"13",X"E5",X"CD",X"6B",X"04",X"E1",
		X"23",X"10",X"EF",X"79",X"E6",X"03",X"EE",X"03",X"C6",X"33",X"32",X"B0",X"42",X"79",X"E6",X"1C",
		X"EE",X"1C",X"0F",X"0F",X"4F",X"C6",X"31",X"32",X"92",X"40",X"0C",X"41",X"21",X"33",X"42",X"36",
		X"1E",X"21",X"13",X"42",X"11",X"E0",X"FF",X"3E",X"16",X"CD",X"57",X"04",X"3E",X"08",X"91",X"28",
		X"06",X"47",X"3E",X"17",X"CD",X"57",X"04",X"36",X"1F",X"3A",X"40",X"50",X"CB",X"77",X"20",X"91",
		X"C1",X"F1",X"C3",X"6D",X"10",X"FF",X"09",X"43",X"4F",X"4E",X"46",X"49",X"47",X"55",X"52",X"41",
		X"54",X"49",X"4F",X"4E",X"FF",X"FF",X"FF",X"04",X"31",X"32",X"33",X"34",X"35",X"36",X"FF",X"FF",
		X"FF",X"06",X"47",X"4C",X"4F",X"42",X"53",X"20",X"50",X"45",X"52",X"20",X"43",X"52",X"45",X"44",
		X"49",X"54",X"FF",X"FF",X"44",X"49",X"46",X"46",X"49",X"43",X"55",X"4C",X"54",X"59",X"20",X"4C",
		X"45",X"56",X"45",X"4C",X"FF",X"FE",X"45",X"41",X"53",X"59",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"48",X"41",X"52",X"44",X"FF",X"FF",X"41",X"54",X"54",X"52",X"41",X"43",
		X"54",X"20",X"4D",X"4F",X"44",X"45",X"20",X"53",X"4F",X"55",X"4E",X"44",X"FF",X"FF",X"4F",X"4E",
		X"20",X"FF",X"FF",X"4F",X"46",X"46",X"FF",X"FF",X"FF",X"0E",X"20",X"54",X"41",X"42",X"4C",X"45",
		X"20",X"4D",X"4F",X"44",X"45",X"4C",X"20",X"FF",X"FF",X"FF",X"0E",X"55",X"50",X"52",X"49",X"47",
		X"48",X"54",X"20",X"4D",X"4F",X"44",X"45",X"4C",X"FF",X"FF",X"F5",X"C5",X"97",X"CD",X"B4",X"02",
		X"CD",X"12",X"06",X"11",X"F1",X"13",X"21",X"86",X"42",X"CD",X"6B",X"04",X"21",X"00",X"40",X"11",
		X"AD",X"4C",X"CD",X"39",X"14",X"21",X"00",X"44",X"13",X"CD",X"39",X"14",X"21",X"00",X"4C",X"13",
		X"CD",X"39",X"14",X"01",X"AD",X"4C",X"3E",X"03",X"21",X"70",X"43",X"11",X"01",X"14",X"F5",X"E5",
		X"CD",X"6B",X"04",X"D5",X"11",X"1F",X"14",X"0A",X"E6",X"0F",X"28",X"03",X"11",X"2C",X"14",X"CD",
		X"6B",X"04",X"11",X"40",X"FF",X"19",X"D1",X"CD",X"6B",X"04",X"D5",X"11",X"1F",X"14",X"0A",X"E6",
		X"F0",X"28",X"03",X"11",X"2C",X"14",X"CD",X"6B",X"04",X"D1",X"E1",X"23",X"23",X"F1",X"03",X"3D",
		X"20",X"CC",X"11",X"13",X"12",X"21",X"07",X"40",X"CD",X"65",X"04",X"CD",X"FB",X"11",X"C1",X"F1",
		X"C9",X"FF",X"09",X"53",X"54",X"41",X"54",X"49",X"43",X"20",X"52",X"41",X"4D",X"FF",X"06",X"FF",
		X"FF",X"34",X"4B",X"20",X"FF",X"FF",X"34",X"4E",X"20",X"FF",X"FF",X"34",X"4C",X"20",X"FF",X"FF",
		X"34",X"50",X"20",X"FF",X"FF",X"34",X"4D",X"20",X"FF",X"FF",X"34",X"52",X"20",X"FF",X"FF",X"FF",
		X"0E",X"4F",X"4B",X"20",X"20",X"20",X"20",X"20",X"FF",X"06",X"FF",X"FF",X"FF",X"FF",X"4E",X"4F",
		X"54",X"20",X"4F",X"4B",X"20",X"FF",X"06",X"FF",X"FF",X"97",X"01",X"04",X"00",X"E5",X"C5",X"F5",
		X"4E",X"77",X"AE",X"EB",X"B6",X"77",X"EB",X"71",X"F1",X"23",X"10",X"F3",X"C1",X"0D",X"20",X"EE",
		X"E1",X"3D",X"FE",X"FE",X"20",X"E4",X"C9",X"F5",X"C5",X"97",X"CD",X"B4",X"02",X"CD",X"12",X"06",
		X"11",X"A4",X"14",X"21",X"86",X"42",X"CD",X"6B",X"04",X"21",X"00",X"20",X"01",X"1F",X"FE",X"CD",
		X"C1",X"14",X"F5",X"21",X"00",X"00",X"01",X"20",X"00",X"CD",X"C1",X"14",X"01",X"FE",X"3F",X"11",
		X"09",X"00",X"3F",X"00",X"00",X"40",X"3F",X"00",X"00",X"80",X"3F",X"00",X"00",X"C0",X"3F",X"00",
		X"00",X"80",X"3F",X"00",X"00",X"40",X"3F",X"00",X"00",X"C0",X"3F",X"00",X"00",X"C0",X"3F",X"00",
		X"00",X"40",X"3F",X"00",X"00",X"FF",X"45",X"50",X"52",X"4F",X"4D",X"20",X"43",X"48",X"45",X"43",
		X"4B",X"FF",X"FF",X"FF",X"FF",X"55",X"32",X"20",X"FF",X"FF",X"FF",X"FF",X"CC",X"33",X"20",X"FF",
		X"FF",X"97",X"86",X"23",X"10",X"FC",X"0D",X"20",X"F9",X"C9",X"F5",X"CD",X"6B",X"04",X"0A",X"C1",
		X"11",X"1F",X"14",X"B8",X"28",X"04",X"11",X"2C",X"14",X"78",X"F5",X"CD",X"6B",X"04",X"3E",X"0B",
		X"32",X"02",X"4C",X"F1",X"CD",X"35",X"04",X"C9",X"F5",X"C5",X"97",X"32",X"3B",X"4C",X"32",X"A7",
		X"4C",X"CD",X"E9",X"05",X"3E",X"06",X"CD",X"1A",X"03",X"3E",X"13",X"CD",X"15",X"03",X"06",X"1E",
		X"CD",X"72",X"03",X"CD",X"FB",X"11",X"C1",X"F1",X"C3",X"6D",X"10",X"F5",X"C5",X"97",X"32",X"08",
		X"4C",X"11",X"AB",X"4C",X"21",X"AA",X"4C",X"3C",X"12",X"77",X"97",X"D5",X"E5",X"CD",X"B4",X"02",
		X"CD",X"12",X"06",X"11",X"06",X"16",X"21",X"86",X"42",X"CD",X"6B",X"04",X"11",X"15",X"16",X"21",
		X"8A",X"43",X"CD",X"6B",X"04",X"11",X"70",X"16",X"21",X"D5",X"42",X"CD",X"6B",X"04",X"11",X"13",
		X"12",X"21",X"07",X"40",X"CD",X"65",X"04",X"E1",X"D1",X"1A",X"E5",X"21",X"95",X"41",X"CD",X"F3",
		X"03",X"E1",X"06",X"70",X"CD",X"65",X"03",X"32",X"C0",X"50",X"3A",X"40",X"50",X"CB",X"77",X"CA",
		X"01",X"16",X"CB",X"6F",X"28",X"2C",X"3A",X"00",X"50",X"CB",X"47",X"28",X"06",X"CB",X"5F",X"28",
		X"11",X"18",X"E4",X"34",X"1A",X"C6",X"01",X"27",X"FE",X"25",X"20",X"03",X"3E",X"01",X"77",X"12",
		X"18",X"C7",X"35",X"1A",X"D6",X"01",X"27",X"A7",X"20",X"05",X"3E",X"18",X"77",X"3E",X"24",X"12",
		X"18",X"B7",X"1A",X"32",X"4D",X"4D",X"7E",X"32",X"4C",X"4D",X"00",X"FE",X"01",X"28",X"18",X"3D",
		X"47",X"3A",X"80",X"50",X"E6",X"1C",X"EE",X"1C",X"0F",X"0F",X"3C",X"4F",X"3E",X"01",X"81",X"10",
		X"FD",X"FE",X"10",X"38",X"02",X"3E",X"0F",X"32",X"4E",X"4D",X"97",X"32",X"A5",X"4E",X"32",X"16",
		X"4C",X"32",X"14",X"4C",X"3C",X"32",X"BB",X"4D",X"32",X"3C",X"4C",X"32",X"37",X"4C",X"D5",X"E5",
		X"CD",X"C3",X"27",X"CD",X"E9",X"05",X"11",X"13",X"12",X"21",X"07",X"40",X"CD",X"65",X"04",X"11",
		X"7D",X"16",X"21",X"28",X"40",X"CD",X"65",X"04",X"32",X"C0",X"50",X"3A",X"40",X"50",X"CB",X"77",
		X"28",X"0A",X"CB",X"6F",X"20",X"F2",X"CD",X"6E",X"06",X"CD",X"B0",X"2E",X"E1",X"D1",X"C3",X"1A",
		X"15",X"C1",X"F1",X"C3",X"6D",X"10",X"FF",X"09",X"4C",X"45",X"56",X"45",X"4C",X"20",X"43",X"48",
		X"45",X"43",X"4B",X"FF",X"FF",X"FF",X"06",X"4D",X"4F",X"56",X"45",X"20",X"4A",X"4F",X"59",X"53",
		X"54",X"49",X"43",X"4B",X"20",X"FF",X"0D",X"55",X"50",X"20",X"FF",X"06",X"4F",X"52",X"20",X"FF",
		X"08",X"44",X"4F",X"57",X"4E",X"FF",X"06",X"FF",X"FE",X"54",X"4F",X"20",X"53",X"45",X"4C",X"45",
		X"43",X"54",X"20",X"4C",X"45",X"56",X"45",X"4C",X"20",X"4E",X"55",X"4D",X"42",X"45",X"52",X"2E",
		X"FF",X"FE",X"48",X"49",X"54",X"20",X"FF",X"0E",X"43",X"41",X"4C",X"4C",X"20",X"FF",X"06",X"54",
		X"4F",X"20",X"53",X"45",X"54",X"55",X"50",X"20",X"4C",X"45",X"56",X"45",X"4C",X"2E",X"FF",X"FF",
		X"FF",X"07",X"4C",X"45",X"56",X"45",X"4C",X"20",X"4E",X"4F",X"3A",X"FF",X"FF",X"FF",X"06",X"59",
		X"41",X"4C",X"50",X"20",X"4F",X"54",X"FF",X"0E",X"20",X"4C",X"4C",X"41",X"43",X"FF",X"06",X"20",
		X"54",X"49",X"48",X"FF",X"FF",X"F5",X"C5",X"CD",X"ED",X"06",X"97",X"32",X"14",X"4C",X"CD",X"B4",
		X"02",X"CD",X"12",X"06",X"32",X"08",X"4C",X"11",X"AB",X"4C",X"21",X"AA",X"4C",X"12",X"77",X"D5",
		X"E5",X"11",X"2D",X"17",X"21",X"86",X"42",X"CD",X"6B",X"04",X"11",X"3C",X"17",X"21",X"8A",X"43",
		X"CD",X"6B",X"04",X"11",X"99",X"17",X"21",X"D5",X"42",X"CD",X"6B",X"04",X"11",X"13",X"12",X"21",
		X"07",X"40",X"CD",X"65",X"04",X"E1",X"D1",X"1A",X"E5",X"21",X"95",X"41",X"CD",X"F3",X"03",X"E1",
		X"06",X"70",X"CD",X"65",X"03",X"32",X"C0",X"50",X"3A",X"40",X"50",X"CB",X"77",X"28",X"36",X"CB",
		X"6F",X"28",X"2C",X"3A",X"00",X"50",X"CB",X"47",X"28",X"06",X"CB",X"5F",X"28",X"10",X"18",X"E5",
		X"34",X"1A",X"C6",X"01",X"27",X"FE",X"23",X"20",X"02",X"97",X"77",X"12",X"18",X"C9",X"35",X"1A",
		X"D6",X"01",X"27",X"FE",X"99",X"20",X"05",X"3E",X"16",X"77",X"3E",X"22",X"12",X"18",X"B8",X"7E",
		X"CD",X"7A",X"09",X"18",X"B2",X"CD",X"ED",X"06",X"C1",X"F1",X"C3",X"6D",X"10",X"FF",X"09",X"53",
		X"4F",X"55",X"4E",X"44",X"20",X"43",X"48",X"45",X"43",X"4B",X"FF",X"FF",X"FF",X"06",X"4D",X"4F",
		X"56",X"45",X"20",X"4A",X"4F",X"59",X"53",X"54",X"49",X"43",X"4B",X"20",X"FF",X"0D",X"55",X"50",
		X"20",X"FF",X"06",X"4F",X"52",X"20",X"FF",X"08",X"44",X"4F",X"57",X"4E",X"FF",X"06",X"FF",X"FE",
		X"54",X"4F",X"20",X"53",X"45",X"4C",X"45",X"43",X"54",X"20",X"53",X"4F",X"55",X"4E",X"44",X"20",
		X"4E",X"55",X"4D",X"42",X"45",X"52",X"2E",X"FF",X"FE",X"48",X"49",X"54",X"20",X"FF",X"0E",X"43",
		X"41",X"4C",X"4C",X"20",X"FF",X"06",X"54",X"4F",X"20",X"45",X"58",X"45",X"43",X"55",X"54",X"45",
		X"20",X"53",X"4F",X"55",X"4E",X"44",X"2E",X"FF",X"FF",X"FF",X"07",X"53",X"4F",X"55",X"4E",X"44",
		X"20",X"4E",X"4F",X"3A",X"FF",X"FF",X"F5",X"C5",X"97",X"CD",X"B4",X"02",X"CD",X"12",X"06",X"11",
		X"44",X"18",X"21",X"86",X"42",X"CD",X"6B",X"04",X"11",X"54",X"18",X"21",X"4A",X"43",X"CD",X"6B",
		X"04",X"11",X"9F",X"18",X"21",X"50",X"43",X"CD",X"6B",X"04",X"11",X"D0",X"18",X"21",X"10",X"41",
		X"CD",X"6B",X"04",X"11",X"13",X"12",X"21",X"07",X"40",X"CD",X"65",X"04",X"97",X"32",X"5A",X"50",
		X"06",X"04",X"11",X"40",X"18",X"21",X"56",X"50",X"1A",X"77",X"13",X"23",X"10",X"FA",X"3A",X"40",
		X"50",X"5F",X"2F",X"E6",X"0F",X"4F",X"3A",X"00",X"50",X"57",X"2F",X"E6",X"0F",X"47",X"CB",X"6B",
		X"20",X"02",X"CB",X"E0",X"CB",X"6A",X"20",X"02",X"CB",X"E8",X"CB",X"63",X"20",X"02",X"CB",X"E1",
		X"CB",X"7A",X"20",X"02",X"CB",X"E9",X"78",X"B1",X"3E",X"0A",X"20",X"01",X"97",X"32",X"5A",X"50",
		X"32",X"C0",X"50",X"78",X"21",X"50",X"47",X"CD",X"0C",X"19",X"79",X"21",X"10",X"45",X"CD",X"0C",
		X"19",X"3A",X"40",X"50",X"CB",X"77",X"20",X"B6",X"CD",X"ED",X"06",X"C1",X"F1",X"C3",X"6D",X"10",
		X"02",X"01",X"00",X"00",X"FF",X"09",X"42",X"55",X"54",X"54",X"4F",X"4E",X"20",X"43",X"48",X"45",
		X"43",X"4B",X"FF",X"FF",X"FF",X"06",X"20",X"20",X"20",X"44",X"45",X"50",X"52",X"45",X"53",X"53",
		X"45",X"44",X"20",X"42",X"55",X"54",X"54",X"4F",X"4E",X"53",X"FF",X"FE",X"20",X"20",X"20",X"41",
		X"52",X"45",X"20",X"48",X"49",X"47",X"48",X"4C",X"49",X"47",X"48",X"54",X"45",X"44",X"2E",X"FF",
		X"FE",X"FF",X"FE",X"FF",X"0D",X"50",X"4C",X"41",X"59",X"45",X"52",X"20",X"31",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"20",X"32",X"FF",X"FF",X"FF",
		X"0C",X"55",X"50",X"FF",X"FE",X"FF",X"FE",X"4C",X"45",X"46",X"54",X"FF",X"FE",X"FF",X"FE",X"52",
		X"49",X"47",X"48",X"54",X"FF",X"FE",X"FF",X"FE",X"44",X"4F",X"57",X"4E",X"FF",X"FE",X"FF",X"FE",
		X"43",X"41",X"4C",X"4C",X"FF",X"FE",X"FF",X"FE",X"43",X"4F",X"49",X"4E",X"49",X"4E",X"FF",X"FF",
		X"FF",X"0C",X"20",X"20",X"20",X"20",X"55",X"50",X"FF",X"FE",X"FF",X"FE",X"20",X"20",X"4C",X"45",
		X"46",X"54",X"FF",X"FE",X"FF",X"FE",X"20",X"52",X"49",X"47",X"48",X"54",X"FF",X"FE",X"FF",X"FE",
		X"20",X"20",X"44",X"4F",X"57",X"4E",X"FF",X"FE",X"FF",X"FE",X"20",X"20",X"43",X"41",X"4C",X"4C",
		X"FF",X"FE",X"FF",X"FE",X"45",X"4E",X"45",X"52",X"47",X"59",X"FF",X"FF",X"C5",X"06",X"06",X"0F",
		X"F5",X"C5",X"3E",X"0C",X"30",X"02",X"3E",X"08",X"11",X"E0",X"FF",X"06",X"06",X"CD",X"57",X"04",
		X"11",X"C2",X"00",X"19",X"C1",X"F1",X"10",X"E7",X"C1",X"C9",X"D5",X"FD",X"21",X"00",X"00",X"7E",
		X"16",X"00",X"5F",X"3E",X"06",X"32",X"00",X"4C",X"FD",X"19",X"2B",X"10",X"F2",X"32",X"C0",X"50",
		X"0D",X"20",X"EC",X"D1",X"FD",X"19",X"FD",X"29",X"FD",X"29",X"FD",X"E5",X"E1",X"CB",X"3C",X"CB",
		X"1D",X"00",X"21",X"5D",X"37",X"E9",X"CD",X"9E",X"19",X"CD",X"C6",X"1A",X"CD",X"C3",X"27",X"32",
		X"C0",X"50",X"CD",X"B0",X"2E",X"3A",X"A5",X"4E",X"FE",X"01",X"28",X"05",X"CD",X"98",X"1A",X"18",
		X"EB",X"CD",X"D4",X"1A",X"3A",X"3A",X"4C",X"FE",X"01",X"20",X"DE",X"CD",X"67",X"37",X"3A",X"36",
		X"4C",X"A7",X"CA",X"93",X"3B",X"97",X"32",X"14",X"4C",X"3C",X"32",X"15",X"4C",X"CD",X"00",X"1A",
		X"18",X"C4",X"11",X"00",X"00",X"ED",X"53",X"10",X"4C",X"ED",X"53",X"12",X"4C",X"C9",X"3A",X"80",
		X"50",X"E6",X"1C",X"EE",X"1C",X"0F",X"0F",X"C6",X"02",X"32",X"92",X"4C",X"32",X"31",X"01",X"3A",
		X"80",X"50",X"E6",X"03",X"EE",X"03",X"C6",X"03",X"21",X"38",X"4C",X"77",X"32",X"9F",X"4C",X"C3",
		X"B0",X"27",X"3A",X"37",X"4C",X"32",X"39",X"4C",X"FE",X"01",X"28",X"04",X"7E",X"32",X"A1",X"4C",
		X"F3",X"DB",X"64",X"3E",X"12",X"00",X"0F",X"47",X"DB",X"01",X"FB",X"97",X"21",X"96",X"4C",X"77",
		X"23",X"10",X"FC",X"32",X"16",X"4C",X"3C",X"32",X"A0",X"4C",X"32",X"A2",X"4C",X"32",X"4C",X"4D",
		X"32",X"4F",X"4D",X"32",X"4D",X"4D",X"32",X"50",X"4D",X"32",X"4E",X"4D",X"32",X"51",X"4D",X"C9",
		X"21",X"36",X"4C",X"E5",X"3E",X"01",X"32",X"4B",X"4D",X"CD",X"5E",X"02",X"97",X"CD",X"BD",X"02",
		X"CD",X"12",X"06",X"11",X"6D",X"1A",X"21",X"2F",X"42",X"CD",X"6B",X"04",X"E1",X"7E",X"E5",X"11",
		X"7F",X"1A",X"21",X"70",X"42",X"FE",X"01",X"28",X"06",X"11",X"89",X"1A",X"21",X"B0",X"42",X"CD",
		X"6B",X"04",X"E1",X"3A",X"40",X"50",X"47",X"CB",X"68",X"0E",X"01",X"28",X"0A",X"7E",X"FE",X"02",
		X"38",X"16",X"CB",X"70",X"20",X"12",X"0C",X"7E",X"91",X"27",X"77",X"79",X"32",X"37",X"4C",X"32",
		X"17",X"4C",X"3E",X"06",X"CD",X"7A",X"09",X"C9",X"32",X"C0",X"50",X"3A",X"03",X"4C",X"3C",X"FE",
		X"0E",X"38",X"02",X"3E",X"03",X"32",X"03",X"4C",X"CD",X"E4",X"04",X"18",X"B0",X"FF",X"06",X"50",
		X"52",X"45",X"53",X"53",X"FF",X"FE",X"FF",X"FE",X"53",X"54",X"41",X"52",X"54",X"FF",X"FF",X"31",
		X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"FF",X"FF",X"31",X"20",X"4F",X"52",X"20",X"32",X"20",
		X"50",X"4C",X"41",X"59",X"45",X"52",X"FF",X"FF",X"97",X"CD",X"BD",X"02",X"3A",X"4B",X"4D",X"01",
		X"51",X"4D",X"21",X"4F",X"4D",X"FE",X"01",X"20",X"06",X"01",X"4E",X"4D",X"21",X"4C",X"4D",X"7E",
		X"34",X"23",X"7E",X"C6",X"01",X"27",X"77",X"3A",X"80",X"50",X"E6",X"1C",X"EE",X"1C",X"0F",X"0F",
		X"3C",X"57",X"0A",X"82",X"02",X"C9",X"21",X"9F",X"4C",X"3A",X"4B",X"4D",X"FE",X"01",X"28",X"02",
		X"23",X"23",X"35",X"C9",X"97",X"CD",X"BD",X"02",X"32",X"A5",X"4E",X"21",X"4B",X"4D",X"3C",X"BE",
		X"11",X"9F",X"4C",X"28",X"03",X"11",X"A1",X"4C",X"1A",X"A7",X"28",X"41",X"3A",X"39",X"4C",X"FE",
		X"02",X"28",X"05",X"97",X"32",X"3A",X"4C",X"C9",X"7E",X"EE",X"03",X"77",X"CD",X"5E",X"02",X"97",
		X"32",X"3A",X"4C",X"3E",X"05",X"CD",X"7A",X"09",X"F5",X"97",X"E5",X"CD",X"BD",X"02",X"11",X"7B",
		X"1B",X"21",X"6F",X"42",X"CD",X"6B",X"04",X"E1",X"7E",X"FE",X"02",X"3E",X"32",X"28",X"01",X"3D",
		X"32",X"90",X"41",X"06",X"B4",X"CD",X"72",X"03",X"F1",X"CD",X"A1",X"03",X"C9",X"CD",X"41",X"1B",
		X"3A",X"39",X"4C",X"3D",X"32",X"39",X"4C",X"FE",X"01",X"28",X"BD",X"3E",X"01",X"32",X"3A",X"4C",
		X"C9",X"E5",X"11",X"66",X"1B",X"21",X"6F",X"42",X"CD",X"6B",X"04",X"E1",X"3E",X"01",X"BE",X"3E",
		X"32",X"C2",X"55",X"1B",X"3D",X"32",X"90",X"41",X"3E",X"11",X"CD",X"7A",X"09",X"06",X"B4",X"CD",
		X"72",X"03",X"CD",X"A1",X"03",X"C9",X"FF",X"0D",X"47",X"41",X"4D",X"45",X"20",X"4F",X"56",X"45",
		X"52",X"FF",X"FE",X"50",X"4C",X"41",X"59",X"45",X"52",X"FF",X"FF",X"FF",X"0E",X"47",X"45",X"54",
		X"20",X"52",X"45",X"41",X"44",X"59",X"FF",X"FE",X"50",X"4C",X"41",X"59",X"45",X"52",X"FF",X"FF",
		X"2A",X"12",X"4C",X"4E",X"23",X"46",X"23",X"E5",X"2A",X"10",X"4C",X"09",X"22",X"10",X"4C",X"C1",
		X"ED",X"43",X"12",X"4C",X"78",X"FE",X"0F",X"C2",X"F0",X"20",X"79",X"FE",X"D8",X"C2",X"F0",X"20",
		X"11",X"B9",X"A8",X"19",X"7C",X"E6",X"3F",X"67",X"CD",X"92",X"19",X"CD",X"F0",X"20",X"D1",X"E9",
		X"13",X"1A",X"E5",X"26",X"00",X"6F",X"E6",X"80",X"28",X"01",X"25",X"19",X"EB",X"E1",X"C3",X"5D",
		X"1C",X"E5",X"23",X"23",X"36",X"00",X"E1",X"C9",X"3A",X"2C",X"4F",X"21",X"00",X"40",X"0E",X"21",
		X"F3",X"ED",X"A2",X"5F",X"07",X"83",X"07",X"83",X"07",X"16",X"00",X"5F",X"0D",X"ED",X"AA",X"FB",
		X"21",X"D8",X"4E",X"19",X"11",X"0B",X"00",X"19",X"7E",X"2B",X"A7",X"20",X"5D",X"3A",X"2C",X"4F",
		X"A7",X"28",X"57",X"E5",X"11",X"FB",X"FF",X"19",X"46",X"23",X"4E",X"23",X"23",X"36",X"00",X"CD",
		X"F9",X"20",X"E1",X"3A",X"35",X"4F",X"A7",X"C0",X"23",X"23",X"35",X"C0",X"3E",X"13",X"CD",X"7A",
		X"09",X"3A",X"29",X"4E",X"77",X"2B",X"36",X"A0",X"2B",X"E5",X"11",X"FA",X"FF",X"19",X"97",X"77",
		X"2B",X"77",X"2B",X"2B",X"E5",X"CD",X"99",X"21",X"E1",X"E5",X"23",X"23",X"23",X"23",X"70",X"23",
		X"71",X"E1",X"2B",X"7E",X"3D",X"07",X"07",X"16",X"00",X"5F",X"21",X"4A",X"2B",X"19",X"5E",X"23",
		X"56",X"E1",X"72",X"2B",X"73",X"1B",X"3E",X"FD",X"18",X"04",X"56",X"2B",X"5E",X"1A",X"FE",X"FF",
		X"CA",X"D1",X"1B",X"FE",X"FE",X"CA",X"C0",X"1B",X"FE",X"FD",X"E5",X"13",X"1A",X"28",X"0A",X"1B",
		X"23",X"23",X"7E",X"FE",X"C0",X"C2",X"E5",X"1C",X"1A",X"E1",X"2B",X"77",X"01",X"FB",X"FF",X"09",
		X"13",X"1A",X"86",X"FE",X"10",X"28",X"33",X"CB",X"7F",X"20",X"3B",X"77",X"23",X"13",X"1A",X"86",
		X"FE",X"0A",X"28",X"40",X"FE",X"FF",X"28",X"44",X"77",X"23",X"13",X"1A",X"86",X"77",X"23",X"13",
		X"1A",X"86",X"77",X"13",X"2B",X"1A",X"86",X"47",X"13",X"23",X"1A",X"86",X"4F",X"13",X"23",X"23",
		X"E5",X"23",X"73",X"23",X"72",X"E1",X"CD",X"F9",X"20",X"C9",X"2B",X"2B",X"7E",X"3C",X"E6",X"0F",
		X"77",X"23",X"23",X"97",X"18",X"C5",X"2B",X"2B",X"7E",X"3D",X"E6",X"0F",X"77",X"23",X"23",X"1A",
		X"C6",X"10",X"18",X"B7",X"2B",X"2B",X"34",X"23",X"23",X"97",X"18",X"BC",X"2B",X"2B",X"35",X"23",
		X"23",X"3E",X"09",X"18",X"B3",X"D5",X"E5",X"7E",X"32",X"2E",X"4F",X"3A",X"14",X"4C",X"FE",X"01",
		X"20",X"09",X"CD",X"3D",X"3C",X"3A",X"30",X"4C",X"4F",X"18",X"43",X"3A",X"2C",X"4F",X"A7",X"20",
		X"3B",X"CD",X"74",X"01",X"3A",X"0D",X"4C",X"4F",X"3E",X"FF",X"32",X"0D",X"4C",X"79",X"2F",X"0E",
		X"80",X"CB",X"77",X"28",X"04",X"CB",X"E1",X"18",X"25",X"CB",X"6F",X"28",X"04",X"CB",X"D9",X"18",
		X"1D",X"E6",X"0F",X"28",X"19",X"CB",X"D1",X"47",X"E6",X"06",X"28",X"06",X"CB",X"57",X"28",X"0E",
		X"18",X"06",X"CB",X"C9",X"CB",X"40",X"28",X"06",X"CB",X"C1",X"18",X"02",X"0E",X"80",X"E1",X"E5",
		X"3A",X"2C",X"4F",X"A7",X"28",X"73",X"11",X"FA",X"FF",X"19",X"5E",X"23",X"56",X"06",X"0B",X"CD",
		X"B4",X"1F",X"A7",X"28",X"64",X"06",X"0B",X"CD",X"AE",X"1F",X"A7",X"28",X"5C",X"23",X"23",X"23",
		X"23",X"23",X"06",X"05",X"CD",X"B4",X"1F",X"A7",X"28",X"28",X"06",X"05",X"CD",X"AE",X"1F",X"A7",
		X"28",X"20",X"3A",X"E3",X"4E",X"CB",X"67",X"20",X"1C",X"E6",X"86",X"FE",X"86",X"28",X"13",X"7E",
		X"A7",X"28",X"0F",X"FE",X"A0",X"28",X"0B",X"FE",X"C0",X"28",X"07",X"3E",X"01",X"32",X"A5",X"4E",
		X"18",X"27",X"3A",X"E3",X"4E",X"FE",X"99",X"20",X"20",X"7E",X"A7",X"28",X"1C",X"FE",X"C0",X"28",
		X"18",X"E6",X"86",X"FE",X"86",X"28",X"12",X"0E",X"C0",X"11",X"F5",X"FF",X"19",X"7E",X"CD",X"23",
		X"05",X"3E",X"0E",X"CD",X"7A",X"09",X"C3",X"74",X"1F",X"E1",X"E5",X"11",X"F8",X"FF",X"19",X"7E",
		X"A7",X"28",X"06",X"E1",X"D1",X"1A",X"C3",X"79",X"1C",X"23",X"7E",X"A7",X"28",X"28",X"79",X"E6",
		X"86",X"FE",X"86",X"3A",X"2E",X"4F",X"20",X"01",X"79",X"E6",X"87",X"F6",X"86",X"4F",X"06",X"04",
		X"E6",X"01",X"20",X"02",X"06",X"FC",X"11",X"07",X"00",X"19",X"CD",X"0F",X"22",X"3A",X"2E",X"4F",
		X"B9",X"28",X"D0",X"C3",X"74",X"1F",X"CD",X"12",X"21",X"3A",X"2C",X"4F",X"A7",X"28",X"15",X"E5",
		X"11",X"07",X"00",X"19",X"CB",X"71",X"20",X"04",X"CB",X"76",X"28",X"04",X"E1",X"C3",X"74",X"1F",
		X"CD",X"C4",X"1F",X"E1",X"2B",X"2B",X"CD",X"DF",X"21",X"22",X"30",X"4F",X"3A",X"2C",X"4F",X"A7",
		X"20",X"32",X"CB",X"6E",X"28",X"2E",X"CB",X"AE",X"E1",X"E5",X"11",X"F6",X"FF",X"19",X"CD",X"B3",
		X"21",X"97",X"77",X"2B",X"77",X"11",X"E0",X"FF",X"19",X"77",X"23",X"77",X"3E",X"06",X"CD",X"23",
		X"05",X"3E",X"0F",X"CD",X"7A",X"09",X"21",X"8B",X"4E",X"35",X"20",X"08",X"3E",X"01",X"32",X"A4",
		X"4E",X"C3",X"C3",X"1D",X"79",X"FE",X"90",X"CA",X"74",X"1F",X"3A",X"2E",X"4F",X"FE",X"90",X"79",
		X"20",X"05",X"0E",X"99",X"C3",X"74",X"1F",X"FE",X"88",X"C2",X"EF",X"1E",X"2A",X"30",X"4F",X"CB",
		X"66",X"CA",X"74",X"1F",X"2B",X"CB",X"76",X"C2",X"74",X"1F",X"23",X"23",X"CB",X"76",X"C2",X"74",
		X"1F",X"E1",X"E5",X"11",X"FB",X"FF",X"19",X"46",X"11",X"FC",X"FF",X"19",X"7E",X"F5",X"2B",X"7E",
		X"22",X"3A",X"4F",X"C5",X"CD",X"F0",X"21",X"3A",X"32",X"4F",X"A1",X"20",X"05",X"C1",X"F1",X"C3",
		X"74",X"1F",X"C1",X"F1",X"23",X"E5",X"96",X"3E",X"04",X"F2",X"AE",X"1E",X"ED",X"44",X"11",X"F8",
		X"FF",X"19",X"5F",X"7E",X"A7",X"28",X"04",X"E1",X"C3",X"74",X"1F",X"3E",X"04",X"CD",X"7A",X"09",
		X"36",X"01",X"23",X"23",X"73",X"23",X"70",X"2A",X"3A",X"4F",X"CD",X"B3",X"21",X"2B",X"2B",X"11",
		X"00",X"04",X"19",X"EB",X"E1",X"E5",X"23",X"23",X"73",X"23",X"72",X"3A",X"62",X"4D",X"D6",X"02",
		X"12",X"21",X"E0",X"FF",X"19",X"77",X"E1",X"CD",X"DF",X"21",X"CB",X"B6",X"C3",X"74",X"1F",X"E6",
		X"86",X"FE",X"86",X"20",X"5F",X"2A",X"30",X"4F",X"CB",X"76",X"20",X"09",X"3A",X"2E",X"4F",X"E6",
		X"86",X"FE",X"86",X"20",X"36",X"3A",X"2C",X"4F",X"CB",X"41",X"28",X"08",X"CB",X"5E",X"28",X"11",
		X"06",X"04",X"18",X"06",X"CB",X"56",X"28",X"16",X"06",X"FC",X"E1",X"E5",X"CD",X"0F",X"22",X"18",
		X"53",X"A7",X"28",X"4E",X"CB",X"56",X"28",X"19",X"79",X"EE",X"01",X"4F",X"18",X"EA",X"A7",X"28",
		X"41",X"CB",X"5E",X"28",X"0C",X"79",X"EE",X"01",X"4F",X"18",X"D5",X"3A",X"2C",X"4F",X"A7",X"28",
		X"31",X"ED",X"5F",X"E6",X"3F",X"FE",X"20",X"38",X"29",X"E6",X"0F",X"FE",X"08",X"0E",X"84",X"38",
		X"1B",X"0C",X"18",X"08",X"FE",X"84",X"20",X"1A",X"CB",X"41",X"28",X"10",X"CB",X"4E",X"28",X"14",
		X"3A",X"2C",X"4F",X"A7",X"28",X"0C",X"79",X"EE",X"01",X"4F",X"18",X"08",X"CB",X"46",X"28",X"04",
		X"18",X"EE",X"0E",X"80",X"E1",X"3A",X"2E",X"4F",X"B9",X"D1",X"1A",X"CA",X"79",X"1C",X"71",X"CD",
		X"40",X"22",X"E5",X"11",X"F5",X"FF",X"19",X"7E",X"07",X"16",X"00",X"5F",X"21",X"9A",X"22",X"19",
		X"5E",X"23",X"56",X"79",X"CD",X"6C",X"22",X"07",X"26",X"00",X"6F",X"19",X"5E",X"23",X"56",X"CD",
		X"92",X"22",X"E1",X"2B",X"72",X"2B",X"73",X"E1",X"1B",X"3E",X"FD",X"C3",X"5E",X"1C",X"3A",X"DE",
		X"4E",X"92",X"18",X"04",X"3A",X"DD",X"4E",X"93",X"CB",X"7F",X"28",X"02",X"ED",X"44",X"B8",X"3E",
		X"00",X"D0",X"3C",X"C9",X"3A",X"14",X"4C",X"A7",X"C0",X"4E",X"23",X"23",X"35",X"C0",X"3A",X"2A",
		X"4E",X"5F",X"ED",X"5F",X"E6",X"3F",X"FE",X"10",X"30",X"01",X"1C",X"73",X"11",X"F3",X"FF",X"19",
		X"7E",X"11",X"0B",X"00",X"19",X"FE",X"01",X"28",X"12",X"FE",X"02",X"28",X"17",X"FE",X"03",X"28",
		X"23",X"FE",X"04",X"28",X"48",X"FE",X"05",X"28",X"3C",X"18",X"FE",X"0E",X"84",X"ED",X"5F",X"E6",
		X"01",X"B1",X"4F",X"C9",X"0E",X"84",X"ED",X"5F",X"E6",X"11",X"20",X"03",X"0E",X"88",X"C9",X"E6",
		X"01",X"B1",X"4F",X"C9",X"7E",X"4F",X"E6",X"86",X"FE",X"86",X"20",X"10",X"11",X"F9",X"FF",X"19",
		X"7E",X"A7",X"C0",X"ED",X"5F",X"E6",X"02",X"C0",X"0E",X"84",X"18",X"02",X"0E",X"86",X"ED",X"5F",
		X"E6",X"01",X"B1",X"4F",X"C9",X"01",X"06",X"0E",X"11",X"0A",X"20",X"18",X"06",X"01",X"02",X"04",
		X"11",X"0B",X"30",X"ED",X"43",X"36",X"4F",X"ED",X"53",X"38",X"4F",X"11",X"F7",X"FF",X"19",X"E5",
		X"CD",X"DF",X"21",X"CB",X"76",X"E1",X"23",X"23",X"23",X"20",X"54",X"ED",X"5F",X"E6",X"06",X"28",
		X"0D",X"ED",X"5F",X"E6",X"3F",X"FE",X"10",X"0E",X"86",X"DA",X"2E",X"20",X"18",X"04",X"0E",X"88",
		X"C9",X"2B",X"3A",X"DD",X"4E",X"96",X"06",X"01",X"38",X"03",X"05",X"ED",X"44",X"4F",X"3A",X"39",
		X"4F",X"B9",X"38",X"26",X"ED",X"5F",X"47",X"11",X"06",X"00",X"19",X"7E",X"CB",X"57",X"20",X"05",
		X"0E",X"84",X"C3",X"2E",X"20",X"E6",X"01",X"4F",X"3A",X"38",X"4F",X"A0",X"20",X"07",X"3E",X"84",
		X"B1",X"EE",X"01",X"4F",X"C9",X"3E",X"84",X"B1",X"4F",X"C9",X"3E",X"84",X"B0",X"4F",X"C9",X"23",
		X"ED",X"5F",X"47",X"3A",X"36",X"4F",X"A0",X"28",X"B8",X"46",X"11",X"05",X"00",X"19",X"7E",X"E6",
		X"86",X"FE",X"86",X"20",X"1D",X"E5",X"11",X"F9",X"FF",X"19",X"7E",X"E1",X"A7",X"4E",X"C0",X"3A",
		X"DE",X"4E",X"90",X"28",X"08",X"ED",X"5F",X"47",X"3A",X"37",X"4F",X"A0",X"C0",X"0E",X"84",X"C3",
		X"2E",X"20",X"3A",X"DE",X"4E",X"90",X"06",X"01",X"30",X"01",X"05",X"3E",X"86",X"B0",X"4F",X"C9",
		X"ED",X"5F",X"E6",X"03",X"3C",X"32",X"0B",X"4C",X"C9",X"E5",X"3A",X"2D",X"4F",X"07",X"07",X"5F",
		X"16",X"00",X"21",X"8C",X"4E",X"19",X"D1",X"1A",X"77",X"23",X"1B",X"1A",X"77",X"23",X"70",X"23",
		X"71",X"C9",X"E5",X"11",X"07",X"00",X"19",X"7E",X"CB",X"67",X"20",X"7B",X"A7",X"28",X"78",X"FE",
		X"C0",X"28",X"74",X"E6",X"86",X"FE",X"86",X"28",X"6E",X"3A",X"2C",X"4F",X"A7",X"20",X"07",X"7E",
		X"E6",X"84",X"FE",X"84",X"28",X"61",X"C5",X"11",X"F6",X"FF",X"19",X"4E",X"23",X"46",X"23",X"23",
		X"E5",X"C5",X"06",X"04",X"21",X"AD",X"4E",X"11",X"0C",X"00",X"7E",X"B9",X"28",X"05",X"19",X"10",
		X"F9",X"18",X"41",X"23",X"C1",X"7E",X"23",X"90",X"0E",X"10",X"28",X"32",X"FE",X"FF",X"0E",X"0C",
		X"20",X"33",X"7E",X"B9",X"38",X"2F",X"11",X"F7",X"FF",X"19",X"7E",X"E1",X"A7",X"28",X"27",X"3A",
		X"2C",X"4F",X"A7",X"28",X"12",X"C1",X"0E",X"C0",X"2B",X"2B",X"2B",X"2B",X"7E",X"CD",X"23",X"05",
		X"3E",X"0E",X"CD",X"7A",X"09",X"18",X"10",X"3E",X"01",X"32",X"A5",X"4E",X"18",X"08",X"7E",X"B9",
		X"30",X"03",X"18",X"D2",X"C1",X"E1",X"C1",X"E1",X"C9",X"7E",X"07",X"07",X"07",X"07",X"06",X"F6",
		X"90",X"ED",X"44",X"47",X"23",X"7E",X"3D",X"4F",X"07",X"07",X"81",X"07",X"07",X"07",X"0E",X"18",
		X"81",X"4F",X"C9",X"7E",X"3D",X"E5",X"26",X"00",X"6F",X"29",X"29",X"29",X"29",X"29",X"29",X"EB",
		X"21",X"00",X"00",X"AF",X"ED",X"52",X"EB",X"E1",X"23",X"7E",X"3D",X"47",X"07",X"07",X"80",X"ED",
		X"44",X"A7",X"28",X"06",X"83",X"5F",X"3E",X"FF",X"8A",X"57",X"21",X"9E",X"43",X"19",X"C9",X"3E",
		X"06",X"96",X"07",X"07",X"07",X"07",X"2B",X"86",X"16",X"00",X"5F",X"21",X"2B",X"4E",X"19",X"C9",
		X"21",X"AD",X"4E",X"11",X"0C",X"00",X"0E",X"08",X"F5",X"96",X"CB",X"7F",X"28",X"02",X"ED",X"44",
		X"A7",X"28",X"0A",X"FE",X"01",X"28",X"06",X"CB",X"39",X"19",X"F1",X"18",X"EB",X"F1",X"C9",X"11",
		X"F6",X"FF",X"19",X"C5",X"7E",X"CD",X"F0",X"21",X"79",X"2F",X"5F",X"3A",X"32",X"4F",X"A3",X"32",
		X"32",X"4F",X"23",X"E5",X"CD",X"DF",X"21",X"CB",X"B6",X"E1",X"11",X"F8",X"FF",X"19",X"36",X"02",
		X"23",X"7E",X"23",X"70",X"CD",X"8C",X"30",X"3A",X"34",X"4F",X"B1",X"32",X"34",X"4F",X"C1",X"C9",
		X"C5",X"E5",X"7E",X"E6",X"86",X"FE",X"86",X"28",X"20",X"3A",X"2E",X"4F",X"E6",X"86",X"FE",X"86",
		X"20",X"17",X"11",X"F6",X"FF",X"19",X"7E",X"CD",X"F0",X"21",X"11",X"F9",X"FF",X"19",X"36",X"00",
		X"11",X"08",X"00",X"19",X"CD",X"DF",X"21",X"CB",X"F6",X"E1",X"C1",X"C9",X"C5",X"06",X"09",X"CB",
		X"77",X"20",X"1C",X"05",X"CB",X"6F",X"20",X"17",X"05",X"FE",X"99",X"28",X"12",X"05",X"CB",X"67",
		X"20",X"0D",X"05",X"CB",X"5F",X"20",X"08",X"05",X"CB",X"57",X"28",X"03",X"E6",X"03",X"47",X"78",
		X"C1",X"C9",X"3E",X"FF",X"BA",X"C0",X"18",X"FE",X"FF",X"FF",X"A6",X"22",X"8E",X"23",X"65",X"24",
		X"3E",X"25",X"04",X"26",X"E1",X"26",X"B9",X"22",X"DE",X"22",X"03",X"23",X"0C",X"23",X"3C",X"23",
		X"4C",X"23",X"5C",X"23",X"15",X"23",X"7B",X"98",X"22",X"0E",X"FD",X"00",X"03",X"00",X"00",X"00",
		X"12",X"FD",X"00",X"03",X"00",X"00",X"00",X"16",X"FD",X"00",X"03",X"00",X"00",X"01",X"1A",X"FC",
		X"00",X"04",X"00",X"00",X"00",X"1E",X"FD",X"00",X"03",X"00",X"00",X"00",X"FE",X"DC",X"0C",X"03",
		X"00",X"FD",X"00",X"00",X"00",X"10",X"03",X"00",X"FD",X"00",X"00",X"00",X"14",X"03",X"00",X"FD",
		X"00",X"00",X"01",X"18",X"04",X"00",X"FC",X"00",X"00",X"00",X"1C",X"03",X"00",X"FD",X"00",X"00",
		X"00",X"FE",X"DC",X"04",X"00",X"FF",X"00",X"FC",X"00",X"00",X"FE",X"F8",X"04",X"00",X"01",X"00",
		X"04",X"00",X"00",X"FE",X"F8",X"24",X"00",X"00",X"00",X"00",X"00",X"16",X"FD",X"24",X"00",X"00",
		X"00",X"00",X"00",X"12",X"FD",X"24",X"00",X"00",X"00",X"00",X"00",X"0C",X"FD",X"24",X"00",X"00",
		X"00",X"00",X"00",X"06",X"FD",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"F1",X"20",X"00",X"00",X"00",
		X"00",X"00",X"02",X"22",X"00",X"00",X"00",X"00",X"00",X"02",X"FE",X"F1",X"24",X"00",X"00",X"00",
		X"00",X"00",X"08",X"FD",X"24",X"00",X"00",X"00",X"00",X"00",X"10",X"28",X"00",X"00",X"00",X"00",
		X"00",X"16",X"2A",X"00",X"00",X"00",X"00",X"00",X"16",X"FE",X"F1",X"04",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FE",X"F8",X"DB",X"65",X"E1",X"D1",X"C1",X"F1",X"FB",X"C3",X"C2",X"19",X"A2",X"23",
		X"DC",X"23",X"98",X"22",X"98",X"22",X"16",X"24",X"98",X"22",X"98",X"22",X"98",X"22",X"1F",X"24",
		X"48",X"24",X"36",X"FE",X"00",X"02",X"00",X"00",X"00",X"3A",X"FE",X"00",X"02",X"00",X"00",X"00",
		X"3E",X"FE",X"00",X"02",X"00",X"00",X"00",X"3A",X"FE",X"00",X"02",X"00",X"00",X"00",X"36",X"FE",
		X"00",X"02",X"00",X"00",X"00",X"3A",X"FE",X"00",X"02",X"00",X"00",X"00",X"3E",X"FE",X"00",X"02",
		X"00",X"00",X"00",X"3A",X"FE",X"00",X"02",X"00",X"00",X"00",X"FE",X"C7",X"34",X"02",X"00",X"FE",
		X"00",X"00",X"00",X"38",X"02",X"00",X"FE",X"00",X"00",X"00",X"3C",X"02",X"00",X"FE",X"00",X"00",
		X"00",X"38",X"02",X"00",X"FE",X"00",X"00",X"00",X"34",X"02",X"00",X"FE",X"00",X"00",X"00",X"38",
		X"02",X"00",X"FE",X"00",X"00",X"00",X"3C",X"02",X"00",X"FE",X"00",X"00",X"00",X"38",X"02",X"00",
		X"FE",X"00",X"00",X"00",X"FE",X"C7",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"F8",X"2C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FD",X"2E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FD",X"2C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"D8",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"79",X"24",X"A5",X"24",X"98",X"22",X"98",X"22",X"D1",X"24",X"27",
		X"25",X"98",X"22",X"98",X"22",X"E1",X"24",X"0A",X"25",X"52",X"FE",X"00",X"02",X"00",X"00",X"00",
		X"4A",X"FD",X"00",X"03",X"00",X"00",X"00",X"4E",X"FD",X"00",X"03",X"00",X"00",X"00",X"56",X"FE",
		X"00",X"02",X"00",X"00",X"00",X"4E",X"FD",X"00",X"03",X"00",X"00",X"00",X"4A",X"FD",X"00",X"03",
		X"00",X"00",X"00",X"FE",X"D5",X"50",X"02",X"00",X"FE",X"00",X"00",X"01",X"48",X"03",X"00",X"FD",
		X"00",X"00",X"00",X"4C",X"03",X"00",X"FD",X"00",X"00",X"00",X"54",X"02",X"00",X"FE",X"00",X"00",
		X"00",X"4C",X"03",X"00",X"FD",X"00",X"00",X"00",X"48",X"03",X"00",X"FD",X"00",X"00",X"00",X"FE",
		X"D5",X"48",X"00",X"00",X"00",X"00",X"00",X"00",X"4C",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",
		X"F1",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"FD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FD",X"46",X"00",X"00",X"00",X"00",X"00",X"00",X"FD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FD",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"D8",X"5C",X"00",X"00",X"00",X"00",X"00",
		X"00",X"5C",X"00",X"00",X"00",X"00",X"00",X"00",X"5C",X"00",X"00",X"00",X"00",X"00",X"00",X"5C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"58",X"00",X"00",X"00",X"00",X"00",X"02",X"58",X"00",
		X"00",X"00",X"00",X"00",X"04",X"58",X"00",X"00",X"00",X"00",X"00",X"02",X"FE",X"EA",X"52",X"25",
		X"77",X"25",X"F2",X"25",X"FB",X"25",X"9C",X"25",X"98",X"22",X"98",X"22",X"98",X"22",X"AC",X"25",
		X"D5",X"25",X"6E",X"FD",X"00",X"03",X"00",X"00",X"00",X"72",X"FD",X"00",X"03",X"00",X"00",X"00",
		X"76",X"FC",X"00",X"04",X"00",X"00",X"01",X"7A",X"FD",X"00",X"03",X"00",X"00",X"00",X"7E",X"FD",
		X"00",X"03",X"00",X"00",X"00",X"FE",X"DC",X"6C",X"03",X"00",X"FD",X"00",X"00",X"00",X"70",X"03",
		X"00",X"FD",X"00",X"00",X"00",X"74",X"04",X"00",X"FC",X"00",X"00",X"01",X"78",X"03",X"00",X"FD",
		X"00",X"00",X"00",X"7C",X"03",X"00",X"FD",X"00",X"00",X"00",X"FE",X"DC",X"64",X"00",X"00",X"00",
		X"00",X"00",X"00",X"68",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"F1",X"60",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FD",X"62",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FD",X"60",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"D8",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"64",X"00",X"FF",X"00",X"FC",X"00",X"00",X"FE",X"F8",X"64",X"00",X"01",X"00",X"04",
		X"00",X"00",X"FE",X"F8",X"18",X"26",X"3D",X"26",X"B8",X"26",X"C1",X"26",X"62",X"26",X"CA",X"26",
		X"98",X"22",X"98",X"22",X"72",X"26",X"9B",X"26",X"92",X"FD",X"00",X"03",X"00",X"00",X"00",X"96",
		X"FD",X"00",X"03",X"00",X"00",X"00",X"9A",X"FC",X"00",X"04",X"00",X"00",X"00",X"9E",X"FD",X"00",
		X"03",X"00",X"00",X"00",X"A2",X"FD",X"00",X"03",X"00",X"00",X"00",X"FE",X"DC",X"90",X"03",X"00",
		X"FD",X"00",X"00",X"00",X"94",X"03",X"00",X"FD",X"00",X"00",X"00",X"98",X"04",X"00",X"FC",X"00",
		X"00",X"00",X"9C",X"03",X"00",X"FD",X"00",X"00",X"00",X"A0",X"03",X"00",X"FD",X"00",X"00",X"00",
		X"FE",X"DC",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"8C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"F1",X"84",X"00",X"00",X"00",X"00",X"00",X"00",X"FD",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FD",X"86",X"00",X"00",X"00",X"00",X"00",X"00",X"FD",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FD",X"84",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"D8",X"A8",X"00",X"00",X"00",X"00",
		X"00",X"00",X"A8",X"00",X"00",X"00",X"00",X"00",X"00",X"A8",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A8",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"88",X"00",X"FF",X"00",X"FC",X"00",X"00",X"FE",
		X"F8",X"88",X"00",X"01",X"00",X"04",X"00",X"00",X"FE",X"F8",X"A4",X"00",X"00",X"00",X"00",X"00",
		X"02",X"A4",X"00",X"00",X"00",X"00",X"00",X"04",X"A4",X"00",X"00",X"00",X"00",X"00",X"02",X"FE",
		X"EA",X"F5",X"26",X"13",X"27",X"87",X"27",X"90",X"27",X"31",X"27",X"99",X"27",X"98",X"22",X"98",
		X"22",X"41",X"27",X"6A",X"27",X"BA",X"FC",X"00",X"04",X"00",X"00",X"00",X"BE",X"FC",X"00",X"04",
		X"00",X"00",X"00",X"C2",X"FC",X"00",X"04",X"00",X"00",X"00",X"BE",X"FC",X"00",X"04",X"00",X"00",
		X"00",X"FE",X"E3",X"B8",X"04",X"00",X"FC",X"00",X"00",X"00",X"BC",X"04",X"00",X"FC",X"00",X"00",
		X"00",X"C0",X"04",X"00",X"FC",X"00",X"00",X"00",X"BC",X"04",X"00",X"FC",X"00",X"00",X"00",X"FE",
		X"E3",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"B4",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",
		X"F1",X"AC",X"00",X"00",X"00",X"00",X"00",X"00",X"FD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FD",X"AE",X"00",X"00",X"00",X"00",X"00",X"00",X"FD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FD",X"AC",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"D8",X"C8",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C8",X"00",X"00",X"00",X"00",X"00",X"00",X"C8",X"00",X"00",X"00",X"00",X"00",X"00",X"C8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"B0",X"00",X"FF",X"00",X"FC",X"00",X"00",X"FE",X"F8",
		X"B0",X"00",X"01",X"00",X"04",X"00",X"00",X"FE",X"F8",X"C4",X"00",X"00",X"00",X"00",X"00",X"02",
		X"C4",X"00",X"00",X"00",X"00",X"00",X"03",X"C4",X"00",X"00",X"00",X"00",X"00",X"02",X"FE",X"EA",
		X"F5",X"C5",X"D5",X"E5",X"F3",X"11",X"5F",X"37",X"21",X"C3",X"27",X"01",X"03",X"06",X"DB",X"64",
		X"C3",X"29",X"37",X"97",X"CD",X"BD",X"02",X"CD",X"C7",X"02",X"06",X"1E",X"CD",X"72",X"03",X"21",
		X"2B",X"4E",X"06",X"AB",X"77",X"23",X"10",X"FC",X"3C",X"32",X"A3",X"4C",X"36",X"0B",X"23",X"36",
		X"55",X"3A",X"16",X"4C",X"A7",X"28",X"14",X"97",X"32",X"32",X"4C",X"3E",X"05",X"32",X"33",X"4C",
		X"21",X"7A",X"10",X"22",X"34",X"4C",X"21",X"DC",X"42",X"36",X"3C",X"3A",X"4B",X"4D",X"FE",X"01",
		X"01",X"3C",X"4C",X"11",X"9C",X"4C",X"21",X"4C",X"4D",X"28",X"09",X"01",X"3D",X"4C",X"11",X"9D",
		X"4C",X"21",X"4F",X"4D",X"1A",X"32",X"9E",X"4C",X"0A",X"32",X"3E",X"4C",X"7E",X"FE",X"19",X"20",
		X"11",X"3A",X"14",X"4C",X"A7",X"7E",X"20",X"0A",X"3A",X"9E",X"4C",X"3C",X"32",X"9E",X"4C",X"3E",
		X"01",X"77",X"11",X"BB",X"30",X"3D",X"07",X"26",X"00",X"6F",X"19",X"7E",X"23",X"66",X"6F",X"CD",
		X"56",X"2E",X"32",X"62",X"4D",X"CD",X"5C",X"2B",X"97",X"32",X"DC",X"46",X"23",X"CD",X"56",X"2E",
		X"32",X"61",X"4D",X"23",X"CD",X"56",X"2E",X"32",X"5F",X"4D",X"23",X"CD",X"56",X"2E",X"32",X"60",
		X"4D",X"23",X"F3",X"DB",X"37",X"3E",X"72",X"00",X"47",X"DB",X"4D",X"3E",X"66",X"00",X"90",X"ED",
		X"44",X"0F",X"47",X"DB",X"32",X"DB",X"46",X"FB",X"11",X"01",X"00",X"78",X"32",X"56",X"4D",X"CD",
		X"56",X"2E",X"23",X"E5",X"D5",X"C5",X"07",X"DC",X"DE",X"2B",X"07",X"DC",X"E3",X"2B",X"21",X"1E",
		X"2C",X"22",X"52",X"4D",X"21",X"12",X"2C",X"06",X"06",X"E5",X"07",X"30",X"0E",X"F5",X"C5",X"D5",
		X"4E",X"23",X"46",X"EB",X"09",X"CD",X"F2",X"2B",X"D1",X"C1",X"F1",X"2A",X"52",X"4D",X"23",X"22",
		X"52",X"4D",X"E1",X"23",X"23",X"10",X"E2",X"C1",X"D1",X"21",X"05",X"00",X"19",X"EB",X"E1",X"10",
		X"BA",X"06",X"06",X"78",X"32",X"56",X"4D",X"3E",X"06",X"90",X"5F",X"07",X"07",X"83",X"16",X"00",
		X"5F",X"ED",X"53",X"57",X"4D",X"C5",X"CD",X"56",X"2E",X"23",X"E5",X"CD",X"3D",X"2C",X"21",X"DE",
		X"2C",X"22",X"52",X"4D",X"21",X"C4",X"2C",X"06",X"05",X"CD",X"8F",X"2C",X"D1",X"EB",X"CD",X"56",
		X"2E",X"EB",X"13",X"D5",X"06",X"08",X"CD",X"8F",X"2C",X"E1",X"C1",X"10",X"C6",X"3E",X"06",X"47",
		X"32",X"5A",X"4D",X"3E",X"E0",X"32",X"5C",X"4D",X"11",X"E6",X"4E",X"ED",X"53",X"5D",X"4D",X"78",
		X"32",X"56",X"4D",X"3E",X"01",X"32",X"59",X"4D",X"3E",X"E6",X"32",X"5B",X"4D",X"C5",X"CD",X"56",
		X"2E",X"23",X"E5",X"CD",X"38",X"2C",X"06",X"05",X"CD",X"EB",X"2C",X"D1",X"EB",X"CD",X"56",X"2E",
		X"EB",X"13",X"D5",X"06",X"08",X"CD",X"EB",X"2C",X"3A",X"5A",X"4D",X"3D",X"32",X"5A",X"4D",X"3A",
		X"5C",X"4D",X"D6",X"28",X"32",X"5C",X"4D",X"E1",X"C1",X"10",X"C4",X"06",X"06",X"78",X"32",X"56",
		X"4D",X"3E",X"06",X"90",X"5F",X"07",X"07",X"83",X"16",X"00",X"5F",X"ED",X"53",X"57",X"4D",X"C5",
		X"CD",X"56",X"2E",X"23",X"E5",X"21",X"59",X"2D",X"22",X"52",X"4D",X"21",X"49",X"2D",X"06",X"08",
		X"CD",X"29",X"2D",X"E1",X"C1",X"10",X"D6",X"01",X"FC",X"2D",X"ED",X"43",X"52",X"4D",X"01",X"F4",
		X"2D",X"ED",X"43",X"54",X"4D",X"CD",X"56",X"2E",X"32",X"32",X"4F",X"32",X"33",X"4F",X"07",X"07",
		X"07",X"07",X"23",X"06",X"04",X"11",X"A6",X"4E",X"C5",X"D5",X"07",X"30",X"7E",X"F5",X"CD",X"56",
		X"2E",X"47",X"23",X"CD",X"56",X"2E",X"23",X"32",X"56",X"4D",X"E5",X"90",X"21",X"56",X"4D",X"CD",
		X"B6",X"2D",X"CD",X"38",X"2E",X"CB",X"D6",X"47",X"21",X"56",X"4D",X"35",X"CD",X"B6",X"2D",X"CD",
		X"38",X"2E",X"CB",X"D6",X"CB",X"DE",X"10",X"F0",X"CB",X"96",X"E1",X"97",X"12",X"13",X"CD",X"56",
		X"2E",X"23",X"32",X"56",X"4D",X"E5",X"47",X"07",X"07",X"80",X"47",X"D6",X"1E",X"ED",X"44",X"F5",
		X"78",X"07",X"07",X"07",X"C6",X"F0",X"12",X"13",X"97",X"12",X"13",X"12",X"13",X"12",X"13",X"ED",
		X"4B",X"54",X"4D",X"0A",X"6F",X"03",X"0A",X"67",X"F1",X"06",X"00",X"4F",X"09",X"7D",X"12",X"13",
		X"7C",X"12",X"13",X"ED",X"4B",X"52",X"4D",X"0A",X"12",X"13",X"3A",X"56",X"4D",X"12",X"13",X"97",
		X"12",X"CD",X"E5",X"2D",X"CD",X"38",X"2E",X"CB",X"F6",X"E1",X"F1",X"D1",X"E5",X"2A",X"54",X"4D",
		X"23",X"23",X"22",X"54",X"4D",X"2A",X"52",X"4D",X"23",X"22",X"52",X"4D",X"21",X"0C",X"00",X"19",
		X"EB",X"E1",X"C1",X"05",X"C2",X"98",X"29",X"CD",X"79",X"2B",X"21",X"D8",X"4E",X"97",X"77",X"23",
		X"36",X"01",X"23",X"36",X"01",X"23",X"77",X"23",X"77",X"23",X"36",X"E6",X"23",X"36",X"18",X"23",
		X"36",X"09",X"23",X"36",X"04",X"23",X"36",X"7B",X"23",X"36",X"23",X"23",X"36",X"A0",X"3A",X"4B",
		X"4D",X"FE",X"01",X"11",X"9C",X"4C",X"21",X"4E",X"4D",X"28",X"06",X"11",X"9D",X"4C",X"21",X"51",
		X"4D",X"3A",X"9E",X"4C",X"12",X"7E",X"FE",X"10",X"38",X"0A",X"3A",X"14",X"4C",X"A7",X"7E",X"20",
		X"03",X"3E",X"0F",X"77",X"11",X"E4",X"35",X"3D",X"07",X"26",X"00",X"6F",X"19",X"7E",X"23",X"66",
		X"6F",X"3A",X"9E",X"4C",X"A7",X"7E",X"28",X"01",X"97",X"01",X"25",X"4E",X"02",X"23",X"7E",X"03",
		X"02",X"03",X"02",X"23",X"7E",X"03",X"02",X"23",X"7E",X"03",X"02",X"23",X"7E",X"03",X"02",X"11",
		X"E6",X"4E",X"C3",X"6A",X"2E",X"3A",X"01",X"4C",X"47",X"23",X"7E",X"12",X"23",X"4E",X"C5",X"E5",
		X"21",X"07",X"00",X"19",X"EB",X"3D",X"07",X"07",X"06",X"00",X"4F",X"21",X"48",X"2B",X"09",X"06",
		X"04",X"7E",X"12",X"23",X"13",X"10",X"FA",X"97",X"12",X"13",X"E1",X"C1",X"79",X"12",X"13",X"3A",
		X"2A",X"4E",X"12",X"13",X"10",X"D3",X"3A",X"9E",X"4C",X"A7",X"28",X"06",X"21",X"27",X"4E",X"35",
		X"23",X"35",X"3A",X"14",X"4C",X"A7",X"20",X"3E",X"97",X"32",X"A3",X"4C",X"3E",X"0B",X"CD",X"0E",
		X"05",X"CD",X"95",X"05",X"CD",X"C4",X"05",X"3A",X"37",X"4C",X"FE",X"02",X"20",X"0B",X"3E",X"0B",
		X"CD",X"16",X"05",X"CD",X"9E",X"05",X"CD",X"CC",X"05",X"3A",X"4B",X"4D",X"FE",X"01",X"3E",X"0E",
		X"32",X"02",X"4C",X"28",X"12",X"CD",X"CC",X"05",X"3A",X"AC",X"4C",X"A7",X"20",X"03",X"CD",X"6E",
		X"06",X"3E",X"01",X"32",X"A3",X"4C",X"C9",X"CD",X"C4",X"05",X"18",X"EC",X"DB",X"65",X"DB",X"64",
		X"E1",X"D1",X"C1",X"F1",X"FB",X"C3",X"B5",X"2A",X"05",X"0B",X"1F",X"24",X"12",X"11",X"E1",X"24",
		X"0A",X"18",X"AC",X"25",X"0C",X"21",X"72",X"26",X"0B",X"2B",X"41",X"27",X"E5",X"CD",X"1A",X"03",
		X"06",X"07",X"3E",X"08",X"11",X"E0",X"FF",X"21",X"81",X"43",X"C5",X"06",X"1A",X"CD",X"57",X"04",
		X"01",X"45",X"03",X"09",X"C1",X"10",X"F3",X"E1",X"C9",X"3E",X"20",X"11",X"01",X"00",X"06",X"1E",
		X"21",X"A1",X"43",X"CD",X"5C",X"04",X"06",X"1E",X"21",X"41",X"40",X"CD",X"5C",X"04",X"3E",X"25",
		X"11",X"E0",X"FF",X"06",X"1A",X"21",X"80",X"43",X"CD",X"57",X"04",X"3E",X"2D",X"06",X"1A",X"21",
		X"9F",X"43",X"CD",X"57",X"04",X"3A",X"A1",X"43",X"FE",X"28",X"3E",X"29",X"28",X"02",X"3E",X"24",
		X"32",X"A0",X"43",X"3A",X"41",X"40",X"FE",X"28",X"3E",X"5C",X"28",X"02",X"3E",X"26",X"32",X"40",
		X"40",X"3A",X"BE",X"43",X"FE",X"20",X"3E",X"5D",X"28",X"02",X"3E",X"2C",X"32",X"BF",X"43",X"3A",
		X"5E",X"40",X"FE",X"20",X"3E",X"5E",X"28",X"02",X"3E",X"2F",X"32",X"5F",X"40",X"C9",X"21",X"A0",
		X"43",X"18",X"03",X"21",X"40",X"40",X"D5",X"19",X"36",X"08",X"11",X"05",X"00",X"19",X"36",X"08",
		X"D1",X"C9",X"E5",X"11",X"01",X"00",X"06",X"05",X"3E",X"03",X"CD",X"5C",X"04",X"E1",X"01",X"E0",
		X"FF",X"09",X"06",X"05",X"3E",X"02",X"CD",X"5C",X"04",X"CD",X"38",X"2E",X"CB",X"CE",X"23",X"CB",
		X"C6",X"C9",X"A0",X"43",X"E0",X"42",X"20",X"42",X"E0",X"41",X"20",X"41",X"60",X"40",X"00",X"03",
		X"06",X"07",X"0A",X"0D",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"19",X"1D",
		X"1D",X"1D",X"1B",X"1A",X"1D",X"1D",X"1D",X"1C",X"11",X"2E",X"2C",X"18",X"03",X"11",X"24",X"2C",
		X"07",X"06",X"03",X"21",X"9E",X"43",X"DC",X"5C",X"2C",X"07",X"06",X"01",X"21",X"1E",X"42",X"DC",
		X"5C",X"2C",X"07",X"06",X"03",X"21",X"1E",X"41",X"DC",X"5C",X"2C",X"C9",X"F5",X"C5",X"3A",X"56",
		X"4D",X"3D",X"4F",X"07",X"07",X"81",X"ED",X"44",X"06",X"00",X"28",X"01",X"05",X"4F",X"09",X"C1",
		X"C5",X"D5",X"CD",X"86",X"2C",X"01",X"E5",X"FF",X"09",X"CD",X"86",X"2C",X"01",X"E5",X"FF",X"09",
		X"D1",X"C1",X"10",X"EC",X"F1",X"C9",X"06",X"05",X"1A",X"77",X"13",X"2B",X"10",X"FA",X"C9",X"C5",
		X"E5",X"07",X"30",X"22",X"F5",X"5E",X"23",X"56",X"3A",X"3E",X"4C",X"A7",X"20",X"0B",X"D5",X"E5",
		X"CD",X"29",X"2E",X"CB",X"6E",X"E1",X"D1",X"28",X"0C",X"CD",X"61",X"2D",X"CD",X"38",X"2E",X"CB",
		X"EE",X"21",X"8B",X"4E",X"34",X"F1",X"2A",X"52",X"4D",X"23",X"22",X"52",X"4D",X"E1",X"23",X"23",
		X"C1",X"10",X"CC",X"C9",X"85",X"43",X"45",X"43",X"05",X"43",X"C5",X"42",X"85",X"42",X"45",X"42",
		X"05",X"42",X"C5",X"41",X"85",X"41",X"45",X"41",X"05",X"41",X"C5",X"40",X"85",X"40",X"01",X"02",
		X"03",X"04",X"05",X"06",X"07",X"08",X"09",X"0A",X"0B",X"0C",X"0D",X"C5",X"07",X"30",X"21",X"F5",
		X"2A",X"5D",X"4D",X"23",X"ED",X"5B",X"59",X"4D",X"73",X"23",X"72",X"23",X"97",X"77",X"23",X"77",
		X"23",X"ED",X"5B",X"5B",X"4D",X"73",X"23",X"72",X"11",X"08",X"00",X"19",X"22",X"5D",X"4D",X"F1",
		X"CD",X"17",X"2D",X"C1",X"10",X"D5",X"C9",X"F5",X"3A",X"59",X"4D",X"3C",X"32",X"59",X"4D",X"3A",
		X"5B",X"4D",X"C6",X"F0",X"32",X"5B",X"4D",X"F1",X"C9",X"C5",X"E5",X"07",X"30",X"0D",X"F5",X"5E",
		X"23",X"56",X"CD",X"95",X"2D",X"CD",X"38",X"2E",X"CB",X"E6",X"F1",X"2A",X"52",X"4D",X"23",X"22",
		X"52",X"4D",X"E1",X"23",X"23",X"C1",X"10",X"E1",X"C9",X"85",X"43",X"05",X"43",X"C5",X"42",X"45",
		X"42",X"C5",X"41",X"45",X"41",X"05",X"41",X"85",X"40",X"01",X"03",X"04",X"06",X"08",X"0A",X"0B",
		X"0D",X"2A",X"57",X"4D",X"19",X"3A",X"61",X"4D",X"77",X"2B",X"3C",X"77",X"11",X"E0",X"FF",X"19",
		X"3C",X"77",X"23",X"3C",X"77",X"11",X"20",X"04",X"19",X"3A",X"9E",X"4C",X"A7",X"3A",X"60",X"4D",
		X"47",X"3A",X"5F",X"4D",X"4F",X"28",X"03",X"01",X"00",X"00",X"70",X"2B",X"71",X"11",X"E0",X"FF",
		X"19",X"71",X"23",X"70",X"C9",X"2A",X"57",X"4D",X"19",X"2B",X"2B",X"7E",X"C6",X"10",X"77",X"11",
		X"E0",X"FF",X"19",X"7E",X"C6",X"11",X"77",X"11",X"00",X"04",X"19",X"3A",X"62",X"4D",X"3D",X"77",
		X"11",X"20",X"00",X"19",X"77",X"C9",X"F5",X"C5",X"D5",X"7E",X"4F",X"07",X"07",X"81",X"D6",X"1E",
		X"ED",X"44",X"06",X"00",X"4F",X"2A",X"54",X"4D",X"7E",X"23",X"66",X"6F",X"09",X"06",X"05",X"3E",
		X"04",X"86",X"77",X"11",X"E0",X"FF",X"19",X"3E",X"05",X"86",X"77",X"11",X"1F",X"00",X"19",X"10",
		X"EE",X"D1",X"C1",X"F1",X"C9",X"F5",X"C5",X"D5",X"E5",X"11",X"FB",X"01",X"CD",X"44",X"01",X"E1",
		X"D1",X"C1",X"F1",X"C9",X"45",X"43",X"85",X"42",X"85",X"41",X"C5",X"40",X"02",X"05",X"09",X"0C",
		X"D5",X"97",X"57",X"5A",X"7E",X"23",X"E5",X"6F",X"26",X"00",X"19",X"EB",X"E1",X"10",X"F5",X"3E",
		X"05",X"32",X"01",X"4C",X"32",X"C0",X"50",X"0D",X"20",X"EA",X"D1",X"19",X"CB",X"24",X"CB",X"24",
		X"CB",X"3C",X"CB",X"3C",X"E5",X"DD",X"E1",X"DD",X"E9",X"21",X"65",X"4D",X"3A",X"4B",X"4D",X"FE",
		X"01",X"28",X"08",X"21",X"C5",X"4D",X"18",X"03",X"21",X"2B",X"4E",X"F5",X"C5",X"E5",X"2A",X"52",
		X"4D",X"46",X"3A",X"56",X"4D",X"D6",X"06",X"ED",X"44",X"07",X"07",X"07",X"07",X"80",X"06",X"00",
		X"4F",X"E1",X"09",X"C1",X"F1",X"C9",X"C5",X"D5",X"0E",X"51",X"F3",X"ED",X"50",X"ED",X"58",X"7E",
		X"0E",X"28",X"ED",X"50",X"ED",X"58",X"FB",X"D1",X"C1",X"C9",X"F5",X"C5",X"D5",X"E5",X"F3",X"21",
		X"7E",X"2E",X"11",X"9C",X"F5",X"01",X"08",X"22",X"DB",X"64",X"DB",X"65",X"18",X"82",X"3E",X"08",
		X"C3",X"32",X"2F",X"3A",X"2E",X"4F",X"FE",X"90",X"3E",X"07",X"C2",X"32",X"2F",X"3E",X"09",X"C3",
		X"32",X"2F",X"3A",X"E3",X"4E",X"FE",X"86",X"3A",X"2E",X"4F",X"28",X"0A",X"FE",X"87",X"CA",X"35",
		X"2F",X"3E",X"00",X"C3",X"32",X"2F",X"FE",X"86",X"CA",X"35",X"2F",X"3E",X"01",X"C3",X"32",X"2F",
		X"3A",X"25",X"4E",X"32",X"0E",X"4C",X"97",X"32",X"A7",X"4C",X"3C",X"32",X"3B",X"4C",X"06",X"1E",
		X"CD",X"72",X"03",X"3A",X"8B",X"4E",X"32",X"C0",X"50",X"A7",X"CA",X"A8",X"2F",X"3A",X"A5",X"4E",
		X"A7",X"C2",X"F0",X"2F",X"3E",X"15",X"CD",X"7A",X"09",X"3A",X"35",X"4F",X"3C",X"E6",X"03",X"32",
		X"35",X"4F",X"3A",X"16",X"4C",X"A7",X"28",X"03",X"CD",X"77",X"11",X"97",X"32",X"2D",X"4F",X"32",
		X"2C",X"4F",X"32",X"34",X"4F",X"3D",X"32",X"0D",X"4C",X"3E",X"0F",X"32",X"32",X"4F",X"CD",X"D8",
		X"1B",X"3A",X"2E",X"4F",X"E6",X"86",X"FE",X"86",X"20",X"0E",X"3A",X"E3",X"4E",X"E6",X"86",X"FE",
		X"86",X"28",X"05",X"3E",X"0A",X"CD",X"7A",X"09",X"3A",X"E3",X"4E",X"FE",X"99",X"CA",X"7E",X"2E",
		X"FE",X"90",X"CA",X"83",X"2E",X"E6",X"86",X"FE",X"86",X"CA",X"92",X"2E",X"FE",X"84",X"20",X"05",
		X"3E",X"10",X"CD",X"7A",X"09",X"3A",X"14",X"4C",X"A7",X"20",X"10",X"3A",X"E3",X"4E",X"CB",X"67",
		X"3A",X"28",X"4E",X"20",X"03",X"3A",X"27",X"4E",X"CD",X"B6",X"06",X"3E",X"01",X"06",X"05",X"F5",
		X"C5",X"32",X"2D",X"4F",X"32",X"2C",X"4F",X"CD",X"D8",X"1B",X"C1",X"F1",X"3C",X"10",X"F0",X"3A",
		X"33",X"4F",X"47",X"3A",X"32",X"4F",X"A0",X"06",X"04",X"0E",X"08",X"F5",X"C5",X"A1",X"C4",X"2D",
		X"30",X"C1",X"F1",X"CB",X"29",X"10",X"F4",X"3A",X"14",X"4C",X"A7",X"20",X"1A",X"97",X"32",X"A3",
		X"4C",X"3A",X"4B",X"4D",X"FE",X"01",X"3E",X"06",X"28",X"05",X"CD",X"16",X"05",X"18",X"03",X"CD",
		X"0E",X"05",X"3E",X"01",X"32",X"A3",X"4C",X"CD",X"A9",X"30",X"CD",X"A9",X"30",X"CD",X"8A",X"03",
		X"C3",X"C3",X"2E",X"CD",X"0E",X"05",X"18",X"20",X"97",X"32",X"3B",X"4C",X"CD",X"23",X"05",X"32",
		X"A3",X"4C",X"3C",X"32",X"A7",X"4C",X"3A",X"14",X"4C",X"A7",X"20",X"0C",X"3A",X"4B",X"4D",X"FE",
		X"01",X"3E",X"06",X"28",X"DE",X"CD",X"16",X"05",X"3E",X"01",X"32",X"A3",X"4C",X"CD",X"ED",X"06",
		X"3E",X"0D",X"CD",X"7A",X"09",X"CD",X"A1",X"03",X"97",X"32",X"A5",X"4E",X"3A",X"4B",X"4D",X"21",
		X"3C",X"4C",X"FE",X"01",X"28",X"03",X"21",X"3D",X"4C",X"36",X"01",X"97",X"32",X"A7",X"4C",X"C9",
		X"97",X"32",X"3B",X"4C",X"3C",X"32",X"A7",X"4C",X"CD",X"ED",X"06",X"3E",X"0C",X"CD",X"7A",X"09",
		X"CD",X"A1",X"03",X"3E",X"01",X"32",X"A5",X"4E",X"3A",X"4B",X"4D",X"21",X"3C",X"4C",X"11",X"65",
		X"4D",X"FE",X"01",X"28",X"06",X"21",X"3D",X"4C",X"11",X"C5",X"4D",X"36",X"00",X"21",X"2B",X"4E",
		X"06",X"60",X"7E",X"12",X"23",X"13",X"10",X"FA",X"97",X"32",X"A7",X"4C",X"C9",X"F5",X"3E",X"04",
		X"90",X"5F",X"07",X"83",X"07",X"07",X"16",X"00",X"5F",X"21",X"A6",X"4E",X"19",X"7E",X"A7",X"20",
		X"05",X"CD",X"82",X"30",X"F1",X"C9",X"FE",X"01",X"20",X"FE",X"23",X"7E",X"23",X"46",X"CD",X"8C",
		X"30",X"11",X"FA",X"FF",X"19",X"7E",X"2B",X"2B",X"BE",X"20",X"1E",X"2B",X"36",X"00",X"E5",X"CD",
		X"82",X"30",X"E1",X"11",X"0A",X"00",X"19",X"5E",X"23",X"56",X"3A",X"62",X"4D",X"3D",X"12",X"21",
		X"E0",X"FF",X"19",X"77",X"3E",X"02",X"CD",X"7A",X"09",X"C1",X"3A",X"34",X"4F",X"B0",X"32",X"34",
		X"4F",X"C9",X"11",X"08",X"00",X"19",X"CD",X"DF",X"21",X"CB",X"F6",X"C9",X"80",X"2B",X"77",X"11",
		X"08",X"00",X"19",X"7E",X"80",X"77",X"FE",X"FC",X"28",X"09",X"FE",X"28",X"C0",X"36",X"00",X"2B",
		X"34",X"23",X"C9",X"36",X"24",X"2B",X"35",X"23",X"C9",X"3A",X"25",X"4E",X"A7",X"C8",X"21",X"0E",
		X"4C",X"35",X"C0",X"3A",X"25",X"4E",X"77",X"CD",X"8A",X"03",X"C9",X"ED",X"30",X"22",X"31",X"57",
		X"31",X"86",X"31",X"B2",X"31",X"E1",X"31",X"16",X"32",X"4B",X"32",X"80",X"32",X"B5",X"32",X"E7",
		X"32",X"1C",X"33",X"51",X"33",X"86",X"33",X"BB",X"33",X"ED",X"33",X"22",X"34",X"57",X"34",X"8C",
		X"34",X"B8",X"34",X"E7",X"34",X"1C",X"35",X"48",X"35",X"7D",X"35",X"B2",X"35",X"0F",X"90",X"05",
		X"05",X"21",X"21",X"21",X"21",X"21",X"21",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",
		X"04",X"04",X"04",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"00",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"01",X"06",X"01",X"01",X"06",X"03",X"01",X"06",X"04",X"01",
		X"06",X"06",X"18",X"94",X"02",X"03",X"C0",X"C0",X"21",X"21",X"21",X"21",X"00",X"40",X"00",X"40",
		X"00",X"E0",X"01",X"50",X"02",X"48",X"04",X"44",X"00",X"08",X"02",X"00",X"00",X"00",X"00",X"20",
		X"01",X"00",X"00",X"08",X"18",X"18",X"19",X"80",X"01",X"80",X"0F",X"01",X"04",X"02",X"04",X"06",
		X"05",X"04",X"06",X"05",X"01",X"04",X"02",X"1B",X"98",X"01",X"01",X"C0",X"21",X"D2",X"D2",X"21",
		X"C0",X"1C",X"47",X"08",X"42",X"A0",X"40",X"A0",X"40",X"08",X"42",X"1C",X"47",X"00",X"80",X"00",
		X"20",X"00",X"80",X"00",X"20",X"00",X"80",X"00",X"00",X"04",X"04",X"20",X"20",X"04",X"04",X"06",
		X"01",X"06",X"06",X"01",X"06",X"06",X"15",X"9C",X"04",X"04",X"21",X"31",X"39",X"39",X"31",X"21",
		X"0F",X"F8",X"81",X"F0",X"00",X"20",X"00",X"20",X"81",X"F0",X"0F",X"F8",X"00",X"01",X"00",X"01",
		X"80",X"01",X"80",X"01",X"00",X"01",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"06",X"04",X"1E",X"A0",X"04",X"06",X"21",X"33",X"33",X"33",X"33",X"21",X"03",X"F8",X"00",X"00",
		X"40",X"00",X"40",X"00",X"00",X"00",X"03",X"F8",X"14",X"01",X"40",X"00",X"00",X"00",X"00",X"00",
		X"44",X"00",X"00",X"01",X"42",X"42",X"42",X"42",X"42",X"42",X"09",X"01",X"06",X"06",X"01",X"06",
		X"06",X"12",X"A4",X"06",X"06",X"2D",X"2D",X"C0",X"C0",X"2D",X"2D",X"47",X"1C",X"47",X"1C",X"00",
		X"E0",X"00",X"E0",X"47",X"1C",X"47",X"1C",X"08",X"00",X"00",X"02",X"00",X"10",X"01",X"01",X"00",
		X"00",X"00",X"00",X"81",X"81",X"C3",X"C3",X"81",X"81",X"0F",X"01",X"06",X"06",X"03",X"04",X"03",
		X"03",X"04",X"04",X"01",X"06",X"01",X"18",X"B4",X"04",X"0E",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"54",X"05",X"12",X"09",X"54",X"05",X"12",X"09",X"54",X"05",X"12",X"09",X"00",X"20",X"40",X"80",
		X"00",X"02",X"40",X"00",X"00",X"20",X"40",X"80",X"18",X"18",X"18",X"18",X"18",X"18",X"0F",X"01",
		X"06",X"02",X"01",X"06",X"05",X"01",X"06",X"05",X"01",X"06",X"02",X"1B",X"AC",X"06",X"06",X"21",
		X"21",X"C0",X"C0",X"C0",X"21",X"02",X"00",X"05",X"00",X"0F",X"A1",X"10",X"61",X"00",X"21",X"00",
		X"1E",X"00",X"00",X"00",X"10",X"01",X"00",X"08",X"02",X"00",X"10",X"00",X"00",X"02",X"02",X"06",
		X"24",X"60",X"40",X"0F",X"01",X"02",X"02",X"02",X"03",X"02",X"03",X"04",X"04",X"04",X"06",X"04",
		X"15",X"B0",X"04",X"04",X"21",X"D2",X"C6",X"C6",X"2B",X"21",X"01",X"F0",X"18",X"E1",X"14",X"81",
		X"17",X"81",X"03",X"20",X"01",X"F0",X"10",X"00",X"04",X"00",X"00",X"00",X"00",X"40",X"00",X"C0",
		X"00",X"00",X"01",X"37",X"37",X"C7",X"C7",X"01",X"0F",X"02",X"03",X"02",X"04",X"05",X"05",X"02",
		X"05",X"02",X"01",X"06",X"06",X"12",X"A8",X"07",X"07",X"C8",X"D0",X"21",X"21",X"21",X"21",X"14",
		X"15",X"08",X"AA",X"04",X"50",X"0A",X"A8",X"01",X"50",X"02",X"AA",X"00",X"40",X"04",X"00",X"00",
		X"20",X"00",X"20",X"00",X"20",X"00",X"00",X"10",X"20",X"01",X"01",X"81",X"80",X"0D",X"01",X"02",
		X"01",X"04",X"06",X"05",X"02",X"04",X"03",X"0F",X"B8",X"06",X"09",X"21",X"D0",X"21",X"21",X"C2",
		X"21",X"08",X"00",X"19",X"C0",X"0C",X"40",X"00",X"42",X"00",X"73",X"00",X"02",X"00",X"00",X"00",
		X"02",X"00",X"20",X"00",X"80",X"00",X"04",X"00",X"01",X"01",X"0C",X"31",X"8C",X"30",X"80",X"0F",
		X"01",X"03",X"02",X"02",X"04",X"03",X"03",X"05",X"04",X"04",X"06",X"05",X"1E",X"BC",X"1F",X"1C",
		X"C0",X"C2",X"C4",X"25",X"35",X"25",X"1F",X"E7",X"1F",X"E1",X"17",X"9C",X"07",X"9C",X"00",X"9C",
		X"00",X"9C",X"00",X"00",X"00",X"12",X"00",X"02",X"08",X"00",X"00",X"02",X"00",X"00",X"00",X"04",
		X"01",X"81",X"01",X"81",X"0F",X"01",X"04",X"04",X"01",X"02",X"01",X"05",X"06",X"06",X"01",X"05",
		X"01",X"0F",X"90",X"05",X"05",X"21",X"33",X"37",X"37",X"23",X"21",X"07",X"FC",X"00",X"E0",X"00",
		X"80",X"00",X"80",X"07",X"E0",X"0F",X"FC",X"00",X"10",X"00",X"10",X"00",X"00",X"00",X"40",X"08",
		X"00",X"00",X"10",X"82",X"69",X"96",X"69",X"86",X"01",X"0F",X"02",X"06",X"02",X"03",X"05",X"03",
		X"02",X"05",X"05",X"01",X"06",X"06",X"18",X"94",X"02",X"03",X"21",X"21",X"D0",X"CC",X"C2",X"21",
		X"02",X"AA",X"05",X"54",X"10",X"FF",X"1E",X"0F",X"1F",X"E1",X"05",X"54",X"00",X"01",X"10",X"00",
		X"02",X"00",X"40",X"20",X"00",X"04",X"00",X"00",X"80",X"00",X"60",X"18",X"06",X"01",X"0F",X"04",
		X"06",X"04",X"03",X"04",X"04",X"02",X"03",X"02",X"01",X"02",X"02",X"1B",X"98",X"01",X"01",X"62",
		X"72",X"72",X"31",X"31",X"21",X"21",X"80",X"21",X"C0",X"21",X"E0",X"01",X"F0",X"01",X"F8",X"01",
		X"FC",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"00",X"00",X"84",X"04",X"04",
		X"01",X"01",X"81",X"0B",X"01",X"06",X"06",X"04",X"06",X"04",X"01",X"03",X"03",X"15",X"9C",X"04",
		X"04",X"21",X"21",X"CC",X"CC",X"21",X"21",X"00",X"70",X"00",X"0E",X"5C",X"07",X"5C",X"07",X"0E",
		X"00",X"01",X"C0",X"00",X"04",X"00",X"80",X"00",X"20",X"00",X"80",X"00",X"20",X"00",X"00",X"80",
		X"B0",X"18",X"18",X"0D",X"01",X"0F",X"05",X"06",X"05",X"03",X"05",X"04",X"02",X"04",X"03",X"01",
		X"02",X"02",X"1E",X"A0",X"04",X"06",X"62",X"6A",X"62",X"70",X"62",X"62",X"0A",X"A1",X"03",X"01",
		X"07",X"E1",X"00",X"FD",X"00",X"51",X"05",X"51",X"00",X"00",X"00",X"12",X"08",X"00",X"01",X"00",
		X"00",X"02",X"00",X"00",X"06",X"C6",X"C6",X"E2",X"E2",X"C2",X"0F",X"01",X"05",X"05",X"02",X"03",
		X"03",X"04",X"06",X"06",X"01",X"06",X"06",X"12",X"A4",X"06",X"06",X"D2",X"D6",X"D6",X"D6",X"D6",
		X"25",X"10",X"E1",X"10",X"81",X"10",X"81",X"10",X"81",X"10",X"81",X"00",X"8C",X"00",X"40",X"00",
		X"04",X"04",X"00",X"00",X"04",X"00",X"40",X"00",X"00",X"64",X"60",X"60",X"60",X"60",X"29",X"0F",
		X"02",X"06",X"06",X"01",X"06",X"06",X"01",X"06",X"01",X"01",X"06",X"06",X"18",X"B4",X"04",X"0E",
		X"70",X"D8",X"CC",X"C6",X"83",X"21",X"81",X"EF",X"00",X"2F",X"00",X"0F",X"80",X"00",X"1F",X"E0",
		X"0F",X"EE",X"02",X"00",X"00",X"40",X"00",X"20",X"20",X"00",X"20",X"08",X"00",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"01",X"06",X"01",X"1B",X"AC",X"06",X"06",X"C0",X"23",X"25",X"29",
		X"31",X"C0",X"03",X"F0",X"03",X"F0",X"03",X"98",X"03",X"38",X"01",X"F8",X"09",X"F8",X"04",X"00",
		X"04",X"00",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"00",X"80",X"81",X"81",X"81",X"81",X"01",
		X"09",X"02",X"06",X"02",X"01",X"06",X"05",X"15",X"B0",X"04",X"04",X"21",X"21",X"62",X"6E",X"6E",
		X"2D",X"02",X"E8",X"02",X"E8",X"0E",X"E1",X"0E",X"01",X"0E",X"01",X"0E",X"0C",X"08",X"00",X"00",
		X"02",X"00",X"00",X"40",X"00",X"41",X"02",X"40",X"10",X"80",X"81",X"26",X"1A",X"1A",X"19",X"0F",
		X"05",X"06",X"05",X"01",X"04",X"01",X"01",X"04",X"01",X"01",X"05",X"01",X"12",X"A8",X"07",X"07",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"1F",X"EF",X"1F",X"EF",X"1F",X"EF",X"1F",X"EF",X"1F",X"EF",
		X"1F",X"EF",X"00",X"10",X"00",X"10",X"00",X"10",X"00",X"10",X"00",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"01",X"06",X"01",X"0F",X"B8",X"06",X"09",X"95",X"7A",X"97",X"7A",
		X"97",X"C0",X"10",X"9C",X"00",X"21",X"10",X"80",X"00",X"21",X"10",X"80",X"10",X"E1",X"06",X"00",
		X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"61",X"66",X"66",X"66",X"66",X"66",
		X"0F",X"01",X"06",X"04",X"01",X"06",X"04",X"01",X"05",X"03",X"01",X"06",X"03",X"1E",X"BC",X"1F",
		X"1C",X"C0",X"7A",X"97",X"9B",X"76",X"DA",X"10",X"E1",X"00",X"21",X"10",X"80",X"10",X"20",X"00",
		X"81",X"10",X"21",X"00",X"40",X"00",X"02",X"00",X"00",X"08",X"00",X"00",X"40",X"00",X"40",X"66",
		X"66",X"66",X"66",X"66",X"66",X"0F",X"01",X"06",X"06",X"01",X"06",X"01",X"01",X"06",X"01",X"01",
		X"06",X"06",X"1E",X"A0",X"04",X"06",X"2D",X"2D",X"21",X"21",X"21",X"C0",X"48",X"02",X"08",X"02",
		X"08",X"02",X"00",X"00",X"00",X"00",X"00",X"7E",X"00",X"00",X"40",X"00",X"00",X"44",X"00",X"07",
		X"00",X"00",X"00",X"00",X"24",X"24",X"24",X"A4",X"00",X"40",X"0E",X"01",X"03",X"03",X"03",X"06",
		X"04",X"03",X"06",X"06",X"08",X"36",X"17",X"36",X"26",X"36",X"35",X"36",X"44",X"36",X"53",X"36",
		X"62",X"36",X"71",X"36",X"80",X"36",X"8F",X"36",X"9E",X"36",X"AD",X"36",X"BC",X"36",X"CB",X"36",
		X"DA",X"36",X"E9",X"36",X"F8",X"36",X"07",X"37",X"01",X"18",X"15",X"20",X"03",X"01",X"28",X"01",
		X"20",X"01",X"18",X"01",X"10",X"01",X"08",X"01",X"17",X"14",X"19",X"03",X"01",X"10",X"02",X"10",
		X"02",X"10",X"02",X"10",X"01",X"10",X"01",X"16",X"13",X"16",X"03",X"01",X"0C",X"03",X"0D",X"03",
		X"0E",X"03",X"0F",X"02",X"10",X"01",X"15",X"12",X"14",X"03",X"02",X"0B",X"04",X"0C",X"04",X"0D",
		X"04",X"0E",X"03",X"0F",X"01",X"14",X"11",X"12",X"03",X"03",X"0A",X"05",X"0B",X"05",X"0C",X"05",
		X"0D",X"04",X"0E",X"01",X"13",X"10",X"10",X"02",X"01",X"09",X"02",X"0A",X"03",X"0B",X"04",X"0C",
		X"05",X"0D",X"01",X"12",X"0F",X"0E",X"02",X"03",X"08",X"04",X"09",X"04",X"0A",X"05",X"0B",X"05",
		X"0C",X"01",X"11",X"0E",X"0C",X"02",X"04",X"07",X"04",X"08",X"04",X"09",X"05",X"0A",X"05",X"0B",
		X"01",X"10",X"0D",X"0A",X"02",X"04",X"06",X"05",X"07",X"05",X"08",X"05",X"09",X"04",X"0A",X"01",
		X"0F",X"0C",X"08",X"02",X"05",X"05",X"05",X"06",X"05",X"07",X"05",X"08",X"05",X"09",X"01",X"0E",
		X"0B",X"06",X"01",X"03",X"04",X"05",X"05",X"05",X"06",X"05",X"07",X"05",X"08",X"01",X"0D",X"0A",
		X"04",X"01",X"02",X"05",X"04",X"05",X"04",X"05",X"05",X"05",X"05",X"05",X"01",X"0C",X"09",X"03",
		X"01",X"03",X"03",X"05",X"04",X"05",X"05",X"04",X"06",X"04",X"07",X"01",X"0B",X"08",X"02",X"01",
		X"03",X"01",X"04",X"02",X"05",X"03",X"04",X"04",X"05",X"05",X"01",X"0A",X"07",X"01",X"01",X"05",
		X"01",X"05",X"01",X"05",X"01",X"05",X"01",X"05",X"01",X"01",X"20",X"20",X"80",X"01",X"05",X"72",
		X"04",X"66",X"01",X"32",X"02",X"40",X"03",X"50",X"01",X"20",X"20",X"14",X"01",X"01",X"10",X"04",
		X"15",X"02",X"36",X"03",X"10",X"05",X"13",X"01",X"20",X"20",X"20",X"01",X"03",X"03",X"02",X"30",
		X"04",X"08",X"01",X"28",X"05",X"12",X"F5",X"C5",X"D5",X"E5",X"F3",X"21",X"16",X"37",X"11",X"AF",
		X"A6",X"01",X"07",X"FF",X"DB",X"21",X"C3",X"2A",X"19",X"D5",X"E5",X"97",X"6F",X"67",X"32",X"A5",
		X"4E",X"32",X"A1",X"4C",X"FD",X"E1",X"3C",X"32",X"3C",X"4C",X"32",X"3D",X"4C",X"FD",X"7E",X"00",
		X"FD",X"23",X"5F",X"16",X"00",X"19",X"10",X"F5",X"0D",X"32",X"C0",X"50",X"20",X"EF",X"D1",X"19",
		X"7C",X"EB",X"E5",X"DD",X"E1",X"11",X"84",X"23",X"D5",X"FD",X"E1",X"FD",X"E9",X"DB",X"32",X"E1",
		X"D1",X"C1",X"F1",X"FB",X"C3",X"03",X"3C",X"3A",X"37",X"4C",X"FE",X"01",X"28",X"26",X"DD",X"21",
		X"93",X"4C",X"21",X"9B",X"4C",X"11",X"44",X"4C",X"06",X"03",X"7E",X"12",X"2B",X"1B",X"10",X"FA",
		X"CD",X"2B",X"3A",X"3A",X"91",X"4C",X"A7",X"20",X"08",X"CD",X"AA",X"37",X"CD",X"B1",X"37",X"18",
		X"06",X"CD",X"B1",X"37",X"CD",X"AA",X"37",X"3A",X"94",X"4C",X"FE",X"01",X"C0",X"97",X"32",X"94",
		X"4C",X"CD",X"0C",X"3B",X"06",X"B4",X"CD",X"72",X"03",X"C9",X"21",X"96",X"4C",X"3E",X"01",X"18",
		X"05",X"21",X"99",X"4C",X"3E",X"02",X"32",X"8A",X"4C",X"CD",X"58",X"02",X"11",X"45",X"4C",X"06",
		X"03",X"7E",X"12",X"23",X"13",X"10",X"FA",X"CD",X"D6",X"37",X"C9",X"DB",X"02",X"DB",X"00",X"F1",
		X"C1",X"D1",X"E1",X"C3",X"3F",X"02",X"3A",X"93",X"4C",X"FE",X"0A",X"28",X"04",X"3C",X"32",X"93",
		X"4C",X"DD",X"21",X"7E",X"4C",X"21",X"45",X"4C",X"11",X"42",X"4C",X"06",X"03",X"7E",X"12",X"23",
		X"13",X"10",X"FA",X"CD",X"2B",X"3A",X"3A",X"91",X"4C",X"A7",X"C8",X"3E",X"01",X"32",X"94",X"4C",
		X"11",X"89",X"4C",X"06",X"03",X"2B",X"7E",X"12",X"1B",X"10",X"FA",X"97",X"12",X"1B",X"12",X"1B",
		X"12",X"CD",X"18",X"38",X"CD",X"D2",X"39",X"C9",X"97",X"CD",X"B4",X"02",X"CD",X"12",X"06",X"32",
		X"8C",X"4C",X"11",X"71",X"3A",X"21",X"86",X"42",X"CD",X"6B",X"04",X"3A",X"8A",X"4C",X"FE",X"01",
		X"3E",X"32",X"20",X"01",X"3D",X"32",X"87",X"41",X"3E",X"0B",X"CD",X"7A",X"09",X"CD",X"A1",X"03",
		X"11",X"A4",X"3A",X"21",X"8A",X"43",X"CD",X"6B",X"04",X"11",X"9B",X"3A",X"21",X"52",X"42",X"CD",
		X"6B",X"04",X"11",X"8C",X"3A",X"21",X"DA",X"42",X"CD",X"6B",X"04",X"3E",X"30",X"32",X"8B",X"4C",
		X"CD",X"B2",X"39",X"3E",X"14",X"32",X"8D",X"4C",X"11",X"90",X"4C",X"3E",X"01",X"32",X"8F",X"4C",
		X"3E",X"41",X"12",X"CD",X"8C",X"39",X"06",X"3C",X"32",X"0A",X"4C",X"CD",X"64",X"39",X"3A",X"8C",
		X"4C",X"FE",X"01",X"C8",X"CD",X"7C",X"02",X"CB",X"6F",X"20",X"3B",X"3A",X"8F",X"4C",X"E6",X"01",
		X"3E",X"14",X"28",X"02",X"3E",X"17",X"CD",X"7A",X"09",X"3A",X"8F",X"4C",X"21",X"83",X"4C",X"85",
		X"6F",X"7C",X"CE",X"00",X"67",X"1A",X"77",X"3A",X"8F",X"4C",X"FE",X"03",X"C8",X"3C",X"32",X"8F",
		X"4C",X"CD",X"7C",X"02",X"CB",X"6F",X"20",X"0B",X"CD",X"64",X"39",X"3A",X"8C",X"4C",X"FE",X"01",
		X"C8",X"18",X"EE",X"CD",X"8C",X"39",X"CD",X"7C",X"02",X"CB",X"5F",X"20",X"0B",X"1A",X"3D",X"FE",
		X"2F",X"20",X"02",X"3E",X"5B",X"12",X"18",X"0F",X"CD",X"7C",X"02",X"CB",X"47",X"20",X"9C",X"1A",
		X"3C",X"FE",X"5C",X"20",X"02",X"3E",X"30",X"12",X"CD",X"8C",X"39",X"3A",X"8D",X"4C",X"FE",X"06",
		X"38",X"05",X"3D",X"3D",X"32",X"8D",X"4C",X"32",X"8E",X"4C",X"CD",X"7C",X"02",X"32",X"C0",X"50",
		X"CB",X"5F",X"28",X"0C",X"CB",X"47",X"28",X"08",X"3E",X"14",X"32",X"8D",X"4C",X"C3",X"7B",X"38",
		X"3A",X"0A",X"4C",X"A7",X"20",X"FA",X"3E",X"01",X"32",X"0A",X"4C",X"10",X"13",X"06",X"3C",X"3A",
		X"8B",X"4C",X"D6",X"01",X"27",X"32",X"8B",X"4C",X"CD",X"B2",X"39",X"3A",X"8B",X"4C",X"A7",X"C8",
		X"21",X"8E",X"4C",X"35",X"20",X"C4",X"3A",X"8D",X"4C",X"FE",X"06",X"38",X"05",X"3D",X"3D",X"32",
		X"8D",X"4C",X"77",X"CD",X"7C",X"02",X"CB",X"5F",X"20",X"0B",X"1A",X"3D",X"FE",X"2F",X"20",X"02",
		X"3E",X"5B",X"12",X"18",X"08",X"1A",X"3C",X"FE",X"5C",X"20",X"02",X"3E",X"30",X"12",X"CD",X"8C",
		X"39",X"C3",X"FA",X"38",X"3A",X"0A",X"4C",X"32",X"C0",X"50",X"A7",X"20",X"F7",X"3E",X"01",X"32",
		X"0A",X"4C",X"10",X"17",X"06",X"3C",X"3A",X"8B",X"4C",X"D6",X"01",X"27",X"32",X"8B",X"4C",X"CD",
		X"B2",X"39",X"A7",X"28",X"01",X"C9",X"3E",X"01",X"32",X"8C",X"4C",X"C9",X"F5",X"C5",X"E5",X"21",
		X"52",X"42",X"3A",X"8F",X"4C",X"FE",X"02",X"20",X"03",X"21",X"12",X"42",X"FE",X"03",X"20",X"03",
		X"21",X"D2",X"41",X"3E",X"09",X"32",X"02",X"4C",X"3A",X"90",X"4C",X"CD",X"1A",X"04",X"E1",X"C1",
		X"F1",X"C9",X"21",X"5A",X"41",X"F5",X"97",X"32",X"08",X"4C",X"3A",X"95",X"4C",X"3C",X"FE",X"0F",
		X"38",X"02",X"3E",X"03",X"32",X"95",X"4C",X"32",X"02",X"4C",X"3A",X"8B",X"4C",X"CD",X"F3",X"03",
		X"F1",X"C9",X"01",X"0A",X"0A",X"DD",X"21",X"48",X"4C",X"21",X"4D",X"4C",X"11",X"4E",X"4C",X"32",
		X"C0",X"50",X"C5",X"06",X"06",X"E5",X"21",X"3F",X"4C",X"1A",X"77",X"13",X"23",X"10",X"FA",X"E1",
		X"1B",X"CD",X"2B",X"3A",X"3A",X"91",X"4C",X"FE",X"01",X"20",X"1D",X"06",X"06",X"7E",X"12",X"2B",
		X"1B",X"10",X"FA",X"23",X"13",X"06",X"06",X"D5",X"11",X"3F",X"4C",X"1A",X"77",X"13",X"23",X"10",
		X"FA",X"D1",X"2B",X"13",X"13",X"13",X"13",X"13",X"13",X"D5",X"11",X"06",X"00",X"19",X"DD",X"19",
		X"D1",X"C1",X"10",X"BB",X"06",X"0A",X"0D",X"C2",X"D5",X"39",X"C9",X"F5",X"D5",X"E5",X"21",X"08",
		X"4C",X"97",X"77",X"32",X"91",X"4C",X"11",X"44",X"4C",X"1A",X"DD",X"96",X"05",X"27",X"F5",X"A7",
		X"28",X"03",X"3E",X"01",X"77",X"F1",X"1B",X"1A",X"DD",X"9E",X"04",X"27",X"F5",X"A7",X"28",X"03",
		X"3E",X"01",X"77",X"F1",X"1B",X"1A",X"DD",X"9E",X"03",X"27",X"F5",X"A7",X"28",X"03",X"3E",X"01",
		X"77",X"F1",X"38",X"09",X"7E",X"A7",X"28",X"05",X"3E",X"01",X"32",X"91",X"4C",X"E1",X"D1",X"F1",
		X"C9",X"FF",X"03",X"47",X"52",X"45",X"41",X"54",X"20",X"53",X"43",X"4F",X"52",X"45",X"FF",X"FE",
		X"50",X"4C",X"41",X"59",X"45",X"52",X"20",X"20",X"20",X"21",X"FF",X"FF",X"FF",X"05",X"54",X"49",
		X"4D",X"45",X"20",X"4C",X"45",X"46",X"54",X"FF",X"09",X"FF",X"FF",X"FF",X"06",X"5F",X"20",X"5F",
		X"20",X"5F",X"FF",X"FF",X"FF",X"06",X"4D",X"4F",X"56",X"45",X"20",X"4A",X"4F",X"59",X"53",X"54",
		X"49",X"43",X"4B",X"20",X"FF",X"0D",X"55",X"50",X"20",X"FF",X"06",X"4F",X"52",X"20",X"FF",X"08",
		X"44",X"4F",X"57",X"4E",X"FF",X"06",X"FF",X"FE",X"54",X"4F",X"20",X"53",X"45",X"4C",X"45",X"43",
		X"54",X"20",X"4C",X"45",X"54",X"54",X"45",X"52",X"53",X"2E",X"FF",X"FE",X"48",X"49",X"54",X"20",
		X"FF",X"0E",X"43",X"41",X"4C",X"4C",X"20",X"FF",X"06",X"54",X"4F",X"20",X"45",X"4E",X"54",X"45",
		X"52",X"20",X"49",X"4E",X"49",X"54",X"49",X"41",X"4C",X"53",X"2E",X"FF",X"FF",X"FF",X"09",X"4D",
		X"4F",X"42",X"20",X"4D",X"41",X"53",X"48",X"45",X"52",X"53",X"FF",X"FF",X"97",X"CD",X"BD",X"02",
		X"CD",X"12",X"06",X"11",X"FD",X"3A",X"21",X"86",X"42",X"CD",X"6B",X"04",X"01",X"01",X"0A",X"11",
		X"4B",X"4C",X"21",X"09",X"43",X"E5",X"CD",X"3E",X"3B",X"21",X"06",X"00",X"19",X"EB",X"E1",X"23",
		X"23",X"3A",X"93",X"4C",X"B9",X"C8",X"79",X"C6",X"01",X"27",X"4F",X"10",X"E8",X"C9",X"C5",X"D5",
		X"3E",X"01",X"32",X"08",X"4C",X"3E",X"0D",X"32",X"02",X"4C",X"79",X"CD",X"F3",X"03",X"3E",X"2E",
		X"CD",X"1A",X"04",X"01",X"C0",X"FF",X"09",X"3E",X"01",X"32",X"08",X"4C",X"3E",X"06",X"32",X"02",
		X"4C",X"CD",X"D9",X"03",X"01",X"60",X"FF",X"09",X"3E",X"0E",X"32",X"02",X"4C",X"06",X"03",X"1B",
		X"1A",X"CD",X"1A",X"04",X"C5",X"01",X"40",X"00",X"09",X"C1",X"10",X"F3",X"D1",X"C1",X"C9",X"E5",
		X"D5",X"C5",X"F5",X"11",X"06",X"53",X"21",X"93",X"3B",X"01",X"04",X"00",X"DB",X"01",X"DB",X"03",
		X"C3",X"C1",X"04",X"3E",X"01",X"32",X"14",X"4C",X"32",X"4B",X"4D",X"CD",X"5E",X"02",X"3A",X"80",
		X"50",X"CB",X"6F",X"3E",X"01",X"28",X"01",X"97",X"32",X"15",X"4C",X"97",X"32",X"31",X"4C",X"3C",
		X"32",X"16",X"4C",X"3E",X"19",X"32",X"4C",X"4D",X"3E",X"10",X"CD",X"EF",X"3B",X"32",X"16",X"4C",
		X"F3",X"DB",X"C9",X"DB",X"CB",X"3E",X"66",X"00",X"D6",X"65",X"47",X"DB",X"DC",X"DB",X"E6",X"FB",
		X"78",X"32",X"31",X"4C",X"32",X"4C",X"4D",X"3E",X"11",X"CD",X"EF",X"3B",X"CD",X"0C",X"3B",X"CD",
		X"12",X"06",X"CD",X"49",X"06",X"CD",X"41",X"3E",X"0E",X"08",X"CD",X"2B",X"03",X"18",X"BC",X"32",
		X"4E",X"4D",X"3E",X"01",X"32",X"4B",X"4D",X"32",X"3C",X"4C",X"32",X"3E",X"4C",X"CD",X"C3",X"27",
		X"C3",X"16",X"37",X"3A",X"00",X"4C",X"47",X"97",X"21",X"18",X"4C",X"11",X"04",X"00",X"77",X"19",
		X"10",X"FC",X"CD",X"E9",X"05",X"CD",X"49",X"06",X"97",X"32",X"A3",X"4C",X"3E",X"09",X"CD",X"0E",
		X"05",X"CD",X"C4",X"05",X"3A",X"17",X"4C",X"FE",X"01",X"28",X"08",X"3E",X"09",X"CD",X"16",X"05",
		X"CD",X"CC",X"05",X"3E",X"01",X"32",X"A3",X"4C",X"CD",X"B0",X"2E",X"97",X"C9",X"F5",X"C5",X"E5",
		X"3A",X"2C",X"4F",X"07",X"07",X"06",X"00",X"4F",X"21",X"18",X"4C",X"09",X"7E",X"A7",X"20",X"48",
		X"E5",X"3A",X"31",X"4C",X"A7",X"21",X"A7",X"3C",X"28",X"08",X"FE",X"01",X"21",X"4B",X"3D",X"28",
		X"01",X"FF",X"CB",X"19",X"09",X"4E",X"23",X"46",X"E1",X"E5",X"23",X"23",X"71",X"23",X"70",X"E1",
		X"E5",X"23",X"23",X"4E",X"23",X"46",X"E1",X"F3",X"DB",X"97",X"0A",X"5F",X"DB",X"C8",X"FB",X"7B",
		X"A7",X"28",X"BD",X"E5",X"3C",X"77",X"03",X"23",X"F3",X"DB",X"97",X"0A",X"5F",X"DB",X"C8",X"FB",
		X"7B",X"77",X"03",X"23",X"71",X"23",X"70",X"E1",X"35",X"28",X"D5",X"23",X"7E",X"32",X"30",X"4C",
		X"CD",X"49",X"03",X"E1",X"C1",X"F1",X"C9",X"B3",X"3C",X"2C",X"3D",X"19",X"3D",X"F4",X"3C",X"FB",
		X"3C",X"0A",X"3D",X"10",X"80",X"05",X"85",X"4B",X"84",X"05",X"80",X"05",X"88",X"19",X"80",X"05",
		X"84",X"1E",X"87",X"05",X"85",X"04",X"80",X"14",X"90",X"08",X"80",X"19",X"85",X"08",X"90",X"1E",
		X"80",X"05",X"84",X"16",X"80",X"0E",X"90",X"2F",X"80",X"05",X"84",X"08",X"80",X"10",X"90",X"14",
		X"80",X"0A",X"85",X"05",X"80",X"0A",X"88",X"10",X"80",X"0A",X"90",X"19",X"80",X"0A",X"90",X"1C",
		X"80",X"23",X"84",X"FF",X"0A",X"80",X"18",X"84",X"64",X"80",X"FF",X"0A",X"80",X"0C",X"84",X"09",
		X"80",X"05",X"88",X"04",X"80",X"12",X"84",X"64",X"80",X"FF",X"05",X"80",X"14",X"84",X"0A",X"87",
		X"14",X"84",X"0A",X"86",X"05",X"85",X"64",X"80",X"FF",X"0A",X"80",X"05",X"84",X"05",X"80",X"05",
		X"88",X"10",X"80",X"05",X"84",X"0A",X"86",X"05",X"84",X"64",X"80",X"FF",X"0A",X"80",X"0C",X"85",
		X"05",X"80",X"05",X"88",X"08",X"80",X"04",X"84",X"05",X"86",X"05",X"87",X"14",X"84",X"05",X"80",
		X"05",X"88",X"08",X"80",X"04",X"85",X"0A",X"86",X"10",X"84",X"FF",X"57",X"3D",X"B2",X"3D",X"FF",
		X"3D",X"C3",X"3D",X"E6",X"3D",X"28",X"3E",X"05",X"80",X"0A",X"85",X"05",X"84",X"0A",X"87",X"05",
		X"85",X"05",X"84",X"0A",X"87",X"05",X"85",X"05",X"84",X"0A",X"87",X"05",X"85",X"05",X"84",X"0A",
		X"87",X"05",X"85",X"05",X"84",X"08",X"87",X"03",X"86",X"02",X"87",X"04",X"86",X"07",X"87",X"05",
		X"80",X"1E",X"85",X"05",X"84",X"04",X"90",X"05",X"80",X"0A",X"84",X"0A",X"86",X"0F",X"85",X"03",
		X"80",X"05",X"88",X"10",X"80",X"05",X"85",X"14",X"80",X"0A",X"85",X"14",X"80",X"05",X"88",X"04",
		X"80",X"05",X"90",X"05",X"80",X"05",X"85",X"0C",X"80",X"08",X"90",X"02",X"80",X"05",X"85",X"FF",
		X"FF",X"FF",X"02",X"80",X"08",X"85",X"30",X"84",X"02",X"80",X"28",X"85",X"28",X"84",X"30",X"85",
		X"FF",X"FF",X"FF",X"05",X"80",X"06",X"85",X"05",X"80",X"05",X"88",X"05",X"80",X"12",X"85",X"05",
		X"80",X"05",X"88",X"05",X"80",X"0C",X"84",X"0C",X"85",X"05",X"80",X"05",X"88",X"05",X"80",X"1E",
		X"84",X"05",X"80",X"FF",X"FF",X"FF",X"05",X"80",X"0A",X"84",X"0A",X"87",X"14",X"84",X"0C",X"80",
		X"37",X"85",X"32",X"84",X"0C",X"80",X"32",X"85",X"0A",X"87",X"05",X"84",X"05",X"80",X"FF",X"05",
		X"80",X"05",X"84",X"05",X"80",X"05",X"88",X"05",X"80",X"0A",X"85",X"05",X"80",X"05",X"88",X"05",
		X"80",X"0F",X"84",X"0A",X"87",X"0A",X"85",X"05",X"84",X"05",X"88",X"10",X"80",X"05",X"84",X"0A",
		X"86",X"28",X"85",X"05",X"80",X"05",X"84",X"FF",X"05",X"80",X"04",X"85",X"05",X"88",X"1C",X"80",
		X"04",X"85",X"28",X"87",X"0A",X"80",X"10",X"84",X"0C",X"84",X"0A",X"86",X"28",X"85",X"40",X"80",
		X"FF",X"21",X"9E",X"43",X"11",X"5C",X"3E",X"CD",X"6B",X"04",X"3A",X"80",X"50",X"E6",X"1C",X"EE",
		X"1C",X"0F",X"0F",X"C6",X"32",X"21",X"DE",X"41",X"CD",X"1A",X"04",X"C9",X"FF",X"0B",X"42",X"4F",
		X"4E",X"55",X"53",X"20",X"47",X"4C",X"4F",X"42",X"20",X"41",X"54",X"20",X"30",X"30",X"30",X"30",
		X"30",X"20",X"50",X"4F",X"49",X"4E",X"54",X"53",X"FF",X"FF",X"97",X"42",X"A7",X"3E",X"1E",X"F6",
		X"09",X"00",X"3F",X"00",X"00",X"40",X"3F",X"3F",X"3F",X"80",X"3F",X"3F",X"3E",X"C0",X"3F",X"3F",
		X"3D",X"80",X"3F",X"3F",X"3B",X"40",X"3F",X"3F",X"37",X"C0",X"3F",X"3F",X"2F",X"C0",X"3F",X"3F",
		X"1F",X"40",X"3F",X"3F",X"00",X"3F",X"FF",X"4D",X"45",X"45",X"54",X"20",X"54",X"48",X"45",X"20",
		X"47",X"4C",X"4F",X"42",X"FF",X"FF",X"4D",X"55",X"4E",X"43",X"48",X"20",X"41",X"4C",X"4C",X"20",
		X"54",X"48",X"45",X"20",X"53",X"4E",X"41",X"43",X"4B",X"53",X"FF",X"FE",X"54",X"4F",X"20",X"43",
		X"4C",X"45",X"41",X"52",X"20",X"54",X"48",X"45",X"20",X"4C",X"45",X"56",X"45",X"4C",X"FF",X"FF",
		X"50",X"55",X"53",X"48",X"20",X"43",X"41",X"4C",X"4C",X"20",X"42",X"55",X"54",X"54",X"4F",X"4E",
		X"FF",X"FE",X"54",X"4F",X"20",X"52",X"49",X"44",X"45",X"20",X"45",X"4C",X"45",X"56",X"41",X"54",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
