library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity spr_rom is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of spr_rom is
	type rom is array(0 to  32767) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"21",
		X"11",X"1F",X"FF",X"FF",X"FF",X"00",X"38",X"88",X"FF",X"FF",X"FF",X"FF",X"11",X"13",X"38",X"23",
		X"4F",X"FF",X"FF",X"04",X"33",X"22",X"11",X"12",X"4F",X"FF",X"00",X"33",X"99",X"21",X"11",X"78",
		X"1F",X"03",X"21",X"88",X"93",X"33",X"4F",X"FF",X"03",X"21",X"29",X"93",X"34",X"FF",X"FF",X"03",
		X"22",X"29",X"91",X"12",X"4F",X"FF",X"00",X"33",X"99",X"22",X"21",X"78",X"1F",X"04",X"44",X"33",
		X"33",X"33",X"4F",X"FF",X"11",X"14",X"43",X"33",X"4F",X"FF",X"FF",X"00",X"44",X"33",X"FF",X"FF",
		X"FF",X"FF",X"00",X"22",X"88",X"8F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"21",
		X"11",X"1F",X"FF",X"FF",X"FF",X"00",X"43",X"88",X"FF",X"FF",X"FF",X"FF",X"00",X"44",X"38",X"83",
		X"3F",X"FF",X"FF",X"02",X"11",X"12",X"22",X"22",X"3F",X"FF",X"01",X"13",X"33",X"31",X"11",X"17",
		X"1F",X"04",X"33",X"33",X"22",X"23",X"3F",X"FF",X"02",X"29",X"98",X"33",X"33",X"FF",X"FF",X"04",
		X"11",X"88",X"92",X"23",X"3F",X"FF",X"04",X"22",X"19",X"93",X"21",X"2A",X"1F",X"04",X"33",X"49",
		X"33",X"34",X"FF",X"FF",X"02",X"24",X"88",X"8F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"21",X"11",X"1F",X"FF",X"FF",X"FF",X"00",X"32",
		X"88",X"FF",X"FF",X"FF",X"FF",X"00",X"43",X"28",X"8F",X"FF",X"FF",X"FF",X"00",X"43",X"33",X"33",
		X"3F",X"FF",X"FF",X"02",X"21",X"12",X"22",X"33",X"3F",X"FF",X"01",X"11",X"32",X"21",X"12",X"27",
		X"1F",X"03",X"39",X"93",X"31",X"13",X"4F",X"FF",X"02",X"29",X"81",X"33",X"33",X"3F",X"FF",X"03",
		X"21",X"18",X"92",X"22",X"3B",X"1F",X"03",X"21",X"19",X"33",X"34",X"FF",X"FF",X"04",X"33",X"23",
		X"34",X"FF",X"FF",X"FF",X"02",X"2F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"21",
		X"11",X"1F",X"FF",X"FF",X"FF",X"00",X"33",X"88",X"FF",X"FF",X"FF",X"FF",X"00",X"33",X"38",X"8F",
		X"FF",X"FF",X"FF",X"04",X"43",X"71",X"33",X"3F",X"FF",X"FF",X"02",X"27",X"13",X"33",X"33",X"3F",
		X"FF",X"01",X"11",X"22",X"11",X"21",X"17",X"1F",X"05",X"49",X"92",X"22",X"22",X"4F",X"FF",X"02",
		X"29",X"18",X"33",X"44",X"3C",X"1F",X"03",X"38",X"19",X"22",X"33",X"FF",X"FF",X"04",X"23",X"99",
		X"44",X"FF",X"FF",X"FF",X"00",X"32",X"2F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"21",X"11",X"1F",X"FF",X"FF",X"FF",X"00",X"33",X"88",X"FF",
		X"FF",X"FF",X"FF",X"00",X"33",X"38",X"88",X"3F",X"FF",X"FF",X"03",X"44",X"33",X"33",X"33",X"5F",
		X"FF",X"03",X"37",X"12",X"22",X"22",X"27",X"1F",X"03",X"71",X"33",X"11",X"83",X"3C",X"1F",X"07",
		X"19",X"93",X"33",X"34",X"FF",X"FF",X"04",X"39",X"99",X"34",X"FF",X"FF",X"FF",X"03",X"21",X"49",
		X"FF",X"FF",X"FF",X"FF",X"00",X"32",X"2F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"00",X"21",X"11",X"1F",X"FF",X"FF",X"FF",X"00",X"08",X"88",X"35",X"5F",X"FF",
		X"FF",X"00",X"43",X"22",X"23",X"44",X"5F",X"FF",X"03",X"77",X"43",X"11",X"13",X"37",X"1F",X"07",
		X"74",X"32",X"22",X"33",X"FF",X"FF",X"07",X"43",X"99",X"44",X"FF",X"FF",X"FF",X"04",X"39",X"99",
		X"FF",X"FF",X"FF",X"FF",X"00",X"32",X"2F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"00",X"11",X"11",X"66",X"66",X"6F",X"FF",X"00",X"77",X"77",X"88",X"22",X"3A",X"1F",X"05",
		X"77",X"71",X"12",X"24",X"FF",X"FF",X"05",X"77",X"33",X"35",X"FF",X"FF",X"FF",X"05",X"39",X"94",
		X"FF",X"FF",X"FF",X"FF",X"00",X"43",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"ED",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",
		X"DA",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"ED",X"AA",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"DA",X"AA",X"AF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"08",X"55",X"ED",X"A2",X"EE",X"AA",X"AA",X"FF",X"00",X"00",X"00",X"00",X"08",X"8E",X"E2",X"22",
		X"EA",X"AA",X"A1",X"FF",X"00",X"00",X"00",X"55",X"55",X"BE",X"22",X"22",X"EE",X"BB",X"B2",X"FF",
		X"00",X"54",X"44",X"BB",X"BB",X"B6",X"22",X"A1",X"1A",X"33",X"FF",X"FF",X"66",X"55",X"77",X"7E",
		X"EE",X"BC",X"62",X"2A",X"A3",X"33",X"FF",X"FF",X"00",X"66",X"66",X"6C",X"CC",X"CC",X"63",X"33",
		X"33",X"33",X"FF",X"FF",X"00",X"00",X"00",X"66",X"6C",X"C6",X"55",X"53",X"33",X"3A",X"AA",X"FF",
		X"00",X"00",X"00",X"00",X"06",X"66",X"65",X"55",X"53",X"EA",X"A1",X"FF",X"00",X"00",X"00",X"00",
		X"06",X"66",X"66",X"65",X"55",X"CB",X"B2",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"66",
		X"66",X"5F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"53",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"63",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"56",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"48",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"04",X"84",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"48",
		X"44",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"84",X"44",X"4F",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"05",X"55",X"44",X"43",X"44",X"44",X"44",X"FF",X"00",X"00",X"00",X"00",
		X"05",X"54",X"43",X"33",X"44",X"44",X"4E",X"FF",X"00",X"00",X"00",X"55",X"55",X"B4",X"33",X"33",
		X"44",X"BB",X"B3",X"FF",X"00",X"54",X"44",X"BB",X"BB",X"B0",X"33",X"4E",X"E4",X"55",X"FF",X"FF",
		X"00",X"55",X"55",X"54",X"44",X"B0",X"03",X"34",X"45",X"55",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"05",X"55",X"55",X"55",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",
		X"55",X"54",X"44",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"55",X"55",X"44",X"4E",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"55",X"0B",X"B3",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"5F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"5F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"55",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"55",X"55",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"55",
		X"55",X"5F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"05",X"55",X"55",X"55",X"55",X"54",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"FF",X"00",X"05",X"55",X"55",X"55",X"50",X"55",X"54",
		X"45",X"FF",X"FF",X"FF",X"00",X"00",X"50",X"00",X"55",X"50",X"05",X"55",X"5F",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"05",X"55",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"55",X"54",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"55",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"00",X"BB",X"BB",X"BF",X"FF",X"FF",X"09",X"9B",X"BE",X"EE",X"FF",X"FF",X"39",X"9E",
		X"16",X"DE",X"EF",X"FF",X"43",X"EE",X"11",X"67",X"EF",X"FF",X"43",X"E5",X"E1",X"67",X"EF",X"FF",
		X"33",X"75",X"71",X"67",X"EF",X"FF",X"43",X"75",X"D1",X"6E",X"EF",X"FF",X"43",X"77",X"11",X"6E",
		X"EF",X"FF",X"38",X"87",X"16",X"BB",X"EF",X"FF",X"08",X"89",X"99",X"BB",X"FF",X"FF",X"00",X"99",
		X"99",X"9F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"BB",X"BB",X"BF",X"FF",X"FF",X"09",X"9B",X"BE",X"EE",X"FF",X"FF",X"39",X"9E",X"16",X"DE",
		X"EF",X"FF",X"23",X"EE",X"11",X"67",X"EF",X"FF",X"23",X"E5",X"E1",X"67",X"EF",X"FF",X"33",X"75",
		X"71",X"67",X"EF",X"FF",X"23",X"75",X"D1",X"6E",X"EF",X"FF",X"23",X"77",X"11",X"6E",X"EF",X"FF",
		X"38",X"87",X"16",X"BB",X"EF",X"FF",X"08",X"89",X"99",X"BB",X"FF",X"FF",X"00",X"99",X"99",X"9F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"BB",
		X"BB",X"BF",X"FF",X"FF",X"09",X"9B",X"BE",X"EE",X"FF",X"FF",X"39",X"9E",X"16",X"DE",X"EF",X"FF",
		X"63",X"EE",X"11",X"67",X"EF",X"FF",X"63",X"E5",X"E1",X"67",X"EF",X"FF",X"33",X"75",X"71",X"67",
		X"EF",X"FF",X"63",X"75",X"D1",X"6E",X"EF",X"FF",X"63",X"77",X"11",X"6E",X"EF",X"FF",X"38",X"87",
		X"16",X"BB",X"EF",X"FF",X"08",X"89",X"99",X"BB",X"FF",X"FF",X"00",X"99",X"99",X"9F",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"AF",X"BB",X"DF",X"AA",X"AF",X"FF",X"FF",
		X"FF",X"FF",X"AA",X"FF",X"BB",X"DF",X"AA",X"AF",X"AA",X"FF",X"AA",X"AF",X"BB",X"DF",X"AA",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"44",X"44",X"FF",X"FF",X"00",X"00",
		X"54",X"42",X"2F",X"FF",X"00",X"00",X"05",X"44",X"33",X"DF",X"00",X"05",X"55",X"3A",X"AA",X"AF",
		X"05",X"54",X"44",X"35",X"69",X"8F",X"65",X"2A",X"12",X"35",X"55",X"FF",X"65",X"22",X"A1",X"35",
		X"33",X"FF",X"06",X"53",X"22",X"65",X"33",X"DF",X"00",X"06",X"66",X"5A",X"AA",X"AF",X"00",X"00",
		X"06",X"56",X"59",X"8F",X"00",X"00",X"55",X"53",X"3F",X"FF",X"00",X"00",X"66",X"55",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"B0",X"9F",X"FF",X"FF",X"FF",
		X"00",X"0B",X"BE",X"99",X"FF",X"FF",X"FF",X"00",X"0B",X"BE",X"99",X"FF",X"FF",X"FF",X"00",X"00",
		X"ED",X"E0",X"FF",X"FF",X"FF",X"00",X"0C",X"CE",X"AA",X"FF",X"FF",X"FF",X"00",X"0C",X"CE",X"AA",
		X"FF",X"FF",X"FF",X"00",X"00",X"C0",X"AF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"B0",X"9F",X"FF",X"FF",X"FF",
		X"00",X"0B",X"BE",X"99",X"FF",X"FF",X"FF",X"00",X"BB",X"AE",X"99",X"9F",X"FF",X"FF",X"00",X"BA",
		X"EE",X"E9",X"9F",X"FF",X"FF",X"00",X"0E",X"ED",X"EE",X"0F",X"FF",X"FF",X"00",X"CB",X"EE",X"E9",
		X"AF",X"FF",X"FF",X"00",X"CC",X"BE",X"9A",X"AF",X"FF",X"FF",X"00",X"0C",X"CE",X"AA",X"FF",X"FF",
		X"FF",X"00",X"00",X"C0",X"AF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"B0",X"9F",X"FF",X"FF",X"FF",
		X"00",X"0B",X"AE",X"99",X"FF",X"FF",X"FF",X"00",X"BA",X"AE",X"79",X"9F",X"FF",X"FF",X"0B",X"AA",
		X"EE",X"E7",X"99",X"FF",X"FF",X"0B",X"AE",X"ED",X"EE",X"79",X"FF",X"FF",X"00",X"EE",X"DD",X"DE",
		X"EF",X"FF",X"FF",X"0C",X"BE",X"ED",X"EE",X"9A",X"FF",X"FF",X"0C",X"BB",X"EE",X"E9",X"AA",X"FF",
		X"FF",X"00",X"CB",X"BE",X"9A",X"AF",X"FF",X"FF",X"00",X"0C",X"BE",X"AA",X"FF",X"FF",X"FF",X"00",
		X"00",X"C0",X"AF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"0A",X"A0",X"77",X"FF",X"FF",X"FF",
		X"00",X"A9",X"9E",X"77",X"7F",X"FF",X"FF",X"0A",X"99",X"9E",X"66",X"67",X"FF",X"FF",X"0A",X"99",
		X"EE",X"E6",X"67",X"FF",X"FF",X"09",X"9E",X"ED",X"EE",X"67",X"FF",X"FF",X"00",X"EE",X"DD",X"DE",
		X"EF",X"FF",X"FF",X"00",X"EE",X"DD",X"DE",X"EF",X"FF",X"FF",X"0A",X"AE",X"ED",X"EE",X"78",X"FF",
		X"FF",X"0A",X"AA",X"EE",X"E7",X"78",X"FF",X"FF",X"0B",X"AA",X"AE",X"77",X"88",X"FF",X"FF",X"00",
		X"BA",X"AE",X"88",X"8F",X"FF",X"FF",X"00",X"0B",X"A0",X"88",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"0A",X"50",X"06",X"7F",X"FF",X"FF",
		X"00",X"A9",X"5E",X"E5",X"67",X"FF",X"FF",X"0A",X"98",X"5E",X"E4",X"56",X"7F",X"FF",X"A9",X"87",
		X"5E",X"E3",X"45",X"67",X"FF",X"98",X"76",X"EE",X"EE",X"34",X"56",X"FF",X"AA",X"AE",X"ED",X"DE",
		X"E7",X"77",X"FF",X"0E",X"EE",X"DD",X"DD",X"EE",X"EF",X"FF",X"0E",X"EE",X"DD",X"DD",X"EE",X"EF",
		X"FF",X"BA",X"7E",X"ED",X"DE",X"E3",X"56",X"FF",X"BA",X"87",X"EE",X"EE",X"45",X"67",X"FF",X"BA",
		X"98",X"6E",X"EA",X"56",X"79",X"FF",X"0B",X"A9",X"8E",X"EA",X"67",X"9F",X"FF",X"00",X"BA",X"9E",
		X"EA",X"79",X"FF",X"FF",X"00",X"0B",X"A0",X"0A",X"9F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"09",X"30",X"04",X"5F",X"FF",X"FF",X"00",X"98",X"3E",X"E3",X"45",X"FF",X"FF",X"09",X"87",
		X"3E",X"E2",X"34",X"5F",X"FF",X"98",X"76",X"3E",X"E1",X"23",X"45",X"FF",X"87",X"65",X"EE",X"EE",
		X"11",X"34",X"FF",X"AA",X"AE",X"ED",X"DE",X"E1",X"13",X"FF",X"0E",X"EE",X"DD",X"DD",X"E6",X"66",
		X"FF",X"0E",X"EE",X"DD",X"DD",X"EE",X"EF",X"FF",X"BB",X"BE",X"DD",X"DD",X"EE",X"EF",X"FF",X"87",
		X"6E",X"ED",X"DE",X"E1",X"11",X"FF",X"98",X"76",X"EE",X"EE",X"23",X"45",X"FF",X"A9",X"87",X"5E",
		X"E2",X"34",X"56",X"FF",X"0A",X"98",X"5E",X"E3",X"45",X"6F",X"FF",X"00",X"A9",X"5E",X"E4",X"56",
		X"FF",X"FF",X"00",X"0A",X"50",X"06",X"6F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"03",X"33",X"33",X"33",X"33",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"02",X"22",X"22",X"22",X"22",X"22",X"32",X"2F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"0C",X"CC",
		X"CC",X"53",X"CC",X"3C",X"CC",X"32",X"22",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"CC",X"CC",X"CC",
		X"33",X"C3",X"3C",X"CC",X"33",X"22",X"2F",X"FF",X"FF",X"00",X"00",X"0C",X"CC",X"CC",X"CC",X"CC",
		X"CC",X"CC",X"CC",X"C3",X"31",X"22",X"FF",X"FF",X"00",X"00",X"CC",X"C2",X"CC",X"33",X"33",X"33",
		X"33",X"33",X"2C",X"33",X"11",X"2F",X"FF",X"00",X"0C",X"CC",X"22",X"C7",X"33",X"33",X"33",X"33",
		X"32",X"22",X"C3",X"31",X"1F",X"FF",X"00",X"CC",X"C3",X"22",X"C7",X"33",X"33",X"33",X"33",X"22",
		X"22",X"2C",X"33",X"3C",X"FF",X"0C",X"CC",X"33",X"22",X"CC",X"33",X"33",X"33",X"32",X"22",X"22",
		X"22",X"CC",X"CC",X"FF",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"E1",X"11",X"22",X"22",
		X"22",X"EC",X"FF",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"71",X"11",X"11",X"22",X"2E",
		X"EE",X"FF",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"77",X"71",X"11",X"11",X"EE",X"EE",
		X"EF",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"33",X"DD",X"77",X"11",X"1E",X"EE",X"EE",X"EF",
		X"00",X"00",X"00",X"00",X"00",X"03",X"33",X"23",X"33",X"D7",X"7C",X"EE",X"EE",X"EE",X"EF",X"00",
		X"00",X"00",X"00",X"00",X"33",X"22",X"12",X"23",X"3D",X"7C",X"EE",X"EE",X"EE",X"EF",X"00",X"00",
		X"00",X"00",X"00",X"32",X"21",X"11",X"22",X"3D",X"77",X"CC",X"CC",X"CC",X"CF",X"00",X"00",X"00",
		X"00",X"03",X"32",X"11",X"11",X"12",X"33",X"D7",X"77",X"77",X"77",X"7F",X"00",X"00",X"00",X"00",
		X"03",X"32",X"11",X"11",X"12",X"33",X"D7",X"77",X"77",X"77",X"7F",X"00",X"00",X"00",X"00",X"00",
		X"32",X"21",X"11",X"22",X"3D",X"77",X"11",X"11",X"11",X"1F",X"00",X"00",X"00",X"00",X"00",X"33",
		X"22",X"12",X"23",X"3D",X"75",X"55",X"55",X"55",X"5F",X"00",X"00",X"00",X"00",X"00",X"03",X"33",
		X"23",X"33",X"D7",X"7E",X"55",X"55",X"55",X"5F",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"33",
		X"DD",X"77",X"EC",X"C5",X"55",X"55",X"5F",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"77",
		X"7E",X"CC",X"CC",X"55",X"55",X"5F",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"7E",X"EC",
		X"CC",X"CC",X"C5",X"55",X"FF",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"C3",X"CC",X"CC",
		X"CC",X"CC",X"5C",X"FF",X"0C",X"CC",X"33",X"CC",X"CC",X"55",X"55",X"55",X"5C",X"CC",X"CC",X"CC",
		X"33",X"CC",X"FF",X"00",X"CC",X"C3",X"CC",X"C7",X"55",X"55",X"55",X"55",X"CC",X"CC",X"C3",X"33",
		X"3C",X"FF",X"00",X"0C",X"CC",X"CC",X"C7",X"55",X"55",X"55",X"55",X"5C",X"CC",X"33",X"35",X"5F",
		X"FF",X"00",X"00",X"CC",X"CC",X"CC",X"55",X"55",X"55",X"55",X"55",X"33",X"33",X"55",X"5F",X"FF",
		X"00",X"00",X"0C",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"33",X"35",X"55",X"FF",X"FF",X"00",
		X"00",X"00",X"CC",X"CC",X"CC",X"C5",X"5C",X"55",X"CC",X"33",X"55",X"5F",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"CC",X"CC",X"CC",X"5C",X"C5",X"CC",X"33",X"55",X"FF",X"FF",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"CC",X"CC",X"CC",X"CC",X"CC",X"33",X"5F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"05",X"55",X"55",X"55",X"55",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"00",X"00",X"00",X"03",X"36",X"66",X"66",X"66",X"66",X"66",X"6F",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"03",X"36",X"66",X"66",X"66",X"66",X"66",X"66",X"6F",X"FF",X"FF",
		X"FF",X"00",X"00",X"00",X"03",X"36",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"33",X"36",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"6F",X"FF",X"FF",X"00",
		X"00",X"33",X"31",X"13",X"33",X"33",X"13",X"33",X"30",X"00",X"06",X"66",X"FF",X"FF",X"06",X"33",
		X"33",X"11",X"11",X"33",X"33",X"13",X"33",X"30",X"00",X"03",X"66",X"6F",X"FF",X"06",X"63",X"31",
		X"11",X"11",X"33",X"33",X"13",X"33",X"33",X"00",X"03",X"36",X"66",X"FF",X"06",X"66",X"11",X"11",
		X"11",X"13",X"33",X"13",X"33",X"33",X"33",X"33",X"33",X"33",X"3F",X"06",X"66",X"61",X"11",X"11",
		X"00",X"00",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"66",X"66",X"66",X"11",X"10",X"00",
		X"06",X"16",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"66",X"66",X"66",X"61",X"00",X"06",X"61",
		X"13",X"66",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"66",X"66",X"66",X"60",X"00",X"63",X"31",X"13",
		X"33",X"6F",X"FF",X"FF",X"FF",X"FF",X"FF",X"66",X"66",X"66",X"66",X"06",X"33",X"21",X"11",X"23",
		X"36",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"06",X"32",X"11",X"11",X"12",X"36",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"1F",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"06",X"32",X"11",X"11",X"12",X"36",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"06",X"33",X"21",X"11",X"23",X"36",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"63",X"33",X"11",X"33",X"6F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"11",X"10",X"06",X"63",X"11",X"66",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"00",X"01",X"11",X"11",X"00",X"06",X"16",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"22",X"21",X"11",X"11",X"00",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"02",X"22",
		X"22",X"21",X"11",X"00",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"02",X"22",
		X"22",X"22",X"33",X"13",X"33",X"30",X"02",X"23",X"3F",X"FF",X"FF",X"00",X"33",X"30",X"22",X"22",
		X"23",X"33",X"13",X"33",X"30",X"02",X"23",X"FF",X"FF",X"FF",X"00",X"11",X"03",X"02",X"22",X"33",
		X"33",X"13",X"33",X"30",X"02",X"2F",X"FF",X"FF",X"FF",X"00",X"21",X"13",X"30",X"23",X"33",X"33",
		X"13",X"33",X"30",X"02",X"FF",X"FF",X"FF",X"FF",X"00",X"02",X"21",X"33",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"22",X"23",X"30",X"00",X"33",X"03",X"3F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"02",X"22",X"30",X"00",X"30",X"03",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"22",X"32",X"22",X"22",X"22",X"22",X"22",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"03",X"33",X"33",X"33",X"33",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"8F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"8F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"8F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"8F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"8F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"8F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"8F",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"8F",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"8F",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"8F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"88",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"88",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"08",X"88",X"88",X"8F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"08",X"88",X"88",X"88",X"88",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"08",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"8F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"08",X"88",X"88",X"88",X"88",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"88",X"88",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"08",
		X"88",X"8F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"88",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"88",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"8F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"8F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"8F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"8F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"8F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"8F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0B",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0B",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0B",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0B",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0B",X"1B",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",
		X"1B",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"BB",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"0B",X"BB",X"BB",X"BF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"0B",X"BB",X"BB",X"BB",X"BB",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"0B",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"BB",X"BF",X"FF",X"00",X"00",X"00",X"00",X"00",X"0B",X"BB",X"BB",X"BB",X"BB",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"BB",X"BB",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"BB",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"1B",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0B",X"1B",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"1B",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"1B",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"1B",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"1B",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"1F",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"1F",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"01",X"11",X"11",X"11",X"11",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"11",X"11",X"11",X"11",X"11",X"1F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"11",
		X"11",X"11",X"FF",X"FF",X"00",X"00",X"00",X"01",X"11",X"11",X"11",X"11",X"11",X"11",X"FF",X"FF",
		X"00",X"00",X"00",X"01",X"11",X"11",X"11",X"11",X"11",X"11",X"1F",X"FF",X"00",X"00",X"00",X"01",
		X"11",X"11",X"11",X"11",X"11",X"11",X"1F",X"FF",X"00",X"00",X"00",X"01",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"FF",X"00",X"00",X"00",X"01",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"FF",
		X"00",X"00",X"00",X"01",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"FF",X"00",X"00",X"00",X"00",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"FF",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"FF",X"00",X"00",X"00",X"00",X"01",X"11",X"11",X"11",X"11",X"11",X"1F",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"11",X"11",X"1F",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"01",X"11",X"11",X"11",X"11",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",
		X"11",X"1F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"1F",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"8F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"88",X"88",X"88",X"8F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"08",X"88",X"88",
		X"88",X"88",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"88",X"88",X"88",X"8F",X"FF",
		X"00",X"00",X"00",X"00",X"08",X"88",X"88",X"88",X"88",X"88",X"8F",X"FF",X"00",X"00",X"00",X"00",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"FF",X"00",X"00",X"00",X"00",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"FF",X"00",X"00",X"00",X"08",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"FF",
		X"00",X"00",X"00",X"08",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"FF",X"00",X"00",X"00",X"08",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"FF",X"00",X"00",X"00",X"08",X"88",X"88",X"88",X"88",
		X"88",X"88",X"8F",X"FF",X"00",X"00",X"00",X"08",X"88",X"88",X"88",X"88",X"88",X"88",X"8F",X"FF",
		X"00",X"00",X"00",X"08",X"88",X"88",X"88",X"88",X"88",X"88",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"88",X"88",X"88",X"88",X"88",X"88",X"FF",X"FF",X"00",X"00",X"00",X"00",X"88",X"88",X"88",X"88",
		X"88",X"8F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"08",X"88",X"88",X"88",X"88",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"88",X"8F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"88",X"8F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"11",X"11",X"11",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"01",X"01",X"11",X"11",X"11",X"11",X"1F",X"FF",X"FF",X"FF",X"FF",X"00",
		X"00",X"00",X"11",X"11",X"18",X"88",X"81",X"11",X"11",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"11",
		X"88",X"81",X"88",X"88",X"11",X"11",X"1F",X"FF",X"FF",X"00",X"00",X"01",X"18",X"88",X"81",X"88",
		X"88",X"11",X"11",X"10",X"01",X"FF",X"00",X"00",X"01",X"18",X"88",X"88",X"88",X"88",X"11",X"11",
		X"11",X"11",X"FF",X"00",X"00",X"11",X"11",X"88",X"18",X"88",X"88",X"11",X"88",X"11",X"1F",X"FF",
		X"00",X"00",X"01",X"18",X"81",X"11",X"18",X"88",X"18",X"81",X"81",X"1F",X"FF",X"00",X"00",X"01",
		X"18",X"81",X"11",X"18",X"81",X"18",X"88",X"81",X"11",X"FF",X"00",X"00",X"01",X"11",X"81",X"18",
		X"81",X"11",X"88",X"88",X"88",X"11",X"FF",X"00",X"00",X"11",X"11",X"11",X"88",X"81",X"18",X"88",
		X"88",X"88",X"81",X"FF",X"00",X"00",X"11",X"11",X"81",X"88",X"81",X"18",X"88",X"88",X"81",X"81",
		X"FF",X"00",X"01",X"11",X"18",X"88",X"88",X"81",X"18",X"88",X"88",X"88",X"11",X"FF",X"00",X"00",
		X"01",X"18",X"88",X"88",X"88",X"11",X"11",X"11",X"18",X"11",X"1F",X"00",X"00",X"01",X"11",X"88",
		X"88",X"88",X"11",X"11",X"11",X"11",X"11",X"FF",X"00",X"00",X"00",X"11",X"81",X"18",X"88",X"88",
		X"11",X"88",X"11",X"11",X"FF",X"00",X"00",X"00",X"11",X"11",X"88",X"88",X"88",X"88",X"88",X"11",
		X"1F",X"FF",X"00",X"00",X"01",X"11",X"11",X"88",X"88",X"88",X"88",X"88",X"81",X"1F",X"FF",X"00",
		X"00",X"00",X"10",X"11",X"11",X"88",X"88",X"88",X"88",X"11",X"11",X"FF",X"00",X"00",X"00",X"00",
		X"01",X"11",X"88",X"88",X"88",X"18",X"11",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"11",X"18",
		X"18",X"88",X"11",X"1F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"01",X"11",X"11",X"11",X"11",
		X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"11",X"11",X"11",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"01",X"FF",X"FF",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"1F",X"FF",
		X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"11",X"1F",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"11",X"1F",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",
		X"30",X"00",X"00",X"11",X"11",X"11",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"33",X"30",X"01",
		X"11",X"11",X"11",X"11",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"03",X"33",X"11",X"BB",X"B1",X"B1",
		X"11",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"03",X"33",X"3B",X"BB",X"B1",X"BB",X"11",X"FF",X"FF",
		X"FF",X"00",X"00",X"00",X"13",X"33",X"3B",X"BB",X"BB",X"4B",X"B1",X"1F",X"FF",X"FF",X"00",X"00",
		X"01",X"11",X"44",X"44",X"BB",X"B4",X"4B",X"B1",X"1F",X"FF",X"FF",X"00",X"00",X"01",X"11",X"B4",
		X"44",X"BB",X"44",X"44",X"4B",X"1F",X"FF",X"FF",X"00",X"00",X"11",X"BB",X"B4",X"44",X"44",X"44",
		X"44",X"41",X"1F",X"FF",X"FF",X"00",X"00",X"11",X"BB",X"BB",X"44",X"44",X"4B",X"44",X"11",X"1F",
		X"FF",X"FF",X"00",X"00",X"11",X"BB",X"BB",X"B4",X"44",X"BB",X"B3",X"33",X"33",X"FF",X"FF",X"00",
		X"01",X"11",X"BB",X"BB",X"BB",X"44",X"4B",X"B3",X"B3",X"33",X"3F",X"FF",X"00",X"00",X"11",X"1B",
		X"BB",X"BB",X"44",X"4B",X"BB",X"B1",X"11",X"33",X"FF",X"00",X"00",X"11",X"11",X"34",X"44",X"44",
		X"44",X"BB",X"B1",X"10",X"03",X"FF",X"00",X"00",X"11",X"13",X"34",X"44",X"44",X"4B",X"BB",X"B1",
		X"1F",X"FF",X"FF",X"00",X"00",X"11",X"33",X"34",X"44",X"44",X"BB",X"B1",X"11",X"FF",X"FF",X"FF",
		X"00",X"00",X"33",X"34",X"44",X"BB",X"BB",X"BB",X"B1",X"11",X"FF",X"FF",X"FF",X"00",X"00",X"33",
		X"3B",X"BB",X"BB",X"BB",X"BB",X"11",X"1F",X"FF",X"FF",X"FF",X"00",X"03",X"30",X"1B",X"BB",X"BB",
		X"B1",X"11",X"11",X"1F",X"FF",X"FF",X"FF",X"00",X"33",X"00",X"11",X"1B",X"BB",X"B1",X"11",X"11",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"01",X"11",X"11",X"11",X"11",X"1F",X"FF",X"FF",X"FF",
		X"FF",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"11",X"11",X"11",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"11",
		X"11",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"11",X"11",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"00",X"00",X"00",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"1F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"0A",
		X"A1",X"1A",X"AA",X"11",X"11",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"AA",X"11",X"11",X"1A",X"AA",
		X"AA",X"FF",X"FF",X"FF",X"00",X"00",X"0A",X"AA",X"11",X"11",X"AA",X"A8",X"8A",X"1F",X"FF",X"FF",
		X"00",X"00",X"08",X"A1",X"11",X"AA",X"AA",X"AA",X"8A",X"A1",X"FF",X"FF",X"00",X"00",X"AA",X"AA",
		X"1A",X"A8",X"A1",X"AA",X"AA",X"AA",X"FF",X"FF",X"00",X"00",X"AA",X"AA",X"AA",X"A8",X"A1",X"AA",
		X"11",X"1A",X"FF",X"FF",X"00",X"00",X"A8",X"81",X"11",X"A8",X"A1",X"AA",X"A1",X"1A",X"FF",X"FF",
		X"00",X"00",X"0A",X"AA",X"AA",X"AA",X"AA",X"11",X"A1",X"1A",X"1F",X"FF",X"00",X"00",X"0A",X"AA",
		X"AA",X"11",X"1A",X"11",X"AA",X"AA",X"1F",X"FF",X"00",X"00",X"0A",X"11",X"A1",X"11",X"1A",X"1A",
		X"11",X"AA",X"AA",X"FF",X"00",X"00",X"A1",X"1A",X"A1",X"11",X"AA",X"A1",X"11",X"AA",X"8A",X"FF",
		X"00",X"00",X"A1",X"1A",X"A1",X"11",X"A8",X"AA",X"AA",X"1A",X"8A",X"FF",X"00",X"00",X"A1",X"11",
		X"AA",X"11",X"A8",X"88",X"8A",X"1A",X"AA",X"FF",X"00",X"00",X"AA",X"1A",X"AA",X"11",X"AA",X"A8",
		X"8A",X"11",X"A1",X"FF",X"00",X"00",X"AA",X"1A",X"AA",X"AA",X"11",X"AA",X"AA",X"11",X"1F",X"FF",
		X"00",X"00",X"AA",X"A8",X"AA",X"AA",X"A1",X"1A",X"A1",X"11",X"FF",X"FF",X"00",X"00",X"0A",X"A8",
		X"AA",X"11",X"AA",X"AA",X"A1",X"11",X"FF",X"FF",X"00",X"00",X"00",X"A8",X"AA",X"11",X"A8",X"8A",
		X"A1",X"AA",X"AF",X"FF",X"00",X"00",X"00",X"AA",X"AA",X"11",X"AA",X"AA",X"1A",X"AA",X"FF",X"FF",
		X"00",X"00",X"00",X"1A",X"AA",X"A1",X"1A",X"A1",X"11",X"AF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"1A",X"AA",X"A1",X"11",X"A1",X"1F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"11",X"A8",X"8A",X"AA",
		X"11",X"1F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"AA",X"AA",X"01",X"1F",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"11",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"11",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"01",X"11",X"00",X"AA",X"01",X"1F",X"FF",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"1A",
		X"AA",X"11",X"FF",X"FF",X"00",X"00",X"00",X"00",X"AA",X"AA",X"A1",X"AA",X"AA",X"A1",X"1F",X"FF",
		X"00",X"00",X"00",X"A1",X"11",X"1A",X"11",X"A1",X"11",X"11",X"1F",X"FF",X"00",X"00",X"00",X"A1",
		X"11",X"AA",X"AA",X"11",X"11",X"11",X"AF",X"FF",X"00",X"00",X"00",X"11",X"AA",X"AA",X"AA",X"AA",
		X"A1",X"11",X"AF",X"FF",X"00",X"00",X"0A",X"AA",X"AA",X"AA",X"AA",X"A8",X"89",X"11",X"AF",X"FF",
		X"00",X"00",X"01",X"AA",X"11",X"AA",X"11",X"AA",X"89",X"91",X"AF",X"FF",X"00",X"00",X"AA",X"1A",
		X"11",X"A8",X"A1",X"99",X"99",X"91",X"AA",X"FF",X"00",X"01",X"1A",X"1A",X"1A",X"AA",X"11",X"99",
		X"11",X"11",X"1A",X"FF",X"00",X"11",X"A1",X"11",X"11",X"19",X"11",X"11",X"11",X"11",X"1A",X"AF",
		X"00",X"11",X"A1",X"AA",X"11",X"19",X"9A",X"11",X"11",X"11",X"AA",X"AF",X"00",X"01",X"AA",X"AA",
		X"11",X"1A",X"99",X"A1",X"11",X"11",X"1A",X"AF",X"00",X"01",X"1A",X"AA",X"11",X"1A",X"AA",X"99",
		X"AA",X"11",X"AA",X"1F",X"00",X"0A",X"1A",X"A1",X"11",X"11",X"AA",X"A9",X"AA",X"AA",X"A1",X"1F",
		X"00",X"0A",X"AA",X"A1",X"11",X"19",X"AA",X"AA",X"99",X"AA",X"11",X"1F",X"00",X"01",X"AA",X"99",
		X"11",X"19",X"AA",X"AA",X"99",X"11",X"11",X"AF",X"00",X"00",X"1A",X"A9",X"11",X"AA",X"AA",X"A9",
		X"A9",X"11",X"11",X"AF",X"00",X"00",X"1A",X"A9",X"91",X"AA",X"AA",X"AA",X"91",X"11",X"1A",X"AF",
		X"00",X"00",X"11",X"1A",X"9A",X"AA",X"AA",X"1A",X"91",X"11",X"AA",X"FF",X"00",X"00",X"A1",X"1A",
		X"11",X"AA",X"A1",X"11",X"91",X"11",X"1A",X"FF",X"00",X"00",X"AA",X"1A",X"11",X"1A",X"A1",X"11",
		X"11",X"11",X"AF",X"FF",X"00",X"00",X"0A",X"1A",X"A1",X"1A",X"AA",X"A1",X"11",X"1A",X"AF",X"FF",
		X"00",X"00",X"0A",X"1A",X"A1",X"AA",X"A8",X"8A",X"11",X"AA",X"AF",X"FF",X"00",X"00",X"0A",X"11",
		X"AA",X"AA",X"A8",X"AA",X"11",X"1A",X"AF",X"FF",X"00",X"00",X"00",X"A1",X"1A",X"AA",X"AA",X"A1",
		X"11",X"1A",X"FF",X"FF",X"00",X"00",X"00",X"AA",X"11",X"AA",X"AA",X"11",X"10",X"AA",X"FF",X"FF",
		X"00",X"00",X"00",X"01",X"11",X"AA",X"11",X"A1",X"0A",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"11",X"AA",X"11",X"11",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"AA",X"A0",X"11",X"11",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"11",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"1F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"1F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"11",X"FF",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"AA",X"AF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"11",X"AF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"00",X"00",
		X"00",X"11",X"00",X"AA",X"01",X"1F",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"10",X"00",X"11",
		X"11",X"1A",X"AA",X"11",X"11",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"0A",X"11",X"AA",X"AA",X"A1",
		X"AA",X"AA",X"A1",X"11",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"AA",X"11",X"11",X"1A",X"11",X"A1",
		X"AA",X"A1",X"1A",X"AF",X"FF",X"FF",X"FF",X"00",X"00",X"0A",X"A1",X"11",X"AA",X"AA",X"11",X"AA",
		X"A1",X"1A",X"AA",X"AF",X"FF",X"FF",X"00",X"00",X"AA",X"11",X"AA",X"AA",X"AA",X"11",X"11",X"11",
		X"1A",X"8A",X"AF",X"FF",X"FF",X"00",X"0A",X"11",X"1A",X"AA",X"AA",X"1A",X"11",X"11",X"11",X"AA",
		X"A1",X"AA",X"AA",X"FF",X"00",X"AA",X"11",X"1A",X"99",X"9A",X"A1",X"11",X"11",X"9A",X"AA",X"1A",
		X"AA",X"AA",X"FF",X"00",X"01",X"1A",X"1A",X"99",X"9A",X"91",X"1A",X"1A",X"AA",X"AA",X"AA",X"AA",
		X"1A",X"1F",X"00",X"11",X"8A",X"1A",X"AA",X"AA",X"11",X"11",X"AA",X"AA",X"AA",X"AA",X"A1",X"11",
		X"AF",X"00",X"11",X"A1",X"1A",X"AA",X"A9",X"11",X"11",X"A1",X"11",X"1A",X"AA",X"11",X"1A",X"AF",
		X"00",X"11",X"11",X"AA",X"AA",X"A9",X"9A",X"11",X"11",X"11",X"11",X"1A",X"11",X"AA",X"FF",X"01",
		X"1A",X"AA",X"AA",X"AA",X"AA",X"99",X"A1",X"A1",X"11",X"11",X"11",X"11",X"AA",X"AF",X"00",X"0A",
		X"1A",X"AA",X"AA",X"AA",X"AA",X"99",X"99",X"A1",X"11",X"11",X"AA",X"AA",X"FF",X"00",X"1A",X"A1",
		X"1A",X"AA",X"AA",X"AA",X"A9",X"A9",X"99",X"91",X"1A",X"AA",X"AF",X"FF",X"00",X"AA",X"A1",X"11",
		X"AA",X"A9",X"AA",X"AA",X"99",X"A9",X"A9",X"9A",X"A1",X"FF",X"FF",X"00",X"AA",X"A1",X"11",X"11",
		X"19",X"AA",X"AA",X"1A",X"AA",X"AA",X"AA",X"11",X"AF",X"FF",X"00",X"AA",X"11",X"11",X"11",X"AA",
		X"AA",X"A9",X"1A",X"A1",X"11",X"9A",X"11",X"AF",X"FF",X"00",X"AA",X"AA",X"11",X"11",X"AA",X"AA",
		X"AA",X"11",X"11",X"1A",X"99",X"99",X"AA",X"FF",X"00",X"0A",X"AA",X"11",X"1A",X"AA",X"AA",X"11",
		X"11",X"11",X"AA",X"9A",X"AA",X"AA",X"FF",X"00",X"11",X"1A",X"A1",X"11",X"AA",X"A1",X"11",X"11",
		X"11",X"1A",X"AA",X"AA",X"AA",X"FF",X"00",X"11",X"AA",X"A1",X"11",X"1A",X"AA",X"11",X"11",X"11",
		X"AA",X"A1",X"1A",X"AA",X"AF",X"00",X"11",X"AA",X"A1",X"11",X"11",X"A1",X"11",X"11",X"1A",X"AA",
		X"11",X"1A",X"A0",X"AF",X"00",X"11",X"1A",X"AA",X"11",X"AA",X"A1",X"AA",X"A9",X"AA",X"A1",X"11",
		X"A0",X"00",X"AF",X"00",X"01",X"1A",X"AA",X"AA",X"AA",X"11",X"1A",X"A9",X"99",X"AA",X"AA",X"00",
		X"00",X"1F",X"00",X"0A",X"11",X"AA",X"AA",X"88",X"A1",X"11",X"1A",X"99",X"1F",X"FF",X"FF",X"FF",
		X"FF",X"00",X"0A",X"AA",X"11",X"AA",X"99",X"11",X"11",X"19",X"9A",X"1F",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"AA",X"A1",X"11",X"99",X"91",X"11",X"11",X"91",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"00",X"0A",X"11",X"11",X"A9",X"9A",X"19",X"AA",X"10",X"1F",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"0A",X"11",X"1A",X"AA",X"99",X"99",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",
		X"A1",X"11",X"AA",X"AA",X"99",X"AF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"0A",
		X"AA",X"AA",X"0A",X"AA",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0A",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"A0",X"00",X"00",X"0A",X"AA",X"00",X"00",
		X"00",X"AF",X"FF",X"FF",X"FF",X"00",X"00",X"0A",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"AF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",
		X"0A",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"0A",X"AA",X"A0",X"AA",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"0A",X"AA",X"10",X"0A",X"AF",X"FF",X"FF",
		X"FF",X"00",X"0A",X"AA",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"AA",X"10",X"01",X"0A",X"00",X"A0",X"AA",X"A0",X"1A",X"AF",X"FF",X"FF",X"FF",X"00",
		X"00",X"0A",X"A0",X"00",X"AA",X"AA",X"00",X"AA",X"A1",X"1A",X"AA",X"AF",X"FF",X"FF",X"00",X"00",
		X"AA",X"00",X"AA",X"AA",X"00",X"00",X"01",X"01",X"1A",X"AA",X"AF",X"FF",X"FF",X"00",X"0A",X"10",
		X"0A",X"AA",X"AA",X"1A",X"00",X"00",X"00",X"AA",X"00",X"A0",X"0A",X"FF",X"00",X"AA",X"00",X"0A",
		X"99",X"9A",X"A1",X"10",X"00",X"00",X"00",X"1A",X"A0",X"0A",X"FF",X"00",X"00",X"0A",X"0A",X"99",
		X"91",X"11",X"1A",X"00",X"00",X"00",X"00",X"AA",X"FF",X"FF",X"00",X"00",X"00",X"0A",X"A1",X"10",
		X"10",X"10",X"00",X"00",X"A0",X"00",X"AA",X"00",X"AF",X"00",X"00",X"00",X"1A",X"11",X"00",X"00",
		X"11",X"00",X"00",X"00",X"00",X"11",X"00",X"AF",X"00",X"00",X"01",X"11",X"10",X"00",X"00",X"01",
		X"11",X"10",X"00",X"00",X"11",X"AF",X"FF",X"01",X"1A",X"A1",X"10",X"AA",X"00",X"00",X"00",X"00",
		X"01",X"11",X"10",X"11",X"AA",X"AF",X"00",X"00",X"01",X"10",X"11",X"00",X"00",X"00",X"00",X"00",
		X"11",X"10",X"AA",X"AF",X"FF",X"00",X"1A",X"A1",X"1A",X"01",X"10",X"00",X"00",X"00",X"00",X"91",
		X"10",X"AA",X"FF",X"FF",X"00",X"AA",X"00",X"00",X"A1",X"10",X"00",X"00",X"00",X"00",X"00",X"90",
		X"A1",X"FF",X"FF",X"00",X"AA",X"11",X"10",X"01",X"10",X"10",X"00",X"00",X"00",X"A0",X"A0",X"10",
		X"AF",X"FF",X"00",X"AA",X"01",X"10",X"00",X"11",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"AF",
		X"FF",X"00",X"AA",X"A0",X"11",X"00",X"11",X"10",X"00",X"00",X"01",X"10",X"09",X"00",X"AA",X"FF",
		X"0A",X"0A",X"A0",X"10",X"0A",X"01",X"11",X"01",X"11",X"01",X"AA",X"11",X"AA",X"AA",X"FF",X"0A",
		X"00",X"1A",X"A0",X"00",X"A0",X"01",X"11",X"11",X"00",X"0A",X"11",X"10",X"AA",X"FF",X"0A",X"00",
		X"AA",X"01",X"11",X"0A",X"00",X"11",X"00",X"00",X"AA",X"11",X"0A",X"AA",X"AF",X"00",X"00",X"AA",
		X"A1",X"01",X"11",X"10",X"00",X"10",X"10",X"01",X"11",X"10",X"00",X"AF",X"00",X"A0",X"00",X"AA",
		X"10",X"A1",X"10",X"AA",X"A9",X"AA",X"01",X"11",X"10",X"00",X"AF",X"0A",X"A0",X"0A",X"AA",X"AA",
		X"AA",X"10",X"0A",X"A1",X"11",X"11",X"11",X"00",X"00",X"AF",X"0A",X"AA",X"00",X"00",X"11",X"11",
		X"00",X"00",X"0A",X"91",X"11",X"10",X"00",X"0A",X"AF",X"00",X"AA",X"0A",X"AA",X"00",X"01",X"11",
		X"11",X"09",X"90",X"00",X"00",X"00",X"AA",X"AF",X"00",X"00",X"00",X"A0",X"0A",X"A0",X"90",X"AA",
		X"A0",X"00",X"00",X"00",X"0A",X"AF",X"FF",X"00",X"0A",X"AA",X"00",X"0A",X"A0",X"00",X"AA",X"AA",
		X"AF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"AA",X"00",X"00",X"00",X"00",X"0A",X"A0",X"00",
		X"00",X"00",X"0A",X"FF",X"FF",X"00",X"00",X"0A",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"AF",X"FF",X"FF",X"00",X"00",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"00",X"AF",X"FF",
		X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"00",X"A0",X"AA",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"0A",X"AF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"A0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0A",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",
		X"00",X"00",X"00",X"AF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"0A",X"00",X"00",X"00",X"A0",X"00",X"AF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"AF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"FF",X"FF",X"FF",X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"FF",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"FF",X"FF",X"FF",
		X"FF",X"A0",X"00",X"A0",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"FF",X"A0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"AF",X"A0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AF",X"FF",X"FF",X"A0",X"0A",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"FF",X"FF",X"FF",X"FF",X"00",X"A0",X"00",X"00",
		X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AF",X"FF",X"FF",X"00",X"A0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"AA",X"AF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"09",X"AA",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0A",X"AA",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0A",X"AF",X"FF",X"FF",X"0A",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"AF",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",
		X"00",X"00",X"00",X"AF",X"00",X"00",X"0A",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"AF",X"00",X"00",X"0A",X"00",X"A0",X"00",X"00",X"0A",X"09",X"99",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"AF",
		X"FF",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FA",X"FF",X"FF",X"FF",
		X"00",X"00",X"AA",X"AF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"00",X"0A",X"00",X"00",X"A9",X"00",X"00",X"00",X"00",X"0A",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"0A",X"00",X"00",X"00",X"00",X"00",X"AF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"AF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"0A",X"AA",X"0A",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"AF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"00",X"00",X"09",X"07",X"70",X"AF",X"FF",X"FF",X"FF",X"00",X"03",X"9A",X"87",X"78",X"DD",
		X"AF",X"FF",X"FF",X"00",X"39",X"A9",X"18",X"81",X"9D",X"EA",X"FF",X"FF",X"03",X"9A",X"99",X"81",
		X"18",X"99",X"DE",X"AF",X"FF",X"39",X"9A",X"99",X"98",X"89",X"99",X"DE",X"EA",X"FF",X"99",X"99",
		X"A9",X"99",X"A9",X"9E",X"ED",X"DD",X"FF",X"99",X"99",X"99",X"AA",X"EE",X"ED",X"DD",X"D9",X"FF",
		X"99",X"88",X"99",X"99",X"ED",X"DD",X"88",X"98",X"FF",X"08",X"22",X"48",X"82",X"42",X"84",X"42",
		X"9F",X"FF",X"00",X"A8",X"98",X"98",X"A8",X"98",X"98",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"09",
		X"05",X"50",X"AF",X"FF",X"FF",X"FF",X"00",X"03",X"9A",X"85",X"58",X"DD",X"AF",X"FF",X"FF",X"00",
		X"39",X"A9",X"78",X"87",X"9D",X"EA",X"FF",X"FF",X"03",X"9A",X"99",X"87",X"78",X"99",X"DE",X"AF",
		X"FF",X"39",X"9A",X"99",X"98",X"89",X"99",X"DE",X"EA",X"FF",X"99",X"99",X"A9",X"99",X"A9",X"9E",
		X"ED",X"DD",X"FF",X"99",X"99",X"99",X"AA",X"EE",X"ED",X"DD",X"D9",X"FF",X"89",X"88",X"99",X"99",
		X"ED",X"DD",X"88",X"99",X"FF",X"09",X"42",X"48",X"82",X"44",X"82",X"24",X"8F",X"FF",X"00",X"89",
		X"8A",X"89",X"89",X"8A",X"89",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"09",X"0B",X"B0",X"AF",X"FF",
		X"FF",X"FF",X"00",X"03",X"9A",X"8B",X"B8",X"DD",X"AF",X"FF",X"FF",X"00",X"39",X"A9",X"B8",X"8B",
		X"9D",X"EA",X"FF",X"FF",X"03",X"9A",X"99",X"8B",X"B8",X"99",X"DE",X"AF",X"FF",X"39",X"9A",X"99",
		X"98",X"89",X"99",X"DE",X"EA",X"FF",X"99",X"99",X"A9",X"99",X"A9",X"9E",X"ED",X"DD",X"FF",X"99",
		X"99",X"99",X"AA",X"EE",X"ED",X"DD",X"D9",X"FF",X"99",X"88",X"99",X"99",X"ED",X"DD",X"88",X"A8",
		X"FF",X"08",X"22",X"84",X"48",X"24",X"84",X"22",X"9F",X"FF",X"00",X"98",X"98",X"98",X"98",X"A8",
		X"98",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"09",X"05",X"50",X"AF",X"FF",X"FF",X"FF",X"00",X"03",
		X"9A",X"85",X"58",X"DD",X"AF",X"FF",X"FF",X"00",X"39",X"A9",X"C8",X"8C",X"9D",X"EA",X"FF",X"FF",
		X"03",X"9A",X"99",X"8C",X"C8",X"99",X"DE",X"AF",X"FF",X"39",X"9A",X"99",X"98",X"89",X"99",X"DE",
		X"EA",X"FF",X"99",X"99",X"A9",X"99",X"A9",X"9E",X"ED",X"DD",X"FF",X"99",X"99",X"99",X"AA",X"EE",
		X"ED",X"DD",X"D8",X"FF",X"89",X"88",X"99",X"99",X"ED",X"DD",X"88",X"99",X"FF",X"09",X"44",X"82",
		X"48",X"24",X"82",X"33",X"8F",X"FF",X"00",X"89",X"89",X"89",X"89",X"89",X"89",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"00",X"00",X"00",X"AB",X"AF",X"FF",X"00",X"00",X"00",X"AB",X"DD",X"DD",X"FF",X"00",X"00",X"AB",
		X"EE",X"EE",X"96",X"FF",X"00",X"AB",X"CE",X"EE",X"CA",X"C6",X"FF",X"AA",X"AA",X"11",X"DB",X"A7",
		X"77",X"FF",X"88",X"89",X"41",X"AA",X"A9",X"88",X"FF",X"00",X"88",X"89",X"99",X"AA",X"86",X"FF",
		X"00",X"00",X"88",X"99",X"9A",X"86",X"FF",X"00",X"00",X"00",X"88",X"99",X"AC",X"FF",X"00",X"00",
		X"00",X"00",X"88",X"AF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"E7",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"DC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"EF",X"FF",X"FF",X"FF",X"00",X"00",X"0D",X"0C",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"76",X"CF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"6C",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"0C",X"CE",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"0C",X"00",
		X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"C0",X"00",X"0D",
		X"00",X"CF",X"FF",X"FF",X"00",X"00",X"0D",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"0D",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"0D",X"0D",
		X"FF",X"FF",X"FF",X"FF",X"00",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"C0",X"00",
		X"CF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"0E",X"FF",X"FF",X"00",X"00",X"07",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"9F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"AF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"50",X"0B",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"AF",X"FF",X"00",X"5F",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"09",X"00",
		X"00",X"5F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"BB",X"DF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"AB",X"BB",X"DF",X"FF",X"00",X"0B",X"BA",X"00",X"00",X"99",
		X"AA",X"AA",X"AD",X"FF",X"00",X"B0",X"0A",X"AA",X"AA",X"BB",X"BB",X"BB",X"BB",X"FF",X"BA",X"BA",
		X"AA",X"DD",X"DD",X"EE",X"EE",X"C7",X"77",X"FF",X"88",X"88",X"88",X"99",X"99",X"99",X"99",X"9A",
		X"AA",X"FF",X"00",X"90",X"03",X"33",X"33",X"33",X"33",X"33",X"38",X"FF",X"00",X"09",X"93",X"00",
		X"00",X"88",X"99",X"99",X"9A",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"89",X"99",X"AF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"99",X"AF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"0C",X"33",X"EB",X"FF",X"FF",
		X"00",X"BC",X"31",X"EB",X"BF",X"FF",X"0A",X"BB",X"31",X"EB",X"BD",X"FF",X"9A",X"BB",X"AA",X"7B",
		X"CC",X"7F",X"AA",X"AB",X"31",X"67",X"CC",X"CF",X"BC",X"C4",X"53",X"16",X"7E",X"EF",X"16",X"A5",
		X"44",X"36",X"A1",X"3F",X"22",X"A4",X"54",X"26",X"A8",X"8F",X"AA",X"A5",X"45",X"16",X"BB",X"BF",
		X"88",X"9A",X"42",X"6B",X"BB",X"AF",X"89",X"9A",X"AA",X"AB",X"BB",X"AF",X"09",X"9A",X"26",X"BA",
		X"BA",X"FF",X"00",X"9A",X"31",X"BA",X"AF",X"FF",X"00",X"0A",X"31",X"BA",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"0A",X"31",X"99",X"FF",X"FF",X"00",X"9A",X"32",X"9B",X"AF",X"FF",X"09",X"94",X"53",X"18",
		X"AA",X"FF",X"92",X"A4",X"45",X"26",X"A8",X"BF",X"36",X"A4",X"54",X"26",X"A1",X"3F",X"1C",X"A4",
		X"52",X"11",X"EC",X"3F",X"CA",X"AB",X"31",X"17",X"CB",X"CF",X"AA",X"BB",X"AA",X"7B",X"CC",X"BF",
		X"AB",X"BB",X"31",X"EB",X"CC",X"CF",X"0B",X"BB",X"31",X"EB",X"B7",X"FF",X"00",X"DC",X"31",X"EB",
		X"EF",X"FF",X"00",X"0D",X"33",X"DE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"08",X"26",X"89",X"FF",X"FF",X"00",X"94",X"54",X"66",X"9F",X"FF",X"09",X"25",X"44",X"16",
		X"A9",X"FF",X"92",X"C4",X"52",X"6B",X"C1",X"9F",X"2C",X"AC",X"AA",X"EE",X"BC",X"2F",X"AA",X"BA",
		X"31",X"7B",X"CC",X"CF",X"AB",X"BB",X"21",X"EB",X"BC",X"CF",X"0D",X"BB",X"21",X"EB",X"BD",X"FF",
		X"00",X"DC",X"23",X"EB",X"7F",X"FF",X"00",X"0D",X"DD",X"DD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"0A",X"21",X"29",X"FF",X"FF",X"00",X"A4",X"54",X"16",
		X"9F",X"FF",X"0A",X"AA",X"42",X"6B",X"B9",X"FF",X"AA",X"BB",X"BB",X"CC",X"CB",X"9F",X"CB",X"BB",
		X"41",X"EB",X"CC",X"CF",X"CC",X"BB",X"31",X"7B",X"BD",X"DF",X"0C",X"CB",X"33",X"EB",X"ED",X"FF",
		X"00",X"CE",X"EE",X"E7",X"EF",X"FF",X"00",X"0D",X"DD",X"D7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"08",X"21",X"1B",
		X"FF",X"FF",X"00",X"AB",X"AA",X"AC",X"CF",X"FF",X"0A",X"AB",X"26",X"EB",X"CC",X"FF",X"BA",X"BB",
		X"26",X"EB",X"BC",X"CF",X"DD",X"AB",X"26",X"EB",X"BE",X"EF",X"0E",X"DE",X"EE",X"EE",X"7E",X"FF",
		X"00",X"DD",X"DD",X"DD",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"0A",X"98",X"EB",
		X"FF",X"FF",X"00",X"AB",X"33",X"EB",X"BF",X"FF",X"09",X"9A",X"26",X"EB",X"BB",X"FF",X"CC",X"CE",
		X"EE",X"EE",X"77",X"EF",X"CC",X"CD",X"DD",X"DD",X"DE",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"07",X"55",X"FF",X"FF",X"77",X"55",X"5F",X"FF",
		X"0A",X"AA",X"FF",X"FF",X"99",X"99",X"9F",X"FF",X"EE",X"98",X"49",X"FF",X"AA",X"99",X"49",X"FF",
		X"7A",X"99",X"89",X"FF",X"99",X"99",X"9F",X"FF",X"07",X"77",X"FF",X"FF",X"DC",X"CC",X"6F",X"FF",
		X"0D",X"CC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"07",X"55",X"FF",X"FF",
		X"75",X"55",X"7F",X"FF",X"0A",X"AA",X"FF",X"FF",X"99",X"99",X"9F",X"FF",X"AA",X"98",X"49",X"FF",
		X"EE",X"99",X"49",X"FF",X"7A",X"99",X"89",X"FF",X"99",X"99",X"9F",X"FF",X"07",X"77",X"FF",X"FF",
		X"CC",X"C6",X"6F",X"FF",X"0C",X"C6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"05",X"57",X"FF",X"FF",X"55",X"77",X"AF",X"FF",X"0A",X"AA",X"FF",X"FF",X"99",X"99",X"9F",X"FF",
		X"AA",X"98",X"49",X"FF",X"AA",X"99",X"49",X"FF",X"EE",X"99",X"89",X"FF",X"99",X"99",X"9F",X"FF",
		X"07",X"77",X"FF",X"FF",X"C6",X"66",X"5F",X"FF",X"0C",X"66",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"05",X"7A",X"FF",X"FF",X"57",X"77",X"AF",X"FF",X"0A",X"AA",X"FF",X"FF",
		X"99",X"99",X"9F",X"FF",X"AA",X"98",X"49",X"FF",X"EE",X"99",X"49",X"FF",X"22",X"99",X"89",X"FF",
		X"99",X"99",X"9F",X"FF",X"07",X"77",X"FF",X"FF",X"66",X"65",X"5F",X"FF",X"06",X"55",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0A",X"7C",X"FF",X"FF",X"A7",X"7C",X"BF",X"FF",
		X"0A",X"AA",X"FF",X"FF",X"99",X"99",X"9F",X"FF",X"EE",X"98",X"49",X"FF",X"22",X"99",X"49",X"FF",
		X"AA",X"99",X"89",X"FF",X"99",X"99",X"9F",X"FF",X"07",X"77",X"FF",X"FF",X"65",X"55",X"DF",X"FF",
		X"05",X"5D",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"07",X"CB",X"FF",X"FF",
		X"7C",X"CB",X"5F",X"FF",X"0A",X"AA",X"FF",X"FF",X"99",X"99",X"9F",X"FF",X"22",X"98",X"49",X"FF",
		X"AA",X"99",X"49",X"FF",X"AA",X"99",X"89",X"FF",X"99",X"99",X"9F",X"FF",X"07",X"77",X"FF",X"FF",
		X"55",X"DD",X"DF",X"FF",X"05",X"DD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"07",X"B5",X"FF",X"FF",X"77",X"7B",X"5F",X"FF",X"0A",X"AA",X"FF",X"FF",X"99",X"99",X"9F",X"FF",
		X"77",X"98",X"49",X"FF",X"AA",X"99",X"49",X"FF",X"AA",X"99",X"89",X"FF",X"99",X"99",X"9F",X"FF",
		X"07",X"77",X"FF",X"FF",X"5D",X"DC",X"CF",X"FF",X"0D",X"CC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"07",X"75",X"FF",X"FF",X"C7",X"75",X"5F",X"FF",X"0A",X"AA",X"FF",X"FF",
		X"99",X"99",X"9F",X"FF",X"AA",X"98",X"49",X"FF",X"AA",X"99",X"49",X"FF",X"AA",X"99",X"89",X"FF",
		X"99",X"99",X"9F",X"FF",X"07",X"77",X"FF",X"FF",X"DD",X"CC",X"CF",X"FF",X"0D",X"CC",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"03",X"22",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"03",X"33",X"33",X"33",X"00",X"01",X"1F",
		X"FF",X"FF",X"03",X"33",X"22",X"22",X"11",X"10",X"AA",X"AA",X"FF",X"FF",X"A3",X"32",X"2D",X"44",
		X"44",X"3A",X"A2",X"2A",X"AF",X"FF",X"CC",X"A3",X"3D",X"66",X"99",X"CD",X"D3",X"3D",X"CF",X"FF",
		X"0C",X"CC",X"CC",X"CC",X"CC",X"C0",X"CD",X"DC",X"FF",X"FF",X"00",X"0D",X"DD",X"DD",X"DD",X"00",
		X"0A",X"AF",X"FF",X"FF",X"00",X"00",X"0C",X"CC",X"CF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"03",X"22",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"03",X"33",X"33",
		X"33",X"00",X"0A",X"AF",X"FF",X"FF",X"03",X"33",X"22",X"22",X"11",X"10",X"A2",X"2A",X"FF",X"FF",
		X"A3",X"32",X"2D",X"44",X"44",X"3D",X"D2",X"2D",X"AF",X"FF",X"CC",X"A3",X"3D",X"66",X"99",X"CD",
		X"DD",X"DD",X"CF",X"FF",X"0C",X"CC",X"CC",X"CC",X"CC",X"C0",X"DA",X"AD",X"FF",X"FF",X"00",X"0D",
		X"DD",X"DD",X"DD",X"00",X"0A",X"AF",X"FF",X"FF",X"00",X"00",X"0C",X"CC",X"CF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"03",X"22",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"03",X"33",X"33",X"33",X"00",X"02",X"2F",X"FF",X"FF",X"03",X"33",X"22",X"22",X"11",X"10",
		X"D2",X"2D",X"FF",X"FF",X"A3",X"32",X"2E",X"44",X"44",X"3D",X"DD",X"DD",X"AF",X"FF",X"CC",X"A3",
		X"3E",X"66",X"99",X"CD",X"DA",X"AD",X"CF",X"FF",X"0C",X"CC",X"CC",X"CC",X"CC",X"C0",X"DA",X"AD",
		X"FF",X"FF",X"00",X"0D",X"DD",X"DD",X"DD",X"00",X"0D",X"DF",X"FF",X"FF",X"00",X"00",X"0C",X"CC",
		X"CF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"03",X"22",X"1F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"03",X"33",X"33",X"33",X"00",X"02",X"2F",X"FF",X"FF",X"03",X"33",
		X"22",X"22",X"11",X"10",X"DD",X"DD",X"FF",X"FF",X"A3",X"32",X"2E",X"44",X"44",X"3D",X"DA",X"AD",
		X"AF",X"FF",X"CC",X"A3",X"3E",X"66",X"99",X"CD",X"DA",X"AD",X"7F",X"FF",X"0C",X"CC",X"CC",X"CC",
		X"CC",X"C0",X"77",X"77",X"FF",X"FF",X"00",X"0D",X"DD",X"DD",X"DD",X"00",X"03",X"3F",X"FF",X"FF",
		X"00",X"00",X"0C",X"CC",X"CF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"03",X"22",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"03",X"33",X"33",X"33",X"00",X"0C",X"CF",
		X"FF",X"FF",X"03",X"33",X"22",X"22",X"11",X"10",X"CA",X"AC",X"FF",X"FF",X"A3",X"32",X"2E",X"44",
		X"44",X"3D",X"DA",X"AD",X"AF",X"FF",X"CC",X"A3",X"3E",X"66",X"99",X"C7",X"77",X"77",X"7F",X"FF",
		X"0C",X"CC",X"CC",X"CC",X"CC",X"C0",X"72",X"27",X"FF",X"FF",X"00",X"0D",X"DD",X"DD",X"DD",X"00",
		X"03",X"3F",X"FF",X"FF",X"00",X"00",X"0C",X"CC",X"CF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"11",X"11",
		X"FF",X"FF",X"01",X"77",X"77",X"1F",X"FF",X"17",X"71",X"17",X"71",X"FF",X"17",X"11",X"11",X"71",
		X"FF",X"17",X"11",X"11",X"71",X"FF",X"17",X"71",X"17",X"71",X"FF",X"01",X"77",X"77",X"1F",X"FF",
		X"00",X"11",X"11",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"11",X"11",X"FF",X"FF",X"01",X"11",X"11",X"1F",X"FF",X"11",X"17",X"71",X"11",X"FF",X"11",X"71",
		X"17",X"11",X"FF",X"11",X"71",X"17",X"11",X"FF",X"11",X"17",X"71",X"11",X"FF",X"01",X"11",X"11",
		X"1F",X"FF",X"00",X"11",X"11",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"00",X"77",X"77",X"FF",X"FF",X"07",X"88",X"88",X"7F",X"FF",X"78",X"89",X"98",X"87",X"FF",
		X"78",X"9A",X"A9",X"87",X"FF",X"78",X"9A",X"A9",X"87",X"FF",X"78",X"89",X"98",X"87",X"FF",X"07",
		X"88",X"88",X"7F",X"FF",X"00",X"77",X"77",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"00",X"88",X"88",X"FF",X"FF",X"08",X"99",X"99",X"8F",X"FF",X"89",X"9A",X"A9",
		X"98",X"FF",X"89",X"AB",X"BA",X"98",X"FF",X"89",X"AB",X"BA",X"98",X"FF",X"89",X"9A",X"A9",X"98",
		X"FF",X"08",X"99",X"99",X"8F",X"FF",X"00",X"88",X"88",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"88",X"88",X"FF",X"FF",X"08",X"99",X"99",X"8F",X"FF",X"89",
		X"9B",X"B9",X"98",X"FF",X"89",X"BD",X"DB",X"98",X"FF",X"89",X"BD",X"DB",X"98",X"FF",X"89",X"9B",
		X"B9",X"98",X"FF",X"08",X"99",X"99",X"8F",X"FF",X"00",X"88",X"88",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"88",X"88",X"FF",X"FF",X"08",X"AA",X"AA",X"8F",
		X"FF",X"8A",X"AC",X"CA",X"A8",X"FF",X"8A",X"CE",X"EC",X"A8",X"FF",X"8A",X"CE",X"EC",X"A8",X"FF",
		X"8A",X"AC",X"CA",X"A8",X"FF",X"08",X"AA",X"AA",X"8F",X"FF",X"00",X"88",X"88",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"99",X"99",X"FF",X"FF",X"09",X"CC",
		X"CC",X"9F",X"FF",X"9C",X"CD",X"DC",X"C9",X"FF",X"9C",X"DE",X"ED",X"C9",X"FF",X"9C",X"DE",X"ED",
		X"C9",X"FF",X"9C",X"CD",X"DC",X"C9",X"FF",X"09",X"CC",X"CC",X"9F",X"FF",X"00",X"99",X"99",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"02",
		X"11",X"FF",X"FF",X"FF",X"00",X"02",X"23",X"33",X"12",X"FF",X"FF",X"02",X"22",X"3E",X"EE",X"E1",
		X"2F",X"FF",X"22",X"23",X"EE",X"55",X"EE",X"11",X"FF",X"AA",X"AE",X"E9",X"55",X"5E",X"EA",X"FF",
		X"0C",X"AE",X"99",X"EE",X"66",X"E3",X"FF",X"0C",X"AE",X"99",X"EE",X"66",X"E3",X"FF",X"22",X"3E",
		X"E8",X"88",X"6E",X"E1",X"FF",X"77",X"77",X"EE",X"88",X"EE",X"CC",X"FF",X"0C",X"CD",X"7E",X"EE",
		X"ED",X"7F",X"FF",X"00",X"0C",X"CD",X"DD",X"CC",X"FF",X"FF",X"00",X"00",X"0C",X"CC",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"66",X"66",
		X"FF",X"FF",X"06",X"77",X"77",X"6F",X"FF",X"67",X"71",X"17",X"76",X"FF",X"67",X"11",X"11",X"76",
		X"FF",X"67",X"11",X"11",X"76",X"FF",X"67",X"71",X"17",X"76",X"FF",X"06",X"77",X"77",X"6F",X"FF",
		X"00",X"66",X"66",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"55",X"55",X"FF",X"FF",X"05",X"11",X"11",X"5F",X"FF",X"51",X"17",X"71",X"15",X"FF",X"51",X"71",
		X"17",X"15",X"FF",X"51",X"71",X"17",X"15",X"FF",X"51",X"17",X"71",X"15",X"FF",X"05",X"11",X"11",
		X"5F",X"FF",X"00",X"55",X"55",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"00",X"77",X"77",X"FF",X"FF",X"07",X"88",X"88",X"7F",X"FF",X"78",X"89",X"98",X"87",X"FF",
		X"78",X"9A",X"A9",X"87",X"FF",X"78",X"9A",X"A9",X"87",X"FF",X"78",X"89",X"98",X"87",X"FF",X"07",
		X"88",X"88",X"7F",X"FF",X"00",X"77",X"77",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"00",X"66",X"66",X"FF",X"FF",X"06",X"99",X"99",X"6F",X"FF",X"69",X"9A",X"A9",
		X"96",X"FF",X"69",X"AB",X"BA",X"96",X"FF",X"69",X"AB",X"BA",X"96",X"FF",X"69",X"9A",X"A9",X"96",
		X"FF",X"06",X"99",X"99",X"6F",X"FF",X"00",X"66",X"66",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"55",X"55",X"FF",X"FF",X"05",X"99",X"99",X"5F",X"FF",X"59",
		X"9B",X"B9",X"95",X"FF",X"59",X"BD",X"DB",X"95",X"FF",X"59",X"BD",X"DB",X"95",X"FF",X"59",X"9B",
		X"B9",X"95",X"FF",X"05",X"99",X"99",X"5F",X"FF",X"00",X"55",X"55",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"77",X"77",X"FF",X"FF",X"07",X"AA",X"AA",X"7F",
		X"FF",X"7A",X"AC",X"CA",X"A7",X"FF",X"7A",X"CE",X"EC",X"A7",X"FF",X"7A",X"CE",X"EC",X"A7",X"FF",
		X"7A",X"AC",X"CA",X"A7",X"FF",X"07",X"AA",X"AA",X"7F",X"FF",X"00",X"77",X"77",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"66",X"66",X"FF",X"FF",X"06",X"CC",
		X"CC",X"6F",X"FF",X"6C",X"CD",X"DC",X"C6",X"FF",X"6C",X"DE",X"ED",X"C6",X"FF",X"6C",X"DE",X"ED",
		X"C6",X"FF",X"6C",X"CD",X"DC",X"C6",X"FF",X"06",X"CC",X"CC",X"6F",X"FF",X"00",X"66",X"66",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"FF",X"1E",X"1F",X"01",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"CC",X"0C",X"CF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"0C",X"CC",X"C2",X"CC",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"0C",
		X"2C",X"22",X"2C",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"C2",X"2C",X"22",X"CC",X"CF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"0C",X"22",X"CC",X"C2",X"2C",X"2C",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"0C",X"CC",X"C2",X"CC",X"C2",X"2C",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"0C",X"22",
		X"C2",X"2C",X"C2",X"2C",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"0C",X"22",X"CC",X"2C",X"CC",X"CC",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"C2",X"2C",X"CC",X"2C",X"CF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"C2",X"CC",X"22",X"2C",X"CF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"0C",
		X"CC",X"C2",X"CC",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"CC",X"0C",X"CF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",X"00",X"04",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"E0",X"00",X"CF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"C0",X"00",X"C0",X"00",X"00",X"CC",X"EF",X"FF",X"FF",X"FF",X"00",X"00",X"CC",X"12",
		X"CC",X"21",X"2C",X"CF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"0C",X"C1",X"22",X"11",X"12",X"2F",
		X"FF",X"FF",X"FF",X"FF",X"00",X"04",X"22",X"22",X"11",X"11",X"C1",X"2F",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"02",X"11",X"11",X"11",X"CC",X"2F",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"11",
		X"11",X"1C",X"C1",X"1F",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"11",X"11",X"12",X"C1",X"2C",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"21",X"11",X"CC",X"11",X"CF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"22",X"1C",X"C1",X"22",X"CC",X"CE",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"C2",
		X"12",X"12",X"12",X"2F",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"0C",X"CC",X"11",X"12",X"22",X"CF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"CC",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"0E",X"00",X"E0",X"EF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"0E",X"00",X"0C",X"00",X"C0",X"00",X"E0",X"0E",X"FF",X"FF",X"FF",
		X"00",X"00",X"C0",X"0C",X"0C",X"C0",X"C0",X"C0",X"CF",X"FF",X"FF",X"FF",X"00",X"00",X"0C",X"CC",
		X"4D",X"C0",X"CC",X"CC",X"FF",X"FF",X"FF",X"FF",X"00",X"0E",X"CC",X"C2",X"DD",X"DD",X"D1",X"CC",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"04",X"D2",X"D2",X"11",X"1C",X"CC",X"FF",X"FF",X"FF",X"FF",
		X"00",X"0E",X"CC",X"C1",X"2D",X"1D",X"CD",X"4C",X"CE",X"FF",X"FF",X"FF",X"00",X"00",X"0C",X"DD",
		X"22",X"DD",X"D2",X"1F",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"0C",X"DD",X"CC",X"CC",X"CD",X"2C",
		X"EF",X"FF",X"FF",X"FF",X"00",X"00",X"0C",X"2D",X"EC",X"CD",X"42",X"CF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"0E",X"0C",X"21",X"2C",X"D1",X"1D",X"CC",X"EF",X"FF",X"FF",X"FF",X"00",X"00",X"CC",X"11",
		X"2C",X"CD",X"2D",X"CC",X"FF",X"FF",X"FF",X"FF",X"00",X"EC",X"CC",X"D2",X"CC",X"22",X"42",X"CC",
		X"CE",X"FF",X"FF",X"FF",X"00",X"00",X"0C",X"CC",X"CC",X"CC",X"CC",X"0C",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"C0",X"00",X"C0",X"CC",X"0C",X"C0",X"EF",X"FF",X"FF",X"FF",X"00",X"0E",X"00",X"0E",
		X"00",X"0C",X"00",X"0E",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"EF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"0E",X"00",X"00",X"C0",X"0C",X"00",X"00",X"EF",X"FF",X"FF",X"FF",X"00",X"00",X"CC",X"0D",
		X"C0",X"CC",X"00",X"0C",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"CC",X"DD",X"C2",X"CC",X"C2",X"CC",
		X"FF",X"FF",X"FF",X"FF",X"04",X"00",X"0C",X"DD",X"DC",X"CC",X"CC",X"D2",X"FF",X"FF",X"FF",X"FF",
		X"00",X"CC",X"02",X"2C",X"CC",X"22",X"2C",X"CD",X"CC",X"FF",X"FF",X"FF",X"00",X"0C",X"CC",X"DC",
		X"2C",X"C2",X"22",X"2C",X"DF",X"FF",X"FF",X"FF",X"00",X"00",X"CD",X"DC",X"22",X"C2",X"22",X"CD",
		X"DD",X"2C",X"EF",X"FF",X"00",X"0C",X"DD",X"CC",X"22",X"CC",X"DC",X"22",X"DD",X"CF",X"FF",X"FF",
		X"EC",X"CC",X"CC",X"C2",X"2C",X"22",X"DC",X"22",X"CD",X"CF",X"FF",X"FF",X"00",X"0C",X"2C",X"CC",
		X"DC",X"22",X"DC",X"2C",X"2C",X"CF",X"FF",X"FF",X"00",X"02",X"22",X"DC",X"DC",X"22",X"DD",X"C2",
		X"DC",X"0C",X"FF",X"FF",X"4C",X"CC",X"CC",X"DC",X"2D",X"CC",X"DC",X"CC",X"DD",X"CF",X"FF",X"FF",
		X"00",X"CC",X"2C",X"DD",X"2C",X"DD",X"DC",X"22",X"DD",X"CF",X"FF",X"FF",X"00",X"02",X"22",X"DC",
		X"C2",X"2C",X"CC",X"22",X"2D",X"CF",X"FF",X"FF",X"00",X"CC",X"CC",X"DC",X"22",X"22",X"2C",X"CD",
		X"DD",X"FF",X"FF",X"FF",X"0E",X"00",X"2C",X"DC",X"2C",X"22",X"22",X"CD",X"CC",X"CC",X"FF",X"FF",
		X"00",X"00",X"0C",X"CD",X"CD",X"22",X"22",X"CC",X"C2",X"00",X"EF",X"FF",X"00",X"0C",X"CC",X"2C",
		X"CD",X"CC",X"CC",X"C2",X"CF",X"FF",X"FF",X"FF",X"00",X"0C",X"C2",X"22",X"CC",X"C2",X"DD",X"C2",
		X"CC",X"FF",X"FF",X"FF",X"00",X"0C",X"C0",X"0C",X"CC",X"22",X"DC",X"00",X"0C",X"FF",X"FF",X"FF",
		X"00",X"44",X"00",X"0C",X"00",X"00",X"C0",X"00",X"00",X"EF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"EF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",
		X"6F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"60",X"03",X"33",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"33",X"33",X"33",X"33",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"03",X"CC",
		X"3C",X"CC",X"33",X"33",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"0C",X"CD",X"DD",X"3C",X"CC",X"33",
		X"3F",X"FF",X"FF",X"FF",X"00",X"00",X"CC",X"DD",X"C3",X"C3",X"C3",X"33",X"3F",X"FF",X"FF",X"FF",
		X"00",X"00",X"CC",X"3D",X"DC",X"C3",X"C3",X"33",X"33",X"FF",X"FF",X"FF",X"00",X"00",X"DC",X"CD",
		X"DD",X"CC",X"3C",X"CC",X"33",X"3F",X"FF",X"FF",X"00",X"0C",X"CD",X"DD",X"DC",X"CC",X"CC",X"CC",
		X"33",X"3F",X"FF",X"FF",X"00",X"0C",X"CC",X"DC",X"C3",X"3C",X"CC",X"CC",X"33",X"3F",X"FF",X"FF",
		X"00",X"03",X"CC",X"DC",X"CD",X"33",X"CC",X"C3",X"33",X"3F",X"FF",X"FF",X"00",X"00",X"CD",X"CD",
		X"3D",X"D3",X"CD",X"CC",X"33",X"FF",X"FF",X"FF",X"00",X"00",X"CC",X"DC",X"DC",X"C3",X"DC",X"C3",
		X"33",X"FF",X"FF",X"FF",X"00",X"00",X"CC",X"DD",X"DC",X"CD",X"DD",X"33",X"33",X"FF",X"FF",X"FF",
		X"00",X"00",X"3C",X"CD",X"DC",X"CD",X"D3",X"C3",X"3F",X"FF",X"FF",X"FF",X"00",X"00",X"0C",X"CD",
		X"CD",X"3D",X"3C",X"C3",X"00",X"06",X"FF",X"FF",X"06",X"00",X"00",X"3C",X"CD",X"DC",X"D3",X"33",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"C0",X"33",X"C3",X"33",X"3F",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"0D",X"33",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"06",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"6F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"03",X"33",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"03",X"33",X"C3",X"33",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"03",
		X"33",X"C3",X"33",X"3F",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"33",X"CC",X"33",X"C3",X"3F",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"03",X"3C",X"CC",X"33",X"3C",X"33",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"03",X"33",X"C3",X"33",X"CC",X"33",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"03",X"33",
		X"33",X"C3",X"33",X"33",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"03",X"3C",X"C3",X"CC",X"CC",X"33",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"3C",X"CC",X"33",X"C3",X"33",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"33",X"3C",X"C3",X"33",X"3F",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"03",
		X"33",X"33",X"33",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"03",X"33",X"3F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"6F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"43",X"40",X"4F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"04",X"40",X"44",X"43",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"03",
		X"34",X"30",X"44",X"4F",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"44",X"30",X"43",X"4F",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"04",X"04",X"43",X"30",X"3F",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"04",X"33",X"04",X"03",X"4F",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"30",X"34",X"44",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"04",X"03",X"3F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"AF",X"FF",X"BB",X"DA",X"FF",X"AA",X"AA",X"FF",
		X"AA",X"AF",X"FF",X"AA",X"AA",X"FF",X"BB",X"DA",X"FF",X"AA",X"AF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BB",X"BC",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"9B",X"CC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0C",X"FF",X"FF",X"FF",X"FF",X"99",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"9C",X"CF",
		X"FF",X"FF",X"FF",X"98",X"8C",X"00",X"00",X"00",X"00",X"00",X"09",X"9C",X"CC",X"FF",X"FF",X"FF",
		X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"08",X"8A",X"AA",X"FF",X"FF",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"8A",X"AF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0A",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"9C",X"CF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"09",X"9C",X"CC",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"8A",X"AA",X"00",X"AA",X"AC",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"8A",
		X"A0",X"00",X"9A",X"CC",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"99",
		X"CC",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"98",X"8C",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"FF",X"00",X"00",X"0C",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"9C",X"CF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"09",X"9C",X"CC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"00",X"08",X"8A",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"8A",X"AF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"0A",
		X"00",X"00",X"00",X"00",X"00",X"0A",X"AA",X"CF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"AC",X"CF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",
		X"9C",X"CF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"88",X"CF",X"FF",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"88",X"8F",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"9C",X"CF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"09",X"9C",X"CC",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"08",X"8A",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"8A",
		X"AF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"70",X"70",X"7F",X"70",X"70",X"7F",X"77",X"77",X"7F",X"77",X"77",X"7F",X"FF",
		X"FF",X"FF",X"77",X"77",X"7F",X"70",X"00",X"7F",X"77",X"77",X"7F",X"77",X"77",X"7F",X"FF",X"FF",
		X"FF",X"77",X"77",X"7F",X"70",X"00",X"7F",X"77",X"77",X"7F",X"77",X"77",X"7F",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"70",X"77",X"7F",X"70",X"70",X"7F",X"77",X"70",X"7F",X"77",X"70",X"7F",X"FF",
		X"FF",X"FF",X"77",X"77",X"7F",X"70",X"00",X"7F",X"77",X"77",X"7F",X"77",X"77",X"7F",X"FF",X"FF",
		X"FF",X"77",X"77",X"7F",X"70",X"00",X"7F",X"77",X"77",X"7F",X"77",X"77",X"7F",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"0E",X"FF",X"ED",X"EF",X"ED",X"EF",X"0E",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"3E",X"2E",X"3E",X"2E",X"3E",X"2F",X"3E",X"2E",X"3E",X"2E",X"3E",X"2F",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AF",X"88",X"88",X"88",X"88",X"66",X"FF",X"44",X"44",X"44",X"43",X"EB",X"7F",
		X"55",X"55",X"54",X"44",X"EB",X"7F",X"88",X"88",X"88",X"43",X"ED",X"DF",X"DD",X"DD",X"DD",X"DD",
		X"DD",X"FF",X"EE",X"EE",X"EE",X"EE",X"EE",X"EF",X"3E",X"2E",X"3E",X"2E",X"3E",X"2F",X"3E",X"2E",
		X"3E",X"2E",X"3E",X"2F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"2E",X"3E",X"2E",X"3E",X"2E",X"3F",X"2E",X"3E",X"2E",X"3E",X"2E",X"3F",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AF",X"88",X"88",X"88",X"88",X"66",X"FF",X"44",X"44",X"44",X"43",X"1B",X"7F",X"55",X"55",
		X"54",X"44",X"1B",X"7F",X"88",X"88",X"88",X"43",X"1D",X"DF",X"DD",X"DD",X"DD",X"DD",X"DD",X"FF",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EF",X"2E",X"3E",X"2E",X"3E",X"2E",X"3F",X"2E",X"3E",X"2E",X"3E",
		X"2E",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"06",X"66",X"66",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"77",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"22",
		X"27",X"77",X"77",X"77",X"77",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"02",X"22",X"26",X"66",X"66",
		X"7F",X"FF",X"FF",X"FF",X"00",X"00",X"06",X"62",X"22",X"22",X"27",X"77",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"06",X"22",X"22",X"22",X"26",X"7F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"22",X"22",X"22",X"26",X"7F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"07",X"72",X"22",X"22",X"26",
		X"7F",X"FF",X"FF",X"FF",X"00",X"00",X"06",X"76",X"72",X"22",X"22",X"22",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"08",X"87",X"22",X"22",X"22",X"7F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"78",X"72",X"22",X"22",X"27",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"72",
		X"22",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"06",X"66",X"66",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"02",X"2F",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"02",X"66",X"66",X"6F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"02",X"77",X"77",X"00",X"00",X"00",X"2F",X"FF",X"FF",X"FF",X"00",X"00",X"77",X"77",
		X"77",X"75",X"52",X"22",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"07",X"66",X"66",X"52",X"22",X"2F",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"75",X"52",X"22",X"22",X"25",X"6F",X"FF",X"FF",X"FF",
		X"00",X"00",X"07",X"62",X"22",X"22",X"22",X"5F",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"07",X"52",
		X"22",X"22",X"22",X"2F",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"07",X"52",X"22",X"22",X"25",X"72",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"22",X"22",X"22",X"25",X"67",X"6F",X"FF",X"FF",X"FF",
		X"00",X"00",X"05",X"22",X"22",X"22",X"58",X"82",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"72",X"22",
		X"22",X"55",X"87",X"22",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"02",X"25",X"55",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"20",X"66",X"66",X"6F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"04",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"4F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"04",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"04",X"4F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"44",
		X"4F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"04",X"44",X"4F",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"04",X"44",X"44",X"4F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"44",X"44",X"44",X"4F",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"44",X"44",X"44",X"4F",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"04",X"44",X"44",X"44",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"04",X"44",X"44",X"44",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"44",X"44",X"44",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"04",X"44",X"4F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",
		X"4F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"4F",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"4F",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"04",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"04",X"40",X"4F",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"43",X"43",X"43",X"4F",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"04",X"32",X"44",X"42",X"30",
		X"4F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"03",X"24",X"33",X"34",X"24",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"44",X"43",X"33",X"33",X"44",X"4F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"03",
		X"33",X"33",X"33",X"33",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"43",X"33",X"33",X"33",X"34",
		X"44",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"04",X"23",X"33",X"33",X"24",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"43",X"24",X"33",X"34",X"23",X"4F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"04",
		X"32",X"43",X"42",X"34",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"04",X"44",X"34",X"34",X"04",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"40",X"40",X"44",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"04",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"08",X"88",X"88",X"8F",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"08",X"77",X"77",X"77",X"88",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"87",X"77",X"66",X"66",X"77",X"8F",X"FF",X"FF",X"FF",X"00",X"00",X"07",X"77",
		X"66",X"64",X"46",X"67",X"88",X"FF",X"FF",X"FF",X"00",X"00",X"07",X"76",X"64",X"44",X"44",X"66",
		X"78",X"FF",X"FF",X"FF",X"00",X"00",X"87",X"66",X"44",X"33",X"34",X"46",X"67",X"FF",X"FF",X"FF",
		X"00",X"00",X"87",X"64",X"43",X"33",X"33",X"44",X"67",X"8F",X"FF",X"FF",X"00",X"00",X"87",X"64",
		X"43",X"33",X"33",X"44",X"67",X"8F",X"FF",X"FF",X"00",X"00",X"87",X"64",X"43",X"33",X"33",X"34",
		X"68",X"8F",X"FF",X"FF",X"00",X"00",X"87",X"64",X"44",X"33",X"33",X"44",X"67",X"8F",X"FF",X"FF",
		X"00",X"00",X"87",X"66",X"44",X"33",X"33",X"44",X"67",X"8F",X"FF",X"FF",X"00",X"00",X"88",X"76",
		X"44",X"34",X"44",X"46",X"67",X"8F",X"FF",X"FF",X"00",X"00",X"08",X"76",X"64",X"44",X"66",X"66",
		X"77",X"FF",X"FF",X"FF",X"00",X"00",X"08",X"87",X"66",X"66",X"67",X"77",X"88",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"88",X"77",X"77",X"77",X"78",X"7F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"08",
		X"88",X"78",X"78",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"88",X"8F",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"3F",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"33",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"03",X"33",X"03",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"30",X"00",X"33",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"03",X"30",X"00",X"33",X"3F",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"33",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"33",X"33",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"03",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"02",X"00",X"00",X"00",X"2F",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"02",X"00",
		X"33",X"33",X"2F",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"23",X"33",X"32",X"23",X"00",
		X"02",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"03",X"32",X"00",X"23",X"33",X"2F",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"03",X"20",X"00",X"22",X"33",X"3F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"03",
		X"30",X"00",X"00",X"23",X"3F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"33",X"20",X"00",X"00",X"02",
		X"3F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"33",X"32",X"00",X"00",X"23",X"3F",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"02",X"22",X"00",X"02",X"33",X"3F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"22",
		X"32",X"22",X"33",X"23",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"02",X"20",X"33",X"33",X"23",X"32",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"33",X"23",X"02",X"2F",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"2F",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"2F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"40",X"03",X"33",X"33",X"4F",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"44",
		X"33",X"32",X"33",X"3F",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"03",X"43",X"20",X"23",X"3F",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"33",X"34",X"00",X"02",X"33",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"44",X"42",X"30",X"00",X"04",X"44",X"44",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"33",
		X"20",X"00",X"00",X"02",X"3F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"33",X"20",X"00",X"00",X"03",
		X"3F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"03",X"22",X"40",X"00",X"23",X"3F",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"03",X"34",X"32",X"32",X"33",X"3F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"44",X"33",X"33",X"33",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"04",X"40",X"33",X"00",X"04",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"44",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"33",X"00",X"00",X"00",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"03",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"33",X"93",X"03",X"33",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"03",X"33",X"33",X"22",X"33",X"33",X"33",X"00",X"3F",X"FF",
		X"00",X"00",X"33",X"33",X"20",X"20",X"22",X"33",X"03",X"FF",X"FF",X"FF",X"00",X"00",X"33",X"33",
		X"00",X"00",X"20",X"20",X"33",X"FF",X"FF",X"FF",X"00",X"00",X"33",X"02",X"00",X"00",X"00",X"02",
		X"33",X"3F",X"FF",X"FF",X"00",X"03",X"93",X"20",X"00",X"00",X"00",X"00",X"23",X"FF",X"FF",X"FF",
		X"00",X"03",X"92",X"02",X"00",X"00",X"00",X"02",X"33",X"03",X"FF",X"FF",X"00",X"03",X"30",X"00",
		X"00",X"00",X"00",X"00",X"22",X"93",X"FF",X"FF",X"00",X"03",X"32",X"00",X"00",X"00",X"00",X"00",
		X"03",X"3F",X"FF",X"FF",X"00",X"03",X"33",X"00",X"00",X"00",X"00",X"02",X"22",X"3F",X"FF",X"FF",
		X"00",X"00",X"33",X"00",X"00",X"00",X"00",X"00",X"23",X"3F",X"FF",X"FF",X"00",X"00",X"33",X"00",
		X"20",X"00",X"00",X"00",X"33",X"3F",X"FF",X"FF",X"00",X"00",X"33",X"22",X"00",X"00",X"00",X"00",
		X"23",X"FF",X"FF",X"FF",X"00",X"00",X"03",X"33",X"22",X"00",X"02",X"32",X"33",X"00",X"3F",X"FF",
		X"00",X"00",X"00",X"03",X"33",X"22",X"23",X"33",X"3F",X"FF",X"FF",X"FF",X"00",X"30",X"03",X"00",
		X"33",X"33",X"33",X"33",X"FF",X"FF",X"FF",X"FF",X"00",X"30",X"03",X"00",X"03",X"03",X"33",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"03",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",
		X"03",X"00",X"3F",X"FF",X"00",X"00",X"00",X"00",X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"03",X"33",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"33",X"13",X"33",X"30",X"00",X"00",X"03",X"FF",X"00",X"00",X"00",X"00",X"31",X"11",X"13",X"11",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"03",X"31",X"01",X"11",X"11",X"3F",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"03",X"30",X"11",X"11",X"13",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"03",
		X"10",X"11",X"11",X"3F",X"FF",X"FF",X"FF",X"FF",X"03",X"00",X"00",X"03",X"31",X"11",X"11",X"33",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"03",X"11",X"11",X"11",X"3F",X"FF",X"FF",X"FF",X"FF",
		X"03",X"00",X"00",X"00",X"31",X"10",X"13",X"3F",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"0A",X"11",X"13",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"03",X"33",X"33",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"03",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"90",X"03",X"3F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"33",X"33",X"33",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"03",
		X"33",X"44",X"43",X"33",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"33",X"44",X"66",X"64",X"43",
		X"3F",X"FF",X"FF",X"FF",X"00",X"00",X"03",X"44",X"36",X"67",X"86",X"44",X"33",X"FF",X"FF",X"FF",
		X"00",X"00",X"03",X"46",X"66",X"77",X"77",X"64",X"33",X"30",X"03",X"FF",X"00",X"00",X"34",X"66",
		X"77",X"88",X"78",X"86",X"44",X"4F",X"FF",X"FF",X"00",X"00",X"34",X"68",X"78",X"11",X"18",X"88",
		X"64",X"33",X"FF",X"FF",X"00",X"03",X"36",X"88",X"81",X"11",X"11",X"88",X"64",X"33",X"FF",X"FF",
		X"00",X"03",X"46",X"88",X"11",X"11",X"11",X"88",X"63",X"33",X"FF",X"FF",X"00",X"03",X"46",X"88",
		X"11",X"11",X"11",X"17",X"64",X"33",X"FF",X"FF",X"00",X"03",X"34",X"88",X"11",X"11",X"11",X"17",
		X"64",X"4F",X"FF",X"FF",X"00",X"03",X"46",X"87",X"81",X"11",X"11",X"87",X"86",X"33",X"FF",X"FF",
		X"00",X"33",X"46",X"67",X"81",X"11",X"18",X"77",X"64",X"4F",X"FF",X"FF",X"00",X"00",X"34",X"68",
		X"88",X"11",X"87",X"76",X"63",X"3F",X"FF",X"FF",X"00",X"00",X"34",X"68",X"78",X"88",X"78",X"64",
		X"43",X"3F",X"FF",X"FF",X"00",X"00",X"33",X"46",X"77",X"77",X"86",X"44",X"43",X"FF",X"FF",X"FF",
		X"00",X"00",X"03",X"34",X"66",X"66",X"64",X"43",X"3F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"33",
		X"44",X"44",X"43",X"33",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"33",X"33",X"33",X"3F",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"02",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"20",
		X"00",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"70",X"7F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"07",X"08",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"7F",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"07",X"00",X"77",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"1F",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"2F",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"02",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"07",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"70",
		X"00",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"70",X"7F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"07",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"7F",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"07",X"00",X"77",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"1F",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"7F",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"07",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"8F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"70",X"00",X"6F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"9F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"06",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"6F",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"08",X"88",X"8F",X"FF",X"FF",X"FF",X"00",X"08",X"88",X"99",X"88",X"8F",X"FF",X"FF",
		X"00",X"88",X"99",X"99",X"99",X"88",X"FF",X"FF",X"08",X"89",X"9A",X"AA",X"A9",X"98",X"8F",X"FF",
		X"08",X"99",X"AA",X"BB",X"AA",X"99",X"8F",X"FF",X"88",X"9A",X"AB",X"BB",X"BA",X"A9",X"88",X"FF",
		X"89",X"9A",X"BB",X"CC",X"BB",X"A9",X"98",X"FF",X"89",X"9A",X"BC",X"CC",X"CB",X"A9",X"98",X"FF",
		X"89",X"9A",X"BC",X"CC",X"CB",X"A9",X"98",X"FF",X"89",X"9A",X"BB",X"CC",X"BB",X"A9",X"98",X"FF",
		X"88",X"9A",X"AB",X"BB",X"BA",X"A9",X"88",X"FF",X"08",X"99",X"AA",X"BB",X"AA",X"99",X"8F",X"FF",
		X"08",X"89",X"9A",X"AA",X"A9",X"98",X"8F",X"FF",X"00",X"88",X"99",X"99",X"99",X"88",X"FF",X"FF",
		X"00",X"08",X"88",X"99",X"88",X"8F",X"FF",X"FF",X"00",X"00",X"08",X"88",X"8F",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"09",X"99",X"9F",X"FF",X"FF",X"FF",X"00",X"09",X"99",X"AA",X"99",X"9F",X"FF",X"FF",
		X"00",X"99",X"AA",X"AA",X"AA",X"99",X"FF",X"FF",X"09",X"9A",X"AB",X"BB",X"BA",X"A9",X"9F",X"FF",
		X"09",X"AA",X"BB",X"CC",X"BB",X"AA",X"9F",X"FF",X"99",X"AB",X"BC",X"CC",X"CB",X"BA",X"99",X"FF",
		X"9A",X"AB",X"CC",X"DD",X"CC",X"BA",X"A9",X"FF",X"9A",X"AB",X"CD",X"DD",X"DC",X"BA",X"A9",X"FF",
		X"9A",X"AB",X"CD",X"DD",X"DC",X"BA",X"A9",X"FF",X"9A",X"AB",X"CC",X"DD",X"CC",X"BA",X"A9",X"FF",
		X"99",X"AB",X"BC",X"CC",X"CB",X"BA",X"99",X"FF",X"09",X"AA",X"BB",X"CC",X"BB",X"AA",X"9F",X"FF",
		X"09",X"9A",X"AB",X"BB",X"BA",X"A9",X"9F",X"FF",X"00",X"99",X"AA",X"AA",X"AA",X"99",X"FF",X"FF",
		X"00",X"09",X"99",X"AA",X"99",X"9F",X"FF",X"FF",X"00",X"00",X"09",X"99",X"9F",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"0A",X"AA",X"AF",X"FF",X"FF",X"FF",X"00",X"0A",X"AA",X"BB",X"AA",X"AF",X"FF",X"FF",
		X"00",X"AA",X"BB",X"BB",X"BB",X"AA",X"FF",X"FF",X"0A",X"AB",X"BC",X"CC",X"CB",X"BA",X"AF",X"FF",
		X"0A",X"BB",X"CC",X"DD",X"CC",X"BB",X"AF",X"FF",X"AA",X"BC",X"CD",X"DD",X"DC",X"CB",X"AA",X"FF",
		X"AB",X"BC",X"DD",X"EE",X"DD",X"CB",X"BA",X"FF",X"AB",X"CC",X"DE",X"EE",X"ED",X"CC",X"BA",X"FF",
		X"AB",X"CC",X"DE",X"EE",X"ED",X"CC",X"BA",X"FF",X"AB",X"BC",X"DD",X"EE",X"DD",X"CB",X"BA",X"FF",
		X"AA",X"BC",X"CD",X"DD",X"DC",X"CB",X"AA",X"FF",X"0A",X"BB",X"CC",X"DD",X"CC",X"BB",X"AF",X"FF",
		X"0A",X"AB",X"BC",X"CC",X"CB",X"BA",X"AF",X"FF",X"00",X"AA",X"BB",X"BB",X"BB",X"AA",X"FF",X"FF",
		X"00",X"0A",X"AA",X"BB",X"AA",X"AF",X"FF",X"FF",X"00",X"00",X"0A",X"AA",X"AF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"0A",X"AA",X"AF",X"FF",X"FF",X"FF",X"00",X"0A",X"AA",X"CC",X"AA",X"AF",X"FF",X"FF",
		X"00",X"AA",X"CC",X"CC",X"CC",X"AA",X"FF",X"FF",X"0A",X"AC",X"CD",X"DD",X"DC",X"CA",X"AF",X"FF",
		X"0A",X"CC",X"DD",X"EE",X"DD",X"CC",X"AF",X"FF",X"AA",X"CD",X"DE",X"EE",X"ED",X"DC",X"AA",X"FF",
		X"AC",X"CD",X"EE",X"EE",X"EE",X"DC",X"CA",X"FF",X"AC",X"CD",X"EE",X"EE",X"EE",X"DC",X"CA",X"FF",
		X"AC",X"CD",X"EE",X"EE",X"EE",X"DC",X"CA",X"FF",X"AC",X"CD",X"EE",X"EE",X"EE",X"DC",X"CA",X"FF",
		X"AA",X"CD",X"DE",X"EE",X"ED",X"DC",X"AA",X"FF",X"0A",X"CC",X"DD",X"EE",X"DD",X"CC",X"AF",X"FF",
		X"0A",X"AC",X"CD",X"DD",X"DC",X"CA",X"AF",X"FF",X"00",X"AA",X"CC",X"CC",X"CC",X"AA",X"FF",X"FF",
		X"00",X"0A",X"AA",X"CC",X"AA",X"AF",X"FF",X"FF",X"00",X"00",X"0A",X"AA",X"AF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"0B",X"BB",X"BF",X"FF",X"FF",X"FF",X"00",X"0B",X"BB",X"EE",X"BB",X"BF",X"FF",X"FF",
		X"00",X"BB",X"EE",X"EE",X"EE",X"BB",X"FF",X"FF",X"0B",X"BE",X"EB",X"BB",X"BE",X"EB",X"BF",X"FF",
		X"0B",X"EE",X"BB",X"66",X"BB",X"EE",X"BF",X"FF",X"BB",X"EB",X"B6",X"66",X"6B",X"BE",X"BB",X"FF",
		X"BE",X"EB",X"66",X"66",X"66",X"BE",X"EB",X"FF",X"BE",X"EB",X"66",X"66",X"66",X"BE",X"EB",X"FF",
		X"BE",X"EB",X"66",X"66",X"66",X"BE",X"EB",X"FF",X"BE",X"EB",X"66",X"66",X"66",X"BE",X"EB",X"FF",
		X"BB",X"EB",X"B6",X"66",X"6B",X"BE",X"BB",X"FF",X"0B",X"EE",X"BB",X"66",X"BB",X"EE",X"BF",X"FF",
		X"0B",X"BE",X"EB",X"BB",X"BE",X"EB",X"BF",X"FF",X"00",X"BB",X"EE",X"EE",X"EE",X"BB",X"FF",X"FF",
		X"00",X"0B",X"BB",X"EE",X"BB",X"BF",X"FF",X"FF",X"00",X"00",X"0B",X"BB",X"BF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"88",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"88",X"88",X"88",X"FF",X"FF",X"FF",X"00",X"08",X"89",X"99",X"98",X"8F",X"FF",X"FF",
		X"00",X"88",X"99",X"AA",X"99",X"88",X"FF",X"FF",X"00",X"89",X"9A",X"AA",X"A9",X"98",X"FF",X"FF",
		X"08",X"89",X"AA",X"BB",X"AA",X"98",X"8F",X"FF",X"08",X"89",X"AB",X"BB",X"BA",X"98",X"8F",X"FF",
		X"08",X"89",X"AB",X"BB",X"BA",X"98",X"8F",X"FF",X"08",X"89",X"AA",X"BB",X"AA",X"98",X"8F",X"FF",
		X"00",X"89",X"9A",X"AA",X"A9",X"98",X"FF",X"FF",X"00",X"88",X"99",X"AA",X"99",X"88",X"FF",X"FF",
		X"00",X"08",X"89",X"99",X"98",X"8F",X"FF",X"FF",X"00",X"00",X"88",X"88",X"88",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"88",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"08",X"88",X"8F",X"FF",X"FF",X"FF",X"00",X"08",X"88",X"00",X"88",X"8F",X"FF",X"FF",
		X"00",X"88",X"00",X"00",X"00",X"88",X"FF",X"FF",X"08",X"80",X"08",X"88",X"80",X"08",X"8F",X"FF",
		X"08",X"00",X"88",X"99",X"88",X"00",X"8F",X"FF",X"88",X"08",X"89",X"99",X"98",X"80",X"88",X"FF",
		X"80",X"08",X"99",X"AA",X"99",X"80",X"08",X"FF",X"80",X"08",X"9A",X"AA",X"A9",X"80",X"08",X"FF",
		X"80",X"08",X"9A",X"AA",X"A9",X"80",X"08",X"FF",X"80",X"08",X"99",X"AA",X"99",X"80",X"08",X"FF",
		X"88",X"08",X"89",X"99",X"98",X"80",X"88",X"FF",X"08",X"00",X"88",X"99",X"88",X"00",X"8F",X"FF",
		X"08",X"80",X"08",X"88",X"80",X"08",X"8F",X"FF",X"00",X"88",X"00",X"00",X"00",X"88",X"FF",X"FF",
		X"00",X"08",X"88",X"00",X"88",X"8F",X"FF",X"FF",X"00",X"00",X"08",X"88",X"8F",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"88",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"88",X"88",X"88",X"FF",X"FF",X"FF",X"00",X"08",X"80",X"00",X"08",X"8F",X"FF",X"FF",
		X"00",X"88",X"00",X"88",X"00",X"88",X"FF",X"FF",X"00",X"80",X"08",X"88",X"80",X"08",X"FF",X"FF",
		X"08",X"80",X"88",X"99",X"88",X"08",X"8F",X"FF",X"08",X"80",X"89",X"99",X"98",X"08",X"8F",X"FF",
		X"08",X"80",X"89",X"99",X"98",X"08",X"8F",X"FF",X"08",X"80",X"88",X"99",X"88",X"08",X"8F",X"FF",
		X"00",X"80",X"08",X"88",X"80",X"08",X"FF",X"FF",X"00",X"88",X"00",X"88",X"00",X"88",X"FF",X"FF",
		X"00",X"08",X"80",X"00",X"08",X"8F",X"FF",X"FF",X"00",X"00",X"88",X"88",X"88",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"88",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"90",X"00",X"09",X"8F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"09",X"FF",X"FF",X"FF",
		X"00",X"9F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"09",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"09",X"FF",X"FF",X"00",X"9F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"09",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"90",X"00",X"09",X"FF",X"FF",X"00",X"09",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"09",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"9F",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"08",X"00",X"09",X"FF",X"FF",X"00",X"00",X"00",X"00",X"08",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"9F",X"FF",X"08",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"80",X"00",X"00",X"00",X"00",X"00",X"08",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"8F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"9F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"80",X"08",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"08",X"00",X"00",X"80",X"8F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"09",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"09",X"00",X"F9",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"09",X"C0",X"CF",X"FF",X"FF",X"FF",X"00",X"00",X"99",X"C7",X"CC",X"FF",X"FF",X"FF",
		X"00",X"09",X"99",X"C7",X"CC",X"CF",X"FF",X"FF",X"00",X"99",X"99",X"C7",X"EC",X"CC",X"FF",X"FF",
		X"09",X"99",X"99",X"E7",X"EE",X"CC",X"CF",X"FF",X"99",X"99",X"99",X"E7",X"EE",X"EC",X"CC",X"FF",
		X"07",X"77",X"77",X"77",X"77",X"77",X"7F",X"FF",X"AA",X"AA",X"AE",X"E7",X"EE",X"CC",X"CC",X"FF",
		X"88",X"88",X"88",X"E7",X"EA",X"AA",X"AA",X"FF",X"08",X"88",X"88",X"67",X"BA",X"AA",X"AF",X"FF",
		X"00",X"88",X"88",X"67",X"BA",X"AA",X"FF",X"FF",X"00",X"08",X"88",X"67",X"BA",X"AF",X"FF",X"FF",
		X"00",X"00",X"88",X"67",X"BA",X"FF",X"FF",X"FF",X"00",X"00",X"08",X"60",X"BF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"09",X"C0",X"DF",X"FF",X"FF",X"FF",X"00",X"00",X"99",X"C7",X"DD",X"FF",X"FF",X"FF",
		X"00",X"09",X"99",X"B7",X"BD",X"DF",X"FF",X"FF",X"00",X"99",X"99",X"B7",X"ED",X"DD",X"FF",X"FF",
		X"09",X"99",X"99",X"E7",X"ED",X"DD",X"DF",X"FF",X"99",X"99",X"99",X"E7",X"BD",X"DD",X"DD",X"FF",
		X"07",X"99",X"99",X"B7",X"CD",X"DD",X"7F",X"FF",X"AA",X"77",X"99",X"B7",X"DD",X"77",X"CC",X"FF",
		X"88",X"AA",X"77",X"B7",X"77",X"CC",X"AA",X"FF",X"08",X"88",X"AA",X"77",X"EE",X"AA",X"AF",X"FF",
		X"00",X"88",X"88",X"67",X"AA",X"AA",X"FF",X"FF",X"00",X"08",X"88",X"67",X"AA",X"AF",X"FF",X"FF",
		X"00",X"00",X"88",X"67",X"AA",X"FF",X"FF",X"FF",X"00",X"00",X"08",X"60",X"AF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"08",X"E0",X"EF",X"FF",X"FF",X"FF",X"00",X"00",X"88",X"E7",X"ED",X"FF",X"FF",X"FF",
		X"00",X"08",X"88",X"E7",X"ED",X"DF",X"FF",X"FF",X"00",X"88",X"88",X"E7",X"BD",X"DD",X"FF",X"FF",
		X"08",X"88",X"88",X"B7",X"BD",X"DD",X"DF",X"FF",X"88",X"88",X"88",X"B7",X"CD",X"DD",X"DD",X"FF",
		X"08",X"88",X"88",X"C7",X"CD",X"DD",X"DF",X"FF",X"B7",X"88",X"88",X"C7",X"DD",X"DD",X"7C",X"FF",
		X"8B",X"78",X"88",X"C7",X"DD",X"D7",X"CB",X"FF",X"08",X"B7",X"88",X"C7",X"DD",X"7C",X"BF",X"FF",
		X"00",X"8B",X"78",X"C7",X"D7",X"EB",X"FF",X"FF",X"00",X"08",X"B7",X"C7",X"7E",X"BF",X"FF",X"FF",
		X"00",X"00",X"8B",X"77",X"DB",X"FF",X"FF",X"FF",X"00",X"00",X"08",X"B0",X"BF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"09",X"C7",X"CF",X"FF",X"FF",X"FF",
		X"00",X"00",X"98",X"C7",X"CC",X"FF",X"FF",X"FF",X"00",X"09",X"88",X"C7",X"CC",X"CF",X"FF",X"FF",
		X"00",X"98",X"88",X"C7",X"CC",X"CC",X"FF",X"FF",X"09",X"88",X"88",X"C7",X"CC",X"CC",X"CF",X"FF",
		X"98",X"88",X"88",X"C7",X"CC",X"CC",X"CC",X"FF",X"88",X"88",X"88",X"C7",X"CC",X"CC",X"CC",X"FF",
		X"08",X"88",X"88",X"C7",X"CC",X"CC",X"CF",X"FF",X"00",X"88",X"88",X"C7",X"CC",X"CC",X"FF",X"FF",
		X"00",X"08",X"88",X"C7",X"CC",X"CF",X"FF",X"FF",X"00",X"00",X"88",X"C7",X"CC",X"FF",X"FF",X"FF",
		X"00",X"00",X"08",X"C7",X"CF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"09",X"0A",X"CF",X"FF",X"FF",X"FF",X"00",X"00",X"98",X"77",X"AC",X"FF",X"FF",X"FF",
		X"00",X"09",X"87",X"C7",X"7A",X"CF",X"FF",X"FF",X"00",X"98",X"78",X"C7",X"C7",X"AC",X"FF",X"FF",
		X"09",X"87",X"88",X"C7",X"BC",X"7A",X"CF",X"FF",X"98",X"78",X"88",X"C7",X"BB",X"C7",X"AC",X"FF",
		X"87",X"88",X"88",X"B7",X"BB",X"BC",X"7A",X"FF",X"08",X"88",X"88",X"B7",X"BB",X"BC",X"CF",X"FF",
		X"88",X"88",X"88",X"B7",X"BB",X"BB",X"CC",X"FF",X"08",X"88",X"88",X"B7",X"BB",X"BB",X"BF",X"FF",
		X"00",X"88",X"88",X"B7",X"BB",X"BB",X"FF",X"FF",X"00",X"08",X"88",X"B7",X"BB",X"BF",X"FF",X"FF",
		X"00",X"00",X"88",X"B7",X"BB",X"FF",X"FF",X"FF",X"00",X"00",X"08",X"B0",X"BF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"09",X"E0",X"CF",X"FF",X"FF",X"FF",X"00",X"00",X"99",X"E7",X"EC",X"FF",X"FF",X"FF",
		X"00",X"09",X"99",X"E7",X"EE",X"CF",X"FF",X"FF",X"00",X"99",X"88",X"77",X"AA",X"EC",X"FF",X"FF",
		X"09",X"88",X"77",X"E7",X"77",X"AA",X"CF",X"FF",X"98",X"77",X"88",X"E7",X"EE",X"77",X"AC",X"FF",
		X"07",X"88",X"88",X"C7",X"EC",X"CC",X"7F",X"FF",X"88",X"88",X"88",X"C7",X"BB",X"CC",X"CC",X"FF",
		X"88",X"88",X"88",X"C7",X"BB",X"BB",X"CC",X"FF",X"08",X"88",X"88",X"C7",X"BB",X"BB",X"BF",X"FF",
		X"00",X"88",X"88",X"C7",X"BB",X"BB",X"FF",X"FF",X"00",X"08",X"88",X"C7",X"BB",X"BF",X"FF",X"FF",
		X"00",X"00",X"88",X"C7",X"BB",X"FF",X"FF",X"FF",X"00",X"00",X"08",X"C0",X"BF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"09",X"C0",X"DF",X"FF",X"FF",X"FF",X"00",X"00",X"99",X"C7",X"DD",X"FF",X"FF",X"FF",
		X"00",X"09",X"9C",X"7D",X"DD",X"DF",X"FF",X"FF",X"00",X"99",X"9C",X"7D",X"DD",X"DD",X"FF",X"FF",
		X"09",X"99",X"E7",X"DD",X"DD",X"DD",X"DF",X"FF",X"99",X"99",X"E7",X"DC",X"BE",X"EB",X"DD",X"FF",
		X"07",X"77",X"77",X"77",X"77",X"77",X"7F",X"FF",X"66",X"66",X"7B",X"BB",X"EE",X"BB",X"CC",X"FF",
		X"88",X"88",X"A7",X"AA",X"AA",X"AA",X"AA",X"FF",X"08",X"88",X"A7",X"AA",X"AA",X"AA",X"AF",X"FF",
		X"00",X"88",X"8A",X"7A",X"AA",X"AA",X"FF",X"FF",X"00",X"08",X"8A",X"7A",X"AA",X"AF",X"FF",X"FF",
		X"00",X"00",X"88",X"A7",X"AA",X"FF",X"FF",X"FF",X"00",X"00",X"08",X"A0",X"AF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"09",X"C0",X"DF",X"FF",X"FF",X"FF",X"00",X"00",X"9C",X"7D",X"DD",X"FF",X"FF",X"FF",
		X"00",X"09",X"C7",X"DD",X"DD",X"DF",X"FF",X"FF",X"00",X"9B",X"7D",X"DD",X"DD",X"DD",X"FF",X"FF",
		X"09",X"B7",X"DD",X"DD",X"DD",X"DD",X"DF",X"FF",X"9B",X"7D",X"DD",X"DC",X"CB",X"BE",X"EE",X"FF",
		X"07",X"77",X"77",X"77",X"77",X"77",X"7F",X"FF",X"B7",X"CC",X"CC",X"CC",X"BB",X"EE",X"EE",X"FF",
		X"8B",X"79",X"99",X"99",X"99",X"99",X"99",X"FF",X"08",X"B7",X"99",X"99",X"99",X"99",X"9F",X"FF",
		X"00",X"9B",X"79",X"99",X"99",X"99",X"FF",X"FF",X"00",X"08",X"B7",X"99",X"99",X"9F",X"FF",X"FF",
		X"00",X"00",X"8B",X"79",X"99",X"FF",X"FF",X"FF",X"00",X"00",X"08",X"B0",X"9F",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"CC",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"0C",X"CC",X"CF",X"FF",X"FF",X"FF",
		X"00",X"00",X"CC",X"CC",X"CC",X"FF",X"FF",X"FF",X"00",X"0C",X"CC",X"CC",X"CC",X"CF",X"FF",X"FF",
		X"00",X"CC",X"CC",X"CC",X"CC",X"CC",X"FF",X"FF",X"0C",X"CC",X"CC",X"CC",X"CC",X"CC",X"CF",X"FF",
		X"07",X"77",X"77",X"77",X"77",X"77",X"7F",X"FF",X"0C",X"CC",X"CC",X"CC",X"CC",X"CC",X"CF",X"FF",
		X"09",X"99",X"99",X"99",X"99",X"99",X"9F",X"FF",X"00",X"99",X"99",X"99",X"99",X"99",X"FF",X"FF",
		X"00",X"09",X"99",X"99",X"99",X"9F",X"FF",X"FF",X"00",X"00",X"99",X"99",X"99",X"FF",X"FF",X"FF",
		X"00",X"00",X"09",X"99",X"9F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"99",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"0C",X"0A",X"CF",X"FF",X"FF",X"FF",X"00",X"00",X"BC",X"C7",X"AC",X"FF",X"FF",X"FF",
		X"00",X"0B",X"BB",X"CC",X"7A",X"CF",X"FF",X"FF",X"00",X"BB",X"BB",X"BB",X"C7",X"AC",X"FF",X"FF",
		X"0B",X"BB",X"BB",X"BB",X"BC",X"7A",X"EF",X"FF",X"BB",X"BB",X"BB",X"BB",X"BB",X"C7",X"AE",X"FF",
		X"07",X"77",X"77",X"77",X"77",X"77",X"7A",X"FF",X"BB",X"BB",X"BB",X"BB",X"CC",X"CC",X"7F",X"FF",
		X"88",X"88",X"88",X"88",X"88",X"87",X"8A",X"FF",X"08",X"88",X"88",X"88",X"88",X"78",X"AF",X"FF",
		X"00",X"88",X"88",X"88",X"87",X"8A",X"FF",X"FF",X"00",X"08",X"88",X"88",X"78",X"AF",X"FF",X"FF",
		X"00",X"00",X"88",X"87",X"8A",X"FF",X"FF",X"FF",X"00",X"00",X"08",X"08",X"AF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"0A",X"C0",X"CF",X"FF",X"FF",X"FF",X"00",X"00",X"AA",X"C7",X"9C",X"FF",X"FF",X"FF",
		X"00",X"0A",X"AA",X"AC",X"79",X"CF",X"FF",X"FF",X"00",X"AA",X"AA",X"AC",X"79",X"EC",X"FF",X"FF",
		X"0A",X"AA",X"AA",X"AC",X"E7",X"9E",X"CF",X"FF",X"AA",X"AA",X"AA",X"AE",X"E7",X"9E",X"EC",X"FF",
		X"07",X"77",X"77",X"77",X"77",X"77",X"7F",X"FF",X"BB",X"BB",X"BB",X"BB",X"EE",X"7E",X"EE",X"FF",
		X"88",X"88",X"88",X"88",X"87",X"8A",X"AA",X"FF",X"08",X"88",X"88",X"88",X"87",X"8A",X"AF",X"FF",
		X"00",X"88",X"88",X"88",X"78",X"AA",X"FF",X"FF",X"00",X"08",X"88",X"88",X"78",X"AF",X"FF",X"FF",
		X"00",X"00",X"88",X"87",X"8A",X"FF",X"FF",X"FF",X"00",X"00",X"08",X"80",X"9F",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"00",X"B2",X"E0",X"00",X"00",X"00",X"00",X"00",X"B2",X"EF",X"FF",X"0B",X"B1",
		X"EE",X"00",X"00",X"00",X"00",X"0B",X"B1",X"EE",X"FF",X"AB",X"B9",X"6E",X"E0",X"00",X"00",X"00",
		X"AB",X"B9",X"6E",X"EF",X"BB",X"41",X"46",X"E0",X"00",X"00",X"00",X"BB",X"41",X"46",X"EF",X"59",
		X"15",X"1A",X"50",X"00",X"00",X"00",X"59",X"15",X"1A",X"5F",X"AA",X"41",X"4D",X"D0",X"00",X"00",
		X"00",X"AA",X"41",X"4D",X"DF",X"AA",X"A9",X"DD",X"B0",X"00",X"00",X"00",X"AA",X"A9",X"DD",X"BF",
		X"0A",X"A5",X"DB",X"00",X"00",X"00",X"00",X"0A",X"A5",X"DB",X"FF",X"00",X"A1",X"A0",X"00",X"0B",
		X"2E",X"00",X"00",X"A1",X"AF",X"FF",X"00",X"00",X"00",X"00",X"AB",X"1E",X"EF",X"FF",X"FF",X"FF",
		X"FF",X"00",X"00",X"00",X"0A",X"BB",X"96",X"EE",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"0B",
		X"B4",X"14",X"6E",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"05",X"91",X"51",X"A5",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"0A",X"A4",X"14",X"DD",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",
		X"0A",X"AA",X"9D",X"DB",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"AA",X"5D",X"BF",X"FF",
		X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"0A",X"1A",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"2E",
		X"3E",X"2E",X"3E",X"2F",X"FF",X"2E",X"3E",X"2E",X"3E",X"2F",X"FF",X"2E",X"3E",X"2E",X"3E",X"2F",
		X"FF",X"EE",X"EE",X"EE",X"EE",X"EF",X"FF",X"99",X"99",X"99",X"99",X"7F",X"FF",X"55",X"55",X"55",
		X"55",X"6C",X"FF",X"EE",X"E4",X"44",X"7E",X"66",X"CF",X"EE",X"E4",X"44",X"7E",X"66",X"CF",X"EE",
		X"E4",X"44",X"77",X"66",X"CF",X"EE",X"E5",X"55",X"55",X"66",X"CF",X"EE",X"E6",X"66",X"66",X"66",
		X"CF",X"EE",X"EB",X"BB",X"BB",X"69",X"AF",X"77",X"77",X"77",X"77",X"77",X"FF",X"DD",X"DD",X"DD",
		X"DD",X"DF",X"FF",X"EE",X"EE",X"EE",X"EE",X"EF",X"FF",X"2E",X"3E",X"2E",X"3E",X"2F",X"FF",X"2E",
		X"3E",X"2E",X"3E",X"2F",X"FF",X"2E",X"3E",X"2E",X"3E",X"2F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3E",X"2E",X"3E",X"2E",X"3F",X"FF",X"3E",X"2E",X"3E",
		X"2E",X"3F",X"FF",X"3E",X"2E",X"3E",X"2E",X"3F",X"FF",X"EE",X"EE",X"EE",X"EE",X"EF",X"FF",X"99",
		X"99",X"99",X"99",X"7F",X"FF",X"55",X"55",X"55",X"55",X"6C",X"FF",X"11",X"E4",X"44",X"7E",X"66",
		X"CF",X"11",X"E4",X"44",X"7E",X"66",X"CF",X"EE",X"E4",X"44",X"77",X"66",X"CF",X"EE",X"E5",X"55",
		X"55",X"66",X"CF",X"11",X"E6",X"66",X"66",X"66",X"CF",X"11",X"EB",X"BB",X"BB",X"69",X"AF",X"77",
		X"77",X"77",X"77",X"77",X"FF",X"DD",X"DD",X"DD",X"DD",X"DF",X"FF",X"EE",X"EE",X"EE",X"EE",X"EF",
		X"FF",X"3E",X"2E",X"3E",X"2E",X"3F",X"FF",X"3E",X"2E",X"3E",X"2E",X"3F",X"FF",X"3E",X"2E",X"3E",
		X"2E",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"B8",X"88",X"88",X"88",
		X"88",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"0B",X"BA",X"88",X"88",X"88",X"88",
		X"88",X"8F",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"0D",X"AA",X"9A",X"AA",X"AA",X"AA",X"66",
		X"66",X"6F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"D9",X"98",X"AA",X"AA",X"AA",X"AA",X"66",
		X"64",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"0D",X"88",X"7A",X"AA",X"AA",X"AA",X"AD",X"34",
		X"4F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"D7",X"76",X"AA",X"AA",X"AA",X"DD",X"53",X"44",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"0D",X"66",X"5A",X"AA",X"AA",X"D7",X"53",X"34",X"7F",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"D5",X"54",X"AA",X"AE",X"E6",X"53",X"13",X"4F",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"44",X"3A",X"AE",X"66",X"43",X"13",X"47",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"D3",X"32",X"DE",X"65",X"43",X"13",X"46",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0D",X"22",X"D7",X"65",X"43",X"13",X"44",X"FF",X"0B",X"D0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"DD",X"D7",X"65",X"43",X"11",X"33",X"6F",X"BB",X"AD",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0D",X"76",X"54",X"43",X"11",X"23",X"6F",X"CA",X"A9",X"D0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"D6",X"54",X"33",X"11",X"23",X"6F",X"BB",X"9A",X"8D",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0D",X"54",X"31",X"11",X"23",X"5F",X"BB",X"C8",X"87",X"D0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"D4",X"31",X"11",X"23",X"5F",X"BB",X"CC",X"77",X"6D",X"00",X"00",X"00",X"00",
		X"00",X"0C",X"DD",X"31",X"11",X"23",X"5F",X"BB",X"CC",X"C6",X"65",X"D0",X"00",X"00",X"00",X"00",
		X"CC",X"BD",X"D1",X"AA",X"23",X"5F",X"BB",X"BC",X"CC",X"55",X"4D",X"00",X"00",X"00",X"00",X"CC",
		X"BA",X"DD",X"A9",X"93",X"5F",X"CB",X"BC",X"CC",X"C4",X"43",X"D0",X"00",X"00",X"0C",X"CB",X"BA",
		X"9D",X"D9",X"88",X"5F",X"0B",X"BC",X"CC",X"CC",X"33",X"2D",X"00",X"00",X"0C",X"CB",X"AA",X"98",
		X"DD",X"87",X"7F",X"0B",X"BC",X"CC",X"CC",X"C2",X"2D",X"D0",X"00",X"CC",X"BB",X"A9",X"98",X"7D",
		X"D7",X"6F",X"0B",X"BB",X"CC",X"CC",X"CC",X"DD",X"7D",X"0C",X"CC",X"BA",X"A9",X"88",X"76",X"DD",
		X"5F",X"0C",X"BB",X"CC",X"CC",X"CC",X"D8",X"76",X"DC",X"CB",X"BA",X"A9",X"88",X"76",X"5D",X"DF",
		X"00",X"BB",X"CC",X"CC",X"CC",X"E8",X"76",X"5D",X"DB",X"AA",X"99",X"87",X"76",X"54",X"DF",X"00",
		X"BB",X"BC",X"CC",X"CE",X"E8",X"76",X"54",X"DD",X"AA",X"98",X"87",X"66",X"54",X"FF",X"00",X"CB",
		X"BC",X"CC",X"CE",X"88",X"76",X"64",X"4D",X"D9",X"98",X"77",X"65",X"5F",X"FF",X"00",X"0B",X"BA",
		X"CC",X"DD",X"88",X"76",X"65",X"44",X"DD",X"98",X"77",X"65",X"5F",X"FF",X"00",X"0C",X"BA",X"AC",
		X"D8",X"88",X"77",X"66",X"5A",X"AD",X"D8",X"76",X"65",X"FF",X"FF",X"00",X"00",X"BA",X"AA",X"A8",
		X"88",X"87",X"76",X"5A",X"99",X"DD",X"76",X"55",X"FF",X"FF",X"00",X"00",X"0A",X"AA",X"A9",X"88",
		X"87",X"77",X"65",X"98",X"8D",X"D6",X"5F",X"FF",X"FF",X"00",X"00",X"00",X"BA",X"A9",X"88",X"88",
		X"67",X"77",X"78",X"77",X"DD",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"0B",X"AA",X"98",X"88",X"88",
		X"77",X"79",X"76",X"6F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"BB",X"AA",X"99",X"88",X"88",
		X"99",X"96",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"AA",X"A9",X"99",X"99",X"99",
		X"9F",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"A9",X"AF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"BB",X"BB",X"BB",X"88",X"8F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"BB",X"BB",X"BB",X"B8",X"88",X"77",X"8F",X"FF",X"FF",X"FF",X"FF",X"00",
		X"00",X"00",X"BB",X"BB",X"BB",X"AA",X"AA",X"88",X"76",X"66",X"9F",X"FF",X"FF",X"FF",X"00",X"00",
		X"0B",X"BB",X"BA",X"AA",X"AA",X"AA",X"AD",X"76",X"55",X"55",X"9F",X"FF",X"FF",X"00",X"00",X"8A",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"9D",X"66",X"54",X"44",X"49",X"FF",X"FF",X"00",X"09",X"87",X"6A",
		X"9A",X"AA",X"AA",X"AA",X"DD",X"65",X"44",X"33",X"34",X"FF",X"FF",X"00",X"0D",X"87",X"65",X"5A",
		X"9A",X"AA",X"A9",X"D7",X"65",X"43",X"32",X"23",X"6F",X"FF",X"00",X"00",X"DD",X"75",X"44",X"1A",
		X"AA",X"A9",X"D7",X"65",X"43",X"11",X"22",X"4F",X"FF",X"00",X"00",X"00",X"DD",X"51",X"12",X"3A",
		X"A9",X"D6",X"65",X"44",X"31",X"12",X"37",X"FF",X"00",X"00",X"00",X"00",X"DD",X"22",X"33",X"4D",
		X"D7",X"65",X"44",X"31",X"12",X"35",X"FF",X"00",X"00",X"00",X"00",X"00",X"DD",X"34",X"4D",X"76",
		X"55",X"44",X"31",X"12",X"35",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"DD",X"4D",X"76",X"54",
		X"44",X"31",X"11",X"35",X"6F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DD",X"66",X"54",X"44",
		X"31",X"11",X"35",X"6F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DD",X"54",X"44",X"16",
		X"12",X"35",X"6F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DD",X"41",X"46",X"66",
		X"35",X"6F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7C",X"DD",X"56",X"67",X"86",
		X"6F",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"76",X"4C",X"DD",X"78",X"89",X"9F",
		X"AD",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"64",X"43",X"3C",X"DD",X"89",X"AF",X"A9",
		X"AD",X"D0",X"00",X"00",X"00",X"00",X"00",X"07",X"54",X"33",X"22",X"1C",X"DD",X"BF",X"99",X"87",
		X"7D",X"D0",X"00",X"00",X"00",X"00",X"B7",X"54",X"33",X"21",X"13",X"4C",X"DF",X"BB",X"87",X"66",
		X"5D",X"D0",X"00",X"00",X"00",X"96",X"54",X"32",X"21",X"33",X"45",X"7F",X"BB",X"CA",X"65",X"54",
		X"4D",X"D0",X"00",X"00",X"75",X"44",X"32",X"11",X"34",X"45",X"8F",X"BB",X"CC",X"CA",X"44",X"33",
		X"1D",X"D0",X"09",X"75",X"43",X"32",X"11",X"34",X"57",X"BF",X"BB",X"BC",X"CC",X"CA",X"31",X"1D",
		X"6D",X"D6",X"65",X"43",X"22",X"11",X"44",X"59",X"FF",X"0B",X"BC",X"CC",X"CC",X"CA",X"1D",X"66",
		X"6D",X"DB",X"43",X"21",X"11",X"45",X"58",X"FF",X"0B",X"BB",X"CC",X"CC",X"CC",X"CD",X"66",X"54",
		X"4D",X"DB",X"21",X"13",X"45",X"7B",X"FF",X"0B",X"BB",X"CC",X"CC",X"CC",X"DD",X"66",X"55",X"43",
		X"5D",X"DB",X"34",X"55",X"9F",X"FF",X"00",X"BB",X"BC",X"CC",X"CC",X"D7",X"76",X"55",X"33",X"67",
		X"8D",X"DB",X"57",X"8F",X"FF",X"00",X"BB",X"BC",X"CC",X"CC",X"D7",X"76",X"55",X"37",X"67",X"88",
		X"9D",X"DB",X"BF",X"FF",X"00",X"0B",X"BB",X"CC",X"CD",X"D8",X"77",X"65",X"54",X"57",X"89",X"9A",
		X"AD",X"DF",X"FF",X"00",X"00",X"BB",X"AC",X"CD",X"88",X"77",X"66",X"55",X"54",X"59",X"AA",X"BB",
		X"CF",X"FF",X"00",X"00",X"BB",X"AA",X"CD",X"88",X"87",X"76",X"66",X"55",X"55",X"5B",X"BC",X"FF",
		X"FF",X"00",X"00",X"0B",X"AA",X"A9",X"98",X"88",X"77",X"76",X"66",X"66",X"66",X"6F",X"FF",X"FF",
		X"00",X"00",X"00",X"AA",X"AA",X"99",X"88",X"88",X"77",X"77",X"77",X"77",X"FF",X"FF",X"FF",X"00",
		X"00",X"00",X"0B",X"AA",X"A9",X"98",X"88",X"88",X"88",X"77",X"8F",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"0A",X"AA",X"AA",X"AA",X"9A",X"A8",X"89",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"0A",X"AA",X"AA",X"AA",X"AF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"88",
		X"88",X"88",X"88",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"0B",X"88",X"88",X"88",
		X"88",X"77",X"77",X"8F",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"0B",X"B8",X"88",X"88",X"88",X"77",
		X"65",X"55",X"66",X"8F",X"FF",X"FF",X"FF",X"00",X"00",X"BB",X"B8",X"88",X"88",X"87",X"76",X"54",
		X"44",X"45",X"68",X"FF",X"FF",X"FF",X"00",X"0B",X"BB",X"B8",X"88",X"88",X"87",X"65",X"33",X"33",
		X"44",X"56",X"8F",X"FF",X"FF",X"00",X"BB",X"BB",X"AA",X"AA",X"AA",X"D7",X"54",X"33",X"33",X"34",
		X"45",X"68",X"FF",X"FF",X"0B",X"BB",X"BA",X"AA",X"AA",X"AA",X"D7",X"54",X"33",X"12",X"33",X"44",
		X"56",X"8F",X"FF",X"0B",X"BB",X"AA",X"AA",X"AA",X"AA",X"E7",X"54",X"31",X"11",X"23",X"34",X"56",
		X"8F",X"FF",X"BB",X"BA",X"AA",X"AA",X"AA",X"AA",X"E7",X"54",X"33",X"11",X"12",X"34",X"45",X"68",
		X"FF",X"BB",X"AA",X"AA",X"AA",X"AA",X"AA",X"E7",X"54",X"33",X"11",X"12",X"34",X"45",X"68",X"FF",
		X"12",X"34",X"56",X"78",X"9A",X"BC",X"D7",X"54",X"43",X"15",X"67",X"89",X"AB",X"CD",X"FF",X"12",
		X"34",X"56",X"78",X"9A",X"BC",X"D7",X"54",X"43",X"15",X"67",X"89",X"AB",X"CD",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"12",X"34",X"56",X"78",X"9A",X"BC",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"12",X"34",X"56",X"78",X"9A",X"BC",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"12",X"34",X"56",X"78",X"9A",X"BC",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"12",X"34",X"56",X"78",X"9A",X"BC",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"12",X"34",X"56",X"78",X"9A",X"BC",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"12",X"34",X"56",X"78",X"9A",X"BC",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"12",
		X"34",X"56",X"78",X"9A",X"BC",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"12",X"34",
		X"56",X"78",X"9A",X"BC",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"12",X"34",X"56",
		X"78",X"9A",X"BC",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"12",X"34",X"56",X"78",
		X"9A",X"BC",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"DD",X"FF",X"12",X"34",X"56",X"78",X"9A",X"BC",X"D8",X"75",X"43",X"35",X"67",X"89",X"AB",X"CD",
		X"FF",X"12",X"34",X"56",X"78",X"9A",X"CC",X"D8",X"65",X"54",X"35",X"67",X"89",X"AB",X"CD",X"FF",
		X"BB",X"CC",X"CC",X"CC",X"CC",X"CC",X"E8",X"66",X"55",X"43",X"44",X"55",X"56",X"8B",X"FF",X"BB",
		X"BC",X"CC",X"CC",X"CC",X"CC",X"E8",X"76",X"65",X"54",X"55",X"55",X"66",X"8B",X"FF",X"0B",X"BB",
		X"CC",X"CC",X"CC",X"CC",X"E8",X"77",X"66",X"55",X"55",X"56",X"68",X"BF",X"FF",X"0B",X"BB",X"BC",
		X"CC",X"CC",X"CC",X"D8",X"77",X"66",X"65",X"55",X"66",X"78",X"BF",X"FF",X"00",X"BB",X"BB",X"CC",
		X"CC",X"CC",X"D8",X"87",X"77",X"66",X"66",X"67",X"8B",X"FF",X"FF",X"00",X"0B",X"BB",X"BB",X"BB",
		X"BB",X"BB",X"88",X"77",X"77",X"77",X"78",X"BF",X"FF",X"FF",X"00",X"00",X"BB",X"BB",X"BB",X"BB",
		X"BB",X"B8",X"87",X"77",X"78",X"8B",X"FF",X"FF",X"FF",X"00",X"00",X"0B",X"BB",X"BB",X"BB",X"BB",
		X"BB",X"88",X"88",X"8B",X"BF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"0B",X"BB",X"CC",X"CC",X"CC",
		X"BB",X"BB",X"BF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"CC",X"CC",X"CC",X"CC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"0A",X"AA",X"AA",X"A9",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"08",X"88",X"76",X"66",X"66",X"67",X"7F",X"FF",X"FF",X"FF",
		X"FF",X"00",X"00",X"00",X"0B",X"88",X"87",X"65",X"55",X"55",X"55",X"67",X"7F",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"88",X"88",X"76",X"54",X"44",X"44",X"44",X"56",X"77",X"FF",X"FF",X"FF",X"00",
		X"00",X"0B",X"88",X"88",X"76",X"54",X"31",X"12",X"33",X"45",X"66",X"6F",X"FF",X"FF",X"00",X"00",
		X"BB",X"88",X"AD",X"76",X"54",X"33",X"11",X"22",X"34",X"5B",X"BC",X"FF",X"FF",X"00",X"00",X"BB",
		X"8A",X"AD",X"86",X"65",X"43",X"11",X"11",X"29",X"AA",X"BB",X"CF",X"FF",X"00",X"0B",X"BB",X"AA",
		X"AD",X"88",X"66",X"54",X"31",X"17",X"89",X"9A",X"AD",X"DF",X"FF",X"00",X"BB",X"BA",X"AA",X"AA",
		X"D8",X"76",X"55",X"33",X"67",X"88",X"9D",X"DB",X"BF",X"FF",X"00",X"BB",X"BA",X"AA",X"AA",X"D8",
		X"76",X"65",X"43",X"67",X"8D",X"DB",X"56",X"9F",X"FF",X"0B",X"BB",X"AA",X"AA",X"AA",X"DD",X"87",
		X"65",X"43",X"5D",X"DB",X"34",X"55",X"8F",X"FF",X"0B",X"BB",X"AA",X"AA",X"AA",X"CD",X"86",X"64",
		X"4D",X"DB",X"21",X"13",X"45",X"7B",X"FF",X"0B",X"BA",X"AA",X"AA",X"AA",X"1D",X"87",X"6D",X"DB",
		X"43",X"21",X"11",X"45",X"59",X"FF",X"BB",X"BA",X"AA",X"AA",X"31",X"1D",X"8D",X"D6",X"65",X"43",
		X"22",X"11",X"44",X"58",X"FF",X"BB",X"AA",X"AA",X"44",X"33",X"1D",X"D0",X"09",X"75",X"43",X"32",
		X"11",X"34",X"57",X"BF",X"BB",X"AA",X"65",X"54",X"4D",X"D0",X"00",X"00",X"75",X"44",X"32",X"11",
		X"34",X"45",X"9F",X"BB",X"87",X"66",X"5D",X"D0",X"00",X"00",X"00",X"96",X"54",X"32",X"21",X"33",
		X"45",X"8F",X"99",X"87",X"7D",X"D0",X"00",X"00",X"00",X"00",X"B7",X"54",X"33",X"21",X"13",X"4C",
		X"DF",X"A9",X"AD",X"D0",X"00",X"00",X"00",X"00",X"00",X"07",X"54",X"33",X"22",X"1C",X"DD",X"BF",
		X"AD",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"64",X"43",X"3C",X"DD",X"89",X"AF",X"D0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"76",X"4C",X"DD",X"78",X"89",X"9F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7C",X"DD",X"56",X"67",X"86",X"5F",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"DD",X"44",X"46",X"66",X"44",X"5F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"DD",X"55",X"54",X"46",X"44",X"45",X"6F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"DD",X"86",X"66",X"55",X"44",X"45",X"55",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DD",X"4D",X"87",X"76",X"65",X"55",X"55",X"66",X"FF",X"00",X"00",X"00",X"00",X"00",X"DD",X"34",
		X"4D",X"88",X"77",X"66",X"66",X"66",X"68",X"FF",X"00",X"00",X"00",X"00",X"DD",X"22",X"33",X"4D",
		X"D8",X"67",X"76",X"66",X"66",X"78",X"FF",X"00",X"00",X"00",X"DD",X"51",X"12",X"3C",X"CC",X"D8",
		X"67",X"77",X"77",X"77",X"8F",X"FF",X"00",X"00",X"DD",X"75",X"44",X"1C",X"CC",X"CC",X"D8",X"87",
		X"77",X"77",X"88",X"8F",X"FF",X"00",X"0D",X"87",X"65",X"5C",X"CC",X"CC",X"CC",X"D8",X"88",X"88",
		X"88",X"88",X"FF",X"FF",X"00",X"09",X"87",X"6C",X"CC",X"CC",X"CC",X"CC",X"DD",X"98",X"88",X"88",
		X"88",X"FF",X"FF",X"00",X"00",X"8B",X"BC",X"CC",X"CC",X"CC",X"CC",X"CD",X"99",X"88",X"88",X"8F",
		X"FF",X"FF",X"00",X"00",X"0B",X"BB",X"BC",X"CC",X"CC",X"CC",X"CD",X"99",X"99",X"99",X"FF",X"FF",
		X"FF",X"00",X"00",X"00",X"BB",X"BB",X"BB",X"CC",X"CC",X"AA",X"99",X"AA",X"9F",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"BB",X"BB",X"BB",X"BA",X"AA",X"AA",X"9F",X"FF",X"FF",X"FF",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"BB",X"BB",X"BB",X"9A",X"AF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"76",X"65",X"55",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"76",X"65",X"54",X"44",X"44",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"99",X"76",
		X"54",X"43",X"33",X"33",X"36",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"09",X"88",X"65",X"43",
		X"33",X"22",X"33",X"76",X"6F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"98",X"86",X"54",X"31",X"11",
		X"11",X"18",X"77",X"DF",X"FF",X"FF",X"FF",X"00",X"00",X"09",X"98",X"76",X"43",X"11",X"11",X"11",
		X"98",X"8D",X"D6",X"FF",X"FF",X"FF",X"00",X"00",X"B9",X"98",X"76",X"43",X"33",X"33",X"1A",X"99",
		X"DD",X"76",X"5F",X"FF",X"FF",X"00",X"0B",X"B9",X"9A",X"D8",X"54",X"44",X"43",X"3A",X"AD",X"D8",
		X"76",X"65",X"FF",X"FF",X"00",X"0B",X"B9",X"AA",X"DD",X"85",X"55",X"54",X"33",X"DD",X"98",X"77",
		X"65",X"FF",X"FF",X"00",X"CB",X"BA",X"AA",X"AE",X"86",X"76",X"65",X"4D",X"D9",X"98",X"77",X"65",
		X"5F",X"FF",X"00",X"BB",X"BA",X"AA",X"AE",X"E8",X"76",X"66",X"DD",X"AA",X"98",X"87",X"66",X"5F",
		X"FF",X"00",X"BB",X"AA",X"AA",X"AA",X"E8",X"77",X"7D",X"DB",X"AA",X"99",X"87",X"76",X"54",X"FF",
		X"0C",X"BB",X"AA",X"AA",X"AA",X"D8",X"88",X"DD",X"CB",X"BA",X"A9",X"88",X"76",X"5D",X"FF",X"0B",
		X"BB",X"AA",X"AA",X"AA",X"DD",X"8D",X"0C",X"CC",X"BA",X"A9",X"88",X"76",X"DD",X"6F",X"0B",X"BA",
		X"AA",X"AA",X"A2",X"2D",X"D0",X"00",X"CC",X"BB",X"A9",X"98",X"7D",X"D7",X"6F",X"0B",X"BA",X"AA",
		X"AA",X"33",X"2D",X"00",X"00",X"0C",X"CB",X"AA",X"98",X"DD",X"87",X"7F",X"CB",X"BA",X"AA",X"A4",
		X"43",X"D0",X"00",X"00",X"0C",X"CB",X"BA",X"9D",X"D9",X"88",X"4F",X"BB",X"AA",X"AA",X"55",X"4D",
		X"00",X"00",X"00",X"00",X"CC",X"BA",X"DD",X"A9",X"93",X"4F",X"BB",X"AA",X"A6",X"65",X"D0",X"00",
		X"00",X"00",X"00",X"CC",X"BD",X"D3",X"AA",X"33",X"4F",X"BB",X"AA",X"77",X"6D",X"00",X"00",X"00",
		X"00",X"00",X"0C",X"DD",X"33",X"33",X"34",X"5F",X"BB",X"A8",X"87",X"D0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"D4",X"44",X"33",X"45",X"5F",X"BB",X"9A",X"8D",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0D",X"54",X"55",X"44",X"55",X"6F",X"CA",X"A9",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"D7",
		X"66",X"65",X"55",X"56",X"6F",X"BC",X"AD",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"77",X"77",
		X"66",X"66",X"66",X"7F",X"0B",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"DD",X"D7",X"67",X"77",
		X"77",X"77",X"8F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"22",X"D8",X"77",X"77",X"77",
		X"77",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D3",X"32",X"DE",X"87",X"77",X"77",X"78",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"44",X"3C",X"CE",X"88",X"77",X"77",X"89",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"D5",X"54",X"CC",X"CE",X"E8",X"88",X"88",X"AF",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"0D",X"66",X"5C",X"CC",X"CC",X"D8",X"88",X"8A",X"9F",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"D7",X"76",X"CC",X"CC",X"CC",X"DD",X"88",X"A9",X"FF",X"FF",X"00",X"00",X"00",
		X"00",X"0D",X"88",X"7C",X"CC",X"CC",X"CC",X"CD",X"AA",X"AF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"D9",X"98",X"CC",X"CC",X"CC",X"CC",X"AA",X"AA",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"0D",X"AA",
		X"9C",X"CC",X"CC",X"CC",X"AA",X"AA",X"AF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"0B",X"BA",X"BB",
		X"BB",X"BB",X"BB",X"BB",X"BF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"BB",X"BB",X"BB",
		X"BB",X"BB",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"88",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"08",X"33",
		X"8F",X"FF",X"FF",X"FF",X"00",X"00",X"08",X"33",X"8F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"88",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"A9",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"09",X"55",
		X"AF",X"FF",X"FF",X"FF",X"00",X"00",X"09",X"55",X"9F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"99",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"88",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"08",X"00",
		X"8F",X"FF",X"FF",X"FF",X"00",X"00",X"08",X"00",X"8F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"88",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"88",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"08",X"33",
		X"8F",X"FF",X"FF",X"FF",X"00",X"00",X"83",X"00",X"38",X"FF",X"FF",X"FF",X"00",X"00",X"83",X"00",
		X"38",X"FF",X"FF",X"FF",X"00",X"00",X"83",X"00",X"38",X"FF",X"FF",X"FF",X"00",X"00",X"83",X"00",
		X"38",X"FF",X"FF",X"FF",X"00",X"00",X"08",X"33",X"8F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"88",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"11",
		X"1F",X"FF",X"FF",X"FF",X"00",X"00",X"11",X"33",X"11",X"FF",X"FF",X"FF",X"00",X"00",X"13",X"33",
		X"31",X"FF",X"FF",X"FF",X"00",X"01",X"13",X"00",X"31",X"1F",X"FF",X"FF",X"00",X"01",X"30",X"00",
		X"03",X"1F",X"FF",X"FF",X"00",X"01",X"30",X"00",X"03",X"1F",X"FF",X"FF",X"00",X"01",X"13",X"00",
		X"31",X"1F",X"FF",X"FF",X"00",X"00",X"13",X"33",X"31",X"FF",X"FF",X"FF",X"00",X"00",X"11",X"33",
		X"11",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"11",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"33",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"33",X"33",
		X"33",X"FF",X"FF",X"FF",X"00",X"03",X"33",X"33",X"33",X"3F",X"FF",X"FF",X"00",X"03",X"30",X"00",
		X"03",X"3F",X"FF",X"FF",X"00",X"33",X"00",X"00",X"00",X"33",X"FF",X"FF",X"00",X"33",X"00",X"00",
		X"00",X"33",X"FF",X"FF",X"00",X"33",X"00",X"00",X"00",X"33",X"FF",X"FF",X"00",X"33",X"00",X"00",
		X"00",X"33",X"FF",X"FF",X"00",X"03",X"30",X"00",X"03",X"3F",X"FF",X"FF",X"00",X"03",X"33",X"33",
		X"33",X"3F",X"FF",X"FF",X"00",X"00",X"33",X"33",X"33",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"33",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"33",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"33",X"33",
		X"33",X"FF",X"FF",X"FF",X"00",X"03",X"38",X"88",X"83",X"3F",X"FF",X"FF",X"00",X"03",X"80",X"00",
		X"08",X"3F",X"FF",X"FF",X"00",X"38",X"00",X"00",X"00",X"83",X"FF",X"FF",X"00",X"38",X"00",X"00",
		X"00",X"83",X"FF",X"FF",X"00",X"38",X"00",X"00",X"00",X"83",X"FF",X"FF",X"00",X"38",X"00",X"00",
		X"00",X"83",X"FF",X"FF",X"00",X"03",X"80",X"00",X"08",X"3F",X"FF",X"FF",X"00",X"03",X"38",X"88",
		X"83",X"3F",X"FF",X"FF",X"00",X"00",X"33",X"33",X"33",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"33",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"88",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"83",X"33",X"38",X"FF",X"FF",X"FF",X"00",X"08",X"30",X"00",
		X"03",X"8F",X"FF",X"FF",X"00",X"83",X"00",X"00",X"00",X"38",X"FF",X"FF",X"00",X"30",X"00",X"00",
		X"00",X"03",X"FF",X"FF",X"08",X"30",X"00",X"11",X"00",X"03",X"8F",X"FF",X"08",X"30",X"01",X"00",
		X"10",X"03",X"8F",X"FF",X"08",X"30",X"01",X"00",X"10",X"03",X"8F",X"FF",X"08",X"30",X"00",X"11",
		X"00",X"03",X"8F",X"FF",X"00",X"30",X"00",X"00",X"00",X"03",X"FF",X"FF",X"00",X"83",X"00",X"00",
		X"00",X"38",X"FF",X"FF",X"00",X"08",X"30",X"00",X"03",X"8F",X"FF",X"FF",X"00",X"00",X"83",X"33",
		X"38",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"88",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"11",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"11",X"11",X"11",X"FF",X"FF",X"FF",X"00",X"01",X"10",X"00",
		X"01",X"1F",X"FF",X"FF",X"00",X"11",X"00",X"00",X"00",X"11",X"FF",X"FF",X"00",X"10",X"00",X"88",
		X"00",X"01",X"FF",X"FF",X"01",X"10",X"08",X"00",X"80",X"01",X"1F",X"FF",X"01",X"10",X"08",X"00",
		X"80",X"01",X"1F",X"FF",X"01",X"10",X"08",X"00",X"80",X"01",X"1F",X"FF",X"01",X"10",X"08",X"00",
		X"80",X"01",X"1F",X"FF",X"00",X"10",X"00",X"88",X"00",X"01",X"FF",X"FF",X"00",X"11",X"00",X"00",
		X"00",X"11",X"FF",X"FF",X"00",X"01",X"10",X"00",X"01",X"1F",X"FF",X"FF",X"00",X"00",X"11",X"11",
		X"11",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"11",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"88",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"88",X"88",
		X"88",X"FF",X"FF",X"FF",X"00",X"08",X"81",X"11",X"18",X"8F",X"FF",X"FF",X"00",X"88",X"10",X"00",
		X"01",X"88",X"FF",X"FF",X"08",X"81",X"00",X"00",X"00",X"18",X"8F",X"FF",X"08",X"10",X"00",X"00",
		X"00",X"11",X"8F",X"FF",X"88",X"10",X"00",X"00",X"00",X"01",X"88",X"FF",X"88",X"10",X"00",X"00",
		X"00",X"01",X"88",X"FF",X"88",X"10",X"00",X"00",X"00",X"01",X"88",X"FF",X"88",X"10",X"00",X"00",
		X"00",X"01",X"88",X"FF",X"08",X"10",X"00",X"00",X"00",X"01",X"8F",X"FF",X"08",X"81",X"00",X"00",
		X"00",X"18",X"8F",X"FF",X"00",X"88",X"10",X"00",X"01",X"88",X"FF",X"FF",X"00",X"08",X"81",X"11",
		X"18",X"8F",X"FF",X"FF",X"00",X"00",X"88",X"88",X"88",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"88",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"88",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"81",X"11",
		X"18",X"FF",X"FF",X"FF",X"00",X"08",X"18",X"88",X"81",X"8F",X"FF",X"FF",X"00",X"81",X"80",X"00",
		X"08",X"18",X"FF",X"FF",X"08",X"18",X"00",X"00",X"00",X"81",X"8F",X"FF",X"01",X"80",X"00",X"00",
		X"00",X"81",X"8F",X"FF",X"81",X"80",X"00",X"00",X"00",X"08",X"18",X"FF",X"81",X"80",X"00",X"00",
		X"00",X"08",X"18",X"FF",X"81",X"80",X"00",X"00",X"00",X"08",X"18",X"FF",X"81",X"80",X"00",X"00",
		X"00",X"08",X"18",X"FF",X"01",X"80",X"00",X"00",X"00",X"08",X"1F",X"FF",X"08",X"18",X"00",X"00",
		X"00",X"81",X"8F",X"FF",X"00",X"81",X"80",X"00",X"08",X"18",X"FF",X"FF",X"00",X"08",X"18",X"88",
		X"81",X"8F",X"FF",X"FF",X"00",X"00",X"81",X"11",X"18",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"88",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"11",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"11",X"88",
		X"11",X"FF",X"FF",X"FF",X"00",X"01",X"88",X"88",X"88",X"1F",X"FF",X"FF",X"00",X"18",X"80",X"00",
		X"08",X"81",X"FF",X"FF",X"01",X"88",X"00",X"00",X"00",X"88",X"1F",X"FF",X"01",X"80",X"00",X"00",
		X"00",X"08",X"1F",X"FF",X"18",X"80",X"00",X"00",X"00",X"08",X"81",X"FF",X"18",X"80",X"00",X"00",
		X"00",X"08",X"81",X"FF",X"18",X"80",X"00",X"00",X"00",X"08",X"81",X"FF",X"18",X"80",X"00",X"00",
		X"00",X"08",X"81",X"FF",X"01",X"80",X"00",X"00",X"00",X"08",X"1F",X"FF",X"01",X"88",X"00",X"00",
		X"00",X"88",X"1F",X"FF",X"00",X"18",X"80",X"00",X"08",X"81",X"FF",X"FF",X"00",X"01",X"88",X"88",
		X"88",X"1F",X"FF",X"FF",X"00",X"00",X"11",X"88",X"11",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"11",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"88",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"88",X"88",
		X"88",X"FF",X"FF",X"FF",X"00",X"08",X"8A",X"AA",X"A8",X"8F",X"FF",X"FF",X"00",X"88",X"A0",X"00",
		X"0A",X"88",X"FF",X"FF",X"08",X"8A",X"00",X"00",X"00",X"A8",X"8F",X"FF",X"08",X"A0",X"00",X"00",
		X"00",X"AA",X"8F",X"FF",X"88",X"A0",X"00",X"00",X"00",X"0A",X"88",X"FF",X"88",X"A0",X"00",X"00",
		X"00",X"0A",X"88",X"FF",X"88",X"A0",X"00",X"00",X"00",X"0A",X"88",X"FF",X"88",X"A0",X"00",X"00",
		X"00",X"0A",X"88",X"FF",X"08",X"A0",X"00",X"00",X"00",X"0A",X"8F",X"FF",X"08",X"8A",X"00",X"00",
		X"00",X"A8",X"8F",X"FF",X"00",X"88",X"A0",X"00",X"0A",X"88",X"FF",X"FF",X"00",X"08",X"8A",X"AA",
		X"A8",X"8F",X"FF",X"FF",X"00",X"00",X"88",X"88",X"88",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"88",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"88",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"8A",X"AA",
		X"A8",X"FF",X"FF",X"FF",X"00",X"08",X"AB",X"BB",X"BA",X"8F",X"FF",X"FF",X"00",X"8A",X"B0",X"00",
		X"0B",X"A8",X"FF",X"FF",X"08",X"AB",X"00",X"00",X"00",X"BA",X"8F",X"FF",X"0A",X"B0",X"00",X"00",
		X"00",X"BB",X"AF",X"FF",X"8A",X"B0",X"00",X"00",X"00",X"0B",X"A8",X"FF",X"8A",X"B0",X"00",X"00",
		X"00",X"0B",X"A8",X"FF",X"8A",X"B0",X"00",X"00",X"00",X"0B",X"A8",X"FF",X"8A",X"B0",X"00",X"00",
		X"00",X"0B",X"A8",X"FF",X"0A",X"B0",X"00",X"00",X"00",X"0B",X"AF",X"FF",X"08",X"AB",X"00",X"00",
		X"00",X"BA",X"8F",X"FF",X"00",X"8A",X"B0",X"00",X"0B",X"A8",X"FF",X"FF",X"00",X"08",X"AB",X"BB",
		X"BA",X"8F",X"FF",X"FF",X"00",X"00",X"8A",X"AA",X"A8",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"88",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"AA",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"AB",X"BB",
		X"BA",X"FF",X"FF",X"FF",X"00",X"0A",X"BC",X"CC",X"CB",X"AF",X"FF",X"FF",X"00",X"AB",X"C0",X"00",
		X"0C",X"BA",X"FF",X"FF",X"0A",X"BC",X"00",X"00",X"00",X"CB",X"AF",X"FF",X"0B",X"C0",X"00",X"00",
		X"00",X"CC",X"BF",X"FF",X"AB",X"C0",X"00",X"00",X"00",X"0C",X"BA",X"FF",X"AB",X"C0",X"00",X"00",
		X"00",X"0C",X"BA",X"FF",X"AB",X"C0",X"00",X"00",X"00",X"0C",X"BA",X"FF",X"AB",X"C0",X"00",X"00",
		X"00",X"0C",X"BA",X"FF",X"0B",X"C0",X"00",X"00",X"00",X"0C",X"BF",X"FF",X"0A",X"BC",X"00",X"00",
		X"00",X"CB",X"AF",X"FF",X"00",X"AB",X"C0",X"00",X"0C",X"BA",X"FF",X"FF",X"00",X"0A",X"BC",X"CC",
		X"CB",X"AF",X"FF",X"FF",X"00",X"00",X"AB",X"BB",X"BA",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"00",X"00",X"AA",X"AA",X"FF",X"FF",X"FF",X"00",X"0A",X"99",X"99",X"AF",X"FF",
		X"FF",X"00",X"A9",X"99",X"88",X"89",X"FF",X"FF",X"0B",X"A9",X"98",X"55",X"58",X"AF",X"FF",X"0A",
		X"99",X"88",X"52",X"56",X"9F",X"FF",X"BA",X"99",X"88",X"52",X"25",X"8A",X"FF",X"AA",X"98",X"65",
		X"53",X"35",X"69",X"FF",X"23",X"45",X"67",X"89",X"AB",X"CD",X"FF",X"23",X"45",X"67",X"89",X"AB",
		X"CD",X"FF",X"23",X"45",X"67",X"89",X"AB",X"CD",X"FF",X"AB",X"BA",X"76",X"54",X"45",X"69",X"FF",
		X"BB",X"BA",X"98",X"55",X"56",X"8A",X"FF",X"0A",X"BA",X"99",X"75",X"56",X"9F",X"FF",X"0B",X"BB",
		X"A9",X"96",X"69",X"AF",X"FF",X"00",X"AB",X"BA",X"A9",X"99",X"FF",X"FF",X"00",X"0A",X"BB",X"AA",
		X"AF",X"FF",X"FF",X"00",X"00",X"BB",X"BB",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"AA",X"AA",X"FF",X"FF",X"FF",X"00",
		X"0A",X"99",X"99",X"AF",X"FF",X"FF",X"00",X"A9",X"99",X"88",X"89",X"FF",X"FF",X"0B",X"A9",X"98",
		X"55",X"58",X"AF",X"FF",X"0A",X"99",X"88",X"52",X"56",X"9F",X"FF",X"BA",X"99",X"88",X"52",X"25",
		X"8A",X"FF",X"AA",X"98",X"65",X"53",X"35",X"69",X"FF",X"87",X"65",X"43",X"21",X"35",X"7B",X"FF",
		X"87",X"65",X"43",X"21",X"35",X"7B",X"FF",X"87",X"65",X"43",X"21",X"35",X"7B",X"FF",X"AB",X"BA",
		X"76",X"54",X"45",X"69",X"FF",X"BB",X"BA",X"98",X"55",X"56",X"8A",X"FF",X"0A",X"BA",X"99",X"75",
		X"56",X"9F",X"FF",X"0B",X"BB",X"A9",X"96",X"69",X"AF",X"FF",X"00",X"AB",X"BA",X"A9",X"99",X"FF",
		X"FF",X"00",X"0A",X"BB",X"AA",X"AF",X"FF",X"FF",X"00",X"00",X"BB",X"BB",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"AA",
		X"AA",X"FF",X"FF",X"FF",X"00",X"0A",X"99",X"99",X"AF",X"FF",X"FF",X"00",X"A9",X"99",X"88",X"89",
		X"FF",X"FF",X"0B",X"A9",X"98",X"55",X"58",X"AF",X"FF",X"0A",X"99",X"88",X"52",X"56",X"9F",X"FF",
		X"BA",X"99",X"88",X"52",X"25",X"8A",X"FF",X"AA",X"98",X"65",X"53",X"35",X"69",X"FF",X"CC",X"BB",
		X"A9",X"87",X"54",X"31",X"FF",X"CC",X"BB",X"A9",X"87",X"54",X"31",X"FF",X"CC",X"BB",X"A9",X"87",
		X"54",X"31",X"FF",X"AB",X"BA",X"76",X"54",X"45",X"69",X"FF",X"BB",X"BA",X"98",X"55",X"56",X"8A",
		X"FF",X"0A",X"BA",X"99",X"75",X"56",X"9F",X"FF",X"0B",X"BB",X"A9",X"96",X"69",X"AF",X"FF",X"00",
		X"AB",X"BA",X"A9",X"99",X"FF",X"FF",X"00",X"0A",X"BB",X"AA",X"AF",X"FF",X"FF",X"00",X"00",X"BB",
		X"BB",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"03",X"30",
		X"FF",X"32",X"13",X"FF",X"31",X"23",X"FF",X"03",X"30",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"10",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"20",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"30",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"40",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"50",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"60",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"70",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"80",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"90",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
