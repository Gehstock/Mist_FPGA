library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_4P is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_4P is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"6E",X"45",X"0B",X"07",X"08",X"09",X"FF",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"0D",X"44",X"0B",X"05",X"09",X"08",X"FF",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"0E",X"10",X"11",X"45",X"03",X"07",X"08",X"09",X"FF",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"12",X"13",X"11",X"44",X"0B",X"05",X"09",X"08",X"FF",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"14",X"15",X"11",X"43",X"0B",X"05",X"08",X"09",X"FF",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"16",X"17",X"11",X"45",X"03",X"04",X"09",X"6D",X"FF",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"18",X"0F",X"11",X"42",X"0A",X"0A",X"0C",X"06",X"FF",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"19",X"1A",X"1B",X"24",X"42",X"0A",X"0A",X"07",X"06",X"FF",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"1C",X"1D",X"1E",X"25",X"42",X"0A",X"0A",X"04",X"06",X"FF",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"1F",X"1D",X"1E",X"25",X"42",X"0A",X"0A",X"05",X"06",X"FF",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"20",X"21",X"22",X"25",X"42",X"0A",X"0A",X"07",X"06",X"FF",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"23",X"45",X"02",X"03",X"07",X"06",X"FF",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"6E",X"44",X"0B",X"0B",X"04",X"06",X"FF",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"6E",X"43",X"0B",X"0B",X"05",X"06",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"08",X"08",X"08",X"08",X"08",X"08",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"08",X"08",X"08",X"08",X"08",X"08",
		X"08",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"88",X"08",X"08",X"08",X"08",X"0A",
		X"08",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"08",X"08",X"08",X"08",X"08",X"0A",
		X"08",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"08",X"08",X"08",X"08",X"08",X"08",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"8A",X"08",X"08",X"08",X"08",X"08",X"08",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"8A",X"08",X"08",X"08",X"08",X"08",X"08",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"08",X"08",X"08",X"08",X"08",X"0A",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"88",X"08",X"08",X"08",X"08",X"08",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"88",X"08",X"08",X"08",X"08",X"08",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"8A",X"08",X"08",X"08",X"08",X"08",X"08",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"08",X"08",X"08",X"08",X"08",X"08",
		X"08",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"88",X"88",X"88",X"08",X"08",X"08",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"8A",X"88",X"08",X"08",X"08",X"08",X"08",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"08",X"08",X"08",X"08",X"08",X"08",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"01",X"71",X"72",X"73",X"74",X"75",X"76",X"3E",X"3F",X"40",X"41",X"4A",X"4C",X"01",X"FF",
		X"FF",X"01",X"71",X"72",X"73",X"74",X"75",X"76",X"3A",X"3B",X"3C",X"3D",X"49",X"01",X"01",X"FF",
		X"FF",X"01",X"71",X"72",X"73",X"74",X"75",X"76",X"36",X"37",X"38",X"39",X"4A",X"01",X"01",X"FF",
		X"FF",X"01",X"71",X"72",X"73",X"74",X"75",X"76",X"32",X"33",X"34",X"35",X"49",X"01",X"4B",X"FF",
		X"FF",X"01",X"71",X"72",X"73",X"74",X"75",X"76",X"2E",X"2F",X"30",X"31",X"46",X"4C",X"01",X"FF",
		X"FF",X"01",X"71",X"72",X"73",X"74",X"75",X"76",X"2A",X"2B",X"2C",X"2D",X"48",X"01",X"01",X"FF",
		X"FF",X"01",X"71",X"72",X"73",X"74",X"75",X"76",X"26",X"27",X"28",X"29",X"47",X"01",X"4C",X"FF",
		X"FF",X"01",X"71",X"72",X"73",X"74",X"75",X"76",X"26",X"27",X"28",X"29",X"47",X"4B",X"01",X"FF",
		X"FF",X"01",X"71",X"72",X"73",X"74",X"75",X"76",X"2A",X"2B",X"2C",X"2D",X"48",X"01",X"01",X"FF",
		X"FF",X"01",X"71",X"72",X"73",X"74",X"75",X"76",X"2E",X"2F",X"30",X"31",X"46",X"01",X"01",X"FF",
		X"FF",X"01",X"71",X"72",X"73",X"74",X"75",X"76",X"32",X"33",X"34",X"35",X"4A",X"4C",X"01",X"FF",
		X"FF",X"01",X"71",X"72",X"73",X"74",X"75",X"76",X"36",X"37",X"38",X"39",X"49",X"01",X"4C",X"FF",
		X"FF",X"01",X"71",X"72",X"73",X"74",X"75",X"76",X"3A",X"3B",X"3C",X"3D",X"4A",X"01",X"01",X"FF",
		X"FF",X"01",X"71",X"72",X"73",X"74",X"75",X"76",X"3E",X"3F",X"40",X"41",X"49",X"01",X"4B",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"80",X"81",X"FF",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"82",X"83",X"84",X"85",X"86",X"81",X"FF",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"8D",X"87",X"88",X"89",X"8A",X"8B",X"8C",X"81",X"FF",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"8E",X"8F",X"90",X"91",X"92",X"C0",X"93",X"94",X"FF",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"95",X"96",X"97",X"98",X"99",X"C1",X"9A",X"9B",X"FF",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"9C",X"9D",X"9E",X"9F",X"A0",X"A1",X"A2",X"A3",X"FF",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"A4",X"AA",X"A5",X"A6",X"A7",X"A8",X"FF",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"A9",X"AA",X"AA",X"AA",X"AB",X"AC",X"A8",X"FF",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"AD",X"AE",X"AA",X"AA",X"AA",X"AF",X"B0",X"B1",X"FF",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"B2",X"B3",X"AE",X"AA",X"AA",X"AA",X"B4",X"B5",X"B1",X"FF",
		X"FF",X"01",X"01",X"01",X"01",X"B6",X"B7",X"B8",X"AE",X"AA",X"AA",X"AA",X"AA",X"B9",X"B1",X"FF",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"BA",X"BB",X"AE",X"AA",X"AA",X"AA",X"AA",X"B9",X"B1",X"FF",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"BC",X"BD",X"AA",X"AA",X"AA",X"AA",X"B9",X"B1",X"FF",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"BE",X"BF",X"AA",X"AA",X"AA",X"B9",X"B1",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"F0",X"F9",X"F8",X"70",X"FC",X"F9",X"FC",X"FF",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"F1",X"70",X"FB",X"F8",X"F9",X"FB",X"F8",X"FF",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"F2",X"F3",X"FE",X"70",X"FB",X"FC",X"FD",X"FF",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"F0",X"FA",X"70",X"FB",X"F9",X"FE",X"FF",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"F4",X"F5",X"F6",X"F8",X"F8",X"FC",X"FF",
		X"FF",X"01",X"01",X"C2",X"C3",X"C4",X"C5",X"C6",X"C7",X"C8",X"C9",X"CA",X"CB",X"F7",X"FD",X"FF",
		X"FF",X"01",X"01",X"CC",X"CD",X"CE",X"CF",X"D0",X"D1",X"D2",X"D3",X"D4",X"D5",X"D6",X"FD",X"FF",
		X"FF",X"01",X"01",X"01",X"01",X"D7",X"D8",X"D9",X"DA",X"DB",X"DC",X"DD",X"DE",X"DF",X"F8",X"FF",
		X"FF",X"01",X"01",X"01",X"E0",X"E1",X"E2",X"E3",X"E4",X"E5",X"E6",X"E7",X"E8",X"E9",X"FB",X"FF",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"EA",X"EB",X"EC",X"ED",X"EE",X"EF",X"FA",X"70",X"FF",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"F4",X"6F",X"F6",X"FB",X"70",X"FA",X"FF",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"F2",X"F3",X"FE",X"F9",X"F8",X"F9",X"FE",X"FF",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"F2",X"F3",X"70",X"FB",X"F8",X"70",X"FC",X"FD",X"FF",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"F1",X"FA",X"F8",X"F9",X"FC",X"FA",X"FB",X"FE",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"8A",X"0A",X"0A",X"8A",X"0A",X"8A",X"0A",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"8A",X"0A",X"0A",X"8A",X"8A",X"0A",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"8A",X"8A",X"0A",X"0A",X"0A",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"8A",X"8A",X"0A",
		X"0A",X"0A",X"0A",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"0A",X"0A",X"0A",X"8A",X"0A",
		X"0A",X"0A",X"0A",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"0A",X"0A",X"0A",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"0A",X"0A",X"0A",
		X"0A",X"0A",X"0A",X"0A",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"01",X"0A",X"8A",X"0A",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"08",X"08",X"08",X"08",X"0A",X"0A",X"8A",X"0A",X"0A",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"8A",X"0A",X"8A",X"8A",X"8A",X"0A",X"0A",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"8A",X"8A",X"0A",X"0A",X"0A",X"8A",X"0A",X"0A",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"8A",X"8A",X"8A",X"8A",X"0A",X"0A",X"0A",X"0A",X"0A",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"8A",X"0A",X"0A",X"0A",X"0A",X"0A",X"8A",X"8A",X"0A",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"55",X"54",X"54",X"54",X"54",X"54",X"53",X"52",X"51",X"FF",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"56",X"57",X"57",X"57",X"58",X"58",X"53",X"52",X"51",X"FF",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"59",X"59",X"53",X"52",X"51",X"FF",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"5B",X"5A",X"5A",X"59",X"59",X"53",X"52",X"51",X"FF",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"59",X"59",X"53",X"52",X"51",X"FF",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"5E",X"5D",X"5C",X"53",X"52",X"51",X"FF",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"5F",X"60",X"53",X"52",X"51",X"FF",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"62",X"61",X"53",X"52",X"51",X"FF",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"63",X"64",X"53",X"52",X"51",X"FF",
		X"FF",X"01",X"01",X"01",X"01",X"65",X"65",X"65",X"65",X"65",X"65",X"65",X"53",X"52",X"51",X"FF",
		X"FF",X"01",X"01",X"01",X"01",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"53",X"52",X"51",X"FF",
		X"FF",X"01",X"01",X"01",X"01",X"67",X"68",X"68",X"68",X"68",X"69",X"6A",X"53",X"52",X"51",X"FF",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"6C",X"6B",X"53",X"52",X"51",X"FF",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"6C",X"6B",X"53",X"52",X"51",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"0A",X"0A",X"0A",X"0A",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"0A",X"0A",X"0A",X"0A",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"0A",X"0A",X"0A",X"0A",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"0A",X"0A",X"0A",X"0A",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"0A",X"0A",X"0A",X"0A",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"0A",X"0A",X"0A",X"0A",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"0A",X"0A",X"0A",X"0A",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"0A",X"0A",X"0A",X"0A",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"0A",X"0A",X"0A",X"0A",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"0A",X"0A",X"0A",X"0A",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"0A",X"0A",X"0A",X"0A",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"0A",X"0A",X"0A",X"0A",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"0A",X"0A",X"0A",X"0A",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"0A",X"0A",X"0A",X"0A",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"07",X"07",X"07",X"07",X"07",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"07",X"07",X"07",X"07",X"07",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"07",X"07",X"07",X"07",X"07",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"07",X"07",X"07",X"07",X"07",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"07",X"07",X"07",X"07",X"07",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"07",X"07",X"07",X"07",X"07",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"07",X"07",X"07",X"07",X"07",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"07",X"07",X"07",X"07",X"07",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"07",X"07",X"07",X"07",X"07",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"07",X"07",X"07",X"07",X"07",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"07",X"07",X"07",X"07",X"07",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"07",X"07",X"07",X"07",X"07",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"07",X"07",X"07",X"07",X"07",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"07",X"07",X"07",X"07",X"07",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"07",X"07",X"07",X"07",X"07",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"07",X"07",X"07",X"07",X"07",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
