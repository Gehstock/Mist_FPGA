library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity travusa_chr_bit3 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of travusa_chr_bit3 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"3F",X"7F",X"70",X"60",X"64",X"6C",X"68",X"00",X"FC",X"FE",X"0E",X"06",X"66",X"F6",X"96",
		X"69",X"6F",X"66",X"60",X"70",X"7F",X"3F",X"00",X"16",X"36",X"26",X"06",X"0E",X"FE",X"FC",X"00",
		X"77",X"67",X"6D",X"7D",X"7B",X"3F",X"1E",X"00",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",
		X"38",X"7D",X"7D",X"6D",X"6F",X"6F",X"67",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"00",X"00",
		X"7F",X"3F",X"00",X"1C",X"3E",X"77",X"63",X"63",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"7F",X"00",X"7D",X"7D",X"00",X"18",X"3B",X"F8",X"F8",X"00",X"80",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BE",X"A0",X"00",X"00",X"00",X"00",
		X"00",X"04",X"04",X"00",X"04",X"04",X"00",X"00",X"28",X"68",X"00",X"40",X"D0",X"00",X"00",X"00",
		X"48",X"C8",X"80",X"AC",X"00",X"94",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"8C",X"80",X"B2",X"A4",X"00",X"00",X"00",X"00",X"06",X"0C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"70",X"C0",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"00",X"00",
		X"00",X"00",X"00",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7E",X"80",X"82",X"82",X"82",X"80",X"00",X"00",X"00",X"00",X"FE",X"80",X"80",X"00",X"00",X"00",
		X"8C",X"98",X"90",X"90",X"B2",X"82",X"82",X"00",X"6C",X"C8",X"80",X"80",X"92",X"82",X"04",X"00",
		X"40",X"DE",X"80",X"80",X"00",X"44",X"58",X"00",X"62",X"C2",X"82",X"82",X"96",X"90",X"90",X"10",
		X"62",X"C2",X"82",X"82",X"96",X"90",X"30",X"00",X"07",X"1C",X"F0",X"80",X"82",X"02",X"06",X"00",
		X"6C",X"C0",X"82",X"82",X"96",X"90",X"20",X"00",X"7C",X"C0",X"82",X"82",X"96",X"90",X"80",X"00",
		X"00",X"00",X"44",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"24",X"64",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0C",X"18",X"B2",X"02",X"06",X"04",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"80",X"80",X"00",X"22",X"22",X"EC",X"00",
		X"6C",X"80",X"92",X"92",X"B6",X"80",X"80",X"00",X"44",X"80",X"82",X"82",X"BE",X"80",X"00",X"00",
		X"7C",X"C0",X"80",X"80",X"82",X"82",X"BE",X"00",X"92",X"92",X"92",X"92",X"B6",X"80",X"80",X"00",
		X"12",X"12",X"12",X"12",X"F6",X"80",X"80",X"00",X"74",X"C4",X"84",X"80",X"92",X"82",X"3C",X"00",
		X"FE",X"00",X"10",X"10",X"F6",X"80",X"80",X"00",X"00",X"00",X"FE",X"80",X"80",X"00",X"00",X"00",
		X"00",X"00",X"7E",X"C0",X"80",X"80",X"80",X"00",X"C2",X"84",X"88",X"00",X"00",X"10",X"F0",X"00",
		X"80",X"80",X"80",X"80",X"BE",X"80",X"80",X"00",X"FC",X"80",X"00",X"FE",X"80",X"00",X"FE",X"00",
		X"FE",X"80",X"80",X"00",X"02",X"02",X"FE",X"00",X"7C",X"80",X"82",X"82",X"BE",X"80",X"00",X"00",
		X"1C",X"20",X"22",X"22",X"EE",X"80",X"80",X"00",X"FC",X"80",X"82",X"82",X"BE",X"80",X"00",X"00",
		X"EC",X"80",X"82",X"02",X"16",X"10",X"F0",X"00",X"60",X"C0",X"84",X"82",X"96",X"90",X"90",X"48",
		X"02",X"02",X"FE",X"80",X"80",X"00",X"02",X"00",X"7E",X"80",X"80",X"80",X"BE",X"80",X"00",X"00",
		X"1E",X"20",X"40",X"C0",X"9E",X"00",X"00",X"00",X"7E",X"80",X"BE",X"80",X"80",X"BE",X"00",X"00",
		X"C2",X"84",X"88",X"00",X"62",X"C0",X"88",X"04",X"0E",X"10",X"E0",X"80",X"86",X"00",X"00",X"00",
		X"87",X"8C",X"98",X"B0",X"A2",X"82",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"7F",X"7F",X"60",X"60",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"DD",X"FF",X"FF",X"FB",X"FF",X"7E",X"FF",X"DF",X"FE",X"FF",X"FF",X"EF",X"7F",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C3",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C3",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FD",X"FB",X"DF",X"FF",X"EE",X"DE",X"FF",X"FF",X"FE",X"FB",X"DF",X"7D",X"F7",X"ED",X"FF",X"FF",
		X"FF",X"F7",X"FF",X"FE",X"D7",X"BE",X"FD",X"5F",X"FE",X"FD",X"BF",X"DF",X"BB",X"F7",X"FD",X"BF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7B",X"FF",X"F6",X"BF",X"FF",X"DB",X"B9",X"FF",X"FF",X"FD",X"7F",X"B7",X"FF",X"FF",X"BB",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C3",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F3",X"20",X"E0",X"90",X"B0",X"78",X"88",X"B0",X"98",
		X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"05",X"1F",X"57",X"FE",X"7D",X"FF",X"DF",X"FB",
		X"62",X"8C",X"7B",X"6B",X"9B",X"76",X"DF",X"ED",X"22",X"1A",X"4D",X"29",X"72",X"85",X"D5",X"78",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0A",X"5A",X"C5",X"63",X"5A",X"A1",X"1F",X"FB",
		X"44",X"1A",X"D6",X"83",X"29",X"70",X"95",X"86",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",
		X"7E",X"3B",X"1F",X"07",X"01",X"00",X"00",X"00",X"FF",X"7F",X"FD",X"AF",X"BB",X"7B",X"1F",X"07",
		X"51",X"B6",X"42",X"D9",X"95",X"46",X"F1",X"90",X"80",X"C0",X"60",X"20",X"80",X"30",X"B8",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"34",X"6C",X"C0",X"18",X"D2",X"86",X"3B",X"E9",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"C0",X"80",X"60",X"20",X"F0",X"A0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"F7",X"FE",X"FF",X"FB",X"FF",X"DF",X"FF",
		X"FF",X"00",X"38",X"7D",X"7D",X"38",X"00",X"FF",X"FF",X"80",X"8E",X"9B",X"9F",X"8E",X"80",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"0F",X"1F",X"7C",X"F8",X"E0",
		X"FF",X"FF",X"FF",X"07",X"00",X"00",X"00",X"00",X"FF",X"3F",X"1F",X"08",X"00",X"00",X"00",X"00",
		X"00",X"80",X"E0",X"E0",X"60",X"70",X"18",X"1C",X"E0",X"83",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"0F",X"1F",X"7C",X"F8",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"0F",X"1F",
		X"7C",X"F8",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"10",X"00",X"0C",X"02",X"01",X"00",X"00",X"00",X"00",X"20",X"88",X"E5",X"F8",X"FF",X"FF",
		X"F8",X"FE",X"FF",X"FF",X"0F",X"0F",X"03",X"01",X"07",X"1F",X"01",X"01",X"00",X"00",X"00",X"00",
		X"1F",X"7C",X"F8",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"0F",X"1F",X"7C",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"60",X"80",X"00",X"00",X"00",X"00",X"80",X"E0",X"78",
		X"C8",X"98",X"64",X"2C",X"C1",X"85",X"AF",X"EE",X"F8",X"E0",X"80",X"00",X"00",X"00",X"E0",X"F0",
		X"00",X"03",X"0F",X"1F",X"7C",X"F8",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"0F",
		X"0F",X"1F",X"7C",X"F8",X"E0",X"80",X"04",X"02",X"38",X"08",X"0E",X"02",X"03",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"E0",X"3C",X"07",X"18",X"D5",X"60",X"2A",X"CF",X"9D",X"03",X"3D",
		X"06",X"04",X"01",X"03",X"03",X"0F",X"1F",X"7C",X"C0",X"E0",X"78",X"B8",X"D8",X"EC",X"F7",X"FB",
		X"FF",X"01",X"E1",X"F1",X"F1",X"E1",X"01",X"FF",X"FF",X"7F",X"3F",X"3F",X"7F",X"FF",X"FF",X"FF",
		X"FF",X"BF",X"9F",X"FF",X"EF",X"F7",X"F9",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"1F",X"87",X"E0",X"FC",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"0F",
		X"77",X"F5",X"A0",X"86",X"34",X"21",X"1B",X"08",X"04",X"07",X"02",X"00",X"03",X"0F",X"1F",X"7C",
		X"24",X"7A",X"B7",X"DF",X"EF",X"99",X"1D",X"1F",X"00",X"03",X"0F",X"1F",X"7C",X"F8",X"E0",X"80",
		X"00",X"00",X"03",X"0F",X"1F",X"7C",X"F8",X"E0",X"F8",X"E0",X"83",X"02",X"00",X"01",X"01",X"00",
		X"FF",X"FF",X"7F",X"3F",X"3F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"03",X"0F",X"1F",X"7C",X"F8",
		X"1F",X"7C",X"F8",X"E0",X"80",X"00",X"00",X"00",X"00",X"0C",X"0C",X"0C",X"04",X"04",X"04",X"04",
		X"00",X"00",X"00",X"00",X"00",X"03",X"0F",X"1F",X"03",X"0F",X"1F",X"7C",X"F8",X"E0",X"80",X"00",
		X"E0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"06",X"06",X"06",X"06",X"06",X"06",X"06",
		X"7C",X"F8",X"E0",X"80",X"00",X"00",X"40",X"40",X"00",X"00",X"00",X"04",X"04",X"04",X"06",X"06",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"80",X"80",X"C1",X"07",X"1F",X"3E",X"F8",X"F0",
		X"0F",X"0F",X"0F",X"0F",X"0E",X"08",X"00",X"01",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",
		X"E0",X"E0",X"E0",X"60",X"60",X"60",X"60",X"60",X"FB",X"FD",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"BF",X"BF",X"BF",X"BF",X"BF",X"FF",X"FF",X"FF",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F8",X"F0",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",X"FB",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"07",X"07",X"07",X"07",X"0F",X"1F",X"1F",X"3F",
		X"60",X"60",X"60",X"60",X"70",X"70",X"78",X"3C",X"0F",X"0F",X"0F",X"07",X"07",X"07",X"07",X"07",
		X"00",X"00",X"00",X"00",X"40",X"40",X"40",X"40",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"0F",
		X"20",X"10",X"30",X"38",X"10",X"00",X"00",X"00",X"FF",X"FF",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F8",X"F8",X"00",X"00",X"02",X"02",X"04",X"00",X"00",X"08",
		X"FF",X"FC",X"F3",X"4F",X"FF",X"FF",X"FF",X"FF",X"E1",X"83",X"3F",X"FF",X"FF",X"FF",X"3F",X"FF",
		X"FF",X"C3",X"10",X"FE",X"FF",X"FF",X"FF",X"FF",X"FB",X"C2",X"00",X"39",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",X"21",X"4C",X"67",X"DF",X"FF",X"FF",X"BF",X"24",X"C0",X"F8",
		X"FF",X"FF",X"FF",X"FF",X"7F",X"BF",X"43",X"0C",X"FF",X"FA",X"FF",X"FF",X"FF",X"FF",X"7D",X"FF",
		X"FF",X"FF",X"FF",X"7F",X"9F",X"EF",X"F7",X"FB",X"7F",X"9F",X"E3",X"FB",X"F8",X"FE",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"7F",X"1F",X"CF",X"E7",X"FF",X"7F",X"1F",X"DF",X"EF",X"F3",X"FD",X"FE",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E0",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"1F",X"03",X"C0",X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"00",X"00",X"80",X"FC",X"FF",
		X"FF",X"FF",X"FF",X"1F",X"03",X"07",X"1F",X"FF",X"1F",X"C7",X"F3",X"F9",X"FC",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"7F",X"1F",X"C7",X"F1",X"3F",X"07",X"C0",X"F8",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"80",X"F8",X"FF",X"FF",X"FF",X"FF",X"7F",X"07",X"00",X"00",X"80",X"FC",
		X"FF",X"FF",X"FF",X"F0",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"FE",X"FE",X"FE",X"FC",X"F0",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"06",X"9E",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"F0",X"F0",X"FF",X"FF",X"FF",X"FF",X"F0",X"F0",X"F0",X"F0",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"FF",X"FF",X"FF",X"FF",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"DE",X"CF",X"C7",X"C3",X"E1",X"F0",X"F8",
		X"FF",X"BF",X"81",X"BF",X"FF",X"A1",X"8D",X"FF",X"FF",X"87",X"B7",X"81",X"FF",X"81",X"BD",X"81",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"D6",X"B9",X"D2",X"C8",X"A0",X"00",
		X"FF",X"7F",X"9F",X"2F",X"0B",X"26",X"88",X"00",X"FF",X"FF",X"EF",X"FB",X"D7",X"EB",X"85",X"00",
		X"00",X"01",X"2B",X"05",X"5F",X"AE",X"5D",X"F7",X"00",X"20",X"E9",X"50",X"B2",X"E5",X"FA",X"AF",
		X"00",X"81",X"51",X"AB",X"D6",X"77",X"DD",X"B6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E3",X"C0",X"DF",X"D7",X"F0",X"C0",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"BF",X"BF",X"3F",X"00",
		X"FF",X"FF",X"BF",X"FF",X"FF",X"FF",X"FF",X"03",X"C7",X"0F",X"FF",X"F9",X"01",X"03",X"FF",X"FF",
		X"93",X"80",X"80",X"81",X"C0",X"80",X"81",X"A0",X"80",X"81",X"FF",X"FF",X"FF",X"00",X"00",X"42",
		X"42",X"42",X"42",X"3C",X"42",X"42",X"42",X"42",X"00",X"44",X"88",X"22",X"22",X"88",X"44",X"00",
		X"00",X"00",X"28",X"42",X"28",X"B4",X"7E",X"FF",X"FF",X"3E",X"6A",X"B4",X"21",X"08",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"F0",X"FF",X"F0",X"E0",X"E0",X"C4",X"00",X"03",X"02",
		X"F0",X"E4",X"E5",X"EF",X"C7",X"83",X"91",X"94",X"A3",X"97",X"E7",X"EF",X"EF",X"EF",X"FF",X"FF",
		X"FF",X"D1",X"C0",X"D0",X"98",X"90",X"00",X"00",X"61",X"21",X"21",X"01",X"01",X"01",X"01",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"07",X"0F",X"4F",X"FF",X"FF",X"FF",
		X"8F",X"83",X"81",X"80",X"80",X"80",X"C0",X"C0",X"FF",X"F7",X"45",X"06",X"3E",X"38",X"10",X"00",
		X"C0",X"E0",X"F8",X"EC",X"FC",X"FD",X"FB",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",
		X"0F",X"8F",X"C3",X"C3",X"83",X"E1",X"F1",X"E1",X"F6",X"4D",X"ED",X"EF",X"9A",X"B6",X"75",X"DD",
		X"F7",X"EF",X"FF",X"FF",X"7F",X"FF",X"FF",X"DF",X"FF",X"FF",X"FB",X"FF",X"77",X"FF",X"FF",X"DF",
		X"00",X"1F",X"20",X"40",X"08",X"18",X"10",X"15",X"00",X"FF",X"00",X"00",X"00",X"00",X"10",X"67",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"08",X"DC",X"00",X"FF",X"00",X"00",X"00",X"00",X"10",X"35",
		X"00",X"F8",X"0C",X"06",X"02",X"02",X"02",X"02",X"12",X"11",X"11",X"13",X"15",X"10",X"11",X"12",
		X"82",X"02",X"02",X"02",X"82",X"82",X"02",X"82",X"13",X"15",X"10",X"08",X"07",X"00",X"00",X"00",
		X"8B",X"51",X"02",X"00",X"FF",X"00",X"00",X"00",X"CC",X"29",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"D3",X"91",X"01",X"00",X"FF",X"00",X"00",X"00",X"02",X"82",X"02",X"22",X"C6",X"0C",X"18",X"10",
		X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"C3",X"3C",X"3C",X"3C",
		X"FF",X"E0",X"C0",X"80",X"80",X"81",X"82",X"84",X"FF",X"07",X"03",X"01",X"01",X"81",X"41",X"21",
		X"FF",X"1F",X"03",X"00",X"60",X"F8",X"00",X"CF",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"1F",X"0F",
		X"72",X"FD",X"FA",X"FE",X"F9",X"FD",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"98",X"B9",X"FD",X"FF",
		X"00",X"00",X"00",X"04",X"95",X"BF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"43",X"EF",X"FF",
		X"FF",X"FF",X"CF",X"97",X"70",X"E8",X"BD",X"17",X"FF",X"FF",X"FF",X"FF",X"00",X"81",X"7A",X"AC",
		X"FF",X"FF",X"FF",X"FF",X"16",X"44",X"6A",X"99",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"E0",X"FF",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"03",X"FF",
		X"EF",X"7F",X"FB",X"BE",X"FD",X"EF",X"FB",X"5B",X"00",X"EF",X"10",X"10",X"10",X"10",X"EF",X"00",
		X"00",X"FC",X"06",X"0A",X"12",X"22",X"82",X"42",X"42",X"00",X"00",X"FF",X"FF",X"E7",X"C3",X"83",
		X"C1",X"E1",X"C0",X"80",X"81",X"C3",X"C7",X"C0",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",
		X"00",X"DA",X"92",X"DA",X"52",X"52",X"DA",X"00",X"00",X"CA",X"AA",X"CA",X"AA",X"AA",X"CE",X"00",
		X"00",X"A4",X"AA",X"AA",X"CA",X"AE",X"AA",X"00",X"00",X"A9",X"AA",X"AA",X"BA",X"AB",X"AA",X"00",
		X"00",X"3B",X"92",X"93",X"91",X"91",X"93",X"00",X"00",X"51",X"51",X"51",X"55",X"51",X"71",X"00",
		X"00",X"4B",X"6A",X"6A",X"5A",X"5A",X"4B",X"00",X"C0",X"81",X"0F",X"08",X"00",X"00",X"00",X"80",
		X"C1",X"80",X"30",X"30",X"30",X"00",X"00",X"71",X"C0",X"81",X"0F",X"01",X"80",X"F0",X"81",X"03",
		X"C1",X"80",X"30",X"30",X"30",X"30",X"41",X"83",X"8F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"01",
		X"E3",X"C3",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"81",X"00",X"00",X"30",X"30",X"30",X"30",X"71",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"03",X"1F",X"E3",X"00",X"00",X"05",X"BF",
		X"00",X"00",X"00",X"00",X"0F",X"70",X"80",X"00",X"38",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EF",X"FD",X"BF",X"F6",X"40",X"40",X"00",X"07",X"F7",X"FA",X"C0",X"00",X"01",X"0E",X"F0",X"00",
		X"80",X"00",X"07",X"38",X"C0",X"00",X"00",X"00",X"3F",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"B7",X"FF",X"EE",X"B2",X"40",X"0C",X"3C",
		X"F7",X"F7",X"FA",X"40",X"00",X"00",X"0F",X"F0",X"D7",X"A0",X"00",X"00",X"0F",X"F0",X"00",X"00",
		X"00",X"00",X"0F",X"F0",X"00",X"00",X"00",X"00",X"0F",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"F3",X"BE",X"F9",X"9F",X"F7",
		X"FF",X"3F",X"3C",X"0C",X"80",X"E1",X"B7",X"FE",X"C0",X"FF",X"3F",X"00",X"00",X"80",X"69",X"FF",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"B5",X"00",X"00",X"00",X"00",X"F8",X"7C",X"7A",X"01",
		X"F8",X"C0",X"C0",X"C3",X"17",X"FD",X"FF",X"DF",X"00",X"06",X"4F",X"77",X"BD",X"FF",X"FF",X"FB",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"01",X"0E",X"F0",X"00",
		X"00",X"00",X"07",X"38",X"C0",X"00",X"02",X"1F",X"0E",X"F0",X"00",X"00",X"05",X"67",X"FE",X"DF",
		X"00",X"03",X"13",X"7F",X"BF",X"FB",X"DF",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"07",X"78",X"C0",X"00",X"00",X"00",X"0F",X"FC",X"3C",X"30",X"07",
		X"00",X"0F",X"F0",X"00",X"00",X"06",X"67",X"7F",X"F0",X"00",X"00",X"02",X"AE",X"7B",X"DF",X"FF",
		X"00",X"04",X"5F",X"FF",X"FF",X"FF",X"BF",X"FB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"F0",X"00",X"00",X"00",X"00",X"0F",X"F0",X"00",X"00",X"05",
		X"00",X"0F",X"FC",X"3C",X"30",X"02",X"CF",X"7E",X"3F",X"C0",X"00",X"00",X"12",X"DF",X"AF",X"FD",
		X"00",X"00",X"00",X"5C",X"FB",X"FF",X"B7",X"FE",X"F0",X"00",X"4A",X"FF",X"EF",X"FF",X"DB",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"F4",X"41",X"C0",X"C8",X"B8",X"B2",X"EF",X"7F",X"FB",
		X"C0",X"3C",X"03",X"00",X"80",X"E8",X"ED",X"B9",X"00",X"00",X"E0",X"1F",X"00",X"00",X"40",X"ED",
		X"00",X"00",X"00",X"80",X"7F",X"3C",X"3C",X"80",X"48",X"24",X"66",X"76",X"EE",X"66",X"25",X"53",
		X"40",X"30",X"18",X"1C",X"8D",X"40",X"D0",X"FC",X"00",X"00",X"00",X"00",X"80",X"60",X"18",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C2",X"E1",X"F0",X"68",X"EC",X"FA",X"BF",X"F7",
		X"00",X"00",X"80",X"60",X"10",X"0C",X"02",X"C1",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"C2",X"A1",X"F3",X"69",X"F8",X"EA",X"FC",X"BF",X"00",X"00",X"80",X"C0",X"A0",X"10",X"08",X"84",
		X"07",X"81",X"C0",X"F0",X"74",X"FE",X"FC",X"EF",X"00",X"00",X"80",X"40",X"20",X"10",X"08",X"04",
		X"84",X"D0",X"FC",X"FA",X"EF",X"BE",X"FF",X"EF",X"60",X"10",X"0C",X"82",X"C1",X"E0",X"A8",X"F8",
		X"00",X"00",X"00",X"00",X"80",X"40",X"30",X"08",X"BF",X"FB",X"EE",X"FE",X"BF",X"FB",X"7D",X"F6",
		X"3C",X"00",X"08",X"EF",X"EE",X"FF",X"BA",X"AF",X"0F",X"00",X"00",X"60",X"B5",X"FE",X"FF",X"EF",
		X"00",X"E0",X"1C",X"03",X"00",X"20",X"70",X"FD",X"00",X"00",X"00",X"80",X"60",X"38",X"3E",X"1D",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"AB",X"CA",X"7D",X"B7",X"DB",X"4A",X"FE",X"65",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"3D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"3C",X"3C",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"6F",X"5F",X"EF",X"8F",X"DF",X"9F",X"7F",X"3F",
		X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F7",X"FB",X"FB",X"FF",X"EF",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"9F",X"1F",X"2F",X"2F",
		X"FF",X"FF",X"FE",X"FC",X"FB",X"FC",X"FF",X"FE",X"1F",X"07",X"8F",X"87",X"CB",X"4E",X"47",X"4F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"F1",X"F0",X"C0",X"C0",X"81",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E1",X"F1",X"FF",X"F4",X"FC",X"E7",X"E7",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0C",X"08",X"30",X"30",X"08",X"0C",X"00",X"00",X"00",X"01",X"03",X"03",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"1C",X"18",X"0C",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"1C",X"18",X"04",X"10",X"00",
		X"00",X"00",X"00",X"20",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"03",X"0F",X"1F",X"3F",X"3F",X"7F",X"7F",X"FF",X"C0",X"F0",X"F8",X"FC",X"FC",X"FE",X"FE",X"FF",
		X"FF",X"7F",X"7F",X"3F",X"3F",X"1F",X"0F",X"03",X"FF",X"FE",X"FE",X"FC",X"FC",X"F8",X"F0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"71",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"40",
		X"00",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"00",X"8E",X"8E",X"8E",X"8E",X"8E",X"8E",X"8E",
		X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"00",X"8E",X"8E",X"8E",X"8E",X"8E",X"8E",X"8E",X"00",
		X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"8E",X"8E",X"8E",X"8E",X"8E",X"8E",X"8E",X"8E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"1E",X"3C",X"1E",X"08",X"00",
		X"00",X"00",X"00",X"60",X"71",X"70",X"60",X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"00",X"00",
		X"00",X"00",X"30",X"71",X"71",X"71",X"71",X"70",X"00",X"00",X"40",X"40",X"00",X"00",X"40",X"40",
		X"00",X"00",X"00",X"01",X"03",X"07",X"0F",X"1F",X"00",X"00",X"80",X"C0",X"E0",X"F0",X"F8",X"FC",
		X"3F",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"FE",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"00",X"FF",X"00",X"FF",X"00",X"00",
		X"FF",X"91",X"00",X"6E",X"6E",X"00",X"91",X"FF",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",
		X"FD",X"A5",X"95",X"FD",X"A5",X"95",X"FD",X"C5",X"B7",X"FF",X"97",X"87",X"FF",X"87",X"CF",X"87",
		X"AD",X"C5",X"FD",X"F5",X"85",X"FD",X"B5",X"85",X"FF",X"87",X"AF",X"C7",X"FF",X"C7",X"BF",X"87",
		X"FD",X"95",X"05",X"6D",X"05",X"05",X"FD",X"55",X"05",X"FD",X"4D",X"45",X"15",X"95",X"FD",X"05",
		X"55",X"05",X"05",X"FD",X"3D",X"0D",X"E5",X"0D",X"05",X"CD",X"9D",X"05",X"05",X"FD",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"FF",X"97",X"87",X"FF",X"07",X"FF",X"87",
		X"FD",X"AD",X"AD",X"FD",X"FD",X"55",X"55",X"05",X"B7",X"CF",X"FF",X"C7",X"BF",X"87",X"BF",X"87",
		X"3D",X"FD",X"05",X"05",X"FD",X"95",X"05",X"6D",X"05",X"05",X"FD",X"75",X"75",X"05",X"8D",X"FD",
		X"05",X"05",X"FD",X"8D",X"05",X"75",X"05",X"05",X"05",X"05",X"FD",X"F5",X"F5",X"05",X"05",X"FD",
		X"FF",X"81",X"00",X"7E",X"7E",X"00",X"81",X"FF",X"7F",X"3F",X"9F",X"CF",X"E7",X"FF",X"A7",X"CF",
		X"FF",X"9E",X"0E",X"6E",X"6E",X"60",X"70",X"FF",X"97",X"FF",X"97",X"87",X"FF",X"47",X"17",X"FF",
		X"F0",X"F7",X"F4",X"F7",X"F4",X"F6",X"F5",X"F4",X"00",X"FF",X"12",X"D5",X"1F",X"B0",X"5E",X"17",
		X"F7",X"F4",X"F7",X"F5",X"F4",X"F7",X"F5",X"F4",X"F0",X"1F",X"F0",X"56",X"1F",X"F0",X"19",X"50",
		X"00",X"FF",X"CF",X"CB",X"88",X"FB",X"CC",X"CB",X"0F",X"EF",X"AF",X"EF",X"2F",X"EF",X"EF",X"6F",
		X"88",X"CF",X"8A",X"F8",X"8F",X"9C",X"EB",X"88",X"2F",X"EF",X"AF",X"2F",X"EF",X"6F",X"AF",X"2F",
		X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"07",X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"F8",X"F8",X"F8",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"13",X"7F",X"13",X"00",X"00",X"00",X"00",X"00",X"40",X"C0",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"73",X"73",X"72",X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"40",
		X"00",X"00",X"30",X"70",X"71",X"73",X"72",X"32",X"00",X"00",X"40",X"40",X"40",X"00",X"00",X"00",
		X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",
		X"00",X"00",X"73",X"72",X"00",X"00",X"73",X"72",X"00",X"00",X"40",X"40",X"00",X"00",X"40",X"40",
		X"00",X"00",X"30",X"70",X"70",X"70",X"73",X"32",X"00",X"00",X"40",X"40",X"00",X"00",X"40",X"40",
		X"00",X"00",X"60",X"60",X"73",X"72",X"60",X"60",X"00",X"00",X"00",X"00",X"40",X"40",X"00",X"00",
		X"00",X"00",X"33",X"73",X"71",X"71",X"73",X"32",X"00",X"00",X"40",X"40",X"00",X"00",X"40",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"31",X"71",X"70",X"70",X"73",X"32",X"00",X"00",X"40",X"40",X"00",X"00",X"40",X"40",
		X"00",X"00",X"73",X"73",X"01",X"03",X"73",X"72",X"00",X"00",X"40",X"40",X"40",X"00",X"40",X"40",
		X"00",X"00",X"33",X"72",X"70",X"70",X"73",X"32",X"00",X"00",X"40",X"40",X"00",X"00",X"40",X"40",
		X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"22",X"36",X"7E",X"FC",X"BC",X"4E",X"36",X"22",
		X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"40",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"F9",X"F8",X"BC",X"F0",X"FC",X"F9",X"F2",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"07",X"00",X"00",X"00",X"00",X"7F",X"FF",X"FF",X"FE",
		X"0F",X"1F",X"1F",X"1F",X"3F",X"3F",X"3F",X"3F",X"FE",X"FC",X"FA",X"FE",X"FE",X"FC",X"FC",X"F9",
		X"00",X"00",X"00",X"00",X"FC",X"43",X"7F",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"F8",
		X"00",X"00",X"00",X"00",X"40",X"6E",X"3A",X"01",X"20",X"0C",X"46",X"82",X"02",X"00",X"48",X"44",
		X"3F",X"3F",X"3F",X"3F",X"1F",X"1F",X"1F",X"0F",X"FF",X"FE",X"FC",X"F8",X"FC",X"FE",X"FF",X"FF",
		X"0F",X"07",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"3F",X"00",X"00",X"00",X"00",
		X"01",X"20",X"42",X"00",X"18",X"1C",X"0E",X"06",X"44",X"48",X"00",X"02",X"82",X"44",X"08",X"3C",
		X"C1",X"FF",X"C3",X"F8",X"00",X"00",X"00",X"00",X"F0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F7",X"F0",X"F4",X"F4",X"F4",X"F4",X"F4",X"F4",X"FF",X"00",X"FF",X"FF",X"F8",X"E0",X"C0",X"83",
		X"F4",X"F4",X"F4",X"F4",X"F4",X"F4",X"F4",X"F0",X"87",X"83",X"C0",X"E0",X"F8",X"FF",X"FF",X"00",
		X"FF",X"00",X"FF",X"FF",X"01",X"01",X"01",X"CF",X"EF",X"0F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",
		X"CF",X"CF",X"01",X"01",X"01",X"FF",X"FF",X"00",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"0F",
		X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"FF",X"FB",X"00",X"00",X"7B",X"03",X"83",X"FF",
		X"B8",X"B8",X"B8",X"BF",X"BF",X"B8",X"B8",X"B8",X"0F",X"07",X"03",X"E3",X"E3",X"03",X"07",X"0F",
		X"BF",X"BF",X"BE",X"BE",X"BE",X"A0",X"A0",X"A0",X"FF",X"07",X"03",X"03",X"73",X"03",X"03",X"03",
		X"BF",X"B7",X"A2",X"A2",X"A2",X"B7",X"BF",X"BC",X"FF",X"FF",X"03",X"03",X"03",X"FF",X"8F",X"C7",
		X"B8",X"B8",X"B9",X"B9",X"B8",X"BC",X"BE",X"BF",X"63",X"33",X"13",X"83",X"C3",X"07",X"0F",X"FF",
		X"B3",X"A3",X"A3",X"A6",X"A6",X"A0",X"A0",X"B0",X"87",X"03",X"03",X"33",X"33",X"63",X"63",X"E7",
		X"3F",X"FF",X"F0",X"80",X"23",X"3F",X"9F",X"8F",X"E0",X"F8",X"78",X"1C",X"0C",X"CC",X"E4",X"F4",
		X"C7",X"E0",X"F0",X"60",X"21",X"03",X"E7",X"FF",X"F4",X"54",X"10",X"00",X"80",X"80",X"C0",X"E0",
		X"EF",X"EF",X"E7",X"E2",X"F0",X"F9",X"FF",X"CF",X"F0",X"E0",X"E0",X"40",X"00",X"00",X"C0",X"E0",
		X"E3",X"7F",X"3F",X"3E",X"00",X"00",X"00",X"00",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",X"FF",X"F1",X"60",X"6E",X"6E",X"00",X"81",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"8F",X"07",X"77",X"77",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"36",X"3C",X"18",X"10",X"00",X"00",X"00",X"00",
		X"86",X"C2",X"42",X"62",X"26",X"3C",X"10",X"00",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",
		X"11",X"18",X"F8",X"38",X"01",X"01",X"83",X"FE",X"0C",X"87",X"C1",X"60",X"30",X"1C",X"07",X"00",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"FC",X"FC",X"FC",X"00",X"00",X"00",X"00",X"0F",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"20",X"00",X"40",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"81",X"01",X"22",
		X"80",X"C0",X"60",X"30",X"10",X"18",X"0C",X"84",X"81",X"E0",X"30",X"18",X"0C",X"06",X"03",X"01",
		X"43",X"46",X"44",X"66",X"22",X"23",X"31",X"11",X"00",X"80",X"80",X"C0",X"40",X"60",X"30",X"18",
		X"11",X"11",X"18",X"08",X"08",X"0C",X"04",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"0F",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"03",X"00",X"00",X"00",X"00",
		X"3F",X"3F",X"BF",X"BF",X"3F",X"00",X"00",X"00",X"03",X"01",X"81",X"FF",X"F0",X"1C",X"06",X"03",
		X"00",X"E0",X"3F",X"00",X"0F",X"38",X"20",X"60",X"F8",X"0F",X"00",X"E0",X"20",X"20",X"20",X"E0",
		X"03",X"00",X"00",X"07",X"0C",X"18",X"10",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"F0",X"00",X"00",X"00",X"00",X"00",X"C0",X"7E",
		X"8F",X"80",X"C0",X"40",X"40",X"70",X"1F",X"00",X"18",X"08",X"08",X"0C",X"FC",X"04",X"00",X"00",
		X"00",X"00",X"00",X"7F",X"41",X"40",X"60",X"3E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"1F",X"0F",X"07",X"03",X"01",X"C1",X"FF",X"E0",X"C0",X"80",X"80",X"80",X"F0",X"FF",X"FF",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"00",X"00",X"00",X"00",X"C0",X"60",X"20",X"30",
		X"06",X"FC",X"00",X"FC",X"07",X"00",X"00",X"F8",X"FC",X"C7",X"7F",X"01",X"00",X"80",X"F0",X"11",
		X"F9",X"0F",X"00",X"80",X"F0",X"1F",X"00",X"00",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"A0",X"90",X"45",X"C3",X"83",X"51",X"78",
		X"F8",X"E0",X"D4",X"DE",X"CE",X"07",X"17",X"CF",X"DC",X"EE",X"76",X"7F",X"7F",X"3F",X"9F",X"9F",
		X"7F",X"BD",X"94",X"41",X"80",X"80",X"C0",X"E2",X"5F",X"BF",X"DF",X"BF",X"CE",X"FE",X"E7",X"FE",
		X"F3",X"EA",X"F1",X"F8",X"F8",X"60",X"70",X"28",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"BF",X"BF",X"3F",X"2F",X"7E",X"6E",X"E4",X"EE",X"0C",X"18",X"78",X"78",X"41",X"C3",X"F2",X"64",
		X"CC",X"BC",X"F8",X"F0",X"F3",X"8E",X"FD",X"FF",X"C5",X"CB",X"0F",X"9F",X"3F",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"F0",X"C7",X"1F",X"7F",
		X"FC",X"F9",X"E3",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"1F",X"03",X"0C",X"1F",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"80",X"00",
		X"1F",X"00",X"00",X"1F",X"00",X"0F",X"1F",X"10",X"80",X"02",X"83",X"9F",X"10",X"10",X"90",X"90",
		X"0F",X"00",X"13",X"1F",X"0C",X"00",X"1F",X"11",X"10",X"10",X"10",X"90",X"9F",X"00",X"80",X"00",
		X"0F",X"00",X"13",X"10",X"1F",X"0F",X"00",X"00",X"80",X"00",X"80",X"80",X"80",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"0F",X"E7",X"F3",X"FB",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"F9",X"FD",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"01",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"C1",X"FC",
		X"FF",X"FF",X"FF",X"FF",X"0F",X"E0",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"E0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"FE",X"FE",X"FC",X"FD",X"F9",X"FB",X"F3",X"F7",
		X"C1",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"C1",X"FC",X"FF",X"FF",X"FF",X"FF",
		X"F7",X"F7",X"F7",X"F7",X"07",X"FF",X"77",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"07",X"77",X"77",X"07",X"07",X"77",X"77",X"07",X"01",X"01",X"01",X"01",X"00",X"01",X"01",X"01",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"0F",
		X"0F",X"0F",X"1F",X"1F",X"00",X"1F",X"1F",X"0F",X"03",X"03",X"07",X"07",X"87",X"E7",X"FF",X"FF",
		X"7E",X"7E",X"7E",X"7E",X"7F",X"7F",X"7F",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"0F",X"0F",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FB",X"FC",X"D0",X"E0",X"40",X"C0",X"80",X"80",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"FF",X"FF",X"FF",X"FF",X"C7",X"01",X"00",X"00",
		X"FC",X"F8",X"F8",X"F8",X"F0",X"F0",X"F1",X"F1",X"00",X"00",X"38",X"7C",X"FE",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"3F",X"3F",X"1F",X"0F",X"07",X"83",X"C3",X"FF",X"FF",X"FF",X"FF",X"FF",X"8F",X"07",X"07",
		X"F1",X"F1",X"F0",X"F8",X"F8",X"F8",X"FC",X"FC",X"FF",X"FF",X"FF",X"FF",X"7F",X"33",X"01",X"01",
		X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"01",X"03",X"C7",X"FF",X"FF",X"FF",X"FF",
		X"E3",X"F3",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"07",X"07",X"8F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"0F",X"0F",X"1F",X"3E",X"04",X"60",X"73",
		X"01",X"00",X"00",X"01",X"00",X"07",X"8F",X"8F",X"FE",X"EE",X"C6",X"C6",X"46",X"06",X"82",X"C2",
		X"C7",X"E0",X"F0",X"60",X"21",X"03",X"E7",X"FF",X"E2",X"42",X"02",X"02",X"82",X"82",X"C2",X"E2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"7F",X"67",X"01",X"01",X"04",X"07",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EF",X"EF",X"E7",X"E2",X"F0",X"F9",X"FF",X"CF",X"F2",X"E2",X"E2",X"42",X"02",X"02",X"C6",X"E6",
		X"E3",X"7F",X"3F",X"3E",X"00",X"00",X"00",X"01",X"E6",X"CE",X"8E",X"1E",X"7E",X"7E",X"FE",X"FE",
		X"00",X"07",X"06",X"05",X"05",X"04",X"07",X"05",X"00",X"F8",X"18",X"E8",X"E8",X"08",X"F8",X"68",
		X"05",X"05",X"04",X"07",X"05",X"05",X"05",X"06",X"68",X"68",X"08",X"F8",X"98",X"68",X"68",X"E8",
		X"00",X"1C",X"3C",X"7C",X"70",X"61",X"73",X"7F",X"00",X"3C",X"7E",X"FF",X"E7",X"C3",X"87",X"9F",
		X"3F",X"1E",X"00",X"3F",X"7F",X"7F",X"60",X"60",X"1E",X"1C",X"00",X"FF",X"FF",X"FF",X"C0",X"C0",
		X"07",X"06",X"05",X"05",X"06",X"07",X"07",X"07",X"F8",X"18",X"E8",X"E8",X"18",X"F8",X"E8",X"E8",
		X"04",X"07",X"06",X"05",X"05",X"06",X"07",X"00",X"08",X"F8",X"D8",X"E8",X"E8",X"18",X"F8",X"00",
		X"70",X"7F",X"3F",X"0F",X"00",X"1C",X"3C",X"7C",X"C0",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",
		X"70",X"60",X"60",X"70",X"7F",X"3F",X"1F",X"00",X"C3",X"C3",X"C3",X"07",X"FF",X"FE",X"FC",X"00",
		X"7F",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"00",X"00",X"00",X"01",X"00",X"00",X"02",X"04",X"02",X"02",X"02",X"82",X"42",X"42",X"22",X"22",
		X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"04",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"42",X"42",X"82",X"02",X"02",X"02",X"02",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"20",X"60",X"E0",X"E0",
		X"08",X"C8",X"28",X"F8",X"08",X"08",X"08",X"08",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",
		X"FF",X"FF",X"FF",X"0F",X"E3",X"F9",X"FC",X"FE",X"7F",X"3F",X"9F",X"CF",X"E7",X"F0",X"FF",X"7F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"C7",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"08",X"08",X"08",X"08",X"FB",X"0B",X"08",X"09",X"60",X"60",X"60",X"00",X"E0",X"E0",X"C0",X"80",
		X"03",X"03",X"00",X"03",X"03",X"00",X"00",X"00",X"E0",X"E0",X"00",X"E0",X"E0",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"01",X"01",X"02",X"00",X"F8",X"E1",X"DF",X"FD",X"FD",X"FE",X"FE",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"7E",X"3F",X"0F",X"03",X"01",X"00",X"00",
		X"FF",X"FF",X"EF",X"E1",X"B8",X"BE",X"4F",X"F2",X"C2",X"82",X"82",X"02",X"42",X"C2",X"82",X"82",
		X"EC",X"FC",X"F9",X"8E",X"C0",X"79",X"30",X"01",X"02",X"06",X"06",X"0E",X"0E",X"1E",X"3E",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"0F",X"0E",X"1E",X"1F",X"37",X"3E",X"3B",
		X"3B",X"1B",X"0B",X"0B",X"1B",X"0B",X"61",X"98",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"04",X"62",X"F2",X"BA",X"78",X"CC",X"A4",X"F2",X"7E",X"7E",X"7E",X"3E",X"3E",X"3E",X"3E",X"1E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"1F",X"10",X"1F",X"00",X"0E",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"1F",X"0E",X"00",X"1F",X"00",X"10",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"1E",X"1E",X"1E",X"0E",X"0E",X"1E",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1E",X"1E",X"1E",X"0E",X"1E",X"0E",X"0E",X"1E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"1F",X"01",X"1F",X"1F",X"00",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"12",X"1F",X"07",X"00",X"11",X"1F",X"0E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"1E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",
		X"62",X"40",X"45",X"62",X"40",X"45",X"66",X"49",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"87",
		X"60",X"40",X"41",X"6E",X"4C",X"40",X"41",X"63",X"BF",X"FF",X"87",X"EF",X"DF",X"87",X"FF",X"87",
		X"FF",X"FF",X"F6",X"E0",X"C0",X"C0",X"C0",X"C0",X"FE",X"0E",X"06",X"22",X"B2",X"92",X"92",X"02",
		X"C0",X"C0",X"F0",X"F0",X"F0",X"E0",X"E0",X"C0",X"46",X"4E",X"1E",X"4E",X"66",X"66",X"46",X"06",
		X"6A",X"40",X"40",X"40",X"41",X"60",X"41",X"60",X"FF",X"87",X"B7",X"86",X"FE",X"8E",X"AE",X"86",
		X"40",X"41",X"6E",X"4C",X"40",X"41",X"63",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"C0",X"C0",X"40",X"20",X"00",X"00",X"02",X"06",X"06",X"06",X"06",X"76",X"0E",X"06",X"62",
		X"14",X"84",X"C4",X"FC",X"FE",X"FF",X"FF",X"FF",X"12",X"92",X"F2",X"62",X"06",X"0E",X"FE",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"00",X"00",X"00",X"00",X"40",X"40",X"C0",X"C0",
		X"0F",X"00",X"03",X"07",X"0F",X"08",X"08",X"07",X"C0",X"00",X"C1",X"C1",X"C2",X"80",X"80",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"78",X"FE",X"8F",X"03",X"01",X"39",X"7C",X"7C",X"00",X"00",X"00",X"00",X"B0",X"B0",X"B0",X"B0",
		X"00",X"07",X"08",X"08",X"0F",X"0F",X"07",X"00",X"00",X"80",X"40",X"42",X"C1",X"C1",X"80",X"00",
		X"09",X"08",X"08",X"0F",X"0F",X"07",X"00",X"00",X"C0",X"40",X"40",X"C0",X"C0",X"80",X"00",X"00",
		X"5C",X"6C",X"39",X"01",X"03",X"8F",X"FE",X"78",X"B0",X"B0",X"B0",X"B0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"7B",X"FF",X"FF",X"EF",X"FF",X"FD",X"FF",X"FF",X"FF",X"F7",X"7F",X"FF",X"FE",
		X"FF",X"FB",X"FF",X"FD",X"DF",X"FF",X"7D",X"FF",X"FF",X"FB",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"FD",X"FF",X"FE",X"BD",X"FF",X"FF",X"DF",
		X"FF",X"FF",X"FD",X"DF",X"BA",X"8F",X"85",X"03",X"FF",X"FF",X"F7",X"FF",X"FC",X"FF",X"DF",X"FF",
		X"03",X"87",X"86",X"7F",X"FD",X"FB",X"EF",X"AF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"C0",X"C0",X"E0",X"E0",X"E0",X"F0",X"F0",X"0F",X"0F",X"07",X"07",X"03",X"03",X"01",X"01",
		X"F0",X"F8",X"F8",X"FC",X"FC",X"FF",X"FF",X"FF",X"01",X"01",X"83",X"C3",X"07",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"F1",X"E0",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",X"80",X"80",X"80",
		X"FC",X"E0",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",
		X"00",X"03",X"0F",X"1E",X"3C",X"38",X"71",X"62",X"00",X"C0",X"F0",X"78",X"3C",X"1C",X"8E",X"46",
		X"62",X"62",X"71",X"38",X"3C",X"1E",X"0F",X"03",X"46",X"46",X"8E",X"1C",X"3C",X"78",X"F0",X"C0",
		X"00",X"00",X"00",X"80",X"80",X"C0",X"E0",X"F8",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"07",
		X"7F",X"3F",X"3F",X"3F",X"1F",X"1F",X"1F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"03",X"03",X"01",X"00",X"02",X"01",X"6A",X"9C",X"AD",X"A5",X"91",X"CB",X"0A",X"0B",
		X"05",X"0C",X"0C",X"1E",X"1E",X"38",X"03",X"1D",X"40",X"82",X"C7",X"75",X"67",X"AD",X"1B",X"9F",
		X"00",X"00",X"03",X"07",X"07",X"0F",X"09",X"0D",X"7D",X"FC",X"E9",X"BF",X"4F",X"62",X"F7",X"A2",
		X"1A",X"1A",X"17",X"35",X"35",X"2F",X"3A",X"37",X"F5",X"2A",X"58",X"B0",X"21",X"93",X"67",X"A7",
		X"00",X"00",X"02",X"02",X"08",X"00",X"10",X"00",X"10",X"40",X"00",X"00",X"00",X"00",X"00",X"05",
		X"00",X"30",X"00",X"00",X"00",X"21",X"01",X"03",X"0D",X"1B",X"3B",X"3F",X"7F",X"5D",X"7F",X"77",
		X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"02",X"00",X"0F",X"1F",X"FF",X"F8",X"C0",X"02",X"17",
		X"04",X"04",X"00",X"00",X"08",X"01",X"03",X"03",X"1F",X"CF",X"6F",X"3F",X"3E",X"84",X"E0",X"F3",
		X"07",X"25",X"03",X"07",X"07",X"21",X"2B",X"08",X"7F",X"3F",X"7F",X"AD",X"BF",X"B5",X"5F",X"EF",
		X"15",X"14",X"06",X"0A",X"03",X"05",X"04",X"01",X"F7",X"E8",X"5F",X"1F",X"0B",X"83",X"C0",X"78",
		X"07",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"FF",X"FF",X"E7",X"81",X"01",X"04",X"07",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"7F",X"1F",X"1F",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FE",X"FE",X"FE",X"FC",X"FC",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"02",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"EE",X"3D",X"7B",X"3D",X"10",X"00",X"00",X"FF",X"FE",X"01",X"23",X"11",X"00",
		X"00",X"00",X"01",X"03",X"06",X"06",X"0C",X"0C",X"22",X"09",X"C4",X"E4",X"22",X"32",X"12",X"12");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
