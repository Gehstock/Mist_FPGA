library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity rom2t35 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of rom2t35 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"49",X"7F",X"49",X"49",X"00",X"36",X"00",X"00",X"24",X"1F",X"24",X"44",X"00",X"1F",X"00",X"00",
		X"41",X"7F",X"41",X"41",X"00",X"3E",X"00",X"00",X"41",X"3E",X"41",X"41",X"00",X"22",X"00",X"00",
		X"70",X"C3",X"FF",X"4A",X"FF",X"FF",X"01",X"FF",X"49",X"7F",X"49",X"49",X"00",X"41",X"00",X"00",
		X"08",X"7F",X"08",X"08",X"00",X"7F",X"00",X"00",X"41",X"3E",X"45",X"41",X"00",X"47",X"00",X"00",
		X"9C",X"CD",X"57",X"01",X"3D",X"84",X"67",X"3D",X"41",X"00",X"41",X"7F",X"00",X"00",X"00",X"00",
		X"01",X"7F",X"01",X"01",X"00",X"01",X"00",X"00",X"3D",X"3D",X"87",X"5F",X"C3",X"87",X"1D",X"FC",
		X"10",X"7F",X"04",X"08",X"00",X"7F",X"00",X"00",X"20",X"7F",X"20",X"18",X"00",X"7F",X"00",X"00",
		X"48",X"7F",X"48",X"48",X"00",X"30",X"00",X"00",X"41",X"3E",X"41",X"41",X"00",X"3E",X"00",X"00",
		X"48",X"7F",X"4A",X"4C",X"00",X"31",X"00",X"00",X"07",X"00",X"7E",X"1E",X"07",X"1E",X"00",X"00",
		X"40",X"40",X"40",X"7F",X"00",X"40",X"00",X"00",X"49",X"32",X"49",X"49",X"00",X"26",X"00",X"00",
		X"06",X"78",X"06",X"01",X"00",X"78",X"00",X"00",X"01",X"7E",X"01",X"01",X"00",X"7E",X"00",X"00",
		X"14",X"63",X"14",X"08",X"00",X"63",X"00",X"00",X"F1",X"CD",X"CD",X"09",X"09",X"CE",X"14",X"C9",
		X"45",X"43",X"51",X"49",X"00",X"61",X"00",X"00",X"10",X"60",X"10",X"0F",X"00",X"60",X"00",X"00",
		X"00",X"00",X"7F",X"21",X"00",X"01",X"00",X"00",X"3E",X"00",X"49",X"45",X"3E",X"51",X"00",X"00",
		X"42",X"00",X"49",X"41",X"66",X"59",X"00",X"00",X"23",X"00",X"49",X"45",X"31",X"49",X"00",X"00",
		X"72",X"00",X"51",X"51",X"4E",X"51",X"00",X"00",X"0C",X"00",X"24",X"14",X"04",X"7F",X"00",X"00",
		X"40",X"00",X"48",X"47",X"60",X"50",X"00",X"00",X"1E",X"00",X"49",X"29",X"46",X"49",X"00",X"00",
		X"31",X"00",X"49",X"49",X"3C",X"4A",X"00",X"00",X"36",X"00",X"49",X"49",X"36",X"49",X"00",X"00",
		X"5F",X"20",X"01",X"21",X"C3",X"3C",X"0B",X"D2",X"A1",X"21",X"C3",X"20",X"40",X"FE",X"AD",X"3A",
		X"7E",X"23",X"00",X"BB",X"00",X"00",X"E9",X"E1",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A9",X"21",X"C3",X"20",X"40",X"FE",X"00",X"00",X"A5",X"21",X"C3",X"20",X"40",X"FE",X"00",X"00",
		X"26",X"26",X"08",X"07",X"12",X"26",X"0E",X"02",X"12",X"26",X"0E",X"02",X"04",X"11",X"1B",X"26",
		X"26",X"04",X"26",X"1C",X"0B",X"0F",X"18",X"00",X"04",X"11",X"26",X"26",X"02",X"12",X"11",X"0E",
		X"1C",X"26",X"0F",X"26",X"00",X"0B",X"04",X"18",X"14",X"0F",X"07",X"12",X"26",X"1B",X"11",X"0E",
		X"02",X"0D",X"04",X"11",X"08",X"03",X"26",X"13",X"12",X"11",X"01",X"26",X"13",X"14",X"0E",X"13",
		X"0B",X"0F",X"18",X"00",X"11",X"04",X"1C",X"26",X"0B",X"0F",X"18",X"00",X"11",X"04",X"1B",X"26",
		X"0A",X"00",X"26",X"E5",X"6F",X"00",X"29",X"29",X"0F",X"26",X"08",X"0E",X"13",X"0D",X"11",X"12",
		X"1A",X"C5",X"13",X"77",X"20",X"01",X"09",X"00",X"19",X"29",X"E1",X"EB",X"08",X"06",X"04",X"D3",
		X"23",X"56",X"23",X"7E",X"6F",X"66",X"CD",X"7A",X"05",X"C1",X"B8",X"C2",X"C9",X"0B",X"23",X"5E",
		X"E6",X"0F",X"CD",X"0F",X"0B",X"E6",X"E6",X"F1",X"0B",X"D3",X"D5",X"7B",X"0F",X"F5",X"0F",X"0F",
		X"3C",X"C3",X"AF",X"09",X"81",X"7D",X"6F",X"27",X"CD",X"0F",X"0B",X"E6",X"C9",X"D1",X"1A",X"C6",
		X"11",X"0E",X"04",X"13",X"26",X"17",X"76",X"F3",X"88",X"7C",X"C3",X"27",X"41",X"1B",X"15",X"26",
		X"30",X"17",X"70",X"11",X"CD",X"0B",X"0A",X"B0",X"3F",X"FE",X"F8",X"C2",X"0E",X"17",X"21",X"04",
		X"01",X"06",X"05",X"FB",X"1A",X"C2",X"CD",X"08",X"0F",X"0E",X"15",X"21",X"C3",X"2A",X"09",X"0D",
		X"20",X"AD",X"0E",X"6F",X"CD",X"01",X"0B",X"EB",X"0A",X"28",X"18",X"C2",X"26",X"08",X"3A",X"00",
		X"20",X"AD",X"99",X"FE",X"53",X"D2",X"CD",X"08",X"32",X"7D",X"20",X"AD",X"26",X"CD",X"3A",X"0B",
		X"0B",X"74",X"13",X"21",X"CD",X"28",X"09",X"F1",X"0A",X"28",X"53",X"CA",X"0E",X"08",X"11",X"15",
		X"62",X"DA",X"DB",X"08",X"E6",X"03",X"C2",X"02",X"18",X"C3",X"3A",X"08",X"20",X"AD",X"02",X"FE",
		X"3E",X"09",X"C3",X"01",X"08",X"7B",X"16",X"CD",X"08",X"6E",X"03",X"DB",X"04",X"E6",X"08",X"CA",
		X"3E",X"20",X"32",X"02",X"20",X"F1",X"16",X"CD",X"DB",X"09",X"E6",X"02",X"3C",X"03",X"E1",X"32",
		X"32",X"3C",X"20",X"E0",X"C6",X"CD",X"00",X"03",X"CD",X"09",X"0B",X"26",X"02",X"DB",X"03",X"E6",
		X"08",X"0E",X"17",X"21",X"11",X"2F",X"0B",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7D",X"E5",X"DD",X"C6",X"24",X"6F",X"B8",X"7E",X"F1",X"CD",X"C3",X"09",X"08",X"BC",X"44",X"4D",
		X"FE",X"81",X"C9",X"81",X"AF",X"CD",X"21",X"03",X"7E",X"23",X"C3",X"B9",X"04",X"B2",X"E6",X"F3",
		X"08",X"06",X"21",X"EF",X"23",X"80",X"08",X"06",X"23",X"00",X"08",X"06",X"21",X"EF",X"23",X"40",
		X"DF",X"09",X"C2",X"05",X"08",X"D9",X"F6",X"21",X"21",X"EF",X"23",X"C0",X"08",X"06",X"06",X"EF",
		X"EF",X"22",X"CD",X"97",X"1C",X"00",X"9F",X"31",X"06",X"22",X"EF",X"05",X"08",X"06",X"ED",X"21",
		X"B4",X"7D",X"B2",X"B3",X"C2",X"A7",X"01",X"5C",X"2A",X"20",X"20",X"A5",X"2A",X"EB",X"20",X"A9",
		X"04",X"D3",X"37",X"C3",X"11",X"08",X"09",X"2D",X"4E",X"21",X"22",X"00",X"20",X"9F",X"C9",X"FB",
		X"3D",X"20",X"E6",X"47",X"FE",X"0F",X"C2",X"0F",X"F1",X"CD",X"C3",X"09",X"08",X"18",X"AD",X"3A",
		X"32",X"78",X"20",X"AD",X"1B",X"C9",X"0F",X"26",X"09",X"28",X"E6",X"78",X"F6",X"F0",X"47",X"09",
		X"13",X"13",X"0D",X"0E",X"CD",X"00",X"0B",X"A7",X"00",X"0B",X"04",X"18",X"26",X"11",X"14",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CD",X"C9",X"4A",X"C4",X"00",X"00",
		X"DF",X"00",X"21",X"DF",X"28",X"10",X"F7",X"CD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"D2",X"CD",X"DF",X"0B",X"10",X"21",X"0E",X"35",X"DF",X"0C",X"10",X"21",X"1E",X"33",X"00",X"20",
		X"28",X"0C",X"F5",X"CD",X"DF",X"10",X"0C",X"21",X"11",X"07",X"0B",X"A0",X"BB",X"CD",X"21",X"09",
		X"00",X"00",X"0C",X"21",X"0E",X"35",X"11",X"07",X"1E",X"33",X"00",X"50",X"D2",X"CD",X"DF",X"0B",
		X"F5",X"CD",X"DF",X"07",X"08",X"21",X"11",X"31",X"0B",X"A0",X"BB",X"CD",X"21",X"09",X"28",X"08",
		X"08",X"21",X"0E",X"35",X"11",X"07",X"0B",X"A0",X"C1",X"00",X"CE",X"CD",X"DF",X"0B",X"00",X"00",
		X"FF",X"FF",X"1A",X"FF",X"00",X"D5",X"A7",X"CD",X"BB",X"CD",X"CD",X"09",X"40",X"4C",X"FF",X"C9",
		X"09",X"BB",X"CD",X"C9",X"1C",X"F3",X"1C",X"0E",X"00",X"0B",X"DF",X"D1",X"00",X"13",X"C2",X"0D",
		X"CD",X"09",X"0B",X"40",X"20",X"CD",X"CD",X"0B",X"1E",X"21",X"11",X"24",X"0B",X"50",X"F1",X"CD",
		X"0B",X"89",X"F1",X"CD",X"C3",X"09",X"0D",X"DB",X"0B",X"48",X"07",X"0E",X"01",X"21",X"11",X"35",
		X"00",X"D1",X"0D",X"13",X"F1",X"C2",X"C9",X"09",X"1A",X"C9",X"00",X"D5",X"A7",X"CD",X"00",X"0B",
		X"0C",X"E2",X"0D",X"10",X"0D",X"25",X"0D",X"3A",X"0C",X"8E",X"0C",X"A3",X"0C",X"B8",X"0C",X"CD",
		X"FF",X"7F",X"80",X"00",X"E3",X"7F",X"80",X"FF",X"00",X"00",X"3E",X"3E",X"00",X"FF",X"3E",X"00",
		X"80",X"C1",X"01",X"01",X"C0",X"FF",X"80",X"20",X"E3",X"C0",X"00",X"C1",X"FF",X"01",X"C0",X"C0",
		X"00",X"02",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"FF",X"02",X"00",X"20",X"00",X"00",
		X"00",X"FF",X"38",X"00",X"FF",X"7C",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"01",X"C6",X"01",X"00",X"00",X"FF",X"EE",X"7C",X"00",X"FF",X"EE",X"00",X"FF",X"C6",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"01",X"00",X"FF",X"00",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"FF",X"F8",X"00",X"FF",X"F8",X"00",X"00",X"FF",X"FF",X"00",X"00",X"F8",X"FC",X"00",X"01",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"20",X"F8",X"00",X"FF",X"20",X"00",X"FF",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"00",X"FF",X"FC",X"00",X"07",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"FF",X"F0",X"00",X"01",X"40",X"FF",X"00",X"FF",X"01",X"00",X"00",X"F0",X"F0",X"01",X"01",
		X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"40",X"40",X"00",X"FF",X"40",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0C",X"86",X"10",X"21",X"C3",X"2E",X"0F",X"F5",X"FF",X"FF",X"FF",X"FF",X"A6",X"11",X"CD",X"10",
		X"0C",X"3A",X"0C",X"4F",X"0C",X"64",X"0C",X"79",X"06",X"EB",X"0C",X"10",X"0C",X"25",X"07",X"E0",
		X"DC",X"00",X"0F",X"F4",X"FF",X"0F",X"00",X"00",X"00",X"00",X"EC",X"EC",X"0F",X"0F",X"00",X"FF",
		X"12",X"F2",X"FF",X"03",X"00",X"00",X"E3",X"E0",X"FA",X"38",X"07",X"17",X"00",X"FF",X"F0",X"00",
		X"FF",X"00",X"00",X"00",X"07",X"00",X"00",X"38",X"01",X"31",X"00",X"FF",X"00",X"00",X"3E",X"1F",
		X"00",X"FF",X"EE",X"00",X"06",X"FA",X"FF",X"07",X"FF",X"FF",X"00",X"00",X"F6",X"F6",X"05",X"05",
		X"78",X"00",X"09",X"F9",X"FF",X"01",X"80",X"00",X"00",X"00",X"FD",X"9C",X"03",X"0B",X"00",X"FF",
		X"1F",X"0F",X"FF",X"00",X"80",X"00",X"03",X"00",X"F1",X"F0",X"00",X"18",X"00",X"FF",X"00",X"80",
		X"02",X"02",X"00",X"FF",X"37",X"00",X"03",X"3D",X"00",X"1C",X"FF",X"FF",X"00",X"00",X"1B",X"1B",
		X"00",X"FF",X"BC",X"80",X"04",X"FC",X"FF",X"00",X"FF",X"03",X"80",X"00",X"FE",X"CE",X"01",X"05",
		X"80",X"C0",X"0F",X"07",X"FF",X"00",X"C0",X"00",X"C0",X"00",X"78",X"78",X"00",X"0C",X"00",X"FF",
		X"05",X"0D",X"01",X"01",X"80",X"FF",X"9B",X"80",X"01",X"00",X"00",X"0E",X"FF",X"FF",X"80",X"80",
		X"00",X"02",X"00",X"FF",X"5E",X"40",X"02",X"7E",X"01",X"86",X"FF",X"01",X"40",X"00",X"CF",X"E7",
		X"00",X"FF",X"C0",X"E0",X"07",X"03",X"FF",X"00",X"FF",X"00",X"60",X"00",X"3C",X"3C",X"00",X"06",
		X"80",X"80",X"3F",X"2F",X"80",X"FF",X"3F",X"80",X"E0",X"00",X"00",X"00",X"00",X"07",X"FF",X"FF",
		X"0D",X"00",X"FF",X"07",X"00",X"00",X"02",X"07",X"FF",X"0D",X"80",X"80",X"0F",X"0F",X"80",X"FF",
		X"86",X"CD",X"C9",X"0C",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"11",X"FF",X"11",X"10",
		X"07",X"20",X"07",X"30",X"07",X"40",X"07",X"50",X"1E",X"7A",X"1E",X"8A",X"1E",X"9A",X"07",X"10",
		X"FF",X"09",X"00",X"00",X"10",X"02",X"00",X"FF",X"80",X"80",X"4E",X"5C",X"00",X"FF",X"24",X"00",
		X"FF",X"27",X"00",X"40",X"24",X"02",X"00",X"FF",X"0C",X"00",X"FF",X"0C",X"40",X"FF",X"1E",X"80",
		X"FF",X"FF",X"80",X"C0",X"03",X"01",X"20",X"FF",X"02",X"00",X"FF",X"04",X"00",X"00",X"03",X"0C",
		X"40",X"FF",X"00",X"00",X"FF",X"02",X"C8",X"FF",X"09",X"90",X"FF",X"04",X"60",X"20",X"04",X"06",
		X"20",X"FF",X"00",X"00",X"FF",X"01",X"C0",X"C0",X"05",X"E8",X"FF",X"04",X"90",X"40",X"00",X"02",
		X"12",X"FF",X"00",X"20",X"FF",X"01",X"20",X"10",X"FF",X"FF",X"FF",X"FF",X"3C",X"F2",X"01",X"00",
		X"3A",X"FF",X"FF",X"5C",X"90",X"09",X"91",X"FF",X"60",X"FF",X"FF",X"18",X"FF",X"FF",X"FF",X"FF",
		X"DF",X"1D",X"C9",X"DF",X"FF",X"FF",X"30",X"30",X"FF",X"89",X"46",X"62",X"FF",X"FF",X"AA",X"CD",
		X"C3",X"F1",X"00",X"08",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3E",X"F5",X"32",X"AA",X"22",X"48",
		X"FF",X"FF",X"EB",X"CD",X"84",X"19",X"C3",X"67",X"FF",X"FF",X"F0",X"FF",X"FF",X"F0",X"60",X"60",
		X"F0",X"F0",X"03",X"03",X"E0",X"FF",X"01",X"E0",X"0A",X"48",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"F0",X"FF",X"0F",X"F0",X"FF",X"01",X"C0",X"C0",X"FF",X"FF",X"FF",X"FF",
		X"07",X"E0",X"FF",X"07",X"C0",X"C0",X"03",X"03",X"FF",X"0F",X"F0",X"F0",X"0F",X"0F",X"E0",X"FF",
		X"1F",X"E0",X"FF",X"1F",X"C0",X"C0",X"0F",X"0F",X"FF",X"FF",X"E0",X"E0",X"1F",X"1F",X"E0",X"FF",
		X"1E",X"41",X"86",X"CD",X"C3",X"0C",X"0D",X"FA",X"80",X"FF",X"07",X"80",X"FF",X"07",X"11",X"FF",
		X"1D",X"21",X"1D",X"31",X"1D",X"41",X"1E",X"31",X"1C",X"B9",X"1C",X"C9",X"1C",X"D9",X"1D",X"11",
		X"FF",X"0F",X"00",X"00",X"06",X"06",X"FF",X"FF",X"80",X"80",X"1F",X"1F",X"00",X"FF",X"0F",X"00",
		X"FF",X"1E",X"00",X"00",X"0C",X"0C",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"1E",X"00",
		X"FF",X"FF",X"00",X"00",X"18",X"18",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"FF",X"07",X"00",X"00",X"01",X"FF",X"00",X"1F",X"C0",X"FF",X"07",X"C0",X"C0",X"07",X"07",
		X"FF",X"00",X"D2",X"FF",X"08",X"53",X"C5",X"F5",X"00",X"00",X"01",X"01",X"00",X"FF",X"01",X"00",
		X"86",X"41",X"47",X"23",X"A7",X"7D",X"9D",X"CA",X"26",X"E5",X"2E",X"0B",X"6E",X"DE",X"F3",X"3A",
		X"80",X"C0",X"0F",X"1F",X"80",X"FF",X"0F",X"80",X"78",X"0D",X"79",X"C3",X"FF",X"0D",X"FF",X"FF",
		X"02",X"00",X"FF",X"00",X"78",X"FF",X"C0",X"A7",X"FF",X"0F",X"00",X"80",X"02",X"0F",X"00",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C1",X"E1",X"C3",X"F1",X"08",X"3F",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3B",X"1F",X"80",X"FF",X"3B",X"80",X"FF",X"31",X"00",X"FF",X"0E",X"00",X"FF",X"1F",X"80",X"00",
		X"FF",X"00",X"CD",X"FF",X"0B",X"26",X"03",X"0E",X"40",X"80",X"40",X"31",X"40",X"FF",X"40",X"00",
		X"C9",X"48",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"9C",X"21",X"11",X"30",X"22",X"51",X"2C",X"CD",
		X"FF",X"FF",X"10",X"21",X"C3",X"2B",X"0E",X"F4",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
