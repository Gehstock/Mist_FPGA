library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity tropical_spr_bit5 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of tropical_spr_bit5 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"07",X"0F",X"0F",X"0F",X"07",X"07",X"07",X"07",X"03",X"01",X"01",X"0F",X"3F",X"7F",X"7F",
		X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"C0",X"C0",X"C0",X"F0",X"FC",X"FE",X"FE",
		X"7F",X"3F",X"0F",X"17",X"16",X"37",X"63",X"01",X"00",X"00",X"08",X"1E",X"0F",X"0F",X"07",X"00",
		X"7E",X"7F",X"7D",X"78",X"78",X"FC",X"FE",X"30",X"B8",X"98",X"18",X"3C",X"3C",X"3C",X"BC",X"BC",
		X"0E",X"06",X"06",X"06",X"03",X"03",X"01",X"01",X"03",X"07",X"01",X"03",X"03",X"03",X"01",X"01",
		X"20",X"20",X"E0",X"60",X"60",X"60",X"60",X"60",X"20",X"20",X"30",X"30",X"30",X"30",X"F0",X"F0",
		X"00",X"00",X"00",X"03",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"03",X"00",X"01",X"07",
		X"00",X"00",X"00",X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"E0",X"C0",X"C0",X"FC",X"FE",
		X"FF",X"FF",X"FF",X"EF",X"EF",X"EF",X"E7",X"F7",X"81",X"B7",X"3F",X"1F",X"0F",X"01",X"00",X"00",
		X"F0",X"F8",X"F8",X"DC",X"8C",X"AE",X"E6",X"F0",X"C0",X"C0",X"C0",X"C0",X"E0",X"E0",X"70",X"F0",
		X"01",X"C3",X"21",X"31",X"78",X"7D",X"7F",X"3C",X"0C",X"0E",X"1A",X"03",X"07",X"07",X"0B",X"0B",
		X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"40",X"40",X"C0",X"40",
		X"0F",X"1F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"1F",X"0F",X"03",X"07",X"0F",X"1F",X"3F",X"3B",
		X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"00",X"00",X"E0",X"F8",X"FC",X"FE",X"FE",
		X"7F",X"7E",X"3C",X"BC",X"BC",X"BC",X"FC",X"BF",X"BF",X"BF",X"7F",X"27",X"07",X"27",X"27",X"33",
		X"60",X"36",X"34",X"18",X"18",X"00",X"00",X"00",X"C0",X"E0",X"F0",X"F8",X"FC",X"FC",X"FE",X"FE",
		X"E0",X"F0",X"F8",X"FC",X"7C",X"3C",X"0E",X"2E",X"6A",X"CB",X"CD",X"E5",X"73",X"79",X"D8",X"18",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"C0",
		X"00",X"01",X"03",X"03",X"03",X"03",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"F8",X"FC",X"FC",X"FC",X"FC",X"FC",X"F8",X"F8",X"F0",X"10",X"7F",X"7F",X"7F",X"FF",X"DF",
		X"80",X"C0",X"E0",X"F0",X"F0",X"B9",X"1F",X"0F",X"87",X"82",X"FE",X"FF",X"FF",X"5F",X"07",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"C0",X"40",X"00",X"00",X"00",X"80",X"C0",X"F0",X"F8",X"FC",
		X"60",X"F8",X"FC",X"FC",X"FE",X"3E",X"7F",X"D9",X"0D",X"06",X"83",X"D0",X"EC",X"BF",X"BE",X"1E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"60",X"20",X"30",X"10",
		X"00",X"00",X"00",X"07",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"07",X"03",X"00",X"38",X"7F",
		X"00",X"00",X"00",X"C0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"C0",X"40",X"C0",X"F0",
		X"0F",X"1F",X"1F",X"3F",X"31",X"05",X"07",X"0F",X"19",X"01",X"09",X"0B",X"1F",X"1F",X"3F",X"3F",
		X"FF",X"FF",X"FF",X"F7",X"F6",X"F7",X"E7",X"EF",X"83",X"ED",X"E8",X"F0",X"A0",X"00",X"80",X"98",
		X"03",X"03",X"03",X"03",X"02",X"02",X"02",X"02",X"01",X"01",X"01",X"01",X"02",X"02",X"02",X"02",
		X"84",X"08",X"08",X"10",X"1C",X"14",X"34",X"2C",X"28",X"E8",X"38",X"38",X"30",X"30",X"70",X"70",
		X"01",X"01",X"03",X"03",X"03",X"03",X"03",X"01",X"01",X"00",X"00",X"06",X"1F",X"3F",X"7F",X"7F",
		X"F0",X"F8",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"F8",X"F0",X"00",X"10",X"F8",X"FC",X"FC",X"FC",
		X"03",X"37",X"16",X"0C",X"0C",X"00",X"01",X"03",X"0F",X"1F",X"3F",X"7F",X"7F",X"FF",X"FF",X"FF",
		X"7E",X"3E",X"1E",X"1C",X"7D",X"7F",X"FE",X"FE",X"3E",X"12",X"00",X"00",X"80",X"80",X"8C",X"98",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"03",
		X"0F",X"1E",X"1E",X"3C",X"3C",X"38",X"78",X"71",X"72",X"F6",X"FC",X"C4",X"CC",X"C8",X"88",X"98",
		X"1F",X"1F",X"3F",X"3F",X"3F",X"3F",X"3F",X"1F",X"1F",X"0F",X"C8",X"FE",X"FE",X"FE",X"FF",X"FB",
		X"00",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"07",X"03",X"02",X"00",X"00",X"00",X"01",X"03",X"07",X"0F",X"1F",
		X"01",X"03",X"07",X"0F",X"0F",X"9D",X"F8",X"F0",X"E1",X"43",X"1F",X"FF",X"FB",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"03",X"07",X"04",X"0D",X"09",
		X"06",X"1F",X"3F",X"3F",X"7F",X"7F",X"FB",X"97",X"8E",X"0C",X"D4",X"B6",X"60",X"E0",X"C0",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"38",X"7A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"3C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"1E",X"1C",X"39",X"3C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"E8",X"EC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"E0",X"E8",X"EC",X"EE",X"E8",X"E0",X"80",X"80",
		X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"00",X"01",X"01",X"01",X"01",X"01",X"01",
		X"00",X"00",X"00",X"00",X"C0",X"D0",X"D8",X"DC",X"D8",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E6",X"E7",X"E7",X"E6",X"E0",X"40",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
		X"E4",X"E0",X"40",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",
		X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"12",X"01",X"0C",X"17",X"45",X"03",X"07",X"0B",X"00",X"41",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"40",X"C0",X"40",X"80",X"C0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"04",X"23",X"05",X"0F",X"13",X"44",X"01",X"03",X"05",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"80",X"C0",X"80",X"C0",X"E0",X"80",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"09",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"04",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"3F",X"0F",X"17",X"16",X"37",X"63",X"01",X"00",X"00",X"08",X"1E",X"0F",X"0F",X"07",X"00",
		X"7E",X"7F",X"7D",X"78",X"78",X"FC",X"FE",X"30",X"B8",X"98",X"18",X"3C",X"3C",X"3C",X"BC",X"BC",
		X"00",X"00",X"00",X"11",X"0F",X"07",X"0F",X"0F",X"0E",X"06",X"06",X"06",X"03",X"03",X"01",X"01",
		X"38",X"98",X"88",X"18",X"10",X"30",X"30",X"20",X"20",X"20",X"E0",X"60",X"60",X"60",X"60",X"60",
		X"01",X"01",X"00",X"02",X"02",X"02",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"B0",X"90",X"90",X"90",X"D0",X"F0",X"70",X"70",X"70",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"0F",X"0F",X"0F",X"0E",X"0E",X"0E",X"0E",X"0F",X"08",X"0B",X"13",X"01",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FD",X"F8",X"FA",X"7E",X"7F",X"1C",X"7C",X"FC",X"FC",X"FE",X"1E",X"07",X"0F",
		X"31",X"39",X"19",X"1D",X"04",X"01",X"00",X"00",X"04",X"07",X"00",X"00",X"01",X"01",X"01",X"00",
		X"F8",X"F8",X"F8",X"FC",X"FC",X"FC",X"FC",X"FC",X"04",X"0C",X"86",X"C6",X"E2",X"F6",X"FE",X"F2",
		X"01",X"05",X"05",X"04",X"02",X"03",X"03",X"03",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",
		X"A0",X"A0",X"80",X"C0",X"70",X"70",X"70",X"70",X"F8",X"F8",X"F8",X"F8",X"FC",X"FC",X"FC",X"FC",
		X"3B",X"5B",X"59",X"5D",X"4D",X"2D",X"2F",X"25",X"15",X"05",X"03",X"01",X"00",X"01",X"01",X"01",
		X"FB",X"F1",X"E1",X"E0",X"E0",X"E0",X"E0",X"F8",X"FE",X"FF",X"FF",X"3F",X"3F",X"3F",X"3F",X"9F",
		X"19",X"09",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"CF",X"37",X"81",X"C0",X"60",X"F0",X"FD",X"FF",X"3F",X"0F",X"01",X"01",X"03",X"00",
		X"1C",X"0E",X"07",X"01",X"04",X"06",X"03",X"03",X"03",X"01",X"01",X"01",X"00",X"00",X"00",X"00",
		X"40",X"40",X"60",X"E0",X"E0",X"F0",X"30",X"F0",X"F8",X"F8",X"F8",X"FC",X"FC",X"FC",X"FE",X"7E",
		X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DF",X"DF",X"5F",X"4F",X"6F",X"A3",X"59",X"3C",X"1E",X"39",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"0F",X"07",X"37",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FF",X"FF",X"BF",X"1F",X"03",X"00",X"F0",X"3C",X"3E",X"7F",X"7F",X"1F",X"0F",X"00",X"01",
		X"0F",X"07",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"18",X"B8",X"FC",X"7C",X"96",X"E6",X"7F",X"7F",X"3F",X"3F",X"1F",X"1F",X"0F",X"0F",X"07",X"07",
		X"FF",X"FF",X"FF",X"FF",X"1F",X"5F",X"7E",X"FE",X"98",X"1E",X"9E",X"BF",X"FA",X"F0",X"F8",X"F9",
		X"F8",X"FC",X"FC",X"7E",X"66",X"76",X"76",X"F2",X"30",X"D8",X"8C",X"00",X"00",X"00",X"00",X"80",
		X"3F",X"3F",X"7F",X"7E",X"78",X"70",X"70",X"E1",X"E1",X"C2",X"C2",X"C4",X"87",X"85",X"8D",X"8B",
		X"98",X"38",X"70",X"40",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"04",X"04",X"04",X"0C",X"0C",X"0C",X"0C",X"1F",X"1F",X"1F",X"1F",X"3F",X"3F",X"3F",X"3F",
		X"20",X"20",X"60",X"60",X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",
		X"DF",X"CF",X"87",X"07",X"1F",X"1F",X"7F",X"FF",X"CF",X"C4",X"C0",X"C0",X"E0",X"E0",X"E3",X"E6",
		X"B8",X"B8",X"B4",X"34",X"68",X"E8",X"90",X"90",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"DC",X"C0",X"80",X"87",X"0C",X"10",X"30",X"40",X"C0",X"80",X"80",X"80",X"00",X"00",X"00",
		X"38",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"03",X"07",X"04",X"04",X"0C",X"0C",X"0F",X"1F",X"1F",X"1F",X"3F",X"3F",X"3F",X"7F",X"7E",
		X"10",X"10",X"30",X"60",X"E0",X"E0",X"C0",X"C0",X"C0",X"80",X"80",X"80",X"00",X"00",X"00",X"00",
		X"FB",X"FB",X"F2",X"E6",X"ED",X"A2",X"32",X"60",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"7F",X"7B",X"FB",X"F0",X"F0",X"C0",X"83",X"04",X"18",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"E0",X"C0",X"80",X"08",X"0C",X"04",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1B",X"1E",X"3C",X"39",X"63",X"67",X"FE",X"FE",X"FC",X"FC",X"F8",X"F8",X"F0",X"F0",X"E0",X"E0",
		X"00",X"40",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"80",X"00",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"02",X"14",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"40",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"0B",X"03",X"16",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"D0",X"90",X"00",X"B0",X"70",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"01",X"0B",X"0D",X"2F",X"3C",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"D0",X"50",X"00",X"80",X"30",X"38",X"78",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"09",X"0B",X"25",X"3F",X"1C",X"07",
		X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"A8",X"88",X"00",X"E8",X"98",X"1C",X"3C",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"19",X"1B",X"15",X"45",X"7F",X"1C",X"03",
		X"00",X"00",X"00",X"00",X"40",X"E0",X"E0",X"A4",X"8C",X"00",X"E0",X"D4",X"8E",X"3E",X"3C",X"F8",
		X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"10",X"3B",X"37",X"2B",X"89",X"FB",X"7F",X"08",X"07",
		X"00",X"40",X"E0",X"E0",X"F0",X"D2",X"D6",X"82",X"00",X"E0",X"93",X"17",X"BF",X"3E",X"7C",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"01",X"04",X"04",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"40",X"30",X"50",X"40",X"50",X"D8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"01",X"04",X"06",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"60",X"40",X"28",X"60",X"68",X"DC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"01",X"05",X"04",X"06",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"60",X"60",X"28",X"28",X"64",X"64",X"44",X"CE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"02",X"0A",X"18",X"18",X"1C",X"3C",X"1F",
		X"00",X"00",X"00",X"00",X"30",X"70",X"60",X"C0",X"E8",X"68",X"44",X"C4",X"C4",X"E4",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0E",X"06",X"16",X"12",X"30",X"31",X"39",X"79",X"3F",
		X"00",X"00",X"00",X"30",X"70",X"60",X"E0",X"E4",X"62",X"62",X"E2",X"E2",X"E2",X"F6",X"F7",X"00",
		X"00",X"00",X"00",X"00",X"04",X"0C",X"1E",X"0A",X"2E",X"24",X"20",X"60",X"71",X"71",X"F1",X"3F",
		X"00",X"00",X"30",X"70",X"60",X"F0",X"B4",X"64",X"62",X"E2",X"E2",X"E2",X"C6",X"CE",X"EF",X"FC",
		X"00",X"00",X"08",X"1C",X"3E",X"1A",X"4E",X"44",X"44",X"40",X"70",X"F1",X"F1",X"F1",X"F3",X"1F",
		X"30",X"70",X"60",X"F0",X"B0",X"34",X"74",X"62",X"62",X"E6",X"E6",X"C6",X"C6",X"8F",X"DE",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"03",X"01",X"00",X"00",
		X"38",X"38",X"7C",X"14",X"5C",X"CC",X"84",X"84",X"80",X"E0",X"E1",X"F1",X"E1",X"E1",X"E3",X"3F",
		X"72",X"F8",X"98",X"B9",X"3D",X"79",X"71",X"72",X"70",X"F0",X"F1",X"E1",X"C3",X"C7",X"EF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"C0",X"C0",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"03",X"03",X"03",X"03",X"07",X"03",X"00",
		X"3C",X"7E",X"3A",X"9E",X"8E",X"8C",X"04",X"00",X"C0",X"E0",X"F0",X"F0",X"E0",X"E1",X"E3",X"3F",
		X"6C",X"5C",X"5C",X"1E",X"3C",X"38",X"7C",X"7C",X"7C",X"78",X"F8",X"F0",X"E1",X"E7",X"F7",X"FF",
		X"00",X"40",X"40",X"40",X"C0",X"A0",X"20",X"20",X"60",X"60",X"60",X"F0",X"F0",X"E0",X"C0",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"80",X"80",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",X"80",X"80",X"80",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"05",
		X"00",X"00",X"00",X"00",X"C0",X"E0",X"E0",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"0D",X"03",
		X"00",X"C0",X"C0",X"D0",X"C0",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"10",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"0D",X"07",
		X"E8",X"E0",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"0C",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"13",X"3A",X"0F",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"04",X"0C",X"FE",
		X"01",X"01",X"01",X"03",X"03",X"03",X"03",X"03",X"03",X"07",X"46",X"E6",X"3C",X"7F",X"1C",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0E",X"3C",X"F6",X"FC",X"2A",
		X"01",X"01",X"01",X"01",X"01",X"01",X"03",X"23",X"43",X"C7",X"66",X"3C",X"1F",X"37",X"C2",X"02",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"82",X"01",X"01",X"02",X"1F",X"FF",X"DE",X"0A",X"05",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"E8",X"EC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"01",X"01",X"01",X"01",X"23",X"43",X"C3",X"83",X"87",X"C7",X"7E",X"3C",X"7F",X"DF",X"0E",X"35",
		X"80",X"80",X"80",X"80",X"80",X"81",X"81",X"80",X"00",X"01",X"03",X"1F",X"FF",X"8B",X"05",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",X"C0",X"80",X"00",X"80",X"C0",X"80",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"E0",X"E4",X"E7",X"E7",X"E7",X"E7",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"01",X"07",X"01",X"03",X"01",X"00",X"02",X"00",X"01",X"06",X"00",X"01",
		X"01",X"01",X"03",X"83",X"83",X"03",X"07",X"07",X"87",X"C7",X"7E",X"DC",X"0E",X"07",X"3F",X"C6",
		X"C0",X"C0",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"07",X"0F",X"1E",X"F1",X"02",X"80",
		X"00",X"00",X"00",X"00",X"60",X"30",X"28",X"30",X"60",X"C0",X"E0",X"F8",X"D0",X"40",X"20",X"00",
		X"00",X"00",X"C0",X"E0",X"30",X"F2",X"F3",X"F3",X"F3",X"F3",X"F3",X"F3",X"F0",X"30",X"C0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"F0",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"00",X"00",X"01",X"00",X"20",X"04",X"00",X"00",X"00",X"00",X"09",X"23",X"01",X"01",X"00",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"30",X"68",X"B0",X"08",X"C4",X"C4",X"E0",
		X"00",X"00",X"04",X"10",X"00",X"00",X"00",X"00",X"09",X"20",X"01",X"00",X"02",X"00",X"11",X"03",
		X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"F0",X"3A",X"54",X"18",X"B0",X"C8",X"A2",
		X"00",X"03",X"05",X"20",X"00",X"00",X"09",X"00",X"00",X"40",X"00",X"00",X"08",X"00",X"44",X"03",
		X"F0",X"A0",X"40",X"F0",X"28",X"F0",X"7C",X"18",X"28",X"74",X"9A",X"30",X"74",X"38",X"D0",X"8C",
		X"01",X"12",X"00",X"09",X"02",X"00",X"20",X"00",X"00",X"08",X"00",X"42",X"00",X"00",X"00",X"00",
		X"F0",X"78",X"E8",X"D8",X"A0",X"68",X"10",X"7C",X"B8",X"0D",X"18",X"68",X"A4",X"6C",X"D2",X"B1",
		X"00",X"01",X"00",X"00",X"09",X"00",X"00",X"01",X"08",X"41",X"02",X"0B",X"07",X"03",X"01",X"42",
		X"48",X"38",X"78",X"E8",X"78",X"20",X"F4",X"78",X"D4",X"60",X"7A",X"AC",X"09",X"A3",X"05",X"4D",
		X"00",X"00",X"04",X"00",X"00",X"04",X"20",X"02",X"01",X"00",X"00",X"00",X"45",X"02",X"13",X"07",
		X"20",X"90",X"78",X"38",X"F0",X"58",X"38",X"50",X"F8",X"E8",X"54",X"C6",X"52",X"09",X"2C",X"9A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"03",X"07",X"07",
		X"00",X"00",X"03",X"1F",X"20",X"00",X"00",X"00",X"00",X"80",X"83",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"C0",X"F8",X"04",X"00",X"00",X"00",X"00",X"01",X"C1",X"FF",X"FF",X"FF",X"FF",X"DF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"C0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",
		X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"10",X"70",X"71",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"7C",X"FF",X"00",X"00",X"00",X"00",X"40",X"40",X"E0",X"FF",X"FF",X"FF",X"FF",X"DF",
		X"00",X"00",X"00",X"00",X"80",X"40",X"20",X"20",X"20",X"20",X"20",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"38",X"79",X"7F",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"1F",X"FF",X"00",X"00",X"00",X"00",X"40",X"40",X"E0",X"FF",X"FF",X"FF",X"FF",X"BF",
		X"00",X"00",X"80",X"C0",X"C0",X"60",X"20",X"20",X"20",X"20",X"20",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"06",X"1E",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"07",X"3F",X"00",X"00",X"00",X"00",X"40",X"40",X"E0",X"FF",X"FF",X"FF",X"FF",X"7F",
		X"00",X"00",X"E0",X"F0",X"78",X"38",X"18",X"18",X"10",X"10",X"30",X"F0",X"E0",X"E0",X"E0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"0F",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"3C",X"7F",X"FF",X"FF",X"FF",X"FF",X"FD",
		X"00",X"00",X"03",X"1F",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"F0",X"F8",X"7C",X"3C",X"1C",X"18",X"18",X"38",X"70",X"E0",X"E0",X"E0",X"C0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"3F",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"39",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",
		X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"F8",X"FE",X"FE",X"3E",X"1C",X"1C",X"1C",X"38",X"30",X"F0",X"E0",X"C0",X"C0",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"0F",X"1F",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"39",X"7F",X"FF",X"FF",X"FF",X"FF",X"E7",
		X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"3F",X"FF",X"3F",X"1F",X"0F",X"0E",X"0E",X"3C",X"7C",X"F8",X"F0",X"E0",X"C0",X"80",
		X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"0F",X"1F",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"12",X"FF",X"FF",X"FF",X"FF",X"FF",X"C7",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"1F",X"FF",X"0F",X"07",X"03",X"03",X"07",X"1F",X"3E",X"FC",X"F8",X"F0",X"E0",X"C0",
		X"00",X"00",X"80",X"E0",X"E0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"3F",X"FF",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"06",X"7E",X"FF",X"FF",X"FF",X"FF",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"07",X"7F",X"0F",X"07",X"03",X"03",X"07",X"0F",X"3F",X"FE",X"FC",X"F8",X"E0",X"C0",
		X"00",X"00",X"F0",X"F8",X"F8",X"F8",X"F0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"06",X"0E",X"0E",X"1F",X"1F",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"C0",
		X"14",X"0C",X"2C",X"38",X"30",X"18",X"18",X"18",X"18",X"18",X"1C",X"1C",X"1C",X"0C",X"0E",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"03",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"28",X"3C",X"38",X"30",X"30",X"20",X"60",X"60",X"60",X"60",X"E0",X"C0",X"C0",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"70",X"7B",X"77",X"2F",X"0F",X"0F",X"0F",X"0F",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"0E",X"FE",X"EE",X"F4",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"70",X"7B",X"77",X"2F",X"0F",X"0F",X"0F",X"0F",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"0E",X"FE",X"EE",X"F4",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"1F",X"3F",X"3F",X"3F",X"2F",X"27",X"67",X"77",X"27",X"01",X"10",
		X"00",X"00",X"00",X"00",X"E0",X"F8",X"FC",X"FC",X"F6",X"F2",X"F2",X"F2",X"EE",X"CC",X"9C",X"78",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"0F",X"0F",X"0F",X"07",X"07",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"01",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"9C",X"0C",X"0C",X"04",X"00",X"00",X"60",X"60",
		X"00",X"00",X"00",X"00",X"03",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"07",X"07",X"00",X"18",
		X"00",X"00",X"00",X"00",X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"C0",X"40",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"03",X"01",X"03",X"02",X"06",X"06",X"06",X"0E",X"07",X"07",X"03",
		X"9C",X"0C",X"0C",X"88",X"08",X"00",X"20",X"E0",X"60",X"60",X"E0",X"E0",X"60",X"60",X"60",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"06",X"00",X"0A",X"08",
		X"0F",X"0F",X"07",X"06",X"07",X"07",X"03",X"39",X"FD",X"FF",X"FF",X"3E",X"3D",X"0D",X"0D",X"0B",
		X"F0",X"F0",X"F0",X"70",X"70",X"E0",X"C0",X"C0",X"C0",X"F0",X"F8",X"F8",X"FC",X"FC",X"DC",X"DC",
		X"3E",X"01",X"03",X"07",X"07",X"03",X"00",X"01",X"03",X"00",X"01",X"01",X"01",X"01",X"00",X"00",
		X"30",X"60",X"40",X"60",X"20",X"A0",X"A0",X"A0",X"E0",X"A0",X"A0",X"A0",X"E0",X"F0",X"F0",X"B0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"03",X"07",X"06",X"05",X"03",X"00",X"00",X"00",X"00",X"08",X"4C",X"20",
		X"3C",X"7C",X"FF",X"FD",X"BD",X"3B",X"3B",X"37",X"17",X"2F",X"2E",X"2C",X"0F",X"5D",X"59",X"B0",
		X"F8",X"10",X"20",X"F0",X"F8",X"F8",X"F0",X"E0",X"C0",X"80",X"30",X"30",X"80",X"80",X"C0",X"C0",
		X"01",X"00",X"01",X"01",X"00",X"00",X"02",X"07",X"01",X"01",X"03",X"03",X"03",X"03",X"03",X"01",
		X"1C",X"8C",X"AC",X"EC",X"88",X"88",X"98",X"18",X"10",X"30",X"30",X"30",X"E0",X"E0",X"60",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"0F",X"3C",
		X"07",X"0F",X"1F",X"1F",X"1F",X"15",X"10",X"08",X"0B",X"03",X"01",X"30",X"F8",X"FF",X"FB",X"C7",
		X"80",X"C0",X"F0",X"A0",X"10",X"20",X"40",X"40",X"20",X"E0",X"D0",X"30",X"F0",X"E0",X"C0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"07",X"00",X"78",X"07",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"04",X"08",X"10",
		X"FC",X"FE",X"7E",X"06",X"DE",X"18",X"90",X"90",X"20",X"20",X"40",X"11",X"10",X"20",X"11",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"0F",X"7F",X"FF",X"FE",X"FE",X"FC",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0D",X"01",X"03",X"26",X"7F",X"CF",X"9F",X"3D",X"3C",X"3C",X"1C",X"00",X"43",X"00",
		X"80",X"00",X"00",X"B0",X"78",X"FC",X"DC",X"DE",X"F6",X"E2",X"E1",X"E4",X"06",X"60",X"E0",X"70",
		X"27",X"33",X"33",X"33",X"17",X"1F",X"11",X"10",X"00",X"08",X"08",X"0C",X"06",X"06",X"07",X"07",
		X"90",X"A0",X"80",X"00",X"80",X"80",X"80",X"80",X"C0",X"C0",X"C0",X"40",X"60",X"60",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"05",X"08",X"04",X"02",X"03",X"01",X"03",X"01",X"00",X"00",X"04",X"0F",X"1B",X"17",X"1F",X"2F",
		X"F8",X"F8",X"A8",X"58",X"F0",X"F0",X"E0",X"A0",X"2E",X"5F",X"B7",X"F3",X"FA",X"FE",X"BC",X"9C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"70",X"18",X"48",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"03",X"03",X"07",X"07",X"07",X"07",X"03",X"01",X"01",X"01",X"01",X"01",X"02",X"02",X"02",
		X"C1",X"C3",X"82",X"82",X"84",X"84",X"00",X"80",X"80",X"80",X"A0",X"A0",X"E0",X"F0",X"F0",X"F0",
		X"00",X"00",X"07",X"3F",X"1F",X"0F",X"1E",X"7E",X"FC",X"F8",X"F0",X"E0",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"1E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"0E",X"1F",X"3F",X"FF",X"FF",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E3",X"FF",X"FF",X"FF",X"FF",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"03",X"03",X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DF",X"DF",X"DF",X"DF",X"3F",X"BF",X"7F",X"78",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"03",X"03",X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"F8",X"FF",X"FF",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"BF",X"BF",X"9F",X"9F",X"3F",X"BF",X"7F",X"78",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"07",X"07",X"07",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"F0",X"FF",X"FE",X"3E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"7F",X"3F",X"3F",X"7F",X"7F",X"FE",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"07",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FD",X"FC",X"FC",X"C0",X"FE",X"FD",X"7D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"7F",X"7F",X"7F",X"FE",X"FC",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"3F",X"3F",X"3F",X"1F",X"1F",X"0F",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F3",X"F7",X"F1",X"F1",X"01",X"FB",X"F7",X"F7",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FE",X"FE",X"FC",X"F8",X"F0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"7C",X"7F",X"3F",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EF",X"DF",X"C7",X"C7",X"07",X"EF",X"DF",X"DE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FE",X"FC",X"F8",X"F0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"F8",X"FF",X"7F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CF",X"9F",X"8F",X"8F",X"0F",X"DF",X"BF",X"BC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FE",X"FC",X"F8",X"F0",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"07",X"07",X"07",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FE",X"FC",X"FC",X"C0",X"FF",X"FE",X"3E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"7F",X"1F",X"1F",X"1F",X"3F",X"FF",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FE",X"F8",X"F0",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"0F",X"0F",X"0F",X"07",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"F9",X"F8",X"F8",X"C0",X"FE",X"FD",X"7D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"7F",X"7F",X"7F",X"FF",X"FC",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FC",X"F8",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"3F",X"3F",X"3F",X"3F",X"3F",X"1F",X"1F",X"1F",X"1E",X"1F",X"0F",X"06",X"00",X"00",
		X"86",X"8C",X"CC",X"C4",X"CC",X"CC",X"DC",X"DC",X"B8",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"07",X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"60",X"F8",X"73",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"07",X"07",X"07",X"03",X"00",X"00",
		X"00",X"00",X"E0",X"E0",X"F1",X"F1",X"F1",X"F1",X"F3",X"F3",X"E0",X"C0",X"80",X"00",X"00",X"00",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"07",X"07",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"C0",X"00",X"00",
		X"07",X"27",X"63",X"77",X"77",X"37",X"17",X"03",X"03",X"03",X"03",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"DC",X"FE",X"FE",X"FE",X"FC",X"F8",X"B0",X"C0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"07",X"07",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"C0",X"00",X"00",
		X"07",X"27",X"63",X"73",X"77",X"37",X"17",X"07",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"DC",X"FE",X"FE",X"FE",X"FC",X"B8",X"B0",X"C0",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"03",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"04",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"00",X"00",X"00",X"00",
		X"1F",X"1F",X"1F",X"0F",X"07",X"17",X"17",X"11",X"01",X"01",X"01",X"11",X"0D",X"00",X"01",X"00",
		X"F8",X"F8",X"78",X"78",X"70",X"08",X"F8",X"0C",X"0C",X"1C",X"1C",X"28",X"C0",X"00",X"00",X"00",
		X"0F",X"0F",X"37",X"77",X"37",X"3F",X"77",X"30",X"38",X"1F",X"1F",X"0F",X"07",X"03",X"13",X"13",
		X"F0",X"F0",X"FC",X"FE",X"F2",X"E6",X"CE",X"5E",X"FE",X"FC",X"F8",X"78",X"70",X"E0",X"88",X"F8",
		X"11",X"01",X"01",X"01",X"0D",X"00",X"00",X"01",X"00",X"00",X"0C",X"0C",X"0C",X"0E",X"0E",X"0F",
		X"8C",X"0C",X"1C",X"1C",X"20",X"80",X"00",X"00",X"00",X"60",X"60",X"60",X"60",X"60",X"60",X"E0",
		X"07",X"07",X"00",X"18",X"7F",X"FF",X"3F",X"0F",X"0F",X"07",X"07",X"03",X"13",X"11",X"01",X"09",
		X"E0",X"C0",X"40",X"F8",X"FE",X"FF",X"7C",X"70",X"70",X"70",X"F0",X"E0",X"48",X"08",X"1C",X"3C",
		X"00",X"01",X"07",X"04",X"04",X"04",X"04",X"04",X"06",X"06",X"07",X"07",X"07",X"07",X"07",X"07",
		X"60",X"60",X"E0",X"C0",X"E0",X"E0",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"E0",X"E0",X"E0",
		X"3F",X"7F",X"7F",X"7F",X"3F",X"1F",X"17",X"17",X"07",X"13",X"13",X"01",X"0C",X"01",X"07",X"03",
		X"FC",X"FE",X"FE",X"7F",X"7B",X"79",X"F8",X"F0",X"B0",X"38",X"08",X"1C",X"FC",X"7C",X"3C",X"9C",
		X"01",X"01",X"01",X"01",X"01",X"05",X"04",X"06",X"06",X"06",X"06",X"07",X"07",X"07",X"07",X"07",
		X"60",X"60",X"60",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"08",X"04",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"03",X"04",X"04",X"04",X"01",X"10",X"30",X"38",X"38",X"1A",X"02",X"00",X"00",X"00",X"02",
		X"D8",X"58",X"18",X"58",X"B0",X"B0",X"B0",X"B0",X"90",X"58",X"D8",X"C8",X"E8",X"E8",X"E8",X"78",
		X"00",X"02",X"02",X"02",X"02",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"90",X"90",X"90",X"D0",X"D0",X"70",X"70",X"70",X"70",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"03",X"03",X"03",X"03",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"F8",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"B0",X"21",X"A3",X"E3",X"47",X"97",X"17",X"07",X"07",X"03",X"10",X"08",X"04",X"02",X"02",X"01",
		X"E0",X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",X"38",X"7C",X"3E",X"3E",X"1E",
		X"09",X"08",X"08",X"08",X"19",X"19",X"1F",X"1F",X"3F",X"3F",X"3E",X"3E",X"3C",X"18",X"00",X"00",
		X"40",X"40",X"C0",X"C0",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"70",X"60",X"30",X"00",X"00",X"00",X"00",X"00",X"60",X"31",X"A1",X"B1",X"00",X"00",X"00",X"00",
		X"0E",X"7E",X"17",X"07",X"03",X"47",X"6F",X"3D",X"FE",X"FE",X"E6",X"FE",X"FF",X"FF",X"7F",X"7F",
		X"C0",X"E0",X"C0",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"E0",X"F0",X"F8",
		X"00",X"07",X"3F",X"7F",X"FF",X"FF",X"7E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"39",X"1F",X"3F",X"FF",X"F8",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FC",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"1F",X"7F",X"2F",X"47",X"25",X"12",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"40",X"C0",X"80",
		X"09",X"01",X"03",X"13",X"13",X"11",X"18",X"0F",X"00",X"06",X"0F",X"0F",X"07",X"07",X"07",X"07",
		X"E0",X"E8",X"B0",X"F0",X"F4",X"C4",X"3C",X"F4",X"EC",X"CC",X"0C",X"08",X"08",X"18",X"90",X"90",
		X"02",X"02",X"02",X"03",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"98",X"F8",X"F8",X"FC",X"FC",X"FC",X"7C",X"7C",X"38",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"F0",X"F8",
		X"0B",X"03",X"00",X"01",X"10",X"30",X"00",X"00",X"00",X"00",X"0C",X"08",X"01",X"01",X"03",X"03",
		X"04",X"0E",X"3E",X"1E",X"E3",X"7F",X"EF",X"FD",X"FD",X"3C",X"00",X"3F",X"BE",X"D8",X"C1",X"C1",
		X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"03",X"03",X"02",X"02",X"02",X"02",X"02",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"70",X"F0",X"30",X"30",X"10",X"10",X"10",X"10",X"30",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"07",X"07",X"07",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"38",X"78",X"F8",X"F8",X"E0",X"CE",X"FE",X"FE",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"7F",X"7F",X"FE",X"F0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"F0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
