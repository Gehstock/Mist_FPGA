library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity nrx_wav_rom is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of nrx_wav_rom is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"80",X"7F",X"7F",X"79",X"6B",X"71",X"7F",X"79",X"95",X"BF",X"D3",X"BE",X"BF",X"B9",X"B5",X"B1",
		X"AD",X"AA",X"A6",X"A3",X"A0",X"9D",X"9A",X"98",X"95",X"93",X"90",X"76",X"20",X"00",X"16",X"01",
		X"0E",X"12",X"1B",X"1F",X"25",X"2A",X"2F",X"34",X"38",X"3C",X"40",X"44",X"47",X"4B",X"4E",X"51",
		X"54",X"56",X"58",X"5A",X"5C",X"68",X"86",X"7E",X"4F",X"66",X"62",X"64",X"67",X"67",X"6A",X"6A",
		X"6D",X"6D",X"6F",X"71",X"81",X"BE",X"FF",X"FD",X"F6",X"FF",X"F7",X"FD",X"F7",X"F9",X"F0",X"ED",
		X"E7",X"E3",X"DD",X"D6",X"AE",X"3E",X"07",X"3E",X"2A",X"38",X"38",X"3D",X"40",X"43",X"46",X"49",
		X"4C",X"4E",X"50",X"52",X"54",X"56",X"61",X"A2",X"FF",X"FD",X"EF",X"FE",X"E8",X"EF",X"E1",X"E3",
		X"D9",X"D8",X"D1",X"CD",X"BC",X"8C",X"5A",X"83",X"D2",X"C4",X"B3",X"BC",X"AC",X"B0",X"A6",X"A7",
		X"A0",X"9F",X"95",X"65",X"01",X"00",X"0E",X"00",X"14",X"12",X"1E",X"20",X"27",X"2A",X"30",X"33",
		X"39",X"43",X"4B",X"3B",X"42",X"47",X"45",X"4D",X"4C",X"57",X"7D",X"AC",X"75",X"55",X"99",X"FA",
		X"FF",X"EC",X"F9",X"C7",X"88",X"4A",X"40",X"67",X"D5",X"FF",X"E5",X"E4",X"E0",X"D7",X"D2",X"B6",
		X"9B",X"BE",X"D0",X"B5",X"BF",X"B1",X"B3",X"AB",X"A9",X"A4",X"9D",X"83",X"5E",X"42",X"23",X"04",
		X"00",X"0F",X"12",X"1B",X"20",X"26",X"2B",X"30",X"34",X"38",X"40",X"4A",X"42",X"41",X"4C",X"49",
		X"51",X"51",X"5D",X"96",X"FF",X"FF",X"ED",X"FA",X"E5",X"E9",X"DD",X"DC",X"D3",X"D1",X"CA",X"C7",
		X"C1",X"BE",X"B9",X"AC",X"6C",X"00",X"00",X"22",X"12",X"28",X"23",X"2F",X"2F",X"37",X"38",X"3E",
		X"40",X"44",X"46",X"49",X"4C",X"4F",X"51",X"56",X"71",X"CD",X"FF",X"F4",X"F9",X"F2",X"E9",X"E8",
		X"DE",X"DC",X"D4",X"D1",X"CA",X"C6",X"C1",X"BC",X"A5",X"4C",X"00",X"16",X"1E",X"1B",X"2B",X"27",
		X"32",X"31",X"39",X"3A",X"40",X"42",X"47",X"48",X"4C",X"4E",X"50",X"52",X"55",X"57",X"5F",X"91",
		X"FB",X"FF",X"EC",X"FF",X"EB",X"EF",X"E4",X"E0",X"C1",X"7A",X"36",X"29",X"32",X"3A",X"3A",X"41",
		X"41",X"46",X"47",X"4B",X"4C",X"4F",X"51",X"53",X"56",X"6B",X"BE",X"FF",X"F6",X"F7",X"FA",X"EA",
		X"ED",X"E1",X"E0",X"D8",X"D5",X"CE",X"CB",X"C5",X"C1",X"BC",X"B8",X"B3",X"AF",X"9A",X"45",X"00",
		X"0A",X"12",X"11",X"20",X"1E",X"29",X"29",X"31",X"33",X"38",X"3A",X"3F",X"41",X"45",X"47",X"4B",
		X"53",X"6E",X"98",X"B6",X"D2",X"E9",X"F5",X"F1",X"E7",X"E4",X"DD",X"D8",X"D2",X"CD",X"C8",X"C3",
		X"BF",X"BA",X"B5",X"A1",X"56",X"00",X"05",X"19",X"15",X"22",X"23",X"2B",X"2D",X"33",X"36",X"3B",
		X"3E",X"42",X"46",X"49",X"4B",X"4D",X"4F",X"54",X"77",X"E0",X"FF",X"EA",X"FA",X"E8",X"E8",X"E0",
		X"DC",X"D6",X"D2",X"C9",X"A2",X"4C",X"14",X"1E",X"29",X"33",X"67",X"B1",X"93",X"3E",X"2F",X"30",
		X"3B",X"3B",X"5C",X"B8",X"FF",X"E1",X"CA",X"B2",X"CC",X"E6",X"C4",X"D1",X"C2",X"C2",X"BA",X"B8",
		X"B2",X"AF",X"AA",X"A7",X"A2",X"8D",X"4D",X"33",X"6F",X"64",X"28",X"00",X"0E",X"12",X"16",X"21",
		X"23",X"2B",X"2D",X"33",X"36",X"3B",X"44",X"7F",X"F4",X"FF",X"D3",X"EA",X"D2",X"D8",X"CB",X"CB",
		X"C2",X"C0",X"B9",X"B5",X"AA",X"84",X"40",X"15",X"06",X"10",X"1C",X"1E",X"28",X"2B",X"31",X"34",
		X"3E",X"74",X"E7",X"FC",X"CF",X"E3",X"CE",X"D2",X"C7",X"C5",X"BF",X"BC",X"B7",X"B3",X"A5",X"79",
		X"59",X"87",X"92",X"97",X"9E",X"97",X"8E",X"59",X"02",X"00",X"13",X"08",X"1D",X"1B",X"27",X"29",
		X"31",X"33",X"39",X"3C",X"44",X"6E",X"D5",X"F6",X"DA",X"ED",X"D8",X"DB",X"D1",X"CF",X"C8",X"C5",
		X"BF",X"BC",X"B7",X"B3",X"AF",X"AB",X"A7",X"A4",X"A0",X"9D",X"9A",X"98",X"95",X"8B",X"63",X"32",
		X"25",X"0D",X"02",X"06",X"0A",X"13",X"1A",X"20",X"26",X"2C",X"31",X"36",X"3A",X"3E",X"42",X"46",
		X"4F",X"84",X"F4",X"FF",X"E0",X"F2",X"DE",X"E0",X"D6",X"D4",X"CD",X"C9",X"C4",X"BF",X"BA",X"B6",
		X"B2",X"AE",X"A8",X"8B",X"2F",X"00",X"0F",X"0E",X"17",X"20",X"24",X"2D",X"30",X"36",X"39",X"3E",
		X"47",X"73",X"CF",X"FD",X"E9",X"E3",X"DE",X"D7",X"D3",X"CD",X"C9",X"C4",X"B7",X"79",X"0D",X"05",
		X"29",X"1B",X"2E",X"2B",X"35",X"36",X"3C",X"3E",X"43",X"45",X"4A",X"5E",X"AB",X"FF",X"FC",X"EB",
		X"EE",X"E2",X"E0",X"D7",X"D3",X"CD",X"C8",X"C3",X"BF",X"BA",X"B6",X"AE",X"84",X"21",X"00",X"1A",
		X"15",X"20",X"25",X"2A",X"2F",X"33",X"38",X"3B",X"40",X"43",X"47",X"4A",X"4D",X"57",X"92",X"FF",
		X"FF",X"E8",X"F7",X"E2",X"E6",X"D9",X"D9",X"D0",X"CE",X"C1",X"93",X"34",X"09",X"20",X"24",X"29",
		X"2F",X"33",X"39",X"3C",X"41",X"4C",X"85",X"F0",X"FF",X"E1",X"EC",X"DC",X"DB",X"D3",X"CF",X"C9",
		X"C3",X"B9",X"8C",X"22",X"00",X"23",X"1B",X"27",X"2B",X"30",X"35",X"3B",X"51",X"8C",X"C9",X"E5",
		X"EE",X"DD",X"DB",X"D4",X"CE",X"C9",X"BC",X"89",X"20",X"01",X"26",X"21",X"3D",X"5C",X"74",X"88",
		X"9A",X"A6",X"AF",X"B4",X"B3",X"93",X"3E",X"12",X"33",X"2F",X"36",X"3A",X"3D",X"41",X"43",X"47",
		X"49",X"4D",X"4F",X"52",X"54",X"5A",X"7A",X"C0",X"F4",X"FF",X"FA",X"F5",X"F0",X"E8",X"E4",X"DD",
		X"D8",X"D2",X"CE",X"C8",X"C4",X"BF",X"BB",X"B7",X"B3",X"AE",X"9E",X"5B",X"00",X"00",X"14",X"11",
		X"1F",X"20",X"29",X"2B",X"31",X"34",X"39",X"3C",X"40",X"43",X"46",X"48",X"4C",X"57",X"84",X"CB",
		X"F3",X"FD",X"F0",X"EB",X"E8",X"E1",X"DE",X"D7",X"D3",X"CD",X"C8",X"C3",X"BE",X"BA",X"B5",X"B1",
		X"AD",X"A9",X"A5",X"A1",X"9E",X"9B",X"98",X"88",X"42",X"00",X"06",X"09",X"03",X"15",X"14",X"20",
		X"22",X"2A",X"2D",X"33",X"36",X"3C",X"3F",X"43",X"45",X"49",X"4E",X"6F",X"C5",X"FF",X"F6",X"EC",
		X"E9",X"E2",X"DD",X"D7",X"D2",X"CD",X"C6",X"A7",X"4D",X"0D",X"32",X"31",X"2A",X"2B",X"33",X"36",
		X"39",X"3D",X"40",X"44",X"46",X"4A",X"4E",X"5D",X"71",X"5A",X"4B",X"5B",X"55",X"5C",X"5A",X"5E",
		X"62",X"75",X"90",X"A7",X"C0",X"D8",X"EF",X"FD",X"FB",X"F8",X"F5",X"ED",X"EA",X"E3",X"DF",X"D9",
		X"D4",X"CF",X"CA",X"C5",X"C0",X"BC",X"B6",X"A6",X"5C",X"00",X"05",X"1E",X"13",X"26",X"22",X"2D",
		X"2D",X"34",X"36",X"3B",X"3D",X"41",X"44",X"47",X"4A",X"60",X"B7",X"FF",X"F1",X"EA",X"ED",X"DE",
		X"E0",X"D5",X"D5",X"CD",X"CB",X"C5",X"C1",X"B3",X"9A",X"A1",X"C0",X"AA",X"AC",X"A6",X"A2",X"9F",
		X"9A",X"98",X"94",X"92",X"88",X"6E",X"4B",X"28",X"00",X"00",X"07",X"02",X"0F",X"13",X"1C",X"20",
		X"27",X"2F",X"4A",X"63",X"42",X"2C",X"45",X"3E",X"46",X"47",X"4E",X"6F",X"B6",X"BD",X"90",X"A9",
		X"DE",X"FF",X"E0",X"E8",X"DD",X"DA",X"D5",X"D0",X"CB",X"C6",X"C1",X"BC",X"B8",X"B3",X"AE",X"9A",
		X"51",X"00",X"03",X"13",X"13",X"1F",X"22",X"2A",X"2D",X"33",X"36",X"3B",X"40",X"5B",X"AF",X"FD",
		X"EE",X"E1",X"E1",X"D6",X"D3",X"CD",X"C9",X"C2",X"AB",X"66",X"22",X"28",X"61",X"8C",X"7B",X"3E",
		X"18",X"33",X"63",X"A9",X"CE",X"DC",X"CE",X"C9",X"C5",X"BE",X"BB",X"B5",X"B1",X"AD",X"A9",X"A3",
		X"88",X"32",X"00",X"08",X"09",X"12",X"1B",X"20",X"2F",X"33",X"2D",X"36",X"3B",X"3D",X"4D",X"7A",
		X"BF",X"E0",X"DC",X"9A",X"67",X"4C",X"36",X"3F",X"43",X"46",X"4C",X"67",X"C0",X"FF",X"F4",X"EC",
		X"EB",X"E0",X"DB",X"CB",X"CC",X"D3",X"C7",X"C4",X"C0",X"BA",X"B6",X"B0",X"AD",X"A9",X"A6",X"A2",
		X"9F",X"9C",X"99",X"97",X"94",X"89",X"54",X"00",X"00",X"0D",X"00",X"0F",X"11",X"1C",X"20",X"2D",
		X"3B",X"34",X"2B",X"3C",X"38",X"40",X"41",X"45",X"48",X"4B",X"55",X"8B",X"F3",X"FF",X"EA",X"F4",
		X"E5",X"E5",X"DC",X"D9",X"D3",X"CE",X"C5",X"A4",X"57",X"1E",X"17",X"23",X"2A",X"2C",X"34",X"37",
		X"53",X"9D",X"EA",X"ED",X"DE",X"DA",X"D5",X"CE",X"CA",X"C4",X"C0",X"BA",X"A8",X"66",X"0D",X"03",
		X"1A",X"1B",X"24",X"29",X"2E",X"33",X"3F",X"6F",X"BF",X"E6",X"CE",X"98",X"89",X"B0",X"E3",X"D6",
		X"C9",X"CA",X"BF",X"BE",X"B0",X"94",X"86",X"AC",X"A4",X"6E",X"21",X"02",X"1A",X"4D",X"72",X"8F",
		X"A8",X"B8",X"C0",X"BC",X"AD",X"7D",X"27",X"03",X"18",X"3B",X"51",X"38",X"19",X"2F",X"30",X"34",
		X"3F",X"62",X"AF",X"E3",X"ED",X"DF",X"CD",X"A2",X"6C",X"53",X"3C",X"52",X"9E",X"DA",X"DA",X"CF",
		X"CA",X"C6",X"BF",X"B4",X"A0",X"B0",X"BC",X"A1",X"7A",X"2C",X"0B",X"06",X"17",X"1C",X"2C",X"5D",
		X"A3",X"CB",X"D8",X"C9",X"AA",X"76",X"67",X"9D",X"BE",X"B3",X"7B",X"40",X"22",X"11",X"1E",X"29",
		X"4D",X"9B",X"CF",X"DB",X"CF",X"C8",X"C0",X"9A",X"60",X"37",X"1F",X"18",X"27",X"2A",X"31",X"35",
		X"3A",X"3E",X"42",X"45",X"4A",X"59",X"7C",X"B7",X"FF",X"FF",X"E5",X"EE",X"DE",X"DF",X"D5",X"D2",
		X"CB",X"C7",X"C1",X"BD",X"B8",X"B5",X"B0",X"AD",X"AA",X"A7",X"A4",X"9F",X"89",X"3A",X"00",X"08",
		X"09",X"0C",X"1A",X"1B",X"25",X"28",X"30",X"32",X"38",X"3B",X"40",X"43",X"46",X"49",X"50",X"6C",
		X"B9",X"FF",X"FB",X"EB",X"EF",X"E2",X"E2",X"D8",X"D3",X"CD",X"CE",X"C5",X"C2",X"BC",X"B8",X"B3",
		X"B0",X"AB",X"A4",X"82",X"2E",X"05",X"1E",X"13",X"12",X"17",X"21",X"24",X"2C",X"2F",X"35",X"38",
		X"3D",X"40",X"44",X"47",X"4B",X"4E",X"51",X"55",X"62",X"8F",X"CC",X"EF",X"FF",X"F7",X"F1",X"EC",
		X"E5",X"E1",X"DA",X"D6",X"D0",X"CB",X"C6",X"C1",X"BD",X"B1",X"7F",X"28",X"04",X"14",X"1D",X"21",
		X"29",X"2D",X"32",X"36",X"3A",X"3E",X"41",X"44",X"48",X"56",X"85",X"AA",X"8B",X"8F",X"C0",X"FC",
		X"F6",X"E3",X"E8",X"DB",X"DA",X"C7",X"9D",X"6A",X"67",X"92",X"C2",X"BD",X"8D",X"53",X"50",X"77",
		X"AB",X"BC",X"CA",X"BE",X"B5",X"8B",X"40",X"13",X"0C",X"1B",X"21",X"25",X"2C",X"2F",X"38",X"54",
		X"A1",X"E2",X"E9",X"DB",X"D6",X"D2",X"CB",X"C7",X"BA",X"93",X"4D",X"24",X"13",X"1D",X"27",X"28",
		X"37",X"5B",X"8C",X"73",X"51",X"4C",X"3D",X"3F",X"40",X"46",X"4D",X"74",X"CA",X"FF",X"F0",X"E9",
		X"E6",X"DD",X"DA",X"D3",X"CF",X"C9",X"C5",X"C0",X"B9",X"9E",X"5B",X"37",X"41",X"2B",X"2C",X"24",
		X"24",X"26",X"2E",X"31",X"35",X"39",X"3D",X"40",X"44",X"49",X"61",X"A6",X"EB",X"F9",X"EE",X"E5",
		X"E3",X"D6",X"BB",X"91",X"9E",X"CD",X"D2",X"C4",X"C4",X"BD",X"B9",X"B4",X"B0",X"AC",X"A8",X"A5",
		X"A1",X"96",X"74",X"32",X"00",X"02",X"0B",X"0B",X"1A",X"1A",X"25",X"28",X"2F",X"32",X"37",X"3A",
		X"3E",X"47",X"74",X"D4",X"FF",X"E4",X"E4",X"DD",X"D7",X"D1",X"C3",X"AE",X"9E",X"99",X"AF",X"CB",
		X"B9",X"B7",X"B5",X"A9",X"91",X"62",X"4E",X"5F",X"97",X"B0",X"AB",X"A5",X"A3",X"9A",X"76",X"36",
		X"2C",X"52",X"60",X"6C",X"75",X"78",X"79",X"76",X"72",X"6B",X"64",X"56",X"2E",X"01",X"11",X"1E",
		X"1E",X"2A",X"2B",X"33",X"36",X"3B",X"3E",X"42",X"49",X"6B",X"B3",X"CE",X"AA",X"A0",X"95",X"8D",
		X"89",X"86",X"86",X"88",X"8C",X"90",X"95",X"9D",X"B5",X"E5",X"ED",X"D5",X"DB",X"CF",X"CE",X"C7",
		X"C4",X"BE",X"BA",X"B5",X"A8",X"8F",X"7A",X"5A",X"19",X"00",X"16",X"18",X"1F",X"27",X"2A",X"31",
		X"35",X"3A",X"3D",X"41",X"45",X"56",X"9C",X"FA",X"FA",X"E4",X"E8",X"DC",X"DA",X"D3",X"D0",X"CA",
		X"C6",X"C1",X"BC",X"B8",X"B3",X"AF",X"AB",X"A6",X"92",X"50",X"05",X"00",X"0C",X"11",X"1B",X"20",
		X"26",X"2B",X"30",X"35",X"39",X"3D",X"4D",X"82",X"C5",X"E6",X"EF",X"D1",X"AA",X"93",X"B3",X"D8",
		X"D1",X"B1",X"7C",X"63",X"80",X"A5",X"A6",X"7F",X"48",X"3C",X"57",X"87",X"9D",X"B4",X"C0",X"C6",
		X"C2",X"BC",X"B8",X"B3",X"AB",X"9C",X"8A",X"7A",X"69",X"54",X"2B",X"00",X"0C",X"1C",X"1A",X"27",
		X"27",X"30",X"32",X"38",X"3B",X"40",X"43",X"49",X"61",X"98",X"C5",X"DF",X"DB",X"A7",X"89",X"91",
		X"BF",X"E1",X"E3",X"DC",X"D4",X"D2",X"CA",X"C7",X"BC",X"99",X"4E",X"1B",X"12",X"1F",X"28",X"2A",
		X"33",X"34",X"3A",X"3C",X"40",X"43",X"47",X"54",X"94",X"F5",X"FF",X"E8",X"EC",X"E1",X"DE",X"D7",
		X"D3",X"CD",X"C8",X"C3",X"BF",X"BA",X"B6",X"B2",X"AC",X"99",X"54",X"00",X"00",X"10",X"12",X"1D",
		X"21",X"29",X"2D",X"34",X"38",X"3C",X"3F",X"43",X"45",X"48",X"4C",X"62",X"A3",X"E7",X"FC",X"F5",
		X"E9",X"E8",X"DE",X"D6",X"B4",X"85",X"65",X"4D",X"46",X"6C",X"A3",X"B4",X"9E",X"71",X"5B",X"46",
		X"39",X"33",X"33",X"3B",X"48",X"7D",X"CB",X"EE",X"E3",X"C4",X"BC",X"D1",X"DB",X"C8",X"C9",X"BF",
		X"B3",X"B2",X"BD",X"B0",X"A4",X"76",X"3F",X"22",X"09",X"0F",X"28",X"52",X"81",X"9C",X"B5",X"B8",
		X"93",X"5B",X"48",X"5B",X"84",X"8B",X"6F",X"40",X"34",X"4E",X"7E",X"8D",X"77",X"4C",X"39",X"2E",
		X"34",X"3D",X"54",X"92",X"BE",X"B0",X"92",X"83",X"76",X"6D",X"69",X"67",X"6A",X"7B",X"B2",X"ED",
		X"EA",X"DA",X"DB",X"D1",X"CE",X"C7",X"C3",X"BE",X"B8",X"9E",X"5C",X"1F",X"0D",X"14",X"22",X"22",
		X"2C",X"2D",X"34",X"37",X"41",X"65",X"AF",X"E0",X"ED",X"E2",X"D9",X"D7",X"C8",X"BE",X"C6",X"C8",
		X"B7",X"A2",X"6A",X"5D",X"7A",X"8C",X"7C",X"4D",X"21",X"14",X"17",X"25",X"26",X"38",X"5D",X"7C",
		X"60",X"4E",X"49",X"41",X"47",X"64",X"AB",X"E3",X"F1",X"E5",X"DD",X"DA",X"D2",X"CF",X"C9",X"C4",
		X"B4",X"83",X"41",X"20",X"16",X"36",X"53",X"50",X"32",X"25",X"37",X"35",X"3D",X"40",X"44",X"47",
		X"4E",X"6F",X"BF",X"F9",X"F9",X"EC",X"E7",X"E2",X"DA",X"D6",X"D0",X"CB",X"BB",X"8E",X"53",X"32",
		X"1A",X"1D",X"2A",X"38",X"65",X"90",X"AB",X"C6",X"D4",X"D6",X"CC",X"C8",X"C3",X"BE",X"BA",X"B6",
		X"B1",X"A5",X"90",X"7B",X"6A",X"58",X"47",X"28",X"04",X"0B",X"1D",X"1B",X"28",X"29",X"31",X"34",
		X"3F",X"5D",X"8C",X"A9",X"BB",X"A9",X"7E",X"71",X"86",X"B3",X"C5",X"B2",X"88",X"78",X"8D",X"B8",
		X"CF",X"D4",X"CB",X"C5",X"BC",X"96",X"62",X"40",X"27",X"1C",X"38",X"69",X"84",X"79",X"57",X"46",
		X"3A",X"32",X"3C",X"64",X"A8",X"D4",X"E8",X"DF",X"D6",X"D4",X"C8",X"B3",X"87",X"68",X"5A",X"6C",
		X"9A",X"A9",X"97",X"6B",X"52",X"3E",X"2D",X"26",X"24",X"2C",X"37",X"5C",X"A3",X"D3",X"E4",X"DB",
		X"D0",X"CF",X"C6",X"C3",X"BC",X"B9",X"B3",X"AD",X"90",X"51",X"35",X"45",X"37",X"20",X"0C",X"20",
		X"24",X"29",X"30",X"38",X"51",X"71",X"89",X"9D",X"A7",X"91",X"63",X"49",X"3B",X"3C",X"44",X"44",
		X"4D",X"6C",X"AD",X"CC",X"BB",X"AC",X"BA",X"E2",X"F4",X"DF",X"E0",X"D5",X"C0",X"A0",X"8B",X"79",
		X"6A",X"63",X"6E",X"A0",X"CB",X"CD",X"B7",X"99",X"94",X"B1",X"C2",X"B1",X"A3",X"7C",X"69",X"85",
		X"9B",X"A3",X"A8",X"A2",X"9F",X"9C",X"96",X"7C",X"3E",X"0A",X"00",X"09",X"1A",X"2C",X"3B",X"48",
		X"56",X"60",X"68",X"5F",X"39",X"22",X"32",X"34",X"38",X"3D",X"40",X"43",X"46",X"52",X"81",X"CD",
		X"F5",X"F8",X"E9",X"E6",X"E0",X"DA",X"D5",X"D0",X"CB",X"C5",X"B5",X"8C",X"62",X"4B",X"43",X"64",
		X"86",X"97",X"AA",X"B1",X"A7",X"7A",X"4C",X"42",X"56",X"73",X"6E",X"50",X"2A",X"23",X"27",X"31",
		X"32",X"39",X"3B",X"40",X"44",X"58",X"95",X"DD",X"F5",X"EF",X"E2",X"E1",X"D8",X"D5",X"C8",X"AD",
		X"90",X"99",X"B8",X"C0",X"AA",X"80",X"60",X"67",X"84",X"95",X"9F",X"A7",X"A1",X"83",X"4A",X"2B",
		X"2C",X"48",X"5A",X"67",X"75",X"76",X"61",X"33",X"20",X"2B",X"47",X"65",X"7C",X"90",X"A0",X"AB",
		X"B4",X"B9",X"BB",X"BA",X"B1",X"8F",X"55",X"30",X"20",X"27",X"31",X"31",X"39",X"3A",X"40",X"4E",
		X"7E",X"BC",X"E0",X"F3",X"E8",X"DF",X"DD",X"D4",X"D0",X"C1",X"B4",X"BC",X"BD",X"9B",X"69",X"44",
		X"45",X"5D",X"6A",X"58",X"34",X"1F",X"2E",X"51",X"72",X"88",X"9E",X"AC",X"B8",X"BE",X"C2",X"BF",
		X"AE",X"7E",X"4C",X"3B",X"48",X"63",X"61",X"47",X"29",X"2E",X"44",X"68",X"87",X"9F",X"B3",X"B4",
		X"96",X"6F",X"5C",X"48",X"3F",X"45",X"6F",X"A0",X"B1",X"A4",X"8A",X"8F",X"AF",X"D7",X"DD",X"D6",
		X"CF",X"CC",X"C3",X"AF",X"81",X"5D",X"44",X"2E",X"23",X"20",X"2A",X"2F",X"33",X"38",X"3B",X"41",
		X"55",X"93",X"D9",X"F1",X"EB",X"DD",X"DB",X"D6",X"D3",X"CA",X"C8",X"C1",X"BE",X"B8",X"B4",X"AF",
		X"A3",X"7D",X"4D",X"30",X"17",X"11",X"2C",X"53",X"69",X"7F",X"8F",X"9A",X"A2",X"A5",X"A6",X"A3",
		X"9E",X"97",X"8E",X"85",X"7B",X"71",X"66",X"5D",X"54",X"4D",X"48",X"44",X"41",X"3F",X"3F",X"41",
		X"43",X"47",X"4D",X"53",X"57",X"4B",X"38",X"40",X"46",X"47",X"56",X"5E",X"51",X"4E",X"68",X"90",
		X"BF",X"C3",X"B3",X"A3",X"A0",X"98",X"9C",X"B3",X"E6",X"F7",X"E8",X"E4",X"DF",X"D8",X"D3",X"CD",
		X"C9",X"C3",X"BF",X"BA",X"B6",X"B1",X"9C",X"67",X"32",X"16",X"08",X"17",X"1D",X"22",X"2E",X"37",
		X"30",X"32",X"3B",X"3A",X"42",X"4F",X"80",X"B9",X"C7",X"B9",X"AE",X"AA",X"A3",X"A1",X"9E",X"9D",
		X"A0",X"B8",X"DD",X"DB",X"CC",X"CE",X"C4",X"C2",X"BB",X"B8",X"B2",X"AF",X"AB",X"A7",X"A1",X"95",
		X"83",X"74",X"61",X"3F",X"0E",X"00",X"0B",X"0E",X"17",X"1D",X"24",X"30",X"44",X"56",X"62",X"5C",
		X"3F",X"34",X"3E",X"40",X"43",X"47",X"4B",X"5D",X"90",X"C0",X"BE",X"B4",X"BD",X"DD",X"F8",X"E9",
		X"E3",X"E0",X"D3",X"BF",X"A5",X"96",X"84",X"79",X"78",X"95",X"BB",X"C7",X"C4",X"BB",X"B9",X"B3",
		X"B0",X"AB",X"A8",X"A4",X"A0",X"95",X"7C",X"64",X"51",X"3D",X"27",X"08",X"00",X"11",X"14",X"1D",
		X"22",X"28",X"2E",X"33",X"38",X"3D",X"49",X"73",X"B3",X"DB",X"EF",X"E7",X"DD",X"DB",X"D2",X"CF",
		X"C8",X"C4",X"BE",X"BB",X"B6",X"B2",X"AE",X"A9",X"9C",X"85",X"70",X"5E",X"4C",X"3C",X"28",X"0D",
		X"07",X"1A",X"1B",X"24",X"28",X"2E",X"33",X"37",X"3C",X"3F",X"43",X"46",X"4A",X"4E",X"59",X"7A",
		X"A4",X"C1",X"DD",X"F1",X"F7",X"EE",X"E8",X"E4",X"DD",X"D8",X"D2",X"CE",X"C8",X"C4",X"BF",X"BA",
		X"B5",X"B0",X"AA",X"91",X"5C",X"3D",X"30",X"10",X"09",X"17",X"1F",X"21",X"2A",X"2D",X"33",X"36",
		X"3B",X"3E",X"42",X"49",X"66",X"A1",X"BF",X"B3",X"AF",X"AB",X"A7",X"A5",X"A2",X"A0",X"A0",X"B1",
		X"D8",X"E5",X"D4",X"D3",X"CC",X"C7",X"C1",X"B3",X"8F",X"62",X"49",X"3F",X"55",X"65",X"5D",X"41",
		X"27",X"24",X"29",X"32",X"34",X"3A",X"3C",X"44",X"5A",X"90",X"BE",X"DB",X"EF",X"E5",X"D6",X"BE",
		X"A2",X"90",X"7F",X"83",X"A0",X"B7",X"B2",X"96",X"79",X"7A",X"8E",X"A2",X"98",X"7A",X"5A",X"4B",
		X"38",X"30",X"28",X"2A",X"2F",X"35",X"3E",X"61",X"99",X"C0",X"DC",X"E7",X"DB",X"D5",X"CA",X"B5",
		X"B4",X"C6",X"BE",X"A6",X"7E",X"63",X"69",X"7B",X"83",X"87",X"8B",X"8A",X"88",X"83",X"78",X"58",
		X"2D",X"17",X"15",X"21",X"26",X"2B",X"33",X"3E",X"47",X"3C",X"44",X"63",X"92",X"B6",X"D0",X"E6",
		X"E8",X"D9",X"BD",X"A6",X"AD",X"C3",X"C4",X"AE",X"86",X"6C",X"56",X"44",X"39",X"30",X"2D",X"2D",
		X"32",X"38",X"40",X"4C",X"59",X"67",X"75",X"84",X"99",X"C3",X"F1",X"EE",X"E0",X"E0",X"D7",X"D3",
		X"CD",X"C8",X"C3",X"BE",X"B2",X"8D",X"56",X"34",X"19",X"12",X"1F",X"24",X"2B",X"38",X"3D",X"33",
		X"3B",X"4D",X"71",X"94",X"91",X"83",X"7B",X"7A",X"85",X"AE",X"D2",X"E4",X"E7",X"DA",X"D7",X"CF",
		X"BF",X"AA",X"B2",X"BD",X"AB",X"89",X"63",X"5B",X"66",X"79",X"7D",X"86",X"87",X"8A",X"89",X"86",
		X"76",X"51",X"30",X"29",X"3A",X"51",X"5C",X"6D",X"78",X"83",X"8B",X"91",X"95",X"97",X"98",X"98",
		X"97",X"94",X"91",X"8D",X"87",X"76",X"51",X"30",X"2A",X"3A",X"51",X"52",X"43",X"32",X"38",X"3C",
		X"40",X"48",X"68",X"9B",X"C0",X"DE",X"EF",X"E8",X"E0",X"DC",X"D6",X"D1",X"CC",X"C6",X"C1",X"BD",
		X"B4",X"96",X"5D",X"3E",X"40",X"42",X"38",X"1F",X"18",X"27",X"29",X"30",X"35",X"39",X"3D",X"40",
		X"4D",X"76",X"A5",X"A6",X"A7",X"BC",X"DE",X"F0",X"DE",X"DD",X"D7",X"D2",X"CD",X"C7",X"C3",X"BD",
		X"B9",X"B4",X"AF",X"A3",X"7D",X"4A",X"2C",X"12",X"09",X"15",X"23",X"34",X"36",X"26",X"2E",X"34",
		X"37",X"3D",X"49",X"71",X"9D",X"A5",X"9B",X"99",X"98",X"97",X"99",X"9A",X"9C",X"9F",X"A2",X"A4",
		X"AB",X"C3",X"DF",X"D6",X"CC",X"CC",X"C3",X"C1",X"BA",X"B7",X"B1",X"AE",X"A5",X"8A",X"5A",X"38",
		X"1E",X"0B",X"0B",X"17",X"1E",X"23",X"2A",X"2E",X"34",X"3B",X"58",X"8E",X"B7",X"D4",X"E6",X"DC",
		X"CC",X"B8",X"A4",X"95",X"8B",X"95",X"B1",X"BF",X"C2",X"BD",X"B7",X"B4",X"AF",X"AA",X"93",X"63",
		X"3A",X"21",X"0A",X"0C",X"17",X"1D",X"23",X"2A",X"2E",X"33",X"37",X"3D",X"51",X"85",X"BA",X"D9",
		X"ED",X"E1",X"D9",X"D4",X"C4",X"AE",X"9B",X"8C",X"7D",X"73",X"74",X"8D",X"A7",X"AA",X"97",X"7C",
		X"77",X"85",X"99",X"95",X"7F",X"61",X"51",X"40",X"36",X"2F",X"2B",X"2C",X"39",X"5E",X"87",X"98",
		X"92",X"82",X"7F",X"78",X"76",X"75",X"75",X"76",X"79",X"7C",X"81",X"90",X"B5",X"D8",X"DD",X"D3",
		X"CD",X"C9",X"C3",X"C0",X"BB",X"B5",X"A0",X"72",X"4A",X"31",X"1F",X"2D",X"3F",X"41",X"32",X"24",
		X"2E",X"39",X"51",X"6E",X"81",X"94",X"99",X"89",X"72",X"72",X"85",X"A0",X"A4",X"96",X"7E",X"74",
		X"69",X"65",X"6B",X"89",X"AB",X"B6",X"AC",X"98",X"99",X"AB",X"C6",X"CF",X"D1",X"C2",X"A7",X"8B",
		X"88",X"96",X"9B",X"8C",X"6C",X"56",X"58",X"69",X"78",X"7F",X"88",X"88",X"7B",X"5A",X"45",X"35",
		X"29",X"26",X"2A",X"31",X"34",X"39",X"3D",X"44",X"51",X"63",X"73",X"84",X"94",X"A6",X"C7",X"EF",
		X"F0",X"E0",X"E1",X"D8",X"D4",X"CE",X"CA",X"C5",X"C0",X"BB",X"B7",X"AE",X"97",X"74",X"5E",X"49",
		X"39",X"2D",X"27",X"34",X"54",X"6E",X"81",X"92",X"9D",X"A6",X"A9",X"AA",X"A8",X"A3",X"99",X"81",
		X"59",X"3E",X"38",X"45",X"51",X"57",X"61",X"67",X"6E",X"72",X"77",X"7A",X"7C",X"7B",X"6D",X"4F",
		X"3A",X"30",X"30",X"39",X"3E",X"54",X"79",X"96",X"AD",X"C0",X"BF",X"AA",X"98",X"8E",X"82",X"7D",
		X"78",X"77",X"77",X"7A",X"85",X"A5",X"CA",X"D8",X"D0",X"BB",X"B7",X"C3",X"CE",X"C3",X"BF",X"BB",
		X"B6",X"B3",X"AE",X"AB",X"A6",X"9B",X"85",X"70",X"5E",X"47",X"24",X"04",X"06",X"13",X"18",X"20",
		X"26",X"2B",X"30",X"35",X"3A",X"4A",X"73",X"9F",X"BB",X"D7",X"E4",X"E1",X"D7",X"D4",X"CD",X"C7",
		X"B8",X"9C",X"93",X"9B",X"93",X"90",X"88",X"7B",X"5D",X"3A",X"2B",X"30",X"41",X"4A",X"55",X"5E",
		X"61",X"53",X"3D",X"36",X"34",X"3B",X"40",X"51",X"75",X"90",X"8F",X"88",X"8E",X"A8",X"C9",X"D6",
		X"CE",X"B9",X"AE",X"A1",X"97",X"8F",X"87",X"83",X"86",X"9D",X"BB",X"C5",X"BA",X"A1",X"93",X"86",
		X"88",X"9D",X"AB",X"A4",X"8B",X"76",X"75",X"83",X"8E",X"84",X"6C",X"55",X"49",X"3B",X"35",X"30",
		X"30",X"34",X"47",X"6C",X"8E",X"A5",X"BB",X"C7",X"C3",X"A9",X"95",X"93",X"A0",X"AA",X"9F",X"85",
		X"6B",X"5D",X"4D",X"47",X"4D",X"68",X"7D",X"7E",X"6F",X"62",X"6A",X"82",X"98",X"A3",X"B0",X"B4",
		X"AB",X"8D",X"74",X"63",X"54",X"4A",X"42",X"3F",X"3E",X"3F",X"43",X"4C",X"62",X"8B",X"AD",X"B8",
		X"B0",X"A5",X"A2",X"9A",X"99",X"A1",X"BE",X"D0",X"D0",X"C8",X"C3",X"BF",X"BA",X"B6",X"B1",X"AE",
		X"A5",X"89",X"58",X"34",X"24",X"26",X"2B",X"22",X"19",X"1F",X"29",X"2A",X"32",X"35",X"3A",X"3D",
		X"41",X"46",X"5A",X"83",X"A8",X"C1",X"DA",X"E4",X"DB",X"C2",X"B9",X"BF",X"D1",X"D0",X"BE",X"A1",
		X"8C",X"7A",X"6A",X"64",X"70",X"87",X"8E",X"84",X"6E",X"63",X"59",X"52",X"54",X"68",X"87",X"9B",
		X"AC",X"B8",X"BB",X"AA",X"8D",X"7B",X"6B",X"5E",X"5A",X"68",X"81",X"8F",X"9C",X"A4",X"A5",X"94",
		X"77",X"66",X"57",X"4C",X"4A",X"5A",X"75",X"81",X"7D",X"6C",X"6A",X"78",X"91",X"A0",X"AD",X"B6",
		X"B5",X"A4",X"86",X"78",X"7A",X"89",X"8F",X"93",X"96",X"95",X"94",X"90",X"8B",X"85",X"80",X"79",
		X"72",X"6C",X"62",X"4C",X"2F",X"21",X"27",X"39",X"47",X"55",X"63",X"6B",X"65",X"54",X"4E",X"4B",
		X"4A",X"4E",X"53",X"5B",X"65",X"73",X"8B",X"B5",X"DA",X"E8",X"E2",X"D6",X"D2",X"C8",X"C3",X"C5",
		X"D4",X"D2",X"C7",X"C6",X"BF",X"BB",X"B5",X"B1",X"AD",X"A8",X"9F",X"8A",X"72",X"5F",X"45",X"21",
		X"06",X"08",X"15",X"1B",X"21",X"27",X"2C",X"31",X"35",X"3A",X"43",X"51",X"5D",X"75",X"9F",X"C4",
		X"D4",X"D0",X"C6",X"C3",X"BB",X"B7",X"BA",X"CE",X"D5",X"CA",X"C6",X"C1",X"BC",X"B8",X"B2",X"AB",
		X"91",X"66",X"4E",X"4D",X"4B",X"3F",X"28",X"15",X"18",X"21",X"27",X"2C",X"32",X"36",X"3B",X"44",
		X"61",X"8C",X"A9",X"C2",X"CD",X"C1",X"B4",X"AC",X"A1",X"9B",X"9E",X"B2",X"C5",X"CC",X"CE",X"C5",
		X"BF",X"AB",X"89",X"71",X"5D",X"4B",X"3F",X"36",X"31",X"2E",X"2F",X"32",X"38",X"3F",X"49",X"54",
		X"63",X"81",X"AA",X"C3",X"C9",X"BF",X"BC",X"C8",X"D8",X"D4",X"CA",X"C2",X"A9",X"94",X"83",X"77",
		X"7A",X"8A",X"91",X"95",X"97",X"92",X"80",X"62",X"4D",X"3C",X"2F",X"27",X"22",X"23",X"29",X"2F",
		X"33",X"39",X"42",X"50",X"5E",X"6C",X"7A",X"88",X"96",X"A2",X"AD",X"B7",X"BE",X"C5",X"C9",X"CB",
		X"CC",X"CA",X"C8",X"C5",X"C9",X"C8",X"BF",X"BD",X"B7",X"B2",X"AD",X"AC",X"A6",X"91",X"6E",X"53",
		X"3E",X"2A",X"1E",X"14",X"13",X"1A",X"26",X"3B",X"59",X"6C",X"80",X"8C",X"89",X"78",X"6E",X"68",
		X"62",X"60",X"5F",X"60",X"63",X"69",X"76",X"95",X"B5",X"C8",X"D9",X"DC",X"D4",X"C7",X"B2",X"99",
		X"89",X"78",X"6B",X"60",X"59",X"5C",X"70",X"85",X"8A",X"7F",X"6F",X"69",X"61",X"5E",X"64",X"7B",
		X"92",X"99",X"90",X"81",X"83",X"92",X"A5",X"A5",X"97",X"82",X"7F",X"89",X"97",X"94",X"85",X"6F",
		X"65",X"58",X"52",X"55",X"69",X"80",X"86",X"7E",X"6F",X"6A",X"64",X"62",X"68",X"81",X"9A",X"A2",
		X"99",X"8B",X"8C",X"9B",X"AD",X"AD",X"9E",X"8A",X"86",X"8E",X"9C",X"9F",X"A4",X"A2",X"9A",X"80",
		X"65",X"54",X"44",X"3A",X"33",X"2F",X"2E",X"30",X"35",X"3D",X"4D",X"6F",X"93",X"AC",X"C3",X"D3",
		X"D7",X"C8",X"B3",X"A5",X"96",X"8A",X"7F",X"79",X"80",X"94",X"A2",X"AA",X"B1",X"B2",X"B1",X"AC",
		X"A5",X"9C",X"93",X"86",X"6F",X"4E",X"35",X"24",X"17",X"18",X"21",X"2E",X"41",X"49",X"41",X"41",
		X"44",X"49",X"51",X"5A",X"65",X"71",X"7D",X"89",X"98",X"B2",X"D8",X"EE",X"EB",X"E1",X"DE",X"D8",
		X"D2",X"CD",X"C8",X"C3",X"BD",X"B8",X"AD",X"92",X"7A",X"7A",X"72",X"6B",X"64",X"5B",X"49",X"2E",
		X"1C",X"17",X"1F",X"27",X"2B",X"33",X"42",X"5D",X"74",X"87",X"99",X"A7",X"B3",X"BB",X"C0",X"C0",
		X"B4",X"9A",X"89",X"86",X"8F",X"95",X"96",X"99",X"98",X"97",X"94",X"8F",X"7F",X"64",X"51",X"43",
		X"38",X"33",X"30",X"32",X"36",X"3D",X"46",X"51",X"5D",X"70",X"93",X"B9",X"D3",X"E7",X"E8",X"DE",
		X"DA",X"D5",X"CF",X"CA",X"C2",X"AE",X"8E",X"76",X"63",X"52",X"46",X"3D",X"38",X"35",X"35",X"38",
		X"3E",X"4B",X"68",X"8A",X"9C",X"9D",X"96",X"9B",X"AC",X"C3",X"CD",X"D2",X"CD",X"C6",X"C3",X"BD",
		X"B9",X"B4",X"AA",X"95",X"73",X"51",X"3E",X"3A",X"3E",X"3F",X"42",X"45",X"44",X"38",X"2A",X"29",
		X"2F",X"35",X"39",X"45",X"60",X"80",X"95",X"AC",X"BB",X"C9",X"D1",X"D1",X"C1",X"AA",X"9B",X"8C",
		X"81",X"7C",X"87",X"97",X"99",X"8F",X"7D",X"79",X"81",X"91",X"98",X"9E",X"A1",X"A2",X"A1",X"9D",
		X"94",X"7E",X"64",X"58",X"5A",X"64",X"68",X"6D",X"71",X"74",X"75",X"6C",X"59",X"4B",X"43",X"3D",
		X"3C",X"3D",X"41",X"49",X"5C",X"7D",X"98",X"A3",X"9F",X"9D",X"AA",X"BF",X"D1",X"D7",X"D6",X"CD",
		X"C9",X"BC",X"A6",X"98",X"9C",X"9A",X"96",X"91",X"8A",X"83",X"7B",X"73",X"62",X"47",X"33",X"2F",
		X"39",X"42",X"41",X"37",X"31",X"3A",X"4E",X"63",X"69",X"65",X"63",X"71",X"89",X"A1",X"B0",X"BF",
		X"C6",X"C3",X"AF",X"A0",X"9E",X"A7",X"AF",X"B0",X"B2",X"AE",X"AB",X"A4",X"9C",X"8B",X"6F",X"58",
		X"51",X"56",X"5D",X"5F",X"64",X"66",X"61",X"51",X"45",X"3F",X"3B",X"3D",X"48",X"63",X"7B",X"8E",
		X"A0",X"AC",X"AE",X"A0",X"95",X"8E",X"87",X"84",X"8A",X"9E",X"AD",X"B6",X"BE",X"C0",X"C0",X"B8",
		X"A4",X"88",X"79",X"77",X"7D",X"79",X"6A",X"57",X"4B",X"42",X"3B",X"38",X"38",X"3B",X"44",X"5A",
		X"78",X"8E",X"A1",X"B0",X"BC",X"C3",X"C7",X"C8",X"C6",X"C0",X"B6",X"9F",X"81",X"70",X"6B",X"6F",
		X"6A",X"5C",X"48",X"3D",X"35",X"31",X"34",X"44",X"5D",X"6C",X"6F",X"6A",X"6C",X"6D",X"70",X"78",
		X"8D",X"A8",X"B5",X"B4",X"A9",X"A3",X"9D",X"98",X"94",X"91",X"8E",X"8C",X"8A",X"89",X"8B",X"99",
		X"AE",X"B8",X"C0",X"C2",X"BE",X"B9",X"B4",X"AE",X"A4",X"97",X"89",X"7B",X"6E",X"61",X"56",X"4C",
		X"40",X"2E",X"18",X"12",X"1A",X"23",X"2C",X"3A",X"47",X"52",X"52",X"4C",X"4D",X"50",X"5D",X"78",
		X"90",X"9B",X"9A",X"97",X"9A",X"9A",X"9D",X"A7",X"BE",X"D0",X"D3",X"C8",X"BA",X"B9",X"C1",X"C8",
		X"BF",X"AB",X"95",X"8E",X"90",X"94",X"89",X"76",X"63",X"5F",X"65",X"6D",X"67",X"5A",X"4D",X"4F",
		X"5B",X"69",X"6A",X"63",X"59",X"57",X"54",X"56",X"58",X"5C",X"62",X"71",X"8C",X"A5",X"B6",X"C5",
		X"CE",X"D2",X"CF",X"C8",X"C1",X"AE",X"92",X"7E",X"6D",X"5E",X"53",X"4B",X"46",X"4A",X"5B",X"6B",
		X"70",X"6A",X"62",X"62",X"60",X"62",X"6B",X"81",X"95",X"9C",X"97",X"8E",X"8B",X"85",X"83",X"80",
		X"7F",X"7F",X"87",X"9A",X"AD",X"B6",X"BF",X"C1",X"BA",X"A5",X"8F",X"7F",X"6F",X"63",X"59",X"55",
		X"5C",X"6B",X"73",X"70",X"64",X"5E",X"5A",X"57",X"57",X"58",X"5A",X"5E",X"63",X"69",X"73",X"87",
		X"A2",X"B5",X"C3",X"CD",X"CF",X"C4",X"AF",X"9E",X"8F",X"81",X"78",X"7A",X"84",X"88",X"8B",X"8D",
		X"8C",X"8A",X"86",X"7F",X"6F",X"59",X"4C",X"4C",X"55",X"59",X"53",X"47",X"44",X"4D",X"5F",X"6D",
		X"79",X"85",X"8E",X"96",X"9B",X"9F",X"A2",X"A2",X"9F",X"92",X"7E",X"73",X"73",X"7D",X"82",X"85",
		X"89",X"87",X"7E",X"6C",X"62",X"5B",X"56",X"54",X"54",X"56",X"5C",X"6E",X"88",X"99",X"9E",X"98",
		X"98",X"A2",X"B4",X"BF",X"C6",X"CB",X"C8",X"BA",X"A2",X"90",X"80",X"72",X"67",X"5E",X"58",X"53",
		X"50",X"4F",X"50",X"53",X"58",X"5D",X"64",X"71",X"8A",X"A2",X"B2",X"C1",X"C8",X"C7",X"B7",X"A5",
		X"9D",X"9F",X"A3",X"A0",X"9E",X"98",X"92",X"8A",X"81",X"79",X"70",X"68",X"5C",X"47",X"33",X"28",
		X"1F",X"1F",X"26",X"32",X"44",X"52",X"52",X"53",X"59",X"5F",X"67",X"6F",X"78",X"82",X"8C",X"95",
		X"9F",X"AD",X"C6",X"DD",X"E3",X"DD",X"D2",X"C8",X"BC",X"B3",X"AD",X"B3",X"B9",X"B7",X"B5",X"AE",
		X"A6",X"9C",X"91",X"85",X"78",X"6C",X"61",X"57",X"4D",X"41",X"2E",X"1D",X"16",X"1A",X"23",X"28",
		X"2E",X"38",X"4C",X"62",X"73",X"80",X"80",X"7D",X"80",X"81",X"85",X"89",X"8E",X"92",X"9C",X"B1",
		X"C6",X"D1",X"DA",X"D8",X"D0",X"CC",X"C7",X"C1",X"BB",X"AC",X"8E",X"72",X"5F",X"4C",X"3F",X"34",
		X"2E",X"2A",X"2A",X"2D",X"32",X"38",X"41",X"4D",X"63",X"82",X"9B",X"AF",X"C0",X"CB",X"CA",X"BB",
		X"B1",X"A7",X"9D",X"97",X"99",X"A4",X"A7",X"A0",X"8F",X"83",X"82",X"89",X"8B",X"82",X"72",X"65",
		X"5D",X"55",X"52",X"4F",X"4F",X"51",X"5E",X"73",X"82",X"85",X"80",X"7C",X"7C",X"7A",X"7B",X"7C",
		X"7E",X"7F",X"82",X"84",X"88",X"95",X"A9",X"B6",X"B5",X"A9",X"A1",X"A2",X"AA",X"AF",X"AE",X"AC",
		X"A5",X"96",X"7E",X"6C",X"65",X"67",X"68",X"66",X"66",X"64",X"64",X"63",X"61",X"59",X"49",X"3F",
		X"3A",X"36",X"36",X"39",X"43",X"57",X"70",X"83",X"95",X"A3",X"AB",X"A6",X"9D",X"98",X"93",X"8F",
		X"8C",X"8A",X"88",X"8C",X"9A",X"AB",X"B4",X"BB",X"BD",X"BD",X"BB",X"B5",X"AA",X"95",X"7D",X"70",
		X"6D",X"6F",X"68",X"5B",X"4C",X"48",X"4E",X"59",X"5C",X"57",X"4F",X"52",X"5E",X"6F",X"77",X"76",
		X"6F",X"6F",X"6F",X"72",X"78",X"89",X"9D",X"AA",X"B6",X"BD",X"BD",X"B1",X"A0",X"95",X"89",X"80",
		X"79",X"72",X"6E",X"6E",X"79",X"87",X"8B",X"86",X"7B",X"7A",X"82",X"8E",X"93",X"98",X"99",X"96",
		X"88",X"77",X"6D",X"63",X"5C",X"57",X"55",X"54",X"55",X"57",X"5B",X"64",X"77",X"8D",X"9C",X"A9",
		X"B2",X"B4",X"AA",X"9B",X"91",X"87",X"7E",X"77",X"73",X"77",X"84",X"8D",X"8B",X"80",X"79",X"7B",
		X"85",X"8C",X"88",X"7D",X"72",X"6D",X"66",X"63",X"61",X"61",X"61",X"63",X"66",X"69",X"6D",X"71",
		X"78",X"85",X"9B",X"AC",X"AF",X"A7",X"A0",X"9B",X"94",X"90",X"8A",X"86",X"81",X"7E",X"7B",X"79",
		X"78",X"77",X"77",X"7F",X"8F",X"9A",X"99",X"8F",X"84",X"7E",X"77",X"74",X"76",X"83",X"8B",X"89",
		X"7E",X"74",X"6E",X"68",X"65",X"62",X"61",X"60",X"61",X"63",X"67",X"72",X"86",X"96",X"9A",X"93",
		X"8C",X"89",X"84",X"83",X"87",X"96",X"9E",X"9C",X"91",X"87",X"88",X"90",X"96",X"90",X"83",X"76",
		X"6E",X"65",X"60",X"62",X"70",X"7A",X"81",X"87",X"8B",X"8E",X"8F",X"8F",X"8E",X"89",X"7B",X"6A",
		X"62",X"64",X"6C",X"70",X"74",X"78",X"7A",X"7D",X"7E",X"80",X"81",X"81",X"7E",X"74",X"66",X"5E",
		X"58",X"55",X"57",X"64",X"76",X"83",X"8F",X"98",X"9E",X"99",X"8E",X"89",X"84",X"81",X"81",X"8B",
		X"9A",X"A3",X"AA",X"AF",X"B1",X"B0",X"AD",X"A9",X"A3",X"9D",X"95",X"8D",X"85",X"7A",X"69",X"55",
		X"4B",X"4A",X"50",X"51",X"4C",X"44",X"41",X"41",X"42",X"47",X"4D",X"56",X"62",X"78",X"92",X"A6",
		X"B6",X"C3",X"C9",X"C4",X"B7",X"B2",X"B4",X"BA",X"BA",X"B9",X"B5",X"AF",X"A7",X"9E",X"94",X"8A",
		X"80",X"76",X"6C",X"63",X"5A",X"4B",X"3A",X"30",X"29",X"25",X"26",X"2C",X"31",X"36",X"3E",X"4A",
		X"57",X"65",X"7A",X"96",X"B1",X"C4",X"D5",X"DF",X"E0",X"D5",X"C9",X"BD",X"B1",X"A6",X"9B",X"91",
		X"87",X"7F",X"78",X"72",X"6E",X"6A",X"68",X"67",X"67",X"69",X"71",X"81",X"8F",X"97",X"9F",X"A3",
		X"A5",X"A5",X"A2",X"9E",X"99",X"92",X"8B",X"83",X"7B",X"73",X"6C",X"66",X"60",X"5B",X"57",X"54",
		X"52",X"51",X"52",X"53",X"55",X"54",X"4D",X"47",X"47",X"47",X"4C",X"56",X"6B",X"7F",X"90",X"A0",
		X"AC",X"B6",X"BD",X"C1",X"BE",X"B1",X"A3",X"9A",X"8F",X"89",X"87",X"8F",X"95",X"93",X"89",X"7E",
		X"78",X"71",X"6E",X"71",X"7D",X"88",X"8F",X"95",X"99",X"9A",X"98",X"8E",X"7E",X"76",X"76",X"7C",
		X"7F",X"80",X"81",X"7F",X"77",X"69",X"61",X"5B",X"57",X"56",X"56",X"58",X"5D",X"6B",X"7E",X"8A",
		X"8D",X"89",X"8A",X"93",X"A1",X"AA",X"B0",X"B4",X"B2",X"A9",X"98",X"8E",X"8B",X"8E",X"8E",X"8C",
		X"8A",X"86",X"83",X"7E",X"79",X"75",X"71",X"6D",X"6A",X"68",X"64",X"5B",X"4E",X"49",X"4C",X"56",
		X"5C",X"5C",X"58",X"57",X"59",X"5C",X"64",X"73",X"88",X"96",X"9B",X"98",X"9A",X"A4",X"B2",X"BA",
		X"C0",X"C3",X"C0",X"B6",X"A4",X"96",X"89",X"7E",X"76",X"76",X"7D",X"80",X"81",X"82",X"80",X"78",
		X"6A",X"63",X"65",X"6D",X"72",X"76",X"7A",X"7A",X"75",X"6A",X"64",X"60",X"5D",X"5C",X"5D",X"60",
		X"63",X"68",X"6E",X"74",X"7B",X"85",X"98",X"AA",X"B1",X"AE",X"A7",X"A9",X"B0",X"B7",X"B4",X"A8",
		X"9A",X"94",X"95",X"97",X"90",X"82",X"72",X"69",X"5F",X"59",X"58",X"60",X"69",X"6F",X"75",X"79",
		X"79",X"71",X"69",X"65",X"61",X"60",X"63",X"70",X"7D",X"82",X"80",X"7B",X"7F",X"89",X"94",X"96",
		X"91",X"88",X"85",X"7F",X"7D",X"7F",X"89",X"94",X"99",X"9E",X"A0",X"A1",X"A0",X"9D",X"99",X"94",
		X"8E",X"84",X"74",X"64",X"5A",X"50",X"4B",X"4B",X"54",X"5F",X"66",X"6F",X"76",X"79",X"74",X"6F",
		X"72",X"7C",X"87",X"8A",X"87",X"81",X"83",X"8C",X"97",X"98",X"93",X"8A",X"86",X"81",X"7D",X"7B",
		X"7A",X"79",X"79",X"7A",X"7C",X"7D",X"81",X"8A",X"9A",X"A4",X"AB",X"B0",X"B2",X"B2",X"AF",X"AA",
		X"A4",X"9D",X"95",X"8C",X"83",X"79",X"70",X"68",X"60",X"5A",X"55",X"50",X"48",X"3C",X"36",X"34",
		X"33",X"37",X"42",X"55",X"64",X"6C",X"6F",X"75",X"82",X"94",X"A3",X"AE",X"B8",X"BD",X"BA",X"AF",
		X"A8",X"A7",X"AC",X"AC",X"A4",X"95",X"8A",X"87",X"8A",X"8A",X"82",X"76",X"6D",X"6D",X"72",X"76",
		X"72",X"69",X"64",X"68",X"71",X"77",X"76",X"6F",X"6C",X"71",X"7C",X"83",X"83",X"7D",X"7A",X"79",
		X"77",X"79",X"80",X"8D",X"96",X"9C",X"A1",X"A3",X"A5",X"A4",X"A2",X"9E",X"9A",X"94",X"8F",X"88",
		X"81",X"7B",X"75",X"70",X"6B",X"63",X"57",X"4B",X"47",X"4B",X"53",X"56",X"54",X"51",X"56",X"61",
		X"70",X"78",X"7B",X"7A",X"7D",X"7F",X"83",X"86",X"8A",X"8D",X"91",X"95",X"98",X"9B",X"9D",X"9F",
		X"A0",X"A1",X"A2",X"A2",X"A1",X"9F",X"A0",X"A8",X"B0",X"B1",X"B2",X"AE",X"A9",X"A2",X"9A",X"91",
		X"88",X"7E",X"75",X"6C",X"63",X"59",X"4A",X"3C",X"36",X"37",X"3D",X"3F",X"3E",X"3B",X"40",X"4C",
		X"5B",X"66",X"6A",X"6B",X"70",X"75",X"7B",X"83",X"93",X"A5",X"AD",X"AD",X"A8",X"AA",X"B0",X"B9",
		X"B9",X"B1",X"A5",X"9C",X"93",X"8B",X"86",X"89",X"8E",X"8E",X"8F",X"8D",X"88",X"7D",X"6F",X"67",
		X"60",X"60",X"67",X"6D",X"71",X"75",X"77",X"75",X"6C",X"67",X"69",X"72",X"79",X"7E",X"83",X"87",
		X"8A",X"8C",X"8C",X"88",X"7D",X"76",X"71",X"6D",X"6B",X"6F",X"7A",X"82",X"83",X"7E",X"7B",X"80",
		X"89",X"91",X"95",X"9A",X"9B",X"98",X"8C",X"84",X"83",X"87",X"8A",X"8A",X"8B",X"8A",X"84",X"78",
		X"70",X"6E",X"73",X"77",X"79",X"7C",X"7C",X"78",X"6F",X"69",X"69",X"71",X"78",X"7C",X"81",X"83",
		X"82",X"7A",X"75",X"72",X"6F",X"6E",X"6E",X"6F",X"72",X"7A",X"88",X"92",X"95",X"92",X"8F",X"8E",
		X"8B",X"8B",X"8F",X"99",X"A1",X"A5",X"A7",X"A7",X"A5",X"A2",X"9D",X"97",X"91",X"8A",X"82",X"7B",
		X"74",X"6E",X"68",X"63",X"5F",X"5A",X"51",X"47",X"42",X"3F",X"3F",X"43",X"4E",X"5E",X"68",X"6D",
		X"6F",X"74",X"79",X"7E",X"84",X"89",X"8F",X"94",X"99",X"9D",X"A3",X"AF",X"BC",X"C3",X"C8",X"C8",
		X"C4",X"B8",X"A7",X"99",X"8C",X"80",X"78",X"77",X"79",X"76",X"6E",X"63",X"5D",X"57",X"53",X"53",
		X"5A",X"65",X"6D",X"74",X"7B",X"7F",X"7C",X"76",X"74",X"71",X"70",X"6F",X"70",X"71",X"73",X"77",
		X"7A",X"80",X"8B",X"99",X"A0",X"9F",X"99",X"96",X"92",X"8E",X"8A",X"87",X"85",X"84",X"8A",X"93",
		X"95",X"90",X"87",X"82",X"7C",X"77",X"73",X"70",X"6E",X"6F",X"76",X"80",X"86",X"8B",X"8F",X"8F",
		X"88",X"7E",X"77",X"72",X"71",X"77",X"7C",X"7F",X"82",X"84",X"85",X"85",X"84",X"83",X"81",X"7F",
		X"79",X"6F",X"67",X"65",X"69",X"6E",X"6D",X"68",X"65",X"68",X"71",X"7A",X"80",X"87",X"8B",X"8B",
		X"85",X"80",X"7D",X"7B",X"7A",X"79",X"7A",X"7B",X"81",X"8D",X"97",X"9D",X"A3",X"A6",X"A8",X"A7",
		X"A6",X"A2",X"9E",X"98",X"8F",X"7F",X"72",X"68",X"5F",X"59",X"55",X"52",X"51",X"52",X"54",X"58",
		X"5D",X"63",X"69",X"6F",X"76",X"7E",X"89",X"99",X"A7",X"AD",X"AB",X"A7",X"A9",X"AF",X"B4",X"B3",
		X"B3",X"AE",X"A5",X"95",X"86",X"7E",X"7B",X"78",X"71",X"66",X"5B",X"55",X"50",X"4D",X"4C",X"4E",
		X"50",X"57",X"64",X"71",X"7B",X"83",X"84",X"82",X"81",X"82",X"82",X"84",X"85",X"86",X"87",X"88",
		X"8A",X"8C",X"94",X"9F",X"A4",X"A1",X"9A",X"94",X"8E",X"89",X"86",X"88",X"8E",X"8F",X"89",X"7F",
		X"79",X"73",X"6E",X"6C",X"6F",X"77",X"7A",X"78",X"72",X"6F",X"6D",X"6B",X"6B",X"6B",X"6D",X"6E",
		X"70",X"72",X"77",X"81",X"8E",X"97",X"9E",X"A3",X"A4",X"9F",X"94",X"8C",X"85",X"7F",X"7A",X"75",
		X"72",X"71",X"76",X"7E",X"82",X"80",X"7A",X"76",X"73",X"71",X"70",X"6F",X"6F",X"71",X"79",X"85",
		X"8D",X"93",X"98",X"9A",X"95",X"8B",X"86",X"85",X"89",X"88",X"83",X"7A",X"75",X"76",X"7B",X"7E",
		X"80",X"82",X"81",X"7B",X"72",X"6D",X"68",X"65",X"63",X"63",X"68",X"72",X"7D",X"84",X"8C",X"91",
		X"95",X"98",X"99",X"96",X"8D",X"84",X"82",X"84",X"88",X"88",X"89",X"88",X"87",X"86",X"84",X"82",
		X"80",X"7E",X"7C",X"7A",X"78",X"74",X"6B",X"64",X"63",X"67",X"6D",X"6F",X"6C",X"69",X"6C",X"74",
		X"7E",X"81",X"80",X"7D",X"81",X"89",X"93",X"98",X"9D",X"9F",X"9E",X"97",X"8F",X"89",X"83",X"7E",
		X"7D",X"83",X"88",X"88",X"83",X"7D",X"7C",X"80",X"86",X"88",X"8A",X"8A",X"8B",X"8A",X"88",X"84",
		X"7A",X"71",X"6E",X"70",X"74",X"73",X"6E",X"69",X"69",X"6F",X"76",X"78",X"77",X"73",X"73",X"73",
		X"74",X"75",X"77",X"79",X"7C",X"7F",X"82",X"85",X"87",X"8A",X"8C",X"8F",X"97",X"A2",X"A8",X"A6",
		X"9F",X"99",X"94",X"8E",X"8B",X"8B",X"8F",X"8F",X"89",X"80",X"78",X"72",X"6D",X"6A",X"6C",X"73",
		X"77",X"7A",X"7D",X"7E",X"7F",X"7F",X"7F",X"7E",X"7D",X"7B",X"75",X"6C",X"66",X"62",X"5F",X"5F",
		X"64",X"6E",X"76",X"7D",X"83",X"88",X"8D",X"90",X"91",X"8D",X"86",X"80",X"7C",X"78",X"75",X"74",
		X"74",X"75",X"7B",X"85",X"8C",X"92",X"97",X"9A",X"9C",X"9C",X"9A",X"93",X"88",X"7F",X"78",X"72",
		X"6E",X"6B",X"69",X"67",X"68",X"69",X"6B",X"6D",X"70",X"74",X"7D",X"89",X"92",X"94",X"91",X"8F",
		X"8E",X"8C",X"8C",X"8F",X"97",X"9B",X"9D",X"9E",X"9D",X"9A",X"94",X"89",X"7D",X"75",X"6D",X"67",
		X"62",X"5F",X"5D",X"5F",X"66",X"6F",X"73",X"73",X"71",X"73",X"7B",X"84",X"89",X"8F",X"92",X"92",
		X"8C",X"85",X"83",X"85",X"89",X"88",X"82",X"7B",X"7A",X"7D",X"82",X"83",X"85",X"86",X"87",X"87",
		X"86",X"85",X"84",X"82",X"7E",X"76",X"6D",X"68",X"64",X"63",X"62",X"62",X"63",X"68",X"72",X"7D",
		X"85",X"8E",X"94",X"97",X"94",X"8F",X"8F",X"92",X"97",X"97",X"92",X"8A",X"85",X"80",X"7C",X"79",
		X"77",X"76",X"75",X"75",X"75",X"76",X"77",X"79",X"7B",X"7D",X"7F",X"84",X"8D",X"96",X"9B",X"A0",
		X"A2",X"A3",X"A2",X"9F",X"9B",X"96",X"90",X"88",X"7C",X"6F",X"66",X"5F",X"5C",X"5E",X"61",X"63",
		X"66",X"67",X"67",X"62",X"60",X"61",X"61",X"64",X"66",X"6A",X"6E",X"73",X"78",X"7F",X"88",X"95",
		X"9F",X"A2",X"A0",X"9E",X"9D",X"9A",X"98",X"95",X"93",X"90",X"8E",X"8B",X"8A",X"8B",X"91",X"94",
		X"95",X"95",X"93",X"90",X"8D",X"89",X"84",X"80",X"7B",X"77",X"72",X"6E",X"6A",X"67",X"64",X"5F",
		X"58",X"52",X"50",X"4F",X"51",X"57",X"62",X"6D",X"76",X"80",X"88",X"8E",X"94",X"97",X"97",X"92",
		X"8F",X"90",X"94",X"98",X"99",X"9A",X"99",X"98",X"95",X"92",X"8E",X"8A",X"85",X"7E",X"74",X"6B",
		X"66",X"61",X"5F",X"5E",X"5E",X"5F",X"62",X"65",X"6A",X"6E",X"73",X"78",X"7E",X"85",X"90",X"9D",
		X"A5",X"AC",X"B1",X"B1",X"AB",X"A1",X"9A",X"93",X"8C",X"87",X"87",X"88",X"85",X"7F",X"76",X"70",
		X"6B",X"68",X"66",X"64",X"64",X"66",X"6D",X"76",X"7B",X"7B",X"79",X"7A",X"80",X"87",X"8B",X"8F",
		X"91",X"91",X"8B",X"84",X"80",X"82",X"85",X"84",X"7F",X"78",X"76",X"78",X"7C",X"7E",X"80",X"81",
		X"82",X"82",X"82",X"80",X"7B",X"74",X"70",X"6C",X"6A",X"6B",X"70",X"78",X"7B",X"7B",X"79",X"7A",
		X"7F",X"87",X"8A",X"89",X"86",X"84",X"83",X"81",X"81",X"80",X"80",X"80",X"81",X"81",X"82",X"83",
		X"84",X"86",X"8D",X"95",X"98",X"95",X"8F",X"8C",X"8E",X"91",X"90",X"8B",X"82",X"7C",X"76",X"75",
		X"79",X"7B",X"79",X"74",X"70",X"70",X"74",X"79",X"7B",X"7D",X"7E",X"7D",X"77",X"72",X"70",X"6E",
		X"6D",X"6C",X"6D",X"6E",X"70",X"72",X"75",X"7C",X"86",X"8E",X"91",X"90",X"8E",X"8D",X"8C",X"8C",
		X"8A",X"89",X"88",X"87",X"85",X"84",X"84",X"83",X"82",X"81",X"81",X"80",X"83",X"8A",X"8F",X"8E",
		X"89",X"84",X"84",X"87",X"8A",X"87",X"80",X"79",X"78",X"7A",X"7C",X"7A",X"75",X"70",X"6D",X"6A",
		X"69",X"6C",X"73",X"7A",X"7B",X"79",X"77",X"7A",X"80",X"85",X"89",X"8C",X"8E",X"8D",X"86",X"81",
		X"80",X"83",X"86",X"84",X"7E",X"79",X"79",X"7D",X"81",X"83",X"85",X"85",X"84",X"7D",X"78",X"74",
		X"71",X"6F",X"6E",X"6F",X"70",X"71",X"73",X"76",X"78",X"7D",X"85",X"8F",X"95",X"9A",X"9E",X"9F",
		X"9B",X"93",X"8E",X"88",X"83",X"80",X"81",X"85",X"86",X"87",X"87",X"85",X"80",X"78",X"74",X"73",
		X"76",X"76",X"73",X"6E",X"6B",X"69",X"68",X"6A",X"70",X"78",X"7E",X"84",X"88",X"8B",X"89",X"84",
		X"82",X"7F",X"7D",X"7C",X"7C",X"7C",X"7E",X"83",X"8A",X"8E",X"91",X"94",X"95",X"96",X"95",X"93",
		X"91",X"8E",X"89",X"81",X"78",X"72",X"70",X"71",X"70",X"6D",X"67",X"65",X"63",X"63",X"65",X"6B",
		X"74",X"7B",X"82",X"87",X"8C",X"8F",X"92",X"93",X"8F",X"89",X"86",X"86",X"89",X"8A",X"86",X"80",
		X"7C",X"79",X"78",X"7C",X"80",X"83",X"86",X"87",X"87",X"81",X"7C",X"79",X"76",X"74",X"75",X"7A",
		X"80",X"81",X"7F",X"7C",X"7B",X"7A",X"79",X"79",X"7A",X"7B",X"7E",X"86",X"8C",X"90",X"94",X"96",
		X"94",X"8E",X"88",X"86",X"87",X"89",X"88",X"88",X"87",X"83",X"7B",X"74",X"71",X"72",X"74",X"74",
		X"76",X"77",X"78",X"79",X"7A",X"79",X"74",X"70",X"70",X"73",X"78",X"7B",X"7F",X"82",X"84",X"85",
		X"86",X"85",X"80",X"7C",X"7A",X"77",X"77",X"78",X"7E",X"84",X"88",X"8B",X"8D",X"8C",X"88",X"83",
		X"82",X"84",X"87",X"87",X"83",X"7E",X"7C",X"79",X"78",X"77",X"77",X"77",X"78",X"79",X"7A",X"7C",
		X"7D",X"7E",X"80",X"83",X"88",X"90",X"95",X"99",X"9C",X"9B",X"97",X"90",X"8A",X"88",X"89",X"88",
		X"86",X"84",X"80",X"7A",X"72",X"6C",X"6B",X"6C",X"6C",X"6A",X"66",X"64",X"64",X"64",X"65",X"67",
		X"6A",X"6D",X"70",X"74",X"78",X"7C",X"80",X"84",X"88",X"8B",X"8F",X"91",X"94",X"96",X"97",X"97",
		X"97",X"97",X"95",X"94",X"92",X"90",X"8F",X"91",X"94",X"95",X"95",X"93",X"90",X"88",X"7E",X"77",
		X"73",X"73",X"71",X"70",X"6F",X"6E",X"6E",X"6D",X"6D",X"6A",X"64",X"61",X"60",X"5F",X"61",X"66",
		X"6F",X"76",X"7C",X"82",X"88",X"8C",X"8F",X"91",X"8F",X"8A",X"86",X"84",X"82",X"81",X"83",X"88",
		X"8B",X"8E",X"8F",X"90",X"90",X"8E",X"8D",X"8A",X"86",X"7F",X"78",X"75",X"76",X"78",X"77",X"73",
		X"6F",X"6F",X"72",X"77",X"79",X"78",X"75",X"77",X"7B",X"81",X"83",X"82",X"7F",X"7F",X"7E",X"7F",
		X"80",X"86",X"8B",X"8F",X"92",X"94",X"94",X"8F",X"89",X"87",X"88",X"89",X"87",X"82",X"7C",X"7A",
		X"7B",X"7D",X"7C",X"78",X"73",X"73",X"75",X"79",X"7A",X"77",X"74",X"73",X"72",X"73",X"73",X"74",
		X"76",X"78",X"7B",X"7D",X"80",X"82",X"85",X"87",X"89",X"8B",X"8E",X"94",X"9A",X"9B",X"98",X"93",
		X"90",X"8B",X"88",X"86",X"87",X"89",X"89",X"88",X"86",X"84",X"82",X"7F",X"7C",X"7A",X"77",X"74",
		X"6E",X"67",X"63",X"60",X"5E",X"5E",X"5F",X"63",X"6B",X"71",X"75",X"75",X"77",X"7D",X"85",X"8B",
		X"8D",X"8B",X"8A",X"8A",X"89",X"8A",X"8C",X"92",X"95",X"94",X"90",X"8C",X"8C",X"8D",X"8F",X"8E",
		X"8E",X"8B",X"86",X"7E",X"79",X"77",X"78",X"78",X"78",X"78",X"78",X"75",X"70",X"6D",X"6B",X"6A",
		X"6A",X"6D",X"74",X"7A",X"7F",X"84",X"87",X"8A",X"8B",X"8D",X"8E",X"8E",X"8D",X"8A",X"83",X"7F",
		X"7B",X"78",X"76",X"77",X"7C",X"7F",X"81",X"84",X"85",X"83",X"7F",X"7B",X"79",X"78",X"78",X"7A",
		X"7F",X"83",X"84",X"81",X"80",X"82",X"86",X"89",X"8B",X"8C",X"8D",X"8D",X"8C",X"8B",X"8A",X"88",
		X"85",X"81",X"79",X"74",X"6F",X"6C",X"6A",X"68",X"68",X"68",X"69",X"6B",X"6E",X"71",X"75",X"79",
		X"7D",X"80",X"84",X"87",X"8A",X"8D",X"8F",X"92",X"98",X"9F",X"A1",X"A3",X"A3",X"A0",X"99",X"91",
		X"8A",X"83",X"7E",X"79",X"78",X"79",X"78",X"77",X"77",X"75",X"70",X"6B",X"69",X"6A",X"6E",X"70",
		X"73",X"75",X"76",X"75",X"72",X"72",X"76",X"7B",X"7E",X"7D",X"7B",X"7C",X"80",X"86",X"89",X"8C",
		X"8E",X"8D",X"8A",X"85",X"83",X"85",X"87",X"87",X"83",X"7F",X"7C",X"7A",X"78",X"77",X"77",X"77",
		X"77",X"78",X"79",X"7C",X"81",X"88",X"8C",X"8F",X"91",X"93",X"93",X"93",X"91",X"8B",X"84",X"80",
		X"7F",X"7F",X"7E",X"7A",X"75",X"73",X"74",X"76",X"78",X"79",X"78",X"74",X"72",X"71",X"71",X"71",
		X"72",X"73",X"75",X"7A",X"81",X"88",X"8C",X"91",X"93",X"95",X"95",X"94",X"91",X"8B",X"85",X"81",
		X"7D",X"7A",X"79",X"7C",X"7E",X"7F",X"80",X"80",X"7E",X"7A",X"77",X"77",X"79",X"7C",X"7E",X"80",
		X"81",X"82",X"82",X"82",X"80",X"7C",X"78",X"76",X"74",X"73",X"73",X"73",X"75",X"78",X"7F",X"84",
		X"88",X"8C",X"8E",X"8D",X"8A",X"87",X"87",X"89",X"8B",X"8C",X"8D",X"8C",X"89",X"83",X"7E",X"7C",
		X"7C",X"7C",X"7A",X"76",X"73",X"71",X"6F",X"6F",X"70",X"71",X"72",X"74",X"76",X"78",X"7A",X"7D",
		X"80",X"85",X"8C",X"92",X"96",X"99",X"9A",X"99",X"93",X"8E",X"8A",X"85",X"81",X"7D",X"7A",X"77",
		X"75",X"73",X"72",X"72",X"72",X"73",X"74",X"75",X"76",X"78",X"7A",X"80",X"87",X"8B",X"8F",X"90",
		X"90",X"8D",X"87",X"84",X"84",X"85",X"85",X"81",X"7C",X"79",X"79",X"7B",X"7C",X"7C",X"7D",X"7C",
		X"79",X"75",X"73",X"74",X"78",X"7A",X"7C",X"7D",X"7E",X"7C",X"79",X"78",X"7A",X"7E",X"80",X"7F",
		X"7C",X"7C",X"7E",X"82",X"85",X"87",X"89",X"89",X"87",X"82",X"80",X"81",X"84",X"85",X"86",X"87",
		X"86",X"82",X"7D",X"7B",X"7B",X"7D",X"7E",X"7F",X"7F",X"80",X"80",X"80",X"7F",X"7D",X"78",X"77",
		X"78",X"7B",X"7D",X"7F",X"80",X"81",X"7F",X"7B",X"7A",X"78",X"77",X"77",X"78",X"79",X"7A",X"7B",
		X"7D",X"7F",X"81",X"84",X"8A",X"90",X"93",X"96",X"97",X"97",X"97",X"96",X"92",X"8B",X"84",X"80",
		X"7F",X"7E",X"7B",X"76",X"71",X"70",X"71",X"73",X"72",X"70",X"6E",X"6F",X"73",X"77",X"78",X"77",
		X"76",X"77",X"77",X"79",X"7A",X"7C",X"7E",X"82",X"87",X"8D",X"90",X"93",X"94",X"94",X"90",X"8C",
		X"88",X"85",X"82",X"7F",X"7D",X"7A",X"79",X"78",X"78",X"77",X"77",X"77",X"7A",X"7F",X"83",X"84",
		X"83",X"81",X"82",X"85",X"88",X"88",X"85",X"81",X"80",X"81",X"83",X"83",X"84",X"83",X"83",X"82",
		X"81",X"7F",X"7E",X"7D",X"7A",X"76",X"72",X"71",X"72",X"74",X"74",X"72",X"71",X"71",X"71",X"72",
		X"73",X"75",X"7A",X"81",X"85",X"87",X"87",X"88",X"8B",X"90",X"92",X"91",X"8D",X"8A",X"88",X"86",
		X"84",X"82",X"80",X"7F",X"7E",X"7E",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7E",X"81",X"86",X"88",
		X"8A",X"8C",X"8C",X"8D",X"8C",X"8B",X"89",X"86",X"83",X"7E",X"78",X"73",X"6F",X"6C",X"6B",X"6C",
		X"70",X"72",X"75",X"78",X"7A",X"7A",X"78",X"77",X"77",X"78",X"79",X"7D",X"83",X"87",X"8A",X"8D",
		X"8F",X"90",X"90",X"8F",X"8C",X"86",X"82",X"7F",X"7C",X"7A",X"7B",X"7E",X"7F",X"81",X"81",X"81",
		X"7F",X"7B",X"7A",X"7A",X"7D",X"7E",X"80",X"81",X"81",X"80",X"7D",X"7B",X"7C",X"7E",X"80",X"80",
		X"80",X"7D",X"7B",X"79",X"78",X"78",X"78",X"79",X"79",X"7A",X"7B",X"7D",X"80",X"85",X"8A",X"8D",
		X"90",X"92",X"92",X"92",X"92",X"90",X"8E",X"8C",X"88",X"82",X"7B",X"78",X"76",X"76",X"74",X"71",
		X"6E",X"6D",X"6C",X"6C",X"6D",X"72",X"76",X"7B",X"7F",X"82",X"83",X"83",X"81",X"81",X"81",X"81",
		X"82",X"85",X"89",X"8B",X"8D",X"8E",X"8E",X"8E",X"8D",X"8A",X"85",X"80",X"7D",X"79",X"77",X"75",
		X"74",X"73",X"72",X"73",X"74",X"75",X"76",X"78",X"7A",X"80",X"85",X"87",X"87",X"86",X"88",X"8B",
		X"8E",X"8E",X"8B",X"87",X"84",X"81",X"7F",X"7D",X"7C",X"7B",X"7C",X"7E",X"81",X"83",X"84",X"85",
		X"86",X"85",X"83",X"7E",X"7B",X"7A",X"7B",X"7B",X"7C",X"7C",X"7C",X"7A",X"77",X"75",X"75",X"78",
		X"7A",X"7A",X"78",X"77",X"79",X"7C",X"7F",X"81",X"83",X"84",X"84",X"81",X"7F",X"7E",X"7E",X"7E",
		X"7D",X"7D",X"7E",X"7E",X"7F",X"80",X"83",X"88",X"8A",X"8B",X"89",X"87",X"86",X"85",X"84",X"85",
		X"88",X"8A",X"8A",X"8A",X"8A",X"89",X"88",X"86",X"83",X"81",X"7E",X"7C",X"7A",X"78",X"77",X"76",
		X"75",X"72",X"6E",X"6C",X"6C",X"6E",X"71",X"71",X"71",X"71",X"72",X"74",X"76",X"7B",X"81",X"86",
		X"88",X"88",X"89",X"8C",X"90",X"92",X"91",X"8F",X"8C",X"8C",X"8E",X"8F",X"8E",X"8D",X"8B",X"87",
		X"82",X"7D",X"79",X"76",X"74",X"72",X"71",X"73",X"77",X"78",X"78",X"77",X"77",X"77",X"78",X"7A",
		X"7D",X"82",X"84",X"87",X"89",X"8A",X"8B",X"8C",X"8C",X"8B",X"8A",X"88",X"84",X"7F",X"7C",X"7B",
		X"7C",X"7A",X"77",X"74",X"73",X"75",X"78",X"79",X"78",X"76",X"76",X"76",X"78",X"79",X"7A",X"7C",
		X"7E",X"82",X"87",X"8A",X"8C",X"8E",X"8F",X"8C",X"89",X"87",X"88",X"89",X"88",X"85",X"80",X"7E",
		X"7E",X"80",X"7F",X"7C",X"79",X"78",X"79",X"7B",X"7B",X"7A",X"78",X"78",X"7A",X"7D",X"7F",X"81",
		X"82",X"83",X"83",X"83",X"83",X"83",X"82",X"82",X"82",X"82",X"81",X"80",X"80",X"7F",X"7E",X"7D",
		X"7C",X"7C",X"7B",X"7B",X"7A",X"79",X"76",X"74",X"74",X"73",X"74",X"76",X"7B",X"7F",X"80",X"81",
		X"81",X"83",X"86",X"89",X"8B",X"8D",X"8E",X"8D",X"8A",X"87",X"85",X"83",X"81",X"7F",X"7E",X"7D",
		X"7C",X"7B",X"7B",X"7B",X"7B",X"7C",X"7F",X"82",X"85",X"88",X"89",X"8A",X"8B",X"8A",X"89",X"88",
		X"87",X"85",X"83",X"81",X"7E",X"7B",X"76",X"73",X"72",X"73",X"74",X"75",X"76",X"76",X"76",X"75",
		X"74",X"75",X"79",X"7C",X"7E",X"81",X"82",X"83",X"81",X"80",X"81",X"84",X"86",X"86",X"84",X"82",
		X"82",X"84",X"85",X"86",X"87",X"87",X"86",X"82",X"80",X"7E",X"7C",X"7B",X"7C",X"7E",X"80",X"81",
		X"7F",X"7D",X"7C",X"7B",X"7A",X"7A",X"7B",X"7E",X"81",X"83",X"83",X"82",X"81",X"81",X"80",X"80",
		X"82",X"85",X"86",X"85",X"82",X"80",X"7F",X"7E",X"7E",X"7F",X"82",X"83",X"82",X"80",X"7F",X"7E",
		X"7D",X"7C",X"7B",X"7B",X"7B",X"7E",X"81",X"82",X"82",X"80",X"7F",X"7E",X"7D",X"7C",X"7C",X"7C",
		X"7D",X"7F",X"83",X"85",X"86",X"88",X"88",X"86",X"82",X"80",X"80",X"81",X"80",X"7E",X"7C",X"7B",
		X"7B",X"7D",X"7D",X"7C",X"7A",X"79",X"78",X"77",X"78",X"7A",X"7D",X"80",X"82",X"84",X"85",X"87",
		X"88",X"88",X"85",X"82",X"7F",X"7D",X"7C",X"7B",X"7A",X"79",X"7A",X"7C",X"7F",X"81",X"83",X"84",
		X"85",X"84",X"82",X"81",X"82",X"83",X"84",X"84",X"84",X"83",X"83",X"83",X"82",X"81",X"7F",X"7B",
		X"78",X"76",X"74",X"74",X"73",X"73",X"74",X"76",X"7A",X"7E",X"81",X"84",X"86",X"88",X"89",X"8A",
		X"8A",X"8A",X"89",X"89",X"88",X"87",X"86",X"84",X"83",X"81",X"7F",X"7D",X"7B",X"79",X"78",X"77",
		X"74",X"72",X"71",X"71",X"71",X"73",X"76",X"7A",X"7C",X"7C",X"7D",X"7E",X"7F",X"81",X"83",X"87",
		X"8A",X"8B",X"8B",X"89",X"8A",X"8C",X"8E",X"8D",X"8A",X"86",X"85",X"85",X"86",X"84",X"81",X"7E",
		X"7D",X"7E",X"7E",X"7D",X"7A",X"78",X"77",X"79",X"7A",X"7A",X"79",X"77",X"78",X"7A",X"7D",X"7E",
		X"7D",X"7C",X"7C",X"7C",X"7D",X"7E",X"81",X"84",X"85",X"87",X"88",X"88",X"88",X"88",X"87",X"86",
		X"84",X"80",X"7E",X"7D",X"7E",X"7E",X"7E",X"7E",X"7E",X"7C",X"79",X"78",X"78",X"7A",X"7B",X"7B",
		X"7C",X"7D",X"7E",X"7F",X"80",X"7F",X"7D",X"7C",X"7B",X"7A",X"7B",X"7B",X"7C",X"7D",X"80",X"83",
		X"86",X"86",X"84",X"83",X"83",X"83",X"83",X"82",X"82",X"82",X"84",X"87",X"88",X"87",X"84",X"83",
		X"82",X"83",X"83",X"81",X"7F",X"7D",X"7E",X"7F",X"80",X"7F",X"7C",X"7B",X"7A",X"79",X"79",X"78",
		X"78",X"78",X"7A",X"7D",X"7E",X"7F",X"7E",X"7E",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",
		X"81",X"82",X"82",X"83",X"84",X"84",X"84",X"84",X"84",X"83",X"83",X"83",X"82",X"82",X"82",X"84",
		X"86",X"86",X"84",X"81",X"80",X"81",X"82",X"81",X"7E",X"7C",X"7B",X"7C",X"7D",X"7D",X"7E",X"7E",
		X"7D",X"7B",X"79",X"79",X"7A",X"7B",X"7C",X"7C",X"7D",X"7D",X"7D",X"7E",X"7E",X"7F",X"80",X"7F",
		X"7E",X"7C",X"7B",X"7C",X"7E",X"7F",X"80",X"81",X"82",X"82",X"83",X"83",X"83",X"83",X"82",X"80",
		X"7E",X"7C",X"7B",X"7B",X"7B",X"7C",X"7E",X"7F",X"7F",X"7E",X"7E",X"80",X"83",X"84",X"86",X"86",
		X"87",X"87",X"88",X"88",X"87",X"86",X"85",X"84",X"82",X"80",X"7D",X"7A",X"77",X"76",X"74",X"74",
		X"74",X"74",X"76",X"79",X"7C",X"7E",X"7F",X"7F",X"81",X"84",X"86",X"88",X"8A",X"8B",X"8C",X"8C",
		X"8B",X"8A",X"89",X"87",X"84",X"82",X"7F",X"7B",X"78",X"76",X"75",X"74",X"75",X"78",X"79",X"79",
		X"78",X"78",X"79",X"79",X"7A",X"7C",X"80",X"82",X"85",X"87",X"88",X"88",X"86",X"84",X"83",X"82",
		X"81",X"80",X"7F",X"7F",X"80",X"82",X"83",X"83",X"81",X"7F",X"7E",X"7D",X"7D",X"7F",X"81",X"83",
		X"84",X"85",X"85",X"83",X"80",X"7E",X"7D",X"7E",X"7E",X"7D",X"7B",X"7A",X"7B",X"7D",X"7E",X"7E",
		X"7D",X"7B",X"7B",X"7A",X"7A",X"7B",X"7E",X"7F",X"81",X"83",X"84",X"84",X"82",X"81",X"80",X"7F",
		X"7E",X"7E",X"7E",X"7E",X"80",X"82",X"84",X"84",X"82",X"81",X"80",X"7F",X"7F",X"7E",X"7E",X"7E",
		X"7E",X"7F",X"81",X"83",X"83",X"82",X"81",X"80",X"7F",X"7E",X"7D",X"7F",X"81",X"81",X"80",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7E",X"7E",X"7E",X"7E",X"7D",X"7D",X"7E",X"7E",X"7F",X"81",X"84",X"84",
		X"84",X"82",X"81",X"80",X"7F",X"7F",X"7E",X"7D",X"7E",X"7F",X"81",X"82",X"83",X"84",X"83",X"82",
		X"7F",X"7E",X"7D",X"7C",X"7B",X"7C",X"7D",X"7E",X"7F",X"80",X"80",X"81",X"81",X"81",X"81",X"80",
		X"7F",X"7D",X"7C",X"7B",X"7B",X"7C",X"7D",X"7E",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",X"7E",X"7C",X"7A",X"7A",
		X"79",X"79",X"7A",X"7C",X"7F",X"81",X"83",X"84",X"85",X"84",X"83",X"82",X"82",X"84",X"85",X"86",
		X"87",X"86",X"85",X"82",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7E",X"7C",X"7B",X"7A",X"79",
		X"79",X"79",X"7C",X"7E",X"7E",X"7E",X"7D",X"7D",X"7D",X"7E",X"7F",X"82",X"84",X"85",X"86",X"87",
		X"88",X"88",X"87",X"86",X"83",X"80",X"7F",X"80",X"80",X"7E",X"7C",X"7B",X"7B",X"7C",X"7D",X"7D",
		X"7C",X"7B",X"7C",X"7D",X"7F",X"7F",X"80",X"81",X"81",X"81",X"82",X"81",X"7F",X"7E",X"7D",X"7C",
		X"7B",X"7C",X"7E",X"80",X"80",X"80",X"7F",X"80",X"82",X"83",X"84",X"83",X"82",X"82",X"83",X"84",
		X"84",X"84",X"81",X"7F",X"7E",X"7E",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",
		X"7E",X"7E",X"7D",X"7D",X"7D",X"7D",X"7C",X"7B",X"79",X"79",X"78",X"79",X"79",X"79",X"7A",X"7B",
		X"7E",X"81",X"83",X"85",X"86",X"87",X"88",X"89",X"89",X"88",X"86",X"84",X"84",X"84",X"84",X"83",
		X"82",X"81",X"7F",X"7C",X"7B",X"7B",X"7B",X"7B",X"7C",X"7C",X"7C",X"7B",X"7A",X"79",X"79",X"7A",
		X"7A",X"7B",X"7D",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"81",X"82",X"82",X"83",X"83",
		X"85",X"87",X"88",X"89",X"89",X"89",X"89",X"88",X"87",X"86",X"84",X"82",X"7F",X"7C",X"79",X"77",
		X"76",X"74",X"74",X"73",X"73",X"74",X"75",X"78",X"7B",X"7C",X"7D",X"7D",X"7F",X"81",X"84",X"85",
		X"84",X"84",X"83",X"83",X"83",X"82",X"82",X"82",X"82",X"81",X"81",X"81",X"83",X"84",X"84",X"84",
		X"83",X"82",X"81",X"81",X"81",X"81",X"82",X"82",X"81",X"81",X"80",X"7E",X"7C",X"7C",X"7C",X"7D",
		X"7C",X"7B",X"7A",X"7B",X"7C",X"7D",X"7E",X"7F",X"7F",X"80",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"80",X"80",X"80",X"7F",X"7E",X"7E",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7C",
		X"7B",X"7C",X"7D",X"7E",X"7F",X"7F",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"81",
		X"81",X"82",X"82",X"83",X"84",X"85",X"86",X"88",X"88",X"89",X"89",X"89",X"89",X"88",X"87",X"85",
		X"84",X"82",X"80",X"7E",X"7B",X"78",X"76",X"74",X"72",X"71",X"71",X"71",X"72",X"73",X"75",X"77",
		X"79",X"7B",X"7D",X"7F",X"81",X"83",X"86",X"89",X"8B",X"8D",X"8E",X"8E",X"8D",X"8A",X"88",X"86",
		X"84",X"82",X"80",X"7F",X"7E",X"7E",X"7F",X"7F",X"7E",X"7D",X"7C",X"7C",X"7D",X"7D",X"7D",X"7E",
		X"7E",X"7E",X"7F",X"7E",X"7D",X"7C",X"7B",X"7A",X"7A",X"79",X"7B",X"7D",X"7E",X"7F",X"80",X"81",
		X"82",X"83",X"83",X"82",X"81",X"80",X"7F",X"7E",X"7E",X"7D",X"7D",X"7D",X"7E",X"7E",X"7F",X"80",
		X"83",X"84",X"84",X"83",X"82",X"82",X"82",X"81",X"81",X"81",X"82",X"83",X"83",X"82",X"80",X"7F",
		X"7E",X"7E",X"7E",X"7E",X"7F",X"80",X"81",X"81",X"81",X"81",X"81",X"80",X"7F",X"7D",X"7C",X"7D",
		X"7E",X"7E",X"7D",X"7C",X"7B",X"7B",X"7B",X"7B",X"7C",X"7E",X"7F",X"7F",X"7F",X"80",X"81",X"83",
		X"83",X"82",X"81",X"81",X"82",X"83",X"84",X"84",X"83",X"83",X"81",X"7F",X"7E",X"7D",X"7D",X"7D",
		X"7C",X"7C",X"7D",X"7F",X"80",X"81",X"80",X"7F",X"7F",X"80",X"81",X"82",X"82",X"83",X"82",X"81",
		X"7F",X"7E",X"7D",X"7D",X"7D",X"7C",X"7C",X"7D",X"7E",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"80",
		X"80",X"82",X"83",X"83",X"83",X"81",X"81",X"80",X"7F",X"7E",X"7E",X"7F",X"80",X"81",X"80",X"80",
		X"7F",X"80",X"81",X"82",X"81",X"7F",X"7E",X"7E",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7E",X"7D",X"7C",X"7B",X"7B",X"7B",X"7B",X"7C",X"7D",X"7E",X"80",X"80",X"80",X"80",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"81",X"82",X"84",X"85",X"84",X"83",X"82",X"82",X"83",
		X"83",X"82",X"81",X"80",X"80",X"81",X"82",X"81",X"81",X"81",X"80",X"80",X"7F",X"7E",X"7C",X"7B",
		X"7B",X"7C",X"7C",X"7D",X"7D",X"7D",X"7D",X"7D",X"7E",X"7D",X"7C",X"7C",X"7D",X"7E",X"7F",X"80",
		X"81",X"81",X"82",X"83",X"83",X"83",X"82",X"82",X"81",X"81",X"7F",X"7E",X"7D",X"7D",X"7C",X"7C",
		X"7D",X"7E",X"7E",X"7E",X"7D",X"7E",X"7F",X"80",X"81",X"82",X"83",X"83",X"84",X"84",X"84",X"83",
		X"81",X"80",X"7F",X"7E",X"7D",X"7C",X"7C",X"7C",X"7B",X"7B",X"7C",X"7D",X"7E",X"7F",X"80",X"80",
		X"81",X"83",X"85",X"86",X"87",X"87",X"87",X"87",X"86",X"85",X"84",X"83",X"82",X"80",X"7D",X"7C",
		X"7B",X"7B",X"7B",X"79",X"78",X"77",X"78",X"7A",X"7A",X"7A",X"79",X"7A",X"7C",X"7D",X"7F",X"7F",
		X"7F",X"80",X"80",X"80",X"81",X"83",X"84",X"84",X"84",X"83",X"83",X"83",X"84",X"84",X"83",X"82",
		X"81",X"81",X"81",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"7E",X"7E",X"7E",X"7F",
		X"80",X"80",X"7E",X"7E",X"7E",X"7E",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",
		X"80",X"80",X"7F",X"7F",X"7F",X"7E",X"7E",X"7E",X"7D",X"7C",X"7B",X"7B",X"7B",X"7C",X"7D",X"7D",
		X"7E",X"7E",X"7E",X"80",X"81",X"82",X"82",X"83",X"83",X"82",X"82",X"81",X"81",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"81",X"82",X"83",X"84",X"84",X"84",X"84",X"84",X"84",X"83",X"83",X"82",
		X"81",X"80",X"7F",X"7D",X"7C",X"7A",X"79",X"78",X"77",X"77",X"77",X"78",X"79",X"7A",X"7C",X"7E",
		X"7E",X"7F",X"80",X"81",X"82",X"83",X"85",X"86",X"87",X"88",X"88",X"88",X"87",X"86",X"85",X"83",
		X"81",X"7F",X"7E",X"7C",X"7B",X"7B",X"7B",X"7B",X"7C",X"7B",X"7B",X"7B",X"7B",X"7B",X"7C",X"7D",
		X"7F",X"80",X"81",X"82",X"82",X"82",X"81",X"81",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"80",X"81",
		X"82",X"81",X"81",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"80",X"81",X"82",X"81",X"81",X"80",
		X"80",X"81",X"80",X"80",X"7F",X"7E",X"7E",X"7E",X"7E",X"7E",X"7D",X"7D",X"7D",X"7D",X"7E",X"7F",
		X"80",X"81",X"82",X"82",X"82",X"82",X"82",X"82",X"81",X"80",X"7F",X"7E",X"7D",X"7D",X"7D",X"7D",
		X"7E",X"7E",X"7D",X"7E",X"7E",X"7F",X"7F",X"7F",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7F",
		X"7F",X"7F",X"80",X"80",X"81",X"81",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"81",X"81",X"82",X"82",X"83",X"83",X"83",X"82",X"82",X"81",X"80",X"7F",X"7D",X"7C",X"7B",
		X"7A",X"7A",X"79",X"79",X"79",X"7A",X"7B",X"7C",X"7C",X"7D",X"7D",X"7D",X"7D",X"7E",X"7E",X"7F",
		X"7F",X"80",X"80",X"81",X"82",X"83",X"84",X"85",X"84",X"84",X"83",X"83",X"83",X"82",X"82",X"82",
		X"81",X"80",X"80",X"80",X"81",X"81",X"81",X"81",X"81",X"80",X"80",X"7F",X"7F",X"7F",X"7E",X"7E",
		X"7D",X"7C",X"7C",X"7C",X"7C",X"7D",X"7D",X"7E",X"7E",X"7D",X"7D",X"7D",X"7E",X"7F",X"7F",X"80",
		X"80",X"7F",X"7F",X"80",X"81",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"81",X"81",X"81",
		X"80",X"7F",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7D",X"7D",X"7C",X"7C",X"7D",X"7D",X"7E",X"7E",
		X"7F",X"7F",X"7F",X"80",X"80",X"82",X"82",X"83",X"83",X"83",X"84",X"84",X"84",X"84",X"83",X"83",
		X"82",X"81",X"80",X"80",X"7E",X"7D",X"7C",X"7B",X"7A",X"79",X"79",X"79",X"79",X"7A",X"7B",X"7C",
		X"7D",X"7E",X"80",X"82",X"83",X"84",X"85",X"85",X"86",X"86",X"86",X"85",X"84",X"82",X"81",X"80",
		X"7F",X"7E",X"7D",X"7D",X"7D",X"7E",X"7E",X"7F",X"7F",X"7F",X"80",X"81",X"81",X"81",X"81",X"81",
		X"81",X"80",X"80",X"7F",X"7F",X"7D",X"7D",X"7C",X"7D",X"7D",X"7D",X"7E",X"7E",X"7F",X"7F",X"7F",
		X"7F",X"80",X"80",X"80",X"7F",X"7F",X"7E",X"7E",X"7E",X"7E",X"7D",X"7E",X"7E",X"7E",X"7F",X"80",
		X"81",X"82",X"83",X"83",X"83",X"83",X"83",X"82",X"82",X"83",X"83",X"83",X"82",X"81",X"80",X"80",
		X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"7E",X"7D",X"7C",X"7C",X"7C",X"7C",X"7C",X"7D",X"7D",X"7E",X"7F",X"7F",X"80",X"80",X"81",X"81",
		X"80",X"80",X"80",X"81",X"81",X"81",X"82",X"82",X"82",X"82",X"81",X"81",X"80",X"7E",X"7E",X"7D",
		X"7D",X"7D",X"7D",X"7E",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"81",X"82",
		X"82",X"82",X"82",X"81",X"81",X"80",X"80",X"7F",X"7F",X"7F",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"7E",X"7F",X"80",X"81",X"81",X"81",X"81",X"81",X"81",X"82",X"82",X"81",X"81",X"81",X"80",X"80",
		X"80",X"7F",X"7F",X"7E",X"7D",X"7D",X"7C",X"7C",X"7C",X"7C",X"7D",X"7E",X"7E",X"7E",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"80",X"81",X"80",X"80",X"80",X"80",X"81",X"81",X"81",X"81",X"81",X"81",X"80",
		X"80",X"80",X"80",X"80",X"80",X"81",X"81",X"80",X"80",X"80",X"7F",X"7E",X"7E",X"7E",X"7E",X"7F",
		X"7F",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"81",X"82",X"82",X"81",X"81",X"80",X"80",X"7F",X"7F",X"7F",X"80",X"80",X"81",X"81",
		X"81",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7E",
		X"7E",X"7E",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7E",
		X"7E",X"7F",X"7F",X"7F",X"7F",X"7E",X"7F",X"7F",X"80",X"80",X"81",X"81",X"80",X"80",X"80",X"80",
		X"80",X"7F",X"7F",X"7F",X"7E",X"7F",X"7F",X"80",X"80",X"80",X"7F",X"80",X"80",X"81",X"81",X"81",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"80",X"80",X"81",X"81",X"80",X"80",X"80",
		X"80",X"80",X"7F",X"7E",X"7E",X"7E",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",
		X"7F",X"7E",X"7E",X"7E",X"7F",X"7F",X"80",X"80",X"81",X"81",X"81",X"80",X"7F",X"7F",X"7F",X"7E",
		X"7F",X"7F",X"80",X"80",X"81",X"81",X"81",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"80",X"80",X"80",
		X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"81",X"80",X"80",X"80",X"80",X"80",
		X"7F",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7E",X"7E",X"7E",
		X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"80",X"80",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"80",X"80",X"80",X"80",
		X"80",X"80",X"81",X"81",X"80",X"80",X"80",X"80",X"81",X"81",X"81",X"81",X"81",X"80",X"80",X"80",
		X"7F",X"7F",X"7E",X"7E",X"7E",X"7E",X"7E",X"7D",X"7D",X"7E",X"7E",X"7E",X"7F",X"7F",X"80",X"80",
		X"80",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"80",X"80",X"80",X"7F",X"7F",
		X"7E",X"7E",X"7E",X"7D",X"7D",X"7D",X"7D",X"7D",X"7C",X"7D",X"7D",X"7D",X"7D",X"7D",X"7E",X"7E",
		X"7E",X"7F",X"7F",X"80",X"80",X"81",X"81",X"82",X"82",X"83",X"83",X"83",X"84",X"84",X"84",X"84",
		X"84",X"84",X"84",X"84",X"84",X"83",X"82",X"82",X"81",X"80",X"7F",X"7E",X"7E",X"7D",X"7C",X"7B",
		X"7B",X"7A",X"7A",X"79",X"79",X"79",X"79",X"7A",X"7A",X"7B",X"7C",X"7D",X"7E",X"7E",X"7F",X"80",
		X"80",X"81",X"81",X"82",X"82",X"83",X"83",X"84",X"84",X"84",X"84",X"84",X"83",X"83",X"82",X"82",
		X"81",X"81",X"81",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"7E",X"7E",X"7E",X"7F",X"7F",X"7F",X"7F",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"7F",X"7F",X"7F",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"80",X"80",X"7F",X"7F",X"7E",X"7E",X"7E",X"7E",X"7E",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"81",X"81",X"82",X"82",X"82",X"82",X"81",X"81",X"81",
		X"80",X"7F",X"7F",X"7E",X"7E",X"7E",X"7D",X"7D",X"7E",X"7E",X"7E",X"7F",X"7F",X"7F",X"7F",X"80",
		X"80",X"81",X"81",X"81",X"82",X"82",X"81",X"81",X"81",X"80",X"80",X"80",X"7F",X"7F",X"7E",X"7E",
		X"7E",X"7E",X"7E",X"7E",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"81",X"81",X"81",X"80",X"80",X"80",X"80",X"80",
		X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7E",X"7E",X"7E",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"7E",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"7D",X"7D",X"7D",X"7E",X"7E",X"7E",X"7E",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"81",X"80",
		X"80",X"81",X"81",X"81",X"81",X"81",X"80",X"80",X"80",X"80",X"81",X"81",X"81",X"81",X"80",X"80",
		X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"7F",X"7F",X"7F",X"7F",X"7E",X"7E",X"7E",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"7F",
		X"7F",X"80",X"80",X"80",X"80",X"80",X"81",X"81",X"81",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"81",X"81",
		X"81",X"81",X"81",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"80",X"7F",X"7F",
		X"7F",X"7F",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",
		X"7F",X"7F",X"7F",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"7F",X"7F",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
