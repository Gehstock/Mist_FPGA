library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity DEVILFISH_ROM_PGM_0 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of DEVILFISH_ROM_PGM_0 is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"AF",X"32",X"01",X"70",X"C3",X"8E",X"00",X"FF",X"C3",X"73",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"77",X"23",X"10",X"FC",X"C9",X"FF",X"FF",X"FF",X"11",X"20",X"00",X"77",X"19",X"10",X"FC",X"C9",
		X"85",X"6F",X"3E",X"00",X"8C",X"67",X"7E",X"C9",X"87",X"E1",X"D5",X"5F",X"16",X"00",X"19",X"5E",
		X"23",X"56",X"EB",X"D1",X"E9",X"FF",X"FF",X"FF",X"00",X"00",X"C3",X"B7",X"01",X"3A",X"0E",X"41",
		X"21",X"02",X"40",X"86",X"23",X"86",X"5F",X"23",X"7E",X"41",X"00",X"00",X"00",X"CD",X"87",X"10",
		X"CD",X"50",X"0C",X"00",X"00",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"21",X"E6",X"43",X"DD",X"7E",X"01",X"77",X"E6",X"0F",X"E7",
		X"C3",X"A7",X"11",X"E5",X"26",X"40",X"3A",X"A0",X"40",X"6F",X"CB",X"7E",X"28",X"0E",X"72",X"2C",
		X"73",X"2C",X"7D",X"FE",X"C0",X"30",X"02",X"3E",X"C0",X"32",X"A0",X"40",X"E1",X"C9",X"21",X"00",
		X"40",X"11",X"01",X"40",X"01",X"FF",X"03",X"36",X"00",X"ED",X"B0",X"3A",X"00",X"78",X"21",X"00",
		X"58",X"11",X"01",X"58",X"01",X"FF",X"00",X"36",X"00",X"ED",X"B0",X"3A",X"00",X"78",X"31",X"00",
		X"44",X"ED",X"56",X"FB",X"21",X"C0",X"40",X"06",X"40",X"3E",X"FF",X"D7",X"32",X"00",X"78",X"3A",
		X"00",X"78",X"AF",X"32",X"01",X"70",X"32",X"04",X"70",X"21",X"00",X"68",X"06",X"08",X"D7",X"CD",
		X"6E",X"10",X"21",X"C0",X"C0",X"22",X"A0",X"40",X"21",X"00",X"50",X"22",X"0B",X"40",X"3E",X"20",
		X"32",X"08",X"40",X"3A",X"00",X"78",X"3A",X"00",X"70",X"47",X"E6",X"01",X"3E",X"10",X"28",X"02",
		X"3E",X"15",X"32",X"17",X"40",X"3E",X"04",X"CB",X"50",X"20",X"02",X"3E",X"03",X"32",X"07",X"40",
		X"78",X"0F",X"0F",X"0F",X"E6",X"01",X"32",X"0F",X"40",X"3A",X"00",X"68",X"E6",X"C0",X"07",X"07",
		X"32",X"00",X"40",X"3A",X"00",X"78",X"21",X"00",X"50",X"11",X"01",X"50",X"01",X"FF",X"03",X"36",
		X"10",X"ED",X"B0",X"3A",X"00",X"78",X"3E",X"01",X"32",X"01",X"70",X"26",X"40",X"FB",X"3A",X"A1",
		X"40",X"6F",X"7E",X"87",X"30",X"05",X"CD",X"54",X"07",X"18",X"F0",X"E6",X"0F",X"4F",X"06",X"00",
		X"36",X"FF",X"23",X"5E",X"36",X"FF",X"2C",X"7D",X"FE",X"C0",X"30",X"02",X"3E",X"C0",X"32",X"A1",
		X"40",X"7B",X"21",X"5F",X"01",X"09",X"5E",X"23",X"56",X"21",X"2B",X"01",X"E5",X"EB",X"E9",X"8A",
		X"02",X"BC",X"02",X"1C",X"03",X"BF",X"03",X"57",X"04",X"10",X"04",X"73",X"04",X"C1",X"06",X"FE",
		X"01",X"C2",X"00",X"02",X"3A",X"F4",X"41",X"A7",X"C0",X"3A",X"2E",X"41",X"FE",X"10",X"DA",X"86",
		X"01",X"3E",X"10",X"32",X"2E",X"41",X"47",X"4F",X"21",X"FD",X"52",X"11",X"E0",X"FF",X"A7",X"28",
		X"05",X"36",X"2C",X"19",X"10",X"FB",X"3E",X"10",X"91",X"C8",X"47",X"CD",X"A4",X"01",X"79",X"77",
		X"19",X"10",X"FC",X"C9",X"3A",X"0D",X"41",X"E6",X"03",X"0E",X"30",X"C8",X"0E",X"21",X"3D",X"C8",
		X"0E",X"28",X"3D",X"C8",X"0E",X"2A",X"C9",X"C3",X"A3",X"07",X"4D",X"52",X"0D",X"52",X"CD",X"51",
		X"4F",X"52",X"0F",X"52",X"CF",X"51",X"51",X"52",X"11",X"52",X"D1",X"51",X"0B",X"52",X"13",X"52",
		X"8F",X"52",X"8F",X"51",X"21",X"EC",X"01",X"3A",X"5F",X"42",X"CB",X"5F",X"28",X"03",X"21",X"F6",
		X"01",X"3A",X"0D",X"41",X"E6",X"03",X"87",X"E7",X"23",X"56",X"5F",X"C9",X"3F",X"38",X"0A",X"34",
		X"52",X"34",X"C2",X"33",X"71",X"2F",X"63",X"38",X"2E",X"34",X"76",X"34",X"E6",X"33",X"72",X"2F",
		X"CD",X"63",X"02",X"CD",X"D4",X"01",X"D5",X"DD",X"E1",X"3A",X"10",X"41",X"A7",X"C8",X"47",X"21",
		X"BA",X"01",X"DD",X"E5",X"D1",X"78",X"3D",X"87",X"4F",X"E7",X"23",X"66",X"6F",X"79",X"87",X"EB",
		X"E7",X"EB",X"CD",X"28",X"02",X"10",X"E8",X"C9",X"1A",X"77",X"13",X"23",X"1A",X"77",X"D5",X"11",
		X"DF",X"FF",X"19",X"D1",X"13",X"1A",X"77",X"23",X"13",X"1A",X"77",X"C9",X"11",X"82",X"02",X"3A",
		X"5F",X"42",X"CB",X"5F",X"28",X"03",X"11",X"86",X"02",X"21",X"CC",X"01",X"3A",X"06",X"40",X"A7",
		X"3E",X"03",X"28",X"03",X"3A",X"5E",X"41",X"87",X"E7",X"23",X"66",X"6F",X"22",X"5C",X"41",X"CD",
		X"28",X"02",X"C9",X"3A",X"5B",X"41",X"A7",X"C2",X"3C",X"02",X"06",X"04",X"21",X"CC",X"01",X"11",
		X"86",X"02",X"78",X"3D",X"87",X"E7",X"23",X"66",X"6F",X"3E",X"4E",X"BE",X"CC",X"28",X"02",X"10",
		X"EB",X"C9",X"4E",X"4F",X"4C",X"4D",X"10",X"10",X"10",X"10",X"A7",X"C2",X"6F",X"01",X"01",X"20",
		X"00",X"2A",X"18",X"40",X"5E",X"23",X"56",X"23",X"EB",X"1A",X"FE",X"FF",X"28",X"05",X"77",X"13",
		X"09",X"18",X"F6",X"13",X"1A",X"FE",X"FF",X"20",X"0E",X"21",X"0A",X"40",X"3A",X"06",X"40",X"A7",
		X"20",X"03",X"21",X"BC",X"40",X"34",X"C9",X"ED",X"53",X"18",X"40",X"C9",X"3A",X"F4",X"41",X"A7",
		X"C0",X"3A",X"64",X"42",X"A7",X"20",X"4A",X"3A",X"5F",X"42",X"E6",X"0F",X"C0",X"3A",X"65",X"42",
		X"FE",X"05",X"20",X"04",X"AF",X"32",X"65",X"42",X"A7",X"28",X"1D",X"3D",X"28",X"1F",X"3D",X"28",
		X"21",X"3D",X"28",X"23",X"11",X"43",X"43",X"21",X"4B",X"50",X"72",X"2C",X"73",X"21",X"AB",X"53",
		X"72",X"2C",X"73",X"21",X"65",X"42",X"34",X"C9",X"11",X"10",X"10",X"18",X"EA",X"11",X"10",X"42",
		X"18",X"E5",X"11",X"10",X"43",X"18",X"E0",X"11",X"42",X"43",X"18",X"DB",X"11",X"43",X"43",X"18",
		X"D6",X"CD",X"F8",X"02",X"21",X"64",X"42",X"34",X"2C",X"36",X"00",X"C9",X"A7",X"C2",X"2D",X"03",
		X"21",X"08",X"51",X"CD",X"6C",X"03",X"21",X"F4",X"52",X"CD",X"6C",X"03",X"C9",X"FE",X"02",X"CA",
		X"5A",X"03",X"FE",X"04",X"CA",X"4C",X"03",X"FE",X"05",X"CA",X"53",X"03",X"2A",X"62",X"42",X"3E",
		X"2F",X"77",X"2C",X"77",X"11",X"DF",X"FF",X"19",X"77",X"2C",X"77",X"C9",X"21",X"08",X"51",X"CD",
		X"6C",X"03",X"C9",X"21",X"F4",X"52",X"CD",X"6C",X"03",X"C9",X"2A",X"60",X"42",X"36",X"37",X"2C",
		X"36",X"38",X"11",X"DF",X"FF",X"19",X"36",X"35",X"2C",X"36",X"36",X"C9",X"3A",X"5F",X"42",X"CB",
		X"5F",X"CA",X"83",X"03",X"36",X"46",X"2C",X"36",X"47",X"11",X"DF",X"FF",X"19",X"36",X"44",X"2C",
		X"36",X"45",X"C9",X"36",X"4A",X"2C",X"36",X"4B",X"11",X"DF",X"FF",X"19",X"36",X"48",X"2C",X"36",
		X"49",X"C9",X"F5",X"3A",X"0D",X"40",X"11",X"A2",X"40",X"0F",X"30",X"03",X"11",X"A5",X"40",X"F1",
		X"C9",X"00",X"01",X"00",X"50",X"01",X"00",X"00",X"02",X"00",X"00",X"03",X"00",X"10",X"00",X"00",
		X"50",X"01",X"00",X"00",X"02",X"00",X"00",X"03",X"00",X"50",X"03",X"00",X"10",X"00",X"00",X"CD",
		X"92",X"03",X"4F",X"87",X"81",X"4F",X"06",X"00",X"21",X"A1",X"03",X"3A",X"0D",X"41",X"A7",X"28",
		X"03",X"21",X"B0",X"03",X"09",X"A7",X"06",X"03",X"1A",X"8E",X"27",X"12",X"13",X"23",X"10",X"F8",
		X"D5",X"3A",X"0D",X"40",X"0F",X"30",X"02",X"3E",X"01",X"CD",X"10",X"04",X"D1",X"1B",X"21",X"AA",
		X"40",X"06",X"03",X"1A",X"BE",X"D8",X"20",X"05",X"1B",X"2B",X"10",X"F7",X"C9",X"CD",X"92",X"03",
		X"21",X"A8",X"40",X"06",X"03",X"1A",X"77",X"13",X"23",X"10",X"FA",X"3E",X"02",X"C3",X"10",X"04",
		X"21",X"A4",X"40",X"DD",X"21",X"61",X"53",X"A7",X"28",X"11",X"21",X"A7",X"40",X"DD",X"21",X"21",
		X"51",X"3D",X"28",X"07",X"21",X"AA",X"40",X"DD",X"21",X"41",X"52",X"11",X"E0",X"FF",X"06",X"03",
		X"0E",X"04",X"7E",X"0F",X"0F",X"0F",X"0F",X"CD",X"42",X"04",X"7E",X"CD",X"42",X"04",X"2B",X"10",
		X"F1",X"C9",X"E6",X"0F",X"28",X"08",X"0E",X"00",X"DD",X"77",X"00",X"DD",X"19",X"C9",X"79",X"A7",
		X"28",X"F6",X"3E",X"10",X"0D",X"18",X"F1",X"F5",X"21",X"A2",X"40",X"A7",X"28",X"09",X"21",X"A5",
		X"40",X"3D",X"28",X"03",X"21",X"A8",X"40",X"36",X"00",X"23",X"36",X"00",X"23",X"36",X"00",X"F1",
		X"C3",X"10",X"04",X"87",X"F5",X"21",X"E0",X"04",X"E6",X"7F",X"5F",X"16",X"00",X"19",X"5E",X"23",
		X"56",X"EB",X"5E",X"23",X"56",X"23",X"EB",X"01",X"E0",X"FF",X"F1",X"38",X"0E",X"FA",X"A5",X"04",
		X"1A",X"FE",X"3F",X"C8",X"D6",X"30",X"77",X"13",X"09",X"18",X"F5",X"1A",X"FE",X"3F",X"C8",X"36",
		X"10",X"13",X"09",X"18",X"F6",X"22",X"B5",X"40",X"ED",X"53",X"B7",X"40",X"EB",X"7B",X"E6",X"1F",
		X"47",X"87",X"C6",X"20",X"6F",X"26",X"40",X"22",X"B9",X"40",X"CB",X"3B",X"CB",X"3B",X"7A",X"E6",
		X"03",X"0F",X"0F",X"B3",X"E6",X"F8",X"4F",X"21",X"00",X"50",X"78",X"85",X"6F",X"11",X"20",X"00",
		X"43",X"36",X"10",X"19",X"10",X"FB",X"2A",X"B9",X"40",X"71",X"3E",X"01",X"32",X"BB",X"40",X"C9",
		X"14",X"05",X"27",X"05",X"3B",X"05",X"48",X"05",X"55",X"05",X"60",X"05",X"6D",X"05",X"7D",X"05",
		X"8D",X"05",X"9E",X"05",X"A8",X"05",X"BA",X"05",X"CF",X"05",X"DC",X"05",X"F2",X"05",X"0B",X"06",
		X"1C",X"06",X"2D",X"06",X"3E",X"06",X"4F",X"06",X"60",X"06",X"71",X"06",X"82",X"06",X"91",X"06",
		X"9C",X"06",X"AF",X"06",X"F4",X"52",X"53",X"45",X"54",X"40",X"46",X"49",X"53",X"48",X"40",X"41",
		X"53",X"40",X"42",X"41",X"49",X"54",X"3F",X"F1",X"52",X"50",X"55",X"53",X"48",X"40",X"53",X"54",
		X"41",X"52",X"54",X"40",X"42",X"55",X"54",X"54",X"4F",X"4E",X"3F",X"94",X"52",X"50",X"4C",X"41",
		X"59",X"45",X"52",X"40",X"4F",X"4E",X"45",X"3F",X"94",X"52",X"50",X"4C",X"41",X"59",X"45",X"52",
		X"40",X"54",X"57",X"4F",X"3F",X"60",X"52",X"48",X"49",X"5B",X"53",X"43",X"4F",X"52",X"45",X"3F",
		X"9F",X"53",X"40",X"43",X"52",X"45",X"44",X"49",X"54",X"40",X"40",X"40",X"3F",X"D1",X"52",X"49",
		X"4E",X"53",X"45",X"52",X"54",X"40",X"40",X"43",X"4F",X"49",X"4E",X"53",X"3F",X"BC",X"52",X"3C",
		X"56",X"49",X"53",X"49",X"4F",X"4E",X"40",X"40",X"31",X"39",X"38",X"34",X"3F",X"78",X"53",X"42",
		X"4F",X"4E",X"55",X"53",X"40",X"40",X"44",X"4F",X"47",X"47",X"49",X"45",X"40",X"3F",X"58",X"51",
		X"30",X"30",X"30",X"40",X"50",X"54",X"53",X"3F",X"D4",X"52",X"4F",X"4E",X"45",X"40",X"50",X"4C",
		X"41",X"59",X"45",X"52",X"40",X"4F",X"4E",X"4C",X"59",X"3F",X"F4",X"52",X"4F",X"4E",X"45",X"40",
		X"4F",X"52",X"40",X"54",X"57",X"4F",X"40",X"50",X"4C",X"41",X"59",X"45",X"52",X"53",X"3F",X"96",
		X"52",X"47",X"41",X"4D",X"45",X"40",X"40",X"4F",X"56",X"45",X"52",X"3F",X"2F",X"53",X"53",X"43",
		X"4F",X"52",X"45",X"40",X"41",X"44",X"56",X"41",X"4E",X"43",X"45",X"40",X"54",X"41",X"42",X"4C",
		X"45",X"3F",X"7D",X"53",X"3C",X"40",X"41",X"52",X"54",X"49",X"43",X"40",X"45",X"4C",X"45",X"43",
		X"54",X"52",X"4F",X"4E",X"49",X"43",X"40",X"4C",X"54",X"44",X"3F",X"52",X"52",X"31",X"30",X"30",
		X"40",X"31",X"35",X"30",X"40",X"3D",X"3D",X"3D",X"50",X"54",X"53",X"3F",X"55",X"52",X"31",X"35",
		X"30",X"40",X"32",X"30",X"30",X"40",X"3D",X"3D",X"3D",X"50",X"54",X"53",X"3F",X"58",X"52",X"32",
		X"30",X"30",X"40",X"32",X"35",X"30",X"40",X"3D",X"3D",X"3D",X"50",X"54",X"53",X"3F",X"5B",X"52",
		X"33",X"30",X"30",X"40",X"33",X"35",X"30",X"40",X"3D",X"3D",X"3D",X"50",X"54",X"53",X"3F",X"CB",
		X"52",X"57",X"45",X"4C",X"4C",X"40",X"44",X"4F",X"4E",X"45",X"40",X"4D",X"55",X"47",X"40",X"3F",
		X"EB",X"51",X"44",X"45",X"56",X"49",X"4C",X"40",X"46",X"49",X"53",X"48",X"40",X"43",X"41",X"4E",
		X"3F",X"ED",X"51",X"4F",X"4E",X"4C",X"59",X"40",X"42",X"45",X"40",X"43",X"41",X"55",X"47",X"48",
		X"54",X"3F",X"EF",X"51",X"57",X"48",X"45",X"4E",X"40",X"43",X"4C",X"41",X"4D",X"50",X"45",X"44",
		X"3F",X"F1",X"51",X"41",X"54",X"40",X"47",X"41",X"54",X"45",X"53",X"3F",X"F8",X"52",X"43",X"41",
		X"54",X"43",X"48",X"40",X"44",X"45",X"56",X"49",X"4C",X"40",X"46",X"49",X"53",X"48",X"3F",X"FA",
		X"52",X"52",X"45",X"54",X"55",X"52",X"4E",X"40",X"54",X"4F",X"40",X"43",X"41",X"42",X"49",X"4E",
		X"3F",X"A7",X"CA",X"CC",X"06",X"3D",X"CA",X"F1",X"06",X"C3",X"2F",X"07",X"21",X"1F",X"51",X"11",
		X"20",X"00",X"3A",X"0D",X"41",X"3C",X"FE",X"06",X"DA",X"DD",X"06",X"3E",X"05",X"47",X"A7",X"28",
		X"06",X"36",X"41",X"19",X"3D",X"20",X"F6",X"3E",X"05",X"90",X"47",X"36",X"10",X"19",X"10",X"FB",
		X"C9",X"3E",X"05",X"CD",X"73",X"04",X"3A",X"02",X"40",X"FE",X"63",X"38",X"02",X"3E",X"63",X"CD",
		X"15",X"07",X"47",X"E6",X"F0",X"28",X"07",X"0F",X"0F",X"0F",X"0F",X"32",X"9F",X"52",X"78",X"E6",
		X"0F",X"32",X"7F",X"52",X"C9",X"47",X"E6",X"0F",X"C6",X"00",X"27",X"4F",X"78",X"E6",X"F0",X"28",
		X"0B",X"0F",X"0F",X"0F",X"0F",X"47",X"AF",X"C6",X"16",X"27",X"10",X"FB",X"81",X"27",X"C9",X"3A",
		X"0E",X"41",X"47",X"4F",X"21",X"7F",X"50",X"11",X"20",X"00",X"A7",X"28",X"0B",X"FE",X"05",X"38",
		X"02",X"06",X"05",X"36",X"40",X"19",X"10",X"FB",X"3E",X"05",X"91",X"C8",X"D8",X"47",X"36",X"10",
		X"19",X"10",X"FB",X"C9",X"3A",X"5F",X"42",X"47",X"E6",X"0F",X"C0",X"11",X"E0",X"FF",X"21",X"E0",
		X"50",X"3A",X"0E",X"40",X"A7",X"28",X"22",X"36",X"02",X"CD",X"94",X"07",X"21",X"40",X"53",X"CD",
		X"92",X"07",X"3A",X"0D",X"40",X"A7",X"21",X"40",X"53",X"28",X"03",X"21",X"E0",X"50",X"CB",X"60",
		X"C8",X"3A",X"06",X"40",X"0F",X"D0",X"C3",X"9B",X"07",X"21",X"E0",X"50",X"CD",X"9B",X"07",X"C3",
		X"6C",X"07",X"36",X"01",X"19",X"36",X"25",X"19",X"36",X"20",X"C9",X"3E",X"10",X"77",X"19",X"77",
		X"19",X"77",X"C9",X"F5",X"C5",X"D5",X"E5",X"DD",X"E5",X"FD",X"E5",X"AF",X"32",X"01",X"70",X"21",
		X"20",X"40",X"11",X"00",X"58",X"01",X"80",X"00",X"ED",X"B0",X"3A",X"00",X"78",X"3A",X"15",X"40",
		X"32",X"16",X"40",X"3A",X"13",X"40",X"32",X"15",X"40",X"2A",X"10",X"40",X"22",X"13",X"40",X"21",
		X"12",X"40",X"3A",X"00",X"70",X"77",X"2B",X"3A",X"00",X"68",X"77",X"2B",X"3A",X"00",X"60",X"77",
		X"21",X"5F",X"42",X"35",X"20",X"02",X"2D",X"34",X"CD",X"17",X"08",X"CD",X"3A",X"08",X"CD",X"7D",
		X"08",X"CD",X"B2",X"08",X"CD",X"CC",X"2A",X"21",X"09",X"08",X"E5",X"3A",X"05",X"40",X"EF",X"E1",
		X"08",X"6B",X"09",X"9D",X"0E",X"A2",X"0F",X"A1",X"0F",X"FD",X"E1",X"DD",X"E1",X"E1",X"D1",X"C1",
		X"3E",X"01",X"32",X"01",X"70",X"F1",X"C9",X"21",X"10",X"40",X"7E",X"23",X"23",X"23",X"B6",X"23",
		X"23",X"2F",X"A6",X"23",X"A6",X"E6",X"03",X"C8",X"CB",X"47",X"C4",X"35",X"08",X"CB",X"4F",X"C8",
		X"21",X"26",X"41",X"34",X"C9",X"21",X"23",X"41",X"34",X"C9",X"21",X"22",X"41",X"7E",X"A7",X"20",
		X"34",X"23",X"B6",X"C8",X"35",X"2B",X"36",X"0F",X"3A",X"00",X"40",X"CB",X"47",X"28",X"17",X"21",
		X"02",X"40",X"7E",X"FE",X"63",X"C8",X"30",X"0B",X"34",X"11",X"01",X"07",X"CF",X"21",X"90",X"58",
		X"CB",X"CE",X"C9",X"36",X"63",X"C9",X"21",X"24",X"41",X"CB",X"46",X"28",X"05",X"36",X"00",X"C3",
		X"4F",X"08",X"36",X"01",X"C9",X"0F",X"0F",X"0F",X"32",X"03",X"60",X"35",X"C9",X"21",X"25",X"41",
		X"7E",X"A7",X"20",X"26",X"23",X"B6",X"C8",X"35",X"2B",X"36",X"0F",X"21",X"02",X"40",X"34",X"34",
		X"34",X"3A",X"00",X"40",X"CB",X"4F",X"20",X"02",X"34",X"34",X"7E",X"FE",X"63",X"C8",X"30",X"C3",
		X"11",X"01",X"07",X"CF",X"21",X"90",X"58",X"CB",X"CE",X"C9",X"0F",X"0F",X"0F",X"32",X"04",X"68",
		X"35",X"C9",X"3A",X"BB",X"40",X"0F",X"D0",X"2A",X"B9",X"40",X"7E",X"E6",X"07",X"20",X"1B",X"EB",
		X"2A",X"B7",X"40",X"7E",X"FE",X"3F",X"28",X"11",X"23",X"22",X"B7",X"40",X"D6",X"30",X"2A",X"B5",
		X"40",X"77",X"01",X"E0",X"FF",X"09",X"22",X"B5",X"40",X"EB",X"35",X"C0",X"AF",X"32",X"BB",X"40",
		X"C9",X"00",X"2A",X"0B",X"40",X"06",X"20",X"3E",X"10",X"D7",X"22",X"0B",X"40",X"21",X"08",X"40",
		X"35",X"C0",X"2D",X"2D",X"36",X"00",X"2D",X"34",X"AF",X"32",X"0A",X"40",X"21",X"2A",X"09",X"CD",
		X"12",X"09",X"11",X"04",X"06",X"CF",X"11",X"00",X"05",X"CF",X"1E",X"02",X"CF",X"AF",X"32",X"BC",
		X"40",X"C9",X"11",X"21",X"40",X"DD",X"21",X"0D",X"41",X"06",X"20",X"7E",X"DD",X"96",X"00",X"12",
		X"23",X"1C",X"EB",X"36",X"00",X"EB",X"1C",X"10",X"F2",X"C9",X"01",X"01",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"06",X"00",X"07",X"07",X"07",X"07",
		X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",
		X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"06",X"06",X"C9",X"00",X"21",X"40",X"0B",X"E5",
		X"3A",X"BC",X"40",X"EF",X"8F",X"0A",X"04",X"0B",X"DB",X"0B",X"E7",X"0B",X"28",X"0C",X"56",X"28",
		X"50",X"0C",X"9B",X"0C",X"B4",X"0C",X"C0",X"0C",X"D0",X"0C",X"ED",X"0C",X"7B",X"0D",X"8B",X"0D",
		X"EC",X"0D",X"B9",X"0F",X"D0",X"0F",X"F8",X"0F",X"31",X"10",X"87",X"10",X"A5",X"10",X"7D",X"0A",
		X"A6",X"09",X"56",X"28",X"37",X"0B",X"00",X"11",X"01",X"00",X"CF",X"11",X"02",X"00",X"CF",X"CD",
		X"1E",X"12",X"CD",X"86",X"12",X"CD",X"8D",X"14",X"CD",X"9D",X"12",X"CD",X"09",X"16",X"CD",X"7A",
		X"13",X"CD",X"07",X"15",X"CD",X"F5",X"14",X"3A",X"02",X"40",X"CD",X"8A",X"16",X"CD",X"F9",X"12",
		X"CD",X"B6",X"16",X"CD",X"41",X"18",X"CD",X"9D",X"18",X"CD",X"74",X"15",X"CD",X"43",X"16",X"CD",
		X"96",X"1E",X"CD",X"8A",X"16",X"CD",X"F2",X"09",X"CD",X"DD",X"27",X"CD",X"C8",X"29",X"CD",X"74",
		X"2A",X"C9",X"00",X"00",X"AF",X"32",X"61",X"41",X"DD",X"21",X"A0",X"42",X"DD",X"7E",X"00",X"A7",
		X"C8",X"CD",X"70",X"1B",X"CD",X"10",X"0A",X"78",X"4F",X"A7",X"CA",X"D4",X"23",X"C3",X"16",X"23",
		X"DD",X"7E",X"03",X"FE",X"C2",X"CA",X"2F",X"0A",X"FE",X"9A",X"CA",X"3F",X"0A",X"FE",X"82",X"CA",
		X"52",X"0A",X"FE",X"42",X"CA",X"62",X"0A",X"FE",X"5A",X"CA",X"72",X"0A",X"06",X"00",X"C9",X"06",
		X"20",X"DD",X"7E",X"04",X"FE",X"7A",X"C8",X"06",X"80",X"FE",X"5A",X"C8",X"06",X"00",X"C9",X"06",
		X"80",X"DD",X"7E",X"04",X"FE",X"9A",X"C8",X"06",X"00",X"FE",X"5A",X"C0",X"CD",X"A0",X"13",X"06",
		X"10",X"C9",X"06",X"10",X"DD",X"7E",X"04",X"FE",X"9A",X"C8",X"06",X"80",X"FE",X"CA",X"C8",X"06",
		X"00",X"C9",X"06",X"20",X"DD",X"7E",X"04",X"FE",X"CA",X"C8",X"06",X"40",X"FE",X"9A",X"C8",X"06",
		X"00",X"C9",X"06",X"40",X"DD",X"7E",X"04",X"FE",X"9A",X"C8",X"06",X"00",X"C9",X"3E",X"34",X"32",
		X"CA",X"50",X"32",X"CE",X"50",X"3D",X"32",X"AA",X"50",X"21",X"BC",X"40",X"34",X"C9",X"C9",X"CD",
		X"8E",X"0A",X"21",X"20",X"40",X"11",X"21",X"40",X"01",X"7F",X"00",X"36",X"00",X"ED",X"B0",X"3A",
		X"00",X"78",X"21",X"00",X"41",X"11",X"01",X"41",X"01",X"1F",X"00",X"36",X"00",X"ED",X"B0",X"21",
		X"A0",X"42",X"11",X"A1",X"42",X"01",X"FF",X"00",X"36",X"00",X"ED",X"B0",X"21",X"02",X"50",X"22",
		X"0B",X"40",X"21",X"08",X"40",X"36",X"20",X"21",X"BC",X"40",X"34",X"AF",X"32",X"06",X"40",X"32",
		X"5F",X"42",X"32",X"0D",X"40",X"32",X"0E",X"40",X"21",X"00",X"68",X"06",X"03",X"D7",X"21",X"80",
		X"58",X"21",X"D0",X"41",X"06",X"10",X"D7",X"06",X"80",X"D7",X"3E",X"FF",X"32",X"00",X"78",X"CD",
		X"F3",X"0A",X"C9",X"21",X"F2",X"05",X"06",X"20",X"AF",X"86",X"23",X"10",X"FC",X"32",X"BD",X"41",
		X"3A",X"00",X"78",X"C9",X"2A",X"0B",X"40",X"06",X"1E",X"3E",X"10",X"D7",X"11",X"02",X"00",X"19",
		X"22",X"0B",X"40",X"21",X"08",X"40",X"35",X"C0",X"21",X"4A",X"09",X"CD",X"12",X"09",X"CD",X"6E",
		X"10",X"21",X"BC",X"40",X"34",X"23",X"36",X"30",X"11",X"01",X"07",X"CF",X"11",X"07",X"06",X"CF",
		X"21",X"4E",X"0B",X"22",X"18",X"40",X"C9",X"21",X"BD",X"40",X"35",X"C0",X"2D",X"36",X"00",X"C9",
		X"3A",X"02",X"40",X"A7",X"C8",X"21",X"05",X"40",X"34",X"AF",X"32",X"0A",X"40",X"C9",X"0E",X"50",
		X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",
		X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",
		X"FF",X"0F",X"50",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"31",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"31",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"FF",X"10",X"50",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"32",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"FF",X"11",X"50",X"30",X"30",X"30",X"30",X"30",X"30",X"30",
		X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",
		X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"FF",X"FF",X"21",X"BD",X"40",X"35",X"C0",
		X"36",X"05",X"11",X"00",X"00",X"CF",X"C9",X"11",X"E0",X"42",X"21",X"01",X"18",X"01",X"20",X"00",
		X"ED",X"B0",X"DD",X"21",X"E0",X"42",X"AF",X"CD",X"76",X"17",X"21",X"E3",X"42",X"36",X"78",X"2C",
		X"36",X"F8",X"11",X"A0",X"42",X"21",X"BD",X"27",X"01",X"20",X"00",X"ED",X"B0",X"21",X"A3",X"42",
		X"36",X"7A",X"2C",X"36",X"EA",X"21",X"BC",X"40",X"34",X"AF",X"32",X"BE",X"40",X"32",X"4F",X"41",
		X"11",X"00",X"06",X"CF",X"CD",X"8C",X"0C",X"C9",X"CD",X"8D",X"14",X"CD",X"07",X"15",X"CD",X"F9",
		X"12",X"CD",X"7A",X"0E",X"CD",X"9D",X"18",X"CD",X"74",X"15",X"CD",X"43",X"16",X"CD",X"96",X"1E",
		X"CD",X"25",X"0E",X"CD",X"40",X"0E",X"CD",X"DD",X"27",X"CD",X"C8",X"29",X"CD",X"74",X"2A",X"C9",
		X"21",X"73",X"2F",X"22",X"18",X"40",X"21",X"02",X"50",X"22",X"0B",X"40",X"21",X"08",X"40",X"36",
		X"20",X"21",X"60",X"40",X"11",X"61",X"40",X"01",X"3F",X"00",X"36",X"00",X"ED",X"B0",X"21",X"BC",
		X"40",X"34",X"2C",X"36",X"30",X"3E",X"4F",X"32",X"C0",X"41",X"3E",X"04",X"32",X"C1",X"41",X"21",
		X"05",X"0E",X"22",X"C2",X"41",X"21",X"60",X"40",X"22",X"C4",X"41",X"C9",X"3A",X"BD",X"41",X"FE",
		X"F0",X"C8",X"21",X"52",X"2E",X"11",X"00",X"40",X"ED",X"B0",X"C9",X"2A",X"0B",X"40",X"06",X"1C",
		X"3E",X"10",X"D7",X"11",X"04",X"00",X"19",X"22",X"0B",X"40",X"21",X"08",X"40",X"35",X"C0",X"21",
		X"BC",X"40",X"34",X"C9",X"21",X"BD",X"40",X"35",X"C0",X"36",X"05",X"11",X"00",X"00",X"CF",X"C9",
		X"11",X"0D",X"06",X"CF",X"11",X"0E",X"06",X"CF",X"21",X"BC",X"40",X"34",X"2C",X"36",X"10",X"C9",
		X"21",X"BD",X"40",X"35",X"C0",X"36",X"20",X"2D",X"34",X"2A",X"C2",X"41",X"ED",X"5B",X"C4",X"41",
		X"01",X"04",X"00",X"ED",X"B0",X"22",X"C2",X"41",X"ED",X"53",X"C4",X"41",X"C9",X"21",X"BD",X"40",
		X"35",X"C0",X"36",X"A0",X"2D",X"34",X"21",X"02",X"50",X"22",X"0B",X"40",X"21",X"08",X"40",X"36",
		X"20",X"16",X"06",X"21",X"C0",X"41",X"5E",X"34",X"CF",X"2A",X"C2",X"41",X"ED",X"5B",X"C4",X"41",
		X"01",X"04",X"00",X"ED",X"B0",X"22",X"C2",X"41",X"ED",X"53",X"C4",X"41",X"3A",X"C1",X"41",X"3D",
		X"C8",X"32",X"C1",X"41",X"21",X"BC",X"40",X"35",X"35",X"C9",X"30",X"30",X"30",X"10",X"10",X"10",
		X"30",X"30",X"30",X"10",X"31",X"10",X"10",X"10",X"10",X"10",X"31",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"32",X"10",X"30",X"30",X"30",X"10",X"10",X"10",X"30",X"30",X"30",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"30",X"10",X"10",X"30",X"10",X"30",X"10",X"10",X"30",X"30",X"33",X"10",X"30",X"10",X"30",X"33",
		X"34",X"30",X"30",X"10",X"10",X"30",X"10",X"30",X"10",X"10",X"30",X"3A",X"5F",X"42",X"CB",X"47",
		X"C0",X"21",X"BD",X"40",X"35",X"C0",X"36",X"B0",X"2D",X"34",X"C9",X"2A",X"0B",X"40",X"06",X"1C",
		X"3E",X"10",X"D7",X"11",X"04",X"00",X"19",X"22",X"0B",X"40",X"21",X"08",X"40",X"35",X"C0",X"21",
		X"60",X"40",X"AF",X"06",X"40",X"D7",X"11",X"14",X"06",X"CF",X"1C",X"CF",X"1C",X"CF",X"1C",X"CF",
		X"1C",X"CF",X"1C",X"CF",X"21",X"38",X"53",X"36",X"4C",X"2C",X"36",X"4D",X"21",X"58",X"53",X"36",
		X"4E",X"2C",X"36",X"4F",X"CD",X"CC",X"0D",X"21",X"BC",X"40",X"34",X"C9",X"01",X"09",X"09",X"21",
		X"49",X"52",X"11",X"2A",X"0D",X"1A",X"77",X"13",X"D5",X"11",X"20",X"00",X"19",X"D1",X"10",X"F5",
		X"06",X"09",X"0D",X"C8",X"D5",X"11",X"E1",X"FE",X"19",X"D1",X"18",X"E9",X"3A",X"5F",X"42",X"CB",
		X"47",X"C0",X"21",X"BD",X"40",X"35",X"C0",X"2D",X"34",X"AF",X"32",X"5F",X"42",X"ED",X"4F",X"3E",
		X"03",X"32",X"5E",X"42",X"C9",X"28",X"04",X"03",X"88",X"48",X"00",X"03",X"88",X"28",X"04",X"02",
		X"A0",X"48",X"00",X"02",X"A0",X"28",X"04",X"04",X"B8",X"48",X"00",X"04",X"B8",X"28",X"04",X"01",
		X"D0",X"48",X"00",X"01",X"D0",X"00",X"DD",X"21",X"A0",X"42",X"CD",X"70",X"1B",X"3A",X"BE",X"40",
		X"A7",X"C0",X"3A",X"A4",X"42",X"FE",X"A8",X"CA",X"A0",X"13",X"FE",X"28",X"CA",X"A0",X"13",X"C9",
		X"3A",X"A0",X"42",X"A7",X"C8",X"DD",X"21",X"A0",X"42",X"0E",X"20",X"3A",X"BE",X"40",X"A7",X"20",
		X"13",X"3A",X"A4",X"42",X"FE",X"22",X"D2",X"60",X"0E",X"0E",X"10",X"3E",X"01",X"32",X"BE",X"40",
		X"79",X"C3",X"13",X"23",X"3A",X"4F",X"41",X"A7",X"C2",X"60",X"0E",X"3A",X"A4",X"42",X"FE",X"A2",
		X"38",X"E7",X"3E",X"01",X"32",X"4F",X"41",X"C3",X"60",X"0E",X"3A",X"A4",X"42",X"FE",X"21",X"C0",
		X"11",X"00",X"43",X"21",X"21",X"18",X"01",X"20",X"00",X"ED",X"B0",X"3E",X"02",X"DD",X"21",X"00",
		X"43",X"CD",X"76",X"17",X"21",X"03",X"43",X"36",X"78",X"2C",X"36",X"02",X"C9",X"21",X"48",X"0F",
		X"E5",X"AF",X"32",X"BC",X"40",X"32",X"5E",X"42",X"3A",X"0A",X"40",X"EF",X"B2",X"0E",X"F7",X"0E",
		X"3A",X"0F",X"21",X"20",X"40",X"11",X"21",X"40",X"01",X"7F",X"00",X"36",X"00",X"ED",X"B0",X"21",
		X"A0",X"42",X"11",X"A1",X"42",X"01",X"FF",X"00",X"36",X"00",X"ED",X"B0",X"21",X"4A",X"09",X"CD",
		X"12",X"09",X"AF",X"32",X"BB",X"40",X"21",X"02",X"50",X"22",X"0B",X"40",X"21",X"09",X"40",X"36",
		X"10",X"2C",X"34",X"AF",X"06",X"06",X"21",X"0B",X"41",X"D7",X"06",X"06",X"21",X"00",X"42",X"D7",
		X"32",X"21",X"42",X"32",X"20",X"42",X"C9",X"2A",X"0B",X"40",X"06",X"1D",X"3E",X"10",X"D7",X"11",
		X"03",X"00",X"19",X"06",X"1D",X"D7",X"19",X"22",X"0B",X"40",X"21",X"09",X"40",X"35",X"C0",X"2C",
		X"34",X"CD",X"6E",X"10",X"AF",X"32",X"0D",X"40",X"11",X"01",X"07",X"CF",X"11",X"01",X"06",X"FF",
		X"1E",X"08",X"CF",X"1C",X"CF",X"3A",X"17",X"40",X"47",X"E6",X"0F",X"32",X"78",X"51",X"78",X"E6",
		X"F0",X"C8",X"0F",X"0F",X"0F",X"0F",X"32",X"98",X"51",X"C9",X"3A",X"02",X"40",X"A7",X"C8",X"3D",
		X"11",X"0A",X"06",X"28",X"01",X"1C",X"CF",X"C9",X"3A",X"11",X"40",X"CB",X"47",X"C2",X"8B",X"0F",
		X"CB",X"4F",X"C8",X"3A",X"02",X"40",X"FE",X"02",X"D8",X"D6",X"02",X"32",X"02",X"40",X"21",X"00",
		X"01",X"22",X"0D",X"40",X"AF",X"32",X"0A",X"40",X"3E",X"03",X"32",X"05",X"40",X"3E",X"01",X"32",
		X"06",X"40",X"11",X"04",X"06",X"CF",X"3A",X"07",X"40",X"32",X"0E",X"41",X"32",X"03",X"42",X"11",
		X"00",X"04",X"CF",X"3A",X"0E",X"40",X"0F",X"D0",X"1C",X"CF",X"C9",X"3A",X"02",X"40",X"A7",X"28",
		X"0A",X"3D",X"32",X"02",X"40",X"21",X"00",X"00",X"C3",X"61",X"0F",X"3E",X"01",X"32",X"05",X"40",
		X"C9",X"C9",X"00",X"3A",X"0A",X"40",X"EF",X"B9",X"0F",X"D0",X"0F",X"F8",X"0F",X"31",X"10",X"87",
		X"10",X"93",X"10",X"A7",X"11",X"56",X"28",X"82",X"29",X"3E",X"36",X"32",X"0B",X"41",X"32",X"00",
		X"42",X"AF",X"32",X"2C",X"41",X"32",X"2D",X"41",X"32",X"2E",X"41",X"CD",X"1C",X"2A",X"34",X"C9",
		X"00",X"AF",X"21",X"20",X"40",X"06",X"80",X"D7",X"CD",X"1C",X"2A",X"34",X"21",X"08",X"40",X"36",
		X"20",X"21",X"00",X"50",X"22",X"0B",X"40",X"AF",X"32",X"2E",X"41",X"32",X"62",X"41",X"32",X"5B",
		X"41",X"21",X"80",X"58",X"06",X"80",X"D7",X"C9",X"2A",X"0B",X"40",X"06",X"20",X"3E",X"10",X"D7",
		X"22",X"0B",X"40",X"21",X"08",X"40",X"35",X"C0",X"21",X"4A",X"09",X"CD",X"12",X"09",X"CD",X"19",
		X"10",X"22",X"18",X"40",X"CD",X"1C",X"2A",X"34",X"C9",X"21",X"27",X"10",X"3A",X"0D",X"41",X"E6",
		X"03",X"87",X"E7",X"23",X"66",X"6F",X"C9",X"9A",X"34",X"1D",X"30",X"87",X"38",X"2C",X"3C",X"70",
		X"2F",X"AF",X"32",X"5F",X"42",X"CD",X"6E",X"10",X"21",X"09",X"40",X"36",X"30",X"CD",X"1C",X"2A",
		X"34",X"3A",X"0E",X"40",X"0F",X"38",X"21",X"11",X"00",X"05",X"CF",X"1E",X"02",X"CF",X"11",X"04",
		X"06",X"CF",X"1E",X"02",X"3A",X"0D",X"40",X"A7",X"28",X"02",X"1E",X"03",X"CF",X"3A",X"06",X"40",
		X"A7",X"C8",X"3E",X"10",X"32",X"B0",X"58",X"C9",X"11",X"01",X"05",X"CF",X"18",X"D9",X"3A",X"0F",
		X"40",X"A7",X"28",X"0A",X"3A",X"0D",X"40",X"A7",X"28",X"04",X"3E",X"00",X"18",X"02",X"3E",X"01",
		X"32",X"06",X"70",X"32",X"07",X"70",X"C9",X"21",X"09",X"40",X"35",X"C0",X"36",X"05",X"11",X"00",
		X"00",X"CF",X"C9",X"00",X"CD",X"6E",X"12",X"11",X"00",X"02",X"CF",X"11",X"02",X"07",X"CF",X"1E",
		X"00",X"CF",X"1E",X"01",X"CF",X"21",X"2E",X"41",X"7E",X"FE",X"10",X"30",X"14",X"3A",X"5F",X"42",
		X"E6",X"07",X"20",X"01",X"34",X"11",X"01",X"00",X"CF",X"AF",X"32",X"62",X"41",X"32",X"0A",X"41",
		X"C9",X"11",X"A0",X"42",X"21",X"BD",X"27",X"01",X"20",X"00",X"ED",X"B0",X"CD",X"1C",X"2A",X"34",
		X"3E",X"10",X"32",X"5C",X"42",X"ED",X"5F",X"E6",X"03",X"47",X"3E",X"01",X"28",X"03",X"07",X"10",
		X"FD",X"32",X"B0",X"58",X"C9",X"3A",X"F4",X"41",X"A7",X"C2",X"27",X"11",X"CD",X"ED",X"28",X"AF",
		X"47",X"21",X"A0",X"42",X"D7",X"06",X"40",X"21",X"60",X"40",X"D7",X"21",X"F1",X"41",X"36",X"1B",
		X"2C",X"36",X"04",X"2C",X"36",X"07",X"2C",X"36",X"01",X"21",X"42",X"50",X"22",X"F5",X"41",X"3E",
		X"FF",X"32",X"F7",X"41",X"AF",X"32",X"B0",X"58",X"3A",X"0D",X"41",X"E6",X"03",X"3C",X"47",X"3E",
		X"01",X"07",X"10",X"FD",X"32",X"A0",X"58",X"3A",X"F3",X"41",X"A7",X"CA",X"34",X"11",X"3D",X"32",
		X"F3",X"41",X"E1",X"C9",X"2A",X"F5",X"41",X"3A",X"F1",X"41",X"A7",X"CA",X"88",X"11",X"47",X"3A",
		X"F2",X"41",X"CD",X"72",X"11",X"3E",X"10",X"77",X"19",X"10",X"FA",X"3A",X"F2",X"41",X"3D",X"CA",
		X"57",X"11",X"32",X"F2",X"41",X"18",X"E0",X"11",X"21",X"00",X"19",X"22",X"F5",X"41",X"21",X"F1",
		X"41",X"7E",X"FE",X"02",X"DA",X"88",X"11",X"D6",X"02",X"77",X"2C",X"36",X"04",X"2C",X"36",X"07",
		X"E1",X"C9",X"11",X"01",X"00",X"FE",X"04",X"C8",X"11",X"20",X"00",X"FE",X"03",X"C8",X"11",X"FF",
		X"FF",X"FE",X"02",X"C8",X"11",X"E0",X"FF",X"C9",X"AF",X"32",X"F1",X"41",X"11",X"13",X"06",X"CF",
		X"21",X"F7",X"41",X"35",X"C2",X"A5",X"11",X"21",X"0D",X"41",X"34",X"AF",X"32",X"F4",X"41",X"32",
		X"10",X"41",X"32",X"0A",X"40",X"E1",X"C9",X"00",X"3A",X"5F",X"42",X"A7",X"20",X"1E",X"3A",X"0D",
		X"40",X"A7",X"20",X"0D",X"3A",X"2C",X"41",X"FE",X"FF",X"28",X"11",X"3C",X"32",X"2C",X"41",X"18",
		X"0B",X"3A",X"2D",X"41",X"FE",X"FF",X"28",X"04",X"3C",X"32",X"2D",X"41",X"00",X"3A",X"F4",X"41",
		X"A7",X"20",X"04",X"11",X"01",X"00",X"CF",X"11",X"02",X"00",X"CF",X"CD",X"1E",X"12",X"CD",X"86",
		X"12",X"CD",X"8D",X"14",X"CD",X"C0",X"12",X"CD",X"9D",X"12",X"CD",X"09",X"16",X"CD",X"7A",X"13",
		X"CD",X"07",X"15",X"CD",X"F5",X"14",X"CD",X"8A",X"16",X"CD",X"F9",X"12",X"CD",X"B6",X"16",X"CD",
		X"41",X"18",X"CD",X"9D",X"18",X"CD",X"74",X"15",X"CD",X"43",X"16",X"CD",X"96",X"1E",X"CD",X"8A",
		X"16",X"CD",X"E4",X"22",X"CD",X"DD",X"27",X"CD",X"C8",X"29",X"CD",X"74",X"2A",X"C9",X"21",X"5B",
		X"41",X"DD",X"21",X"A0",X"42",X"7E",X"A7",X"C8",X"2C",X"7E",X"DD",X"BE",X"11",X"C0",X"2C",X"7E",
		X"DD",X"BE",X"10",X"C0",X"CD",X"7C",X"12",X"3A",X"66",X"41",X"A7",X"20",X"10",X"3A",X"B0",X"58",
		X"E6",X"DF",X"32",X"B0",X"58",X"3E",X"01",X"32",X"A0",X"58",X"32",X"66",X"41",X"21",X"09",X"40",
		X"35",X"35",X"3E",X"90",X"BE",X"DA",X"A5",X"11",X"21",X"10",X"41",X"34",X"AF",X"32",X"09",X"40",
		X"32",X"5B",X"41",X"32",X"5E",X"41",X"32",X"66",X"41",X"DD",X"36",X"08",X"04",X"C9",X"21",X"38",
		X"00",X"06",X"50",X"AF",X"86",X"23",X"10",X"FC",X"32",X"F0",X"41",X"C9",X"3A",X"06",X"40",X"A7",
		X"C8",X"11",X"04",X"03",X"CF",X"C9",X"3A",X"F4",X"41",X"A7",X"C2",X"E5",X"10",X"3A",X"10",X"41",
		X"FE",X"09",X"C0",X"21",X"09",X"40",X"35",X"C2",X"A5",X"11",X"C3",X"E5",X"10",X"3A",X"08",X"51",
		X"FE",X"46",X"CA",X"B9",X"12",X"FE",X"4A",X"CA",X"B9",X"12",X"3A",X"F4",X"52",X"FE",X"46",X"28",
		X"03",X"FE",X"4A",X"C0",X"11",X"05",X"02",X"CF",X"C9",X"11",X"04",X"02",X"CF",X"C3",X"AA",X"12",
		X"3A",X"0F",X"41",X"0F",X"D8",X"21",X"A4",X"40",X"3A",X"0D",X"40",X"0F",X"30",X"03",X"21",X"A7",
		X"40",X"3A",X"17",X"40",X"47",X"7E",X"E6",X"0F",X"07",X"07",X"07",X"07",X"4F",X"2D",X"7E",X"E6",
		X"F0",X"0F",X"0F",X"0F",X"0F",X"B1",X"B8",X"D8",X"21",X"0E",X"41",X"34",X"11",X"02",X"07",X"CF",
		X"2C",X"36",X"01",X"21",X"90",X"58",X"CB",X"C6",X"C9",X"DD",X"21",X"E0",X"42",X"06",X"06",X"DD",
		X"7E",X"00",X"A7",X"C4",X"0E",X"13",X"11",X"20",X"00",X"DD",X"19",X"10",X"F2",X"C9",X"DD",X"7E",
		X"0D",X"A7",X"20",X"53",X"DD",X"36",X"0F",X"02",X"3A",X"0C",X"41",X"A7",X"28",X"03",X"DD",X"34",
		X"0F",X"3A",X"0F",X"41",X"A7",X"DD",X"34",X"0F",X"28",X"03",X"DD",X"34",X"0F",X"3A",X"0D",X"40",
		X"A7",X"3A",X"2D",X"41",X"20",X"03",X"3A",X"2C",X"41",X"FE",X"2F",X"38",X"0A",X"DD",X"34",X"0F",
		X"FE",X"6F",X"38",X"03",X"DD",X"34",X"0F",X"DD",X"7E",X"17",X"A7",X"28",X"03",X"DD",X"34",X"0F",
		X"DD",X"7E",X"0F",X"FE",X"08",X"38",X"04",X"DD",X"36",X"0F",X"08",X"DD",X"7E",X"07",X"A7",X"C8",
		X"DD",X"35",X"0F",X"DD",X"35",X"0F",X"C9",X"DD",X"36",X"0F",X"03",X"3D",X"CA",X"18",X"13",X"3D",
		X"CA",X"18",X"13",X"DD",X"36",X"0F",X"04",X"C3",X"18",X"13",X"DD",X"21",X"A0",X"42",X"DD",X"7E",
		X"00",X"A7",X"C8",X"3A",X"2E",X"41",X"A7",X"C8",X"CD",X"09",X"14",X"3A",X"0F",X"40",X"A7",X"28",
		X"09",X"3A",X"0D",X"40",X"A7",X"3A",X"11",X"40",X"20",X"03",X"3A",X"10",X"40",X"E6",X"10",X"C8",
		X"DD",X"66",X"10",X"DD",X"6E",X"11",X"DD",X"7E",X"04",X"CB",X"57",X"28",X"08",X"E6",X"03",X"28",
		X"04",X"11",X"E0",X"FF",X"19",X"23",X"DD",X"7E",X"03",X"CB",X"57",X"28",X"49",X"E6",X"03",X"28",
		X"45",X"22",X"60",X"42",X"11",X"02",X"02",X"CF",X"21",X"2E",X"41",X"35",X"3E",X"01",X"32",X"C0",
		X"58",X"C9",X"3A",X"06",X"40",X"A7",X"C8",X"ED",X"5F",X"E6",X"07",X"C8",X"3A",X"F0",X"41",X"FE",
		X"F4",X"C8",X"3A",X"02",X"40",X"FE",X"05",X"38",X"06",X"ED",X"5F",X"32",X"FC",X"43",X"C9",X"3A",
		X"5F",X"42",X"E6",X"50",X"C0",X"3A",X"02",X"40",X"A7",X"28",X"05",X"3D",X"32",X"02",X"40",X"C9",
		X"3C",X"3C",X"32",X"02",X"40",X"C9",X"2B",X"18",X"B8",X"CD",X"70",X"1B",X"DD",X"66",X"10",X"DD",
		X"6E",X"11",X"7E",X"FE",X"10",X"C2",X"8B",X"14",X"23",X"7E",X"FE",X"10",X"C2",X"8B",X"14",X"11",
		X"DF",X"FF",X"19",X"7E",X"FE",X"10",X"C2",X"8B",X"14",X"23",X"7E",X"FE",X"10",X"C2",X"8B",X"14",
		X"DD",X"7E",X"04",X"CB",X"57",X"CA",X"4E",X"14",X"E6",X"03",X"CA",X"4E",X"14",X"19",X"7E",X"FE",
		X"10",X"C2",X"8B",X"14",X"23",X"7E",X"FE",X"10",X"C2",X"8B",X"14",X"C3",X"69",X"14",X"DD",X"7E",
		X"03",X"CB",X"57",X"C8",X"E6",X"03",X"C8",X"23",X"7E",X"FE",X"10",X"C2",X"8B",X"14",X"11",X"20",
		X"00",X"19",X"7E",X"FE",X"10",X"C2",X"8B",X"14",X"C9",X"DD",X"7E",X"03",X"CB",X"57",X"C8",X"E6",
		X"03",X"C8",X"23",X"7E",X"FE",X"10",X"C2",X"8B",X"14",X"11",X"20",X"00",X"19",X"7E",X"FE",X"10",
		X"C2",X"8B",X"14",X"19",X"7E",X"FE",X"10",X"C2",X"8B",X"14",X"C9",X"E1",X"C9",X"DD",X"21",X"A0",
		X"42",X"06",X"08",X"FD",X"21",X"60",X"40",X"DD",X"CB",X"00",X"46",X"20",X"10",X"DD",X"7E",X"01",
		X"A7",X"20",X"0A",X"FD",X"36",X"00",X"00",X"FD",X"36",X"03",X"00",X"18",X"28",X"3A",X"0D",X"40",
		X"A7",X"CA",X"E1",X"14",X"3A",X"0F",X"40",X"A7",X"CA",X"E1",X"14",X"DD",X"7E",X"04",X"3C",X"FD",
		X"77",X"00",X"DD",X"7E",X"03",X"3D",X"FD",X"77",X"03",X"DD",X"7E",X"09",X"FD",X"77",X"01",X"DD",
		X"7E",X"08",X"FD",X"77",X"02",X"11",X"20",X"00",X"DD",X"19",X"1E",X"04",X"FD",X"19",X"10",X"B7",
		X"C9",X"DD",X"7E",X"04",X"3D",X"FD",X"77",X"00",X"FD",X"77",X"00",X"DD",X"7E",X"03",X"3C",X"FD",
		X"77",X"03",X"C3",X"C9",X"14",X"3A",X"5F",X"42",X"A7",X"C0",X"3A",X"5E",X"42",X"E6",X"03",X"FE",
		X"03",X"C0",X"11",X"00",X"02",X"CF",X"C9",X"00",X"DD",X"21",X"A0",X"42",X"DD",X"7E",X"00",X"A7",
		X"28",X"22",X"DD",X"7E",X"18",X"FE",X"30",X"28",X"03",X"C3",X"34",X"15",X"DD",X"86",X"0A",X"DD",
		X"77",X"09",X"3A",X"5F",X"42",X"E6",X"05",X"20",X"0B",X"DD",X"34",X"0A",X"DD",X"7E",X"0A",X"E6",
		X"03",X"DD",X"77",X"0A",X"00",X"DD",X"21",X"E0",X"42",X"06",X"06",X"11",X"20",X"00",X"DD",X"7E",
		X"00",X"A7",X"20",X"05",X"DD",X"19",X"10",X"F6",X"C9",X"DD",X"CB",X"0A",X"7E",X"20",X"18",X"DD",
		X"CB",X"07",X"7E",X"20",X"EF",X"3A",X"5F",X"42",X"E6",X"05",X"20",X"0B",X"DD",X"34",X"0A",X"DD",
		X"7E",X"0A",X"E6",X"03",X"DD",X"77",X"0A",X"DD",X"7E",X"0A",X"E6",X"03",X"DD",X"86",X"18",X"DD",
		X"77",X"09",X"18",X"D0",X"DD",X"21",X"E0",X"42",X"06",X"06",X"DD",X"7E",X"00",X"A7",X"28",X"0E",
		X"DD",X"7E",X"05",X"E6",X"0C",X"28",X"63",X"DD",X"7E",X"04",X"E6",X"07",X"28",X"08",X"11",X"20",
		X"00",X"DD",X"19",X"10",X"E5",X"C9",X"CD",X"70",X"1B",X"DD",X"66",X"10",X"DD",X"6E",X"11",X"7E",
		X"FE",X"37",X"20",X"EA",X"3E",X"10",X"CD",X"41",X"03",X"DD",X"36",X"1A",X"FF",X"DD",X"7E",X"0D",
		X"FE",X"02",X"30",X"12",X"DD",X"36",X"18",X"27",X"DD",X"36",X"09",X"27",X"DD",X"36",X"07",X"81",
		X"DD",X"36",X"1F",X"10",X"18",X"C8",X"00",X"DD",X"7E",X"07",X"E6",X"7F",X"FE",X"02",X"28",X"BE",
		X"DD",X"36",X"1F",X"10",X"3C",X"F6",X"80",X"DD",X"77",X"07",X"E6",X"7F",X"FE",X"01",X"20",X"1E",
		X"DD",X"36",X"18",X"26",X"DD",X"36",X"09",X"26",X"18",X"A4",X"DD",X"7E",X"05",X"E6",X"03",X"28",
		X"9D",X"DD",X"7E",X"03",X"18",X"94",X"22",X"62",X"42",X"11",X"01",X"02",X"CF",X"C9",X"DD",X"36",
		X"18",X"27",X"DD",X"36",X"09",X"27",X"C3",X"8E",X"15",X"DD",X"21",X"A0",X"42",X"CD",X"70",X"1B",
		X"DD",X"66",X"10",X"DD",X"6E",X"11",X"7E",X"FE",X"46",X"28",X"03",X"FE",X"4A",X"C0",X"DD",X"CB",
		X"03",X"56",X"28",X"06",X"DD",X"7E",X"03",X"E6",X"03",X"C0",X"DD",X"CB",X"04",X"56",X"28",X"06",
		X"DD",X"7E",X"04",X"E6",X"03",X"C0",X"CD",X"F6",X"15",X"3E",X"02",X"32",X"C0",X"58",X"21",X"2E",
		X"41",X"34",X"C9",X"DD",X"21",X"E0",X"42",X"06",X"06",X"DD",X"CB",X"07",X"7E",X"C2",X"58",X"16",
		X"11",X"20",X"00",X"DD",X"19",X"10",X"F2",X"C9",X"DD",X"35",X"1F",X"20",X"F3",X"DD",X"34",X"02",
		X"DD",X"7E",X"02",X"FE",X"02",X"CA",X"7C",X"16",X"DD",X"36",X"1F",X"10",X"1E",X"00",X"DD",X"7E",
		X"18",X"FE",X"27",X"28",X"02",X"1E",X"04",X"DD",X"73",X"18",X"18",X"D4",X"DD",X"36",X"02",X"00",
		X"DD",X"7E",X"07",X"E6",X"7F",X"DD",X"77",X"07",X"18",X"C6",X"DD",X"21",X"E0",X"42",X"AF",X"32",
		X"0A",X"41",X"11",X"20",X"00",X"06",X"06",X"DD",X"36",X"0E",X"00",X"DD",X"CB",X"00",X"46",X"20",
		X"0B",X"DD",X"CB",X"01",X"46",X"20",X"05",X"DD",X"19",X"10",X"EC",X"C9",X"21",X"0A",X"41",X"34",
		X"DD",X"36",X"0E",X"01",X"18",X"F1",X"11",X"00",X"01",X"CF",X"21",X"0B",X"41",X"7E",X"A7",X"20",
		X"02",X"36",X"2F",X"21",X"2C",X"41",X"3A",X"0D",X"40",X"A7",X"28",X"03",X"21",X"2D",X"41",X"7E",
		X"FE",X"3A",X"3E",X"06",X"30",X"09",X"7E",X"FE",X"28",X"3E",X"05",X"30",X"02",X"3E",X"04",X"21",
		X"0A",X"41",X"BE",X"C8",X"D8",X"21",X"5D",X"42",X"34",X"3A",X"5C",X"42",X"BE",X"C0",X"36",X"00",
		X"2D",X"36",X"D0",X"3E",X"10",X"32",X"4B",X"50",X"32",X"4C",X"50",X"32",X"AB",X"53",X"32",X"AC",
		X"53",X"3E",X"E0",X"32",X"64",X"42",X"3A",X"0B",X"41",X"FE",X"36",X"28",X"22",X"DD",X"21",X"E0",
		X"42",X"11",X"20",X"00",X"06",X"06",X"DD",X"7E",X"0E",X"A7",X"20",X"0E",X"3A",X"06",X"40",X"A7",
		X"28",X"06",X"ED",X"5F",X"CB",X"47",X"28",X"1D",X"18",X"62",X"DD",X"19",X"10",X"E8",X"C9",X"00",
		X"DD",X"21",X"E0",X"42",X"11",X"E0",X"42",X"CD",X"48",X"17",X"DD",X"21",X"00",X"43",X"11",X"00",
		X"43",X"CD",X"8F",X"17",X"C9",X"DD",X"E5",X"D1",X"CD",X"9C",X"17",X"21",X"01",X"18",X"01",X"20",
		X"00",X"ED",X"B0",X"3E",X"35",X"21",X"0B",X"41",X"96",X"21",X"B6",X"17",X"47",X"3A",X"0D",X"41",
		X"A7",X"28",X"11",X"21",X"BF",X"17",X"FE",X"01",X"28",X"0A",X"21",X"C8",X"17",X"FE",X"02",X"28",
		X"03",X"21",X"D1",X"17",X"78",X"E7",X"47",X"87",X"80",X"21",X"F5",X"17",X"E7",X"7E",X"DD",X"77",
		X"08",X"23",X"7E",X"DD",X"77",X"0D",X"23",X"7E",X"DD",X"77",X"18",X"C9",X"DD",X"E5",X"D1",X"CD",
		X"9C",X"17",X"21",X"21",X"18",X"01",X"20",X"00",X"ED",X"B0",X"18",X"B7",X"21",X"0B",X"41",X"35",
		X"7E",X"23",X"FE",X"1B",X"20",X"03",X"36",X"01",X"C9",X"FE",X"12",X"20",X"03",X"36",X"02",X"C9",
		X"FE",X"09",X"C0",X"36",X"03",X"C9",X"00",X"00",X"01",X"01",X"02",X"00",X"00",X"00",X"03",X"01",
		X"01",X"01",X"00",X"02",X"03",X"00",X"01",X"02",X"01",X"02",X"01",X"01",X"03",X"00",X"00",X"03",
		X"01",X"02",X"01",X"00",X"03",X"00",X"01",X"01",X"02",X"03",X"02",X"03",X"00",X"01",X"01",X"00",
		X"03",X"00",X"02",X"03",X"02",X"01",X"00",X"02",X"03",X"01",X"01",X"03",X"02",X"03",X"00",X"01",
		X"02",X"03",X"00",X"01",X"03",X"03",X"00",X"04",X"02",X"01",X"04",X"04",X"02",X"08",X"01",X"03",
		X"08",X"01",X"00",X"00",X"58",X"F0",X"04",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"00",X"00",X"58",X"00",X"08",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"DD",X"21",X"60",X"43",X"06",X"02",X"00",X"DD",X"7E",X"00",X"A7",X"20",X"08",X"11",
		X"20",X"00",X"DD",X"19",X"10",X"F2",X"C9",X"AF",X"DD",X"77",X"17",X"3A",X"0B",X"41",X"FE",X"08",
		X"38",X"ED",X"DD",X"7E",X"03",X"21",X"A3",X"42",X"56",X"BA",X"38",X"1C",X"DD",X"7E",X"17",X"F6",
		X"11",X"DD",X"77",X"17",X"DD",X"7E",X"04",X"21",X"A4",X"42",X"56",X"BA",X"38",X"14",X"DD",X"7E",
		X"17",X"F6",X"44",X"DD",X"77",X"17",X"18",X"C7",X"DD",X"7E",X"17",X"F6",X"22",X"DD",X"77",X"17",
		X"18",X"E2",X"DD",X"7E",X"17",X"F6",X"88",X"DD",X"77",X"17",X"C3",X"4F",X"18",X"DD",X"21",X"E0",
		X"42",X"FD",X"21",X"30",X"41",X"3E",X"06",X"32",X"09",X"40",X"21",X"98",X"19",X"E5",X"DD",X"7E",
		X"00",X"A7",X"C8",X"DD",X"7E",X"06",X"A7",X"C0",X"DD",X"CB",X"07",X"7E",X"C0",X"DD",X"7E",X"1A",
		X"A7",X"C4",X"55",X"19",X"DD",X"7E",X"0F",X"FD",X"BE",X"00",X"C4",X"16",X"19",X"FD",X"6E",X"01",
		X"FD",X"66",X"02",X"29",X"FD",X"75",X"01",X"FD",X"74",X"02",X"FD",X"6E",X"03",X"FD",X"66",X"04",
		X"ED",X"6A",X"FD",X"75",X"03",X"FD",X"74",X"04",X"D0",X"FD",X"34",X"01",X"20",X"03",X"FD",X"34",
		X"02",X"DD",X"7E",X"05",X"0F",X"DA",X"6C",X"1D",X"0F",X"DA",X"96",X"1D",X"0F",X"DA",X"3F",X"1D",
		X"CD",X"15",X"1C",X"DD",X"7E",X"04",X"E6",X"0F",X"FE",X"08",X"CA",X"AD",X"19",X"FE",X"00",X"CA",
		X"AD",X"19",X"DD",X"34",X"04",X"C9",X"FD",X"77",X"00",X"07",X"07",X"21",X"31",X"19",X"E7",X"FD",
		X"77",X"01",X"23",X"7E",X"FD",X"77",X"02",X"23",X"7E",X"FD",X"77",X"03",X"23",X"FD",X"77",X"04",
		X"C9",X"55",X"55",X"55",X"55",X"D5",X"6A",X"D5",X"6A",X"A5",X"94",X"A5",X"94",X"AD",X"B5",X"AD",
		X"B5",X"6D",X"DB",X"6D",X"DB",X"6D",X"DB",X"6D",X"DB",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"3A",X"5F",X"42",X"CB",X"47",X"C0",X"DD",X"35",X"1A",X"C0",X"DD",
		X"7E",X"0D",X"FE",X"02",X"30",X"0D",X"DD",X"36",X"18",X"04",X"DD",X"36",X"09",X"04",X"DD",X"36",
		X"07",X"00",X"C9",X"DD",X"7E",X"18",X"FE",X"04",X"28",X"11",X"DD",X"36",X"07",X"01",X"DD",X"36",
		X"18",X"04",X"DD",X"36",X"09",X"04",X"DD",X"36",X"1A",X"20",X"C9",X"DD",X"36",X"18",X"08",X"DD",
		X"36",X"09",X"08",X"DD",X"36",X"07",X"00",X"C9",X"3A",X"09",X"40",X"3D",X"C8",X"32",X"09",X"40",
		X"11",X"20",X"00",X"DD",X"19",X"11",X"05",X"00",X"FD",X"19",X"C3",X"AA",X"18",X"CD",X"C5",X"19",
		X"CD",X"CE",X"1B",X"CD",X"AE",X"1C",X"CD",X"F7",X"1C",X"DD",X"7E",X"12",X"E6",X"0B",X"20",X"21",
		X"3E",X"04",X"C3",X"29",X"1B",X"CD",X"70",X"1B",X"DD",X"66",X"10",X"DD",X"6E",X"11",X"AF",X"DD",
		X"77",X"12",X"DD",X"77",X"13",X"DD",X"77",X"14",X"DD",X"77",X"15",X"DD",X"77",X"16",X"4D",X"44",
		X"C9",X"DD",X"7E",X"17",X"A7",X"C2",X"97",X"1B",X"3A",X"5B",X"41",X"A7",X"20",X"2D",X"DD",X"E5",
		X"E1",X"7D",X"FE",X"20",X"28",X"25",X"FE",X"40",X"28",X"21",X"ED",X"5F",X"21",X"5F",X"42",X"86",
		X"CB",X"47",X"28",X"17",X"DD",X"7E",X"12",X"E6",X"0F",X"4F",X"07",X"07",X"07",X"07",X"B1",X"4F",
		X"ED",X"5F",X"CB",X"47",X"79",X"CA",X"A0",X"1B",X"C3",X"AB",X"1B",X"DD",X"66",X"04",X"DD",X"6E",
		X"03",X"CD",X"A3",X"1A",X"EB",X"3A",X"A4",X"42",X"67",X"3A",X"A3",X"42",X"6F",X"CD",X"A3",X"1A",
		X"EB",X"22",X"50",X"41",X"ED",X"53",X"52",X"41",X"21",X"FF",X"FF",X"22",X"54",X"41",X"DD",X"CB",
		X"12",X"46",X"CA",X"51",X"1A",X"3E",X"01",X"32",X"58",X"41",X"2A",X"50",X"41",X"2D",X"CD",X"B0",
		X"1A",X"DD",X"CB",X"12",X"4E",X"CA",X"64",X"1A",X"3E",X"02",X"32",X"58",X"41",X"2A",X"50",X"41",
		X"2C",X"CD",X"B0",X"1A",X"DD",X"CB",X"12",X"56",X"CA",X"77",X"1A",X"3E",X"04",X"32",X"58",X"41",
		X"2A",X"50",X"41",X"25",X"CD",X"B0",X"1A",X"DD",X"CB",X"12",X"5E",X"28",X"0C",X"3E",X"08",X"32",
		X"58",X"41",X"2A",X"50",X"41",X"24",X"CD",X"B0",X"1A",X"00",X"DD",X"7E",X"12",X"32",X"63",X"41",
		X"CD",X"C0",X"1D",X"DD",X"7E",X"12",X"21",X"63",X"41",X"BE",X"C2",X"E1",X"19",X"3A",X"59",X"41",
		X"C3",X"29",X"1B",X"CB",X"3D",X"CB",X"3D",X"CB",X"3D",X"CB",X"3C",X"CB",X"3C",X"CB",X"3C",X"C9",
		X"22",X"56",X"41",X"DD",X"E5",X"FD",X"E5",X"DD",X"21",X"52",X"41",X"FD",X"21",X"56",X"41",X"CD",
		X"E3",X"1A",X"FD",X"E1",X"DD",X"E1",X"EB",X"2A",X"54",X"41",X"A7",X"ED",X"52",X"D8",X"CC",X"DC",
		X"1A",X"ED",X"53",X"54",X"41",X"3A",X"58",X"41",X"32",X"59",X"41",X"C9",X"ED",X"5F",X"CB",X"47",
		X"C8",X"EB",X"C9",X"DD",X"7E",X"00",X"FD",X"46",X"00",X"90",X"D2",X"F2",X"1A",X"78",X"DD",X"46",
		X"00",X"90",X"CD",X"0B",X"1B",X"E5",X"DD",X"7E",X"01",X"FD",X"46",X"01",X"90",X"D2",X"05",X"1B",
		X"78",X"DD",X"46",X"01",X"90",X"CD",X"0B",X"1B",X"C1",X"09",X"C9",X"67",X"5F",X"2E",X"00",X"55",
		X"0E",X"08",X"29",X"D2",X"17",X"1B",X"19",X"0D",X"C2",X"12",X"1B",X"C9",X"DD",X"7E",X"12",X"A6",
		X"32",X"59",X"41",X"C2",X"89",X"1A",X"23",X"18",X"F3",X"00",X"DD",X"77",X"05",X"0F",X"38",X"08",
		X"0F",X"38",X"0F",X"0F",X"38",X"16",X"18",X"1E",X"DD",X"7E",X"16",X"DD",X"77",X"06",X"DD",X"35",
		X"03",X"C9",X"DD",X"7E",X"15",X"DD",X"77",X"06",X"DD",X"34",X"03",X"C9",X"DD",X"7E",X"14",X"DD",
		X"77",X"06",X"DD",X"35",X"04",X"C9",X"DD",X"7E",X"13",X"DD",X"77",X"06",X"DD",X"34",X"04",X"C9",
		X"01",X"02",X"04",X"08",X"02",X"04",X"08",X"01",X"04",X"08",X"01",X"02",X"08",X"01",X"02",X"04",
		X"26",X"14",X"DD",X"6E",X"04",X"7D",X"2F",X"6F",X"C5",X"06",X"02",X"7D",X"E6",X"F8",X"CB",X"27",
		X"6F",X"7C",X"17",X"67",X"10",X"F5",X"DD",X"77",X"10",X"DD",X"7E",X"03",X"E6",X"F8",X"0F",X"0F",
		X"0F",X"B5",X"DD",X"77",X"11",X"C1",X"C9",X"ED",X"5F",X"CB",X"47",X"DD",X"7E",X"17",X"28",X"0B",
		X"0F",X"38",X"13",X"0F",X"38",X"16",X"0F",X"38",X"19",X"18",X"1D",X"07",X"38",X"1A",X"07",X"38",
		X"11",X"07",X"38",X"08",X"18",X"00",X"21",X"60",X"1B",X"C3",X"1C",X"1B",X"21",X"64",X"1B",X"C3",
		X"1C",X"1B",X"21",X"68",X"1B",X"C3",X"1C",X"1B",X"21",X"6C",X"1B",X"C3",X"1C",X"1B",X"00",X"11",
		X"C0",X"FF",X"69",X"60",X"19",X"7E",X"CD",X"87",X"27",X"28",X"0D",X"FE",X"31",X"28",X"26",X"DD",
		X"7E",X"12",X"E6",X"F7",X"DD",X"77",X"12",X"C9",X"23",X"7E",X"CD",X"87",X"27",X"28",X"0D",X"FE",
		X"32",X"28",X"18",X"DD",X"7E",X"12",X"E6",X"F7",X"DD",X"77",X"12",X"C9",X"DD",X"7E",X"12",X"F6",
		X"08",X"DD",X"77",X"12",X"C9",X"DD",X"36",X"13",X"01",X"18",X"DD",X"DD",X"7E",X"13",X"F6",X"02",
		X"DD",X"77",X"13",X"18",X"E7",X"DD",X"7E",X"04",X"FE",X"EF",X"D8",X"DD",X"7E",X"0F",X"A7",X"20",
		X"11",X"DD",X"7E",X"19",X"D6",X"20",X"DD",X"77",X"19",X"28",X"02",X"E1",X"C9",X"DD",X"36",X"04",
		X"01",X"C9",X"DD",X"7E",X"19",X"D6",X"40",X"DD",X"77",X"19",X"28",X"F1",X"E1",X"C9",X"DD",X"7E",
		X"04",X"FE",X"01",X"C0",X"DD",X"7E",X"0F",X"A7",X"20",X"11",X"DD",X"7E",X"19",X"D6",X"10",X"DD",
		X"77",X"19",X"28",X"02",X"E1",X"C9",X"DD",X"36",X"04",X"EF",X"C9",X"DD",X"7E",X"19",X"D6",X"20",
		X"DD",X"77",X"19",X"28",X"F1",X"E1",X"C9",X"00",X"11",X"20",X"00",X"69",X"60",X"19",X"7E",X"CD",
		X"87",X"27",X"28",X"0D",X"FE",X"31",X"28",X"26",X"DD",X"7E",X"12",X"E6",X"FB",X"DD",X"77",X"12",
		X"C9",X"23",X"7E",X"CD",X"87",X"27",X"28",X"0D",X"FE",X"32",X"28",X"18",X"DD",X"7E",X"12",X"E6",
		X"FB",X"DD",X"77",X"12",X"C9",X"DD",X"7E",X"12",X"F6",X"04",X"DD",X"77",X"12",X"C9",X"DD",X"36",
		X"14",X"01",X"18",X"DD",X"DD",X"7E",X"14",X"F6",X"02",X"DD",X"77",X"14",X"18",X"E7",X"11",X"FF",
		X"FF",X"69",X"60",X"19",X"7E",X"CD",X"87",X"27",X"28",X"0D",X"FE",X"34",X"28",X"29",X"DD",X"7E",
		X"12",X"E6",X"FE",X"DD",X"77",X"12",X"C9",X"11",X"E0",X"FF",X"19",X"7E",X"CD",X"87",X"27",X"28",
		X"0D",X"FE",X"33",X"28",X"18",X"DD",X"7E",X"12",X"E6",X"FE",X"DD",X"77",X"12",X"C9",X"DD",X"7E",
		X"12",X"F6",X"01",X"DD",X"77",X"12",X"C9",X"DD",X"36",X"16",X"01",X"18",X"DA",X"DD",X"7E",X"16",
		X"F6",X"02",X"DD",X"77",X"16",X"18",X"E7",X"69",X"60",X"23",X"23",X"7E",X"CD",X"87",X"27",X"28",
		X"0D",X"FE",X"34",X"28",X"29",X"DD",X"7E",X"12",X"E6",X"FD",X"DD",X"77",X"12",X"C9",X"11",X"E0",
		X"FF",X"19",X"7E",X"CD",X"87",X"27",X"28",X"0D",X"FE",X"33",X"28",X"18",X"DD",X"7E",X"12",X"E6",
		X"FD",X"DD",X"77",X"12",X"C9",X"DD",X"7E",X"12",X"F6",X"02",X"DD",X"77",X"12",X"C9",X"DD",X"36",
		X"15",X"01",X"18",X"DA",X"DD",X"7E",X"15",X"F6",X"02",X"DD",X"77",X"15",X"C3",X"25",X"1D",X"CD",
		X"3E",X"1C",X"DD",X"7E",X"04",X"E6",X"0F",X"FE",X"08",X"28",X"08",X"FE",X"00",X"28",X"04",X"DD",
		X"35",X"04",X"C9",X"CD",X"C5",X"19",X"CD",X"67",X"1C",X"CD",X"AE",X"1C",X"CD",X"F7",X"1C",X"DD",
		X"7E",X"12",X"E6",X"07",X"C2",X"E1",X"19",X"3E",X"08",X"C3",X"29",X"1B",X"DD",X"7E",X"03",X"E6",
		X"0F",X"FE",X"08",X"28",X"08",X"FE",X"00",X"28",X"04",X"DD",X"35",X"03",X"C9",X"CD",X"C5",X"19",
		X"CD",X"AE",X"1C",X"CD",X"CE",X"1B",X"CD",X"67",X"1C",X"DD",X"7E",X"12",X"E6",X"0D",X"C2",X"E1",
		X"19",X"3E",X"02",X"C3",X"29",X"1B",X"DD",X"7E",X"03",X"E6",X"0F",X"FE",X"08",X"28",X"08",X"FE",
		X"00",X"28",X"04",X"DD",X"34",X"03",X"C9",X"CD",X"C5",X"19",X"CD",X"F7",X"1C",X"CD",X"CE",X"1B",
		X"CD",X"67",X"1C",X"DD",X"7E",X"12",X"E6",X"0E",X"C2",X"E1",X"19",X"3E",X"01",X"C3",X"29",X"1B",
		X"3A",X"59",X"41",X"0F",X"DA",X"D4",X"1D",X"0F",X"DA",X"ED",X"1D",X"0F",X"DA",X"06",X"1E",X"0F",
		X"DA",X"1F",X"1E",X"C9",X"DD",X"7E",X"03",X"D6",X"0C",X"57",X"DD",X"5E",X"04",X"CD",X"58",X"1E",
		X"C0",X"DD",X"7E",X"12",X"E6",X"FE",X"CD",X"38",X"1E",X"DD",X"77",X"12",X"C9",X"DD",X"7E",X"03",
		X"C6",X"0C",X"57",X"DD",X"5E",X"04",X"CD",X"58",X"1E",X"C0",X"DD",X"7E",X"12",X"E6",X"FD",X"CD",
		X"38",X"1E",X"DD",X"77",X"12",X"C9",X"DD",X"56",X"03",X"DD",X"7E",X"04",X"D6",X"0C",X"5F",X"CD",
		X"58",X"1E",X"C0",X"DD",X"7E",X"12",X"E6",X"FB",X"CD",X"38",X"1E",X"DD",X"77",X"12",X"C9",X"DD",
		X"56",X"03",X"DD",X"7E",X"04",X"C6",X"0C",X"5F",X"CD",X"58",X"1E",X"C0",X"DD",X"7E",X"12",X"E6",
		X"F7",X"CD",X"38",X"1E",X"DD",X"77",X"12",X"C9",X"DD",X"6E",X"05",X"CB",X"45",X"20",X"0D",X"CB",
		X"4D",X"20",X"0C",X"CB",X"55",X"20",X"0B",X"CB",X"5D",X"20",X"0A",X"C9",X"F6",X"02",X"C9",X"F6",
		X"01",X"C9",X"F6",X"08",X"C9",X"F6",X"04",X"C9",X"DD",X"E5",X"EB",X"DD",X"21",X"E0",X"42",X"06",
		X"06",X"DD",X"7E",X"03",X"BC",X"28",X"09",X"3D",X"BC",X"28",X"05",X"3C",X"3C",X"BC",X"20",X"0F",
		X"DD",X"7E",X"04",X"BD",X"28",X"14",X"3D",X"BD",X"28",X"10",X"3C",X"3C",X"BD",X"28",X"0B",X"11",
		X"20",X"00",X"DD",X"19",X"10",X"DB",X"DD",X"E1",X"EB",X"C9",X"DD",X"7E",X"02",X"FE",X"03",X"C2",
		X"7F",X"1E",X"DD",X"E1",X"EB",X"C9",X"DD",X"21",X"E0",X"42",X"06",X"06",X"DD",X"7E",X"00",X"A7",
		X"28",X"0C",X"DD",X"CB",X"07",X"7E",X"20",X"06",X"DD",X"7E",X"06",X"A7",X"20",X"08",X"11",X"20",
		X"00",X"DD",X"19",X"10",X"E7",X"C9",X"DD",X"7E",X"05",X"E6",X"7F",X"DD",X"77",X"05",X"DD",X"7E",
		X"0D",X"FE",X"02",X"D2",X"AE",X"22",X"DD",X"7E",X"06",X"E6",X"03",X"FE",X"03",X"CA",X"3C",X"22",
		X"DD",X"7E",X"07",X"A7",X"C2",X"81",X"1F",X"DD",X"7E",X"02",X"EF",X"DF",X"1E",X"02",X"1F",X"DD",
		X"36",X"19",X"16",X"DD",X"7E",X"05",X"E6",X"03",X"28",X"0C",X"DD",X"35",X"04",X"DD",X"35",X"04",
		X"DD",X"34",X"02",X"C3",X"AE",X"1E",X"DD",X"34",X"03",X"DD",X"34",X"03",X"DD",X"34",X"02",X"C3",
		X"AE",X"1E",X"3A",X"5F",X"42",X"CB",X"47",X"C2",X"AE",X"1E",X"DD",X"7E",X"05",X"0F",X"30",X"19",
		X"DD",X"35",X"03",X"DD",X"35",X"19",X"20",X"96",X"DD",X"36",X"06",X"00",X"DD",X"34",X"04",X"DD",
		X"34",X"04",X"DD",X"36",X"02",X"00",X"C3",X"AE",X"1E",X"0F",X"30",X"1A",X"DD",X"34",X"03",X"DD",
		X"35",X"19",X"C2",X"AE",X"1E",X"DD",X"36",X"06",X"00",X"DD",X"34",X"04",X"DD",X"34",X"04",X"DD",
		X"36",X"02",X"00",X"C3",X"AE",X"1E",X"0F",X"30",X"1A",X"DD",X"35",X"04",X"DD",X"35",X"19",X"C2",
		X"AE",X"1E",X"DD",X"36",X"06",X"00",X"DD",X"35",X"03",X"DD",X"35",X"03",X"DD",X"36",X"02",X"00",
		X"C3",X"AE",X"1E",X"0F",X"D2",X"AE",X"1E",X"DD",X"34",X"04",X"DD",X"35",X"19",X"C2",X"AE",X"1E",
		X"DD",X"36",X"06",X"00",X"DD",X"35",X"03",X"DD",X"35",X"03",X"DD",X"36",X"02",X"00",X"C3",X"AE",
		X"1E",X"CD",X"87",X"1F",X"C3",X"AE",X"1E",X"DD",X"7E",X"05",X"0F",X"DA",X"25",X"21",X"0F",X"DA",
		X"BF",X"21",X"0F",X"DA",X"9B",X"20",X"16",X"8C",X"1E",X"8D",X"0E",X"8F",X"DD",X"7E",X"02",X"EF",
		X"BE",X"1F",X"C9",X"1F",X"E6",X"1F",X"00",X"20",X"6F",X"20",X"DD",X"73",X"1D",X"DD",X"71",X"1E",
		X"DD",X"7E",X"18",X"DD",X"72",X"18",X"DD",X"36",X"1B",X"00",X"DD",X"77",X"1C",X"C9",X"DD",X"36",
		X"0A",X"80",X"CD",X"AA",X"1F",X"DD",X"34",X"02",X"C9",X"3A",X"5F",X"42",X"CB",X"47",X"C0",X"DD",
		X"34",X"04",X"DD",X"7E",X"04",X"E6",X"0F",X"FE",X"00",X"28",X"03",X"FE",X"08",X"C0",X"DD",X"36",
		X"19",X"08",X"DD",X"34",X"02",X"C9",X"DD",X"35",X"19",X"C0",X"DD",X"36",X"19",X"30",X"DD",X"7E",
		X"04",X"C6",X"04",X"DD",X"77",X"04",X"DD",X"7E",X"1D",X"DD",X"77",X"18",X"DD",X"34",X"02",X"C9",
		X"DD",X"35",X"19",X"28",X"10",X"DD",X"7E",X"19",X"E6",X"07",X"C0",X"DD",X"7E",X"0A",X"3C",X"E6",
		X"81",X"DD",X"77",X"0A",X"C9",X"CD",X"36",X"20",X"DD",X"7E",X"04",X"C6",X"04",X"DD",X"77",X"04",
		X"DD",X"36",X"1B",X"00",X"DD",X"36",X"0A",X"80",X"DD",X"36",X"19",X"00",X"DD",X"7E",X"1E",X"DD",
		X"77",X"18",X"DD",X"34",X"02",X"C9",X"DD",X"36",X"19",X"30",X"3A",X"0D",X"40",X"A7",X"3A",X"2D",
		X"41",X"20",X"03",X"3A",X"2C",X"41",X"FE",X"7F",X"30",X"1A",X"FE",X"4F",X"30",X"0B",X"DD",X"34",
		X"1B",X"DD",X"7E",X"1B",X"FE",X"04",X"C8",X"E1",X"C9",X"DD",X"34",X"1B",X"DD",X"7E",X"1B",X"FE",
		X"03",X"C8",X"E1",X"C9",X"DD",X"34",X"1B",X"DD",X"7E",X"1B",X"FE",X"02",X"C8",X"E1",X"C9",X"3A",
		X"5F",X"42",X"CB",X"47",X"C0",X"DD",X"34",X"04",X"DD",X"7E",X"04",X"E6",X"0F",X"FE",X"00",X"28",
		X"03",X"FE",X"08",X"C0",X"DD",X"36",X"02",X"00",X"DD",X"36",X"06",X"00",X"DD",X"36",X"0A",X"00",
		X"DD",X"7E",X"1C",X"DD",X"77",X"18",X"DD",X"36",X"19",X"00",X"C9",X"16",X"0C",X"1E",X"0D",X"0E",
		X"0F",X"DD",X"7E",X"02",X"EF",X"BE",X"1F",X"AF",X"20",X"BB",X"20",X"D5",X"20",X"0C",X"21",X"3A",
		X"5F",X"42",X"CB",X"47",X"C0",X"DD",X"35",X"04",X"C3",X"D2",X"1F",X"DD",X"35",X"19",X"C0",X"DD",
		X"36",X"19",X"60",X"DD",X"7E",X"04",X"D6",X"04",X"DD",X"77",X"04",X"DD",X"7E",X"1D",X"DD",X"77",
		X"18",X"DD",X"34",X"02",X"C9",X"DD",X"35",X"19",X"CA",X"EB",X"20",X"DD",X"7E",X"19",X"E6",X"07",
		X"C0",X"DD",X"7E",X"0A",X"3C",X"E6",X"81",X"DD",X"77",X"0A",X"C9",X"CD",X"36",X"20",X"DD",X"7E",
		X"04",X"D6",X"04",X"DD",X"77",X"04",X"DD",X"36",X"1B",X"00",X"DD",X"36",X"0A",X"80",X"DD",X"36",
		X"19",X"00",X"DD",X"7E",X"1E",X"DD",X"77",X"18",X"DD",X"34",X"02",X"C9",X"3A",X"5F",X"42",X"CB",
		X"47",X"C0",X"DD",X"35",X"04",X"DD",X"7E",X"04",X"E6",X"0F",X"FE",X"00",X"CA",X"84",X"20",X"FE",
		X"08",X"C0",X"C3",X"84",X"20",X"16",X"10",X"1E",X"11",X"0E",X"13",X"DD",X"7E",X"02",X"EF",X"BE",
		X"1F",X"39",X"21",X"56",X"21",X"70",X"21",X"A6",X"21",X"3A",X"5F",X"42",X"CB",X"47",X"C0",X"DD",
		X"35",X"03",X"DD",X"7E",X"03",X"E6",X"0F",X"FE",X"00",X"28",X"03",X"FE",X"08",X"C0",X"DD",X"36",
		X"19",X"08",X"DD",X"34",X"02",X"C9",X"DD",X"35",X"19",X"C0",X"DD",X"36",X"19",X"60",X"DD",X"7E",
		X"03",X"D6",X"04",X"DD",X"77",X"03",X"DD",X"7E",X"1D",X"DD",X"77",X"18",X"DD",X"34",X"02",X"C9",
		X"DD",X"35",X"19",X"28",X"10",X"DD",X"7E",X"19",X"E6",X"07",X"C0",X"DD",X"7E",X"0A",X"3C",X"E6",
		X"81",X"DD",X"77",X"0A",X"C9",X"CD",X"36",X"20",X"DD",X"7E",X"03",X"D6",X"04",X"DD",X"77",X"03",
		X"DD",X"36",X"1B",X"00",X"DD",X"36",X"0A",X"80",X"DD",X"36",X"19",X"00",X"DD",X"7E",X"1E",X"DD",
		X"77",X"18",X"DD",X"34",X"02",X"C9",X"3A",X"5F",X"42",X"CB",X"47",X"C0",X"DD",X"35",X"03",X"DD",
		X"7E",X"03",X"E6",X"0F",X"FE",X"00",X"CA",X"84",X"20",X"FE",X"08",X"C0",X"C3",X"84",X"20",X"16",
		X"13",X"1E",X"11",X"0E",X"13",X"DD",X"7E",X"02",X"EF",X"BE",X"1F",X"D3",X"21",X"DF",X"21",X"F9",
		X"21",X"23",X"22",X"3A",X"5F",X"42",X"CB",X"47",X"C0",X"DD",X"34",X"03",X"C3",X"42",X"21",X"DD",
		X"35",X"19",X"C0",X"DD",X"36",X"19",X"60",X"DD",X"7E",X"03",X"C6",X"04",X"DD",X"77",X"03",X"DD",
		X"7E",X"1D",X"DD",X"77",X"18",X"DD",X"34",X"02",X"C9",X"DD",X"35",X"19",X"CA",X"02",X"22",X"C3",
		X"75",X"21",X"CD",X"36",X"20",X"DD",X"7E",X"03",X"C6",X"04",X"DD",X"77",X"03",X"DD",X"36",X"1B",
		X"00",X"DD",X"36",X"0A",X"80",X"DD",X"36",X"19",X"00",X"DD",X"7E",X"1E",X"DD",X"77",X"18",X"DD",
		X"34",X"02",X"C9",X"3A",X"5F",X"42",X"CB",X"47",X"C0",X"DD",X"34",X"03",X"DD",X"7E",X"03",X"E6",
		X"0F",X"FE",X"00",X"CA",X"84",X"20",X"FE",X"08",X"C0",X"C3",X"84",X"20",X"DD",X"7E",X"07",X"A7",
		X"28",X"36",X"CD",X"48",X"22",X"C3",X"AE",X"1E",X"DD",X"7E",X"05",X"0F",X"38",X"18",X"0F",X"38",
		X"1E",X"0F",X"38",X"09",X"16",X"94",X"1E",X"95",X"0E",X"97",X"C3",X"9C",X"1F",X"16",X"14",X"1E",
		X"15",X"0E",X"17",X"C3",X"A1",X"20",X"16",X"18",X"1E",X"19",X"0E",X"1B",X"C3",X"2B",X"21",X"16",
		X"1B",X"1E",X"19",X"0E",X"18",X"C3",X"C5",X"21",X"CD",X"7E",X"22",X"C3",X"AE",X"1E",X"DD",X"7E",
		X"05",X"0F",X"38",X"18",X"0F",X"38",X"1E",X"0F",X"38",X"09",X"16",X"9C",X"1E",X"9D",X"0E",X"9F",
		X"C3",X"9C",X"1F",X"16",X"1C",X"1E",X"1D",X"0E",X"1F",X"C3",X"A1",X"20",X"16",X"20",X"1E",X"21",
		X"0E",X"23",X"C3",X"2B",X"21",X"16",X"23",X"1E",X"21",X"0E",X"20",X"C3",X"C5",X"21",X"DD",X"7E",
		X"07",X"A7",X"28",X"25",X"3D",X"28",X"13",X"DD",X"7E",X"06",X"E6",X"03",X"20",X"06",X"CD",X"48",
		X"22",X"C3",X"AE",X"1E",X"CD",X"87",X"1F",X"C3",X"AE",X"1E",X"DD",X"7E",X"06",X"E6",X"03",X"FE",
		X"03",X"20",X"0D",X"CD",X"7E",X"22",X"C3",X"AE",X"1E",X"DD",X"36",X"06",X"00",X"C3",X"AE",X"1E",
		X"C3",X"D7",X"1E",X"C9",X"00",X"DD",X"21",X"A0",X"42",X"DD",X"7E",X"00",X"A7",X"C8",X"AF",X"32",
		X"61",X"41",X"3A",X"0F",X"40",X"A7",X"C2",X"2F",X"23",X"3A",X"10",X"40",X"47",X"E6",X"80",X"4F",
		X"78",X"E6",X"20",X"07",X"B1",X"4F",X"78",X"E6",X"04",X"07",X"07",X"07",X"B1",X"4F",X"78",X"E6",
		X"08",X"07",X"B1",X"4F",X"A7",X"C8",X"06",X"80",X"07",X"DA",X"56",X"23",X"06",X"40",X"07",X"DA",
		X"56",X"23",X"06",X"20",X"07",X"DA",X"9D",X"23",X"06",X"10",X"07",X"DA",X"9D",X"23",X"C9",X"3A",
		X"0D",X"40",X"A7",X"CA",X"F9",X"22",X"3A",X"10",X"40",X"E6",X"40",X"07",X"4F",X"3A",X"11",X"40",
		X"47",X"E6",X"20",X"07",X"B1",X"4F",X"78",X"E6",X"08",X"07",X"B1",X"4F",X"78",X"E6",X"04",X"07",
		X"07",X"07",X"B1",X"C3",X"13",X"23",X"78",X"32",X"60",X"41",X"CD",X"EA",X"23",X"3A",X"61",X"41",
		X"A7",X"CA",X"D4",X"23",X"3A",X"62",X"41",X"5F",X"E6",X"A0",X"20",X"0B",X"AF",X"32",X"BE",X"41",
		X"3A",X"60",X"41",X"32",X"62",X"41",X"C9",X"3A",X"60",X"41",X"BB",X"20",X"12",X"3A",X"BE",X"41",
		X"A7",X"C8",X"3D",X"32",X"BE",X"41",X"20",X"01",X"C9",X"CB",X"47",X"C2",X"E4",X"22",X"C9",X"3A",
		X"60",X"41",X"32",X"62",X"41",X"3E",X"08",X"32",X"BE",X"41",X"C3",X"E4",X"22",X"78",X"32",X"60",
		X"41",X"CD",X"A5",X"25",X"3A",X"61",X"41",X"A7",X"CA",X"D4",X"23",X"3A",X"62",X"41",X"5F",X"E6",
		X"30",X"20",X"0B",X"AF",X"32",X"BE",X"41",X"3A",X"60",X"41",X"32",X"62",X"41",X"C9",X"3A",X"60",
		X"41",X"BB",X"C2",X"8F",X"23",X"3A",X"BE",X"41",X"A7",X"C8",X"3D",X"32",X"BE",X"41",X"20",X"B9",
		X"32",X"BE",X"41",X"C9",X"AF",X"32",X"BE",X"41",X"3A",X"62",X"41",X"A7",X"C8",X"4F",X"E6",X"30",
		X"C2",X"A5",X"25",X"79",X"E6",X"C0",X"C2",X"EA",X"23",X"C9",X"DD",X"7E",X"04",X"E6",X"07",X"FE",
		X"02",X"CA",X"21",X"24",X"CD",X"0E",X"24",X"C0",X"DD",X"7E",X"04",X"E6",X"07",X"FE",X"02",X"D2",
		X"08",X"24",X"3E",X"10",X"32",X"62",X"41",X"C9",X"3E",X"20",X"32",X"62",X"41",X"C9",X"CB",X"79",
		X"C2",X"1A",X"24",X"11",X"02",X"00",X"CD",X"43",X"24",X"C9",X"11",X"FF",X"FF",X"CD",X"43",X"24",
		X"C9",X"CB",X"79",X"C2",X"99",X"24",X"DD",X"7E",X"03",X"E6",X"07",X"FE",X"02",X"CA",X"38",X"24",
		X"FE",X"04",X"D2",X"04",X"25",X"C3",X"AB",X"24",X"11",X"02",X"00",X"CD",X"89",X"25",X"C0",X"CD",
		X"F1",X"24",X"C9",X"DD",X"66",X"10",X"DD",X"6E",X"11",X"19",X"7E",X"CD",X"87",X"27",X"28",X"09",
		X"FE",X"34",X"28",X"05",X"FE",X"33",X"C2",X"7A",X"24",X"11",X"E0",X"FF",X"19",X"7E",X"CD",X"87",
		X"27",X"C8",X"FE",X"33",X"C8",X"11",X"40",X"00",X"19",X"7E",X"CD",X"87",X"27",X"28",X"03",X"FE",
		X"34",X"C0",X"3E",X"20",X"32",X"62",X"41",X"E1",X"E1",X"C9",X"11",X"E0",X"FF",X"19",X"7E",X"CD",
		X"87",X"27",X"28",X"03",X"FE",X"34",X"C0",X"19",X"7E",X"CD",X"87",X"27",X"28",X"03",X"FE",X"33",
		X"C0",X"3E",X"10",X"32",X"62",X"41",X"E1",X"E1",X"C9",X"DD",X"7E",X"03",X"E6",X"07",X"FE",X"02",
		X"CA",X"7E",X"25",X"FE",X"04",X"D2",X"04",X"25",X"C3",X"AB",X"24",X"DD",X"66",X"10",X"DD",X"6E",
		X"11",X"7E",X"FE",X"34",X"CA",X"4E",X"25",X"CD",X"87",X"27",X"C0",X"11",X"E0",X"FF",X"19",X"7E",
		X"FE",X"33",X"CA",X"74",X"25",X"CD",X"87",X"27",X"C0",X"23",X"7E",X"FE",X"33",X"20",X"0D",X"11",
		X"20",X"00",X"19",X"7E",X"FE",X"34",X"CA",X"6A",X"25",X"C3",X"7C",X"25",X"CD",X"87",X"27",X"C0",
		X"11",X"20",X"00",X"19",X"7E",X"CD",X"87",X"27",X"C0",X"DD",X"36",X"18",X"30",X"CD",X"F1",X"24",
		X"C9",X"00",X"3E",X"01",X"32",X"61",X"41",X"DD",X"34",X"03",X"CB",X"71",X"C0",X"DD",X"35",X"03",
		X"DD",X"35",X"03",X"C9",X"DD",X"66",X"10",X"DD",X"6E",X"11",X"7E",X"FE",X"34",X"28",X"3F",X"CD",
		X"87",X"27",X"C0",X"11",X"E0",X"FF",X"19",X"7E",X"FE",X"33",X"28",X"27",X"CD",X"87",X"27",X"C0",
		X"11",X"20",X"00",X"19",X"23",X"7E",X"FE",X"34",X"28",X"40",X"CD",X"87",X"27",X"C0",X"11",X"E0",
		X"FF",X"19",X"7E",X"FE",X"33",X"28",X"45",X"CD",X"87",X"27",X"C0",X"DD",X"36",X"18",X"30",X"CD",
		X"F1",X"24",X"C9",X"11",X"20",X"00",X"19",X"7E",X"FE",X"34",X"28",X"02",X"18",X"26",X"DD",X"36",
		X"18",X"2C",X"DD",X"36",X"09",X"2C",X"DD",X"7E",X"04",X"E6",X"F8",X"C6",X"02",X"DD",X"77",X"04",
		X"3A",X"5F",X"42",X"E6",X"03",X"C0",X"CD",X"F1",X"24",X"C9",X"DD",X"36",X"18",X"2D",X"DD",X"36",
		X"09",X"2D",X"18",X"E2",X"CD",X"F1",X"24",X"DD",X"36",X"18",X"30",X"C9",X"18",X"F6",X"11",X"FF",
		X"FF",X"CD",X"89",X"25",X"C0",X"CD",X"F1",X"24",X"C9",X"DD",X"66",X"10",X"DD",X"6E",X"11",X"19",
		X"7E",X"CD",X"87",X"27",X"28",X"03",X"FE",X"34",X"C0",X"11",X"E0",X"FF",X"19",X"7E",X"CD",X"87",
		X"27",X"C8",X"FE",X"33",X"C9",X"DD",X"7E",X"03",X"E6",X"07",X"FE",X"02",X"CA",X"DC",X"25",X"CD",
		X"C9",X"25",X"C0",X"DD",X"7E",X"03",X"E6",X"07",X"FE",X"02",X"D2",X"C3",X"25",X"3E",X"40",X"32",
		X"62",X"41",X"C9",X"3E",X"80",X"32",X"62",X"41",X"C9",X"CB",X"69",X"CA",X"D5",X"25",X"11",X"20",
		X"00",X"CD",X"F6",X"26",X"C9",X"11",X"C0",X"FF",X"CD",X"F6",X"26",X"C9",X"CB",X"69",X"CA",X"12",
		X"26",X"00",X"DD",X"7E",X"04",X"FE",X"19",X"30",X"17",X"DD",X"7E",X"03",X"FE",X"50",X"38",X"03",
		X"FE",X"5F",X"D8",X"DD",X"7E",X"04",X"FE",X"03",X"D2",X"00",X"26",X"DD",X"36",X"04",X"F3",X"C9",
		X"DD",X"7E",X"04",X"E6",X"07",X"FE",X"02",X"CA",X"C7",X"26",X"FE",X"04",X"D2",X"44",X"27",X"C3",
		X"42",X"26",X"DD",X"7E",X"04",X"FE",X"DC",X"38",X"17",X"DD",X"7E",X"03",X"FE",X"50",X"38",X"03",
		X"FE",X"5F",X"D8",X"DD",X"7E",X"04",X"FE",X"F2",X"DA",X"30",X"26",X"DD",X"36",X"04",X"01",X"C9",
		X"DD",X"7E",X"04",X"E6",X"07",X"FE",X"02",X"CA",X"D2",X"26",X"FE",X"04",X"D2",X"44",X"27",X"C3",
		X"42",X"26",X"DD",X"66",X"10",X"DD",X"6E",X"11",X"7E",X"FE",X"31",X"28",X"4C",X"CD",X"87",X"27",
		X"C0",X"23",X"7E",X"CD",X"87",X"27",X"C0",X"11",X"DF",X"FF",X"19",X"7E",X"FE",X"31",X"CA",X"A2",
		X"26",X"CD",X"87",X"27",X"C0",X"23",X"7E",X"CD",X"87",X"27",X"C0",X"CD",X"AB",X"26",X"DD",X"36",
		X"18",X"30",X"C9",X"DD",X"36",X"18",X"2A",X"DD",X"36",X"09",X"2A",X"DD",X"7E",X"03",X"E6",X"F8",
		X"C6",X"02",X"DD",X"77",X"03",X"3A",X"5F",X"42",X"E6",X"03",X"C0",X"CD",X"AB",X"26",X"C9",X"DD",
		X"36",X"18",X"2B",X"DD",X"36",X"09",X"2B",X"18",X"E2",X"23",X"7E",X"FE",X"32",X"28",X"D4",X"C3",
		X"BD",X"26",X"23",X"7E",X"FE",X"32",X"28",X"E7",X"C3",X"C5",X"26",X"3E",X"01",X"32",X"61",X"41",
		X"DD",X"34",X"04",X"CB",X"61",X"C0",X"DD",X"35",X"04",X"DD",X"35",X"04",X"C9",X"CD",X"AB",X"26",
		X"DD",X"36",X"18",X"30",X"C9",X"18",X"F6",X"11",X"20",X"00",X"CD",X"DD",X"26",X"C0",X"CD",X"AB",
		X"26",X"C9",X"11",X"C0",X"FF",X"CD",X"DD",X"26",X"C0",X"CD",X"AB",X"26",X"C9",X"DD",X"66",X"10",
		X"DD",X"6E",X"11",X"19",X"7E",X"FE",X"31",X"28",X"04",X"CD",X"87",X"27",X"C0",X"23",X"7E",X"CD",
		X"87",X"27",X"C8",X"FE",X"32",X"C9",X"DD",X"66",X"10",X"DD",X"6E",X"11",X"19",X"7E",X"CD",X"87",
		X"27",X"28",X"09",X"FE",X"31",X"28",X"05",X"FE",X"32",X"C2",X"28",X"27",X"23",X"7E",X"CD",X"87",
		X"27",X"C8",X"FE",X"32",X"C8",X"2B",X"2B",X"7E",X"CD",X"87",X"27",X"28",X"03",X"FE",X"31",X"C0",
		X"3E",X"80",X"32",X"62",X"41",X"E1",X"E1",X"C9",X"23",X"7E",X"CD",X"87",X"27",X"28",X"03",X"FE",
		X"31",X"C0",X"23",X"7E",X"CD",X"87",X"27",X"28",X"03",X"FE",X"32",X"C0",X"3E",X"40",X"32",X"62",
		X"41",X"E1",X"E1",X"C9",X"DD",X"66",X"10",X"DD",X"6E",X"11",X"7E",X"FE",X"31",X"CA",X"99",X"26",
		X"CD",X"87",X"27",X"C0",X"23",X"7E",X"CD",X"87",X"27",X"C0",X"11",X"DF",X"FF",X"19",X"7E",X"FE",
		X"31",X"CA",X"99",X"26",X"CD",X"87",X"27",X"C0",X"23",X"7E",X"CD",X"87",X"27",X"C0",X"19",X"7E",
		X"FE",X"31",X"CA",X"A2",X"26",X"CD",X"87",X"27",X"C0",X"23",X"7E",X"CD",X"87",X"27",X"C0",X"DD",
		X"36",X"18",X"30",X"CD",X"AB",X"26",X"C9",X"FE",X"10",X"C8",X"FE",X"2F",X"C8",X"FE",X"4C",X"C8",
		X"FE",X"4D",X"C8",X"FE",X"4E",X"C8",X"FE",X"4F",X"C8",X"FE",X"44",X"C8",X"FE",X"45",X"C8",X"FE",
		X"46",X"C8",X"FE",X"47",X"C8",X"FE",X"35",X"C8",X"FE",X"36",X"C8",X"FE",X"37",X"C8",X"FE",X"38",
		X"C8",X"FE",X"48",X"C8",X"FE",X"49",X"C8",X"FE",X"4A",X"C8",X"FE",X"4B",X"C9",X"01",X"00",X"00",
		X"C2",X"7A",X"00",X"00",X"00",X"04",X"30",X"00",X"00",X"00",X"00",X"00",X"01",X"52",X"1B",X"00",
		X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FD",X"21",X"A0",
		X"42",X"FD",X"7E",X"00",X"A7",X"C8",X"FD",X"7E",X"01",X"A7",X"C0",X"DD",X"21",X"E0",X"42",X"06",
		X"06",X"DD",X"7E",X"00",X"A7",X"28",X"57",X"DD",X"7E",X"06",X"A7",X"C2",X"4E",X"28",X"DD",X"7E",
		X"03",X"C6",X"07",X"FD",X"96",X"03",X"38",X"46",X"FE",X"0A",X"30",X"42",X"DD",X"7E",X"04",X"C6",
		X"07",X"FD",X"96",X"04",X"38",X"38",X"FE",X"0A",X"30",X"34",X"FD",X"36",X"02",X"00",X"FD",X"36",
		X"0C",X"0F",X"FD",X"36",X"00",X"00",X"FD",X"36",X"01",X"01",X"FD",X"36",X"18",X"34",X"FD",X"36",
		X"0A",X"00",X"AF",X"21",X"80",X"58",X"C5",X"06",X"80",X"D7",X"C1",X"3E",X"01",X"32",X"80",X"58",
		X"21",X"BC",X"40",X"3A",X"06",X"40",X"A7",X"28",X"03",X"21",X"0A",X"40",X"34",X"C9",X"11",X"20",
		X"00",X"DD",X"19",X"10",X"9C",X"C9",X"CD",X"8D",X"14",X"DD",X"21",X"A0",X"42",X"DD",X"36",X"08",
		X"07",X"DD",X"7E",X"0A",X"DD",X"86",X"18",X"DD",X"77",X"09",X"DD",X"7E",X"03",X"FE",X"10",X"DA",
		X"8A",X"28",X"3A",X"5F",X"42",X"CB",X"47",X"C2",X"7D",X"28",X"DD",X"35",X"03",X"CB",X"67",X"C0",
		X"DD",X"7E",X"0A",X"3C",X"E6",X"03",X"DD",X"77",X"0A",X"C9",X"00",X"AF",X"32",X"80",X"58",X"21",
		X"A0",X"42",X"06",X"00",X"D7",X"3A",X"06",X"40",X"A7",X"20",X"05",X"21",X"BC",X"40",X"34",X"C9",
		X"3A",X"0D",X"40",X"A7",X"C2",X"F8",X"28",X"3A",X"0E",X"41",X"A7",X"CA",X"14",X"29",X"3D",X"32",
		X"0E",X"41",X"CD",X"ED",X"28",X"3A",X"0E",X"40",X"A7",X"28",X"2C",X"3A",X"21",X"42",X"A7",X"20",
		X"26",X"21",X"0D",X"40",X"36",X"01",X"21",X"00",X"42",X"11",X"10",X"42",X"01",X"06",X"00",X"ED",
		X"B0",X"21",X"0B",X"41",X"11",X"00",X"42",X"01",X"06",X"00",X"ED",X"B0",X"21",X"10",X"42",X"11",
		X"0B",X"41",X"01",X"06",X"00",X"ED",X"B0",X"21",X"0A",X"40",X"36",X"01",X"C9",X"3A",X"0A",X"41",
		X"21",X"0B",X"41",X"86",X"32",X"0B",X"41",X"C9",X"3A",X"0E",X"41",X"A7",X"CA",X"21",X"29",X"3D",
		X"32",X"0E",X"41",X"CD",X"ED",X"28",X"3A",X"20",X"42",X"A7",X"20",X"DB",X"21",X"0D",X"40",X"36",
		X"00",X"C3",X"C6",X"28",X"21",X"20",X"42",X"36",X"01",X"21",X"0A",X"40",X"34",X"CD",X"2E",X"29",
		X"C9",X"21",X"21",X"42",X"36",X"01",X"21",X"0A",X"40",X"34",X"CD",X"2E",X"29",X"C9",X"21",X"02",
		X"50",X"22",X"0B",X"40",X"21",X"08",X"40",X"36",X"20",X"2C",X"36",X"70",X"AF",X"32",X"BF",X"40",
		X"21",X"A0",X"42",X"11",X"A1",X"42",X"36",X"00",X"01",X"FF",X"00",X"ED",X"B0",X"21",X"60",X"40",
		X"11",X"61",X"40",X"01",X"3F",X"00",X"36",X"00",X"ED",X"B0",X"C9",X"2A",X"0B",X"40",X"06",X"1C",
		X"3E",X"10",X"D7",X"11",X"04",X"00",X"19",X"22",X"0B",X"40",X"21",X"08",X"40",X"35",X"C0",X"3E",
		X"01",X"32",X"BF",X"40",X"11",X"02",X"06",X"3A",X"0D",X"40",X"83",X"5F",X"CF",X"11",X"0C",X"06",
		X"CF",X"C9",X"CD",X"C0",X"29",X"21",X"09",X"40",X"35",X"C0",X"11",X"0C",X"07",X"CF",X"21",X"0D",
		X"40",X"7E",X"A7",X"20",X"16",X"3A",X"0E",X"40",X"A7",X"CA",X"BA",X"29",X"3A",X"21",X"42",X"A7",
		X"C2",X"BA",X"29",X"21",X"0D",X"40",X"36",X"01",X"C3",X"C6",X"28",X"3A",X"20",X"42",X"A7",X"C2",
		X"BA",X"29",X"21",X"0D",X"40",X"36",X"00",X"C3",X"C6",X"28",X"3E",X"01",X"32",X"05",X"40",X"C9",
		X"3A",X"BF",X"40",X"A7",X"CC",X"5B",X"29",X"C9",X"FD",X"21",X"A0",X"42",X"FD",X"7E",X"00",X"A7",
		X"C8",X"FD",X"7E",X"01",X"A7",X"C0",X"DD",X"21",X"E0",X"42",X"06",X"06",X"DD",X"7E",X"00",X"A7",
		X"28",X"32",X"DD",X"7E",X"06",X"A7",X"28",X"2C",X"DD",X"7E",X"01",X"A7",X"20",X"26",X"DD",X"7E",
		X"03",X"C6",X"07",X"FD",X"96",X"03",X"38",X"1C",X"FE",X"0A",X"30",X"18",X"DD",X"7E",X"04",X"C6",
		X"07",X"FD",X"96",X"04",X"38",X"0E",X"FE",X"0A",X"30",X"0A",X"DD",X"7E",X"02",X"FE",X"03",X"28",
		X"17",X"C3",X"1A",X"28",X"11",X"20",X"00",X"DD",X"19",X"10",X"C1",X"C9",X"21",X"0A",X"40",X"3A",
		X"06",X"40",X"A7",X"C0",X"21",X"BC",X"40",X"C9",X"3A",X"06",X"40",X"A7",X"28",X"06",X"DD",X"5E",
		X"0D",X"16",X"03",X"CF",X"DD",X"36",X"00",X"00",X"DD",X"36",X"01",X"01",X"DD",X"36",X"02",X"00",
		X"DD",X"36",X"0C",X"08",X"DD",X"36",X"18",X"38",X"DD",X"36",X"0A",X"00",X"3E",X"04",X"32",X"C0",
		X"58",X"3A",X"5B",X"41",X"A7",X"C2",X"14",X"2A",X"ED",X"5F",X"E6",X"03",X"32",X"5E",X"41",X"3E",
		X"01",X"32",X"5B",X"41",X"3A",X"B0",X"58",X"F6",X"20",X"32",X"B0",X"58",X"3E",X"05",X"32",X"A8",
		X"42",X"C3",X"14",X"2A",X"DD",X"21",X"E0",X"42",X"06",X"06",X"DD",X"7E",X"01",X"A7",X"28",X"2D",
		X"DD",X"7E",X"18",X"DD",X"86",X"0A",X"DD",X"77",X"09",X"DD",X"7E",X"0C",X"E6",X"07",X"FE",X"04",
		X"C2",X"96",X"2A",X"DD",X"34",X"08",X"DD",X"35",X"0C",X"C2",X"AD",X"2A",X"DD",X"36",X"0C",X"08",
		X"DD",X"34",X"02",X"DD",X"7E",X"02",X"FE",X"04",X"28",X"0B",X"DD",X"34",X"0A",X"11",X"20",X"00",
		X"DD",X"19",X"10",X"C6",X"C9",X"DD",X"36",X"00",X"00",X"DD",X"36",X"01",X"00",X"DD",X"36",X"02",
		X"00",X"DD",X"36",X"03",X"00",X"DD",X"36",X"04",X"00",X"C3",X"AD",X"2A",X"3E",X"01",X"32",X"06",
		X"68",X"32",X"07",X"68",X"00",X"3A",X"05",X"40",X"FE",X"03",X"28",X"0D",X"AF",X"32",X"A0",X"58",
		X"32",X"B0",X"58",X"32",X"80",X"58",X"32",X"C0",X"58",X"21",X"C5",X"2D",X"DD",X"21",X"90",X"58",
		X"FD",X"21",X"F1",X"58",X"CD",X"F9",X"2B",X"21",X"03",X"2D",X"DD",X"21",X"A0",X"58",X"FD",X"21",
		X"F2",X"58",X"CD",X"88",X"2B",X"21",X"0D",X"2D",X"DD",X"21",X"B0",X"58",X"FD",X"21",X"F3",X"58",
		X"CD",X"88",X"2B",X"21",X"50",X"2F",X"DD",X"21",X"C0",X"58",X"FD",X"21",X"F4",X"58",X"CD",X"F9",
		X"2B",X"21",X"68",X"2F",X"DD",X"21",X"80",X"58",X"FD",X"21",X"F0",X"58",X"CD",X"F9",X"2B",X"06",
		X"00",X"21",X"F3",X"58",X"CD",X"63",X"2B",X"21",X"F2",X"58",X"CD",X"63",X"2B",X"21",X"F4",X"58",
		X"CD",X"63",X"2B",X"21",X"F0",X"58",X"CD",X"63",X"2B",X"21",X"F1",X"58",X"CD",X"63",X"2B",X"CB",
		X"40",X"20",X"09",X"3E",X"FF",X"32",X"FA",X"58",X"32",X"00",X"78",X"C9",X"3A",X"FA",X"58",X"32",
		X"00",X"78",X"C9",X"7E",X"A7",X"C8",X"CB",X"C0",X"32",X"FA",X"58",X"C9",X"85",X"6F",X"3E",X"00",
		X"8C",X"67",X"7E",X"C9",X"78",X"87",X"CD",X"6C",X"2B",X"5F",X"23",X"56",X"EB",X"C9",X"E1",X"87",
		X"CD",X"6C",X"2B",X"5F",X"23",X"56",X"EB",X"E9",X"DD",X"7E",X"00",X"A7",X"CA",X"FF",X"2B",X"4F",
		X"06",X"08",X"1E",X"80",X"7B",X"A1",X"20",X"05",X"CB",X"3B",X"10",X"F8",X"C9",X"DD",X"7E",X"02",
		X"A3",X"20",X"09",X"DD",X"73",X"02",X"05",X"CD",X"74",X"2B",X"18",X"0C",X"DD",X"35",X"0C",X"C2",
		X"F2",X"2B",X"DD",X"6E",X"06",X"DD",X"66",X"07",X"7E",X"23",X"DD",X"75",X"06",X"DD",X"74",X"07",
		X"FE",X"F0",X"38",X"13",X"21",X"B2",X"2B",X"E5",X"E6",X"0F",X"CA",X"F3",X"2C",X"AF",X"FD",X"77",
		X"00",X"DD",X"77",X"00",X"C3",X"FF",X"2B",X"47",X"07",X"07",X"07",X"E6",X"07",X"21",X"A3",X"2D",
		X"CD",X"6C",X"2B",X"DD",X"77",X"0C",X"78",X"E6",X"1F",X"21",X"AB",X"2D",X"CD",X"6C",X"2B",X"DD",
		X"77",X"0E",X"DD",X"7E",X"0E",X"FD",X"77",X"00",X"C9",X"DD",X"7E",X"00",X"A7",X"20",X"23",X"DD",
		X"7E",X"02",X"A7",X"3E",X"00",X"FD",X"77",X"00",X"C8",X"DD",X"36",X"00",X"00",X"DD",X"36",X"02",
		X"00",X"DD",X"36",X"0D",X"00",X"DD",X"36",X"0E",X"FF",X"DD",X"36",X"0F",X"00",X"FD",X"36",X"00",
		X"00",X"C9",X"4F",X"06",X"08",X"1E",X"80",X"7B",X"A1",X"20",X"05",X"CB",X"3B",X"10",X"F8",X"C9",
		X"DD",X"7E",X"02",X"A3",X"20",X"3F",X"DD",X"73",X"02",X"05",X"78",X"07",X"07",X"07",X"4F",X"06",
		X"00",X"E5",X"09",X"DD",X"E5",X"D1",X"13",X"13",X"13",X"01",X"08",X"00",X"ED",X"B0",X"E1",X"DD",
		X"7E",X"06",X"E6",X"7F",X"DD",X"77",X"0C",X"DD",X"7E",X"04",X"DD",X"77",X"0E",X"DD",X"7E",X"09",
		X"47",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"DD",X"77",X"0B",X"E6",X"08",X"20",X"07",X"DD",X"70",
		X"0F",X"DD",X"36",X"0D",X"00",X"DD",X"35",X"0C",X"20",X"5A",X"DD",X"7E",X"08",X"A7",X"28",X"10",
		X"DD",X"35",X"08",X"20",X"0B",X"7B",X"2F",X"DD",X"A6",X"00",X"DD",X"77",X"00",X"C3",X"F9",X"2B",
		X"DD",X"7E",X"06",X"E6",X"7F",X"DD",X"77",X"0C",X"DD",X"CB",X"06",X"7E",X"28",X"16",X"DD",X"7E",
		X"05",X"ED",X"44",X"DD",X"77",X"05",X"DD",X"CB",X"00",X"46",X"DD",X"CB",X"0D",X"C6",X"28",X"24",
		X"DD",X"CB",X"0D",X"86",X"DD",X"7E",X"04",X"DD",X"86",X"07",X"DD",X"77",X"04",X"DD",X"77",X"0E",
		X"DD",X"7E",X"09",X"DD",X"86",X"0A",X"DD",X"77",X"09",X"47",X"DD",X"7E",X"0B",X"E6",X"08",X"20",
		X"03",X"DD",X"70",X"0F",X"DD",X"7E",X"0E",X"DD",X"86",X"05",X"DD",X"77",X"0E",X"6F",X"26",X"00",
		X"DD",X"7E",X"03",X"E6",X"70",X"28",X"08",X"0F",X"0F",X"0F",X"0F",X"47",X"29",X"10",X"FD",X"FD",
		X"75",X"00",X"C9",X"DD",X"6E",X"06",X"DD",X"66",X"07",X"7E",X"DD",X"77",X"06",X"23",X"7E",X"DD",
		X"77",X"07",X"C9",X"24",X"2E",X"D5",X"2D",X"05",X"2E",X"D5",X"2D",X"05",X"2E",X"52",X"2E",X"02",
		X"2F",X"02",X"2F",X"4A",X"2D",X"38",X"2E",X"19",X"2D",X"6A",X"6B",X"6A",X"6B",X"64",X"62",X"64",
		X"62",X"6A",X"6B",X"6A",X"6B",X"64",X"62",X"64",X"62",X"6A",X"6B",X"6A",X"6B",X"70",X"6E",X"6B",
		X"67",X"64",X"47",X"4B",X"70",X"6E",X"64",X"47",X"4B",X"70",X"6E",X"73",X"00",X"73",X"60",X"67",
		X"6B",X"6E",X"70",X"6E",X"73",X"00",X"73",X"F0",X"19",X"2D",X"6B",X"6E",X"6B",X"6E",X"70",X"6E",
		X"6B",X"49",X"47",X"64",X"67",X"69",X"67",X"6A",X"6B",X"8B",X"6B",X"6E",X"6B",X"6E",X"70",X"6E",
		X"6B",X"49",X"47",X"64",X"67",X"69",X"67",X"6A",X"89",X"67",X"6B",X"6E",X"70",X"6E",X"73",X"70",
		X"6E",X"6B",X"69",X"62",X"64",X"66",X"A7",X"6B",X"6E",X"00",X"6E",X"00",X"6E",X"6B",X"49",X"47",
		X"6B",X"49",X"47",X"73",X"73",X"70",X"8E",X"75",X"87",X"70",X"5E",X"70",X"5E",X"70",X"73",X"00",
		X"73",X"70",X"6E",X"70",X"6B",X"6E",X"69",X"6B",X"6C",X"6E",X"6B",X"89",X"62",X"64",X"66",X"67",
		X"F0",X"4A",X"2D",X"01",X"03",X"05",X"0A",X"14",X"28",X"50",X"00",X"FF",X"03",X"11",X"1F",X"2B",
		X"37",X"42",X"4D",X"57",X"60",X"69",X"72",X"7A",X"81",X"88",X"8F",X"95",X"9B",X"A1",X"A6",X"AB",
		X"B0",X"B5",X"B9",X"BD",X"C1",X"40",X"20",X"F4",X"87",X"00",X"0A",X"FF",X"FF",X"40",X"20",X"FF",
		X"90",X"00",X"01",X"FF",X"FF",X"A0",X"6E",X"73",X"6E",X"73",X"00",X"73",X"69",X"00",X"49",X"00",
		X"49",X"6B",X"6E",X"73",X"00",X"53",X"00",X"53",X"75",X"00",X"55",X"00",X"55",X"B7",X"6E",X"73",
		X"6E",X"73",X"00",X"53",X"00",X"53",X"75",X"00",X"55",X"00",X"55",X"77",X"6E",X"72",X"57",X"55",
		X"6E",X"50",X"52",X"73",X"FF",X"A0",X"8B",X"66",X"00",X"66",X"68",X"00",X"68",X"66",X"00",X"66",
		X"8B",X"66",X"00",X"66",X"8F",X"8D",X"8B",X"66",X"00",X"66",X"6F",X"6D",X"8B",X"6D",X"4A",X"48",
		X"66",X"6A",X"AB",X"FF",X"6E",X"50",X"52",X"93",X"52",X"50",X"6E",X"50",X"52",X"93",X"6E",X"50",
		X"52",X"93",X"52",X"50",X"6E",X"77",X"93",X"FF",X"6B",X"69",X"6B",X"69",X"6B",X"62",X"64",X"67",
		X"6B",X"69",X"6B",X"69",X"8B",X"8E",X"6B",X"69",X"6B",X"69",X"6B",X"62",X"64",X"67",X"6A",X"69",
		X"67",X"FF",X"6B",X"6E",X"6B",X"6E",X"8B",X"87",X"89",X"8B",X"8C",X"00",X"6C",X"6B",X"6C",X"6B",
		X"A9",X"80",X"82",X"86",X"89",X"6C",X"6B",X"6C",X"6B",X"8C",X"70",X"6E",X"6C",X"6B",X"6C",X"69",
		X"6B",X"6E",X"70",X"6E",X"70",X"6E",X"87",X"8B",X"8E",X"73",X"67",X"73",X"67",X"93",X"97",X"95",
		X"93",X"72",X"00",X"72",X"70",X"6E",X"6C",X"69",X"67",X"00",X"67",X"60",X"62",X"64",X"66",X"87",
		X"49",X"4B",X"4C",X"4E",X"50",X"52",X"53",X"55",X"87",X"49",X"4B",X"4C",X"4E",X"50",X"52",X"53",
		X"55",X"67",X"6E",X"6B",X"69",X"67",X"6B",X"69",X"00",X"69",X"60",X"67",X"69",X"67",X"92",X"47",
		X"49",X"4B",X"4C",X"4E",X"50",X"52",X"47",X"92",X"47",X"49",X"4B",X"4C",X"4E",X"50",X"52",X"47",
		X"72",X"70",X"6E",X"6C",X"6B",X"72",X"67",X"62",X"70",X"72",X"67",X"69",X"6B",X"6E",X"73",X"6B",
		X"6E",X"73",X"6B",X"6E",X"73",X"6B",X"6E",X"73",X"92",X"00",X"92",X"00",X"92",X"69",X"6C",X"72",
		X"6B",X"6C",X"70",X"8E",X"8B",X"00",X"8B",X"00",X"8B",X"8F",X"92",X"73",X"72",X"73",X"72",X"70",
		X"6E",X"6C",X"69",X"6B",X"6C",X"72",X"70",X"6E",X"66",X"69",X"6C",X"6B",X"69",X"A7",X"80",X"F0",
		X"52",X"2E",X"A0",X"8E",X"70",X"6E",X"93",X"00",X"93",X"8E",X"70",X"6E",X"95",X"00",X"95",X"8E",
		X"73",X"75",X"77",X"75",X"73",X"72",X"93",X"90",X"AE",X"00",X"8E",X"70",X"6E",X"93",X"00",X"93",
		X"8E",X"70",X"6E",X"95",X"92",X"8E",X"73",X"75",X"77",X"75",X"73",X"72",X"93",X"00",X"93",X"00",
		X"B3",X"78",X"75",X"72",X"6E",X"70",X"6E",X"72",X"6E",X"73",X"00",X"93",X"75",X"97",X"6E",X"78",
		X"75",X"78",X"70",X"6E",X"77",X"75",X"73",X"00",X"73",X"00",X"73",X"70",X"B3",X"F0",X"02",X"2F",
		X"40",X"20",X"F4",X"87",X"FE",X"01",X"FF",X"FF",X"20",X"70",X"FB",X"87",X"00",X"02",X"FF",X"FF",
		X"40",X"20",X"FB",X"87",X"00",X"07",X"FF",X"FF",X"88",X"40",X"ED",X"0A",X"03",X"10",X"4E",X"FF",
		X"00",X"00",X"00",X"E4",X"52",X"39",X"3F",X"3F",X"3F",X"FF",X"05",X"51",X"3F",X"10",X"3F",X"3F",
		X"3F",X"10",X"3F",X"10",X"10",X"3F",X"10",X"3F",X"3F",X"3F",X"10",X"3F",X"10",X"10",X"3F",X"FF",
		X"06",X"51",X"3F",X"10",X"10",X"3F",X"10",X"10",X"3F",X"10",X"10",X"3F",X"10",X"3C",X"3C",X"3F",
		X"10",X"3F",X"10",X"10",X"3F",X"FF",X"07",X"51",X"3F",X"10",X"10",X"3F",X"10",X"10",X"3A",X"3B",
		X"39",X"3E",X"10",X"3D",X"3D",X"3F",X"10",X"3A",X"3B",X"10",X"3F",X"FF",X"C8",X"50",X"3F",X"3F",
		X"3F",X"10",X"3F",X"3F",X"3F",X"10",X"10",X"3A",X"3E",X"10",X"10",X"3F",X"3F",X"3F",X"10",X"10",
		X"3A",X"3F",X"3F",X"FF",X"0A",X"51",X"3F",X"10",X"3F",X"10",X"3F",X"3F",X"3F",X"10",X"3F",X"3F",
		X"3F",X"10",X"3F",X"3F",X"3F",X"FF",X"0B",X"51",X"3F",X"3C",X"3F",X"10",X"3C",X"3C",X"3F",X"10",
		X"10",X"3F",X"10",X"10",X"10",X"10",X"3F",X"FF",X"0C",X"51",X"3F",X"3D",X"3F",X"10",X"3F",X"3D",
		X"3D",X"10",X"10",X"3F",X"10",X"10",X"3F",X"3F",X"3F",X"FF",X"0D",X"51",X"3F",X"10",X"3F",X"10",
		X"3F",X"3F",X"3F",X"10",X"3F",X"3F",X"3F",X"10",X"10",X"10",X"3F",X"FF",X"FF",X"02",X"50",X"21",
		X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",
		X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"FF",
		X"03",X"50",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"31",X"10",X"10",
		X"10",X"10",X"10",X"21",X"10",X"10",X"10",X"31",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"FF",X"04",X"50",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"32",X"10",X"10",X"10",X"10",X"10",X"21",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"FF",X"05",X"50",X"21",X"21",X"21",X"10",X"10",X"21",X"21",X"10",
		X"10",X"21",X"21",X"21",X"21",X"21",X"21",X"10",X"10",X"21",X"10",X"10",X"21",X"21",X"21",X"10",
		X"10",X"21",X"21",X"10",X"10",X"21",X"21",X"21",X"FF",X"46",X"50",X"21",X"33",X"10",X"21",X"21",
		X"10",X"10",X"21",X"21",X"10",X"10",X"10",X"21",X"10",X"10",X"21",X"10",X"10",X"21",X"10",X"21",
		X"10",X"10",X"21",X"21",X"33",X"34",X"21",X"FF",X"47",X"50",X"21",X"10",X"10",X"21",X"21",X"10",
		X"10",X"21",X"21",X"21",X"21",X"21",X"21",X"10",X"10",X"21",X"10",X"10",X"21",X"21",X"21",X"10",
		X"10",X"21",X"21",X"10",X"10",X"21",X"FF",X"48",X"50",X"21",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"21",X"FF",X"49",X"50",X"21",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"21",X"FF",X"0A",X"50",X"21",X"21",X"21",X"21",X"21",X"10",X"10",X"21",X"21",
		X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"10",X"10",X"21",X"21",X"21",X"21",X"10",
		X"10",X"21",X"21",X"21",X"21",X"21",X"21",X"FF",X"0B",X"50",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"21",X"21",X"21",X"21",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"21",
		X"10",X"21",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"FF",X"0C",X"50",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"21",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"21",X"10",X"21",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"FF",X"0D",X"50",
		X"21",X"21",X"21",X"21",X"21",X"10",X"10",X"10",X"10",X"10",X"21",X"10",X"10",X"2E",X"2E",X"2E",
		X"2E",X"2E",X"2E",X"10",X"10",X"21",X"10",X"21",X"10",X"10",X"21",X"21",X"21",X"21",X"21",X"21",
		X"FF",X"4E",X"50",X"21",X"10",X"10",X"10",X"10",X"21",X"10",X"10",X"21",X"10",X"10",X"2E",X"10",
		X"10",X"10",X"10",X"2E",X"10",X"10",X"21",X"21",X"21",X"10",X"10",X"21",X"21",X"21",X"21",X"FF",
		X"4F",X"50",X"21",X"10",X"10",X"10",X"10",X"21",X"33",X"34",X"21",X"10",X"10",X"2E",X"10",X"10",
		X"10",X"10",X"2E",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"21",X"FF",X"50",
		X"50",X"21",X"10",X"10",X"21",X"21",X"21",X"10",X"10",X"21",X"10",X"10",X"2E",X"10",X"10",X"10",
		X"10",X"2E",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"21",X"FF",X"51",X"50",
		X"21",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"21",X"10",X"10",X"2E",X"10",X"10",X"10",X"10",
		X"2E",X"21",X"21",X"21",X"21",X"21",X"10",X"10",X"21",X"10",X"10",X"21",X"FF",X"52",X"50",X"21",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"21",X"10",X"10",X"2E",X"2E",X"2E",X"2E",X"2E",X"2E",
		X"21",X"21",X"21",X"21",X"21",X"10",X"10",X"21",X"33",X"10",X"21",X"FF",X"13",X"50",X"21",X"21",
		X"21",X"10",X"10",X"21",X"21",X"21",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"21",X"21",X"10",X"10",X"21",X"10",X"10",X"21",X"21",X"21",X"FF",X"14",
		X"50",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"21",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"FF",X"15",X"50",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"21",X"21",X"21",X"21",X"21",
		X"21",X"21",X"21",X"10",X"10",X"21",X"21",X"21",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"FF",X"16",X"50",X"21",X"21",X"21",X"21",X"21",X"33",X"10",X"21",X"10",
		X"21",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"21",X"21",X"10",X"10",X"10",X"21",X"21",X"21",
		X"21",X"21",X"10",X"10",X"21",X"21",X"21",X"FF",X"57",X"50",X"21",X"10",X"10",X"10",X"10",X"21",
		X"10",X"21",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"21",X"21",X"10",X"10",X"10",X"21",X"10",
		X"10",X"10",X"21",X"10",X"10",X"21",X"FF",X"58",X"50",X"21",X"10",X"10",X"10",X"10",X"21",X"10",
		X"21",X"33",X"10",X"21",X"21",X"21",X"10",X"10",X"21",X"21",X"10",X"10",X"21",X"21",X"10",X"10",
		X"10",X"21",X"10",X"10",X"21",X"FF",X"59",X"50",X"21",X"10",X"10",X"21",X"21",X"21",X"21",X"21",
		X"10",X"10",X"21",X"21",X"21",X"33",X"10",X"21",X"21",X"10",X"10",X"21",X"21",X"10",X"10",X"10",
		X"21",X"33",X"10",X"21",X"FF",X"1A",X"50",X"21",X"21",X"21",X"10",X"10",X"21",X"21",X"21",X"21",
		X"21",X"10",X"10",X"21",X"21",X"21",X"10",X"10",X"21",X"21",X"10",X"10",X"21",X"21",X"21",X"21",
		X"21",X"21",X"10",X"10",X"21",X"21",X"21",X"FF",X"1B",X"50",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"31",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"FF",X"1C",X"50",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"FF",X"1D",X"50",
		X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",
		X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",
		X"FF",X"FF",X"71",X"6B",X"70",X"6A",X"6F",X"69",X"6E",X"68",X"6D",X"67",X"6C",X"66",X"65",X"60",
		X"62",X"5D",X"64",X"5F",X"63",X"5E",X"62",X"5D",X"61",X"5C",X"5B",X"55",X"5A",X"54",X"59",X"53",
		X"58",X"52",X"57",X"51",X"56",X"50",X"71",X"6B",X"70",X"7D",X"6F",X"69",X"6E",X"68",X"6D",X"7C",
		X"6C",X"66",X"65",X"60",X"62",X"5D",X"64",X"5F",X"63",X"5E",X"62",X"5D",X"61",X"5C",X"7B",X"77",
		X"7A",X"76",X"59",X"75",X"58",X"74",X"79",X"73",X"78",X"72",X"81",X"EC",X"DE",X"EB",X"F0",X"80",
		X"EF",X"EA",X"FE",X"E9",X"ED",X"E8",X"E7",X"E2",X"E6",X"E1",X"E5",X"62",X"62",X"E0",X"E4",X"DF",
		X"E3",X"DE",X"DD",X"96",X"DC",X"96",X"DB",X"D8",X"DA",X"D7",X"D9",X"82",X"84",X"7E",X"81",X"EC",
		X"DE",X"DE",X"0B",X"1A",X"EF",X"0F",X"DE",X"0E",X"DE",X"FF",X"FE",X"FA",X"FD",X"F9",X"E5",X"5D",
		X"5D",X"E0",X"FC",X"F8",X"FB",X"DE",X"F7",X"F3",X"F6",X"F3",X"F5",X"F2",X"F4",X"F1",X"DE",X"82",
		X"84",X"7E",X"C1",X"96",X"96",X"BE",X"C0",X"BD",X"BF",X"BC",X"96",X"BB",X"96",X"BA",X"B9",X"B5",
		X"B8",X"B4",X"AF",X"AF",X"AE",X"AE",X"B7",X"B3",X"B6",X"B2",X"B1",X"81",X"B0",X"81",X"AF",X"AB",
		X"AE",X"AA",X"AD",X"81",X"AC",X"81",X"96",X"D4",X"C1",X"D3",X"D6",X"D2",X"D5",X"D1",X"C1",X"D0",
		X"C1",X"96",X"CF",X"CB",X"CE",X"CA",X"AF",X"AF",X"AE",X"AE",X"CD",X"C9",X"CC",X"C8",X"C7",X"81",
		X"C6",X"81",X"AF",X"C3",X"AE",X"C2",X"C5",X"81",X"C4",X"81",X"02",X"50",X"30",X"30",X"30",X"30",
		X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",
		X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"FF",X"03",X"50",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"31",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"31",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"FF",
		X"04",X"50",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"FF",X"05",X"50",X"30",X"30",X"30",X"10",X"10",X"30",X"30",X"30",X"30",X"30",X"30",
		X"10",X"10",X"30",X"30",X"30",X"30",X"10",X"10",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",
		X"10",X"10",X"30",X"30",X"30",X"FF",X"46",X"50",X"30",X"10",X"10",X"30",X"10",X"10",X"10",X"10",
		X"30",X"10",X"10",X"30",X"30",X"30",X"30",X"10",X"10",X"30",X"30",X"30",X"30",X"30",X"30",X"30",
		X"30",X"33",X"34",X"30",X"FF",X"47",X"50",X"30",X"10",X"10",X"30",X"30",X"30",X"30",X"30",X"30",
		X"10",X"10",X"10",X"10",X"31",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"30",X"FF",X"48",X"50",X"30",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"32",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"30",X"FF",X"49",X"50",X"30",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"30",X"30",X"30",X"30",X"30",X"30",X"10",X"10",X"30",X"30",X"10",X"10",X"30",X"30",X"30",X"30",
		X"30",X"FF",X"0A",X"50",X"30",X"30",X"30",X"30",X"30",X"10",X"10",X"30",X"30",X"30",X"30",X"10",
		X"10",X"30",X"30",X"30",X"30",X"30",X"30",X"10",X"10",X"30",X"30",X"33",X"10",X"30",X"30",X"30",
		X"30",X"30",X"30",X"30",X"FF",X"0B",X"50",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"30",X"10",
		X"10",X"30",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"30",X"30",X"10",X"10",X"10",X"10",X"10",X"FF",X"0C",X"50",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"30",X"10",X"10",X"30",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"30",X"30",X"10",X"10",X"10",X"10",X"10",X"FF",X"0D",X"50",X"30",X"30",X"30",
		X"30",X"30",X"10",X"10",X"30",X"10",X"10",X"30",X"10",X"10",X"2E",X"2E",X"2E",X"2E",X"2E",X"2E",
		X"10",X"10",X"30",X"10",X"10",X"30",X"30",X"30",X"10",X"10",X"30",X"30",X"30",X"FF",X"4E",X"50",
		X"30",X"30",X"30",X"33",X"10",X"30",X"10",X"10",X"30",X"10",X"10",X"2E",X"10",X"10",X"10",X"10",
		X"2E",X"10",X"10",X"30",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"30",X"FF",X"4F",X"50",X"30",
		X"30",X"30",X"10",X"10",X"30",X"30",X"30",X"30",X"10",X"10",X"2E",X"10",X"10",X"10",X"10",X"2E",
		X"10",X"10",X"30",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"30",X"FF",X"50",X"50",X"30",X"30",
		X"30",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"2E",X"10",X"10",X"10",X"10",X"2E",X"10",
		X"10",X"30",X"33",X"10",X"30",X"30",X"30",X"10",X"10",X"30",X"FF",X"51",X"50",X"30",X"30",X"30",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"2E",X"10",X"10",X"10",X"10",X"2E",X"10",X"10",
		X"30",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"30",X"FF",X"52",X"50",X"30",X"30",X"30",X"30",
		X"30",X"10",X"10",X"30",X"30",X"10",X"10",X"2E",X"2E",X"2E",X"2E",X"2E",X"2E",X"10",X"10",X"30",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"30",X"FF",X"13",X"50",X"30",X"30",X"30",X"30",X"30",
		X"30",X"30",X"10",X"10",X"30",X"30",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"30",X"10",X"10",X"30",X"30",X"30",X"10",X"10",X"30",X"30",X"30",X"FF",X"14",X"50",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"30",X"30",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"FF",X"15",
		X"50",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"30",X"30",X"30",X"30",X"30",X"30",
		X"30",X"30",X"30",X"30",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"FF",X"16",X"50",X"30",X"30",X"30",X"10",X"10",X"30",X"30",X"10",X"10",X"30",X"30",X"30",
		X"30",X"30",X"30",X"30",X"10",X"10",X"30",X"33",X"10",X"30",X"30",X"30",X"30",X"30",X"30",X"10",
		X"10",X"30",X"30",X"30",X"FF",X"57",X"50",X"30",X"10",X"10",X"30",X"30",X"10",X"10",X"10",X"31",
		X"10",X"10",X"10",X"10",X"10",X"30",X"30",X"30",X"10",X"10",X"30",X"30",X"30",X"30",X"30",X"30",
		X"10",X"10",X"30",X"FF",X"58",X"50",X"30",X"10",X"10",X"30",X"30",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"30",X"FF",X"59",X"50",X"30",X"33",X"34",X"30",X"30",X"10",X"10",X"30",X"30",X"30",X"30",
		X"30",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"30",X"FF",X"1A",X"50",X"30",X"30",X"30",X"10",X"10",X"30",X"30",X"10",X"10",X"30",X"30",X"30",
		X"30",X"30",X"10",X"10",X"30",X"30",X"30",X"30",X"30",X"30",X"33",X"34",X"30",X"30",X"30",X"10",
		X"10",X"30",X"30",X"30",X"FF",X"1B",X"50",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"31",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"FF",X"1C",X"50",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"FF",X"1D",X"50",X"30",X"30",X"30",
		X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",
		X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"FF",X"FF",X"9B",
		X"95",X"9A",X"94",X"99",X"5D",X"98",X"5D",X"97",X"93",X"96",X"92",X"91",X"8D",X"90",X"62",X"5D",
		X"5D",X"62",X"8C",X"8F",X"8B",X"8E",X"8A",X"89",X"83",X"88",X"82",X"87",X"81",X"86",X"80",X"85",
		X"7F",X"84",X"7E",X"A9",X"A3",X"A8",X"A2",X"A7",X"5D",X"A6",X"5D",X"A5",X"93",X"A4",X"A1",X"91",
		X"8D",X"90",X"62",X"5D",X"5D",X"62",X"8C",X"8F",X"9F",X"A0",X"9E",X"89",X"83",X"88",X"82",X"87",
		X"81",X"9D",X"80",X"9C",X"7F",X"84",X"7E",X"02",X"50",X"28",X"28",X"28",X"28",X"28",X"28",X"28",
		X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",
		X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"FF",X"03",X"50",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"31",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"28",X"28",X"28",
		X"28",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"FF",X"04",X"50",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"28",X"28",X"28",X"28",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"FF",
		X"05",X"50",X"28",X"28",X"28",X"10",X"10",X"28",X"10",X"10",X"28",X"28",X"28",X"10",X"10",X"28",
		X"28",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"28",X"28",X"28",X"28",X"33",X"10",X"28",
		X"28",X"28",X"FF",X"46",X"50",X"28",X"10",X"10",X"28",X"10",X"10",X"28",X"28",X"28",X"10",X"10",
		X"28",X"28",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"28",X"28",X"28",X"28",X"10",X"10",
		X"28",X"FF",X"47",X"50",X"28",X"10",X"10",X"28",X"10",X"10",X"28",X"28",X"28",X"10",X"10",X"28",
		X"28",X"33",X"10",X"28",X"28",X"28",X"28",X"10",X"10",X"28",X"28",X"28",X"28",X"10",X"10",X"28",
		X"FF",X"48",X"50",X"28",X"10",X"10",X"28",X"10",X"10",X"10",X"10",X"28",X"10",X"10",X"28",X"28",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"28",X"FF",
		X"49",X"50",X"28",X"10",X"10",X"28",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"28",X"28",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"28",X"FF",X"0A",
		X"50",X"28",X"28",X"28",X"10",X"10",X"28",X"28",X"28",X"10",X"10",X"10",X"10",X"10",X"28",X"28",
		X"10",X"10",X"10",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"10",X"10",X"28",X"28",
		X"28",X"FF",X"0B",X"50",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"28",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"28",X"28",X"28",X"10",
		X"10",X"10",X"10",X"10",X"FF",X"0C",X"50",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"28",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"31",X"10",X"10",X"10",X"10",X"10",X"10",X"FF",X"0D",X"50",X"28",X"28",X"28",X"28",X"28",X"28",
		X"28",X"28",X"10",X"10",X"28",X"10",X"10",X"2E",X"2E",X"2E",X"2E",X"2E",X"2E",X"10",X"10",X"28",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"28",X"28",X"28",X"FF",X"4E",X"50",X"28",X"28",X"28",
		X"28",X"28",X"28",X"10",X"10",X"28",X"10",X"10",X"2E",X"10",X"10",X"10",X"10",X"2E",X"10",X"10",
		X"28",X"10",X"10",X"28",X"28",X"28",X"28",X"28",X"28",X"FF",X"4F",X"50",X"28",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"28",X"10",X"10",X"2E",X"10",X"10",X"10",X"10",X"2E",X"10",X"10",X"28",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"28",X"FF",X"50",X"50",X"28",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"28",X"10",X"10",X"2E",X"10",X"10",X"10",X"10",X"2E",X"10",X"10",X"28",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"28",X"FF",X"51",X"50",X"28",X"10",X"10",X"28",X"28",X"28",
		X"28",X"28",X"28",X"10",X"10",X"2E",X"10",X"10",X"10",X"10",X"2E",X"10",X"10",X"28",X"28",X"28",
		X"28",X"28",X"28",X"10",X"10",X"28",X"FF",X"12",X"50",X"28",X"28",X"28",X"10",X"10",X"28",X"28",
		X"28",X"28",X"28",X"28",X"10",X"10",X"2E",X"2E",X"2E",X"2E",X"2E",X"2E",X"10",X"10",X"31",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"28",X"28",X"28",X"FF",X"13",X"50",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"31",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"FF",X"14",X"50",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"32",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"28",X"10",X"10",X"28",X"28",X"28",X"10",X"10",X"10",X"10",X"10",X"FF",
		X"15",X"50",X"28",X"28",X"28",X"10",X"10",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"10",
		X"10",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"28",
		X"28",X"28",X"FF",X"56",X"50",X"28",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"28",X"FF",X"57",X"50",X"28",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"28",X"28",X"28",X"28",X"28",X"28",
		X"FF",X"58",X"50",X"28",X"28",X"28",X"28",X"10",X"10",X"28",X"28",X"28",X"28",X"28",X"28",X"28",
		X"10",X"10",X"28",X"28",X"28",X"28",X"28",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"28",X"FF",
		X"59",X"50",X"28",X"10",X"10",X"28",X"33",X"10",X"28",X"10",X"10",X"10",X"28",X"10",X"10",X"10",
		X"10",X"31",X"10",X"10",X"10",X"28",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"28",X"FF",X"1A",
		X"50",X"28",X"28",X"28",X"28",X"28",X"28",X"10",X"10",X"28",X"28",X"28",X"28",X"28",X"10",X"10",
		X"10",X"10",X"32",X"10",X"10",X"10",X"28",X"28",X"28",X"28",X"28",X"28",X"10",X"10",X"28",X"28",
		X"28",X"FF",X"1B",X"50",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"28",X"28",X"28",X"28",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"FF",X"1C",X"50",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"28",X"10",X"10",X"28",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"FF",X"1D",X"50",X"28",X"28",X"28",X"28",X"28",X"28",
		X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",
		X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"FF",X"FF",X"42",X"50",X"2A",X"2A",
		X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",
		X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"FF",X"43",X"50",X"2A",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"2A",X"FF",X"04",X"50",X"2A",X"2A",X"2A",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"2A",X"2A",X"2A",X"FF",X"05",X"50",X"10",
		X"10",X"10",X"10",X"10",X"2A",X"2A",X"10",X"10",X"2A",X"2A",X"10",X"10",X"2A",X"2A",X"2A",X"2A",
		X"2A",X"2A",X"10",X"10",X"2A",X"2A",X"10",X"10",X"2A",X"2A",X"10",X"10",X"10",X"10",X"10",X"FF",
		X"06",X"50",X"10",X"10",X"10",X"10",X"10",X"2A",X"2A",X"10",X"10",X"2A",X"2A",X"33",X"10",X"2A",
		X"2A",X"2A",X"2A",X"2A",X"2A",X"10",X"10",X"2A",X"2A",X"10",X"10",X"2A",X"2A",X"10",X"10",X"10",
		X"10",X"10",X"FF",X"07",X"50",X"2A",X"2A",X"2A",X"33",X"10",X"2A",X"2A",X"10",X"10",X"2A",X"2A",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"31",X"10",X"10",X"2A",X"2A",X"10",X"10",X"2A",X"2A",
		X"33",X"10",X"2A",X"2A",X"2A",X"FF",X"48",X"50",X"2A",X"10",X"10",X"2A",X"2A",X"10",X"10",X"2A",
		X"2A",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"2A",X"2A",X"10",X"10",X"2A",
		X"2A",X"10",X"10",X"2A",X"FF",X"49",X"50",X"2A",X"10",X"10",X"2A",X"2A",X"10",X"10",X"2A",X"2A",
		X"2A",X"2A",X"2A",X"2A",X"10",X"10",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"10",X"10",X"2A",X"2A",
		X"10",X"10",X"2A",X"FF",X"0A",X"50",X"2A",X"2A",X"2A",X"10",X"10",X"2A",X"2A",X"10",X"10",X"2A",
		X"2A",X"2A",X"2A",X"2A",X"2A",X"10",X"10",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"10",X"10",X"2A",
		X"2A",X"10",X"10",X"2A",X"2A",X"2A",X"FF",X"0B",X"50",X"10",X"10",X"10",X"10",X"10",X"2A",X"2A",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"2A",X"2A",X"10",X"10",X"10",X"10",X"10",X"FF",X"0C",X"50",X"10",X"10",X"10",X"10",
		X"10",X"2A",X"2A",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"2A",X"2A",X"10",X"10",X"10",X"10",X"10",X"FF",X"0D",X"50",X"2A",
		X"2A",X"2A",X"10",X"10",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"10",X"10",X"2E",X"2E",X"2E",X"2E",
		X"2E",X"2E",X"10",X"10",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"10",X"10",X"2A",X"2A",X"2A",X"FF",
		X"4E",X"50",X"2A",X"10",X"10",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"10",X"10",X"2E",X"10",X"10",
		X"10",X"10",X"2E",X"10",X"10",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"10",X"10",X"2A",X"FF",X"4F",
		X"50",X"2A",X"10",X"10",X"10",X"10",X"10",X"10",X"2A",X"2A",X"10",X"10",X"2E",X"10",X"10",X"10",
		X"10",X"2E",X"10",X"10",X"2A",X"2A",X"10",X"10",X"10",X"31",X"10",X"10",X"2A",X"FF",X"50",X"50",
		X"2A",X"10",X"10",X"10",X"10",X"10",X"10",X"2A",X"2A",X"10",X"10",X"2E",X"10",X"10",X"10",X"10",
		X"2E",X"10",X"10",X"2A",X"2A",X"10",X"10",X"10",X"10",X"10",X"10",X"2A",X"FF",X"51",X"50",X"2A",
		X"33",X"10",X"2A",X"2A",X"10",X"10",X"2A",X"2A",X"10",X"10",X"2E",X"10",X"10",X"10",X"10",X"2E",
		X"10",X"10",X"2A",X"2A",X"10",X"10",X"2A",X"2A",X"10",X"10",X"2A",X"FF",X"12",X"50",X"2A",X"2A",
		X"2A",X"10",X"10",X"2A",X"2A",X"10",X"10",X"2A",X"2A",X"10",X"10",X"2E",X"2E",X"2E",X"2E",X"2E",
		X"2E",X"10",X"10",X"2A",X"2A",X"33",X"10",X"2A",X"2A",X"10",X"10",X"2A",X"2A",X"2A",X"FF",X"13",
		X"50",X"10",X"10",X"10",X"10",X"10",X"2A",X"2A",X"10",X"10",X"2A",X"2A",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"2A",X"2A",X"10",X"10",X"2A",X"2A",X"10",X"10",X"10",X"10",
		X"10",X"FF",X"14",X"50",X"10",X"10",X"10",X"10",X"10",X"2A",X"2A",X"10",X"10",X"31",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"2A",X"2A",X"10",
		X"10",X"10",X"10",X"10",X"FF",X"15",X"50",X"2A",X"2A",X"2A",X"10",X"10",X"2A",X"2A",X"10",X"10",
		X"10",X"10",X"10",X"10",X"2A",X"2A",X"10",X"10",X"2A",X"2A",X"10",X"10",X"10",X"10",X"10",X"10",
		X"2A",X"2A",X"10",X"10",X"2A",X"2A",X"2A",X"FF",X"56",X"50",X"2A",X"10",X"10",X"2A",X"2A",X"2A",
		X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"10",X"10",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",
		X"2A",X"2A",X"2A",X"10",X"10",X"2A",X"FF",X"57",X"50",X"2A",X"10",X"10",X"2A",X"2A",X"2A",X"2A",
		X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"10",X"10",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",
		X"2A",X"2A",X"10",X"10",X"2A",X"FF",X"58",X"50",X"2A",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"31",X"10",X"10",X"10",
		X"10",X"10",X"10",X"2A",X"FF",X"59",X"50",X"2A",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"2A",X"FF",X"5A",X"50",X"2A",X"10",X"10",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",
		X"2A",X"10",X"10",X"2A",X"2A",X"10",X"10",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"33",
		X"10",X"2A",X"FF",X"5B",X"50",X"2A",X"10",X"10",X"10",X"10",X"10",X"10",X"31",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"2A",X"FF",X"5C",X"50",X"2A",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"2A",
		X"FF",X"5D",X"50",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",
		X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
