library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity tron_sp_bits_2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of tron_sp_bits_2 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",
		X"00",X"77",X"22",X"00",X"00",X"77",X"22",X"00",X"00",X"22",X"77",X"00",X"00",X"22",X"77",X"00",
		X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"00",X"22",X"00",
		X"00",X"00",X"22",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"22",X"00",X"00",
		X"00",X"22",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"22",X"00",X"22",X"77",X"22",X"00",X"22",X"77",
		X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",
		X"77",X"00",X"66",X"00",X"77",X"00",X"66",X"00",X"00",X"00",X"62",X"00",X"00",X"00",X"77",X"00",
		X"22",X"66",X"22",X"77",X"22",X"66",X"22",X"77",X"00",X"22",X"77",X"22",X"00",X"22",X"77",X"22",
		X"00",X"22",X"77",X"22",X"00",X"22",X"77",X"22",X"00",X"66",X"22",X"00",X"00",X"66",X"22",X"00",
		X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"22",X"00",X"22",X"77",X"22",X"00",X"22",X"77",
		X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",
		X"77",X"00",X"66",X"00",X"77",X"00",X"66",X"00",X"00",X"00",X"62",X"00",X"00",X"00",X"77",X"00",
		X"22",X"66",X"22",X"77",X"22",X"66",X"22",X"77",X"00",X"22",X"77",X"22",X"00",X"22",X"77",X"22",
		X"00",X"22",X"77",X"22",X"00",X"22",X"77",X"22",X"00",X"66",X"22",X"00",X"00",X"66",X"22",X"00",
		X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",
		X"CC",X"77",X"00",X"00",X"CC",X"77",X"CC",X"00",X"00",X"22",X"77",X"77",X"00",X"22",X"77",X"77",
		X"CC",X"22",X"77",X"77",X"CC",X"22",X"77",X"77",X"77",X"22",X"22",X"77",X"77",X"22",X"22",X"27",
		X"72",X"22",X"22",X"0C",X"22",X"22",X"22",X"CC",X"77",X"22",X"72",X"77",X"77",X"22",X"77",X"77",
		X"CC",X"22",X"27",X"22",X"CC",X"22",X"77",X"27",X"CC",X"22",X"27",X"77",X"CC",X"22",X"22",X"77",
		X"77",X"77",X"22",X"CC",X"77",X"77",X"22",X"00",X"77",X"22",X"22",X"77",X"77",X"22",X"22",X"77",
		X"CC",X"22",X"77",X"22",X"CC",X"22",X"77",X"22",X"00",X"27",X"77",X"77",X"00",X"77",X"77",X"77",
		X"00",X"CC",X"77",X"CC",X"00",X"CC",X"77",X"CC",X"CC",X"00",X"55",X"00",X"CC",X"00",X"55",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"A0",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0A",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",
		X"00",X"00",X"A0",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",
		X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"00",X"00",X"00",X"BC",X"00",X"00",X"0C",X"BB",X"00",X"00",X"0C",X"BB",X"00",
		X"00",X"0C",X"BB",X"00",X"00",X"0C",X"BB",X"00",X"00",X"00",X"BC",X"00",X"00",X"00",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"BC",X"00",
		X"00",X"00",X"BC",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"01",X"11",X"02",X"00",X"11",X"11",X"22",X"00",X"12",X"31",X"1C",X"00",X"1A",
		X"31",X"A1",X"00",X"12",X"31",X"00",X"00",X"12",X"31",X"00",X"00",X"12",X"31",X"11",X"11",X"1A",
		X"31",X"DD",X"DD",X"12",X"31",X"DD",X"DD",X"12",X"31",X"DD",X"DD",X"12",X"31",X"DD",X"DD",X"1A",
		X"31",X"DD",X"DD",X"12",X"31",X"DD",X"DD",X"12",X"31",X"DD",X"DD",X"12",X"31",X"DD",X"22",X"12",
		X"31",X"DD",X"33",X"1A",X"31",X"DD",X"D3",X"12",X"31",X"DD",X"D3",X"12",X"31",X"DD",X"33",X"12",
		X"31",X"DD",X"33",X"12",X"31",X"DD",X"D3",X"1A",X"31",X"DD",X"D3",X"12",X"31",X"DD",X"33",X"12",
		X"31",X"DA",X"22",X"12",X"31",X"DD",X"DD",X"1A",X"31",X"11",X"11",X"12",X"31",X"00",X"00",X"12",
		X"31",X"00",X"00",X"1A",X"11",X"00",X"00",X"12",X"11",X"00",X"00",X"11",X"01",X"00",X"00",X"01",
		X"01",X"11",X"11",X"11",X"11",X"DD",X"DD",X"DD",X"13",X"33",X"33",X"33",X"11",X"11",X"11",X"11",
		X"2A",X"2A",X"22",X"22",X"11",X"11",X"11",X"11",X"11",X"33",X"33",X"33",X"01",X"33",X"22",X"31",
		X"00",X"11",X"23",X"11",X"00",X"DD",X"33",X"D0",X"00",X"DD",X"D3",X"10",X"00",X"DD",X"D3",X"10",
		X"00",X"DD",X"33",X"10",X"00",X"DD",X"D3",X"10",X"21",X"DD",X"D3",X"10",X"2C",X"DD",X"33",X"10",
		X"33",X"11",X"23",X"10",X"33",X"33",X"22",X"10",X"33",X"33",X"33",X"10",X"33",X"1A",X"1A",X"10",
		X"2C",X"DD",X"DD",X"10",X"21",X"DD",X"DD",X"10",X"00",X"DD",X"DD",X"10",X"00",X"11",X"11",X"11",
		X"01",X"33",X"33",X"31",X"11",X"33",X"33",X"33",X"11",X"11",X"11",X"11",X"2A",X"2A",X"22",X"22",
		X"11",X"11",X"11",X"11",X"13",X"33",X"33",X"33",X"11",X"DD",X"DD",X"DD",X"01",X"11",X"11",X"11",
		X"55",X"00",X"00",X"55",X"5A",X"00",X"00",X"CC",X"C5",X"00",X"00",X"CC",X"C5",X"00",X"00",X"CC",
		X"C5",X"00",X"00",X"C6",X"55",X"00",X"00",X"CC",X"5A",X"00",X"00",X"CC",X"C5",X"00",X"22",X"CC",
		X"C5",X"22",X"22",X"CC",X"C5",X"22",X"C2",X"C6",X"55",X"22",X"7C",X"CC",X"5A",X"22",X"7C",X"CC",
		X"C5",X"2C",X"77",X"CC",X"C5",X"C7",X"77",X"CC",X"C5",X"77",X"57",X"C6",X"55",X"77",X"55",X"CC",
		X"5A",X"75",X"55",X"CC",X"C5",X"55",X"55",X"CC",X"C5",X"55",X"55",X"CC",X"C5",X"55",X"55",X"C6",
		X"55",X"55",X"55",X"CC",X"5A",X"75",X"55",X"CC",X"C5",X"77",X"55",X"CC",X"C5",X"C7",X"57",X"CC",
		X"C5",X"C7",X"77",X"C6",X"55",X"CC",X"CC",X"CC",X"5A",X"07",X"22",X"CC",X"C5",X"07",X"22",X"CC",
		X"55",X"07",X"77",X"CC",X"55",X"07",X"0C",X"5C",X"05",X"07",X"00",X"55",X"05",X"07",X"00",X"05",
		X"55",X"C2",X"52",X"25",X"55",X"C2",X"52",X"25",X"5C",X"C5",X"CC",X"55",X"A5",X"55",X"55",X"5A",
		X"CC",X"6C",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"55",X"66",X"66",X"6A",X"05",X"CC",X"CC",X"CC",
		X"00",X"55",X"CC",X"55",X"00",X"55",X"77",X"50",X"00",X"55",X"55",X"C0",X"00",X"55",X"55",X"C7",
		X"00",X"5C",X"55",X"C2",X"00",X"C7",X"55",X"C2",X"00",X"7C",X"55",X"C2",X"00",X"C7",X"55",X"C2",
		X"00",X"C7",X"55",X"C2",X"00",X"7C",X"55",X"C2",X"00",X"C7",X"55",X"C2",X"00",X"5C",X"55",X"C2",
		X"00",X"55",X"55",X"C7",X"00",X"55",X"55",X"C0",X"00",X"55",X"77",X"50",X"00",X"55",X"CC",X"55",
		X"05",X"CC",X"CC",X"CC",X"55",X"66",X"66",X"6A",X"CC",X"CC",X"CC",X"CC",X"CC",X"6C",X"CC",X"CC",
		X"A5",X"55",X"55",X"5A",X"5C",X"C5",X"CC",X"55",X"55",X"C2",X"52",X"25",X"55",X"CC",X"5C",X"C5",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"0A",X"F0",X"00",
		X"00",X"FA",X"3F",X"00",X"00",X"59",X"33",X"00",X"00",X"55",X"93",X"90",X"00",X"55",X"59",X"00",
		X"00",X"53",X"AA",X"00",X"00",X"33",X"A5",X"00",X"00",X"39",X"55",X"00",X"00",X"99",X"55",X"00",
		X"00",X"55",X"55",X"F0",X"00",X"33",X"99",X"00",X"00",X"93",X"99",X"00",X"00",X"39",X"A9",X"00",
		X"00",X"93",X"AA",X"00",X"00",X"93",X"53",X"00",X"00",X"33",X"33",X"50",X"00",X"33",X"3A",X"00",
		X"00",X"33",X"3F",X"00",X"00",X"33",X"F0",X"00",X"00",X"33",X"00",X"00",X"00",X"30",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"05",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"02",X"00",X"EE",X"22",X"23",X"0E",X"EE",X"22",
		X"32",X"2E",X"EE",X"00",X"23",X"00",X"E0",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",
		X"00",X"22",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"02",X"E2",X"00",
		X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"22",X"00",
		X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"20",X"00",X"00",X"22",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"23",X"00",
		X"00",X"00",X"22",X"00",X"00",X"00",X"02",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"02",
		X"00",X"00",X"00",X"02",X"00",X"00",X"A0",X"00",X"00",X"00",X"AA",X"33",X"00",X"00",X"2A",X"B3",
		X"00",X"00",X"22",X"B3",X"00",X"00",X"22",X"B3",X"00",X"00",X"72",X"B3",X"00",X"00",X"A7",X"B3",
		X"00",X"00",X"AA",X"B3",X"00",X"00",X"0A",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",
		X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"20",X"00",X"00",X"02",X"20",X"00",X"00",X"22",X"00",
		X"00",X"00",X"23",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"02",X"20",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"22",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"22",X"00",X"00",X"02",X"20",X"00",
		X"00",X"02",X"00",X"00",X"DD",X"20",X"00",X"00",X"D6",X"20",X"00",X"00",X"D6",X"00",X"00",X"00",
		X"D6",X"DD",X"00",X"00",X"D7",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"0D",X"DD",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"02",X"00",X"00",
		X"00",X"02",X"20",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"22",X"20",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"07",X"CF",X"00",X"00",X"FF",X"7C",X"00",X"00",X"FF",X"7C",X"00",X"00",X"FF",X"7C",
		X"00",X"00",X"FF",X"7C",X"00",X"00",X"07",X"CF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"7C",X"00",X"00",X"00",X"7C",X"00",
		X"00",X"00",X"07",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",
		X"00",X"00",X"0F",X"C7",X"00",X"00",X"07",X"7C",X"00",X"00",X"FF",X"7C",X"00",X"00",X"FF",X"7C",
		X"00",X"00",X"FF",X"7C",X"00",X"00",X"FF",X"CF",X"00",X"00",X"07",X"FF",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"70",X"00",
		X"00",X"00",X"77",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"70",X"00",
		X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",
		X"00",X"00",X"07",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F7",
		X"00",X"00",X"0F",X"CF",X"00",X"00",X"0F",X"7C",X"00",X"00",X"7F",X"7C",X"00",X"00",X"FF",X"7C",
		X"00",X"00",X"FF",X"7C",X"00",X"00",X"FF",X"CF",X"00",X"00",X"0F",X"FF",X"00",X"00",X"00",X"70",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"70",X"00",
		X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"0F",X"CF",X"00",X"00",X"FF",X"7C",X"00",X"00",X"FF",X"7C",X"00",X"00",X"7F",X"7C",
		X"00",X"00",X"FF",X"7C",X"00",X"00",X"FF",X"CF",X"00",X"00",X"0F",X"FF",X"00",X"00",X"00",X"77",
		X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"2C",X"00",X"00",
		X"00",X"0C",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"F7",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"0F",X"FF",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"0F",X"CF",X"00",X"00",X"FF",X"7C",X"00",X"00",X"FF",X"7C",X"00",X"00",X"FF",X"7C",
		X"00",X"00",X"7F",X"7C",X"00",X"00",X"FF",X"CF",X"00",X"00",X"0F",X"F7",X"00",X"00",X"00",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"70",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"C7",X"00",X"00",X"00",X"CC",X"00",X"00",
		X"00",X"7C",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"FF",X"CF",X"00",X"00",X"0F",X"7C",X"00",X"00",X"0F",X"7C",X"00",X"00",X"0F",X"7C",
		X"00",X"00",X"07",X"7C",X"00",X"00",X"0F",X"CF",X"00",X"00",X"0F",X"FF",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"70",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"C7",X"00",X"00",X"00",X"CC",X"00",X"00",
		X"00",X"7C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"FF",X"CF",X"00",X"00",X"0F",X"7C",X"00",X"00",X"0F",X"7C",X"00",X"00",X"0F",X"7C",
		X"00",X"00",X"07",X"7C",X"00",X"00",X"0F",X"CF",X"00",X"00",X"0F",X"FF",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C7",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",
		X"0C",X"00",X"00",X"00",X"07",X"77",X"00",X"00",X"00",X"77",X"00",X"FF",X"00",X"07",X"FF",X"F7",
		X"00",X"00",X"FF",X"CF",X"00",X"00",X"FF",X"7C",X"00",X"00",X"FF",X"7C",X"00",X"00",X"FF",X"7C",
		X"00",X"00",X"0F",X"7C",X"00",X"00",X"0F",X"CF",X"00",X"00",X"07",X"FF",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"7C",X"00",X"00",X"F0",X"CC",X"70",X"0F",X"F7",
		X"7C",X"77",X"FF",X"FF",X"07",X"77",X"FF",X"CF",X"00",X"00",X"FF",X"7C",X"00",X"00",X"FF",X"7C",
		X"00",X"00",X"0F",X"7C",X"00",X"00",X"0F",X"7C",X"00",X"00",X"0F",X"CF",X"00",X"00",X"00",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"F0",X"00",X"00",X"FF",X"FF",X"07",X"00",X"FC",X"CF",X"CC",X"77",X"FC",X"CF",
		X"CC",X"77",X"FC",X"CF",X"07",X"00",X"FC",X"CF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"0F",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"30",X"00",X"EE",X"39",X"93",X"33",X"EE",X"E9",X"99",
		X"E9",X"99",X"99",X"99",X"9E",X"9E",X"99",X"EE",X"9C",X"E9",X"99",X"99",X"EC",X"99",X"99",X"99",
		X"EC",X"99",X"99",X"33",X"9C",X"E9",X"E9",X"EE",X"93",X"EE",X"E9",X"99",X"30",X"EE",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"3E",X"33",X"00",X"00",
		X"9E",X"99",X"00",X"00",X"EE",X"EE",X"00",X"00",X"E9",X"99",X"00",X"00",X"E9",X"33",X"00",X"00",
		X"33",X"EE",X"00",X"00",X"EE",X"99",X"00",X"00",X"E9",X"33",X"00",X"00",X"33",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"33",X"00",X"EE",X"39",X"9E",X"33",X"EE",X"E9",X"9E",
		X"E9",X"99",X"99",X"EE",X"9E",X"9E",X"99",X"99",X"9C",X"E9",X"99",X"99",X"EC",X"99",X"99",X"93",
		X"EC",X"99",X"99",X"33",X"9C",X"E9",X"E9",X"99",X"93",X"EE",X"E9",X"EE",X"30",X"EE",X"33",X"9E",
		X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"93",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"99",X"00",X"00",X"33",X"33",X"00",X"00",X"9E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"93",X"00",X"00",X"00",X"30",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",
		X"E9",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"9E",X"33",X"00",X"00",X"99",X"E9",X"00",X"00",
		X"33",X"EE",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"9E",X"00",X"00",
		X"00",X"9E",X"00",X"00",X"00",X"E3",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"4E",X"E0",X"00",X"00",X"44",X"EE",X"00",
		X"00",X"04",X"E9",X"99",X"00",X"00",X"EE",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"04",X"EE",X"00",
		X"00",X"44",X"EE",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"E9",X"00",
		X"00",X"00",X"99",X"00",X"00",X"40",X"00",X"00",X"00",X"4E",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"9E",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"EE",X"00",X"00",X"04",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"9E",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9E",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",
		X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",
		X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",
		X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"EE",X"40",X"00",X"00",X"E9",X"40",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",
		X"00",X"00",X"40",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"09",X"E0",X"00",X"99",X"0F",X"E9",X"00",X"EE",X"CC",X"CC",X"E0",
		X"EE",X"EE",X"CC",X"E0",X"EE",X"CC",X"CC",X"E0",X"EC",X"CC",X"CC",X"FF",X"EC",X"CC",X"CC",X"FF",
		X"EC",X"CC",X"CC",X"FF",X"EC",X"CC",X"CC",X"FF",X"EE",X"CC",X"CC",X"E0",X"EE",X"EE",X"CC",X"E0",
		X"EE",X"CC",X"CC",X"E0",X"99",X"0F",X"E9",X"00",X"00",X"09",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"EE",X"00",X"00",X"9E",X"EE",X"00",X"00",X"9E",X"EE",X"00",
		X"00",X"9E",X"CE",X"00",X"00",X"9E",X"CE",X"00",X"00",X"9E",X"CE",X"00",X"00",X"9E",X"CE",X"00",
		X"00",X"0C",X"CE",X"00",X"00",X"0C",X"CE",X"00",X"00",X"0C",X"CE",X"00",X"00",X"FC",X"CE",X"00",
		X"00",X"EC",X"CE",X"00",X"00",X"EC",X"CE",X"00",X"00",X"EC",X"CE",X"00",X"00",X"EC",X"CE",X"00",
		X"00",X"EC",X"CE",X"00",X"00",X"EC",X"CE",X"00",X"00",X"EC",X"CC",X"00",X"00",X"9C",X"CC",X"00",
		X"00",X"EC",X"CC",X"00",X"00",X"E9",X"CC",X"00",X"00",X"09",X"CC",X"00",X"00",X"0E",X"1C",X"00",
		X"00",X"0E",X"CC",X"00",X"00",X"0E",X"CC",X"00",X"00",X"0E",X"EE",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"70",X"00",X"FF",X"0F",X"74",X"00",X"77",X"CC",X"CC",X"70",
		X"77",X"77",X"CC",X"70",X"77",X"CC",X"CC",X"70",X"7C",X"CC",X"CC",X"FF",X"7C",X"CC",X"CC",X"FF",
		X"7C",X"CC",X"CC",X"FF",X"7C",X"CC",X"CC",X"FF",X"77",X"CC",X"CC",X"70",X"77",X"77",X"CC",X"70",
		X"77",X"CC",X"CC",X"70",X"FF",X"0F",X"74",X"00",X"00",X"0F",X"70",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"70",X"00",X"00",X"00",X"77",X"00",X"00",X"F7",X"77",X"00",X"00",X"F7",X"77",X"00",
		X"00",X"F7",X"C7",X"00",X"00",X"F7",X"C7",X"00",X"00",X"F7",X"C7",X"00",X"00",X"F7",X"C7",X"00",
		X"00",X"0C",X"C7",X"00",X"00",X"0C",X"C7",X"00",X"00",X"0C",X"C7",X"00",X"00",X"FC",X"C7",X"00",
		X"00",X"7C",X"C7",X"00",X"00",X"7C",X"C7",X"00",X"00",X"7C",X"C7",X"00",X"00",X"7C",X"C7",X"00",
		X"00",X"7C",X"C7",X"00",X"00",X"7C",X"C7",X"00",X"00",X"7C",X"CC",X"00",X"00",X"4C",X"CC",X"00",
		X"00",X"7C",X"CC",X"00",X"00",X"74",X"CC",X"00",X"00",X"04",X"CC",X"00",X"00",X"07",X"4C",X"00",
		X"00",X"07",X"CC",X"00",X"00",X"07",X"CC",X"00",X"00",X"07",X"77",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"31",X"31",X"31",X"00",X"13",X"13",X"13",X"00",X"31",X"31",X"31",X"00",X"11",X"11",X"11",
		X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"01",X"11",X"11",X"11",X"01",X"11",X"11",X"11",
		X"01",X"11",X"11",X"11",X"01",X"11",X"11",X"11",X"11",X"11",X"11",X"10",X"11",X"11",X"11",X"10",
		X"11",X"11",X"11",X"10",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",
		X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"53",X"53",X"53",X"00",X"35",X"35",X"35",X"00",X"53",X"53",X"53",X"00",X"35",X"35",X"35",
		X"00",X"53",X"53",X"53",X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",
		X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",
		X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",
		X"03",X"33",X"33",X"33",X"03",X"33",X"33",X"33",X"03",X"33",X"33",X"33",X"03",X"33",X"33",X"33",
		X"13",X"13",X"13",X"10",X"31",X"31",X"31",X"30",X"13",X"13",X"13",X"00",X"31",X"31",X"31",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"B5",X"B5",X"B5",X"00",X"5B",X"5B",X"5B",X"00",X"B5",X"B5",X"B5",X"00",X"5B",X"5B",X"5B",
		X"00",X"B5",X"B5",X"B5",X"00",X"5B",X"5B",X"5B",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",
		X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",
		X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",
		X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",
		X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",
		X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"35",X"35",X"35",
		X"00",X"53",X"53",X"53",X"00",X"35",X"35",X"35",X"00",X"53",X"53",X"53",X"05",X"35",X"35",X"35",
		X"0B",X"DB",X"DB",X"DB",X"00",X"BD",X"BD",X"BD",X"00",X"DB",X"DB",X"DB",X"00",X"BD",X"BD",X"BD",
		X"00",X"DB",X"DB",X"DB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",
		X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",
		X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",
		X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",
		X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",
		X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"B5",X"B5",X"B5",X"00",X"5B",X"5B",X"5B",
		X"00",X"B5",X"B5",X"B5",X"00",X"5B",X"5B",X"5B",X"00",X"B5",X"B5",X"B5",X"00",X"5B",X"5B",X"5B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DF",X"DF",X"DF",X"00",X"FD",X"FD",X"FD",X"00",X"DF",X"DF",X"DF",X"00",X"FD",X"FD",X"FD",X"00",
		X"DD",X"DD",X"DD",X"D0",X"DD",X"DD",X"DD",X"D0",X"DD",X"DD",X"DD",X"D0",X"DD",X"DD",X"DD",X"D0",
		X"0D",X"DD",X"DD",X"DD",X"0D",X"DD",X"DD",X"DD",X"0D",X"DD",X"DD",X"DD",X"0D",X"DD",X"DD",X"DD",
		X"00",X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",
		X"00",X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",X"BD",X"BD",X"BD",
		X"00",X"DB",X"DB",X"DB",X"00",X"BD",X"BD",X"BD",X"00",X"DB",X"DB",X"DB",X"00",X"BD",X"BD",X"BD",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",
		X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"F0",
		X"FF",X"FF",X"FF",X"F0",X"FF",X"FF",X"FF",X"F0",X"0F",X"FF",X"FF",X"FF",X"0F",X"FF",X"FF",X"FF",
		X"0F",X"FF",X"FF",X"FF",X"0F",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",
		X"00",X"FF",X"FF",X"FF",X"00",X"DF",X"DF",X"DF",X"00",X"FD",X"FD",X"FD",X"00",X"DF",X"DF",X"DF",
		X"06",X"60",X"60",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"66",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"66",X"50",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"05",X"05",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"05",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"44",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"44",X"04",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"40",X"00",X"00",
		X"06",X"60",X"60",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"66",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"50",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"55",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"44",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"44",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",
		X"00",X"7F",X"00",X"00",X"00",X"A0",X"00",X"02",X"00",X"00",X"A0",X"79",X"00",X"B0",X"7F",X"00",
		X"00",X"00",X"00",X"09",X"00",X"A0",X"00",X"0A",X"00",X"00",X"00",X"50",X"00",X"F0",X"90",X"00",
		X"A0",X"07",X"09",X"00",X"0A",X"A0",X"90",X"A0",X"79",X"09",X"09",X"02",X"00",X"E0",X"20",X"90",
		X"00",X"00",X"0B",X"05",X"00",X"A0",X"A0",X"E0",X"00",X"09",X"00",X"02",X"00",X"E0",X"00",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"07",X"00",X"00",X"00",X"90",X"07",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",
		X"00",X"70",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"07",X"11",X"00",X"00",
		X"03",X"99",X"00",X"00",X"03",X"99",X"00",X"00",X"03",X"99",X"00",X"00",X"03",X"79",X"00",X"00",
		X"03",X"79",X"00",X"00",X"03",X"79",X"07",X"00",X"03",X"79",X"00",X"00",X"03",X"93",X"00",X"00",
		X"03",X"93",X"00",X"00",X"03",X"93",X"00",X"07",X"04",X"93",X"00",X"00",X"44",X"44",X"00",X"00",
		X"44",X"43",X"00",X"00",X"44",X"93",X"00",X"00",X"04",X"93",X"00",X"07",X"03",X"93",X"00",X"00",
		X"03",X"93",X"00",X"00",X"03",X"79",X"00",X"00",X"07",X"79",X"07",X"00",X"00",X"79",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"11",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"70",X"00",X"77",X"55",X"50",X"00",X"55",
		X"5C",X"00",X"00",X"CC",X"5C",X"00",X"00",X"CC",X"5C",X"00",X"00",X"CC",X"5C",X"00",X"00",X"CC",
		X"5C",X"00",X"00",X"CC",X"5C",X"00",X"00",X"CC",X"5C",X"00",X"00",X"CC",X"5C",X"00",X"00",X"CC",
		X"5C",X"00",X"00",X"CC",X"5C",X"00",X"00",X"CC",X"55",X"00",X"50",X"55",X"00",X"00",X"C5",X"00",
		X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"5C",X"CC",X"55",X"CC",
		X"5C",X"C5",X"00",X"CC",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"00",
		X"00",X"55",X"CC",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"50",X"00",X"00",X"CC",X"50",X"00",
		X"00",X"CC",X"50",X"00",X"00",X"CC",X"50",X"00",X"00",X"C5",X"50",X"00",X"00",X"50",X"00",X"00",
		X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",
		X"00",X"00",X"05",X"05",X"00",X"00",X"5C",X"05",X"00",X"00",X"5C",X"05",X"00",X"00",X"5C",X"05",
		X"00",X"00",X"5C",X"05",X"00",X"00",X"5C",X"05",X"00",X"00",X"5C",X"05",X"00",X"00",X"05",X"05",
		X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",
		X"00",X"50",X"00",X"00",X"00",X"C5",X"50",X"00",X"00",X"CC",X"50",X"00",X"00",X"CC",X"50",X"00",
		X"00",X"CC",X"50",X"00",X"00",X"55",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
