library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity bg_map is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of bg_map is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"0B",X"09",X"0A",X"0B",X"09",X"0A",X"0B",X"09",X"0A",X"0B",X"09",X"0A",X"02",X"00",
		X"00",X"05",X"06",X"00",X"05",X"06",X"07",X"05",X"06",X"00",X"05",X"06",X"00",X"05",X"06",X"00",
		X"00",X"03",X"0D",X"09",X"0C",X"04",X"07",X"03",X"0D",X"09",X"0C",X"0D",X"09",X"0C",X"04",X"00",
		X"00",X"00",X"00",X"07",X"03",X"0D",X"08",X"0C",X"04",X"07",X"05",X"06",X"00",X"05",X"06",X"00",
		X"00",X"01",X"0B",X"08",X"0C",X"04",X"00",X"05",X"06",X"07",X"03",X"0D",X"09",X"0C",X"04",X"00",
		X"00",X"05",X"06",X"07",X"03",X"0D",X"09",X"0C",X"0D",X"08",X"0C",X"04",X"07",X"00",X"00",X"00",
		X"00",X"05",X"06",X"07",X"05",X"06",X"00",X"05",X"06",X"00",X"03",X"0D",X"08",X"0A",X"02",X"00",
		X"00",X"03",X"0D",X"08",X"0C",X"0D",X"09",X"0C",X"0D",X"09",X"0C",X"04",X"07",X"05",X"06",X"00",
		X"00",X"05",X"06",X"00",X"05",X"06",X"00",X"05",X"06",X"00",X"05",X"06",X"07",X"05",X"06",X"00",
		X"00",X"03",X"0D",X"09",X"0C",X"0D",X"09",X"0C",X"0D",X"09",X"0C",X"0D",X"08",X"0C",X"04",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"0B",X"09",X"0A",X"0B",X"09",X"0A",X"0B",X"09",X"0A",X"0B",X"09",X"0A",X"02",X"00",
		X"00",X"03",X"0D",X"08",X"0C",X"0D",X"08",X"0C",X"04",X"07",X"05",X"06",X"07",X"05",X"06",X"00",
		X"00",X"03",X"0D",X"08",X"0C",X"04",X"07",X"03",X"0D",X"08",X"0C",X"0D",X"08",X"0C",X"04",X"00",
		X"00",X"05",X"06",X"07",X"03",X"0D",X"08",X"0C",X"04",X"07",X"03",X"0D",X"08",X"0C",X"04",X"00",
		X"00",X"03",X"0D",X"08",X"0C",X"0D",X"08",X"0C",X"0D",X"08",X"0C",X"0D",X"08",X"0C",X"04",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"03",X"0D",X"08",X"0A",X"02",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"0B",X"08",X"0C",X"04",X"07",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"03",X"0D",X"08",X"0A",X"02",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"0B",X"08",X"0C",X"0D",X"08",X"0A",X"02",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"0B",X"09",X"0A",X"0B",X"09",X"0A",X"0B",X"09",X"0A",X"0B",X"09",X"0A",X"02",X"00",
		X"00",X"03",X"0D",X"09",X"0C",X"0D",X"08",X"0A",X"0B",X"08",X"0A",X"0B",X"09",X"0C",X"04",X"00",
		X"00",X"03",X"0D",X"09",X"0C",X"0D",X"09",X"0C",X"04",X"00",X"03",X"0D",X"09",X"0C",X"04",X"00",
		X"00",X"03",X"0D",X"09",X"0A",X"0B",X"08",X"0C",X"0D",X"09",X"0C",X"0D",X"09",X"0C",X"04",X"00",
		X"00",X"00",X"00",X"00",X"03",X"04",X"07",X"03",X"0D",X"08",X"0A",X"02",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"0D",X"08",X"0C",X"0D",X"09",X"0C",X"04",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"04",X"00",X"00",X"00",X"00",X"05",X"06",X"00",X"00",X"00",X"00",
		X"00",X"01",X"0B",X"09",X"0C",X"04",X"00",X"00",X"00",X"00",X"03",X"0D",X"09",X"0A",X"02",X"00",
		X"00",X"03",X"0D",X"08",X"0C",X"04",X"00",X"00",X"00",X"00",X"03",X"0D",X"09",X"0C",X"04",X"00",
		X"00",X"03",X"0D",X"08",X"0C",X"04",X"00",X"00",X"00",X"00",X"03",X"0D",X"08",X"0C",X"04",X"00",
		X"00",X"00",X"00",X"00",X"03",X"0D",X"09",X"0A",X"0B",X"09",X"0C",X"04",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"0D",X"08",X"0A",X"0B",X"08",X"0C",X"04",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"0B",X"09",X"0A",X"0B",X"09",X"0A",X"0B",X"09",X"0A",X"0B",X"09",X"0A",X"02",X"00",
		X"00",X"03",X"0D",X"09",X"0C",X"0D",X"09",X"0C",X"0D",X"09",X"0C",X"0D",X"09",X"0C",X"04",X"00",
		X"00",X"01",X"0B",X"08",X"0A",X"0B",X"08",X"0A",X"0B",X"08",X"0A",X"0B",X"08",X"0A",X"02",X"00",
		X"00",X"03",X"0D",X"09",X"0C",X"0D",X"09",X"0C",X"0D",X"09",X"0C",X"0D",X"09",X"0C",X"04",X"00",
		X"00",X"01",X"0B",X"08",X"0A",X"0B",X"08",X"0C",X"0D",X"08",X"0A",X"0B",X"08",X"0A",X"02",X"00",
		X"00",X"03",X"0D",X"09",X"0C",X"0D",X"09",X"0C",X"0D",X"09",X"0C",X"0D",X"09",X"0C",X"04",X"00",
		X"00",X"03",X"0D",X"08",X"0A",X"0B",X"08",X"0A",X"0B",X"08",X"0A",X"0B",X"08",X"0C",X"04",X"00",
		X"00",X"03",X"0D",X"09",X"0C",X"0D",X"09",X"0C",X"0D",X"09",X"0C",X"0D",X"09",X"0C",X"04",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"0B",X"09",X"0A",X"0B",X"09",X"0A",X"0B",X"09",X"0A",X"0B",X"09",X"0A",X"02",X"00",
		X"00",X"03",X"0D",X"09",X"0A",X"0B",X"09",X"0A",X"0B",X"09",X"0A",X"0B",X"08",X"0C",X"04",X"00",
		X"00",X"01",X"0B",X"09",X"0A",X"0B",X"09",X"0C",X"0D",X"09",X"0C",X"04",X"07",X"05",X"06",X"00",
		X"00",X"03",X"0D",X"09",X"0A",X"0B",X"09",X"0A",X"0B",X"09",X"0A",X"02",X"07",X"05",X"06",X"00",
		X"00",X"03",X"0D",X"09",X"0A",X"0B",X"09",X"0A",X"0B",X"09",X"0C",X"0D",X"08",X"0C",X"04",X"00",
		X"00",X"03",X"0D",X"09",X"0C",X"0D",X"09",X"0A",X"0B",X"09",X"0A",X"02",X"07",X"05",X"06",X"00",
		X"00",X"03",X"0D",X"09",X"0A",X"0B",X"09",X"0A",X"0B",X"09",X"0C",X"04",X"07",X"05",X"06",X"00",
		X"00",X"03",X"0D",X"09",X"0A",X"0B",X"09",X"0A",X"0B",X"09",X"0C",X"04",X"07",X"05",X"06",X"00",
		X"00",X"05",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"0B",X"08",X"0C",X"04",X"00",
		X"00",X"05",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"06",X"00",X"05",X"06",X"00",
		X"00",X"05",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"06",X"00",X"05",X"06",X"00",
		X"00",X"03",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"0D",X"09",X"0C",X"04",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"0B",X"09",X"0A",X"02",X"00",X"01",X"0B",X"09",X"0A",X"02",X"00",
		X"00",X"01",X"0B",X"09",X"0C",X"04",X"07",X"01",X"0B",X"09",X"0C",X"04",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"0D",X"08",X"0A",X"02",X"07",X"01",X"0B",X"09",X"0A",X"02",X"00",
		X"00",X"01",X"0B",X"09",X"0C",X"04",X"07",X"03",X"0D",X"08",X"0C",X"04",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"0B",X"08",X"0C",X"04",X"00",X"03",X"0D",X"09",X"0A",X"02",X"00",
		X"00",X"01",X"0B",X"09",X"0C",X"04",X"00",X"03",X"0D",X"09",X"0C",X"04",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"0D",X"09",X"0A",X"02",X"07",X"01",X"0B",X"09",X"0A",X"02",X"00",
		X"00",X"01",X"0B",X"09",X"0C",X"04",X"07",X"03",X"0D",X"08",X"0C",X"04",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"0B",X"08",X"0A",X"02",X"07",X"03",X"0D",X"09",X"0A",X"02",X"00",
		X"00",X"01",X"0B",X"09",X"0C",X"04",X"00",X"03",X"0D",X"08",X"0C",X"04",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
