library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_SND_1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_SND_1 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"80",X"13",X"80",X"18",X"02",X"02",X"02",X"03",X"03",X"03",X"1D",X"0C",X"09",X"07",X"1E",X"00",
		X"00",X"00",X"19",X"5D",X"0C",X"5D",X"0C",X"5D",X"0C",X"07",X"28",X"00",X"03",X"81",X"0B",X"14",
		X"00",X"23",X"81",X"0B",X"15",X"00",X"25",X"81",X"0B",X"16",X"00",X"27",X"81",X"01",X"06",X"00",
		X"00",X"81",X"03",X"03",X"81",X"E8",X"21",X"67",X"07",X"19",X"D5",X"0A",X"F4",X"01",X"F9",X"01",
		X"18",X"01",X"01",X"01",X"01",X"01",X"01",X"1D",X"0A",X"09",X"09",X"1E",X"00",X"00",X"00",X"07",
		X"08",X"00",X"03",X"81",X"0B",X"FC",X"FF",X"23",X"81",X"0B",X"FE",X"FF",X"25",X"81",X"0B",X"FE",
		X"FF",X"27",X"81",X"01",X"03",X"03",X"81",X"EC",X"1A",X"D5",X"0A",X"F4",X"01",X"F9",X"01",X"1E",
		X"0A",X"09",X"09",X"07",X"76",X"00",X"03",X"81",X"0B",X"FC",X"FF",X"23",X"81",X"0B",X"FE",X"FF",
		X"25",X"81",X"0B",X"FE",X"FF",X"27",X"81",X"0B",X"FC",X"FF",X"31",X"81",X"0B",X"FE",X"FF",X"33",
		X"81",X"0B",X"FE",X"FF",X"35",X"81",X"01",X"03",X"03",X"81",X"DD",X"1D",X"00",X"00",X"00",X"07",
		X"08",X"00",X"03",X"81",X"0B",X"FC",X"FF",X"31",X"81",X"0B",X"FE",X"FF",X"33",X"81",X"0B",X"FE",
		X"FF",X"35",X"81",X"01",X"03",X"03",X"81",X"EC",X"21",X"67",X"07",X"19",X"FF",X"0F",X"00",X"02",
		X"80",X"00",X"1E",X"00",X"00",X"00",X"18",X"03",X"02",X"02",X"03",X"03",X"03",X"07",X"07",X"00",
		X"03",X"81",X"14",X"E9",X"08",X"0B",X"9C",X"FF",X"23",X"81",X"0B",X"EC",X"FF",X"25",X"81",X"0B",
		X"FB",X"FF",X"27",X"81",X"03",X"03",X"81",X"EA",X"10",X"1D",X"03",X"03",X"03",X"14",X"30",X"09",
		X"1D",X"05",X"08",X"03",X"14",X"30",X"09",X"1D",X"07",X"07",X"03",X"14",X"30",X"09",X"1D",X"07",
		X"06",X"03",X"14",X"30",X"09",X"1D",X"07",X"05",X"03",X"14",X"30",X"09",X"1D",X"06",X"03",X"06",
		X"14",X"30",X"09",X"1D",X"06",X"05",X"06",X"14",X"30",X"09",X"1D",X"03",X"03",X"06",X"14",X"30",
		X"09",X"1D",X"03",X"03",X"04",X"14",X"30",X"09",X"1D",X"03",X"03",X"04",X"14",X"30",X"09",X"15",
		X"07",X"0A",X"00",X"05",X"81",X"13",X"05",X"81",X"15",X"19",X"D5",X"06",X"F4",X"05",X"F9",X"03",
		X"1D",X"09",X"09",X"09",X"1E",X"00",X"00",X"00",X"07",X"3C",X"00",X"03",X"81",X"01",X"03",X"03",
		X"81",X"FB",X"21",X"67",X"07",X"19",X"12",X"00",X"15",X"00",X"20",X"00",X"1D",X"09",X"0B",X"09",
		X"1E",X"00",X"00",X"00",X"07",X"05",X"00",X"05",X"81",X"13",X"05",X"81",X"10",X"19",X"50",X"00",
		X"60",X"00",X"00",X"02",X"1D",X"09",X"0B",X"04",X"1E",X"00",X"00",X"00",X"07",X"05",X"00",X"05",
		X"81",X"13",X"05",X"81",X"10",X"18",X"02",X"02",X"02",X"02",X"02",X"02",X"06",X"1F",X"29",X"81",
		X"06",X"F7",X"2A",X"81",X"1D",X"10",X"00",X"00",X"06",X"38",X"2F",X"81",X"06",X"01",X"30",X"81",
		X"01",X"06",X"FF",X"05",X"81",X"01",X"03",X"05",X"81",X"FB",X"06",X"4F",X"05",X"81",X"01",X"03",
		X"05",X"81",X"FB",X"1D",X"00",X"00",X"00",X"01",X"21",X"67",X"07",X"18",X"03",X"03",X"03",X"03",
		X"03",X"03",X"19",X"FF",X"0F",X"FF",X"0F",X"FF",X"0F",X"1A",X"FF",X"0F",X"FF",X"0F",X"FF",X"0F",
		X"22",X"D5",X"09",X"16",X"10",X"08",X"A0",X"E4",X"09",X"B5",X"0A",X"69",X"0B",X"35",X"0C",X"B1",
		X"0C",X"2D",X"0D",X"06",X"01",X"80",X"01",X"C9",X"01",X"D4",X"01",X"C9",X"01",X"D1",X"02",X"D4",
		X"01",X"C8",X"01",X"D4",X"01",X"C8",X"01",X"CB",X"05",X"D4",X"01",X"80",X"01",X"C9",X"01",X"D4",
		X"01",X"C9",X"01",X"D1",X"02",X"D4",X"01",X"C8",X"01",X"D4",X"01",X"C8",X"01",X"CB",X"03",X"C4",
		X"01",X"80",X"01",X"C4",X"01",X"80",X"01",X"C9",X"01",X"CC",X"01",X"D5",X"01",X"80",X"01",X"D4",
		X"01",X"80",X"01",X"D4",X"01",X"80",X"01",X"C9",X"01",X"CC",X"01",X"D5",X"01",X"80",X"01",X"D4",
		X"02",X"80",X"01",X"80",X"01",X"A9",X"01",X"AC",X"01",X"B9",X"01",X"80",X"01",X"B9",X"01",X"BC",
		X"01",X"C9",X"01",X"80",X"01",X"C9",X"01",X"CC",X"01",X"D9",X"01",X"80",X"01",X"D9",X"01",X"DC",
		X"01",X"E9",X"02",X"E9",X"02",X"E9",X"02",X"E9",X"01",X"E9",X"01",X"E9",X"01",X"E9",X"01",X"E4",
		X"01",X"E6",X"01",X"E1",X"01",X"E4",X"02",X"E6",X"01",X"D9",X"01",X"D9",X"01",X"DB",X"01",X"DC",
		X"01",X"D9",X"01",X"DB",X"02",X"E1",X"01",X"E9",X"01",X"E1",X"01",X"D9",X"02",X"DB",X"02",X"D9",
		X"01",X"80",X"01",X"D9",X"02",X"D9",X"02",X"D9",X"02",X"D9",X"01",X"D9",X"01",X"D9",X"01",X"D9",
		X"01",X"D4",X"01",X"D6",X"01",X"D1",X"01",X"D4",X"02",X"D6",X"01",X"C9",X"01",X"C9",X"01",X"CB",
		X"01",X"CC",X"01",X"C9",X"01",X"CB",X"02",X"D1",X"01",X"C9",X"01",X"D1",X"01",X"C9",X"02",X"CB",
		X"02",X"C9",X"02",X"80",X"00",X"02",X"80",X"01",X"C4",X"02",X"80",X"02",X"C4",X"01",X"80",X"01",
		X"C4",X"01",X"C8",X"01",X"CB",X"05",X"C4",X"02",X"80",X"01",X"C4",X"02",X"80",X"02",X"C4",X"01",
		X"80",X"01",X"C4",X"01",X"C8",X"01",X"CB",X"03",X"C4",X"01",X"80",X"01",X"C4",X"03",X"80",X"01",
		X"C5",X"01",X"80",X"01",X"C4",X"01",X"80",X"01",X"C4",X"03",X"80",X"01",X"C5",X"01",X"80",X"01",
		X"C4",X"02",X"80",X"01",X"80",X"01",X"A9",X"01",X"AC",X"01",X"B9",X"01",X"80",X"01",X"B9",X"01",
		X"BC",X"01",X"C9",X"01",X"80",X"01",X"C9",X"01",X"CC",X"01",X"D9",X"01",X"80",X"01",X"D9",X"01",
		X"DC",X"01",X"E9",X"02",X"D9",X"02",X"D9",X"02",X"D9",X"01",X"D9",X"01",X"D9",X"01",X"D9",X"04",
		X"80",X"02",X"D9",X"01",X"D5",X"01",X"D5",X"01",X"80",X"01",X"D5",X"02",X"80",X"02",X"D4",X"01",
		X"80",X"01",X"D4",X"01",X"80",X"02",X"D4",X"02",X"D4",X"01",X"80",X"01",X"C9",X"02",X"C9",X"02",
		X"C9",X"02",X"C9",X"01",X"C9",X"01",X"C9",X"01",X"C9",X"01",X"80",X"01",X"C9",X"02",X"80",X"02",
		X"C9",X"01",X"C4",X"01",X"C5",X"01",X"80",X"01",X"C5",X"02",X"80",X"02",X"C4",X"01",X"80",X"01",
		X"C4",X"01",X"80",X"02",X"C4",X"02",X"C4",X"02",X"80",X"01",X"80",X"01",X"C9",X"01",X"D4",X"01",
		X"C9",X"01",X"D1",X"02",X"D4",X"01",X"C8",X"01",X"D4",X"01",X"C8",X"01",X"CB",X"05",X"D4",X"01",
		X"80",X"01",X"C9",X"01",X"D4",X"01",X"C9",X"01",X"D1",X"02",X"D4",X"01",X"C8",X"01",X"D4",X"01",
		X"C8",X"01",X"CB",X"03",X"C4",X"01",X"80",X"01",X"C4",X"01",X"80",X"01",X"C9",X"01",X"CC",X"01",
		X"D5",X"01",X"80",X"01",X"D4",X"01",X"80",X"01",X"D4",X"01",X"80",X"01",X"C9",X"01",X"CC",X"01",
		X"D5",X"01",X"80",X"01",X"D4",X"02",X"80",X"01",X"80",X"01",X"A9",X"01",X"AC",X"01",X"B9",X"01",
		X"80",X"01",X"B9",X"01",X"BC",X"01",X"C9",X"01",X"80",X"01",X"C9",X"01",X"CC",X"01",X"D9",X"01",
		X"80",X"01",X"D9",X"01",X"DC",X"01",X"E9",X"02",X"CC",X"02",X"CC",X"02",X"CC",X"02",X"CC",X"01",
		X"E9",X"01",X"E4",X"01",X"E6",X"01",X"E1",X"01",X"E4",X"02",X"E6",X"01",X"D9",X"01",X"D9",X"01",
		X"DB",X"01",X"DC",X"01",X"D9",X"01",X"DB",X"02",X"E1",X"01",X"E9",X"01",X"E1",X"01",X"D9",X"02",
		X"DB",X"02",X"D9",X"01",X"80",X"01",X"D9",X"02",X"BC",X"02",X"BC",X"02",X"BC",X"02",X"BC",X"01",
		X"D9",X"01",X"D4",X"01",X"D6",X"01",X"D1",X"01",X"D4",X"02",X"D6",X"01",X"C9",X"01",X"C9",X"01",
		X"CB",X"01",X"CC",X"01",X"C9",X"01",X"CB",X"02",X"D1",X"01",X"C9",X"01",X"D1",X"01",X"C9",X"02",
		X"CB",X"02",X"C9",X"02",X"80",X"02",X"B9",X"02",X"C1",X"02",X"C1",X"02",X"B9",X"02",X"BB",X"02",
		X"C2",X"02",X"C2",X"02",X"B4",X"02",X"B9",X"02",X"C1",X"02",X"C1",X"02",X"B9",X"02",X"BB",X"02",
		X"C2",X"02",X"C2",X"02",X"B4",X"04",X"B5",X"02",X"B4",X"02",X"B4",X"04",X"B5",X"02",X"B4",X"02",
		X"80",X"02",X"99",X"02",X"80",X"02",X"A9",X"02",X"80",X"02",X"B9",X"02",X"80",X"02",X"C9",X"02",
		X"80",X"02",X"C9",X"02",X"C9",X"02",X"C9",X"02",X"C9",X"02",X"D1",X"02",X"D1",X"02",X"D1",X"02",
		X"D1",X"02",X"CC",X"02",X"CC",X"02",X"D1",X"02",X"D1",X"02",X"D1",X"02",X"D2",X"02",X"D1",X"02",
		X"80",X"02",X"B9",X"02",X"B9",X"02",X"B9",X"02",X"B9",X"02",X"C1",X"02",X"C1",X"02",X"C1",X"02",
		X"C1",X"02",X"BC",X"02",X"BC",X"02",X"C1",X"02",X"C1",X"02",X"C1",X"02",X"C2",X"02",X"C1",X"02",
		X"80",X"02",X"A9",X"02",X"B9",X"02",X"B9",X"02",X"A9",X"02",X"AB",X"02",X"B8",X"02",X"B8",X"02",
		X"A4",X"02",X"A9",X"02",X"B9",X"02",X"B9",X"02",X"A9",X"02",X"AB",X"02",X"B8",X"02",X"B8",X"02",
		X"A4",X"04",X"A5",X"02",X"A4",X"02",X"A4",X"04",X"A5",X"02",X"A4",X"02",X"80",X"02",X"99",X"02",
		X"80",X"02",X"A9",X"02",X"80",X"02",X"B9",X"02",X"80",X"02",X"C9",X"02",X"80",X"02",X"C6",X"02",
		X"C6",X"02",X"C6",X"02",X"C6",X"02",X"C9",X"02",X"C9",X"02",X"C9",X"02",X"C9",X"02",X"C9",X"02",
		X"C9",X"02",X"C9",X"02",X"C9",X"02",X"C9",X"02",X"C8",X"02",X"C9",X"02",X"80",X"02",X"B6",X"02",
		X"B6",X"02",X"B6",X"02",X"B6",X"02",X"C9",X"02",X"C9",X"02",X"C9",X"02",X"C9",X"02",X"C9",X"02",
		X"C9",X"02",X"C9",X"02",X"C9",X"02",X"B9",X"02",X"B8",X"02",X"B9",X"02",X"A0",X"02",X"80",X"02",
		X"B4",X"02",X"B4",X"02",X"80",X"02",X"80",X"02",X"B4",X"02",X"B4",X"02",X"80",X"02",X"80",X"02",
		X"B4",X"02",X"B4",X"02",X"80",X"02",X"80",X"02",X"B4",X"02",X"B4",X"02",X"80",X"08",X"80",X"08",
		X"80",X"08",X"80",X"08",X"80",X"02",X"C3",X"02",X"C3",X"02",X"C3",X"02",X"C3",X"02",X"C4",X"02",
		X"C4",X"02",X"C4",X"02",X"C4",X"02",X"C5",X"02",X"C5",X"02",X"C4",X"02",X"C4",X"02",X"C4",X"02",
		X"C4",X"04",X"80",X"02",X"B3",X"02",X"B3",X"02",X"B3",X"02",X"B3",X"02",X"B4",X"02",X"B4",X"02",
		X"B4",X"02",X"B4",X"02",X"B5",X"02",X"B5",X"02",X"B4",X"02",X"B4",X"02",X"B4",X"02",X"B4",X"04",
		X"80",X"18",X"02",X"02",X"02",X"02",X"02",X"02",X"1A",X"FF",X"00",X"80",X"00",X"00",X"00",X"1E",
		X"08",X"08",X"00",X"07",X"0A",X"00",X"05",X"81",X"07",X"4F",X"01",X"03",X"81",X"01",X"03",X"03",
		X"81",X"FB",X"07",X"4F",X"01",X"03",X"81",X"0B",X"C0",X"FF",X"33",X"81",X"0B",X"C0",X"FF",X"31",
		X"81",X"01",X"03",X"03",X"81",X"FB",X"0B",X"40",X"00",X"33",X"81",X"0B",X"40",X"00",X"31",X"81",
		X"06",X"02",X"00",X"81",X"03",X"05",X"81",X"D0",X"10",X"18",X"03",X"03",X"03",X"03",X"03",X"03",
		X"06",X"00",X"00",X"81",X"19",X"FF",X"0F",X"FF",X"0F",X"FF",X"0F",X"1A",X"FF",X"0F",X"FF",X"0F",
		X"FF",X"0F",X"22",X"F8",X"0D",X"21",X"67",X"07",X"08",X"55",X"07",X"0E",X"12",X"0E",X"16",X"0E",
		X"1A",X"0E",X"1E",X"0E",X"22",X"0E",X"0A",X"02",X"C1",X"04",X"C3",X"02",X"BC",X"02",X"C1",X"06",
		X"C3",X"00",X"08",X"80",X"08",X"80",X"08",X"80",X"08",X"80",X"08",X"80",X"08",X"80",X"08",X"80",
		X"08",X"80",X"08",X"80",X"08",X"80",X"19",X"32",X"00",X"35",X"00",X"40",X"00",X"1D",X"09",X"0B",
		X"09",X"1E",X"00",X"00",X"00",X"07",X"2D",X"00",X"05",X"81",X"13",X"05",X"81",X"21",X"67",X"07",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
