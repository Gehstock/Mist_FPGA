library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity LLANDER_PROG_ROM_0 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of LLANDER_PROG_ROM_0 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"6B",X"20",X"13",X"62",X"A9",X"80",X"85",X"5D",X"24",X"97",X"30",X"0F",X"A9",X"00",X"85",X"22",
		X"85",X"97",X"24",X"5D",X"10",X"4C",X"20",X"13",X"62",X"D0",X"28",X"A5",X"22",X"D0",X"21",X"20",
		X"13",X"62",X"A9",X"F0",X"A2",X"08",X"20",X"5F",X"79",X"A2",X"00",X"86",X"23",X"86",X"A4",X"86",
		X"A5",X"A9",X"11",X"85",X"63",X"A9",X"20",X"A6",X"98",X"D0",X"01",X"4A",X"85",X"22",X"D0",X"03",
		X"20",X"35",X"62",X"20",X"A9",X"73",X"A2",X"2C",X"A0",X"CA",X"A5",X"21",X"F0",X"04",X"A2",X"A0",
		X"A0",X"C3",X"A5",X"22",X"29",X"20",X"F0",X"04",X"A2",X"00",X"A0",X"F0",X"8E",X"00",X"40",X"8C",
		X"01",X"40",X"A2",X"40",X"A0",X"04",X"A5",X"86",X"4A",X"90",X"04",X"A2",X"42",X"A0",X"84",X"86",
		X"28",X"84",X"27",X"A5",X"22",X"29",X"20",X"D0",X"2D",X"20",X"95",X"67",X"20",X"39",X"65",X"20",
		X"67",X"65",X"20",X"AD",X"65",X"A5",X"22",X"29",X"10",X"D0",X"1B",X"24",X"22",X"10",X"1D",X"A5",
		X"62",X"29",X"0F",X"F0",X"0B",X"A5",X"29",X"85",X"27",X"A5",X"2A",X"85",X"28",X"20",X"95",X"75",
		X"20",X"D6",X"68",X"4C",X"CE",X"60",X"20",X"7E",X"68",X"4C",X"CE",X"60",X"20",X"9D",X"66",X"24",
		X"22",X"50",X"18",X"A5",X"23",X"D0",X"0B",X"A5",X"86",X"29",X"0F",X"C9",X"08",X"D0",X"03",X"20",
		X"09",X"65",X"20",X"9E",X"68",X"20",X"FF",X"67",X"4C",X"CE",X"60",X"20",X"9F",X"79",X"A0",X"DE",
		X"A9",X"4B",X"A2",X"06",X"20",X"A6",X"7E",X"AD",X"00",X"20",X"29",X"02",X"F0",X"FE",X"20",X"2D",
		X"65",X"A0",X"02",X"A2",X"F0",X"A5",X"86",X"4A",X"90",X"04",X"A2",X"E1",X"A0",X"42",X"8E",X"03",
		X"40",X"8C",X"02",X"40",X"8D",X"00",X"30",X"E6",X"86",X"A2",X"00",X"AD",X"00",X"20",X"29",X"04",
		X"D0",X"02",X"A2",X"20",X"A9",X"1F",X"20",X"53",X"79",X"20",X"E6",X"62",X"20",X"14",X"64",X"24",
		X"22",X"30",X"37",X"50",X"1F",X"20",X"32",X"6B",X"20",X"3C",X"63",X"20",X"71",X"6B",X"20",X"1B",
		X"75",X"A5",X"01",X"C9",X"10",X"D0",X"02",X"A9",X"0F",X"4A",X"09",X"01",X"AA",X"A9",X"30",X"20",
		X"53",X"79",X"D0",X"0D",X"A9",X"20",X"A2",X"00",X"20",X"53",X"79",X"A5",X"22",X"29",X"20",X"D0",
		X"09",X"20",X"68",X"6C",X"20",X"4F",X"6D",X"20",X"1C",X"71",X"A5",X"22",X"F0",X"5B",X"20",X"AB",
		X"62",X"24",X"22",X"30",X"33",X"70",X"55",X"A2",X"00",X"A5",X"86",X"29",X"10",X"D0",X"02",X"A2",
		X"10",X"A9",X"0F",X"20",X"5F",X"79",X"2C",X"00",X"24",X"30",X"06",X"A9",X"40",X"85",X"25",X"D0",
		X"04",X"06",X"25",X"B0",X"0D",X"24",X"5D",X"10",X"0C",X"20",X"13",X"62",X"A9",X"10",X"85",X"22",
		X"D0",X"03",X"4C",X"40",X"60",X"4C",X"62",X"60",X"24",X"62",X"50",X"0E",X"24",X"5C",X"10",X"04",
		X"24",X"5D",X"30",X"06",X"20",X"68",X"6C",X"20",X"4F",X"6D",X"A5",X"86",X"4A",X"B0",X"E6",X"E6",
		X"56",X"10",X"E2",X"06",X"56",X"A5",X"62",X"85",X"5D",X"4C",X"08",X"60",X"A5",X"5D",X"30",X"28",
		X"20",X"AA",X"64",X"24",X"97",X"30",X"0C",X"A5",X"8D",X"C9",X"05",X"90",X"03",X"4C",X"01",X"60",
		X"4C",X"62",X"60",X"2C",X"05",X"24",X"30",X"06",X"A9",X"40",X"85",X"68",X"D0",X"F2",X"06",X"68",
		X"90",X"EE",X"A9",X"64",X"85",X"56",X"D0",X"E8",X"20",X"E0",X"6B",X"A5",X"5D",X"85",X"62",X"0A",
		X"D0",X"07",X"A0",X"00",X"A9",X"50",X"20",X"13",X"63",X"20",X"90",X"6B",X"20",X"94",X"76",X"A2",
		X"00",X"86",X"AF",X"86",X"B0",X"86",X"B1",X"A0",X"0A",X"96",X"57",X"88",X"10",X"FB",X"A9",X"20",
		X"20",X"53",X"79",X"06",X"22",X"A9",X"01",X"85",X"56",X"A9",X"0A",X"85",X"61",X"A9",X"41",X"85",
		X"63",X"D0",X"AD",X"8D",X"00",X"3E",X"A2",X"08",X"86",X"02",X"BD",X"0E",X"78",X"95",X"06",X"BD",
		X"B3",X"4B",X"95",X"0C",X"CA",X"D0",X"F3",X"86",X"60",X"86",X"61",X"A5",X"74",X"85",X"5F",X"A9",
		X"11",X"85",X"63",X"10",X"53",X"A5",X"74",X"29",X"03",X"85",X"33",X"18",X"69",X"01",X"29",X"03",
		X"85",X"34",X"A5",X"74",X"4A",X"4A",X"29",X"0F",X"C9",X"0F",X"D0",X"02",X"A9",X"04",X"20",X"9E",
		X"62",X"85",X"35",X"49",X"0F",X"20",X"9E",X"62",X"85",X"36",X"A2",X"03",X"BD",X"13",X"78",X"95",
		X"5E",X"BD",X"0F",X"78",X"95",X"07",X"BD",X"AE",X"55",X"95",X"11",X"CA",X"10",X"EE",X"A9",X"00",
		X"AA",X"A0",X"07",X"96",X"9C",X"88",X"10",X"FB",X"A9",X"40",X"85",X"22",X"A9",X"0F",X"20",X"5F",
		X"79",X"A9",X"10",X"85",X"02",X"20",X"BE",X"62",X"A2",X"00",X"A0",X"0E",X"96",X"4F",X"88",X"10",
		X"FB",X"CA",X"A0",X"07",X"96",X"79",X"88",X"10",X"FB",X"A9",X"40",X"85",X"4E",X"60",X"C9",X"04",
		X"B0",X"04",X"69",X"01",X"09",X"0A",X"60",X"11",X"11",X"22",X"11",X"2C",X"04",X"24",X"10",X"2D",
		X"06",X"24",X"90",X"2D",X"E6",X"23",X"A5",X"23",X"29",X"03",X"85",X"23",X"A5",X"02",X"0A",X"0A",
		X"85",X"67",X"A9",X"00",X"A2",X"03",X"95",X"03",X"CA",X"10",X"FB",X"85",X"66",X"A6",X"23",X"BD",
		X"A7",X"62",X"85",X"63",X"BD",X"E2",X"62",X"AA",X"A9",X"F0",X"4C",X"5F",X"79",X"A9",X"40",X"85",
		X"24",X"60",X"08",X"04",X"02",X"01",X"20",X"6B",X"79",X"D0",X"07",X"24",X"97",X"70",X"03",X"20",
		X"09",X"63",X"A6",X"B6",X"F0",X"05",X"C6",X"B6",X"20",X"09",X"63",X"A6",X"B8",X"F0",X"09",X"C6",
		X"B8",X"20",X"09",X"63",X"C6",X"99",X"D0",X"F9",X"60",X"A5",X"98",X"0A",X"AA",X"BD",X"2A",X"63",
		X"BC",X"2B",X"63",X"A2",X"FF",X"86",X"97",X"F8",X"18",X"65",X"AD",X"AA",X"98",X"65",X"AE",X"D8",
		X"90",X"03",X"A9",X"99",X"AA",X"85",X"AE",X"86",X"AD",X"60",X"00",X"09",X"50",X"04",X"00",X"06",
		X"50",X"07",X"00",X"09",X"00",X"11",X"00",X"13",X"50",X"15",X"00",X"18",X"A5",X"56",X"F0",X"01",
		X"60",X"A5",X"23",X"C9",X"03",X"F0",X"03",X"4C",X"D4",X"63",X"A5",X"66",X"18",X"65",X"03",X"85",
		X"66",X"A5",X"67",X"65",X"04",X"85",X"67",X"4A",X"4A",X"29",X"1F",X"85",X"02",X"A0",X"00",X"A5",
		X"03",X"A6",X"04",X"F0",X"0A",X"E8",X"D0",X"0B",X"C9",X"C0",X"90",X"07",X"88",X"30",X"04",X"C9",
		X"41",X"90",X"F9",X"84",X"05",X"24",X"97",X"10",X"5A",X"20",X"04",X"64",X"0A",X"0A",X"0A",X"0A",
		X"A0",X"00",X"29",X"F0",X"F0",X"25",X"90",X"01",X"88",X"18",X"65",X"03",X"AA",X"98",X"65",X"04",
		X"10",X"0A",X"C9",X"FC",X"B0",X"0E",X"A9",X"FC",X"A2",X"00",X"F0",X"08",X"C9",X"04",X"90",X"04",
		X"A9",X"03",X"A2",X"E0",X"85",X"04",X"86",X"03",X"4C",X"FE",X"63",X"A5",X"05",X"F0",X"1E",X"A5",
		X"06",X"F0",X"05",X"A9",X"00",X"AA",X"F0",X"11",X"A5",X"03",X"05",X"04",X"F0",X"0F",X"A9",X"50",
		X"A2",X"00",X"24",X"04",X"10",X"03",X"A9",X"B0",X"CA",X"86",X"04",X"85",X"03",X"A5",X"03",X"05",
		X"04",X"85",X"06",X"60",X"24",X"97",X"10",X"FB",X"20",X"04",X"64",X"F0",X"F6",X"18",X"65",X"67",
		X"85",X"67",X"AA",X"4A",X"4A",X"29",X"1F",X"85",X"02",X"A5",X"23",X"D0",X"11",X"E8",X"F0",X"06",
		X"E0",X"42",X"D0",X"0A",X"A9",X"10",X"85",X"02",X"0A",X"0A",X"85",X"67",X"90",X"D5",X"A2",X"00",
		X"A0",X"06",X"D0",X"5D",X"A2",X"00",X"2C",X"06",X"24",X"10",X"01",X"CA",X"2C",X"07",X"24",X"10",
		X"01",X"E8",X"8A",X"60",X"24",X"22",X"50",X"04",X"A5",X"56",X"D0",X"44",X"A5",X"84",X"4A",X"4A",
		X"AA",X"4A",X"85",X"37",X"A0",X"00",X"E4",X"82",X"B0",X"1A",X"A5",X"84",X"38",X"E5",X"82",X"A0",
		X"0F",X"90",X"11",X"C5",X"37",X"90",X"0D",X"A5",X"82",X"A4",X"84",X"20",X"C0",X"70",X"8A",X"4A",
		X"4A",X"4A",X"4A",X"A8",X"84",X"01",X"A0",X"00",X"A5",X"85",X"C9",X"4B",X"90",X"08",X"E6",X"83",
		X"C6",X"84",X"C6",X"84",X"84",X"85",X"24",X"97",X"10",X"04",X"A5",X"22",X"D0",X"02",X"84",X"01",
		X"60",X"A9",X"00",X"F8",X"85",X"39",X"86",X"38",X"84",X"37",X"A5",X"AC",X"38",X"E5",X"37",X"A8",
		X"A5",X"AD",X"E5",X"38",X"AA",X"A5",X"AE",X"E5",X"39",X"B0",X"14",X"24",X"97",X"10",X"29",X"A9",
		X"40",X"85",X"97",X"A9",X"00",X"85",X"AC",X"85",X"AD",X"85",X"AE",X"85",X"8D",X"F0",X"0A",X"84",
		X"AC",X"86",X"AD",X"85",X"AE",X"05",X"AD",X"F0",X"E2",X"18",X"A0",X"02",X"A2",X"00",X"B5",X"A1",
		X"75",X"37",X"95",X"A1",X"E8",X"88",X"10",X"F6",X"D8",X"60",X"A0",X"00",X"A5",X"56",X"F0",X"49",
		X"24",X"97",X"10",X"46",X"A5",X"86",X"4A",X"90",X"1A",X"A5",X"02",X"C9",X"08",X"90",X"0A",X"F0",
		X"12",X"C9",X"19",X"B0",X"04",X"C6",X"02",X"D0",X"07",X"18",X"69",X"01",X"29",X"1F",X"85",X"02",
		X"20",X"BC",X"62",X"A5",X"5F",X"D0",X"04",X"85",X"5E",X"F0",X"02",X"C6",X"5F",X"A5",X"02",X"C9",
		X"08",X"D0",X"16",X"A5",X"56",X"C9",X"3C",X"B0",X"0A",X"24",X"5C",X"30",X"06",X"A5",X"61",X"C9",
		X"10",X"B0",X"09",X"A9",X"10",X"85",X"01",X"C6",X"56",X"60",X"84",X"01",X"84",X"56",X"60",X"04",
		X"04",X"02",X"82",X"04",X"08",X"02",X"82",X"07",X"F0",X"A2",X"02",X"B5",X"5E",X"85",X"37",X"B5",
		X"5F",X"A0",X"05",X"4A",X"66",X"37",X"88",X"D0",X"FA",X"85",X"38",X"B5",X"5E",X"38",X"E5",X"37",
		X"95",X"5E",X"B5",X"5F",X"E5",X"38",X"95",X"5F",X"CA",X"CA",X"10",X"DF",X"60",X"46",X"73",X"90",
		X"FC",X"AD",X"00",X"20",X"4A",X"90",X"FA",X"60",X"2E",X"A5",X"4F",X"0A",X"85",X"8C",X"0A",X"85",
		X"8B",X"24",X"4E",X"70",X"0D",X"A9",X"E2",X"A2",X"51",X"20",X"D5",X"7E",X"A9",X"BA",X"A2",X"51",
		X"D0",X"0B",X"A9",X"BC",X"A2",X"4B",X"20",X"D5",X"7E",X"A9",X"F0",X"A2",X"44",X"A4",X"27",X"84",
		X"2D",X"A4",X"28",X"84",X"2E",X"D0",X"2B",X"24",X"4E",X"50",X"1C",X"A2",X"A1",X"20",X"9E",X"65",
		X"A9",X"FE",X"A2",X"52",X"20",X"92",X"65",X"24",X"22",X"70",X"01",X"60",X"A2",X"A3",X"20",X"9E",
		X"65",X"A9",X"0E",X"A2",X"53",X"D0",X"0B",X"A9",X"16",X"A2",X"54",X"20",X"D5",X"7E",X"A9",X"EE",
		X"A2",X"53",X"18",X"65",X"8C",X"A8",X"8A",X"69",X"00",X"A2",X"0A",X"4C",X"A6",X"7E",X"A9",X"00",
		X"85",X"37",X"85",X"39",X"85",X"3A",X"86",X"38",X"A0",X"37",X"4C",X"DC",X"7E",X"20",X"84",X"66",
		X"A0",X"0D",X"A9",X"00",X"85",X"3E",X"85",X"40",X"20",X"A4",X"7E",X"A5",X"27",X"85",X"29",X"A5",
		X"28",X"85",X"2A",X"A5",X"02",X"C9",X"09",X"B0",X"06",X"20",X"6E",X"66",X"4C",X"C9",X"7E",X"A2",
		X"04",X"A0",X"04",X"C6",X"3E",X"C6",X"40",X"C9",X"10",X"90",X"0E",X"C9",X"19",X"90",X"06",X"A2",
		X"00",X"E6",X"40",X"F0",X"08",X"29",X"0F",X"10",X"09",X"A0",X"00",X"E6",X"3E",X"20",X"F9",X"67",
		X"29",X"07",X"86",X"3D",X"84",X"3F",X"20",X"6E",X"66",X"84",X"37",X"85",X"38",X"A0",X"00",X"B1",
		X"37",X"0A",X"85",X"39",X"C8",X"B1",X"37",X"29",X"0F",X"09",X"20",X"2A",X"85",X"3A",X"24",X"4E",
		X"50",X"05",X"A5",X"39",X"18",X"90",X"18",X"88",X"B1",X"39",X"0A",X"85",X"64",X"C8",X"B1",X"39",
		X"29",X"0F",X"09",X"20",X"2A",X"85",X"65",X"20",X"37",X"66",X"A5",X"39",X"18",X"69",X"02",X"85",
		X"64",X"A5",X"3A",X"69",X"00",X"85",X"65",X"A0",X"00",X"B1",X"64",X"91",X"27",X"C8",X"B1",X"64",
		X"C9",X"A0",X"90",X"08",X"C9",X"F0",X"B0",X"17",X"88",X"4C",X"F8",X"74",X"45",X"3F",X"91",X"27",
		X"C8",X"B1",X"64",X"91",X"27",X"C8",X"B1",X"64",X"45",X"3D",X"91",X"27",X"C8",X"D0",X"DA",X"45",
		X"3F",X"91",X"27",X"88",X"B1",X"27",X"45",X"3D",X"91",X"27",X"C8",X"C8",X"D0",X"CB",X"0A",X"85",
		X"8B",X"24",X"4E",X"50",X"07",X"69",X"F4",X"A8",X"A9",X"4D",X"D0",X"05",X"69",X"A2",X"A8",X"A9",
		X"4B",X"69",X"00",X"60",X"A5",X"08",X"A6",X"07",X"20",X"EF",X"6C",X"85",X"10",X"84",X"0F",X"A5",
		X"0A",X"A6",X"09",X"20",X"EF",X"6C",X"84",X"0D",X"09",X"A0",X"85",X"0E",X"60",X"A5",X"01",X"F0",
		X"FB",X"A5",X"8B",X"24",X"4E",X"50",X"03",X"18",X"69",X"12",X"AA",X"BC",X"72",X"67",X"BD",X"71",
		X"67",X"24",X"3E",X"10",X"03",X"20",X"F9",X"67",X"85",X"3D",X"98",X"24",X"40",X"10",X"03",X"20",
		X"F9",X"67",X"85",X"3F",X"A5",X"01",X"A0",X"74",X"20",X"EF",X"70",X"A8",X"A5",X"86",X"4A",X"90",
		X"01",X"C8",X"A5",X"01",X"18",X"69",X"10",X"0A",X"0A",X"0A",X"90",X"02",X"A9",X"F0",X"85",X"8F",
		X"84",X"39",X"98",X"A4",X"3F",X"20",X"EF",X"70",X"86",X"3A",X"A5",X"3D",X"20",X"F9",X"67",X"A8",
		X"A5",X"39",X"20",X"EF",X"70",X"86",X"39",X"A5",X"3E",X"45",X"40",X"10",X"06",X"20",X"28",X"67",
		X"4C",X"09",X"67",X"20",X"09",X"67",X"4C",X"28",X"67",X"A0",X"00",X"A5",X"3A",X"18",X"65",X"3D",
		X"10",X"01",X"88",X"85",X"19",X"84",X"1A",X"A2",X"00",X"A5",X"39",X"18",X"65",X"3F",X"10",X"01",
		X"CA",X"85",X"1B",X"86",X"1C",X"4C",X"4A",X"67",X"A5",X"3A",X"20",X"F9",X"67",X"A2",X"00",X"18",
		X"65",X"3D",X"10",X"01",X"CA",X"85",X"19",X"86",X"1A",X"A5",X"39",X"20",X"F9",X"67",X"A2",X"00",
		X"18",X"65",X"3F",X"10",X"01",X"CA",X"85",X"1B",X"86",X"1C",X"A5",X"3E",X"45",X"40",X"10",X"1E",
		X"A5",X"19",X"F0",X"0B",X"20",X"F9",X"67",X"85",X"19",X"A5",X"1A",X"49",X"FF",X"85",X"1A",X"A5",
		X"1B",X"F0",X"0B",X"20",X"F9",X"67",X"85",X"1B",X"A5",X"1C",X"49",X"FF",X"85",X"1C",X"4C",X"43",
		X"78",X"00",X"F9",X"02",X"FA",X"03",X"FA",X"04",X"FB",X"05",X"FB",X"06",X"FC",X"06",X"FD",X"07",
		X"FE",X"07",X"00",X"00",X"FC",X"01",X"FC",X"01",X"FC",X"02",X"FD",X"03",X"FD",X"03",X"FE",X"04",
		X"FF",X"04",X"FF",X"04",X"00",X"A0",X"3C",X"A9",X"55",X"20",X"A4",X"7E",X"A9",X"A4",X"20",X"EB",
		X"67",X"A0",X"01",X"A9",X"9D",X"18",X"20",X"5A",X"7B",X"A2",X"02",X"20",X"AA",X"7E",X"A0",X"01",
		X"A9",X"9C",X"20",X"ED",X"67",X"A9",X"AD",X"20",X"EB",X"67",X"A9",X"AF",X"20",X"F4",X"67",X"20",
		X"D1",X"7E",X"A9",X"A6",X"20",X"F4",X"67",X"20",X"D1",X"7E",X"A9",X"A9",X"20",X"F4",X"67",X"A9",
		X"55",X"A0",X"AA",X"20",X"A4",X"7E",X"A5",X"9B",X"0A",X"69",X"60",X"20",X"E3",X"67",X"A5",X"9A",
		X"0A",X"69",X"5A",X"A8",X"A9",X"55",X"69",X"00",X"4C",X"C9",X"7E",X"A0",X"02",X"18",X"20",X"5A",
		X"7B",X"4C",X"D1",X"7E",X"A0",X"03",X"4C",X"59",X"7B",X"49",X"FF",X"18",X"69",X"01",X"60",X"A2");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
