//============================================================================
// 
//  Time Pilot '84 main PCB replica
//  Copyright (C) 2020 Ace
//
//  Permission is hereby granted, free of charge, to any person obtaining a
//  copy of this software and associated documentation files (the "Software"),
//  to deal in the Software without restriction, including without limitation
//  the rights to use, copy, modify, merge, publish, distribute, sublicense,
//  and/or sell copies of the Software, and to permit persons to whom the 
//  Software is furnished to do so, subject to the following conditions:
//
//  The above copyright notice and this permission notice shall be included in
//  all copies or substantial portions of the Software.
//
//  THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
//  IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
//  FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
//  AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
//  LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING
//  FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER
//  DEALINGS IN THE SOFTWARE.
//
//============================================================================

//Module declaration, I/O ports
module TimePilot84_CPU(
	input         reset,
	input         clk_49m, //Actual frequency: 49.152MHz
	output  [3:0] red, green, blue, //12-bit RGB, 4 bits per color
	output        video_hsync, video_vsync, video_csync, //CSync not needed for MISTer
	output        video_hblank, video_vblank,
	
	input   [7:0] sndbrd_D,
	output  [7:0] cpubrd_D,
	output        cpubrd_A5, cpubrd_A6,
	output        n_sda, n_son,
	output        in5, ioen,
	
	input         is_set3, //Flag to remap primary CPU address space for Time Pilot '84 Set 3
	output [15:0] main_cpu_rom_addr,
	input   [7:0] main_cpu_rom_do,	
	output [12:0] sub_cpu_rom_addr,
	input   [7:0] sub_cpu_rom_do,
	output [12:0] sp_rom_addr,
	input  [31:0] sp_rom_do
);

//Assign active high HBlank and VBlank outputs
assign video_hblank = hblk;
assign video_vblank = vblk;

//Output IN5, IOEN to sound board
assign in5 = n_in5;
assign ioen = n_ioen;

//Output primary MC6809E address lines A5 and A6 to sound board
assign cpubrd_A5 = mA[5];
assign cpubrd_A6 = mA[6];

//Assign CPU board data output to sound board
assign cpubrd_D = mD_out;

//------------------------------------------------- Abstracted logic modelling -------------------------------------------------//

/*Some of Time Pilot '84's original logic was found to be extremely unstable when using a 1:1 chip-level logic model. The result*/
/*of this was that the game would produce inconsistent visual errors every time this source code would be recompiled. The code  */
/*presented in this section of the CPU board model is an abstracted equivalent of the original logic adjusted to match the      */
/*timings of the signals generated by the original logic.                                                                       */
/*See the included PDF in the "docs" folder to learn more about the logic this section abstracts.                               */

//Partial abstraction of Time Pilot '84's primary CPU address decoding - this replaces the 74LS138 at 3A and half of the 74LS139
//at 7F.
//Time Pilot '84 (Set 3) has everything but its ROMs relocated to completely different locations in the primary MC6809E's address
//space - this abstraction includes extra logic using an external flag to remap the address space for this particular variant of
//the game.
wire n_mcpu_ram_en = is_set3 ? n_mcpu_ram_en_set3 : n_mcpu_ram_en_set1;
wire n_ioen = is_set3 ? ~((mA[15:4] == 12'h1A0 | mA[15:4] == 12'h1A2 | mA[15:4] == 12'h1A4 | mA[15:4] == 12'h1A6) & m_rw & meq):
                        ~((mA[15:4] == 12'h280 | mA[15:4] == 12'h282 | mA[15:4] == 12'h284 | mA[15:4] == 12'h286) & m_rw & meq);
wire n_in5 = is_set3 ? ~((mA[15:8] == 8'h1C) & m_rw & meq) : ~((mA[15:8] == 8'h30) & m_rw & meq);
wire n_latch_en = is_set3 ? ~((mA[15:8] == 8'h1C) & ~m_rw & meq) : ~((mA[15:8] == 8'h30) & ~m_rw & meq);
assign n_sda = is_set3 ? ~((mA[15:4] == 12'h1E8) & ~m_rw & meq) : ~((mA[15:8] == 8'h3A) & ~m_rw & meq);
assign n_son = is_set3 ? ~((mA[15:8] == 8'h1E) & ~m_rw & meq) : ~((mA[15:8] == 8'h38) & ~m_rw & meq);
wire xscroll_lat = is_set3 ? ~((mA[15:8] == 8'h1F) & ~m_rw & meq) : ~((mA[15:8] == 8'h3C) & ~m_rw & meq);
wire yscroll_lat = is_set3 ? ~((mA[15:4] == 12'h1F8) & ~m_rw & meq) : ~((mA[15:8] == 8'h3E) & ~m_rw & meq);
wire n_col0 = is_set3 ? ~((mA[15:8] == 8'h1A) & ~m_rw & meq) : ~((mA[15:8] == 8'h28) & ~m_rw & meq);
wire n_mafr = is_set3 ? ~((mA[15:8] == 8'h18) & ~m_rw & meq) : ~((mA[15:8] == 8'h20) & ~m_rw & meq);

//Signal to the video hardware when to draw the HUD - these signals are active when the horizontal counter is above 504 and below
//138 for the bottom HUD, and above 507 and below 284 for the top HUD.
//The PCB generates this signal by latching the signal used to enable the scroll registers (labelled scroll_lat in this
//implementation) on the falling edge of h2 (bit 1 of the horizontal counter) through the 74LS174 at 3G, then again latched twice
//through the 74LS377 at 2G on the rising edge of the pixel clock whenever the horizontal counter's 2 least significant bits are
//both set to 1 (this is the n_ld signal), first for the bottom HUD, then again for the top HUD.
wire bottom_hud_en = ({n_h256, h128, h64, h32, h16, h8, h4, h2, h1} > 504 || {n_h256, h128, h64, h32, h16, h8, h4, h2, h1} < 138);
wire top_hud_en = ({n_h256, h128, h64, h32, h16, h8, h4, h2, h1} > 507 || {n_h256, h128, h64, h32, h16, h8, h4, h2, h1} < 284);

//Generate HBlank (active high) while the horizontal counter is between 138 and 268
//While the Konami 082 custom chip generates VBlank, HBlank is generated externally using discrete logic, in this case, a
//combination of the 74LS74 at 4A and half of the 74LS74 at 4B
wire hblk = ({n_h256, h128, h64, h32, h16, h8, h4, h2, h1} > 137 && {n_h256, h128, h64, h32, h16, h8, h4, h2, h1} < 269);

//Output video signal from color PROMs, otherwise output black if in HBlank or VBlank
//This is normally achieved on the PCB by disabling the output of the 74LS157 at 3D when in HBlank and clearing the outputs of the
//74LS174 at 3C when in VBlank.
assign red = (hblk | vblk) ? 4'h0 : prom_red;
assign green = (hblk | vblk) ? 4'h0 : prom_green;
assign blue = (hblk | vblk) ? 4'h0 : prom_blue;

//------------------------------------------------- Chip-level logic modelling -------------------------------------------------//

//Konami 083 custom chip 1/2 - this one shifts the pixel data from character ROMs
k083 u1G
(
	.CK(clk2x),
	.LOAD(ld),
	.FLIP(charrom_flip),
	.DB0i(charrom_D),
	.DSH0(char_lut_A[1:0])
);

//Latch VCOL lines for character lookup PROM and color address bus bits A[6:4]
wire vcol0, vcol1;
ls174 u2B
(
	.d({1'b0, mD_out[3], mD_out[4], mD_out[2:0]}),
	.clk(n_col0),
	.mr(n_res),
	.q({1'bZ, vcol0, vcol1, color_A[6:4]})
);

//Latch SH and SF busses
wire [3:0] SH, SF;
ls273 u2E
(
	.d({SS, SH[0], SH[1], SH[2], SH[3]}),
	.clk(clk2x),
	.res(1'b1),
	.q({SH, SF[0], SF[1], SF[2], SF[3]})
);

//Latch S and SS busses
wire [3:0] S, SS;
ls273 u2F
(
	.d({S[0], S[1], S[2], S[3], char_lut_D}),
	.clk(clk2x),
	.res(1'b1),
	.q({SS[0], SS[1], SS[2], SS[3], S})
);

//Latch address lines A[5:2] for character lookup PROM, load for character ROM 083 custom chip
wire charrom_flip;
ls377 u2G
(
	.d({char_flip, 3'b000, charram1_Dl2}),
	.clk(clk2x),
	.e(n_ld),
	.q({charrom_flip, 3'bZZZ, char_lut_A[5:2]}) //Q[6:4] and D[6:4] would be responsible for generating the top
	                                            //and bottom HUD signals on the PCB
);

//Generate primary MC6809E VBlank IRQ clear and H/V flip signals
wire vrev, hrev, vblk_irq_clr;
ls259 u3B
(
	.d(mD_out[0]),
	.n_clr(n_res),
	.n_g(n_latch_en),
	.s(mA[2:0]),
	.q({2'bZZ, vrev, hrev, 3'bZZZ, vblk_irq_clr})
);

//Latch address lines A7 and A[3:0] for color PROMs, enable to draw bottom HUD
ls174 u3C
(
	.d({1'b0, char_spr_D[0], char_spr_D[2:1], char_spr_D[3], ch_sp_sel}), //D7 is the input to latch the bottom HUD enable signal
	.clk(clk2),
	.mr(1), //This is wired to the active-low VBlank output of the 082 custom chip, but is unnecessary with the abstracted handling of
	        //blanking in this implementation
	.q({1'bZ, color_A[0], color_A[2:1], color_A[3], color_A[7]}) //Bottom HUD enable is output from Q7
);

//Multiplex character and sprite data
wire [3:0] char_spr_D;
ls157 u3D
(
	.i0({sprite_D[0], sprite_D[2], sprite_D[3], sprite_D[1]}),
	.i1({char_D[0], char_D[2], char_D[3], char_D[1]}),
	.n_e(0), //The PCB clears this mux using HBlank, but this was found to cut a line off from the video output during testing and is
	         //abstracted instead
	.s(ch_sp_sel),
	.z({char_spr_D[0], char_spr_D[2], char_spr_D[3], char_spr_D[1]})
);

//Multiplex lower 2 bits of character data
wire [3:0] char_D;
ls153 u3E
(
	.i_a({S[0], SS[0], SH[0], SF[0]}),
	.i_b({S[1], SS[1], SH[1], SF[1]}),
	.n_e(2'b00),
	.s({char_sel1, char_sel0}),
	.z(char_D[1:0])
);

//Multiplex upper 2 bits of character data
ls153 u3F
(
	.i_a({S[2], SS[2], SH[2], SF[2]}),
	.i_b({S[3], SS[3], SH[3], SF[3]}),
	.n_e(2'b00),
	.s({char_sel1, char_sel0}),
	.z(char_D[3:2])
);

//Latch lowest 4 bits of already-latched character RAM data output
//The HUD signal would be latched from D[4] to Q[4] but has been omitted as this is part of the logic used to signal that the game is
//drawing the top and bottom HUDs, which has been abstracted
wire [3:0] charram1_Dl2;
ls174 u3G
(
	.d({2'b00, charram1_Dlat[3:0]}),
	.clk(n_h2),
	.mr(1'b1),
	.q({2'bZZ, charram1_Dl2})
);

//Latch address lines A[11:4] for character ROMs
ls273 u3H
(
	.d({charram0_Dlat[4], charram0_Dlat[5], charram0_Dlat[6], charram0_Dlat[7], charram0_Dlat[0], charram0_Dlat[1], charram0_Dlat[2], charram0_Dlat[3]}),
	.clk(n_h2),
	.res(1'b1),
	.q({charrom_A[8], charrom_A[9], charrom_A[10], charrom_A[11], charrom_A[4], charrom_A[5], charrom_A[6], charrom_A[7]})
);

//Generate lower 4 address lines for character ROMs
ls86 u3J
(
	.a1(ha2l),
	.b1(char_hflip),
	.y1(charrom_A[3]),
	.a2(va2l),
	.b2(char_vflip),
	.y2(charrom_A[1]),
	.a3(char_vflip),
	.b3(va1l),
	.y3(charrom_A[0]),
	.a4(va4l),
	.b4(char_vflip),
	.y4(charrom_A[2])
);

//The 74LS74s at 4A and 4B are part of the HBlank logic and logic to signal the game is drawing the bottom HUD - both are omitted
//as the signals have been abstracted
//See supplemental documentation included in the "docs" folder for more information

//Latch primary MC6809E data bus for Y scroll register (labelleed J and SHF1/SHF0 in the schematics)
wire [7:2] J;
wire shf0, shf1;
ls374 u4C
(
	.d({mD_out[3], mD_out[7], mD_out[0], mD_out[2], mD_out[6], mD_out[1], mD_out[5:4]}),
	.clk(xscroll_lat),
	.out_ctl(scroll_lat),
	.q({J[3], J[7], shf0, J[2], J[6], shf1, J[5:4]})
);

//Latch primary MC6809E data bus for X scroll register (labelled L in the schematics)
wire [7:0] L;
ls374 u4D
(
	.d({mD_out[2], mD_out[0], mD_out[3], mD_out[7], mD_out[4], mD_out[6:5], mD_out[1]}),
	.clk(yscroll_lat),
	.out_ctl(scroll_lat),
	.q({L[2], L[0], L[3], L[7], L[4], L[6:5], L[1]})
);

//Multiplex address lines A[3:0] for character RAM
ls157 u4E
(
	.i0({mA[2], mA[3], mA[1:0]}),
	.i1({ha[5], ha[6], ha[4:3]}),
	.n_e(1'b0),
	.s(n_h2),
	.z({charram_A[2], charram_A[3], charram_A[1:0]})
);

//Character RAM bank 1
wire [10:0] charram_A;
wire [7:0] charram1_D;
spram #(8, 11) u4F
(
	.clk(h1),
	.we(~n_charram1_we & ~n_charram1_en & n_charram_oe),
	.addr(charram_A),
	.data(mD_out),
	.q(charram1_D)
);

//Latch data output from character RAM bank 1
wire [7:0] charram1_Dlat;
ls273 u4G
(
	.d({charram1_D[7:6], charram1_D[4], charram1_D[5], charram1_D[3:0]}),
	.clk(h2),
	.res(1'b1),
	.q({charram1_Dlat[7:6], charram1_Dlat[4], charram1_Dlat[5], charram1_Dlat[3:0]})
);

//Latch data output from character RAM bank 0
wire [7:0] charram0_Dlat;
ls273 u4H
(
	.d({charram0_D[4], charram0_D[5], charram0_D[6], charram0_D[7], charram0_D[0], charram0_D[1], charram0_D[2], charram0_D[3]}),
	.clk(h2),
	.res(1'b1),
	.q({charram0_Dlat[4], charram0_Dlat[5], charram0_Dlat[6], charram0_Dlat[7], charram0_Dlat[0], charram0_Dlat[1], charram0_Dlat[2], charram0_Dlat[3]})
);

//Latch character ROM address lines A[3:0], character ROM address line A12, character ROM chip enable, character H/V flip bits
wire n_charrom0_ce, char_hflip, char_vflip, va1l, va2l, va4l, ha2l;
ls273 u4J
(
	.d({charram1_Dlat[5:4], charram1_Dlat[6], charram1_Dlat[7], va1, va2, va4, ha[2]}),
	.clk(n_h2),
	.res(1'b1),
	.q({n_charrom0_ce, charrom_A[12], char_hflip, char_vflip, va1l, va2l, va4l, ha2l})
);

//XOR horizontal counter bits [5:2] with HREV
wire h4x, h8x, h16x, h32x;
ls86 u5A
(
	.a1(h4),
	.b1(hrev),
	.y1(h4x),
	.a2(h16),
	.b2(hrev),
	.y2(h16x),
	.a3(hrev),
	.b3(h32),
	.y3(h32x),
	.a4(hrev),
	.b4(h8),
	.y4(h8x)
);

//XOR horizontal counter bits 6 and 7 with HREV, invert bit 3 of the horizontal counter and XOR 128H with !256H
wire h64x, h128x, h128_256, n_h8;
ls86 u5B
(
	.a1(h64),
	.b1(hrev),
	.y1(h64x),
	.a2(n_h256),
	.b2(h128),
	.y2(h128_256),
	.a3(h8),
	.b3(1'b0),
	.y3(n_h8),
	.a4(hrev),
	.b4(h128),
	.y4(h128x)
);

//Sum XORed horizontal counter bits [5:2] with X scroll register bits [5:2]
wire [7:2] ha;
wire ha_carry;
ls283 u5C
(
	.a({h32x, h16x, h8x, h4x}),
	.b(J[5:2]),
	.c_in(scroll_lat),
	.sum(ha[5:2]),
	.c_out(ha_carry)
);

//Sum XORed vertical counter bits [3:0] with Y scroll register bits [3:0]
wire va1, va2, va4, va8, va_carry;
ls283 u5D
(
	.a({v8x, v4x, v2x, v1x}),
	.b(L[3:0]),
	.c_in(scroll_lat),
	.sum({va8, va4, va2, va1}),
	.c_out(va_carry)
);

//Multiplex address lines A[7:4] for character RAM
ls157 u5E
(
	.i0({mA[6], mA[7], mA[5:4]}),
	.i1({va16, va32, va8, ha[7]}),
	.n_e(1'b0),
	.s(n_h2),
	.z({charram_A[6], charram_A[7], charram_A[5:4]})
);

//Character RAM bank 0
wire [7:0] charram0_D;
spram #(8, 11) u5F
(
	.clk(h1),
	.we(~n_charram0_we & ~n_charram0_en & n_charram_oe),
	.addr(charram_A),
	.data(mD_out),
	.q(charram0_D)
);

//Generate read enable lines for character RAM banks and chip enable for character RAM bank 0
wire charram0_rd, charram1_rd, n_charram0_en;
ls27 u5G
(
	.a1(n_m_rw),
	.b1(n_h2),
	.c1(n_vr2),
	.y1(charram1_rd),
	.a2(n_h2),
	.b2(n_m_rw),
	.c2(n_vr1),
	.y2(charram0_rd),
	.a3(charram0_we),
	.b3(charram0_rd),
	.c3(1'b0),
	.y3(n_charram0_en)
);

//5H and 5J are 74LS245s used to send data to/from character RAM and the primary MC6809E - not needed for this implementation

//Konami 082 custom chip - responsible for all video timings
wire vblk, h1, h2, h4, h8, h16, h32, h64, h128, n_h256, v1, v2, v4, v8, v16, v32, v64, v128;
k082 u6A
(
	.clk(pixel_clk),
	.n_vsync(video_vsync),
	.sync(video_csync),
	.n_hsync(video_hsync),
	.vblk(vblk),
	//The active-low VBlank output, n_vblk, is used by the PCB to clear the latch addressing the lower 4 bits of
	//the color PROMs at 3C but can be omitted from this implementation as blanking is handled differently to the PCB
	.h1(h1),
	.h2(h2),
	.h4(h4),
	.h8(h8),
	.h16(h16),
	.h32(h32),
	.h64(h64),
	.h128(h128),
	.n_h256(n_h256),
	.v1(v1),
	.v2(v2),
	.v4(v4),
	.v8(v8),
	.v16(v16),
	.v32(v32),
	.v64(v64),
	.v128(v128)
);

//Sum XORed horizontal counter bits [7:6] with X scroll register bits [7:6]
//Upper 2 adders unused, pull inputs low
ls283 u6C
(
	.a({2'b00, h128x, h64x}),
	.b({2'b00, J[7:6]}),
	.c_in(ha_carry),
	.sum({2'bZZ, ha[7:6]})
);

//Sum XORed vertical counter bits [7:4] with Y scroll register bits [7:4]
wire va16, va32, va64, va128;
ls283 u6D
(
	.a({v128x, v64x, v32x, v16x}),
	.b(L[7:4]),
	.c_in(va_carry),
	.sum({va128, va64, va32, va16})
);

//Multiplex address lines A[10:8] and output enable for character RAM
wire n_charram_oe;
ls157 u6E
(
	.i0({mA[10], n_m_rw, mA[9:8]}),
	.i1({scroll_lat, 1'b0, va128, va64}),
	.n_e(1'b0),
	.s(n_h2),
	.z({charram_A[10], n_charram_oe, charram_A[9:8]})
);

//Invert combined output enable signal for shared RAM, write enables for character RAM banks, read/write output from primary MC6809E,
//generate redundant CLK2
//Inverter 1 inverts the character ROM chip enable to select which of the two character ROMs to enable - this has been replaced with
//direct multiplexing
wire n_charram0_we, n_charram1_we, n_sharedram_oe, clk2x, n_m_rw;
ls04 u6F
(
	.a2(charram0_we),
	.y2(n_charram0_we),
	.a3(charram1_we),
	.y3(n_charram1_we),
	.a4(sharedram_oe),
	.y4(n_sharedram_oe),
	.a5(n_clk2),
	.y5(clk2x),
	.a6(m_rw),
	.y6(n_m_rw)
);

//Generate write enables for both character RAM banks and chip enable for character RAM bank 1
wire charram0_we, charram1_we, n_charram1_en;
ls27 u6G
(
	.a1(n_vr2),
	.b1(charram0_wr1),
	.c1(m_rw),
	.y1(charram1_we),
	.a2(charram1_we),
	.b2(charram1_rd),
	.c2(1'b0),
	.y2(n_charram1_en),
	.a3(charram0_wr1),
	.b3(n_vr1),
	.c3(m_rw),
	.y3(charram0_we)
);

//Latch vertical counter bits from 082 custom chip
wire [7:0] vcnt_lat;
ls273 u7B
(
	.d({v128, v64, v8, v4, v2, v1, v32, v16}),
	.clk(n_h256),
	.res(1'b1),
	.q({vcnt_lat[7:6], vcnt_lat[3:0], vcnt_lat[5:4]})
);

//XOR latched vertical counter bits [3:0] with VREV
wire v1x, v2x, v4x, v8x;
ls86 u7C
(
	.a1(vcnt_lat[1]),
	.b1(vrev),
	.y1(v2x),
	.a2(vcnt_lat[0]),
	.b2(vrev),
	.y2(v1x),
	.a3(vrev),
	.b3(vcnt_lat[3]),
	.y3(v8x),
	.a4(vrev),
	.b4(vcnt_lat[2]),
	.y4(v4x)
);

//XOR latched vertical counter bits [7:4] with VREV
wire v16x, v32x, v64x, v128x;
ls86 u7D
(
	.a1(vcnt_lat[5]),
	.b1(vrev),
	.y1(v32x),
	.a2(vcnt_lat[4]),
	.b2(vrev),
	.y2(v16x),
	.a3(vrev),
	.b3(vcnt_lat[7]),
	.y3(v128x),
	.a4(vrev),
	.b4(vcnt_lat[6]),
	.y4(v64x)
);

//Multiplex address lines A[3:0] for shared RAM
ls157 u7E
(
	.i0({mA[2], mA[3], mA[1:0]}),
	.i1({sA[2], sA[3], sA[1:0]}),
	.n_e(1'b0),
	.s(n_h2),
	.z({sharedram_A[2], sharedram_A[3], sharedram_A[1:0]})
);

//Generate write enables for sprite RAM
//The second half of this chip generates latch signals for X and Y scroll registers, sound data and IRQ triggers for the sound
//PCB - this can be ignored as the logic has been abstracted
wire n_spriteram0_we, n_spriteram1_we;
ls139 u7F
(
	.n_e({n_spriteram_dec_en, 1'b1}),
	.a0({sA[1], 1'b0}),
	.a1({sprram_en0, 1'b0}),
	.o1({n_spriteram0_we, n_spriteram1_we, 2'bZZ})
);

//Generate sprite RAM address line A8, write 1 for character RAM bank 0, sprite RAM decoder enable, enable for sprite RAM bank 1
wire charram0_wr1, n_spriteram_dec_en, sprram_en1;
ls32 u7G
(
	.a1(sA[9]),
	.b1(h2),
	.y1(spriteram_A[8]),
	.a2(n_h2),
	.b2(h1d),
	.y2(charram0_wr1),
	.a3(h2),
	.b3(n_ora),
	.y3(n_spriteram_dec_en),
	.a4(sprram_en0),
	.b4(s_rw),
	.y4(sprram_en1)
);

//Invert all clocks and bit 1 of the horizontal counter output from the 082 custom chip
//Gates 1 and 6 part of circuit to drive 18.432MHz crystal on the original PCB and gate 5
//inverts this clock, omit these gates
wire n_h2, clk1, clk2;
ls368 u8A
(
	.n_g1(0),
	.a2(h2),
	.y2(n_h2),
	.a3(n_clk2),
	.y3(clk2),
	.a4(n_clk1),
	.y4(clk1)
);

//Sprite RAM bank 0 (upper 4 bits)
wire [15:0] spriteram_D;
wire [9:0] spriteram_A;
spram #(4, 10) u8B
(
	.clk(pixel_clk),
	.we(~n_spriteram0_we & ~n_spriteram0_en),
	.addr(spriteram_A),
	.data(sD_out[7:4]),
	.q(spriteram_D[7:4])
);

//Sprite RAM bank 1 (upper 4 bits)
spram #(4, 10) u8C
(
	.clk(pixel_clk),
	.we(~n_spriteram1_we & ~n_spriteram1_en),
	.addr(spriteram_A),
	.data(sD_out[7:4]),
	.q(spriteram_D[15:12])
);

//Multiplex address lines A[3:0] for sprite RAM
ls157 u8D
(
	.i0({h32, h64, h16, h4}),
	.i1({sA[3], sA[4], sA[2], sA[0]}),
	.n_e(1'b0),
	.s(n_h2),
	.z({spriteram_A[2], spriteram_A[3], spriteram_A[1:0]})
);

//Multiplex address lines A[7:4] for shared RAM
ls157 u8E
(
	.i0({mA[6], mA[7], mA[5:4]}),
	.i1({sA[6], sA[7], sA[5:4]}),
	.n_e(1'b0),
	.s(n_h2),
	.z({sharedram_A[6], sharedram_A[7], sharedram_A[5:4]})
);

//Generate enable lines for shared RAM data bus multiplexing and LD0 signal for 502 custom chip
wire n_mcpu_sharedram_en, n_scpu_sharedram_en, n_ld0;
ls10 u8F
(
	.a1(n_h2),
	.b1(n_sharedram_rd),
	.c1(scr),
	.y1(n_scpu_sharedram_en),
	.a2(n_sharedram_rd),
	.b2(mcr),
	.c2(h2),
	.y2(n_mcpu_sharedram_en),
	.a3(h4),
	.b3(h2),
	.c3(h1),
	.y3(n_ld0)
);

//NAND shared RAM output enable with inverted latched H1 bit of horizontal counter, generate read
//enable for shared RAM and active-low LD signal, enable for watchdog timer reset
wire sharedram_h1, n_sharedram_rd, n_ld, watchdog_timer_rst;
ls00 u8G
(
	.a1(n_h1d),
	.b1(n_sharedram_oe),
	.y1(sharedram_h1),
	.a2(sharedram_h1),
	.b2(n_sharedram_oe),
	.y2(n_sharedram_rd),
	.a3(0), //Keep watchdog permanently disabled to prevent the risk of inappopriate resets or reset loops
	.b3(watchdog_timer_trig),
	.y3(watchdog_timer_rst),
	.a4(h1),
	.b4(h2),
	.y4(n_ld)
);

//Clock divider
//The PCB uses a 74LS107 located at 9A to divide 18.432MHz by 3 to obtain the required 6.144MHz pixel
//clock - this implementation replaces the 74LS107 by a 74LS163 to divide a faster 49.152MHz clock by
//4 for clocking PROMs and the sprite line buffer RAM at 12.288MHz and by 8 to obtain the 6.144MHz
//pixel clock
wire clk_12m, pixel_clk, n_clk1, n_clk2;
ls163 u9A
(
	.n_clr(1'b1),
	.clk(clk_49m),
	.din(4'h0),
	.enp(1'b1),
	.ent(1'b1),
	.n_load(1'b1),
	.q({1'bZ, pixel_clk, clk_12m, 1'bZ})
);
assign n_clk1 = ~pixel_clk;
assign n_clk2 = ~pixel_clk;

//Sprite RAM bank 0 (lower 4 bits)
spram #(4, 10) u9B
(
	.clk(pixel_clk),
	.we(~n_spriteram0_we & ~n_spriteram0_en),
	.addr(spriteram_A),
	.data(sD_out[3:0]),
	.q(spriteram_D[3:0])
);

//Sprite RAM bank 1 (lower 4 bits)
spram #(4, 10) u9C
(
	.clk(pixel_clk),
	.we(~n_spriteram1_we & ~n_spriteram1_en),
	.addr(spriteram_A),
	.data(sD_out[3:0]),
	.q(spriteram_D[11:8])
);

//Multiplex address lines A[7:4] for sprite RAM
ls157 u9D
(
	.i0({2'b11, h128, h128_256}),
	.i1({sA[7], sA[8], sA[6:5]}),
	.n_e(1'b0),
	.s(n_h2),
	.z({spriteram_A[6], spriteram_A[7], spriteram_A[5:4]})
);

//Multiplex output enable lines and address lines A[10:8] for shared RAM
wire sharedram_oe;
ls157 u9E
(
	.i0({mA[10], m_rw, mA[9:8]}),
	.i1({sA[10], s_rw, sA[9:8]}),
	.n_e(1'b0),
	.s(n_h2),
	.z({sharedram_A[10], sharedram_oe, sharedram_A[9:8]})
);

//Multplex data from CPUs to shared RAM (handled by the 74LS245s at 10G and 10F on the PCB)
wire [7:0] sharedram_Din = h2 ? mD_out : sD_out;

//Shared RAM for the two MC6809E CPUs
wire [10:0] sharedram_A;
wire [7:0] sharedram_D;
spram #(8, 11) u9F
(
	.clk(h1),
	.we(~n_sharedram_we),
	.addr(sharedram_A),
	.data(sharedram_Din),
	.q(sharedram_D)
);

//More address decoding for both MC6809Es (sprite RAM enables for secondary MC6809E, shared RAM
//and character RAM enables for primary MC6809E)
wire n_spriteram0_en, n_spriteram1_en, n_mcr, n_vr2, n_vr1;
ls139 u9G
(
	.n_e({n_mcpu_ram_en, n_spriteram_dec_en}),
	.a0({mA[11], sA[1]}),
	.a1({mA[12], sprram_en1}),
	.o0({n_spriteram0_en, n_spriteram1_en, 2'bZZ}),
	.o1({1'bZ, n_mcr, n_vr2, n_vr1})
);

//Konami 503 custom chip - generates sprite addresses for lower half of sprite ROMs, sprite
//data + collision control and enables for sprite write and 083 custom chip
wire csobj, k083_ctl, n_cara, n_ocoll;
k503 u11A
(
	.OB(spriteram_D[7:0]),
	.VCNT(vcnt_lat),
	.H4(h4),
	.H8(n_h8),
	.LD(n_ld),
	.OCS(csobj),
	.NE83(k083_ctl),
	.ODAT(n_cara),
	.OCOL(n_ocoll),
	.R(spriterom_A[5:0])
);

//Latch address lines A[12:6] and chip enables for sprite ROMs from sprite RAM bank 1
wire n_spriterom0_en;
ls273 u11C
(
	.d({spriteram_D[12], spriteram_D[13], spriteram_D[14], spriteram_D[15], spriteram_D[11:8]}),
	.clk(n_cara),
	.res(1'b1),
	.q({spriterom_A[10], spriterom_A[11], spriterom_A[12], n_spriterom0_en, spriterom_A[9:6]})
);

//11D is a 74LS244 used to buffer bits [12:5] of the address bus from the secondary MC6809E, not needed for this implementation

//11E is a 74LS367 used to buffer bits [4:0] of the address bus from the secondary MC6809E and its R/W signal, not needed for this
//implementation

//11F is a 74LS245 used to buffer the data bus from the secondary MC6809E, not needed for this implementation

//11G is a 74LS244 used to buffer bits [12:5] of the address bus from the primary MC6809E, not needed for this implementation

//11H is a 74LS367 used to buffer bits [4:0] of the address bus from the primary MC6809E and its R/W signal, not needed for this
//implementation

//11J is a 74LS245 used to buffer the data bus from the primary MC6809E, not needed for this implementation

//Generate upper half of sprite line buffer bank 0 address bus
ls163 u12C
(
	.n_clr(n_sprite_lbuff0_clr),
	.clk(clk2),
	.din(spriteram_D[15:12]),
	.enp(sprite_lbuff0_carry),
	.ent(sprite_lbuff0_carry),
	.n_load(n_sprite_lbuff0_ld),
	.q(sprite_lbuff0_A[7:4])
);

//Latch address lines A[7:4] for sprite lookup PROM, enable for sprite line buffer, XORed SHFx signals
//latch SCROLL again twice
wire shf0_l, shf1_l, sprite_lbuff_sel, sprrom_flip;
ls377 u12D
(
	.d({spriteram_D[3:0], shf0_rev, shf1_rev, csobj, k083_ctl}),
	.clk(clk2),
	.e(n_ocoll),
	.q({sprite_lut_A[7:4], shf0_l, shf1_l, sprite_lbuff_sel, sprrom_flip})
);

//Secondary CPU - Motorola MC6809E (uses modified version of John E. Kent's CPU09 by B. Cuzeau)
wire [15:0] sA;
wire [7:0] sD_out;
wire s_rw;
cpu09 u12E
(
	.clk(se),
	.ce(1),
	.rst(~n_res),
	.rw(s_rw),
	.addr(sA),
	.data_in(sD_in),
	.data_out(sD_out),
	.halt(0),
	.irq(~n_sirq),
	.firq(0),
	.nmi(0)
);
//Multiplex data inputs to secondary MC6809E
wire [7:0] sD_in =
		~n_rom5_en                         ? sub_cpu_rom_do:
//		~n_rom5_en                         ? eprom5_D:
		~n_scpu_sharedram_en               ? sharedram_D:
		~n_spriteram1_en & n_spriteram1_we ? spriteram_D[15:8]:
		~n_spriteram0_en & n_spriteram0_we ? spriteram_D[7:0]:
		~n_beam_en                         ? vcnt_lat:
		8'hFF;

//Primary CPU - Motorola MC6809E (uses modified version of John E. Kent's CPU09 by B. Cuzeau)
wire [15:0] mA;
wire [7:0] mD_out;
wire m_rw;
cpu09 u12G
(
	.clk(me),
	.ce(1),
	.rst(~n_res),
	.rw(m_rw),
	.addr(mA),
	.data_in(mD_in),
	.data_out(mD_out),
	.halt(0),
	.irq(~n_mirq),
	.firq(0),
	.nmi(0)
);
//Multiplex data inputs to primary MC6809E
wire [7:0] mD_in =
		sndbrd_dir                       ? sndbrd_D:
		(~n_charram0_en & ~n_charram_oe) ? charram0_D:
		(~n_charram1_en & ~n_charram_oe) ? charram1_D:
		~n_mcpu_sharedram_en             ? sharedram_D:
//		~n_rom1_en                       ? eprom1_D:
//		~n_rom2_en                       ? eprom2_D:
//		~n_rom3_en                       ? eprom3_D:
//		~n_rom4_en                       ? eprom4_D:
		~n_rom1_en                       ? main_cpu_rom_do:
		~n_rom2_en                       ? main_cpu_rom_do:
		~n_rom3_en                       ? main_cpu_rom_do:
		~n_rom4_en                       ? main_cpu_rom_do:
		8'hFF;

//Address decoding for primary MC6809E (1/2)
wire n_rom1_en, n_rom2_en, n_rom3_en, n_rom4_en, n_mcpu_ram_en_set1, n_mcpu_ram_en_set3;
ls138 u12J
(
	.n_e1(1'b0),
	.n_e2(1'b0),
	.e3(meq),
	.a(mA[15:13]),
	//o[0] is usually unused and o[1] is chained into the 74LS138 at 3A for further address decoding.
	//o[0] is used here at it spans the entire address space taking up by shared RAM and character RAM
	//for Time Pilot '84 (Set 3).
	.o({n_rom4_en, n_rom3_en, n_rom2_en, n_rom1_en, 1'bZ, n_mcpu_ram_en_set1, 1'bZ, n_mcpu_ram_en_set3})
);

//Generate lower half of sprite line buffer bank 0 address bus
wire sprite_lbuff0_carry;
ls163 u13C
(
	.n_clr(n_sprite_lbuff0_clr),
	.clk(clk2),
	.din(spriteram_D[11:8]),
	.enp(1'b1),
	.ent(1'b1),
	.n_load(n_sprite_lbuff0_ld),
	.q(sprite_lbuff0_A[3:0]),
	.rco(sprite_lbuff0_carry)
);

//Sprite line buffer bank 0
wire [7:0] sprite_lbuff0_A;
wire [3:0] sprite_lbuff0_D;
spram #(4, 10) u13D
(
	.clk(clk_12m),
	.we(~clk2 & ~n_sprite_lbuff0_en),
	.addr({2'b00, sprite_lbuff0_A}),
	.data(sprite_lbuff_Do[3:0]),
	.q(sprite_lbuff0_D)
);

//Address decoding for secondary MC6809E
wire n_rom5_en, n_scr, n_ora, n_scpu_irq, n_beam_en, n_safr;
ls138 u13E
(
	.n_e1(1'b0),
	.n_e2(1'b0),
	.e3(seq),
	.a(sA[15:13]),
	.o({n_rom5_en, 2'bZZ, n_scr, n_ora, n_scpu_irq, n_beam_en, n_safr})
);

//Invert E and Q clocks for secondary MC6809E, MCR and SCR
//Inverter 5 inverts the chip enable for sprite ROMs - this is not required here and has
//been omitted
wire scr, se, sq, ld, mcr;
ls04 u13F
(
	.a1(n_scr),
	.y1(scr),
	.a2(n_sq),
	.y2(sq),
	.a3(n_se),
	.y3(se),
	.a4(n_ld),
	.y4(ld),
	.a6(n_mcr),
	.y6(mcr)
);

//NAND horizontal counter bits [6:4], sound board direction signal, watchdog timer + power-on reset
wire res, n_h32_128, sndbrd_dir;
ls10 u13G
(
	.a1(h32),
	.b1(h128),
	.c1(h64),
	.y1(n_h32_128),
	.a2(1), //This is usually connected to !IN6, which is a signal that serves no real purpose on the PCB
	.b2(n_ioen),
	.c2(n_in5),
	.y2(sndbrd_dir),
	.a3(n_watchdog_timer),
	.b3(n_por_timer_out),
	.c3(reset),
	.y3(res)
);

//Invert reset line for the entire PCB, E and Q clocks for primary MC6809E, power-on reset timer output,
//watchdog timer output
wire n_res, me, mq, sprite_lbuff_h, n_por_timer_out, n_watchdog_timer;
ls04 u13H
(
	.a1(res),
	.y1(n_res),
	.a2(n_me),
	.y2(me),
	.a3(n_mq),
	.y3(mq),
	.a4(sprite_lbuff_l),
	.y4(sprite_lbuff_h),
	.a5(por_timer_out),
	.y5(n_por_timer_out),
	.a6(watchdog_timer),
	.y6(n_watchdog_timer)
);

//Generate the following signals:
//VBlank IRQ for primary MC6809E, latch for scrolling/static screen area
wire n_mirq, scroll_lat;
ls74 u13J
(
	.n_pre1(vblk_irq_clr),
	.n_clr1(1'b1),
	.clk1(vblk),
	.d1(1'b0),
	.q1(n_mirq),
	.n_pre2(1'b1),
	.n_clr2(1'b1),
	.clk2(h16),
	.d2(scroll),
	.n_q2(scroll_lat)
);

//Generate upper half of sprite line buffer bank 1 address bus
ls163 u14C
(
	.n_clr(n_sprite_lbuff1_clr),
	.clk(clk2),
	.din(spriteram_D[15:12]),
	.enp(sprite_lbuff1_carry),
	.ent(sprite_lbuff1_carry),
	.n_load(n_sprite_lbuff1_ld),
	.q(sprite_lbuff1_A[7:4])
);

//Sprite line buffer bank 1
wire [7:0] sprite_lbuff1_A;
wire [3:0] sprite_lbuff1_D;
spram #(4, 10) u14D
(
	.clk(clk_12m),
	.we(~clk2 & ~n_sprite_lbuff1_en),
	.addr({2'b00, sprite_lbuff1_A}),
	.data(sprite_lbuff_Do[7:4]),
	.q(sprite_lbuff1_D)
);

//Invert H256 signal for Konami 502, XOR shf0 and shf1 with inverted HREV, generate character flip signal
wire shf1_rev, h256, char_flip, shf0_rev;
ls86 u14E
(
	.a1(shf1),
	.b1(n_hrev),
	.y1(shf1_rev),
	.a2(n_h256),
	.b2(0),
	.y2(h256),
	.a3(n_hrev),
	.b3(char_hflip),
	.y3(char_flip),
	.a4(n_hrev),
	.b4(shf0),
	.y4(shf0_rev)
);

//Generate VBlank interrupt and clear signal for secondary MC6809E
wire n_sirq, s_vblk_irq_clr;
ls74 u14F
(
	.n_pre1(s_vblk_irq_clr),
	.n_clr1(1),
	.clk1(vblk),
	.d1(0),
	.q1(n_sirq),
	.n_pre2(1),
	.n_clr2(n_res),
	.clk2(n_scpu_irq),
	.d2(sD_out[0]),
	.q2(s_vblk_irq_clr)
);

//Generate E and Q clocks for both MC6809Es
wire n_me, n_mq, n_se, n_sq;
ls74 u14G
(
	.n_pre1(1),
	.n_clr1(1),
	.clk1(clk2),
	.d1(h2),
	.q1(n_mq),
	.n_q1(n_sq),
	.n_pre2(1),
	.n_clr2(1),
	.clk2(clk2),
	.d2(n_mq),
	.q2(n_me),
	.n_q2(n_se)
);

//Watchdog timer
wire watchdog_timer_fb, watchdog_timer;
ls293 u14H
(
	.clk1(vblk),
	.clk2(watchdog_timer_fb),
	.clr1(watchdog_timer_rst),
	.clr2(watchdog_timer_rst),
	.q({watchdog_timer, 2'bZZ, watchdog_timer_fb})
);

//Latch least significant bit of horizontal counter, latch for watchdog timer
wire h1d, n_h1d, watchdog_lat;
ls74 u14J
(
	.n_pre1(1),
	.n_clr1(1),
	.clk1(n_clk1),
	.d1(h1),
	.q1(h1d),
	.n_q1(n_h1d),
	.n_pre2(watchdog_lat_pre),
	.n_clr2(n_res),
	.clk2(n_safr),
	.d2(watchdog_safr),
	.q2(watchdog_lat)
);

//Generate lower half of sprite line buffer bank 1 address bus
wire sprite_lbuff1_carry;
ls163 u15C
(
	.n_clr(n_sprite_lbuff1_clr),
	.clk(clk2),
	.din(spriteram_D[11:8]),
	.enp(1),
	.ent(1),
	.n_load(n_sprite_lbuff1_ld),
	.q(sprite_lbuff1_A[3:0]),
	.rco(sprite_lbuff1_carry)
);

//Konami 502 custom chip, responsible for generating sprites (sits between sprite ROMs and the sprite line buffer)
wire [7:0] sprite_lbuff_Do;
wire [4:0] sprite_D;
wire sprite_lbuff_l, sprite_lbuff_dec0, sprite_lbuff_dec1;
k502 u15D
(
	.CK1(clk1),
	.CK2(k502_ck2),
	.LD0(n_ld0),
	.H2(h2),
	.H256(h256),
	.SPAL(sprite_lut_D),
	.SPLBi({sprite_lbuff1_D, sprite_lbuff0_D}),
	.SPLBo(sprite_lbuff_Do),
	.OSEL(sprite_lbuff_l),
	.OLD(sprite_lbuff_dec1),
	.OCLR(sprite_lbuff_dec0),
	.COL(sprite_D)
);

//Generate inverted HREV signal, background mux select signals, sprite RAM write select signal
wire n_hrev, vmux0, vmux1, sprram_en0;
ls02 u15F
(
	.a1(hrev),
	.b1(0),
	.y1(n_hrev),
	.a2(shf1_l),
	.b2(top_hud_en),
	.y2(vmux1),
	.a3(shf0_l),
	.b3(top_hud_en),
	.y3(vmux0),
	.a4(s_rw),
	.b4(h1d),
	.y4(sprram_en0)
);

//Generate character data select lines, combined EQ clocks for each CPU
wire char_sel0, char_sel1, meq, seq;
ls32 u15G
(
	.a1(vmux1),
	.b1(bottom_hud_en),
	.y1(char_sel1),
	.a2(n_sq),
	.b2(n_se),
	.y2(meq),
	.a3(n_me),
	.b3(n_mq),
	.y3(seq),
	.a4(bottom_hud_en),
	.b4(vmux0),
	.y4(char_sel0)
);

//15H contains an NE555 timer which takes approximately 326ms to pull the board out of reset.  Model this as a
//32-bit counter that pulls the core out of reset when its value reaches 1998221
reg [31:0] por_timer = 0;
always_ff @(posedge pixel_clk) begin
	if(por_timer < 1998221)
		por_timer <= por_timer + 1;
end
wire por_timer_out = (por_timer < 1998220);

//Generate watchdog latch preset, watchdog timer trigger, sprite RAM address line A9, watchdog latch SAFR input
wire watchdog_lat_pre, watchdog_timer_trig, watchdog_safr;
ls32 u15J
(
	.a1(n_sq),
	.b1(n_mafr),
	.y1(watchdog_lat_pre),
	.a2(n_mafr),
	.b2(watchdog_lat),
	.y2(watchdog_timer_trig),
	.a3(sA[10]),
	.b3(h2),
	.y3(spriteram_A[9]),
	.a4(0),
	.b4(n_safr),
	.y4(watchdog_safr)
);

//Konami 083 custom chip 2/2 - this one shifts the pixel data from sprite ROMs
k083 u16A
(
	.CK(clk2),
	.LOAD(ld),
	.FLIP(sprrom_flip),
	.DB0i(spriterom_D[7:0]),
	.DB1i(spriterom_D[15:8]),
	.DSH0(sprite_lut_A[1:0]),
	.DSH1(sprite_lut_A[3:2])
);

//Generate load and clear signals for 74LS163s generating addresses for sprite line buffer
wire n_sprite_lbuff0_ld, n_sprite_lbuff1_ld, n_sprite_lbuff0_clr, n_sprite_lbuff1_clr;
ls139 u16D
(
	.n_e({n_ld, n_ocoll}),
	.a0({sprite_lbuff_dec0, sprite_lbuff_dec1}),
	.a1({sprite_lbuff_dec1, 1'b0}),
	.o0({2'bZZ, n_sprite_lbuff1_ld, n_sprite_lbuff0_ld}),
	.o1({1'bZ, n_sprite_lbuff0_clr, n_sprite_lbuff1_clr, 1'bZ})
);

//Generate clock for 502 custom chip, select line for character/sprite MUX, color MUX enable
wire k502_ck2, ch_sp_sel, n_sharedram_we, color_mux;
ls32 u16E
(
	.a1(1'b0),
	.b1(clk2),
	.y1(k502_ck2),
	.a2(sprite_D[4]),
	.b2(color_mux),
	.y2(ch_sp_sel),
	.a3(sharedram_en),
	.b3(sharedram_h1),
	.y3(n_sharedram_we),
	.a4(top_hud_en),
	.b4(bottom_hud_en),
	.y4(color_mux)
);

//Generate combined shared RAM enable, sprite line buffer enables, scroll data to be latched
wire sharedram_en, n_sprite_lbuff0_en, n_sprite_lbuff1_en, scroll;
ls08 u16F
(
	.a1(n_mcpu_sharedram_en),
	.b1(n_scpu_sharedram_en),
	.y1(sharedram_en),
	.a2(sprite_lbuff_l),
	.b2(sprite_lbuff_sel),
	.y2(n_sprite_lbuff0_en),
	.a3(sprite_lbuff_h),
	.b3(sprite_lbuff_sel),
	.y3(n_sprite_lbuff1_en),
	.a4(n_h256),
	.b4(n_h32_128),
	.y4(scroll)
);


//ROMs
//Primary CPU ROM
/*
wire [7:0] eprom1_D;
wire [7:0] eprom2_D;
wire [7:0] eprom3_D;
wire [7:0] eprom4_D;
wire [7:0] eprom5_D;


cpu1_rom u7J(
	.clk(mq),
	.addr(mA[12:0]),
	.data(eprom1_D)
);

cpu2_rom u8J(
	.clk(mq),
	.addr(mA[12:0]),
	.data(eprom2_D)
);

cpu3_rom u9J(
	.clk(mq),
	.addr(mA[12:0]),
	.data(eprom3_D)
);

cpu4_rom u10J(
	.clk(mq),
	.addr(mA[12:0]),
	.data(eprom4_D)
);*/

assign main_cpu_rom_addr = mA[15:0];

//Secondary CPU ROM
/*
sub_rom u10D(
	.clk(sq),
	.addr(sA[12:0]),
	.data(eprom5_D)
);*/
assign sub_cpu_rom_addr = sA[12:0];

//Character ROM
//Multiplex character and sprite ROM data outputs.
//The PCB connects these signals directly to the chip enable signals on the EPROMs at 2J (character) and 12A/13A (sprite) and
//invert them through one inverter at 6F (character) and 13F (sprite) for the second set of character ROMs (3J) and sprite
//ROMs (14A/15A).
wire [7:0] charrom_D =  ~n_charrom0_ce ? eprom7_D : eprom8_D;
wire [12:0] charrom_A;
wire [7:0] eprom7_D;
wire [7:0] eprom8_D;
char_rom1 u2J(
	.clk(pixel_clk),
	.addr(charrom_A),
	.data(eprom7_D)
);

char_rom2 u1J(
	.clk(pixel_clk),
	.addr(charrom_A),
	.data(eprom8_D)
);

//Sprite ROM
//wire [15:0] spriterom_D = ~n_spriterom0_en ? {eprom11_D, eprom9_D} : {eprom12_D, eprom10_D};
assign sp_rom_addr = spriterom_A;
wire [15:0] spriterom_D =  ~n_spriterom0_en ? sp_rom_do[15:0] : sp_rom_do[31:16];

//Sprite ROM 1/4
wire [12:0] spriterom_A;
//wire [7:0] eprom9_D;
//wire [7:0] eprom10_D;
//wire [7:0] eprom11_D;
//wire [7:0] eprom12_D;
/*
spr_rom1  u12A(
	.clk(pixel_clk),
	.addr(spriterom_A),
	.data(eprom9_D)
);

spr_rom2  u13A(
	.clk(pixel_clk),
	.addr(spriterom_A),
	.data(eprom10_D)
);

spr_rom3  u14A(
	.clk(pixel_clk),
	.addr(spriterom_A),
	.data(eprom11_D)
);

spr_rom4  u15A(
	.clk(pixel_clk),
	.addr(spriterom_A),
	.data(eprom12_D)
);*/

//PROMS
//Color
wire [7:0] color_A;
wire [3:0] prom_red;
wire [3:0] prom_green;
wire [3:0] prom_blue;
pal_r u2C(
	.clk(clk_12m),
	.addr(color_A),
	.data(prom_red)
);

pal_g u2D(
	.clk(clk_12m),
	.addr(color_A),
	.data(prom_green)
);

pal_b u1E(
	.clk(clk_12m),
	.addr(color_A),
	.data(prom_blue)
);

//Character lookup PROM
wire [5:0] char_lut_A;
wire [3:0] char_lut_D;
char_lut u1F(
	.clk(clk_12m),
	.addr({vcol1, vcol0, char_lut_A}),
	.data(char_lut_D)
);

//Sprite lookup PROM
wire [7:0] sprite_lut_A;
wire [3:0] sprite_lut_D;
sprite_lut u16C(
	.clk(clk_12m),
	.addr(sprite_lut_A),
	.data(sprite_lut_D)
);

endmodule
