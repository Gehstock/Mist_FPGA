library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity MoonWar_program1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of MoonWar_program1 is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"F3",X"AF",X"D3",X"4D",X"ED",X"47",X"DB",X"61",X"CB",X"47",X"C2",X"00",X"02",X"DB",X"60",
		X"CB",X"47",X"C2",X"65",X"06",X"DD",X"21",X"5D",X"01",X"18",X"68",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"D3",X"4D",X"F5",X"3A",X"00",X"40",X"B7",X"C2",X"1D",X"05",
		X"F1",X"C3",X"0B",X"1B",X"07",X"00",X"F8",X"B9",X"00",X"01",X"00",X"00",X"0D",X"20",X"FD",X"10",
		X"FB",X"DB",X"66",X"3E",X"01",X"01",X"41",X"01",X"11",X"47",X"82",X"ED",X"41",X"0D",X"ED",X"51",
		X"0C",X"0C",X"ED",X"41",X"0C",X"ED",X"41",X"0C",X"0C",X"0C",X"ED",X"59",X"0E",X"51",X"3D",X"28",
		X"EA",X"01",X"00",X"00",X"0D",X"20",X"FD",X"10",X"FB",X"DB",X"67",X"AF",X"D3",X"40",X"D3",X"50",
		X"DD",X"E9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"18",X"3B",X"01",X"C0",X"08",X"21",X"00",X"00",X"16",X"08",X"7E",X"09",X"AF",X"ED",X"4F",X"32",
		X"00",X"10",X"15",X"20",X"F5",X"0E",X"7F",X"16",X"20",X"7B",X"E6",X"20",X"47",X"ED",X"78",X"CB",
		X"0B",X"0D",X"15",X"20",X"F4",X"3E",X"80",X"01",X"57",X"80",X"ED",X"79",X"05",X"0D",X"CB",X"0F",
		X"30",X"F8",X"0E",X"47",X"ED",X"79",X"0D",X"CB",X"0F",X"30",X"F9",X"18",X"C5",X"3E",X"01",X"ED",
		X"47",X"AF",X"01",X"00",X"10",X"86",X"23",X"0D",X"C2",X"45",X"01",X"10",X"F8",X"FE",X"FF",X"C2",
		X"55",X"01",X"1C",X"DD",X"E9",X"ED",X"57",X"A7",X"C2",X"02",X"01",X"18",X"FE",X"1E",X"00",X"21",
		X"00",X"00",X"DD",X"21",X"69",X"01",X"C3",X"41",X"01",X"21",X"00",X"10",X"DD",X"21",X"73",X"01",
		X"C3",X"41",X"01",X"21",X"00",X"20",X"DD",X"21",X"7D",X"01",X"C3",X"41",X"01",X"21",X"00",X"30",
		X"DD",X"21",X"87",X"01",X"C3",X"41",X"01",X"21",X"00",X"C0",X"DD",X"21",X"91",X"01",X"C3",X"41",
		X"01",X"DD",X"21",X"98",X"01",X"C3",X"79",X"00",X"2A",X"75",X"00",X"ED",X"4B",X"77",X"00",X"36",
		X"55",X"2B",X"ED",X"A1",X"E2",X"AA",X"01",X"23",X"18",X"F5",X"16",X"AA",X"31",X"FF",X"FF",X"ED",
		X"4B",X"77",X"00",X"7A",X"2F",X"AE",X"20",X"16",X"72",X"2B",X"ED",X"A1",X"EA",X"CB",X"01",X"7A",
		X"FE",X"55",X"28",X"25",X"31",X"01",X"00",X"16",X"55",X"18",X"E4",X"39",X"18",X"E5",X"57",X"ED",
		X"57",X"CB",X"0F",X"38",X"01",X"76",X"1E",X"12",X"7A",X"E6",X"0F",X"CA",X"02",X"01",X"1D",X"7A",
		X"E6",X"F0",X"CA",X"02",X"01",X"1D",X"C3",X"02",X"01",X"ED",X"57",X"CB",X"0F",X"1E",X"20",X"D2",
		X"B1",X"02",X"C3",X"02",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"01",X"48",X"10",X"ED",X"78",X"0C",X"ED",X"78",X"0C",X"ED",X"78",X"0C",X"0C",X"ED",X"78",X"0C",
		X"ED",X"78",X"0C",X"ED",X"78",X"0C",X"3E",X"01",X"ED",X"79",X"01",X"48",X"00",X"ED",X"78",X"0C",
		X"ED",X"78",X"0C",X"ED",X"78",X"21",X"00",X"50",X"11",X"00",X"70",X"06",X"10",X"78",X"3D",X"D3",
		X"4B",X"3E",X"80",X"77",X"12",X"4E",X"CB",X"0F",X"30",X"F9",X"AF",X"DB",X"4E",X"3E",X"08",X"32",
		X"00",X"50",X"32",X"00",X"70",X"AF",X"DB",X"4E",X"23",X"13",X"10",X"E1",X"06",X"0D",X"11",X"00",
		X"A0",X"21",X"FE",X"5F",X"3E",X"80",X"25",X"77",X"4E",X"24",X"37",X"CB",X"15",X"CB",X"14",X"19",
		X"CB",X"0F",X"10",X"F2",X"21",X"11",X"11",X"11",X"11",X"11",X"31",X"00",X"88",X"0E",X"10",X"06",
		X"10",X"E5",X"E5",X"E5",X"E5",X"10",X"FA",X"19",X"F1",X"3B",X"3B",X"0D",X"20",X"F1",X"DB",X"4C",
		X"AF",X"DB",X"4E",X"AF",X"DB",X"61",X"E6",X"02",X"28",X"FE",X"21",X"00",X"50",X"11",X"00",X"70",
		X"3E",X"F0",X"ED",X"47",X"01",X"4B",X"00",X"ED",X"57",X"ED",X"79",X"0E",X"00",X"79",X"70",X"12",
		X"48",X"2F",X"46",X"47",X"B1",X"20",X"F6",X"ED",X"57",X"D6",X"10",X"ED",X"47",X"20",X"E5",X"18",
		X"FE",X"DD",X"21",X"B8",X"02",X"C3",X"79",X"00",X"21",X"FF",X"5F",X"11",X"00",X"00",X"DD",X"21",
		X"C5",X"02",X"C3",X"95",X"03",X"01",X"00",X"00",X"21",X"00",X"40",X"DD",X"21",X"D2",X"02",X"C3",
		X"76",X"03",X"21",X"00",X"40",X"11",X"55",X"00",X"DD",X"21",X"DF",X"02",X"C3",X"95",X"03",X"21",
		X"FF",X"5F",X"11",X"AA",X"55",X"DD",X"21",X"EC",X"02",X"C3",X"95",X"03",X"21",X"00",X"40",X"11",
		X"FF",X"AA",X"DD",X"21",X"F9",X"02",X"C3",X"95",X"03",X"21",X"FF",X"5F",X"11",X"00",X"FF",X"DD",
		X"21",X"06",X"03",X"C3",X"95",X"03",X"79",X"B0",X"C2",X"C1",X"03",X"DD",X"21",X"12",X"03",X"C3",
		X"79",X"00",X"21",X"FF",X"87",X"11",X"00",X"00",X"DD",X"21",X"1F",X"03",X"C3",X"95",X"03",X"01",
		X"00",X"00",X"21",X"00",X"80",X"DD",X"21",X"2C",X"03",X"C3",X"76",X"03",X"21",X"00",X"84",X"DD",
		X"21",X"36",X"03",X"C3",X"76",X"03",X"21",X"00",X"80",X"11",X"55",X"00",X"DD",X"21",X"43",X"03",
		X"C3",X"8F",X"03",X"21",X"FF",X"87",X"11",X"AA",X"55",X"DD",X"21",X"50",X"03",X"C3",X"8F",X"03",
		X"21",X"00",X"80",X"11",X"FF",X"AA",X"DD",X"21",X"5D",X"03",X"C3",X"8F",X"03",X"21",X"FF",X"87",
		X"11",X"00",X"FF",X"DD",X"21",X"6A",X"03",X"C3",X"8F",X"03",X"79",X"B0",X"C2",X"6C",X"03",X"DD",
		X"21",X"42",X"04",X"C3",X"79",X"00",X"16",X"00",X"72",X"7E",X"AA",X"B0",X"47",X"23",X"72",X"7E",
		X"AA",X"B1",X"4F",X"2B",X"15",X"C2",X"78",X"03",X"36",X"00",X"23",X"36",X"00",X"DD",X"E9",X"D9",
		X"01",X"00",X"08",X"18",X"04",X"D9",X"01",X"00",X"20",X"D9",X"7E",X"AA",X"B0",X"47",X"73",X"7E",
		X"AB",X"B0",X"47",X"CB",X"43",X"C2",X"AA",X"03",X"2B",X"3E",X"23",X"78",X"41",X"4F",X"D9",X"0D",
		X"C2",X"B7",X"03",X"05",X"CA",X"BB",X"03",X"D9",X"C3",X"9A",X"03",X"D9",X"78",X"41",X"4F",X"DD",
		X"E9",X"21",X"22",X"04",X"11",X"01",X"00",X"78",X"A2",X"C2",X"E8",X"03",X"79",X"A3",X"C3",X"E8",
		X"03",X"EB",X"29",X"EB",X"D2",X"C7",X"03",X"11",X"00",X"40",X"1D",X"FD",X"7E",X"00",X"C2",X"DA",
		X"03",X"15",X"C2",X"DA",X"03",X"C3",X"B8",X"02",X"08",X"7E",X"23",X"D9",X"6F",X"D9",X"7E",X"23",
		X"D9",X"67",X"11",X"1F",X"00",X"06",X"03",X"08",X"B7",X"28",X"07",X"36",X"FC",X"23",X"36",X"3F",
		X"18",X"05",X"36",X"84",X"23",X"36",X"21",X"19",X"10",X"EE",X"06",X"24",X"B7",X"28",X"07",X"36",
		X"FF",X"23",X"36",X"FF",X"18",X"05",X"36",X"80",X"23",X"36",X"01",X"19",X"10",X"EE",X"D9",X"C3",
		X"D1",X"03",X"8D",X"50",X"4D",X"4A",X"0D",X"44",X"CD",X"56",X"15",X"44",X"55",X"4A",X"95",X"50",
		X"D5",X"56",X"89",X"50",X"49",X"4A",X"09",X"44",X"C9",X"56",X"11",X"44",X"51",X"4A",X"91",X"50",
		X"D1",X"56",X"21",X"00",X"60",X"16",X"01",X"42",X"AF",X"4F",X"5F",X"ED",X"47",X"ED",X"57",X"D3",
		X"4B",X"36",X"FF",X"72",X"36",X"00",X"7E",X"BB",X"20",X"FE",X"ED",X"57",X"3C",X"ED",X"47",X"FE",
		X"10",X"20",X"0B",X"CB",X"12",X"30",X"E0",X"DD",X"21",X"87",X"04",X"C3",X"79",X"00",X"79",X"CB",
		X"1F",X"CB",X"18",X"CB",X"19",X"59",X"ED",X"57",X"FE",X"08",X"38",X"D1",X"3E",X"08",X"CB",X"08",
		X"CB",X"13",X"3D",X"20",X"F9",X"18",X"C6",X"1E",X"00",X"DD",X"21",X"CA",X"04",X"21",X"00",X"60",
		X"01",X"01",X"01",X"7B",X"D3",X"4B",X"78",X"32",X"00",X"40",X"71",X"79",X"DD",X"E9",X"AE",X"20",
		X"FE",X"77",X"78",X"A1",X"28",X"02",X"3E",X"80",X"57",X"DB",X"4E",X"AA",X"17",X"38",X"FE",X"CB",
		X"00",X"30",X"E0",X"CB",X"01",X"30",X"DC",X"DD",X"23",X"DD",X"23",X"DD",X"23",X"3E",X"10",X"83",
		X"5F",X"30",X"D0",X"DD",X"21",X"FA",X"04",X"C3",X"79",X"00",X"00",X"18",X"D1",X"B0",X"18",X"CE",
		X"2F",X"18",X"18",X"AF",X"18",X"21",X"A0",X"18",X"C5",X"78",X"18",X"C2",X"A8",X"18",X"18",X"2F",
		X"18",X"EB",X"2F",X"18",X"0F",X"A8",X"18",X"B6",X"78",X"18",X"0C",X"A0",X"18",X"09",X"AF",X"18",
		X"AD",X"2F",X"18",X"E2",X"B0",X"18",X"00",X"2F",X"18",X"A4",X"ED",X"5E",X"3E",X"07",X"ED",X"47",
		X"DD",X"21",X"85",X"1A",X"3E",X"FF",X"D3",X"4F",X"47",X"31",X"FF",X"43",X"DB",X"4E",X"1F",X"CB",
		X"10",X"78",X"EE",X"55",X"28",X"03",X"FB",X"18",X"FE",X"D3",X"4F",X"06",X"FF",X"31",X"FF",X"43",
		X"DB",X"4D",X"DB",X"4E",X"1F",X"CB",X"10",X"78",X"EE",X"20",X"CA",X"79",X"00",X"DB",X"4C",X"18",
		X"FE",X"AF",X"D3",X"4F",X"DB",X"4E",X"31",X"40",X"40",X"DB",X"65",X"CB",X"7F",X"20",X"FA",X"CD",
		X"65",X"1E",X"CD",X"DE",X"CB",X"F3",X"21",X"F8",X"05",X"7E",X"B7",X"CA",X"85",X"1A",X"CD",X"C6",
		X"05",X"06",X"00",X"11",X"00",X"CF",X"CD",X"E4",X"05",X"CD",X"C6",X"05",X"E5",X"5E",X"23",X"56",
		X"23",X"46",X"23",X"E5",X"21",X"00",X"00",X"E5",X"E5",X"E5",X"39",X"CD",X"9F",X"05",X"11",X"CF",
		X"00",X"CD",X"B9",X"05",X"E1",X"E1",X"E1",X"E1",X"E3",X"DB",X"65",X"CB",X"7F",X"20",X"16",X"DB",
		X"48",X"CB",X"7F",X"20",X"F4",X"E5",X"5E",X"23",X"56",X"23",X"46",X"AF",X"12",X"13",X"10",X"FC",
		X"E1",X"D1",X"C3",X"5C",X"05",X"E1",X"DB",X"65",X"CB",X"7F",X"20",X"FA",X"C3",X"49",X"05",X"E5",
		X"D5",X"C5",X"1A",X"13",X"E6",X"F0",X"4F",X"1A",X"13",X"07",X"07",X"07",X"07",X"E6",X"0F",X"B1",
		X"77",X"23",X"05",X"10",X"ED",X"C1",X"D1",X"E1",X"C9",X"C5",X"D5",X"E5",X"53",X"1E",X"00",X"CD",
		X"A0",X"2F",X"E1",X"D1",X"C1",X"C9",X"C5",X"D5",X"E5",X"01",X"C0",X"19",X"11",X"00",X"44",X"21",
		X"00",X"46",X"ED",X"B0",X"01",X"00",X"02",X"AF",X"12",X"13",X"0D",X"C2",X"D8",X"05",X"10",X"F8",
		X"E1",X"D1",X"C1",X"C9",X"EB",X"CD",X"68",X"2F",X"EB",X"4E",X"CD",X"EE",X"2F",X"13",X"23",X"47",
		X"7E",X"B7",X"78",X"C2",X"E9",X"05",X"23",X"C9",X"43",X"72",X"65",X"64",X"69",X"74",X"73",X"00",
		X"BA",X"F8",X"02",X"43",X"68",X"75",X"74",X"65",X"20",X"31",X"00",X"BC",X"F8",X"08",X"43",X"68",
		X"75",X"74",X"65",X"20",X"32",X"00",X"C4",X"F8",X"08",X"43",X"68",X"75",X"74",X"65",X"20",X"33",
		X"00",X"CC",X"F8",X"08",X"50",X"6C",X"61",X"79",X"73",X"00",X"D4",X"F8",X"06",X"54",X"6F",X"74",
		X"61",X"6C",X"20",X"53",X"63",X"6F",X"72",X"65",X"00",X"DA",X"F8",X"0C",X"54",X"6F",X"74",X"61",
		X"6C",X"20",X"53",X"65",X"63",X"6F",X"6E",X"64",X"73",X"20",X"6F",X"66",X"20",X"50",X"6C",X"61",
		X"79",X"00",X"E6",X"F8",X"0C",X"48",X"69",X"67",X"68",X"20",X"53",X"63",X"6F",X"72",X"65",X"73",
		X"00",X"F2",X"F8",X"06",X"00",X"31",X"86",X"F8",X"CD",X"65",X"1E",X"CD",X"99",X"CB",X"21",X"ED",
		X"06",X"11",X"20",X"00",X"CD",X"C5",X"06",X"11",X"20",X"80",X"CD",X"C5",X"06",X"11",X"08",X"10",
		X"CD",X"C5",X"06",X"11",X"10",X"D0",X"CD",X"C5",X"06",X"21",X"A0",X"47",X"CD",X"5C",X"1E",X"21",
		X"A0",X"55",X"CD",X"5C",X"1E",X"11",X"08",X"20",X"DB",X"61",X"CD",X"CB",X"06",X"DB",X"60",X"CD",
		X"CB",X"06",X"DB",X"62",X"CD",X"CB",X"06",X"DB",X"63",X"CD",X"CB",X"06",X"DB",X"64",X"CD",X"CB",
		X"06",X"11",X"08",X"90",X"DB",X"48",X"CD",X"CA",X"06",X"DB",X"49",X"CD",X"CA",X"06",X"DB",X"4A",
		X"CD",X"CA",X"06",X"18",X"D0",X"06",X"00",X"C3",X"E4",X"05",X"2F",X"0E",X"08",X"21",X"35",X"07",
		X"1F",X"38",X"03",X"21",X"37",X"07",X"F5",X"D5",X"C5",X"CD",X"C5",X"06",X"C1",X"D1",X"F1",X"21",
		X"20",X"00",X"19",X"EB",X"0D",X"20",X"E6",X"21",X"00",X"0F",X"19",X"EB",X"C9",X"5A",X"50",X"55",
		X"20",X"44",X"49",X"50",X"20",X"53",X"57",X"49",X"54",X"43",X"48",X"45",X"53",X"00",X"56",X"46",
		X"42",X"20",X"53",X"57",X"49",X"54",X"43",X"48",X"45",X"53",X"00",X"31",X"20",X"20",X"20",X"32",
		X"20",X"20",X"20",X"33",X"20",X"20",X"20",X"34",X"20",X"20",X"20",X"35",X"20",X"20",X"20",X"36",
		X"20",X"20",X"20",X"37",X"20",X"20",X"20",X"38",X"00",X"30",X"3D",X"4F",X"46",X"46",X"20",X"20",
		X"7F",X"3D",X"4F",X"4E",X"00",X"7F",X"00",X"30",X"00",X"78",X"21",X"00",X"44",X"54",X"5D",X"36",
		X"01",X"23",X"73",X"23",X"01",X"FD",X"1B",X"EB",X"ED",X"B0",X"21",X"00",X"45",X"54",X"5D",X"06",
		X"20",X"36",X"FF",X"23",X"10",X"FB",X"01",X"80",X"02",X"09",X"EB",X"01",X"7F",X"18",X"ED",X"B0",
		X"CD",X"99",X"CB",X"CD",X"86",X"07",X"21",X"00",X"44",X"11",X"01",X"44",X"01",X"FF",X"1B",X"36",
		X"FF",X"ED",X"B0",X"21",X"00",X"81",X"11",X"01",X"81",X"01",X"FF",X"06",X"36",X"11",X"ED",X"B0",
		X"CD",X"86",X"07",X"C3",X"3A",X"07",X"DB",X"49",X"CB",X"47",X"20",X"FA",X"DB",X"49",X"CB",X"47",
		X"28",X"FA",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"09",X"05",X"17",X"05",
		X"00",X"9D",X"12",X"5C",X"08",X"CD",X"13",X"01",X"48",X"08",X"5C",X"08",X"CD",X"13",X"02",X"D1",
		X"15",X"5C",X"08",X"CD",X"13",X"03",X"6F",X"14",X"C8",X"19",X"66",X"1A",X"04",X"72",X"08",X"5C",
		X"08",X"CD",X"13",X"05",X"79",X"15",X"5C",X"08",X"CD",X"13",X"06",X"A9",X"15",X"C8",X"19",X"66",
		X"1A",X"07",X"13",X"15",X"5C",X"08",X"CD",X"13",X"08",X"86",X"10",X"BA",X"10",X"5E",X"12",X"09",
		X"D0",X"13",X"5C",X"08",X"CD",X"13",X"FF",X"FF",X"2C",X"13",X"2C",X"13",X"37",X"13",X"37",X"13",
		X"4C",X"13",X"4C",X"13",X"41",X"13",X"41",X"13",X"00",X"00",X"48",X"08",X"57",X"13",X"6D",X"13",
		X"57",X"13",X"6D",X"13",X"81",X"13",X"97",X"13",X"B1",X"13",X"B1",X"13",X"CD",X"13",X"00",X"00",
		X"6C",X"08",X"34",X"14",X"38",X"14",X"3D",X"14",X"43",X"14",X"4A",X"14",X"52",X"14",X"65",X"14",
		X"65",X"14",X"00",X"00",X"7E",X"08",X"02",X"0F",X"04",X"40",X"0C",X"60",X"14",X"50",X"24",X"48",
		X"44",X"44",X"84",X"42",X"84",X"42",X"FC",X"7E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"0F",X"06",X"00",X"0A",X"20",X"12",X"30",X"24",X"48",
		X"44",X"44",X"84",X"42",X"84",X"42",X"7C",X"7A",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"0F",X"06",X"00",X"0A",X"20",X"12",X"30",X"22",X"28",
		X"42",X"24",X"84",X"42",X"FC",X"42",X"00",X"42",X"00",X"3E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"0F",X"07",X"00",X"09",X"20",X"12",X"30",X"22",X"28",
		X"42",X"24",X"82",X"22",X"7C",X"42",X"00",X"42",X"00",X"7A",X"00",X"06",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"0F",X"07",X"80",X"08",X"80",X"11",X"10",X"21",X"18",
		X"42",X"24",X"62",X"22",X"1C",X"42",X"00",X"42",X"00",X"42",X"00",X"32",X"00",X"0C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"0F",X"07",X"C0",X"08",X"40",X"10",X"80",X"21",X"08",
		X"42",X"14",X"32",X"22",X"0C",X"22",X"00",X"42",X"00",X"62",X"00",X"12",X"00",X"0C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"0F",X"07",X"C0",X"08",X"40",X"10",X"80",X"21",X"08",
		X"22",X"14",X"1A",X"12",X"04",X"22",X"00",X"42",X"00",X"42",X"00",X"22",X"00",X"14",X"00",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"0F",X"07",X"C0",X"08",X"40",X"10",X"40",X"20",X"80",
		X"11",X"0C",X"0A",X"12",X"04",X"22",X"00",X"42",X"00",X"42",X"00",X"42",X"00",X"24",X"00",X"18",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"0F",X"07",X"C0",X"08",X"20",X"10",X"40",X"10",X"80",
		X"09",X"04",X"06",X"0A",X"00",X"12",X"00",X"22",X"00",X"42",X"00",X"42",X"00",X"24",X"00",X"18",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"0F",X"07",X"C0",X"08",X"20",X"10",X"20",X"10",X"40",
		X"08",X"84",X"07",X"0A",X"00",X"12",X"00",X"22",X"00",X"42",X"00",X"82",X"00",X"44",X"00",X"28",
		X"00",X"10",X"00",X"00",X"00",X"00",X"02",X"0F",X"07",X"C0",X"08",X"20",X"08",X"10",X"08",X"20",
		X"04",X"C0",X"05",X"06",X"02",X"1A",X"00",X"22",X"00",X"42",X"00",X"82",X"00",X"44",X"00",X"28",
		X"00",X"10",X"00",X"00",X"00",X"00",X"02",X"0F",X"07",X"C0",X"08",X"20",X"08",X"10",X"04",X"20",
		X"04",X"C0",X"03",X"06",X"02",X"0A",X"00",X"32",X"00",X"42",X"00",X"82",X"00",X"84",X"00",X"48",
		X"00",X"30",X"00",X"00",X"00",X"00",X"02",X"0F",X"07",X"C0",X"08",X"20",X"04",X"10",X"04",X"18",
		X"02",X"E0",X"03",X"00",X"00",X"06",X"00",X"1A",X"00",X"72",X"00",X"82",X"00",X"84",X"00",X"48",
		X"00",X"50",X"00",X"60",X"00",X"00",X"02",X"0F",X"07",X"C0",X"04",X"20",X"02",X"10",X"02",X"18",
		X"02",X"60",X"03",X"80",X"00",X"00",X"00",X"0E",X"00",X"32",X"00",X"C2",X"00",X"84",X"00",X"88",
		X"00",X"90",X"00",X"60",X"00",X"40",X"02",X"0F",X"03",X"C0",X"02",X"20",X"02",X"10",X"02",X"08",
		X"02",X"3C",X"01",X"C0",X"00",X"00",X"00",X"00",X"00",X"3E",X"00",X"C2",X"00",X"84",X"00",X"88",
		X"00",X"90",X"00",X"A0",X"00",X"C0",X"02",X"0F",X"03",X"C0",X"02",X"20",X"01",X"10",X"01",X"08",
		X"01",X"3C",X"01",X"C0",X"00",X"00",X"00",X"00",X"00",X"1E",X"01",X"E2",X"01",X"04",X"01",X"08",
		X"01",X"10",X"00",X"A0",X"00",X"C0",X"02",X"0F",X"01",X"C0",X"01",X"20",X"01",X"10",X"01",X"08",
		X"01",X"04",X"01",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"FE",X"01",X"04",X"01",X"08",
		X"01",X"10",X"01",X"20",X"01",X"C0",X"02",X"0F",X"00",X"C0",X"00",X"A0",X"01",X"10",X"01",X"08",
		X"01",X"04",X"01",X"E2",X"00",X"1E",X"00",X"00",X"00",X"00",X"01",X"E0",X"01",X"1C",X"02",X"08",
		X"02",X"10",X"02",X"20",X"03",X"C0",X"02",X"0F",X"00",X"C0",X"00",X"A0",X"00",X"90",X"00",X"88",
		X"00",X"84",X"00",X"C2",X"00",X"3E",X"00",X"00",X"00",X"00",X"01",X"C0",X"02",X"3C",X"02",X"08",
		X"02",X"10",X"02",X"20",X"03",X"C0",X"02",X"0F",X"00",X"40",X"00",X"A0",X"00",X"90",X"00",X"88",
		X"00",X"84",X"00",X"C2",X"00",X"72",X"00",X"0E",X"00",X"00",X"03",X"80",X"02",X"70",X"02",X"08",
		X"02",X"10",X"04",X"20",X"07",X"C0",X"02",X"0F",X"00",X"00",X"00",X"30",X"00",X"48",X"00",X"44",
		X"00",X"82",X"00",X"82",X"00",X"62",X"00",X"1A",X"00",X"06",X"01",X"00",X"02",X"E0",X"04",X"18",
		X"04",X"10",X"08",X"20",X"07",X"C0",X"02",X"0F",X"00",X"00",X"00",X"20",X"00",X"50",X"00",X"48",
		X"00",X"84",X"00",X"82",X"00",X"62",X"00",X"12",X"00",X"0A",X"03",X"06",X"04",X"C0",X"04",X"20",
		X"08",X"10",X"08",X"20",X"07",X"C0",X"02",X"0F",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"28",
		X"00",X"44",X"00",X"82",X"00",X"62",X"00",X"12",X"00",X"0A",X"03",X"06",X"04",X"80",X"08",X"60",
		X"08",X"10",X"08",X"20",X"07",X"C0",X"02",X"0F",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"28",
		X"00",X"44",X"00",X"82",X"00",X"42",X"00",X"22",X"00",X"12",X"07",X"0E",X"09",X"80",X"08",X"40",
		X"10",X"20",X"10",X"20",X"0F",X"C0",X"02",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",
		X"00",X"34",X"00",X"42",X"00",X"42",X"00",X"22",X"00",X"12",X"06",X"0A",X"09",X"04",X"10",X"80",
		X"10",X"40",X"08",X"20",X"07",X"C0",X"02",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",
		X"00",X"34",X"00",X"42",X"00",X"82",X"00",X"42",X"04",X"22",X"0A",X"12",X"11",X"0C",X"20",X"80",
		X"10",X"40",X"08",X"20",X"07",X"C0",X"02",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",
		X"00",X"14",X"00",X"22",X"00",X"42",X"00",X"42",X"04",X"22",X"0A",X"12",X"31",X"14",X"20",X"88",
		X"10",X"80",X"08",X"40",X"07",X"C0",X"02",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0C",X"00",X"12",X"00",X"62",X"00",X"42",X"0C",X"22",X"32",X"22",X"42",X"14",X"21",X"08",
		X"10",X"80",X"08",X"40",X"07",X"C0",X"02",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"00",X"1A",X"00",X"62",X"00",X"42",X"1C",X"22",X"62",X"22",X"42",X"24",X"21",X"18",
		X"11",X"10",X"09",X"00",X"07",X"00",X"02",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0E",X"00",X"32",X"00",X"42",X"3C",X"42",X"42",X"22",X"42",X"24",X"22",X"28",
		X"11",X"10",X"09",X"00",X"07",X"00",X"02",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"3E",X"00",X"42",X"FC",X"42",X"84",X"42",X"42",X"24",X"22",X"28",
		X"12",X"30",X"0A",X"20",X"06",X"00",X"02",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"06",X"3C",X"7A",X"C4",X"42",X"84",X"42",X"44",X"44",X"24",X"48",
		X"14",X"50",X"0C",X"60",X"04",X"00",X"02",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"7E",X"84",X"42",X"84",X"42",X"44",X"44",X"24",X"48",
		X"14",X"50",X"0C",X"60",X"04",X"40",X"02",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"00",X"BC",X"7E",X"84",X"42",X"84",X"42",X"44",X"44",X"24",X"48",
		X"14",X"90",X"08",X"A0",X"00",X"C0",X"02",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"F8",X"00",X"84",X"00",X"84",X"7E",X"84",X"42",X"48",X"84",X"28",X"88",
		X"18",X"90",X"08",X"A0",X"00",X"C0",X"02",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"40",X"00",X"B8",X"00",X"84",X"00",X"84",X"70",X"88",X"8C",X"48",X"84",X"28",X"88",
		X"11",X"10",X"01",X"20",X"01",X"C0",X"02",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"00",X"B0",X"00",X"8C",X"00",X"84",X"00",X"88",X"60",X"88",X"98",X"48",X"84",X"31",X"08",
		X"11",X"10",X"02",X"20",X"03",X"C0",X"02",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"60",X"00",X"90",X"00",X"88",X"00",X"84",X"00",X"88",X"60",X"88",X"90",X"50",X"88",X"21",X"08",
		X"02",X"10",X"02",X"20",X"03",X"C0",X"02",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"70",X"00",X"8C",X"00",X"84",X"00",X"84",X"00",X"88",X"40",X"90",X"B0",X"50",X"88",X"21",X"08",
		X"02",X"10",X"04",X"20",X"07",X"C0",X"02",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",
		X"58",X"00",X"84",X"00",X"84",X"00",X"84",X"00",X"88",X"00",X"90",X"E0",X"61",X"10",X"02",X"08",
		X"04",X"10",X"04",X"20",X"07",X"C0",X"02",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",
		X"48",X"00",X"84",X"00",X"84",X"00",X"88",X"00",X"90",X"00",X"A0",X"C0",X"41",X"20",X"02",X"10",
		X"04",X"10",X"08",X"20",X"07",X"C0",X"02",X"0F",X"00",X"00",X"00",X"00",X"10",X"00",X"28",X"00",
		X"48",X"00",X"84",X"00",X"84",X"00",X"88",X"00",X"90",X"00",X"E1",X"C0",X"02",X"20",X"04",X"10",
		X"08",X"10",X"08",X"20",X"07",X"C0",X"02",X"0F",X"00",X"00",X"00",X"00",X"10",X"00",X"28",X"00",
		X"44",X"00",X"84",X"00",X"88",X"00",X"90",X"00",X"A0",X"00",X"C1",X"80",X"02",X"40",X"0C",X"20",
		X"10",X"20",X"08",X"20",X"07",X"C0",X"02",X"0F",X"00",X"00",X"08",X"00",X"14",X"00",X"24",X"00",
		X"42",X"00",X"82",X"00",X"8C",X"00",X"90",X"00",X"A0",X"00",X"C1",X"80",X"06",X"40",X"08",X"40",
		X"10",X"20",X"08",X"20",X"07",X"C0",X"02",X"0F",X"00",X"00",X"08",X"00",X"14",X"00",X"24",X"00",
		X"42",X"00",X"82",X"00",X"8C",X"00",X"B0",X"00",X"C0",X"00",X"01",X"80",X"1E",X"40",X"20",X"40",
		X"10",X"40",X"08",X"20",X"07",X"C0",X"02",X"0F",X"00",X"00",X"0C",X"00",X"12",X"00",X"22",X"00",
		X"42",X"00",X"86",X"00",X"98",X"00",X"E0",X"00",X"00",X"00",X"03",X"00",X"1C",X"80",X"20",X"80",
		X"10",X"40",X"08",X"40",X"07",X"C0",X"02",X"0F",X"06",X"00",X"0A",X"00",X"12",X"00",X"22",X"00",
		X"42",X"00",X"86",X"00",X"F8",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"78",X"80",X"20",X"80",
		X"10",X"80",X"08",X"80",X"07",X"80",X"02",X"0F",X"06",X"00",X"0A",X"00",X"11",X"00",X"21",X"00",
		X"41",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"41",X"00",X"21",X"00",
		X"11",X"00",X"08",X"80",X"07",X"80",X"02",X"0F",X"07",X"00",X"09",X"00",X"11",X"00",X"21",X"00",
		X"41",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"41",X"00",X"21",X"00",
		X"11",X"00",X"09",X"00",X"07",X"00",X"02",X"0F",X"07",X"80",X"08",X"80",X"11",X"00",X"21",X"00",
		X"41",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"41",X"00",X"21",X"00",
		X"11",X"00",X"0A",X"00",X"06",X"00",X"02",X"0F",X"07",X"80",X"08",X"80",X"10",X"80",X"20",X"80",
		X"78",X"80",X"07",X"00",X"00",X"00",X"00",X"00",X"F8",X"00",X"86",X"00",X"42",X"00",X"22",X"00",
		X"12",X"00",X"0A",X"00",X"06",X"00",X"02",X"0F",X"07",X"80",X"08",X"80",X"10",X"80",X"20",X"80",
		X"1C",X"80",X"03",X"80",X"00",X"00",X"E0",X"00",X"98",X"00",X"84",X"00",X"42",X"00",X"22",X"00",
		X"12",X"00",X"0A",X"00",X"04",X"00",X"02",X"0F",X"07",X"C0",X"08",X"20",X"10",X"40",X"38",X"40",
		X"06",X"80",X"01",X"00",X"C0",X"00",X"B0",X"00",X"8C",X"00",X"82",X"00",X"42",X"00",X"24",X"00",
		X"14",X"00",X"0C",X"00",X"00",X"00",X"02",X"0F",X"07",X"C0",X"08",X"20",X"10",X"20",X"08",X"40",
		X"06",X"80",X"C1",X"00",X"A0",X"00",X"90",X"00",X"8C",X"00",X"82",X"00",X"42",X"00",X"24",X"00",
		X"18",X"00",X"00",X"00",X"00",X"00",X"02",X"0F",X"07",X"C0",X"08",X"20",X"10",X"20",X"0C",X"20",
		X"02",X"40",X"C1",X"C0",X"A0",X"00",X"90",X"00",X"8C",X"00",X"82",X"00",X"42",X"00",X"2C",X"00",
		X"10",X"00",X"00",X"00",X"00",X"00",X"02",X"0F",X"07",X"C0",X"08",X"20",X"08",X"10",X"04",X"20",
		X"02",X"20",X"E1",X"C0",X"90",X"00",X"88",X"00",X"84",X"00",X"82",X"00",X"44",X"00",X"28",X"00",
		X"10",X"00",X"00",X"00",X"00",X"00",X"02",X"0F",X"07",X"C0",X"08",X"20",X"04",X"10",X"02",X"10",
		X"41",X"20",X"A0",X"C0",X"90",X"00",X"88",X"00",X"84",X"00",X"84",X"00",X"48",X"00",X"30",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"0F",X"07",X"C0",X"08",X"20",X"04",X"10",X"02",X"08",
		X"61",X"30",X"90",X"C0",X"88",X"00",X"84",X"00",X"82",X"00",X"84",X"00",X"58",X"00",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"0F",X"07",X"C0",X"04",X"20",X"02",X"10",X"21",X"08",
		X"51",X"10",X"90",X"A0",X"88",X"40",X"84",X"00",X"84",X"00",X"88",X"00",X"70",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"0F",X"03",X"C0",X"02",X"20",X"02",X"10",X"21",X"08",
		X"51",X"08",X"88",X"90",X"88",X"60",X"84",X"00",X"84",X"00",X"98",X"00",X"60",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"0F",X"01",X"C0",X"01",X"20",X"01",X"10",X"31",X"08",
		X"48",X"84",X"88",X"9C",X"88",X"60",X"84",X"00",X"88",X"00",X"B0",X"00",X"40",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"0F",X"01",X"C0",X"01",X"20",X"11",X"10",X"28",X"88",
		X"48",X"84",X"88",X"84",X"84",X"78",X"84",X"00",X"B8",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"0F",X"00",X"C0",X"08",X"A0",X"18",X"90",X"28",X"88",
		X"48",X"84",X"84",X"42",X"84",X"7E",X"84",X"00",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"0F",X"00",X"40",X"0C",X"60",X"14",X"50",X"24",X"48",
		X"44",X"44",X"84",X"42",X"84",X"46",X"BC",X"78",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FA",X"10",X"FA",X"10",X"FA",X"10",X"18",X"11",X"18",X"11",
		X"18",X"11",X"36",X"11",X"36",X"11",X"36",X"11",X"18",X"11",X"18",X"11",X"18",X"11",X"FA",X"10",
		X"FA",X"10",X"FA",X"10",X"54",X"11",X"54",X"11",X"54",X"11",X"72",X"11",X"72",X"11",X"72",X"11",
		X"54",X"11",X"54",X"11",X"54",X"11",X"00",X"00",X"86",X"10",X"90",X"11",X"90",X"11",X"AE",X"11",
		X"AE",X"11",X"CE",X"11",X"CE",X"11",X"EC",X"11",X"EC",X"11",X"0A",X"12",X"0A",X"12",X"24",X"12",
		X"24",X"12",X"3E",X"12",X"3E",X"12",X"48",X"12",X"48",X"12",X"48",X"12",X"48",X"12",X"48",X"12",
		X"48",X"12",X"48",X"12",X"3E",X"12",X"3E",X"12",X"3E",X"12",X"3E",X"12",X"52",X"12",X"52",X"12",
		X"52",X"12",X"52",X"12",X"5E",X"12",X"00",X"00",X"BA",X"10",X"02",X"0E",X"40",X"20",X"20",X"40",
		X"10",X"80",X"3F",X"C0",X"46",X"C0",X"FF",X"40",X"C1",X"40",X"D9",X"40",X"D1",X"40",X"C1",X"40",
		X"FF",X"40",X"81",X"40",X"A5",X"80",X"FF",X"00",X"02",X"0E",X"42",X"00",X"22",X"00",X"12",X"00",
		X"3F",X"C0",X"46",X"C0",X"FF",X"40",X"C1",X"40",X"D9",X"40",X"D1",X"40",X"C1",X"40",X"FF",X"40",
		X"81",X"40",X"A5",X"80",X"FF",X"00",X"02",X"0E",X"28",X"00",X"14",X"00",X"0A",X"00",X"3F",X"C0",
		X"46",X"C0",X"FF",X"40",X"C1",X"40",X"D9",X"40",X"D1",X"40",X"C1",X"40",X"FF",X"40",X"81",X"40",
		X"A5",X"80",X"FF",X"00",X"02",X"0E",X"04",X"20",X"04",X"40",X"04",X"80",X"3F",X"C0",X"46",X"C0",
		X"FF",X"40",X"C1",X"40",X"D9",X"40",X"D1",X"40",X"C1",X"40",X"FF",X"40",X"81",X"40",X"A5",X"80",
		X"FF",X"00",X"02",X"0E",X"00",X"A0",X"01",X"40",X"02",X"80",X"3F",X"C0",X"46",X"C0",X"FF",X"40",
		X"C1",X"40",X"D9",X"40",X"D1",X"40",X"C1",X"40",X"FF",X"40",X"81",X"40",X"A5",X"80",X"FF",X"00",
		X"02",X"0E",X"00",X"00",X"20",X"40",X"10",X"80",X"2D",X"C0",X"46",X"C0",X"7F",X"00",X"C1",X"40",
		X"D9",X"40",X"C1",X"40",X"C1",X"00",X"EF",X"40",X"81",X"40",X"A1",X"80",X"7F",X"00",X"02",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"21",X"00",X"17",X"00",X"4C",X"C0",X"AB",X"00",X"C0",X"40",
		X"81",X"00",X"41",X"40",X"C0",X"00",X"AD",X"00",X"00",X"40",X"A4",X"80",X"E9",X"00",X"02",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"12",X"00",X"0C",X"00",X"2A",X"80",X"40",X"40",X"00",X"00",
		X"41",X"40",X"40",X"00",X"A4",X"00",X"00",X"40",X"A5",X"00",X"54",X"00",X"02",X"0E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"2A",X"00",X"44",X"40",X"10",X"00",X"41",X"00",
		X"50",X"00",X"24",X"00",X"12",X"40",X"00",X"00",X"04",X"00",X"02",X"0C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"28",X"00",X"44",X"80",X"10",X"00",X"45",X"00",X"10",X"00",
		X"00",X"00",X"04",X"00",X"02",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"28",X"00",X"44",X"80",X"10",X"00",X"45",X"00",X"10",X"00",X"00",X"00",X"04",X"00",X"01",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"30",X"01",X"08",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"10",X"01",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"3C",X"3C",X"18",X"01",X"01",
		X"00",X"01",X"0A",X"10",X"02",X"0E",X"10",X"10",X"10",X"08",X"0E",X"02",X"10",X"01",X"0A",X"10",
		X"00",X"2E",X"10",X"10",X"10",X"28",X"2E",X"00",X"10",X"01",X"0A",X"10",X"00",X"6C",X"10",X"10",
		X"10",X"28",X"6C",X"00",X"10",X"01",X"0A",X"10",X"00",X"E8",X"10",X"10",X"10",X"28",X"E8",X"00",
		X"10",X"01",X"0A",X"10",X"80",X"E0",X"10",X"10",X"10",X"20",X"E0",X"80",X"10",X"E9",X"12",X"E9",
		X"12",X"E9",X"12",X"F0",X"12",X"F0",X"12",X"F0",X"12",X"F8",X"12",X"F8",X"12",X"F8",X"12",X"01",
		X"13",X"01",X"13",X"01",X"13",X"0B",X"13",X"0B",X"13",X"0B",X"13",X"15",X"13",X"15",X"13",X"15",
		X"13",X"20",X"13",X"20",X"13",X"20",X"13",X"15",X"13",X"15",X"13",X"15",X"13",X"0B",X"13",X"0B",
		X"13",X"0B",X"13",X"01",X"13",X"01",X"13",X"01",X"13",X"F8",X"12",X"F8",X"12",X"F8",X"12",X"F0",
		X"12",X"F0",X"12",X"F0",X"12",X"00",X"00",X"9D",X"12",X"01",X"05",X"00",X"00",X"00",X"00",X"10",
		X"01",X"06",X"00",X"00",X"00",X"10",X"10",X"10",X"01",X"07",X"00",X"00",X"28",X"10",X"10",X"10",
		X"28",X"01",X"08",X"00",X"00",X"6C",X"10",X"10",X"10",X"28",X"44",X"01",X"08",X"00",X"82",X"EE",
		X"10",X"10",X"10",X"28",X"C6",X"01",X"09",X"00",X"82",X"EE",X"10",X"10",X"10",X"28",X"C6",X"82",
		X"01",X"0A",X"10",X"82",X"EE",X"10",X"10",X"10",X"28",X"C6",X"82",X"10",X"01",X"09",X"08",X"09",
		X"0A",X"14",X"6B",X"14",X"28",X"48",X"08",X"01",X"08",X"00",X"41",X"2A",X"14",X"6B",X"14",X"2A",
		X"41",X"01",X"09",X"08",X"48",X"28",X"14",X"6B",X"14",X"0A",X"09",X"08",X"01",X"09",X"08",X"49",
		X"2A",X"14",X"2A",X"14",X"2A",X"49",X"08",X"02",X"0A",X"01",X"00",X"10",X"10",X"0C",X"60",X"03",
		X"80",X"05",X"40",X"09",X"20",X"02",X"80",X"0E",X"E0",X"10",X"10",X"01",X"00",X"02",X"09",X"00",
		X"00",X"30",X"18",X"80",X"20",X"03",X"90",X"11",X"10",X"09",X"20",X"10",X"10",X"0E",X"E0",X"11",
		X"10",X"02",X"0A",X"00",X"00",X"08",X"08",X"13",X"84",X"01",X"00",X"01",X"00",X"20",X"42",X"10",
		X"04",X"20",X"02",X"08",X"08",X"30",X"06",X"02",X"0C",X"10",X"10",X"23",X"88",X"01",X"00",X"01",
		X"00",X"00",X"02",X"00",X"00",X"40",X"08",X"00",X"00",X"20",X"00",X"00",X"08",X"08",X"00",X"00",
		X"20",X"02",X"0D",X"02",X"00",X"80",X"01",X"10",X"00",X"00",X"00",X"00",X"02",X"40",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"08",X"00",X"00",X"00",X"80",X"01",X"01",X"00",
		X"04",X"14",X"04",X"14",X"0D",X"14",X"0D",X"14",X"15",X"14",X"15",X"14",X"1C",X"14",X"1C",X"14",
		X"23",X"14",X"23",X"14",X"2B",X"14",X"2B",X"14",X"2B",X"14",X"2B",X"14",X"23",X"14",X"23",X"14",
		X"1C",X"14",X"1C",X"14",X"15",X"14",X"15",X"14",X"0D",X"14",X"0D",X"14",X"04",X"14",X"04",X"14",
		X"00",X"00",X"D0",X"13",X"01",X"07",X"10",X"00",X"00",X"99",X"00",X"00",X"10",X"01",X"06",X"00",
		X"10",X"00",X"54",X"00",X"10",X"01",X"05",X"00",X"00",X"10",X"38",X"10",X"01",X"05",X"00",X"00",
		X"28",X"10",X"28",X"01",X"06",X"00",X"44",X"00",X"10",X"00",X"44",X"01",X"07",X"82",X"00",X"00",
		X"10",X"00",X"00",X"82",X"01",X"02",X"18",X"18",X"01",X"03",X"10",X"38",X"10",X"01",X"04",X"18",
		X"3C",X"3C",X"18",X"01",X"05",X"38",X"7C",X"7C",X"7C",X"38",X"01",X"06",X"3C",X"7E",X"7E",X"7E",
		X"7E",X"3C",X"01",X"07",X"38",X"7C",X"FE",X"FE",X"FE",X"7C",X"38",X"01",X"08",X"3C",X"7E",X"FF",
		X"FF",X"FF",X"FF",X"7E",X"3C",X"01",X"08",X"3C",X"7E",X"DB",X"FF",X"FF",X"BD",X"42",X"3C",X"8B",
		X"14",X"8B",X"14",X"8B",X"14",X"8B",X"14",X"9F",X"14",X"9F",X"14",X"9F",X"14",X"9F",X"14",X"B3",
		X"14",X"B3",X"14",X"B3",X"14",X"B3",X"14",X"00",X"00",X"6F",X"14",X"02",X"09",X"01",X"00",X"00",
		X"00",X"01",X"00",X"13",X"90",X"28",X"28",X"40",X"04",X"B6",X"DA",X"40",X"04",X"2B",X"68",X"02",
		X"09",X"00",X"00",X"00",X"00",X"01",X"00",X"13",X"90",X"28",X"28",X"40",X"04",X"9B",X"6A",X"40",
		X"04",X"26",X"C8",X"02",X"09",X"00",X"00",X"01",X"00",X"00",X"00",X"13",X"90",X"28",X"28",X"40",
		X"04",X"AD",X"B2",X"40",X"04",X"2D",X"A8",X"DB",X"14",X"DB",X"14",X"DB",X"14",X"DB",X"14",X"F7",
		X"14",X"F7",X"14",X"F7",X"14",X"F7",X"14",X"00",X"00",X"C7",X"14",X"02",X"0D",X"02",X"00",X"04",
		X"00",X"02",X"00",X"04",X"00",X"02",X"00",X"55",X"00",X"A8",X"A8",X"05",X"50",X"02",X"00",X"01",
		X"00",X"02",X"00",X"01",X"00",X"02",X"00",X"02",X"0D",X"01",X"00",X"00",X"01",X"01",X"00",X"00",
		X"80",X"01",X"00",X"02",X"A8",X"55",X"54",X"2A",X"80",X"01",X"00",X"02",X"00",X"01",X"00",X"02",
		X"00",X"01",X"00",X"71",X"15",X"71",X"15",X"68",X"15",X"68",X"15",X"5E",X"15",X"5E",X"15",X"53",
		X"15",X"53",X"15",X"3B",X"15",X"3B",X"15",X"53",X"15",X"53",X"15",X"5E",X"15",X"5E",X"15",X"68",
		X"15",X"68",X"15",X"71",X"15",X"71",X"15",X"00",X"00",X"13",X"15",X"02",X"0B",X"1C",X"00",X"22",
		X"00",X"41",X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"41",X"00",X"22",
		X"00",X"1C",X"00",X"01",X"09",X"00",X"00",X"1C",X"22",X"41",X"41",X"41",X"22",X"1C",X"01",X"08",
		X"00",X"00",X"00",X"1C",X"22",X"22",X"22",X"1C",X"01",X"07",X"00",X"00",X"00",X"00",X"1C",X"14",
		X"1C",X"01",X"06",X"00",X"00",X"00",X"00",X"00",X"08",X"95",X"15",X"95",X"15",X"95",X"15",X"95",
		X"15",X"95",X"15",X"95",X"15",X"9F",X"15",X"9F",X"15",X"9F",X"15",X"9F",X"15",X"9F",X"15",X"9F",
		X"15",X"00",X"00",X"79",X"15",X"01",X"08",X"10",X"08",X"10",X"AA",X"55",X"08",X"10",X"08",X"01",
		X"08",X"08",X"10",X"08",X"55",X"AA",X"10",X"08",X"10",X"BD",X"15",X"BD",X"15",X"C2",X"15",X"C2",
		X"15",X"C7",X"15",X"C7",X"15",X"CC",X"15",X"CC",X"15",X"00",X"00",X"A9",X"15",X"01",X"03",X"22",
		X"57",X"8A",X"01",X"03",X"42",X"AF",X"12",X"01",X"03",X"8A",X"57",X"22",X"01",X"03",X"12",X"AF",
		X"42",X"05",X"16",X"05",X"16",X"10",X"16",X"10",X"16",X"1B",X"16",X"1B",X"16",X"26",X"16",X"26",
		X"16",X"31",X"16",X"31",X"16",X"3C",X"16",X"3C",X"16",X"46",X"16",X"46",X"16",X"4F",X"16",X"4F",
		X"16",X"59",X"16",X"59",X"16",X"64",X"16",X"64",X"16",X"6F",X"16",X"6F",X"16",X"7A",X"16",X"7A",
		X"16",X"00",X"00",X"D1",X"15",X"01",X"09",X"FF",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"FF",
		X"01",X"09",X"7F",X"C1",X"81",X"81",X"81",X"81",X"81",X"83",X"FE",X"01",X"09",X"3F",X"21",X"E1",
		X"81",X"81",X"81",X"87",X"84",X"FC",X"01",X"09",X"1F",X"11",X"11",X"F1",X"81",X"8F",X"88",X"88",
		X"F8",X"01",X"09",X"0F",X"09",X"09",X"09",X"FF",X"90",X"90",X"90",X"F0",X"01",X"08",X"00",X"0F",
		X"09",X"F9",X"99",X"9F",X"90",X"F0",X"01",X"07",X"00",X"00",X"FF",X"99",X"99",X"99",X"FF",X"01",
		X"08",X"00",X"F0",X"90",X"9F",X"99",X"F9",X"09",X"0F",X"01",X"09",X"F0",X"90",X"90",X"90",X"FF",
		X"09",X"09",X"09",X"0F",X"01",X"09",X"E0",X"A0",X"A0",X"FC",X"24",X"3F",X"05",X"05",X"07",X"01",
		X"09",X"C0",X"C0",X"FE",X"42",X"42",X"42",X"7F",X"03",X"03",X"01",X"09",X"80",X"FF",X"81",X"81",
		X"81",X"81",X"81",X"FF",X"01",X"2D",X"FD",X"21",X"73",X"40",X"FD",X"36",X"19",X"04",X"CD",X"B0",
		X"28",X"CD",X"0B",X"28",X"D9",X"3A",X"EE",X"43",X"CB",X"3F",X"CB",X"3F",X"E6",X"3F",X"CB",X"27",
		X"5F",X"16",X"00",X"21",X"1E",X"18",X"19",X"19",X"19",X"46",X"23",X"4E",X"23",X"5E",X"23",X"56",
		X"D5",X"23",X"5E",X"23",X"56",X"DD",X"E5",X"DD",X"21",X"77",X"40",X"DD",X"7E",X"0B",X"80",X"6F",
		X"DD",X"7E",X"11",X"81",X"67",X"DD",X"E1",X"DD",X"72",X"0F",X"DD",X"73",X"0E",X"D1",X"DD",X"72",
		X"09",X"DD",X"73",X"08",X"DD",X"75",X"0B",X"DD",X"74",X"11",X"D9",X"DD",X"CB",X"14",X"DE",X"DD",
		X"36",X"15",X"FF",X"78",X"FE",X"00",X"20",X"05",X"21",X"DE",X"19",X"18",X"0F",X"21",X"B8",X"19",
		X"DD",X"36",X"15",X"0A",X"DD",X"CB",X"14",X"9E",X"DD",X"CB",X"14",X"D6",X"DD",X"75",X"12",X"DD",
		X"74",X"13",X"DD",X"CB",X"00",X"CE",X"DD",X"E5",X"E1",X"FD",X"E5",X"CD",X"D1",X"2B",X"FD",X"E1",
		X"DD",X"CB",X"00",X"D6",X"DD",X"E5",X"CD",X"F1",X"C6",X"CD",X"18",X"C7",X"CD",X"4B",X"28",X"DD",
		X"E1",X"DD",X"CB",X"00",X"7E",X"20",X"28",X"DD",X"CB",X"14",X"7E",X"C2",X"9D",X"17",X"DD",X"CB",
		X"14",X"6E",X"20",X"12",X"DD",X"35",X"15",X"20",X"0D",X"AF",X"DD",X"77",X"09",X"DD",X"77",X"08",
		X"DD",X"77",X"0F",X"DD",X"77",X"0E",X"DD",X"E5",X"3E",X"01",X"CD",X"40",X"28",X"18",X"D0",X"DD",
		X"E5",X"CD",X"34",X"3B",X"E1",X"11",X"0B",X"00",X"19",X"7E",X"D6",X"02",X"77",X"11",X"06",X"00",
		X"19",X"7E",X"D6",X"02",X"77",X"23",X"01",X"C8",X"19",X"71",X"23",X"70",X"DD",X"E5",X"CD",X"4B",
		X"28",X"DD",X"E1",X"DD",X"7E",X"00",X"B7",X"28",X"0E",X"21",X"66",X"1A",X"DD",X"7E",X"04",X"DD",
		X"46",X"05",X"BD",X"20",X"04",X"78",X"BC",X"28",X"14",X"DD",X"CB",X"14",X"5E",X"20",X"03",X"CD",
		X"AA",X"20",X"DD",X"E5",X"3E",X"01",X"CD",X"40",X"28",X"DD",X"E1",X"18",X"D6",X"3A",X"C1",X"43",
		X"FE",X"20",X"30",X"09",X"DD",X"E5",X"CD",X"4B",X"28",X"DD",X"E1",X"18",X"F0",X"CD",X"BD",X"28",
		X"DD",X"CB",X"14",X"5E",X"28",X"0A",X"21",X"F3",X"43",X"7E",X"35",X"CD",X"9E",X"C5",X"18",X"10",
		X"DD",X"CB",X"14",X"56",X"28",X"0A",X"21",X"ED",X"43",X"7E",X"CB",X"FF",X"35",X"CD",X"9E",X"C5",
		X"CD",X"4B",X"28",X"18",X"FB",X"06",X"0F",X"FD",X"21",X"A7",X"40",X"C5",X"FD",X"CB",X"00",X"56",
		X"C4",X"EC",X"17",X"01",X"30",X"00",X"FD",X"09",X"C1",X"10",X"F0",X"C9",X"FD",X"CB",X"14",X"46",
		X"C8",X"FD",X"66",X"13",X"FD",X"6E",X"12",X"5E",X"23",X"56",X"EB",X"56",X"23",X"5E",X"1C",X"DD",
		X"7E",X"11",X"FD",X"96",X"11",X"3C",X"F8",X"BB",X"D0",X"DD",X"7E",X"0B",X"FD",X"96",X"0B",X"F8",
		X"CB",X"22",X"CB",X"22",X"CB",X"22",X"14",X"BA",X"D0",X"FD",X"CB",X"00",X"F6",X"C9",X"06",X"FB",
		X"00",X"00",X"00",X"FC",X"07",X"FB",X"64",X"00",X"05",X"FC",X"07",X"FC",X"C7",X"00",X"14",X"FC",
		X"09",X"FC",X"29",X"01",X"2D",X"FC",X"0A",X"FC",X"87",X"01",X"4E",X"FC",X"0B",X"FD",X"E2",X"01",
		X"79",X"FC",X"0C",X"FD",X"38",X"02",X"AD",X"FC",X"0C",X"FD",X"89",X"02",X"E9",X"FC",X"0D",X"FE",
		X"D4",X"02",X"2C",X"FD",X"0E",X"FF",X"17",X"03",X"77",X"FD",X"0F",X"00",X"53",X"03",X"C7",X"FD",
		X"0F",X"01",X"87",X"03",X"1E",X"FE",X"0F",X"02",X"B2",X"03",X"78",X"FE",X"10",X"03",X"D3",X"03",
		X"D7",X"FE",X"10",X"04",X"EC",X"03",X"39",X"FF",X"10",X"05",X"FB",X"03",X"9C",X"FF",X"10",X"06",
		X"00",X"04",X"00",X"00",X"10",X"07",X"FB",X"03",X"64",X"00",X"10",X"08",X"EC",X"03",X"C7",X"00",
		X"10",X"09",X"D3",X"03",X"29",X"01",X"0F",X"0A",X"B2",X"03",X"87",X"01",X"0F",X"0B",X"87",X"03",
		X"E2",X"01",X"0F",X"0C",X"53",X"03",X"38",X"02",X"0E",X"0D",X"17",X"03",X"89",X"02",X"0D",X"0E",
		X"D4",X"02",X"D4",X"02",X"0D",X"0F",X"89",X"02",X"17",X"03",X"0C",X"0F",X"38",X"02",X"53",X"03",
		X"0B",X"0F",X"E2",X"01",X"87",X"03",X"0A",X"0F",X"87",X"01",X"B2",X"03",X"08",X"0F",X"29",X"01",
		X"D3",X"03",X"07",X"0F",X"C2",X"00",X"EC",X"03",X"07",X"0F",X"64",X"00",X"FB",X"03",X"06",X"0F",
		X"00",X"00",X"00",X"04",X"05",X"0F",X"9C",X"FF",X"FB",X"03",X"04",X"0F",X"39",X"FF",X"EC",X"03",
		X"03",X"0F",X"D7",X"FE",X"D3",X"03",X"02",X"0F",X"79",X"FE",X"B2",X"03",X"01",X"0F",X"1E",X"FE",
		X"87",X"03",X"00",X"0E",X"C8",X"FD",X"53",X"03",X"FF",X"0E",X"77",X"FD",X"17",X"03",X"FE",X"0E",
		X"2C",X"FD",X"D4",X"02",X"FE",X"0C",X"E9",X"FC",X"89",X"02",X"FE",X"0B",X"AD",X"FC",X"38",X"02",
		X"FE",X"0A",X"79",X"FC",X"E2",X"01",X"FD",X"0A",X"4E",X"FC",X"87",X"01",X"FD",X"09",X"2D",X"FC",
		X"29",X"01",X"FD",X"07",X"14",X"FC",X"C7",X"00",X"FC",X"07",X"05",X"FC",X"64",X"00",X"FC",X"06",
		X"00",X"FC",X"00",X"00",X"FC",X"05",X"05",X"FC",X"9C",X"FF",X"FC",X"03",X"14",X"FC",X"39",X"FF",
		X"FC",X"03",X"2D",X"FC",X"D7",X"FE",X"FC",X"01",X"4E",X"FC",X"79",X"FE",X"FD",X"00",X"79",X"FC",
		X"1E",X"FE",X"FD",X"00",X"AD",X"FC",X"C8",X"FD",X"FE",X"FF",X"E9",X"FC",X"77",X"FD",X"FE",X"FE",
		X"2C",X"FD",X"2C",X"FD",X"FE",X"FD",X"77",X"FD",X"E9",X"FC",X"FF",X"FC",X"C7",X"FD",X"AD",X"FC",
		X"00",X"FB",X"1E",X"FE",X"79",X"FC",X"02",X"FB",X"78",X"FE",X"4E",X"FC",X"04",X"FB",X"D7",X"FE",
		X"2D",X"FC",X"05",X"FB",X"39",X"FF",X"14",X"FC",X"05",X"FB",X"9C",X"FF",X"05",X"FC",X"09",X"1A",
		X"0F",X"1A",X"15",X"1A",X"1B",X"1A",X"21",X"1A",X"00",X"00",X"9E",X"19",X"F5",X"19",X"FA",X"19",
		X"FF",X"19",X"04",X"1A",X"00",X"00",X"AC",X"19",X"F2",X"19",X"F2",X"19",X"69",X"1A",X"70",X"1A",
		X"77",X"1A",X"7E",X"1A",X"00",X"00",X"BC",X"19",X"27",X"1A",X"32",X"1A",X"3B",X"1A",X"45",X"1A",
		X"51",X"1A",X"45",X"1A",X"51",X"1A",X"5B",X"1A",X"66",X"1A",X"00",X"00",X"D8",X"19",X"F2",X"19",
		X"F2",X"19",X"F2",X"19",X"F2",X"19",X"EC",X"19",X"00",X"00",X"E6",X"19",X"01",X"04",X"40",X"E0",
		X"E0",X"40",X"01",X"01",X"40",X"01",X"03",X"40",X"80",X"40",X"01",X"03",X"A0",X"40",X"40",X"01",
		X"03",X"40",X"20",X"40",X"01",X"03",X"40",X"40",X"A0",X"01",X"04",X"80",X"40",X"40",X"20",X"01",
		X"04",X"00",X"C0",X"60",X"00",X"01",X"04",X"00",X"60",X"C0",X"00",X"01",X"04",X"20",X"40",X"40",
		X"80",X"01",X"04",X"40",X"40",X"40",X"40",X"01",X"09",X"10",X"6C",X"54",X"AA",X"54",X"AA",X"54",
		X"6C",X"10",X"01",X"07",X"00",X"00",X"08",X"28",X"1C",X"10",X"08",X"01",X"08",X"00",X"28",X"40",
		X"10",X"04",X"48",X"00",X"10",X"01",X"0A",X"08",X"54",X"18",X"6A",X"96",X"60",X"16",X"58",X"20",
		X"10",X"01",X"08",X"08",X"40",X"10",X"02",X"80",X"20",X"02",X"48",X"01",X"09",X"00",X"10",X"01",
		X"40",X"00",X"00",X"00",X"81",X"08",X"01",X"01",X"00",X"01",X"05",X"90",X"00",X"00",X"00",X"90",
		X"01",X"05",X"40",X"10",X"00",X"80",X"20",X"01",X"05",X"60",X"00",X"90",X"00",X"60",X"01",X"05",
		X"20",X"80",X"00",X"10",X"40",X"F3",X"31",X"40",X"40",X"DB",X"60",X"CB",X"4F",X"C2",X"3A",X"07",
		X"21",X"86",X"F8",X"06",X"34",X"36",X"00",X"23",X"10",X"FB",X"21",X"00",X"40",X"01",X"00",X"04",
		X"AF",X"77",X"23",X"0D",X"20",X"FB",X"10",X"F9",X"CD",X"0B",X"1B",X"21",X"F2",X"F8",X"11",X"73",
		X"43",X"06",X"1E",X"7E",X"23",X"E6",X"F0",X"4F",X"7E",X"23",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",
		X"B1",X"12",X"13",X"10",X"EE",X"DB",X"49",X"2F",X"21",X"B5",X"F8",X"77",X"23",X"77",X"CD",X"E9",
		X"1A",X"CD",X"BF",X"1D",X"CD",X"92",X"1C",X"CD",X"B5",X"1E",X"CD",X"92",X"1C",X"CD",X"B0",X"2D",
		X"CA",X"CE",X"1A",X"CD",X"E9",X"1A",X"CD",X"BA",X"1C",X"F3",X"E1",X"22",X"D1",X"43",X"32",X"D3",
		X"43",X"31",X"40",X"40",X"CD",X"6A",X"29",X"DD",X"21",X"43",X"40",X"CD",X"B0",X"28",X"CD",X"0B",
		X"28",X"CD",X"7B",X"2B",X"2A",X"D1",X"43",X"3A",X"D3",X"43",X"E9",X"ED",X"73",X"5E",X"F8",X"31",
		X"5E",X"F8",X"F5",X"C5",X"D5",X"E5",X"DD",X"E5",X"DB",X"65",X"CB",X"7F",X"C2",X"31",X"05",X"3A",
		X"E1",X"43",X"B7",X"CC",X"AB",X"23",X"CD",X"60",X"1B",X"3A",X"E1",X"43",X"B7",X"20",X"1D",X"2A",
		X"AE",X"F8",X"7C",X"B5",X"28",X"19",X"DB",X"44",X"E6",X"C0",X"FE",X"40",X"20",X"11",X"7E",X"CB",
		X"7F",X"20",X"09",X"23",X"D3",X"44",X"CB",X"77",X"28",X"05",X"18",X"E6",X"21",X"00",X"00",X"22",
		X"AE",X"F8",X"DD",X"E1",X"E1",X"D1",X"C1",X"F1",X"ED",X"7B",X"5E",X"F8",X"D3",X"4C",X"ED",X"45",
		X"21",X"8E",X"F8",X"46",X"23",X"56",X"23",X"5E",X"23",X"0E",X"41",X"CB",X"80",X"CB",X"C2",X"ED",
		X"51",X"0D",X"ED",X"41",X"0C",X"CB",X"82",X"ED",X"51",X"0D",X"ED",X"59",X"0C",X"0C",X"06",X"03",
		X"79",X"0C",X"51",X"5E",X"23",X"4F",X"7E",X"23",X"ED",X"79",X"79",X"4A",X"ED",X"59",X"14",X"14",
		X"10",X"F1",X"0D",X"3E",X"00",X"06",X"04",X"B6",X"23",X"ED",X"79",X"E6",X"C0",X"C6",X"40",X"10",
		X"F6",X"C9",X"06",X"06",X"21",X"D4",X"F8",X"CD",X"A1",X"32",X"3A",X"E9",X"43",X"FE",X"02",X"CC",
		X"A1",X"32",X"CD",X"57",X"1C",X"01",X"0D",X"00",X"11",X"B5",X"43",X"21",X"85",X"1C",X"ED",X"B0",
		X"CD",X"7C",X"2E",X"2A",X"CF",X"43",X"AF",X"32",X"E1",X"43",X"3C",X"32",X"B1",X"F8",X"CD",X"51",
		X"3A",X"21",X"B5",X"43",X"11",X"C2",X"43",X"01",X"0D",X"00",X"ED",X"B0",X"3E",X"02",X"77",X"3A",
		X"E9",X"43",X"FE",X"02",X"28",X"04",X"AF",X"32",X"C3",X"43",X"CD",X"63",X"36",X"FB",X"AF",X"32",
		X"E4",X"43",X"32",X"F0",X"43",X"32",X"F3",X"43",X"32",X"ED",X"43",X"32",X"5E",X"F9",X"32",X"FD",
		X"43",X"3E",X"40",X"32",X"C0",X"43",X"32",X"C1",X"43",X"CD",X"CA",X"28",X"DD",X"CB",X"00",X"7E",
		X"28",X"0A",X"CD",X"57",X"C8",X"21",X"BF",X"43",X"36",X"10",X"18",X"D1",X"3E",X"3C",X"CD",X"40",
		X"28",X"CD",X"6A",X"29",X"21",X"B6",X"43",X"7E",X"C6",X"99",X"27",X"77",X"08",X"3A",X"BF",X"43",
		X"B7",X"CC",X"57",X"C8",X"08",X"E5",X"21",X"BF",X"43",X"36",X"10",X"E1",X"08",X"CD",X"70",X"1C",
		X"7E",X"B7",X"C2",X"EA",X"1B",X"08",X"20",X"F5",X"CD",X"70",X"1C",X"CD",X"3F",X"31",X"CD",X"70",
		X"1C",X"CD",X"3F",X"31",X"C3",X"CE",X"1A",X"21",X"00",X"00",X"22",X"AF",X"43",X"22",X"B1",X"43",
		X"22",X"B3",X"43",X"22",X"B7",X"F8",X"22",X"B8",X"F8",X"21",X"98",X"C0",X"22",X"AE",X"F8",X"C9",
		X"E5",X"21",X"B5",X"43",X"11",X"C2",X"43",X"06",X"0D",X"1A",X"4E",X"EB",X"12",X"71",X"EB",X"23",
		X"13",X"10",X"F6",X"E1",X"C9",X"01",X"03",X"00",X"FF",X"00",X"15",X"00",X"00",X"00",X"01",X"10",
		X"40",X"40",X"06",X"05",X"2A",X"88",X"F8",X"23",X"36",X"28",X"2B",X"CB",X"CE",X"DB",X"65",X"CB",
		X"47",X"28",X"04",X"3E",X"01",X"18",X"22",X"CD",X"83",X"1D",X"CD",X"9F",X"1D",X"C2",X"E3",X"1A",
		X"2A",X"88",X"F8",X"CB",X"4E",X"20",X"E6",X"10",X"DB",X"C9",X"6F",X"CD",X"F9",X"1C",X"CB",X"4D",
		X"3E",X"01",X"28",X"05",X"CD",X"F9",X"1C",X"3E",X"02",X"32",X"E9",X"43",X"2A",X"88",X"F8",X"CB",
		X"C6",X"E1",X"C3",X"A2",X"1B",X"E5",X"21",X"00",X"00",X"39",X"CD",X"E8",X"1C",X"77",X"06",X"02",
		X"11",X"78",X"D5",X"CD",X"A0",X"2F",X"E1",X"C9",X"3A",X"BB",X"F8",X"0F",X"0F",X"0F",X"0F",X"E6",
		X"0F",X"4F",X"3A",X"BA",X"F8",X"E6",X"F0",X"B1",X"C9",X"CD",X"E8",X"1C",X"C6",X"99",X"27",X"4F",
		X"E6",X"F0",X"32",X"BA",X"F8",X"79",X"07",X"07",X"07",X"07",X"E6",X"F0",X"32",X"BB",X"F8",X"C9",
		X"7E",X"B7",X"C8",X"C5",X"E5",X"35",X"78",X"3D",X"87",X"87",X"87",X"5F",X"16",X"00",X"21",X"BC",
		X"F8",X"19",X"06",X"08",X"CD",X"A1",X"32",X"E1",X"E5",X"11",X"05",X"00",X"19",X"7E",X"57",X"3C",
		X"E6",X"03",X"77",X"ED",X"78",X"E6",X"0F",X"CB",X"1A",X"17",X"4F",X"06",X"00",X"21",X"63",X"1D",
		X"09",X"7E",X"CB",X"42",X"28",X"04",X"07",X"07",X"07",X"07",X"E6",X"0F",X"C6",X"00",X"27",X"57",
		X"CD",X"E8",X"1C",X"FE",X"99",X"28",X"09",X"82",X"27",X"30",X"02",X"3E",X"99",X"CD",X"FF",X"1C",
		X"E1",X"C1",X"C9",X"11",X"11",X"22",X"22",X"33",X"33",X"44",X"44",X"55",X"55",X"66",X"66",X"77",
		X"77",X"AA",X"AA",X"EE",X"EE",X"00",X"11",X"11",X"22",X"00",X"55",X"00",X"77",X"00",X"21",X"11",
		X"21",X"11",X"32",X"C5",X"21",X"B2",X"F8",X"CD",X"E8",X"1C",X"F5",X"01",X"62",X"03",X"CD",X"10",
		X"1D",X"23",X"0C",X"10",X"F9",X"CD",X"E8",X"1C",X"C1",X"B8",X"C4",X"D5",X"1C",X"C1",X"C9",X"CD",
		X"E8",X"1C",X"2E",X"00",X"B7",X"28",X"08",X"FE",X"01",X"2E",X"01",X"28",X"02",X"2E",X"03",X"DB",
		X"49",X"2F",X"A5",X"C9",X"2A",X"AE",X"F8",X"7C",X"B5",X"C0",X"EB",X"22",X"AE",X"F8",X"C9",X"CD",
		X"65",X"1E",X"AF",X"32",X"EC",X"43",X"CD",X"47",X"CB",X"CD",X"40",X"2F",X"90",X"0C",X"BE",X"1F",
		X"31",X"39",X"38",X"31",X"20",X"53",X"54",X"45",X"52",X"4E",X"20",X"45",X"6C",X"65",X"63",X"74",
		X"72",X"6F",X"6E",X"69",X"63",X"73",X"2C",X"20",X"49",X"6E",X"63",X"2E",X"00",X"CD",X"D5",X"1C",
		X"CD",X"95",X"2E",X"CD",X"05",X"1F",X"1C",X"1F",X"58",X"1F",X"38",X"1F",X"77",X"1F",X"21",X"73",
		X"43",X"3E",X"01",X"32",X"40",X"40",X"11",X"38",X"18",X"D5",X"E5",X"7E",X"23",X"B6",X"23",X"B6",
		X"E1",X"E5",X"20",X"04",X"E1",X"D1",X"18",X"35",X"21",X"40",X"40",X"06",X"02",X"CD",X"A0",X"2F",
		X"13",X"E1",X"06",X"06",X"CD",X"AA",X"2F",X"13",X"AF",X"4E",X"CD",X"EE",X"2F",X"13",X"23",X"4E",
		X"CD",X"EE",X"2F",X"13",X"23",X"4E",X"CD",X"EE",X"2F",X"23",X"D1",X"7A",X"C6",X"10",X"57",X"3A",
		X"40",X"40",X"C6",X"01",X"27",X"32",X"40",X"40",X"FE",X"11",X"C2",X"09",X"1E",X"21",X"00",X"46",
		X"CD",X"5C",X"1E",X"21",X"00",X"5B",X"CD",X"5C",X"1E",X"21",X"80",X"5D",X"3E",X"FF",X"06",X"40",
		X"77",X"23",X"10",X"FC",X"C9",X"21",X"00",X"81",X"01",X"00",X"07",X"AF",X"77",X"23",X"0D",X"20",
		X"FB",X"10",X"F9",X"F3",X"ED",X"73",X"40",X"40",X"31",X"00",X"60",X"06",X"E0",X"11",X"00",X"00",
		X"D5",X"D5",X"D5",X"D5",X"D5",X"D5",X"D5",X"D5",X"D5",X"D5",X"D5",X"D5",X"D5",X"D5",X"D5",X"D5",
		X"10",X"EE",X"ED",X"7B",X"40",X"40",X"FB",X"DB",X"49",X"CB",X"57",X"20",X"13",X"DB",X"63",X"CB",
		X"7F",X"28",X"0D",X"3A",X"B5",X"43",X"FE",X"02",X"20",X"06",X"3E",X"FF",X"32",X"EC",X"43",X"C9",
		X"AF",X"32",X"EC",X"43",X"C9",X"CD",X"F5",X"1E",X"CD",X"E8",X"1C",X"28",X"21",X"3D",X"28",X"0F",
		X"CD",X"B4",X"CB",X"CD",X"05",X"1F",X"CF",X"1F",X"1C",X"20",X"F6",X"1F",X"39",X"20",X"C9",X"CD",
		X"AB",X"CB",X"CD",X"05",X"1F",X"8F",X"1F",X"1C",X"20",X"B1",X"1F",X"39",X"20",X"C9",X"CD",X"A2",
		X"CB",X"CD",X"05",X"1F",X"4D",X"20",X"7C",X"20",X"60",X"20",X"93",X"20",X"D9",X"11",X"9A",X"C0",
		X"CD",X"B4",X"1D",X"D9",X"C9",X"21",X"C0",X"5B",X"01",X"C0",X"02",X"AF",X"77",X"23",X"0D",X"C2",
		X"FC",X"1E",X"10",X"F8",X"C9",X"E1",X"54",X"5D",X"01",X"08",X"00",X"09",X"E5",X"EB",X"DB",X"60",
		X"E6",X"C0",X"07",X"07",X"07",X"4F",X"09",X"7E",X"23",X"66",X"6F",X"E9",X"CD",X"40",X"2F",X"90",
		X"28",X"00",X"4D",X"4F",X"4F",X"4E",X"20",X"57",X"41",X"52",X"20",X"48",X"69",X"67",X"68",X"20",
		X"53",X"63",X"6F",X"72",X"65",X"73",X"00",X"C9",X"CD",X"40",X"2F",X"90",X"20",X"00",X"53",X"63",
		X"6F",X"72",X"65",X"20",X"65",X"6C",X"65",X"76",X"65",X"73",X"20",X"64",X"75",X"20",X"4D",X"4F",
		X"4F",X"4E",X"20",X"57",X"41",X"52",X"00",X"C9",X"CD",X"40",X"2F",X"90",X"28",X"00",X"48",X"24",
		X"68",X"65",X"20",X"4D",X"4F",X"4F",X"4E",X"20",X"57",X"41",X"52",X"20",X"70",X"75",X"6E",X"6B",
		X"74",X"7A",X"61",X"68",X"6C",X"00",X"C9",X"CD",X"40",X"2F",X"90",X"38",X"00",X"4D",X"4F",X"4F",
		X"4E",X"20",X"57",X"41",X"52",X"20",X"52",X"65",X"63",X"6F",X"72",X"64",X"73",X"00",X"C9",X"CD",
		X"40",X"2F",X"90",X"14",X"BE",X"50",X"75",X"73",X"68",X"20",X"31",X"20",X"50",X"6C",X"61",X"79",
		X"65",X"72",X"20",X"53",X"74",X"61",X"72",X"74",X"20",X"42",X"75",X"74",X"74",X"6F",X"6E",X"00",
		X"C9",X"CD",X"40",X"2F",X"90",X"24",X"BE",X"50",X"6F",X"75",X"73",X"73",X"65",X"72",X"20",X"62",
		X"6F",X"75",X"74",X"6F",X"6E",X"20",X"73",X"74",X"61",X"72",X"74",X"20",X"31",X"00",X"C9",X"CD",
		X"40",X"2F",X"90",X"04",X"BE",X"50",X"75",X"73",X"68",X"20",X"31",X"20",X"6F",X"72",X"20",X"32",
		X"20",X"50",X"6C",X"61",X"79",X"65",X"72",X"20",X"53",X"74",X"61",X"72",X"74",X"20",X"42",X"75",
		X"74",X"74",X"6F",X"6E",X"00",X"C9",X"CD",X"40",X"2F",X"90",X"04",X"BE",X"50",X"72",X"65",X"73",
		X"73",X"65",X"72",X"20",X"6C",X"65",X"20",X"62",X"6F",X"75",X"74",X"6F",X"6E",X"20",X"73",X"74",
		X"61",X"72",X"74",X"20",X"31",X"20",X"6F",X"75",X"20",X"32",X"00",X"C9",X"CD",X"40",X"2F",X"90",
		X"38",X"BE",X"53",X"74",X"61",X"72",X"74",X"6B",X"6E",X"6F",X"65",X"70",X"66",X"65",X"20",X"64",
		X"72",X"25",X"65",X"63",X"6B",X"65",X"6E",X"00",X"C9",X"CD",X"40",X"2F",X"90",X"44",X"BE",X"50",
		X"75",X"6C",X"73",X"61",X"72",X"20",X"53",X"74",X"61",X"72",X"74",X"00",X"C9",X"CD",X"40",X"2F",
		X"90",X"58",X"BE",X"49",X"6E",X"73",X"65",X"72",X"74",X"20",X"43",X"6F",X"69",X"6E",X"00",X"C9",
		X"CD",X"40",X"2F",X"90",X"30",X"BE",X"49",X"6E",X"74",X"72",X"6F",X"64",X"75",X"69",X"72",X"65",
		X"20",X"75",X"6E",X"65",X"20",X"70",X"69",X"65",X"63",X"65",X"00",X"C9",X"CD",X"40",X"2F",X"90",
		X"48",X"BE",X"4D",X"25",X"6E",X"7A",X"65",X"20",X"65",X"69",X"6E",X"77",X"65",X"72",X"66",X"65",
		X"6E",X"00",X"C9",X"CD",X"40",X"2F",X"90",X"48",X"BE",X"50",X"6F",X"6E",X"67",X"61",X"20",X"6C",
		X"61",X"20",X"6D",X"6F",X"6E",X"65",X"64",X"61",X"00",X"C9",X"FD",X"21",X"77",X"40",X"FD",X"7E",
		X"0B",X"C6",X"04",X"DD",X"96",X"0B",X"D2",X"BB",X"20",X"ED",X"44",X"47",X"FD",X"7E",X"11",X"C6",
		X"04",X"DD",X"96",X"11",X"D2",X"C9",X"20",X"ED",X"44",X"4F",X"16",X"00",X"3E",X"0F",X"B9",X"38",
		X"03",X"B8",X"30",X"07",X"CB",X"38",X"CB",X"39",X"14",X"18",X"F3",X"79",X"07",X"07",X"07",X"07",
		X"B0",X"CB",X"22",X"D5",X"5F",X"16",X"00",X"21",X"99",X"21",X"19",X"19",X"7E",X"23",X"66",X"6F",
		X"E5",X"7B",X"0F",X"0F",X"0F",X"0F",X"5F",X"D5",X"D1",X"21",X"99",X"21",X"19",X"19",X"5E",X"23",
		X"56",X"E1",X"3A",X"B8",X"43",X"B7",X"28",X"18",X"F2",X"15",X"21",X"CB",X"2A",X"CB",X"1B",X"CB",
		X"2C",X"CB",X"1D",X"18",X"0B",X"47",X"CB",X"25",X"CB",X"14",X"CB",X"23",X"CB",X"12",X"10",X"F6",
		X"F1",X"F5",X"B7",X"28",X"0B",X"47",X"CB",X"2A",X"CB",X"1B",X"CB",X"2C",X"CB",X"1D",X"10",X"F6",
		X"FD",X"7E",X"0B",X"C6",X"04",X"DD",X"BE",X"0B",X"DC",X"8F",X"21",X"FD",X"7E",X"11",X"C6",X"04",
		X"DD",X"BE",X"11",X"EB",X"DC",X"8F",X"21",X"EB",X"F1",X"F5",X"B7",X"20",X"22",X"E5",X"F5",X"CD",
		X"18",X"C7",X"CD",X"18",X"C7",X"F1",X"E1",X"DD",X"CB",X"14",X"46",X"28",X"0A",X"DD",X"CB",X"14",
		X"6E",X"28",X"04",X"DD",X"CB",X"00",X"FE",X"CD",X"8F",X"21",X"EB",X"CD",X"8F",X"21",X"EB",X"DD",
		X"74",X"07",X"DD",X"75",X"06",X"DD",X"72",X"0D",X"DD",X"73",X"0C",X"F1",X"E6",X"0E",X"4F",X"06",
		X"00",X"21",X"99",X"23",X"09",X"5E",X"23",X"56",X"21",X"8E",X"21",X"E5",X"EB",X"E9",X"C9",X"F5",
		X"7C",X"2F",X"67",X"7D",X"2F",X"6F",X"23",X"F1",X"C9",X"00",X"00",X"FF",X"3F",X"00",X"10",X"1C",
		X"07",X"00",X"04",X"8F",X"02",X"C7",X"01",X"4E",X"01",X"00",X"01",X"CA",X"00",X"A4",X"00",X"87",
		X"00",X"72",X"00",X"61",X"00",X"54",X"00",X"49",X"00",X"00",X"00",X"A1",X"16",X"73",X"0B",X"12",
		X"06",X"A7",X"03",X"6A",X"02",X"B5",X"01",X"44",X"01",X"FA",X"00",X"C7",X"00",X"A1",X"00",X"86",
		X"00",X"71",X"00",X"60",X"00",X"53",X"00",X"48",X"00",X"00",X"00",X"B9",X"05",X"A8",X"05",X"19",
		X"04",X"DD",X"02",X"0D",X"02",X"85",X"01",X"29",X"01",X"EA",X"00",X"BC",X"00",X"9A",X"00",X"81",
		X"00",X"6D",X"00",X"5E",X"00",X"51",X"00",X"47",X"00",X"00",X"00",X"06",X"02",X"BB",X"02",X"84",
		X"02",X"0C",X"02",X"9D",X"01",X"46",X"01",X"04",X"01",X"D2",X"00",X"AD",X"00",X"90",X"00",X"7A",
		X"00",X"68",X"00",X"5A",X"00",X"4E",X"00",X"45",X"00",X"00",X"00",X"EA",X"00",X"6E",X"01",X"89",
		X"01",X"6A",X"01",X"D5",X"00",X"06",X"01",X"DB",X"00",X"B7",X"00",X"9A",X"00",X"83",X"00",X"70",
		X"00",X"61",X"00",X"55",X"00",X"4A",X"00",X"42",X"00",X"00",X"00",X"7C",X"00",X"D2",X"00",X"F8",
		X"00",X"FA",X"00",X"E8",X"00",X"CE",X"00",X"B4",X"00",X"9C",X"00",X"87",X"00",X"75",X"00",X"66",
		X"00",X"59",X"00",X"4F",X"00",X"46",X"00",X"3E",X"00",X"00",X"00",X"49",X"00",X"82",X"00",X"A3",
		X"00",X"AF",X"00",X"AC",X"00",X"A1",X"00",X"92",X"00",X"83",X"00",X"75",X"00",X"67",X"00",X"5C",
		X"00",X"51",X"00",X"49",X"00",X"41",X"00",X"3A",X"00",X"00",X"00",X"2E",X"00",X"55",X"00",X"6F",
		X"00",X"7D",X"00",X"81",X"00",X"7D",X"00",X"76",X"00",X"6D",X"00",X"63",X"00",X"5A",X"00",X"51",
		X"00",X"49",X"00",X"42",X"00",X"3C",X"00",X"36",X"00",X"00",X"00",X"1F",X"00",X"3A",X"00",X"4F",
		X"00",X"5C",X"00",X"62",X"00",X"62",X"00",X"5F",X"00",X"5B",X"00",X"54",X"00",X"4E",X"00",X"48",
		X"00",X"42",X"00",X"3C",X"00",X"37",X"00",X"32",X"00",X"00",X"00",X"16",X"00",X"2A",X"00",X"3A",
		X"00",X"45",X"00",X"4B",X"00",X"4E",X"00",X"4D",X"00",X"4B",X"00",X"48",X"00",X"43",X"00",X"3F",
		X"00",X"3A",X"00",X"36",X"00",X"32",X"00",X"2E",X"00",X"00",X"00",X"10",X"00",X"1F",X"00",X"2B",
		X"00",X"34",X"00",X"3B",X"00",X"3E",X"00",X"3F",X"00",X"3E",X"00",X"3D",X"00",X"3A",X"00",X"37",
		X"00",X"34",X"00",X"30",X"00",X"2D",X"00",X"2A",X"00",X"00",X"00",X"0C",X"00",X"17",X"00",X"17",
		X"00",X"29",X"00",X"2E",X"00",X"32",X"00",X"34",X"00",X"34",X"00",X"33",X"00",X"32",X"00",X"30",
		X"00",X"2E",X"00",X"2B",X"00",X"29",X"00",X"26",X"00",X"00",X"00",X"09",X"00",X"12",X"00",X"1A",
		X"00",X"20",X"00",X"25",X"00",X"29",X"00",X"2B",X"00",X"2C",X"00",X"2C",X"00",X"2B",X"00",X"2A",
		X"00",X"28",X"00",X"26",X"00",X"25",X"00",X"23",X"00",X"00",X"00",X"07",X"00",X"0E",X"00",X"15",
		X"00",X"1A",X"00",X"1E",X"00",X"21",X"00",X"24",X"00",X"25",X"00",X"25",X"00",X"25",X"00",X"24",
		X"00",X"24",X"00",X"22",X"00",X"21",X"00",X"1F",X"00",X"00",X"00",X"06",X"00",X"0C",X"00",X"11",
		X"00",X"15",X"00",X"19",X"00",X"1C",X"00",X"1E",X"00",X"1F",X"00",X"20",X"00",X"20",X"00",X"20",
		X"00",X"1F",X"00",X"1F",X"00",X"1E",X"00",X"1C",X"00",X"00",X"00",X"05",X"00",X"09",X"00",X"0E",
		X"00",X"12",X"00",X"15",X"00",X"17",X"00",X"19",X"00",X"1B",X"00",X"1C",X"00",X"1C",X"00",X"1C",
		X"00",X"1C",X"00",X"1B",X"00",X"1B",X"00",X"1A",X"00",X"80",X"3C",X"66",X"3D",X"7C",X"3D",X"92",
		X"3D",X"A8",X"3D",X"A8",X"3D",X"A8",X"3D",X"A8",X"3D",X"A8",X"3D",X"DD",X"21",X"BB",X"23",X"ED",
		X"4B",X"9B",X"F8",X"CD",X"BB",X"23",X"ED",X"43",X"9B",X"F8",X"C9",X"0A",X"03",X"26",X"00",X"87",
		X"6F",X"11",X"CA",X"23",X"19",X"7E",X"23",X"66",X"6F",X"E9",X"EA",X"23",X"F5",X"23",X"F6",X"23",
		X"01",X"24",X"0D",X"24",X"17",X"24",X"23",X"24",X"2F",X"24",X"40",X"24",X"4A",X"24",X"56",X"24",
		X"64",X"24",X"7D",X"24",X"8D",X"24",X"A2",X"24",X"B5",X"24",X"0B",X"21",X"00",X"00",X"22",X"9D",
		X"F8",X"22",X"9F",X"F8",X"C9",X"C9",X"0A",X"03",X"6F",X"87",X"9F",X"67",X"09",X"44",X"4D",X"DD",
		X"E9",X"0A",X"03",X"6F",X"0A",X"03",X"67",X"35",X"20",X"EC",X"03",X"DD",X"E9",X"0A",X"03",X"6F",
		X"0A",X"03",X"67",X"5E",X"C3",X"26",X"24",X"0A",X"03",X"6F",X"0A",X"03",X"67",X"5E",X"23",X"56",
		X"C3",X"35",X"24",X"0A",X"03",X"5F",X"0A",X"03",X"6F",X"0A",X"03",X"67",X"73",X"DD",X"E9",X"0A",
		X"03",X"5F",X"0A",X"03",X"57",X"0A",X"03",X"6F",X"0A",X"03",X"67",X"73",X"23",X"72",X"DD",X"E9",
		X"0A",X"03",X"6F",X"0A",X"03",X"67",X"5E",X"C3",X"59",X"24",X"0A",X"03",X"6F",X"0A",X"03",X"67",
		X"5E",X"23",X"56",X"C3",X"6A",X"24",X"0A",X"03",X"5F",X"0A",X"03",X"6F",X"0A",X"03",X"67",X"7E",
		X"83",X"77",X"DD",X"E9",X"0A",X"03",X"5F",X"0A",X"03",X"57",X"0A",X"03",X"6F",X"0A",X"03",X"67",
		X"E5",X"7E",X"23",X"66",X"6F",X"19",X"EB",X"E1",X"73",X"23",X"72",X"DD",X"E9",X"0A",X"03",X"5F",
		X"0A",X"03",X"6F",X"0A",X"03",X"67",X"CB",X"2E",X"1D",X"20",X"FB",X"DD",X"E9",X"0A",X"03",X"5F",
		X"0A",X"03",X"6F",X"0A",X"03",X"67",X"23",X"CB",X"2E",X"2B",X"CB",X"1E",X"23",X"1D",X"20",X"F7",
		X"DD",X"E9",X"0A",X"03",X"5F",X"0A",X"03",X"6F",X"0A",X"03",X"67",X"0A",X"77",X"23",X"03",X"1D",
		X"C2",X"AB",X"24",X"DD",X"E9",X"0A",X"03",X"87",X"C3",X"A4",X"24",X"63",X"2A",X"AE",X"F8",X"7C",
		X"B5",X"C0",X"EB",X"22",X"AE",X"F8",X"C9",X"DD",X"21",X"73",X"40",X"DD",X"36",X"00",X"80",X"21",
		X"A3",X"40",X"F9",X"CD",X"0B",X"28",X"3A",X"B5",X"43",X"FE",X"01",X"3E",X"DD",X"28",X"02",X"3E",
		X"EE",X"32",X"EB",X"43",X"21",X"56",X"F9",X"22",X"5A",X"F9",X"21",X"00",X"00",X"22",X"58",X"F9",
		X"DD",X"36",X"0B",X"6C",X"DD",X"36",X"11",X"64",X"AF",X"CD",X"B8",X"26",X"DD",X"36",X"00",X"02",
		X"DD",X"CB",X"14",X"C6",X"FD",X"E5",X"DD",X"E5",X"E1",X"CD",X"D1",X"2B",X"DD",X"CB",X"00",X"E6",
		X"CD",X"EF",X"CB",X"FD",X"E1",X"CD",X"28",X"28",X"01",X"FF",X"FF",X"DD",X"21",X"77",X"40",X"DD",
		X"CB",X"00",X"7E",X"C2",X"E1",X"26",X"FD",X"E5",X"CD",X"EF",X"CB",X"FD",X"E1",X"DD",X"7E",X"15",
		X"B7",X"28",X"03",X"DD",X"35",X"15",X"3A",X"E1",X"43",X"B7",X"28",X"4E",X"2A",X"E2",X"43",X"7E",
		X"23",X"22",X"E2",X"43",X"B7",X"CA",X"D4",X"C9",X"4F",X"E6",X"C0",X"79",X"28",X"38",X"E6",X"3F",
		X"47",X"21",X"EE",X"43",X"DD",X"CB",X"00",X"7E",X"C2",X"E1",X"26",X"CB",X"79",X"28",X"02",X"34",
		X"34",X"CB",X"71",X"28",X"02",X"35",X"35",X"C5",X"7E",X"CB",X"3F",X"CB",X"3F",X"CD",X"B8",X"26",
		X"CD",X"4B",X"28",X"DD",X"21",X"77",X"40",X"DD",X"7E",X"15",X"B7",X"28",X"03",X"DD",X"35",X"15",
		X"C1",X"10",X"CE",X"C3",X"1B",X"25",X"E6",X"17",X"18",X"30",X"CD",X"AD",X"26",X"DB",X"48",X"CD",
		X"2A",X"C7",X"28",X"02",X"DB",X"4A",X"2F",X"57",X"A8",X"F6",X"80",X"A2",X"42",X"08",X"21",X"FE",
		X"43",X"DB",X"49",X"2F",X"E6",X"08",X"BE",X"77",X"28",X"0F",X"CB",X"5F",X"28",X"0B",X"CD",X"4E",
		X"3F",X"3A",X"EE",X"43",X"C6",X"7F",X"32",X"EE",X"43",X"08",X"C5",X"CB",X"77",X"C2",X"65",X"26",
		X"DD",X"36",X"09",X"00",X"DD",X"36",X"08",X"00",X"DD",X"36",X"0F",X"00",X"DD",X"36",X"0E",X"00",
		X"DD",X"36",X"07",X"00",X"DD",X"36",X"06",X"00",X"DD",X"36",X"0D",X"00",X"DD",X"36",X"0C",X"00",
		X"06",X"00",X"CB",X"7F",X"F5",X"C4",X"FB",X"25",X"F1",X"06",X"01",X"CB",X"6F",X"F5",X"C4",X"FB",
		X"25",X"F1",X"3E",X"01",X"CD",X"40",X"28",X"C1",X"C3",X"1B",X"25",X"FD",X"7E",X"19",X"B7",X"C0",
		X"78",X"FE",X"01",X"20",X"29",X"3A",X"ED",X"43",X"CD",X"60",X"26",X"FE",X"04",X"38",X"09",X"D9",
		X"11",X"FA",X"C0",X"CD",X"BC",X"24",X"D9",X"C9",X"CD",X"CB",X"27",X"D0",X"3A",X"ED",X"43",X"3C",
		X"32",X"ED",X"43",X"CB",X"FF",X"CD",X"9A",X"C5",X"CD",X"67",X"3A",X"C3",X"58",X"26",X"3A",X"F3",
		X"43",X"CD",X"60",X"26",X"FE",X"04",X"38",X"0F",X"3A",X"C1",X"43",X"FE",X"1F",X"D0",X"D9",X"11",
		X"C1",X"C0",X"CD",X"BC",X"24",X"D9",X"C9",X"CD",X"CB",X"27",X"D0",X"3A",X"F3",X"43",X"3C",X"32",
		X"F3",X"43",X"CD",X"9A",X"C5",X"CD",X"90",X"3B",X"FD",X"21",X"86",X"16",X"CD",X"28",X"28",X"C9",
		X"FE",X"FF",X"C0",X"AF",X"C9",X"3A",X"EE",X"43",X"CB",X"3F",X"CB",X"3F",X"E6",X"3F",X"CB",X"27",
		X"5F",X"16",X"00",X"21",X"1E",X"18",X"19",X"19",X"19",X"23",X"23",X"5E",X"23",X"56",X"06",X"05",
		X"CB",X"2A",X"CB",X"1B",X"10",X"FA",X"DD",X"73",X"06",X"DD",X"72",X"07",X"23",X"5E",X"23",X"56",
		X"06",X"05",X"CB",X"2A",X"CB",X"1B",X"10",X"FA",X"DD",X"73",X"0C",X"DD",X"72",X"0D",X"DD",X"CB",
		X"00",X"D6",X"DD",X"CB",X"00",X"DE",X"DD",X"CB",X"00",X"E6",X"C3",X"F2",X"25",X"3A",X"EE",X"43",
		X"CB",X"3F",X"CB",X"3F",X"B9",X"CA",X"D8",X"26",X"CD",X"DE",X"C5",X"4F",X"21",X"00",X"00",X"16",
		X"00",X"5F",X"19",X"29",X"29",X"29",X"29",X"29",X"11",X"86",X"08",X"19",X"22",X"56",X"F9",X"21",
		X"56",X"F9",X"DD",X"75",X"12",X"DD",X"74",X"13",X"DD",X"7E",X"00",X"F6",X"03",X"DD",X"77",X"00",
		X"C9",X"CD",X"E3",X"3A",X"3E",X"09",X"32",X"E4",X"43",X"FD",X"36",X"04",X"01",X"CD",X"4B",X"28",
		X"3E",X"0A",X"32",X"F0",X"43",X"DD",X"21",X"A3",X"40",X"11",X"30",X"00",X"3E",X"08",X"DD",X"36",
		X"04",X"01",X"DD",X"CB",X"00",X"7E",X"28",X"04",X"DD",X"36",X"00",X"81",X"DD",X"19",X"3D",X"20",
		X"ED",X"CD",X"4B",X"28",X"21",X"A3",X"40",X"01",X"00",X"80",X"71",X"23",X"10",X"FC",X"DD",X"21",
		X"A3",X"40",X"3E",X"08",X"08",X"DD",X"E5",X"E1",X"01",X"00",X"30",X"71",X"23",X"10",X"FC",X"DD",
		X"36",X"00",X"81",X"DD",X"E5",X"E1",X"11",X"2E",X"00",X"19",X"DD",X"75",X"02",X"DD",X"74",X"03",
		X"11",X"04",X"00",X"DD",X"19",X"DD",X"CB",X"00",X"CE",X"CD",X"A5",X"27",X"FD",X"7E",X"0F",X"80",
		X"DD",X"77",X"0B",X"FD",X"7E",X"15",X"81",X"DD",X"77",X"11",X"21",X"C8",X"19",X"DD",X"75",X"12",
		X"DD",X"74",X"13",X"11",X"2C",X"00",X"DD",X"19",X"21",X"8E",X"27",X"DD",X"74",X"FF",X"DD",X"75",
		X"FE",X"08",X"3D",X"20",X"AF",X"3E",X"2D",X"CD",X"40",X"28",X"FD",X"7E",X"01",X"B7",X"28",X"05",
		X"CD",X"4B",X"28",X"18",X"F5",X"FD",X"36",X"00",X"00",X"CD",X"4B",X"28",X"18",X"F7",X"FD",X"CB",
		X"04",X"D6",X"FD",X"E5",X"DD",X"E1",X"11",X"04",X"00",X"DD",X"19",X"CD",X"AA",X"20",X"3E",X"02",
		X"CD",X"40",X"28",X"18",X"ED",X"08",X"57",X"08",X"01",X"02",X"02",X"CB",X"52",X"20",X"0C",X"CB",
		X"4A",X"20",X"02",X"06",X"06",X"CB",X"42",X"C8",X"0E",X"06",X"C9",X"01",X"04",X"07",X"CB",X"4A",
		X"20",X"02",X"06",X"01",X"CB",X"42",X"C8",X"78",X"41",X"4F",X"C9",X"21",X"EB",X"27",X"E5",X"D1",
		X"7E",X"23",X"66",X"6F",X"E5",X"E1",X"B4",X"C8",X"7E",X"B7",X"28",X"06",X"13",X"13",X"D5",X"E1",
		X"18",X"EE",X"E5",X"DD",X"E1",X"DD",X"36",X"00",X"80",X"37",X"C9",X"A3",X"40",X"D3",X"40",X"03",
		X"41",X"33",X"41",X"63",X"41",X"93",X"41",X"C3",X"41",X"F3",X"41",X"23",X"42",X"53",X"42",X"83",
		X"42",X"B3",X"42",X"E3",X"42",X"13",X"43",X"43",X"43",X"00",X"00",X"D9",X"DD",X"E5",X"E1",X"22",
		X"88",X"F8",X"AF",X"CB",X"C6",X"23",X"77",X"23",X"77",X"23",X"77",X"23",X"E5",X"77",X"06",X"15",
		X"23",X"77",X"10",X"FC",X"DD",X"E1",X"D9",X"C9",X"21",X"00",X"00",X"39",X"31",X"86",X"F8",X"FD",
		X"E5",X"FD",X"2A",X"88",X"F8",X"FD",X"22",X"8C",X"F8",X"FD",X"75",X"02",X"FD",X"74",X"03",X"C9",
		X"FD",X"2A",X"88",X"F8",X"FD",X"77",X"01",X"FD",X"36",X"00",X"82",X"21",X"00",X"00",X"39",X"31",
		X"86",X"F8",X"FD",X"2A",X"88",X"F8",X"FD",X"75",X"02",X"FD",X"74",X"03",X"2A",X"8C",X"F8",X"7C",
		X"B5",X"28",X"10",X"FD",X"2A",X"8C",X"F8",X"21",X"00",X"00",X"22",X"8C",X"F8",X"FD",X"22",X"88",
		X"F8",X"18",X"04",X"FD",X"2A",X"88",X"F8",X"01",X"30",X"00",X"FD",X"09",X"FD",X"E5",X"E1",X"01",
		X"73",X"43",X"B7",X"ED",X"42",X"38",X"04",X"FD",X"21",X"43",X"40",X"FD",X"CB",X"00",X"46",X"28",
		X"E6",X"FD",X"22",X"88",X"F8",X"FD",X"E5",X"E1",X"11",X"04",X"00",X"19",X"E5",X"CD",X"4E",X"2C",
		X"E1",X"CD",X"D1",X"2B",X"FD",X"2A",X"88",X"F8",X"FD",X"66",X"03",X"FD",X"6E",X"02",X"F9",X"C9",
		X"D9",X"D1",X"01",X"30",X"00",X"DD",X"E5",X"E1",X"09",X"F9",X"D5",X"D9",X"C9",X"D9",X"DD",X"E5",
		X"E1",X"06",X"05",X"AF",X"77",X"2B",X"10",X"FC",X"D9",X"C9",X"CD",X"65",X"1E",X"CD",X"3B",X"CB",
		X"CD",X"10",X"C3",X"CD",X"89",X"29",X"CD",X"99",X"C7",X"FB",X"FD",X"21",X"E4",X"28",X"CD",X"28",
		X"28",X"C3",X"EB",X"28",X"FD",X"21",X"73",X"28",X"C3",X"C7",X"24",X"DD",X"21",X"73",X"40",X"DD",
		X"CB",X"00",X"7E",X"C8",X"21",X"E4",X"43",X"3A",X"BF",X"43",X"B6",X"C8",X"3A",X"E1",X"43",X"B7",
		X"28",X"09",X"CD",X"83",X"1D",X"CD",X"9F",X"1D",X"C2",X"E3",X"1A",X"FD",X"2A",X"88",X"F8",X"FD",
		X"7E",X"01",X"B7",X"C2",X"64",X"29",X"CD",X"72",X"C5",X"FD",X"36",X"01",X"06",X"FD",X"CB",X"00",
		X"CE",X"CD",X"5F",X"C7",X"30",X"07",X"FD",X"21",X"B3",X"29",X"CD",X"28",X"28",X"21",X"F4",X"43",
		X"34",X"7E",X"FE",X"09",X"20",X"2E",X"AF",X"77",X"06",X"0C",X"21",X"E6",X"F8",X"3A",X"E1",X"43",
		X"B7",X"20",X"21",X"CD",X"A1",X"32",X"CD",X"37",X"C0",X"21",X"FD",X"43",X"34",X"7E",X"FE",X"28",
		X"38",X"12",X"3E",X"1A",X"77",X"21",X"BF",X"43",X"7E",X"FE",X"99",X"28",X"07",X"C6",X"01",X"27",
		X"77",X"CD",X"7B",X"C5",X"CD",X"4B",X"28",X"C3",X"EB",X"28",X"21",X"73",X"40",X"06",X"0F",X"11",
		X"2C",X"00",X"AF",X"77",X"23",X"23",X"23",X"23",X"77",X"19",X"10",X"F7",X"21",X"43",X"40",X"22",
		X"88",X"F8",X"21",X"00",X"00",X"22",X"8C",X"F8",X"C9",X"21",X"00",X"08",X"11",X"07",X"00",X"3A",
		X"BE",X"43",X"E6",X"0F",X"BE",X"28",X"07",X"3E",X"FF",X"BE",X"C8",X"19",X"18",X"F1",X"23",X"01",
		X"07",X"00",X"11",X"F7",X"43",X"ED",X"B0",X"C9",X"2A",X"AE",X"F8",X"7C",X"B5",X"C0",X"EB",X"22",
		X"AE",X"F8",X"C9",X"CD",X"8B",X"3E",X"21",X"E4",X"43",X"34",X"CD",X"B0",X"28",X"CD",X"0B",X"28",
		X"CD",X"A4",X"2A",X"CD",X"07",X"2A",X"DD",X"CB",X"14",X"C6",X"DD",X"CB",X"00",X"CE",X"DD",X"E5",
		X"E1",X"FD",X"E5",X"CD",X"D1",X"2B",X"FD",X"E1",X"DD",X"CB",X"00",X"D6",X"DD",X"E5",X"3E",X"09",
		X"CD",X"40",X"28",X"3E",X"01",X"CD",X"40",X"28",X"DD",X"E1",X"DD",X"CB",X"00",X"76",X"20",X"21",
		X"CD",X"AA",X"20",X"DD",X"E5",X"DD",X"22",X"F1",X"43",X"CD",X"15",X"C8",X"30",X"07",X"FD",X"21",
		X"FC",X"C9",X"CD",X"28",X"28",X"18",X"DC",X"2A",X"F7",X"43",X"DD",X"75",X"12",X"DD",X"74",X"13",
		X"C9",X"21",X"00",X"00",X"39",X"31",X"86",X"F8",X"E5",X"DD",X"E5",X"21",X"BF",X"43",X"7E",X"3D",
		X"27",X"77",X"CD",X"34",X"3B",X"E1",X"11",X"0B",X"00",X"19",X"7E",X"D6",X"04",X"77",X"11",X"06",
		X"00",X"19",X"7E",X"D6",X"06",X"77",X"23",X"3A",X"F9",X"43",X"4F",X"3A",X"FA",X"43",X"47",X"71",
		X"23",X"70",X"23",X"36",X"01",X"23",X"36",X"01",X"3A",X"BE",X"43",X"FA",X"51",X"2A",X"C6",X"04",
		X"27",X"F5",X"E6",X"0F",X"4F",X"06",X"01",X"CD",X"C3",X"2E",X"F1",X"CB",X"3F",X"CB",X"3F",X"CB",
		X"3F",X"CB",X"3F",X"28",X"06",X"4F",X"06",X"02",X"CD",X"C3",X"2E",X"CD",X"E8",X"C6",X"CD",X"E8",
		X"C6",X"CD",X"E8",X"C6",X"E1",X"F9",X"2A",X"FB",X"43",X"DD",X"7E",X"04",X"BD",X"20",X"06",X"DD",
		X"7E",X"05",X"BC",X"28",X"0E",X"CD",X"AA",X"20",X"DD",X"E5",X"3E",X"01",X"CD",X"40",X"28",X"DD",
		X"E1",X"18",X"E3",X"CD",X"BD",X"28",X"21",X"E4",X"43",X"35",X"2A",X"88",X"F8",X"CB",X"86",X"CD",
		X"4B",X"28",X"18",X"F6",X"3A",X"E1",X"43",X"B7",X"C2",X"62",X"2B",X"CD",X"7C",X"2E",X"17",X"17",
		X"17",X"E6",X"03",X"CA",X"48",X"2B",X"3D",X"CA",X"55",X"2B",X"3D",X"28",X"68",X"18",X"45",X"DD",
		X"70",X"0B",X"DD",X"71",X"11",X"CD",X"7C",X"2E",X"E6",X"0F",X"08",X"3A",X"BE",X"43",X"FE",X"07",
		X"38",X"02",X"3E",X"07",X"47",X"08",X"CB",X"27",X"F6",X"01",X"10",X"FA",X"F6",X"10",X"6F",X"CD",
		X"7C",X"2E",X"26",X"00",X"B7",X"F2",X"EB",X"2A",X"CD",X"8F",X"21",X"DD",X"75",X"08",X"DD",X"74",
		X"09",X"CD",X"7C",X"2E",X"26",X"00",X"B7",X"F2",X"FD",X"2A",X"CD",X"8F",X"21",X"DD",X"75",X"0E",
		X"DD",X"74",X"0F",X"C9",X"06",X"09",X"CD",X"7C",X"2E",X"FE",X"CD",X"D2",X"06",X"2B",X"4F",X"FE",
		X"28",X"30",X"06",X"11",X"E0",X"C0",X"CD",X"A8",X"29",X"FE",X"B4",X"38",X"A2",X"11",X"D9",X"C0",
		X"CD",X"A8",X"29",X"18",X"9A",X"06",X"C0",X"CD",X"7C",X"2E",X"FE",X"CD",X"D2",X"27",X"2B",X"4F",
		X"FE",X"28",X"30",X"06",X"11",X"CB",X"C0",X"CD",X"A8",X"29",X"FE",X"B4",X"DA",X"BF",X"2A",X"11",
		X"D2",X"C0",X"CD",X"A8",X"29",X"C3",X"BF",X"2A",X"0E",X"09",X"CD",X"7C",X"2E",X"FE",X"C0",X"30",
		X"F9",X"47",X"C3",X"BF",X"2A",X"0E",X"CD",X"CD",X"7C",X"2E",X"FE",X"C0",X"30",X"F9",X"47",X"C3",
		X"BF",X"2A",X"DD",X"36",X"0B",X"A0",X"DD",X"36",X"11",X"CD",X"DD",X"36",X"08",X"80",X"DD",X"36",
		X"09",X"FF",X"DD",X"36",X"0E",X"80",X"DD",X"36",X"0E",X"FF",X"C9",X"F3",X"ED",X"73",X"8A",X"F8",
		X"31",X"40",X"F8",X"F5",X"08",X"F5",X"C5",X"D5",X"E5",X"DD",X"E5",X"FD",X"E5",X"DB",X"4E",X"1F",
		X"38",X"22",X"CD",X"03",X"C1",X"21",X"B5",X"F8",X"7E",X"23",X"46",X"A8",X"4F",X"DB",X"49",X"2F",
		X"77",X"2B",X"70",X"A1",X"E6",X"E0",X"2B",X"87",X"D2",X"AF",X"2B",X"34",X"C3",X"A6",X"2B",X"C2",
		X"A6",X"2B",X"18",X"03",X"CD",X"D2",X"2C",X"FD",X"E1",X"DD",X"E1",X"E1",X"D1",X"C1",X"F1",X"08",
		X"3E",X"01",X"D3",X"4F",X"3E",X"3F",X"ED",X"47",X"ED",X"5E",X"F1",X"ED",X"7B",X"8A",X"F8",X"FB",
		X"C9",X"E5",X"FD",X"E1",X"CB",X"46",X"CA",X"ED",X"2B",X"CB",X"86",X"E5",X"23",X"7E",X"D3",X"4B",
		X"23",X"5E",X"23",X"56",X"23",X"7E",X"23",X"66",X"6F",X"CD",X"07",X"2D",X"E1",X"CB",X"4E",X"C8",
		X"CB",X"8E",X"E5",X"11",X"0B",X"00",X"19",X"7E",X"11",X"06",X"00",X"19",X"56",X"5F",X"23",X"EB",
		X"06",X"90",X"CD",X"68",X"2F",X"FD",X"77",X"01",X"EB",X"7E",X"23",X"66",X"6F",X"7E",X"23",X"66",
		X"6F",X"7E",X"CB",X"7F",X"28",X"19",X"23",X"E6",X"7F",X"47",X"7E",X"23",X"4F",X"EB",X"3A",X"EC",
		X"43",X"B7",X"CA",X"2A",X"2C",X"ED",X"42",X"C3",X"2E",X"2C",X"09",X"C3",X"2E",X"2C",X"EB",X"FD",
		X"75",X"04",X"FD",X"74",X"05",X"FD",X"73",X"02",X"FD",X"72",X"03",X"CD",X"07",X"2D",X"E1",X"DB",
		X"4E",X"CB",X"7F",X"C8",X"CB",X"FE",X"FD",X"E5",X"DD",X"E1",X"CD",X"D5",X"17",X"C9",X"CB",X"56",
		X"C8",X"E5",X"FD",X"E1",X"11",X"06",X"00",X"19",X"1E",X"C2",X"16",X"06",X"FD",X"7E",X"0B",X"BA",
		X"38",X"03",X"BB",X"38",X"06",X"CD",X"74",X"2D",X"C3",X"85",X"2C",X"5E",X"23",X"56",X"23",X"4E",
		X"23",X"46",X"EB",X"09",X"EB",X"2B",X"73",X"23",X"72",X"23",X"4E",X"23",X"46",X"EB",X"09",X"EB",
		X"2B",X"73",X"23",X"72",X"23",X"1E",X"CF",X"16",X"06",X"FD",X"7E",X"11",X"BA",X"38",X"03",X"BB",
		X"38",X"06",X"CD",X"74",X"2D",X"C3",X"B2",X"2C",X"5E",X"23",X"56",X"23",X"4E",X"23",X"46",X"EB",
		X"09",X"EB",X"2B",X"73",X"23",X"72",X"23",X"4E",X"23",X"46",X"EB",X"09",X"EB",X"2B",X"73",X"23",
		X"72",X"23",X"5E",X"23",X"56",X"13",X"13",X"EB",X"7E",X"23",X"B6",X"2B",X"C2",X"C5",X"2C",X"23",
		X"23",X"7E",X"23",X"66",X"6F",X"EB",X"72",X"2B",X"73",X"3E",X"07",X"FD",X"B6",X"00",X"FD",X"77",
		X"00",X"C9",X"21",X"43",X"40",X"06",X"11",X"11",X"30",X"00",X"CB",X"4E",X"28",X"09",X"23",X"35",
		X"2B",X"20",X"04",X"CB",X"8E",X"CB",X"C6",X"19",X"10",X"F0",X"C9",X"2A",X"86",X"F8",X"7C",X"B5",
		X"28",X"0E",X"01",X"77",X"43",X"11",X"30",X"00",X"19",X"E5",X"B7",X"ED",X"42",X"E1",X"38",X"03",
		X"21",X"77",X"40",X"22",X"86",X"F8",X"C9",X"CB",X"7A",X"C0",X"06",X"00",X"7E",X"23",X"3D",X"CA",
		X"47",X"2D",X"3A",X"EC",X"43",X"B7",X"7E",X"23",X"C2",X"31",X"2D",X"01",X"1E",X"00",X"EB",X"08",
		X"1A",X"13",X"77",X"23",X"1A",X"13",X"77",X"23",X"36",X"00",X"08",X"09",X"3D",X"C2",X"1F",X"2D",
		X"C9",X"01",X"E2",X"FF",X"EB",X"08",X"1A",X"13",X"77",X"2B",X"1A",X"13",X"77",X"2B",X"36",X"00",
		X"08",X"09",X"3D",X"C2",X"35",X"2D",X"C9",X"3A",X"EC",X"43",X"B7",X"7E",X"23",X"C2",X"62",X"2D",
		X"01",X"1F",X"00",X"EB",X"08",X"1A",X"13",X"77",X"23",X"36",X"00",X"08",X"09",X"3D",X"C2",X"54",
		X"2D",X"C9",X"01",X"E1",X"FF",X"EB",X"08",X"1A",X"13",X"77",X"2B",X"36",X"00",X"08",X"09",X"3D",
		X"C2",X"66",X"2D",X"C9",X"FD",X"CB",X"14",X"46",X"20",X"0A",X"E1",X"FD",X"36",X"00",X"01",X"FD",
		X"CB",X"14",X"FE",X"C9",X"FD",X"CB",X"14",X"6E",X"28",X"05",X"FD",X"35",X"15",X"28",X"EB",X"36",
		X"00",X"23",X"36",X"00",X"23",X"7E",X"23",X"2F",X"4F",X"7E",X"2F",X"47",X"03",X"70",X"2B",X"71",
		X"23",X"23",X"36",X"00",X"23",X"1D",X"CB",X"78",X"C2",X"AD",X"2D",X"1E",X"06",X"73",X"23",X"C9",
		X"2A",X"AF",X"43",X"22",X"E6",X"43",X"3A",X"B1",X"43",X"32",X"E8",X"43",X"21",X"00",X"00",X"22",
		X"AF",X"43",X"22",X"B0",X"43",X"2A",X"CF",X"43",X"E5",X"21",X"18",X"2E",X"22",X"E2",X"43",X"22",
		X"CF",X"43",X"3E",X"FF",X"32",X"E1",X"43",X"01",X"0D",X"00",X"11",X"B5",X"43",X"21",X"0B",X"2E",
		X"ED",X"B0",X"AF",X"32",X"E4",X"43",X"32",X"F0",X"43",X"32",X"F3",X"43",X"32",X"ED",X"43",X"32",
		X"EE",X"43",X"CD",X"CA",X"28",X"E1",X"F5",X"22",X"CF",X"43",X"CD",X"7C",X"2E",X"2A",X"E6",X"43",
		X"22",X"AF",X"43",X"2A",X"E7",X"43",X"22",X"B0",X"43",X"F1",X"C9",X"01",X"01",X"30",X"00",X"02",
		X"28",X"28",X"28",X"00",X"01",X"08",X"40",X"40",X"B0",X"84",X"90",X"00",X"00",X"FF",X"4C",X"C6",
		X"02",X"C6",X"02",X"C6",X"02",X"FF",X"FF",X"81",X"02",X"C4",X"02",X"C4",X"02",X"C4",X"02",X"C3",
		X"FF",X"00",X"87",X"01",X"44",X"01",X"44",X"01",X"44",X"01",X"FF",X"FF",X"91",X"02",X"44",X"02",
		X"44",X"02",X"44",X"02",X"5F",X"02",X"C4",X"02",X"C4",X"00",X"5F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"02",X"FF",X"FF",X"02",X"FF",X"02",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"9F",X"C3",X"00",
		X"A2",X"FF",X"10",X"FF",X"10",X"02",X"45",X"02",X"45",X"02",X"C4",X"02",X"FF",X"10",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"E5",X"2A",X"CF",X"43",
		X"54",X"5D",X"29",X"19",X"29",X"19",X"29",X"29",X"29",X"29",X"19",X"11",X"53",X"31",X"19",X"22",
		X"CF",X"43",X"7C",X"E1",X"C9",X"AF",X"32",X"E0",X"43",X"11",X"00",X"D5",X"21",X"AF",X"43",X"06",
		X"06",X"CD",X"A0",X"2F",X"3A",X"E9",X"43",X"FE",X"02",X"C0",X"11",X"B0",X"D5",X"21",X"B2",X"43",
		X"06",X"06",X"CD",X"A0",X"2F",X"C9",X"3A",X"B5",X"43",X"FE",X"02",X"21",X"B2",X"43",X"C8",X"21",
		X"AF",X"43",X"C9",X"3E",X"FF",X"32",X"E0",X"43",X"1E",X"04",X"CD",X"B6",X"2E",X"23",X"23",X"23",
		X"CB",X"38",X"08",X"04",X"2B",X"1D",X"10",X"FC",X"08",X"30",X"08",X"CB",X"21",X"CB",X"21",X"CB",
		X"21",X"CB",X"21",X"CD",X"F2",X"2E",X"79",X"86",X"27",X"77",X"D0",X"2B",X"1D",X"C8",X"0E",X"01",
		X"18",X"F1",X"08",X"7B",X"FE",X"02",X"20",X"19",X"7E",X"E6",X"0F",X"81",X"27",X"E6",X"F0",X"28",
		X"10",X"D9",X"CD",X"20",X"2F",X"3A",X"BD",X"43",X"3C",X"B8",X"CC",X"13",X"2F",X"32",X"BD",X"43",
		X"D9",X"08",X"C9",X"21",X"B6",X"43",X"7E",X"C6",X"01",X"27",X"77",X"CD",X"14",X"3E",X"AF",X"C9",
		X"06",X"0A",X"DB",X"61",X"E6",X"F8",X"C8",X"06",X"0F",X"CB",X"5F",X"C0",X"06",X"14",X"CB",X"67",
		X"C0",X"06",X"1E",X"CB",X"6F",X"C0",X"06",X"28",X"CB",X"77",X"C0",X"06",X"32",X"CB",X"7F",X"C0",
		X"E1",X"46",X"23",X"5E",X"23",X"56",X"23",X"EB",X"CD",X"68",X"2F",X"EB",X"4E",X"CB",X"B9",X"CD",
		X"EE",X"2F",X"47",X"3A",X"EC",X"43",X"B7",X"20",X"03",X"13",X"18",X"01",X"1B",X"23",X"7E",X"B7",
		X"78",X"C2",X"4C",X"2F",X"23",X"E9",X"06",X"90",X"3A",X"EC",X"43",X"B7",X"3E",X"07",X"20",X"15",
		X"A5",X"B0",X"D3",X"4B",X"CB",X"3C",X"CB",X"1D",X"CB",X"3C",X"CB",X"1D",X"CB",X"3C",X"CB",X"1D",
		X"01",X"00",X"64",X"09",X"C9",X"A5",X"B0",X"CB",X"DF",X"D3",X"4B",X"CB",X"3C",X"CB",X"1D",X"CB",
		X"3C",X"CB",X"1D",X"CB",X"3C",X"CB",X"1D",X"44",X"4D",X"21",X"FF",X"7F",X"B7",X"ED",X"42",X"C9",
		X"C5",X"06",X"00",X"EB",X"CD",X"68",X"2F",X"EB",X"08",X"C1",X"CB",X"81",X"78",X"3D",X"20",X"02",
		X"CB",X"C1",X"7E",X"CB",X"40",X"20",X"09",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"2B",
		X"23",X"E6",X"0F",X"20",X"08",X"CB",X"41",X"20",X"06",X"3E",X"20",X"18",X"0A",X"CB",X"C1",X"C6",
		X"30",X"FE",X"3A",X"38",X"02",X"C6",X"07",X"E5",X"C5",X"4F",X"08",X"CD",X"EE",X"2F",X"08",X"C1",
		X"E1",X"3A",X"EC",X"43",X"B7",X"20",X"03",X"13",X"18",X"01",X"1B",X"10",X"BF",X"C9",X"D5",X"E5",
		X"32",X"5C",X"F9",X"06",X"09",X"C5",X"CD",X"46",X"C7",X"01",X"C8",X"35",X"C5",X"CD",X"32",X"C7",
		X"E1",X"7E",X"B7",X"F2",X"20",X"30",X"06",X"03",X"0E",X"20",X"C5",X"CD",X"46",X"C7",X"C1",X"D5",
		X"C5",X"3A",X"EC",X"43",X"B7",X"28",X"05",X"CD",X"3B",X"C7",X"18",X"03",X"CD",X"32",X"C7",X"D1",
		X"EB",X"3E",X"09",X"F5",X"F3",X"3A",X"5C",X"F9",X"D3",X"4B",X"3A",X"EC",X"43",X"B7",X"28",X"13",
		X"1A",X"E6",X"7F",X"13",X"77",X"2B",X"36",X"00",X"E5",X"01",X"E1",X"FF",X"C5",X"CD",X"32",X"C7",
		X"E1",X"18",X"11",X"1A",X"E6",X"7F",X"13",X"77",X"23",X"36",X"00",X"E5",X"01",X"1F",X"00",X"C5",
		X"CD",X"32",X"C7",X"E1",X"FB",X"F1",X"3D",X"28",X"03",X"F5",X"18",X"C8",X"E1",X"D1",X"3A",X"5C",
		X"F9",X"C9",X"E5",X"32",X"5C",X"F9",X"79",X"FE",X"20",X"20",X"02",X"0E",X"0A",X"06",X"06",X"C5",
		X"CD",X"46",X"C7",X"01",X"FC",X"30",X"C5",X"CD",X"32",X"C7",X"E1",X"EB",X"06",X"06",X"C5",X"F3",
		X"3A",X"5C",X"F9",X"D3",X"4B",X"3A",X"EC",X"43",X"B7",X"28",X"11",X"1A",X"13",X"77",X"2B",X"36",
		X"00",X"E5",X"01",X"E1",X"FF",X"C5",X"CD",X"32",X"C7",X"E1",X"18",X"0F",X"1A",X"13",X"77",X"23",
		X"36",X"00",X"E5",X"01",X"1F",X"00",X"C5",X"CD",X"32",X"C7",X"E1",X"FB",X"C1",X"05",X"28",X"03",
		X"C5",X"18",X"CC",X"E1",X"C9",X"3E",X"01",X"F5",X"78",X"FE",X"00",X"20",X"02",X"F1",X"C9",X"7E",
		X"CB",X"40",X"20",X"0A",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"18",X"03",X"E6",X"0F",
		X"23",X"4F",X"F1",X"F5",X"B7",X"28",X"10",X"79",X"B7",X"28",X"05",X"F1",X"AF",X"F5",X"18",X"07",
		X"78",X"FE",X"01",X"28",X"02",X"0E",X"20",X"C5",X"D5",X"EB",X"C5",X"CD",X"66",X"2F",X"C1",X"EB",
		X"CD",X"62",X"30",X"D1",X"3E",X"05",X"83",X"5F",X"C1",X"05",X"18",X"BC",X"06",X"09",X"09",X"09",
		X"09",X"06",X"02",X"06",X"02",X"02",X"02",X"07",X"06",X"09",X"01",X"02",X"04",X"0F",X"0F",X"01",
		X"02",X"01",X"09",X"06",X"09",X"09",X"0F",X"01",X"01",X"01",X"0F",X"08",X"0E",X"01",X"01",X"0E",
		X"07",X"08",X"0E",X"09",X"09",X"06",X"0F",X"01",X"01",X"02",X"02",X"02",X"06",X"09",X"06",X"09",
		X"09",X"06",X"06",X"09",X"07",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"21",X"CD",
		X"B6",X"2E",X"E5",X"23",X"23",X"EB",X"21",X"DA",X"F8",X"0E",X"03",X"06",X"0C",X"1A",X"E6",X"0F",
		X"28",X"06",X"CD",X"A1",X"32",X"3D",X"20",X"FA",X"05",X"1A",X"E6",X"F0",X"28",X"07",X"CD",X"A1",
		X"32",X"D6",X"10",X"20",X"F9",X"05",X"1B",X"0D",X"20",X"E3",X"0E",X"0A",X"11",X"73",X"43",X"E1",
		X"E5",X"D5",X"06",X"03",X"1A",X"BE",X"38",X"11",X"20",X"04",X"13",X"23",X"10",X"F6",X"D1",X"21",
		X"06",X"00",X"19",X"EB",X"E1",X"0D",X"20",X"E8",X"C9",X"D1",X"D5",X"06",X"00",X"0D",X"28",X"14",
		X"21",X"00",X"00",X"09",X"29",X"09",X"29",X"E5",X"19",X"2B",X"54",X"5D",X"01",X"06",X"00",X"09",
		X"EB",X"C1",X"ED",X"B8",X"D1",X"E1",X"06",X"03",X"7E",X"23",X"12",X"13",X"10",X"FA",X"EB",X"E5",
		X"CD",X"65",X"1E",X"CD",X"BD",X"CB",X"CD",X"05",X"1F",X"BC",X"32",X"F9",X"32",X"DB",X"32",X"18",
		X"33",X"08",X"06",X"01",X"21",X"B5",X"43",X"CD",X"AA",X"2F",X"CD",X"05",X"1F",X"37",X"33",X"FF",
		X"33",X"9B",X"33",X"79",X"34",X"CD",X"40",X"2F",X"90",X"78",X"62",X"5F",X"5F",X"5F",X"00",X"CD",
		X"05",X"1F",X"55",X"35",X"EC",X"34",X"9B",X"35",X"06",X"36",X"06",X"00",X"21",X"78",X"60",X"CD",
		X"68",X"2F",X"EB",X"E1",X"E5",X"06",X"03",X"36",X"20",X"23",X"10",X"FB",X"E1",X"3E",X"FF",X"32",
		X"B6",X"43",X"06",X"03",X"0E",X"51",X"C5",X"DB",X"48",X"CD",X"2A",X"C7",X"28",X"02",X"DB",X"4A",
		X"2F",X"CB",X"7F",X"20",X"F2",X"AF",X"CD",X"2A",X"C7",X"28",X"02",X"3E",X"08",X"CD",X"EE",X"2F",
		X"D5",X"E5",X"3E",X"06",X"CD",X"40",X"28",X"E1",X"D1",X"C1",X"3A",X"B6",X"43",X"3D",X"32",X"B6",
		X"43",X"28",X"42",X"DB",X"48",X"CD",X"2A",X"C7",X"28",X"02",X"DB",X"4A",X"2F",X"CB",X"7F",X"28",
		X"49",X"3E",X"FA",X"32",X"B6",X"43",X"71",X"C5",X"3A",X"EC",X"43",X"B7",X"01",X"40",X"00",X"28",
		X"03",X"01",X"C0",X"FF",X"D5",X"EB",X"09",X"EB",X"AF",X"CD",X"2A",X"C7",X"28",X"02",X"3E",X"08",
		X"F6",X"90",X"0E",X"5F",X"CD",X"EE",X"2F",X"D1",X"C1",X"23",X"3A",X"EC",X"43",X"B7",X"13",X"28",
		X"02",X"1B",X"1B",X"10",X"91",X"21",X"73",X"43",X"11",X"F2",X"F8",X"06",X"1E",X"7E",X"23",X"12",
		X"13",X"07",X"07",X"07",X"07",X"12",X"13",X"10",X"F4",X"C9",X"3A",X"EE",X"43",X"CB",X"3F",X"CB",
		X"3F",X"CB",X"3F",X"E6",X"1F",X"C6",X"41",X"FE",X"5B",X"38",X"02",X"3E",X"20",X"4F",X"C3",X"06",
		X"32",X"F5",X"C5",X"D5",X"E5",X"16",X"00",X"58",X"1D",X"19",X"0E",X"10",X"7E",X"E6",X"F0",X"81",
		X"27",X"77",X"30",X"03",X"2B",X"10",X"F5",X"E1",X"D1",X"C1",X"F1",X"C9",X"CD",X"40",X"2F",X"90",
		X"28",X"08",X"43",X"6F",X"6E",X"67",X"72",X"61",X"74",X"75",X"6C",X"61",X"74",X"69",X"6F",X"6E",
		X"73",X"20",X"50",X"6C",X"61",X"79",X"65",X"72",X"20",X"00",X"C9",X"CD",X"40",X"2F",X"90",X"20",
		X"08",X"46",X"65",X"6C",X"69",X"63",X"69",X"74",X"61",X"74",X"69",X"6F",X"6E",X"73",X"2C",X"20",
		X"6A",X"6F",X"75",X"65",X"75",X"72",X"20",X"00",X"C9",X"CD",X"40",X"2F",X"90",X"20",X"08",X"47",
		X"6C",X"25",X"65",X"63",X"6B",X"77",X"25",X"65",X"6E",X"73",X"63",X"68",X"65",X"20",X"53",X"70",
		X"69",X"65",X"6C",X"65",X"72",X"20",X"00",X"C9",X"CD",X"40",X"2F",X"90",X"20",X"08",X"46",X"65",
		X"6C",X"69",X"63",X"69",X"74",X"61",X"63",X"69",X"6F",X"6E",X"65",X"73",X"20",X"6A",X"75",X"67",
		X"61",X"64",X"6F",X"72",X"20",X"00",X"C9",X"CD",X"40",X"2F",X"90",X"08",X"20",X"59",X"6F",X"75",
		X"20",X"68",X"61",X"76",X"65",X"20",X"6A",X"6F",X"69",X"6E",X"65",X"64",X"20",X"74",X"68",X"65",
		X"20",X"61",X"73",X"74",X"72",X"6F",X"6E",X"61",X"75",X"74",X"73",X"00",X"CD",X"40",X"2F",X"90",
		X"0C",X"30",X"69",X"6E",X"20",X"74",X"68",X"65",X"20",X"4D",X"4F",X"4F",X"4E",X"20",X"57",X"41",
		X"52",X"20",X"68",X"61",X"6C",X"6C",X"20",X"6F",X"66",X"20",X"66",X"61",X"6D",X"65",X"00",X"CD",
		X"40",X"2F",X"90",X"18",X"50",X"45",X"6E",X"74",X"65",X"72",X"20",X"79",X"6F",X"75",X"72",X"20",
		X"69",X"6E",X"69",X"74",X"69",X"61",X"6C",X"73",X"3A",X"00",X"C9",X"CD",X"40",X"2F",X"90",X"08",
		X"20",X"56",X"6F",X"75",X"73",X"20",X"65",X"74",X"65",X"73",X"20",X"61",X"75",X"20",X"74",X"61",
		X"62",X"6C",X"65",X"61",X"75",X"20",X"64",X"27",X"68",X"6F",X"6E",X"6E",X"65",X"75",X"72",X"00",
		X"CD",X"40",X"2F",X"90",X"0C",X"30",X"64",X"65",X"73",X"20",X"61",X"73",X"74",X"72",X"6F",X"6E",
		X"61",X"75",X"74",X"65",X"73",X"20",X"64",X"75",X"20",X"4D",X"4F",X"4F",X"4E",X"20",X"57",X"41",
		X"52",X"2E",X"00",X"CD",X"40",X"2F",X"90",X"18",X"50",X"54",X"61",X"70",X"65",X"72",X"20",X"76",
		X"6F",X"73",X"20",X"69",X"6E",X"69",X"74",X"69",X"61",X"6C",X"65",X"73",X"3A",X"00",X"C9",X"CD",
		X"40",X"2F",X"90",X"20",X"20",X"53",X"69",X"65",X"20",X"68",X"61",X"62",X"65",X"6E",X"20",X"64",
		X"69",X"65",X"20",X"68",X"24",X"65",X"63",X"68",X"73",X"74",X"65",X"00",X"CD",X"40",X"2F",X"90",
		X"14",X"30",X"61",X"73",X"74",X"72",X"6F",X"6E",X"61",X"75",X"74",X"69",X"73",X"63",X"68",X"65",
		X"20",X"61",X"75",X"73",X"7A",X"65",X"69",X"63",X"68",X"6E",X"75",X"6E",X"67",X"00",X"CD",X"40",
		X"2F",X"90",X"30",X"40",X"69",X"6D",X"20",X"4D",X"4F",X"4F",X"4E",X"20",X"57",X"41",X"52",X"20",
		X"65",X"72",X"6C",X"61",X"6E",X"67",X"74",X"2E",X"00",X"CD",X"40",X"2F",X"90",X"18",X"52",X"49",
		X"68",X"72",X"65",X"20",X"69",X"6E",X"69",X"74",X"69",X"61",X"6C",X"65",X"6E",X"20",X"65",X"69",
		X"6E",X"67",X"65",X"62",X"65",X"6E",X"3A",X"00",X"C9",X"CD",X"40",X"2F",X"90",X"04",X"20",X"55",
		X"73",X"74",X"65",X"64",X"20",X"68",X"61",X"20",X"69",X"6E",X"67",X"72",X"65",X"73",X"61",X"64",
		X"6F",X"20",X"65",X"6E",X"20",X"6C",X"61",X"20",X"73",X"61",X"6C",X"61",X"00",X"CD",X"40",X"2F",
		X"90",X"10",X"30",X"64",X"65",X"20",X"6C",X"61",X"20",X"66",X"61",X"6D",X"61",X"20",X"64",X"65",
		X"20",X"61",X"73",X"74",X"72",X"6F",X"6E",X"61",X"75",X"74",X"61",X"73",X"00",X"CD",X"40",X"2F",
		X"90",X"40",X"40",X"64",X"65",X"20",X"4D",X"4F",X"4F",X"4E",X"20",X"57",X"41",X"52",X"2E",X"00",
		X"CD",X"40",X"2F",X"90",X"18",X"52",X"45",X"6E",X"74",X"72",X"65",X"20",X"73",X"75",X"73",X"20",
		X"69",X"6E",X"69",X"63",X"69",X"61",X"6C",X"65",X"73",X"3A",X"00",X"C9",X"CD",X"40",X"2F",X"90",
		X"08",X"80",X"5A",X"75",X"72",X"20",X"23",X"6E",X"64",X"65",X"72",X"75",X"6E",X"67",X"20",X"64",
		X"65",X"73",X"20",X"62",X"75",X"73",X"63",X"68",X"73",X"74",X"61",X"62",X"65",X"6E",X"73",X"00",
		X"CD",X"40",X"2F",X"90",X"08",X"90",X"72",X"61",X"64",X"20",X"64",X"72",X"65",X"68",X"65",X"6E",
		X"2C",X"20",X"64",X"61",X"6E",X"6E",X"20",X"61",X"75",X"66",X"20",X"46",X"49",X"52",X"45",X"00",
		X"CD",X"40",X"2F",X"90",X"08",X"A0",X"64",X"72",X"25",X"65",X"63",X"6B",X"65",X"6E",X"2C",X"20",
		X"75",X"6D",X"20",X"69",X"68",X"6E",X"20",X"7A",X"75",X"20",X"73",X"70",X"65",X"69",X"63",X"68",
		X"65",X"72",X"6E",X"00",X"C9",X"CD",X"40",X"2F",X"90",X"08",X"80",X"4D",X"6F",X"76",X"65",X"20",
		X"77",X"68",X"65",X"65",X"6C",X"20",X"74",X"6F",X"20",X"63",X"68",X"61",X"6E",X"67",X"65",X"20",
		X"6C",X"65",X"74",X"74",X"65",X"72",X"00",X"CD",X"40",X"2F",X"90",X"08",X"90",X"74",X"68",X"65",
		X"6E",X"20",X"70",X"72",X"65",X"73",X"73",X"20",X"46",X"49",X"52",X"45",X"20",X"74",X"6F",X"20",
		X"73",X"74",X"6F",X"72",X"65",X"20",X"69",X"74",X"2E",X"00",X"C9",X"CD",X"40",X"2F",X"90",X"04",
		X"80",X"54",X"6F",X"75",X"72",X"6E",X"65",X"72",X"20",X"6C",X"61",X"20",X"72",X"6F",X"75",X"65",
		X"20",X"70",X"6F",X"75",X"72",X"20",X"63",X"68",X"61",X"6E",X"67",X"65",X"72",X"00",X"CD",X"40",
		X"2F",X"90",X"04",X"90",X"6C",X"61",X"20",X"6C",X"65",X"74",X"74",X"72",X"65",X"2C",X"20",X"70",
		X"75",X"69",X"73",X"20",X"61",X"70",X"70",X"75",X"79",X"65",X"72",X"20",X"73",X"75",X"72",X"00",
		X"CD",X"40",X"2F",X"90",X"04",X"A0",X"46",X"49",X"52",X"45",X"20",X"70",X"6F",X"75",X"72",X"20",
		X"6C",X"65",X"20",X"6D",X"65",X"74",X"74",X"72",X"65",X"20",X"65",X"6E",X"20",X"6D",X"65",X"6D",
		X"6F",X"69",X"72",X"65",X"00",X"C9",X"CD",X"40",X"2F",X"90",X"04",X"80",X"50",X"61",X"72",X"61",
		X"20",X"63",X"61",X"6D",X"62",X"69",X"61",X"72",X"20",X"6C",X"65",X"20",X"6C",X"65",X"74",X"72",
		X"61",X"2C",X"20",X"67",X"69",X"72",X"65",X"00",X"CD",X"40",X"2F",X"90",X"04",X"90",X"6C",X"61",
		X"20",X"72",X"75",X"65",X"64",X"61",X"2C",X"20",X"6C",X"75",X"65",X"67",X"6F",X"20",X"6F",X"70",
		X"72",X"69",X"6D",X"61",X"20",X"46",X"49",X"52",X"45",X"00",X"CD",X"40",X"2F",X"90",X"04",X"A0",
		X"70",X"61",X"72",X"61",X"20",X"61",X"6C",X"6D",X"61",X"63",X"65",X"6E",X"61",X"72",X"6C",X"61",
		X"2E",X"00",X"C9",X"CD",X"65",X"1E",X"CD",X"BD",X"CB",X"CD",X"92",X"C8",X"3A",X"E9",X"43",X"3D",
		X"06",X"08",X"28",X"02",X"06",X"0E",X"C5",X"78",X"FE",X"0E",X"CC",X"EB",X"3E",X"CD",X"05",X"1F",
		X"A2",X"36",X"B1",X"36",X"C1",X"36",X"CF",X"36",X"08",X"06",X"01",X"21",X"B5",X"43",X"CD",X"AA",
		X"2F",X"C1",X"CB",X"40",X"3E",X"0F",X"28",X"02",X"3E",X"05",X"C5",X"CD",X"40",X"28",X"C1",X"10",
		X"D5",X"C9",X"CD",X"40",X"2F",X"90",X"60",X"50",X"50",X"6C",X"61",X"79",X"65",X"72",X"20",X"00",
		X"C9",X"CD",X"40",X"2F",X"90",X"60",X"50",X"53",X"70",X"69",X"65",X"6C",X"65",X"72",X"20",X"00",
		X"C9",X"CD",X"40",X"2F",X"90",X"60",X"50",X"4A",X"6F",X"75",X"65",X"72",X"20",X"00",X"C9",X"CD",
		X"40",X"2F",X"90",X"60",X"50",X"4A",X"75",X"67",X"61",X"64",X"6F",X"72",X"20",X"00",X"C9",X"00",
		X"3E",X"41",X"5D",X"51",X"5D",X"41",X"3E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"00",X"10",X"14",X"14",X"14",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"14",X"00",X"3A",X"46",X"42",X"42",X"46",X"3A",X"00",X"14",X"00",X"3C",
		X"42",X"42",X"42",X"42",X"3C",X"00",X"14",X"00",X"42",X"42",X"42",X"42",X"42",X"3C",X"00",X"18",
		X"24",X"28",X"10",X"29",X"46",X"46",X"39",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"08",X"10",X"10",X"10",X"10",X"10",X"08",X"04",X"10",X"08",X"04",X"04",X"04",X"04",X"04",
		X"08",X"10",X"00",X"00",X"08",X"2A",X"1C",X"1C",X"2A",X"08",X"00",X"00",X"00",X"08",X"08",X"3E",
		X"08",X"08",X"00",X"00",X"80",X"00",X"00",X"00",X"18",X"18",X"08",X"10",X"00",X"00",X"00",X"00",
		X"00",X"3E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"18",X"00",
		X"00",X"01",X"02",X"04",X"08",X"10",X"20",X"40",X"1C",X"22",X"41",X"41",X"41",X"41",X"41",X"22",
		X"1C",X"08",X"18",X"08",X"08",X"08",X"08",X"08",X"08",X"1C",X"3E",X"41",X"01",X"01",X"3E",X"40",
		X"40",X"40",X"7F",X"3E",X"41",X"01",X"01",X"1E",X"01",X"01",X"41",X"3E",X"02",X"06",X"0A",X"12",
		X"22",X"7F",X"02",X"02",X"02",X"7F",X"40",X"40",X"40",X"7E",X"01",X"01",X"41",X"3E",X"3E",X"41",
		X"40",X"40",X"7E",X"41",X"41",X"41",X"3E",X"7F",X"01",X"02",X"02",X"04",X"04",X"08",X"08",X"08",
		X"3E",X"41",X"41",X"41",X"3E",X"41",X"41",X"41",X"3E",X"3E",X"41",X"41",X"41",X"3F",X"01",X"01",
		X"41",X"3E",X"00",X"00",X"00",X"18",X"18",X"00",X"00",X"18",X"18",X"98",X"18",X"00",X"00",X"18",
		X"18",X"08",X"10",X"00",X"02",X"04",X"08",X"10",X"20",X"10",X"08",X"04",X"02",X"00",X"00",X"00",
		X"3E",X"00",X"3E",X"00",X"00",X"00",X"20",X"10",X"08",X"04",X"02",X"04",X"08",X"10",X"20",X"1C",
		X"22",X"02",X"02",X"04",X"08",X"08",X"00",X"08",X"3E",X"41",X"4F",X"49",X"49",X"4F",X"40",X"40",
		X"3F",X"3E",X"41",X"41",X"41",X"7F",X"41",X"41",X"41",X"41",X"7E",X"41",X"41",X"41",X"7E",X"41",
		X"41",X"41",X"7E",X"3E",X"41",X"40",X"40",X"40",X"40",X"40",X"41",X"3E",X"7E",X"41",X"41",X"41",
		X"41",X"41",X"41",X"41",X"7E",X"7F",X"40",X"40",X"40",X"7C",X"40",X"40",X"40",X"7F",X"7F",X"40",
		X"40",X"40",X"7C",X"40",X"40",X"40",X"40",X"3E",X"41",X"40",X"40",X"47",X"41",X"41",X"41",X"3F",
		X"41",X"41",X"41",X"41",X"7F",X"41",X"41",X"41",X"41",X"1C",X"08",X"08",X"08",X"08",X"08",X"08",
		X"08",X"1C",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"41",X"3E",X"41",X"42",X"44",X"48",X"50",
		X"68",X"44",X"42",X"41",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"7F",X"41",X"63",X"55",
		X"49",X"41",X"41",X"41",X"41",X"41",X"41",X"61",X"51",X"49",X"45",X"43",X"41",X"41",X"41",X"3E",
		X"41",X"41",X"41",X"41",X"41",X"41",X"41",X"3E",X"7E",X"41",X"41",X"41",X"7E",X"40",X"40",X"40",
		X"40",X"3E",X"41",X"41",X"41",X"41",X"41",X"45",X"42",X"3D",X"7E",X"41",X"41",X"41",X"7E",X"48",
		X"44",X"42",X"41",X"3E",X"41",X"40",X"40",X"3E",X"01",X"01",X"41",X"3E",X"7F",X"08",X"08",X"08",
		X"08",X"08",X"08",X"08",X"08",X"41",X"41",X"41",X"41",X"41",X"41",X"41",X"41",X"3E",X"41",X"41",
		X"41",X"22",X"22",X"14",X"14",X"08",X"08",X"41",X"41",X"41",X"41",X"41",X"49",X"55",X"63",X"41",
		X"41",X"41",X"22",X"14",X"08",X"14",X"22",X"41",X"41",X"41",X"41",X"22",X"14",X"08",X"08",X"08",
		X"08",X"08",X"7F",X"01",X"02",X"04",X"08",X"10",X"20",X"40",X"7F",X"3C",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"3C",X"00",X"00",X"40",X"20",X"10",X"08",X"04",X"02",X"01",X"3C",X"04",X"04",
		X"04",X"04",X"04",X"04",X"04",X"3C",X"08",X"14",X"22",X"41",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"18",X"18",X"10",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"3A",X"46",X"42",X"42",X"46",X"3A",X"40",X"40",X"40",X"5C",X"62",X"42",
		X"42",X"62",X"5C",X"00",X"00",X"00",X"3C",X"42",X"40",X"40",X"42",X"3C",X"02",X"02",X"02",X"3A",
		X"46",X"42",X"42",X"46",X"3A",X"00",X"00",X"00",X"3C",X"42",X"7E",X"40",X"40",X"3C",X"0C",X"12",
		X"10",X"10",X"38",X"10",X"10",X"10",X"10",X"BA",X"46",X"42",X"42",X"46",X"3A",X"02",X"42",X"3C",
		X"40",X"40",X"40",X"7C",X"42",X"42",X"42",X"42",X"42",X"00",X"08",X"00",X"08",X"08",X"08",X"08",
		X"08",X"08",X"84",X"04",X"04",X"04",X"04",X"04",X"04",X"44",X"38",X"40",X"40",X"40",X"44",X"48",
		X"50",X"70",X"48",X"44",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"00",X"00",X"00",
		X"76",X"49",X"49",X"49",X"49",X"49",X"00",X"00",X"00",X"7C",X"42",X"42",X"42",X"42",X"42",X"00",
		X"00",X"00",X"3C",X"42",X"42",X"42",X"42",X"3C",X"DC",X"62",X"42",X"42",X"62",X"5C",X"40",X"40",
		X"40",X"BA",X"46",X"42",X"42",X"46",X"3A",X"02",X"02",X"02",X"00",X"00",X"00",X"5C",X"62",X"40",
		X"40",X"40",X"40",X"00",X"00",X"00",X"3C",X"42",X"30",X"0C",X"42",X"3C",X"00",X"10",X"10",X"7C",
		X"10",X"10",X"10",X"10",X"10",X"00",X"00",X"00",X"42",X"42",X"42",X"42",X"42",X"3C",X"00",X"00",
		X"00",X"44",X"44",X"44",X"44",X"28",X"10",X"00",X"00",X"00",X"41",X"41",X"41",X"49",X"49",X"36",
		X"00",X"00",X"00",X"42",X"24",X"18",X"18",X"24",X"42",X"C2",X"42",X"42",X"42",X"46",X"3A",X"02",
		X"42",X"3C",X"00",X"00",X"00",X"7E",X"04",X"08",X"10",X"20",X"7E",X"0C",X"10",X"10",X"10",X"20",
		X"10",X"10",X"10",X"0C",X"08",X"08",X"08",X"00",X"00",X"08",X"08",X"08",X"00",X"18",X"04",X"04",
		X"04",X"02",X"04",X"04",X"04",X"18",X"30",X"49",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"55",
		X"2A",X"55",X"2A",X"55",X"2A",X"55",X"2A",X"55",X"00",X"00",X"00",X"00",X"24",X"66",X"66",X"66",
		X"00",X"21",X"9F",X"F8",X"F5",X"3E",X"FF",X"BE",X"38",X"09",X"D3",X"4D",X"77",X"21",X"D3",X"3A",
		X"22",X"9B",X"F8",X"F1",X"D3",X"4C",X"C9",X"21",X"9F",X"F8",X"F5",X"3E",X"0E",X"BE",X"38",X"09",
		X"D3",X"4D",X"77",X"21",X"7D",X"3A",X"22",X"9B",X"F8",X"F1",X"D3",X"4C",X"C9",X"0E",X"04",X"97",
		X"F8",X"00",X"05",X"06",X"06",X"0E",X"03",X"8E",X"F8",X"92",X"92",X"92",X"0F",X"03",X"91",X"F8",
		X"32",X"00",X"32",X"00",X"32",X"00",X"06",X"04",X"AB",X"F8",X"06",X"32",X"A9",X"F8",X"01",X"0B",
		X"15",X"00",X"91",X"F8",X"0B",X"17",X"00",X"93",X"F8",X"0B",X"29",X"00",X"95",X"F8",X"03",X"A9",
		X"F8",X"EC",X"07",X"32",X"00",X"91",X"F8",X"03",X"AB",X"F8",X"DF",X"06",X"FA",X"A9",X"F8",X"01",
		X"0B",X"0A",X"00",X"91",X"F8",X"0B",X"0D",X"00",X"93",X"F8",X"0B",X"0F",X"00",X"95",X"F8",X"03",
		X"A9",X"F8",X"EC",X"0E",X"03",X"8E",X"F8",X"00",X"00",X"00",X"0E",X"04",X"98",X"F8",X"00",X"00",
		X"00",X"00",X"00",X"21",X"9F",X"F8",X"F5",X"3E",X"16",X"BE",X"38",X"09",X"D3",X"4D",X"77",X"21",
		X"F9",X"3A",X"22",X"9B",X"F8",X"F1",X"D3",X"4C",X"C9",X"0E",X"04",X"97",X"F8",X"00",X"06",X"07",
		X"06",X"0E",X"03",X"8E",X"F8",X"90",X"90",X"90",X"06",X"10",X"A9",X"F8",X"07",X"AC",X"00",X"91",
		X"F8",X"0F",X"02",X"93",X"F8",X"14",X"00",X"0A",X"00",X"06",X"19",X"AB",X"F8",X"01",X"0A",X"05",
		X"93",X"F8",X"0A",X"1E",X"95",X"F8",X"03",X"AB",X"F8",X"F3",X"0A",X"FC",X"91",X"F8",X"03",X"A9",
		X"F8",X"DF",X"02",X"9F",X"21",X"9F",X"F8",X"F5",X"3E",X"13",X"BE",X"38",X"09",X"D3",X"4D",X"77",
		X"21",X"4A",X"3B",X"22",X"9B",X"F8",X"F1",X"D3",X"4C",X"C9",X"0E",X"03",X"8E",X"F8",X"82",X"80",
		X"80",X"0E",X"04",X"97",X"F8",X"03",X"05",X"06",X"07",X"0F",X"03",X"91",X"F8",X"01",X"00",X"01",
		X"00",X"05",X"00",X"0E",X"03",X"8E",X"F8",X"92",X"90",X"90",X"06",X"37",X"AB",X"F8",X"06",X"06",
		X"A9",X"F8",X"01",X"03",X"A9",X"F8",X"FB",X"0B",X"01",X"00",X"91",X"F8",X"03",X"AB",X"F8",X"EE",
		X"0E",X"03",X"8E",X"F8",X"00",X"00",X"00",X"0E",X"04",X"97",X"F8",X"00",X"00",X"00",X"00",X"00",
		X"21",X"9F",X"F8",X"F5",X"3E",X"0F",X"BE",X"38",X"09",X"D3",X"4D",X"77",X"21",X"A6",X"3B",X"22",
		X"9B",X"F8",X"F1",X"D3",X"4C",X"C9",X"0E",X"03",X"8E",X"F8",X"92",X"92",X"92",X"0E",X"04",X"97",
		X"F8",X"00",X"06",X"07",X"06",X"0F",X"03",X"91",X"F8",X"00",X"01",X"10",X"02",X"20",X"03",X"06",
		X"28",X"AB",X"F8",X"01",X"0B",X"16",X"00",X"91",X"F8",X"0B",X"1F",X"00",X"93",X"F8",X"0B",X"14",
		X"00",X"95",X"F8",X"03",X"AB",X"F8",X"EC",X"0F",X"03",X"91",X"F8",X"00",X"01",X"10",X"02",X"20",
		X"03",X"06",X"37",X"AB",X"F8",X"01",X"0B",X"2A",X"00",X"91",X"F8",X"0B",X"33",X"00",X"93",X"F8",
		X"0B",X"28",X"00",X"95",X"F8",X"03",X"AB",X"F8",X"EC",X"06",X"23",X"AB",X"F8",X"01",X"0B",X"F5",
		X"FF",X"91",X"F8",X"0B",X"F5",X"FF",X"93",X"F8",X"0B",X"F5",X"FF",X"95",X"F8",X"03",X"AB",X"F8",
		X"EC",X"0E",X"03",X"8E",X"F8",X"00",X"00",X"00",X"0E",X"04",X"97",X"F8",X"00",X"00",X"00",X"00",
		X"00",X"21",X"9F",X"F8",X"F5",X"3E",X"12",X"BE",X"38",X"09",X"D3",X"4D",X"77",X"21",X"37",X"3C",
		X"22",X"9B",X"F8",X"F1",X"D3",X"4C",X"C9",X"0F",X"03",X"91",X"F8",X"14",X"00",X"2D",X"00",X"5A",
		X"00",X"0E",X"03",X"8E",X"F8",X"92",X"92",X"92",X"0E",X"04",X"97",X"F8",X"00",X"06",X"05",X"07",
		X"06",X"04",X"AB",X"F8",X"06",X"50",X"A9",X"F8",X"01",X"0B",X"08",X"00",X"91",X"F8",X"0B",X"11",
		X"00",X"93",X"F8",X"0B",X"2F",X"00",X"95",X"F8",X"03",X"A9",X"F8",X"EC",X"03",X"AB",X"F8",X"E4",
		X"0E",X"03",X"8E",X"F8",X"00",X"00",X"00",X"0E",X"04",X"97",X"F8",X"00",X"00",X"00",X"00",X"00",
		X"21",X"9F",X"F8",X"F5",X"3E",X"11",X"BE",X"38",X"09",X"D3",X"4D",X"77",X"21",X"F6",X"3C",X"22",
		X"9B",X"F8",X"F1",X"D3",X"4C",X"C9",X"06",X"06",X"AB",X"F8",X"0F",X"03",X"91",X"F8",X"2C",X"01",
		X"C8",X"00",X"64",X"00",X"0E",X"04",X"97",X"F8",X"00",X"07",X"06",X"05",X"02",X"5E",X"06",X"08",
		X"AB",X"F8",X"0F",X"03",X"91",X"F8",X"58",X"02",X"90",X"01",X"C8",X"00",X"0E",X"04",X"97",X"F8",
		X"00",X"06",X"06",X"05",X"02",X"46",X"06",X"0A",X"AB",X"F8",X"0F",X"03",X"91",X"F8",X"84",X"03",
		X"58",X"02",X"2C",X"01",X"0E",X"04",X"97",X"F8",X"00",X"06",X"05",X"04",X"02",X"2E",X"06",X"0C",
		X"AB",X"F8",X"0F",X"03",X"91",X"F8",X"E2",X"04",X"20",X"03",X"90",X"01",X"0E",X"04",X"97",X"F8",
		X"00",X"05",X"05",X"04",X"02",X"16",X"06",X"04",X"AB",X"F8",X"0F",X"03",X"91",X"F8",X"96",X"00",
		X"64",X"00",X"32",X"00",X"0E",X"04",X"97",X"F8",X"00",X"07",X"07",X"07",X"04",X"AB",X"F8",X"A7",
		X"F8",X"0A",X"01",X"9F",X"F8",X"0E",X"03",X"8E",X"F8",X"92",X"92",X"92",X"04",X"A7",X"F8",X"A9",
		X"F8",X"01",X"0B",X"0C",X"00",X"91",X"F8",X"0B",X"08",X"00",X"93",X"F8",X"0B",X"04",X"00",X"95",
		X"F8",X"03",X"A9",X"F8",X"EC",X"04",X"A7",X"F8",X"A9",X"F8",X"0A",X"FE",X"A9",X"F8",X"01",X"0B",
		X"F7",X"FF",X"91",X"F8",X"0B",X"FA",X"FF",X"93",X"F8",X"0B",X"FD",X"FF",X"95",X"F8",X"03",X"A9",
		X"F8",X"EC",X"03",X"AB",X"F8",X"C6",X"0E",X"03",X"8E",X"F8",X"00",X"00",X"00",X"0E",X"04",X"97",
		X"F8",X"00",X"00",X"00",X"00",X"00",X"21",X"9F",X"F8",X"F5",X"3E",X"08",X"BE",X"38",X"09",X"D3",
		X"4D",X"77",X"21",X"96",X"3C",X"22",X"9B",X"F8",X"F1",X"D3",X"4C",X"C9",X"21",X"9F",X"F8",X"F5",
		X"3E",X"06",X"BE",X"38",X"09",X"D3",X"4D",X"77",X"21",X"AE",X"3C",X"22",X"9B",X"F8",X"F1",X"D3",
		X"4C",X"C9",X"21",X"9F",X"F8",X"F5",X"3E",X"04",X"BE",X"38",X"09",X"D3",X"4D",X"77",X"21",X"C6",
		X"3C",X"22",X"9B",X"F8",X"F1",X"D3",X"4C",X"C9",X"21",X"9F",X"F8",X"F5",X"3E",X"02",X"BE",X"38",
		X"09",X"D3",X"4D",X"77",X"21",X"DE",X"3C",X"22",X"9B",X"F8",X"F1",X"D3",X"4C",X"C9",X"21",X"9F",
		X"F8",X"F5",X"3E",X"14",X"BE",X"38",X"09",X"D3",X"4D",X"77",X"21",X"EA",X"3D",X"22",X"9B",X"F8",
		X"F1",X"D3",X"4C",X"C9",X"21",X"9F",X"F8",X"F5",X"3E",X"15",X"BE",X"38",X"09",X"D3",X"4D",X"77",
		X"21",X"04",X"3E",X"22",X"9B",X"F8",X"F1",X"D3",X"4C",X"C9",X"0E",X"04",X"97",X"F8",X"00",X"06",
		X"06",X"06",X"0E",X"03",X"8E",X"F8",X"92",X"92",X"92",X"0F",X"03",X"91",X"F8",X"E8",X"03",X"4C",
		X"04",X"B0",X"04",X"00",X"0B",X"F6",X"FF",X"91",X"F8",X"0B",X"F5",X"FF",X"93",X"F8",X"0B",X"F4",
		X"FF",X"95",X"F8",X"00",X"21",X"9F",X"F8",X"F5",X"3E",X"34",X"BE",X"38",X"09",X"D3",X"4D",X"77",
		X"21",X"2A",X"3E",X"22",X"9B",X"F8",X"F1",X"D3",X"4C",X"C9",X"0E",X"04",X"97",X"F8",X"00",X"07",
		X"07",X"07",X"0E",X"03",X"8E",X"F8",X"92",X"92",X"92",X"0F",X"03",X"91",X"F8",X"C8",X"00",X"3C",
		X"00",X"28",X"00",X"06",X"14",X"AB",X"F8",X"06",X"14",X"A9",X"F8",X"01",X"0B",X"14",X"00",X"91",
		X"F8",X"0B",X"06",X"00",X"93",X"F8",X"0B",X"04",X"00",X"95",X"F8",X"03",X"A9",X"F8",X"EC",X"06",
		X"14",X"A9",X"F8",X"01",X"0B",X"EC",X"FF",X"91",X"F8",X"0B",X"FA",X"FF",X"93",X"F8",X"0B",X"FC",
		X"FF",X"95",X"F8",X"03",X"A9",X"F8",X"EC",X"03",X"AB",X"F8",X"CC",X"0E",X"03",X"8E",X"F8",X"00",
		X"00",X"00",X"0E",X"04",X"97",X"F8",X"00",X"00",X"00",X"00",X"00",X"21",X"9F",X"F8",X"F5",X"3E",
		X"10",X"BE",X"38",X"09",X"D3",X"4D",X"77",X"21",X"A1",X"3E",X"22",X"9B",X"F8",X"F1",X"D3",X"4C",
		X"C9",X"0E",X"04",X"97",X"F8",X"00",X"07",X"06",X"06",X"0E",X"03",X"8E",X"F8",X"92",X"92",X"92",
		X"06",X"03",X"A9",X"F8",X"06",X"1E",X"AB",X"F8",X"0F",X"03",X"91",X"F8",X"B0",X"04",X"BC",X"04",
		X"C7",X"04",X"0B",X"F4",X"FF",X"91",X"F8",X"0B",X"F5",X"FF",X"93",X"F8",X"0B",X"F6",X"FF",X"95",
		X"F8",X"01",X"01",X"03",X"AB",X"F8",X"EB",X"03",X"A9",X"F8",X"D9",X"0E",X"03",X"8E",X"F8",X"00",
		X"00",X"00",X"0E",X"04",X"97",X"F8",X"00",X"00",X"00",X"00",X"00",X"21",X"9F",X"F8",X"F5",X"3E",
		X"17",X"BE",X"38",X"09",X"D3",X"4D",X"77",X"21",X"01",X"3F",X"22",X"9B",X"F8",X"F1",X"D3",X"4C",
		X"C9",X"0E",X"04",X"97",X"F8",X"00",X"07",X"07",X"07",X"0E",X"03",X"8E",X"F8",X"92",X"92",X"92",
		X"06",X"03",X"A9",X"F8",X"0F",X"03",X"91",X"F8",X"2C",X"01",X"90",X"01",X"C8",X"00",X"06",X"3C",
		X"AB",X"F8",X"01",X"03",X"AB",X"F8",X"FB",X"0F",X"03",X"91",X"F8",X"84",X"03",X"BC",X"02",X"20",
		X"03",X"06",X"28",X"AB",X"F8",X"01",X"03",X"AB",X"F8",X"FB",X"03",X"A9",X"F8",X"D6",X"0E",X"03",
		X"8E",X"F8",X"00",X"00",X"00",X"0E",X"04",X"97",X"F8",X"00",X"00",X"00",X"00",X"00",X"21",X"9F",
		X"F8",X"F5",X"3E",X"13",X"BE",X"38",X"09",X"D3",X"4D",X"77",X"21",X"64",X"3F",X"22",X"9B",X"F8",
		X"F1",X"D3",X"4C",X"C9",X"0E",X"03",X"8E",X"F8",X"82",X"82",X"82",X"0F",X"03",X"91",X"F8",X"80",
		X"02",X"00",X"02",X"00",X"03",X"0E",X"04",X"97",X"F8",X"00",X"07",X"07",X"07",X"06",X"32",X"AB",
		X"F8",X"01",X"0B",X"07",X"00",X"91",X"F8",X"0B",X"0B",X"00",X"93",X"F8",X"0B",X"04",X"00",X"95",
		X"F8",X"01",X"03",X"AB",X"F8",X"EC",X"0E",X"03",X"8E",X"F8",X"00",X"00",X"00",X"0E",X"04",X"97",
		X"F8",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"7B",X"2B",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
