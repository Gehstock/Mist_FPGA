`define BUILD_DATE "190212"
`define BUILD_TIME "175138"
