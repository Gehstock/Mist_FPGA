library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity pickin_program is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of pickin_program is
	type rom is array(0 to  24575) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"C3",X"D0",X"0E",X"3A",X"FE",X"70",X"FE",X"01",X"3E",X"50",X"32",X"F7",X"71",X"C8",X"3A",X"FE",
		X"70",X"FE",X"02",X"3E",X"40",X"32",X"F7",X"71",X"C8",X"3E",X"30",X"32",X"F7",X"71",X"C9",X"C6",
		X"01",X"27",X"32",X"F7",X"71",X"C9",X"00",X"08",X"02",X"11",X"00",X"1A",X"00",X"00",X"00",X"01",
		X"80",X"58",X"04",X"10",X"00",X"10",X"12",X"08",X"F5",X"C5",X"D5",X"E5",X"DD",X"E5",X"FD",X"E5",
		X"D9",X"C5",X"D5",X"E5",X"08",X"F5",X"AF",X"32",X"00",X"A0",X"3A",X"00",X"B8",X"F3",X"3E",X"01",
		X"32",X"A0",X"72",X"CD",X"FB",X"2E",X"CD",X"DF",X"0B",X"CD",X"E7",X"02",X"CD",X"4D",X"08",X"CD",
		X"F1",X"09",X"3A",X"A6",X"72",X"FE",X"00",X"28",X"04",X"3D",X"32",X"A6",X"72",X"3A",X"91",X"72",
		X"FE",X"00",X"28",X"01",X"3C",X"32",X"91",X"72",X"11",X"00",X"98",X"21",X"80",X"75",X"01",X"20",
		X"00",X"ED",X"B0",X"CD",X"B2",X"0D",X"3A",X"76",X"72",X"3C",X"32",X"76",X"72",X"CD",X"27",X"0A",
		X"3A",X"79",X"72",X"3C",X"32",X"79",X"72",X"CD",X"62",X"0A",X"3A",X"7C",X"72",X"3C",X"32",X"7C",
		X"72",X"CD",X"A9",X"0A",X"DD",X"21",X"42",X"70",X"CD",X"1C",X"0A",X"DD",X"21",X"43",X"70",X"CD",
		X"1C",X"0A",X"DD",X"21",X"CA",X"72",X"CD",X"1C",X"0A",X"3A",X"5C",X"70",X"FE",X"01",X"CA",X"3F",
		X"02",X"3A",X"FA",X"71",X"FE",X"01",X"28",X"34",X"3A",X"F6",X"71",X"FE",X"00",X"20",X"11",X"3A",
		X"F7",X"71",X"FE",X"00",X"20",X"0A",X"3A",X"FD",X"71",X"FE",X"00",X"20",X"03",X"C3",X"FC",X"00",
		X"AF",X"3A",X"F6",X"71",X"DE",X"01",X"27",X"32",X"F6",X"71",X"3A",X"F7",X"71",X"DE",X"00",X"27",
		X"32",X"F7",X"71",X"3A",X"FD",X"71",X"DE",X"00",X"27",X"32",X"FD",X"71",X"3A",X"52",X"70",X"FE",
		X"0A",X"28",X"06",X"3C",X"32",X"52",X"70",X"18",X"24",X"AF",X"32",X"52",X"70",X"21",X"E2",X"70",
		X"06",X"09",X"CD",X"80",X"02",X"23",X"10",X"FA",X"21",X"BF",X"72",X"CD",X"80",X"02",X"21",X"C0",
		X"72",X"CD",X"80",X"02",X"21",X"C3",X"72",X"CD",X"80",X"02",X"CD",X"0E",X"0C",X"3A",X"62",X"70",
		X"FE",X"00",X"20",X"45",X"3A",X"63",X"70",X"FE",X"01",X"28",X"22",X"3A",X"A6",X"72",X"FE",X"00",
		X"20",X"37",X"21",X"13",X"70",X"DD",X"21",X"88",X"75",X"FD",X"21",X"80",X"75",X"CD",X"5F",X"03",
		X"DD",X"21",X"98",X"75",X"FD",X"21",X"80",X"75",X"CD",X"5F",X"03",X"18",X"1C",X"21",X"BD",X"72",
		X"DD",X"21",X"88",X"75",X"FD",X"21",X"80",X"75",X"CD",X"5F",X"03",X"21",X"BE",X"72",X"DD",X"21",
		X"98",X"75",X"FD",X"21",X"80",X"75",X"CD",X"5F",X"03",X"3A",X"42",X"70",X"FE",X"00",X"C2",X"29",
		X"02",X"3A",X"5D",X"70",X"FE",X"01",X"CA",X"29",X"02",X"3A",X"13",X"70",X"FE",X"01",X"CA",X"29",
		X"02",X"CD",X"19",X"03",X"3A",X"8D",X"72",X"FE",X"01",X"28",X"58",X"3A",X"0D",X"73",X"2F",X"E6",
		X"01",X"32",X"0D",X"73",X"3A",X"00",X"B8",X"AF",X"32",X"45",X"70",X"11",X"0C",X"00",X"ED",X"53",
		X"4D",X"70",X"DD",X"21",X"88",X"75",X"FD",X"21",X"34",X"70",X"CD",X"B1",X"04",X"3E",X"02",X"32",
		X"45",X"70",X"DD",X"21",X"98",X"75",X"FD",X"21",X"84",X"72",X"CD",X"B1",X"04",X"DD",X"21",X"90",
		X"75",X"FD",X"21",X"34",X"70",X"CD",X"BA",X"03",X"3A",X"D0",X"72",X"FE",X"00",X"28",X"11",X"47",
		X"DD",X"21",X"D1",X"72",X"C5",X"CD",X"6D",X"02",X"C1",X"11",X"09",X"00",X"DD",X"19",X"10",X"F4",
		X"CD",X"64",X"0C",X"CD",X"57",X"0C",X"CD",X"0D",X"0C",X"11",X"18",X"00",X"3A",X"FD",X"70",X"FE",
		X"03",X"20",X"03",X"11",X"3C",X"00",X"ED",X"53",X"4D",X"70",X"DD",X"21",X"80",X"75",X"FD",X"21",
		X"20",X"70",X"3E",X"01",X"32",X"BA",X"72",X"3A",X"62",X"70",X"FE",X"00",X"CC",X"12",X"05",X"AF",
		X"32",X"BA",X"72",X"CD",X"A6",X"03",X"CD",X"32",X"2D",X"DD",X"21",X"80",X"75",X"FD",X"21",X"20",
		X"70",X"CD",X"B7",X"02",X"DD",X"21",X"88",X"75",X"FD",X"21",X"34",X"70",X"CD",X"B7",X"02",X"CD",
		X"3F",X"09",X"3A",X"00",X"B8",X"CD",X"78",X"09",X"3A",X"00",X"B8",X"3E",X"00",X"32",X"A0",X"72",
		X"3A",X"00",X"B8",X"CD",X"D7",X"0D",X"3E",X"01",X"32",X"00",X"A0",X"ED",X"56",X"F1",X"08",X"E1",
		X"D1",X"C1",X"D9",X"FD",X"E1",X"DD",X"E1",X"E1",X"D1",X"C1",X"F1",X"FB",X"C9",X"DD",X"7E",X"05",
		X"FE",X"00",X"28",X"08",X"FE",X"D0",X"38",X"04",X"CD",X"1A",X"20",X"C9",X"DD",X"34",X"05",X"C9",
		X"7E",X"FE",X"00",X"C8",X"FE",X"FF",X"C8",X"3C",X"77",X"C9",X"3E",X"FF",X"CD",X"35",X"27",X"E5",
		X"CD",X"F0",X"26",X"3E",X"07",X"CD",X"35",X"27",X"E1",X"ED",X"5B",X"65",X"70",X"19",X"C5",X"3A",
		X"82",X"75",X"47",X"3A",X"67",X"70",X"80",X"32",X"82",X"75",X"3A",X"83",X"75",X"47",X"3A",X"68",
		X"70",X"80",X"32",X"83",X"75",X"C1",X"C9",X"FD",X"7E",X"00",X"FE",X"00",X"C8",X"DD",X"7E",X"02",
		X"3D",X"DD",X"77",X"06",X"DD",X"7E",X"03",X"DD",X"77",X"07",X"C9",X"3A",X"03",X"70",X"E6",X"80",
		X"FE",X"80",X"C8",X"3A",X"02",X"70",X"E6",X"80",X"FE",X"80",X"C0",X"C9",X"3E",X"3A",X"32",X"80",
		X"75",X"3E",X"01",X"32",X"14",X"70",X"C9",X"3A",X"14",X"70",X"FE",X"00",X"C8",X"3A",X"14",X"70",
		X"3C",X"32",X"14",X"70",X"FE",X"11",X"20",X"0A",X"3E",X"3A",X"32",X"80",X"75",X"AF",X"32",X"14",
		X"70",X"C9",X"FE",X"09",X"38",X"08",X"3A",X"80",X"75",X"3C",X"32",X"80",X"75",X"C9",X"3A",X"80",
		X"75",X"FE",X"33",X"C8",X"3D",X"32",X"80",X"75",X"C9",X"3A",X"BD",X"72",X"FE",X"00",X"C0",X"3A",
		X"BE",X"72",X"FE",X"00",X"C0",X"DD",X"21",X"80",X"75",X"FD",X"21",X"90",X"75",X"CD",X"6C",X"03",
		X"38",X"27",X"CD",X"82",X"03",X"38",X"22",X"3A",X"61",X"70",X"FE",X"01",X"28",X"15",X"3E",X"01",
		X"32",X"62",X"70",X"3A",X"20",X"70",X"FE",X"00",X"28",X"09",X"CD",X"00",X"24",X"2A",X"AD",X"72",
		X"CD",X"C1",X"1E",X"3E",X"01",X"32",X"61",X"70",X"C9",X"3E",X"00",X"32",X"61",X"70",X"C9",X"00",
		X"CD",X"6C",X"03",X"D8",X"CD",X"82",X"03",X"D8",X"3E",X"01",X"77",X"C9",X"DD",X"7E",X"02",X"CD",
		X"98",X"03",X"80",X"FD",X"BE",X"02",X"D8",X"FD",X"7E",X"02",X"CD",X"98",X"03",X"80",X"DD",X"BE",
		X"02",X"C9",X"DD",X"7E",X"03",X"CD",X"98",X"03",X"80",X"FD",X"BE",X"03",X"D8",X"FD",X"7E",X"03",
		X"CD",X"98",X"03",X"80",X"DD",X"BE",X"03",X"C9",X"F5",X"06",X"0B",X"3A",X"20",X"70",X"FE",X"00",
		X"28",X"02",X"06",X"0A",X"F1",X"C9",X"3A",X"62",X"70",X"FE",X"00",X"C8",X"3A",X"92",X"75",X"3C",
		X"32",X"82",X"75",X"3A",X"93",X"75",X"32",X"83",X"75",X"C9",X"DD",X"7E",X"02",X"32",X"C6",X"72",
		X"DD",X"7E",X"03",X"32",X"C7",X"72",X"3A",X"4B",X"70",X"FE",X"01",X"28",X"0D",X"DD",X"7E",X"02",
		X"47",X"3A",X"49",X"70",X"80",X"DD",X"77",X"02",X"18",X"0B",X"3A",X"49",X"70",X"47",X"DD",X"7E",
		X"02",X"90",X"DD",X"77",X"02",X"3A",X"4A",X"70",X"47",X"3A",X"4C",X"70",X"FE",X"01",X"28",X"09",
		X"DD",X"7E",X"03",X"80",X"DD",X"77",X"03",X"18",X"07",X"DD",X"7E",X"03",X"90",X"DD",X"77",X"03",
		X"CD",X"A1",X"17",X"28",X"27",X"CD",X"BD",X"17",X"28",X"22",X"CD",X"69",X"17",X"28",X"1D",X"CD",
		X"85",X"17",X"28",X"18",X"3A",X"94",X"72",X"FE",X"01",X"28",X"0C",X"E5",X"21",X"49",X"70",X"7E",
		X"23",X"86",X"E1",X"FE",X"00",X"28",X"05",X"AF",X"32",X"A7",X"72",X"C9",X"21",X"66",X"0E",X"22",
		X"00",X"73",X"21",X"77",X"0E",X"22",X"02",X"73",X"3A",X"A7",X"72",X"3C",X"32",X"A7",X"72",X"FE",
		X"07",X"20",X"0C",X"3A",X"00",X"B8",X"AF",X"32",X"A7",X"72",X"CD",X"2E",X"0C",X"18",X"26",X"CD",
		X"FB",X"2E",X"E6",X"03",X"47",X"32",X"49",X"70",X"CD",X"FB",X"2E",X"E6",X"03",X"32",X"4A",X"70",
		X"B0",X"FE",X"00",X"28",X"EA",X"CD",X"FB",X"2E",X"E6",X"01",X"32",X"4B",X"70",X"CD",X"FB",X"2E",
		X"E6",X"01",X"32",X"4C",X"70",X"CD",X"A4",X"04",X"3A",X"62",X"70",X"FE",X"00",X"CA",X"BA",X"03",
		X"3A",X"82",X"75",X"E6",X"FC",X"32",X"82",X"75",X"3A",X"83",X"75",X"3C",X"E6",X"FC",X"32",X"83",
		X"75",X"3E",X"00",X"32",X"5B",X"70",X"32",X"62",X"70",X"3E",X"40",X"32",X"A6",X"72",X"CD",X"DB",
		X"02",X"C3",X"BA",X"03",X"3A",X"C6",X"72",X"DD",X"77",X"02",X"3A",X"C7",X"72",X"DD",X"77",X"03",
		X"C9",X"FD",X"7E",X"01",X"E6",X"20",X"FE",X"20",X"CC",X"53",X"05",X"FD",X"7E",X"01",X"E6",X"40",
		X"FE",X"40",X"CC",X"B3",X"05",X"FD",X"7E",X"01",X"E6",X"10",X"FE",X"10",X"CC",X"10",X"06",X"FD",
		X"7E",X"01",X"E6",X"08",X"FE",X"08",X"CC",X"6D",X"06",X"FD",X"7E",X"05",X"3C",X"FD",X"77",X"05",
		X"FE",X"02",X"C0",X"AF",X"FD",X"77",X"05",X"3A",X"45",X"70",X"FE",X"02",X"28",X"04",X"CD",X"02",
		X"05",X"C9",X"3A",X"98",X"75",X"3D",X"32",X"98",X"75",X"FE",X"3B",X"C0",X"3E",X"3F",X"32",X"98",
		X"75",X"C9",X"3A",X"88",X"75",X"3D",X"32",X"88",X"75",X"FE",X"2A",X"C0",X"3E",X"2F",X"32",X"88",
		X"75",X"C9",X"3A",X"02",X"70",X"E6",X"78",X"FE",X"00",X"20",X"04",X"32",X"22",X"70",X"C9",X"3A",
		X"22",X"70",X"FE",X"FF",X"28",X"04",X"3C",X"32",X"22",X"70",X"3A",X"03",X"70",X"E6",X"20",X"FE",
		X"20",X"CC",X"53",X"05",X"3A",X"03",X"70",X"E6",X"40",X"FE",X"40",X"CC",X"B3",X"05",X"3A",X"03",
		X"70",X"E6",X"10",X"FE",X"10",X"CC",X"10",X"06",X"3A",X"03",X"70",X"E6",X"08",X"FE",X"08",X"CC",
		X"6D",X"06",X"C9",X"CD",X"8F",X"05",X"C2",X"5C",X"07",X"CD",X"62",X"07",X"3A",X"BA",X"72",X"FE",
		X"01",X"20",X"13",X"3A",X"B6",X"72",X"CD",X"C5",X"06",X"FE",X"FF",X"28",X"01",X"3C",X"32",X"B6",
		X"72",X"FE",X"05",X"D4",X"08",X"07",X"DD",X"35",X"03",X"3E",X"37",X"CD",X"AA",X"06",X"78",X"3D",
		X"47",X"C8",X"C5",X"CD",X"8F",X"05",X"C1",X"C2",X"5C",X"07",X"DD",X"35",X"03",X"18",X"EF",X"11",
		X"07",X"03",X"CD",X"FE",X"18",X"2B",X"7E",X"CD",X"42",X"07",X"C0",X"11",X"07",X"06",X"CD",X"FE",
		X"18",X"2B",X"7E",X"CD",X"42",X"07",X"C0",X"11",X"07",X"0C",X"CD",X"FE",X"18",X"2B",X"7E",X"CD",
		X"42",X"07",X"C9",X"CD",X"EF",X"05",X"C2",X"5C",X"07",X"CD",X"62",X"07",X"3A",X"BA",X"72",X"FE",
		X"01",X"20",X"13",X"3A",X"B7",X"72",X"CD",X"C5",X"06",X"FE",X"FF",X"28",X"01",X"3C",X"32",X"B7",
		X"72",X"FE",X"05",X"D4",X"08",X"07",X"DD",X"34",X"03",X"3E",X"77",X"CD",X"AA",X"06",X"78",X"3D",
		X"47",X"C8",X"C5",X"CD",X"EF",X"05",X"C1",X"C2",X"5C",X"07",X"DD",X"34",X"03",X"18",X"EF",X"11",
		X"10",X"03",X"CD",X"FE",X"18",X"7E",X"CD",X"42",X"07",X"C0",X"11",X"10",X"06",X"CD",X"FE",X"18",
		X"7E",X"CD",X"42",X"07",X"C0",X"11",X"10",X"0C",X"CD",X"FE",X"18",X"7E",X"CD",X"42",X"07",X"C9",
		X"CD",X"4C",X"06",X"C2",X"5C",X"07",X"CD",X"62",X"07",X"3A",X"BA",X"72",X"FE",X"01",X"20",X"13",
		X"3A",X"B8",X"72",X"CD",X"C5",X"06",X"FE",X"FF",X"28",X"01",X"3C",X"32",X"B8",X"72",X"FE",X"05",
		X"D4",X"20",X"07",X"DD",X"34",X"02",X"3E",X"B9",X"CD",X"AA",X"06",X"78",X"3D",X"47",X"C8",X"C5",
		X"CD",X"4C",X"06",X"C1",X"C2",X"5C",X"07",X"DD",X"34",X"02",X"18",X"EF",X"11",X"03",X"10",X"CD",
		X"FE",X"18",X"7E",X"CD",X"42",X"07",X"C0",X"11",X"06",X"10",X"CD",X"FE",X"18",X"7E",X"CD",X"42",
		X"07",X"C0",X"11",X"0C",X"10",X"CD",X"FE",X"18",X"7E",X"CD",X"42",X"07",X"C9",X"CD",X"D5",X"06",
		X"C2",X"5C",X"07",X"CD",X"62",X"07",X"3A",X"BA",X"72",X"FE",X"01",X"20",X"13",X"3A",X"B9",X"72",
		X"CD",X"C5",X"06",X"FE",X"FF",X"28",X"01",X"3C",X"32",X"B9",X"72",X"FE",X"05",X"D4",X"20",X"07",
		X"DD",X"35",X"02",X"3E",X"39",X"CD",X"AA",X"06",X"78",X"3D",X"47",X"C8",X"C5",X"CD",X"D5",X"06",
		X"C1",X"C2",X"5C",X"07",X"DD",X"35",X"02",X"18",X"EF",X"C9",X"C5",X"47",X"3A",X"20",X"70",X"FE",
		X"00",X"28",X"04",X"78",X"D6",X"15",X"47",X"3A",X"CD",X"72",X"FE",X"06",X"78",X"38",X"01",X"3C",
		X"32",X"80",X"75",X"C1",X"C9",X"F5",X"AF",X"32",X"B6",X"72",X"32",X"B7",X"72",X"32",X"B8",X"72",
		X"32",X"B9",X"72",X"F1",X"C9",X"11",X"03",X"07",X"CD",X"FE",X"18",X"AF",X"11",X"20",X"00",X"ED",
		X"5A",X"7E",X"CD",X"42",X"07",X"C0",X"11",X"06",X"07",X"CD",X"FE",X"18",X"AF",X"11",X"20",X"00",
		X"ED",X"5A",X"7E",X"CD",X"42",X"07",X"C0",X"11",X"0C",X"07",X"CD",X"FE",X"18",X"AF",X"11",X"20",
		X"00",X"ED",X"5A",X"7E",X"CD",X"42",X"07",X"C9",X"3A",X"94",X"72",X"FE",X"01",X"C8",X"DD",X"7E",
		X"02",X"C5",X"CD",X"38",X"07",X"DD",X"7E",X"02",X"E6",X"F8",X"80",X"C1",X"DD",X"77",X"02",X"C9",
		X"3A",X"94",X"72",X"FE",X"01",X"C8",X"DD",X"7E",X"03",X"C5",X"CD",X"38",X"07",X"DD",X"7E",X"03",
		X"E6",X"F8",X"80",X"C1",X"DD",X"77",X"03",X"C9",X"E6",X"07",X"06",X"00",X"FE",X"04",X"D8",X"06",
		X"08",X"C9",X"E5",X"5F",X"FD",X"7E",X"00",X"FE",X"01",X"20",X"05",X"01",X"08",X"00",X"18",X"04",
		X"ED",X"4B",X"4D",X"70",X"21",X"D3",X"07",X"7B",X"ED",X"B1",X"E1",X"C9",X"3E",X"01",X"FD",X"77",
		X"04",X"C9",X"3A",X"94",X"72",X"FE",X"01",X"28",X"3D",X"3A",X"FD",X"70",X"FE",X"03",X"28",X"33",
		X"FD",X"7E",X"02",X"FE",X"07",X"38",X"2F",X"FE",X"08",X"28",X"40",X"FE",X"10",X"38",X"24",X"06",
		X"02",X"3A",X"4D",X"70",X"FE",X"0C",X"C0",X"3A",X"FE",X"70",X"FE",X"01",X"C8",X"E5",X"3A",X"FE",
		X"70",X"21",X"0D",X"73",X"86",X"E1",X"06",X"02",X"FE",X"09",X"D8",X"06",X"04",X"FE",X"11",X"D0",
		X"06",X"03",X"C9",X"06",X"01",X"C9",X"FD",X"7E",X"03",X"FE",X"00",X"28",X"07",X"AF",X"FD",X"77",
		X"03",X"06",X"01",X"C9",X"3E",X"01",X"FD",X"77",X"03",X"F1",X"C9",X"FD",X"7E",X"03",X"FE",X"02",
		X"28",X"0A",X"FD",X"7E",X"03",X"3C",X"FD",X"77",X"03",X"06",X"02",X"C9",X"3E",X"00",X"FD",X"77",
		X"03",X"F1",X"C9",X"40",X"41",X"42",X"43",X"44",X"45",X"FF",X"FE",X"CB",X"CA",X"C9",X"C8",X"A4",
		X"A5",X"A6",X"A7",X"A0",X"A1",X"A2",X"A3",X"9C",X"9D",X"9E",X"9F",X"54",X"55",X"56",X"57",X"58",
		X"59",X"5A",X"5B",X"5C",X"5D",X"5E",X"5F",X"60",X"61",X"62",X"63",X"64",X"65",X"66",X"67",X"68",
		X"69",X"6A",X"6B",X"6C",X"6D",X"6E",X"6F",X"70",X"71",X"72",X"73",X"74",X"75",X"76",X"77",X"00",
		X"C9",X"3A",X"11",X"70",X"FE",X"01",X"28",X"0D",X"FE",X"02",X"28",X"13",X"FE",X"03",X"28",X"19",
		X"FE",X"04",X"28",X"1F",X"C9",X"3A",X"82",X"75",X"3C",X"3C",X"3C",X"32",X"82",X"75",X"C9",X"3A",
		X"82",X"75",X"3D",X"3D",X"3D",X"32",X"82",X"75",X"C9",X"3A",X"83",X"75",X"3D",X"3D",X"3D",X"32",
		X"83",X"75",X"C9",X"3A",X"83",X"75",X"3C",X"3C",X"3C",X"32",X"83",X"75",X"C9",X"CD",X"88",X"08",
		X"CD",X"A5",X"08",X"CD",X"C2",X"08",X"CD",X"DF",X"08",X"3A",X"07",X"70",X"E6",X"08",X"FE",X"08",
		X"C0",X"3A",X"00",X"70",X"FE",X"00",X"C0",X"3A",X"53",X"70",X"FE",X"00",X"C0",X"3A",X"02",X"70",
		X"E6",X"04",X"FE",X"04",X"3E",X"01",X"28",X"0C",X"3A",X"04",X"70",X"E6",X"04",X"FE",X"04",X"3E",
		X"02",X"28",X"01",X"C9",X"32",X"00",X"70",X"C9",X"3A",X"02",X"70",X"E6",X"01",X"47",X"3A",X"03",
		X"70",X"E6",X"01",X"B8",X"C8",X"3A",X"03",X"70",X"E6",X"01",X"FE",X"01",X"C0",X"3E",X"01",X"0E",
		X"01",X"CD",X"FC",X"08",X"C9",X"3A",X"02",X"70",X"E6",X"02",X"47",X"3A",X"03",X"70",X"E6",X"02",
		X"B8",X"C8",X"3A",X"03",X"70",X"E6",X"02",X"FE",X"02",X"C0",X"3E",X"02",X"0E",X"02",X"CD",X"FC",
		X"08",X"C9",X"3A",X"04",X"70",X"E6",X"01",X"47",X"3A",X"05",X"70",X"E6",X"01",X"B8",X"C8",X"3A",
		X"05",X"70",X"E6",X"01",X"FE",X"01",X"C0",X"3E",X"06",X"0E",X"05",X"CD",X"FC",X"08",X"C9",X"3A",
		X"04",X"70",X"E6",X"02",X"47",X"3A",X"05",X"70",X"E6",X"02",X"B8",X"C8",X"3A",X"05",X"70",X"E6",
		X"02",X"FE",X"02",X"C0",X"3E",X"0E",X"0E",X"0A",X"CD",X"FC",X"08",X"C9",X"F5",X"CD",X"71",X"09",
		X"21",X"5F",X"37",X"CD",X"CF",X"0B",X"AF",X"32",X"7C",X"72",X"F1",X"47",X"3A",X"07",X"70",X"E6",
		X"01",X"FE",X"01",X"78",X"28",X"01",X"87",X"21",X"01",X"70",X"86",X"77",X"FE",X"02",X"D4",X"22",
		X"09",X"C9",X"21",X"01",X"70",X"7E",X"FE",X"02",X"D8",X"3A",X"00",X"70",X"FE",X"90",X"C8",X"C6",
		X"01",X"27",X"32",X"00",X"70",X"21",X"01",X"70",X"35",X"35",X"CD",X"3F",X"09",X"18",X"E3",X"3A",
		X"07",X"70",X"E6",X"08",X"FE",X"08",X"20",X"0A",X"21",X"7F",X"89",X"11",X"42",X"58",X"CD",X"49",
		X"19",X"C9",X"3A",X"00",X"70",X"E6",X"0F",X"32",X"7F",X"88",X"3A",X"00",X"70",X"CB",X"0F",X"CB",
		X"0F",X"CB",X"0F",X"CB",X"0F",X"E6",X"0F",X"32",X"9F",X"88",X"C9",X"01",X"01",X"01",X"00",X"01",
		X"00",X"79",X"21",X"08",X"70",X"86",X"77",X"C9",X"3A",X"5E",X"70",X"FE",X"01",X"28",X"06",X"3A",
		X"02",X"70",X"32",X"03",X"70",X"AF",X"32",X"05",X"A0",X"18",X"08",X"3E",X"07",X"D3",X"08",X"3E",
		X"1F",X"D3",X"09",X"3E",X"0E",X"D3",X"08",X"DB",X"0C",X"2F",X"CD",X"CF",X"09",X"47",X"3A",X"53",
		X"70",X"FE",X"00",X"78",X"20",X"09",X"E6",X"07",X"47",X"3A",X"02",X"70",X"E6",X"F8",X"B0",X"32",
		X"02",X"70",X"3A",X"04",X"70",X"32",X"05",X"70",X"3E",X"0F",X"D3",X"08",X"DB",X"0C",X"2F",X"32",
		X"04",X"70",X"3A",X"00",X"A8",X"2F",X"32",X"07",X"70",X"3E",X"01",X"32",X"05",X"A0",X"C9",X"47",
		X"3A",X"00",X"A8",X"2F",X"CB",X"07",X"E6",X"01",X"4F",X"3A",X"0B",X"70",X"A1",X"32",X"0D",X"70",
		X"FE",X"01",X"28",X"02",X"78",X"C9",X"3A",X"04",X"70",X"E6",X"F8",X"4F",X"78",X"E6",X"07",X"B1",
		X"C9",X"21",X"04",X"A0",X"FD",X"21",X"08",X"70",X"FD",X"7E",X"00",X"FE",X"00",X"28",X"16",X"FD",
		X"34",X"01",X"FD",X"7E",X"01",X"FE",X"10",X"38",X"0C",X"FE",X"20",X"38",X"0B",X"FD",X"35",X"00",
		X"AF",X"FD",X"77",X"01",X"C9",X"AF",X"77",X"C9",X"3E",X"01",X"77",X"C9",X"DD",X"7E",X"00",X"FE",
		X"00",X"C8",X"3C",X"DD",X"77",X"00",X"C9",X"2A",X"74",X"72",X"11",X"02",X"00",X"19",X"7E",X"FE",
		X"FF",X"CA",X"EC",X"0A",X"3A",X"7E",X"72",X"47",X"3A",X"76",X"72",X"B8",X"C0",X"AF",X"32",X"76",
		X"72",X"2A",X"74",X"72",X"11",X"05",X"53",X"AF",X"32",X"06",X"A0",X"CD",X"18",X"0B",X"3E",X"0F",
		X"D3",X"08",X"3E",X"01",X"32",X"06",X"A0",X"2A",X"74",X"72",X"11",X"03",X"00",X"19",X"22",X"74",
		X"72",X"C9",X"2A",X"77",X"72",X"11",X"02",X"00",X"19",X"7E",X"FE",X"FF",X"CA",X"EC",X"0A",X"3A",
		X"7E",X"72",X"47",X"3A",X"79",X"72",X"B8",X"C0",X"AF",X"32",X"79",X"72",X"2A",X"7A",X"72",X"11",
		X"02",X"00",X"19",X"7E",X"FE",X"FF",X"20",X"16",X"2A",X"77",X"72",X"11",X"0D",X"53",X"AF",X"32",
		X"05",X"A0",X"CD",X"18",X"0B",X"3E",X"0F",X"D3",X"08",X"3E",X"01",X"32",X"05",X"A0",X"2A",X"77",
		X"72",X"11",X"03",X"00",X"19",X"22",X"77",X"72",X"C9",X"3A",X"F7",X"72",X"FE",X"00",X"28",X"04",
		X"CD",X"9F",X"0C",X"C9",X"2A",X"7A",X"72",X"11",X"02",X"00",X"19",X"7E",X"FE",X"FF",X"C8",X"3E",
		X"02",X"47",X"3A",X"7C",X"72",X"B8",X"C0",X"AF",X"32",X"7C",X"72",X"2A",X"7A",X"72",X"11",X"15",
		X"53",X"AF",X"32",X"05",X"A0",X"CD",X"1E",X"0B",X"3E",X"0F",X"D3",X"08",X"3E",X"01",X"32",X"05",
		X"A0",X"2A",X"7A",X"72",X"11",X"03",X"00",X"19",X"22",X"7A",X"72",X"C9",X"3A",X"7F",X"72",X"FE",
		X"00",X"C8",X"3A",X"A2",X"72",X"FE",X"01",X"C8",X"21",X"29",X"34",X"CD",X"89",X"0B",X"21",X"C0",
		X"30",X"CD",X"A3",X"0B",X"AF",X"32",X"76",X"72",X"32",X"79",X"72",X"3A",X"F7",X"72",X"2F",X"E6",
		X"01",X"32",X"F7",X"72",X"CD",X"F7",X"0D",X"C9",X"3A",X"F7",X"72",X"FE",X"01",X"C8",X"3E",X"06",
		X"D3",X"08",X"3E",X"07",X"D3",X"09",X"3E",X"07",X"D3",X"08",X"3E",X"38",X"D3",X"09",X"0E",X"00",
		X"D5",X"CD",X"3C",X"0B",X"D1",X"EB",X"0E",X"08",X"CD",X"7C",X"0B",X"C9",X"C5",X"E5",X"7E",X"FE",
		X"00",X"20",X"0E",X"23",X"7E",X"FE",X"00",X"20",X"08",X"23",X"7E",X"FE",X"00",X"20",X"02",X"18",
		X"10",X"E1",X"C1",X"06",X"03",X"79",X"D3",X"08",X"7E",X"CD",X"66",X"0B",X"23",X"0C",X"10",X"F5",
		X"C9",X"E1",X"C1",X"F1",X"F1",X"C9",X"E5",X"87",X"26",X"00",X"6F",X"11",X"1D",X"53",X"19",X"7E",
		X"D3",X"09",X"0C",X"79",X"D3",X"08",X"23",X"7E",X"D3",X"09",X"E1",X"C9",X"06",X"06",X"79",X"D3",
		X"08",X"0C",X"7E",X"D3",X"09",X"23",X"10",X"F6",X"C9",X"E5",X"2A",X"74",X"72",X"D5",X"11",X"02",
		X"00",X"19",X"D1",X"7E",X"E1",X"FE",X"FF",X"C0",X"CD",X"D7",X"0B",X"AF",X"32",X"76",X"72",X"22",
		X"74",X"72",X"C9",X"E5",X"2A",X"77",X"72",X"D5",X"11",X"02",X"00",X"19",X"D1",X"7E",X"E1",X"FE",
		X"FF",X"C0",X"CD",X"D7",X"0B",X"AF",X"32",X"79",X"72",X"22",X"77",X"72",X"C9",X"E5",X"2A",X"7A",
		X"72",X"D5",X"11",X"02",X"00",X"19",X"D1",X"7E",X"E1",X"FE",X"FF",X"C0",X"CD",X"D7",X"0B",X"AF",
		X"32",X"7C",X"72",X"22",X"7A",X"72",X"C9",X"3A",X"53",X"70",X"FE",X"01",X"C8",X"F1",X"C9",X"3A",
		X"02",X"70",X"FE",X"A5",X"C0",X"3E",X"04",X"08",X"21",X"AB",X"8B",X"11",X"B8",X"52",X"CD",X"6B",
		X"23",X"21",X"AC",X"8B",X"11",X"CD",X"52",X"CD",X"6B",X"23",X"21",X"AD",X"8B",X"11",X"E3",X"52",
		X"CD",X"6B",X"23",X"21",X"AE",X"8B",X"11",X"F6",X"52",X"CD",X"6B",X"23",X"C9",X"C9",X"3A",X"63",
		X"70",X"FE",X"00",X"C8",X"3A",X"C3",X"72",X"E6",X"03",X"FE",X"00",X"28",X"05",X"FE",X"02",X"28",
		X"07",X"C9",X"3E",X"21",X"32",X"85",X"75",X"C9",X"3E",X"2C",X"32",X"85",X"75",X"C9",X"E5",X"D5",
		X"C5",X"2A",X"C8",X"72",X"11",X"04",X"00",X"19",X"22",X"C8",X"72",X"11",X"94",X"0C",X"AF",X"E5",
		X"ED",X"52",X"E1",X"20",X"06",X"21",X"84",X"0C",X"22",X"C8",X"72",X"11",X"49",X"70",X"01",X"04",
		X"00",X"ED",X"B0",X"C1",X"D1",X"E1",X"C9",X"3A",X"CD",X"72",X"3C",X"FE",X"0D",X"20",X"01",X"AF",
		X"32",X"CD",X"72",X"C9",X"3A",X"CE",X"72",X"3C",X"FE",X"03",X"32",X"CE",X"72",X"C0",X"AF",X"32",
		X"CE",X"72",X"3A",X"90",X"75",X"FE",X"33",X"20",X"06",X"3E",X"36",X"32",X"90",X"75",X"C9",X"3D",
		X"32",X"90",X"75",X"C9",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"00",X"3A",X"F7",X"72",X"FE",X"00",X"C8",X"CD",X"BD",X"0B",X"C9",X"3A",
		X"F7",X"72",X"FE",X"01",X"C0",X"AF",X"32",X"05",X"A0",X"ED",X"5B",X"00",X"73",X"0E",X"00",X"CD",
		X"4D",X"0D",X"28",X"27",X"ED",X"53",X"00",X"73",X"FE",X"FE",X"28",X"33",X"06",X"3E",X"CD",X"59",
		X"0D",X"ED",X"5B",X"02",X"73",X"0E",X"02",X"CD",X"4D",X"0D",X"28",X"23",X"ED",X"53",X"02",X"73",
		X"FE",X"FE",X"28",X"1B",X"06",X"3C",X"CD",X"59",X"0D",X"18",X"14",X"ED",X"5B",X"04",X"73",X"0E",
		X"04",X"CD",X"4D",X"0D",X"28",X"09",X"ED",X"53",X"04",X"73",X"06",X"3B",X"CD",X"59",X"0D",X"3E",
		X"01",X"32",X"05",X"A0",X"AF",X"32",X"06",X"A0",X"ED",X"5B",X"06",X"73",X"0E",X"00",X"CD",X"4D",
		X"0D",X"28",X"0F",X"ED",X"53",X"06",X"73",X"FE",X"FE",X"28",X"3C",X"06",X"3E",X"CD",X"53",X"0D",
		X"18",X"35",X"3A",X"BF",X"72",X"FE",X"00",X"20",X"2E",X"ED",X"5B",X"08",X"73",X"13",X"ED",X"53",
		X"08",X"73",X"1B",X"1A",X"FE",X"FF",X"20",X"08",X"21",X"0E",X"0E",X"22",X"08",X"73",X"18",X"17",
		X"FE",X"FE",X"28",X"13",X"06",X"08",X"DD",X"21",X"EA",X"5F",X"FE",X"01",X"28",X"04",X"DD",X"21",
		X"E1",X"5F",X"0E",X"06",X"CD",X"7E",X"0D",X"3E",X"01",X"32",X"06",X"A0",X"C9",X"1A",X"FE",X"FF",
		X"C8",X"13",X"C9",X"DD",X"21",X"5F",X"0E",X"18",X"04",X"DD",X"21",X"F3",X"5F",X"87",X"26",X"00",
		X"6F",X"11",X"1D",X"53",X"19",X"79",X"D3",X"08",X"7E",X"D3",X"09",X"0C",X"79",X"D3",X"08",X"23",
		X"7E",X"D3",X"09",X"3E",X"07",X"D3",X"08",X"78",X"D3",X"09",X"0E",X"08",X"06",X"06",X"79",X"DD",
		X"23",X"D3",X"08",X"DD",X"7E",X"00",X"D3",X"09",X"0C",X"10",X"F3",X"C9",X"11",X"76",X"0E",X"ED",
		X"53",X"00",X"73",X"ED",X"53",X"02",X"73",X"11",X"85",X"0E",X"ED",X"53",X"04",X"73",X"11",X"5E",
		X"0E",X"ED",X"53",X"06",X"73",X"11",X"93",X"0E",X"ED",X"53",X"08",X"73",X"3E",X"00",X"32",X"F7",
		X"72",X"C9",X"3A",X"0D",X"70",X"FE",X"01",X"C9",X"06",X"08",X"DD",X"21",X"00",X"98",X"DD",X"7E",
		X"02",X"3C",X"DD",X"77",X"02",X"DD",X"7E",X"03",X"3D",X"DD",X"77",X"03",X"DD",X"23",X"DD",X"23",
		X"DD",X"23",X"DD",X"23",X"10",X"E8",X"C9",X"3A",X"94",X"72",X"FE",X"01",X"C8",X"3A",X"9E",X"72",
		X"FE",X"01",X"C8",X"3A",X"F7",X"72",X"FE",X"01",X"C8",X"3A",X"62",X"70",X"FE",X"01",X"C8",X"AF",
		X"32",X"92",X"75",X"32",X"93",X"75",X"C9",X"3A",X"F7",X"72",X"FE",X"00",X"C8",X"3A",X"FD",X"70",
		X"FE",X"03",X"C8",X"3E",X"78",X"32",X"92",X"75",X"3E",X"E0",X"32",X"93",X"75",X"C9",X"01",X"FE",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"00",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"FE",X"FE",X"00",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"01",X"FE",X"FE",X"FE",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"00",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"00",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"01",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"FE",X"FE",X"FE",X"FE",X"00",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FF",X"3E",
		X"1F",X"1F",X"1F",X"FF",X"1E",X"00",X"0B",X"0C",X"0D",X"00",X"00",X"01",X"FE",X"FE",X"FE",X"FE",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"20",X"FE",X"FE",X"00",X"FF",X"1D",X"1C",
		X"1B",X"1A",X"19",X"FE",X"00",X"FF",X"25",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"FE",X"FE",X"FE",X"FF",X"19",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"FE",X"FF",X"3F",X"3F",X"FD",X"63",X"65",X"6B",X"FD",X"6F",X"75",X"4D",X"DC",X"6F",X"8D",X"22",
		X"79",X"09",X"05",X"6F",X"75",X"7F",X"ED",X"0B",X"6C",X"61",X"BE",X"4F",X"EF",X"6F",X"ED",X"67",
		X"7D",X"77",X"75",X"67",X"FD",X"5B",X"F9",X"7F",X"FD",X"6F",X"F9",X"7D",X"6D",X"63",X"4D",X"4F",
		X"AF",X"32",X"00",X"A0",X"32",X"03",X"A0",X"F3",X"3C",X"06",X"08",X"21",X"00",X"70",X"AF",X"4F",
		X"77",X"23",X"0D",X"20",X"FB",X"10",X"F8",X"31",X"F0",X"77",X"CD",X"8C",X"0D",X"CD",X"9F",X"19",
		X"ED",X"56",X"3E",X"01",X"32",X"00",X"A0",X"FB",X"21",X"3A",X"55",X"11",X"80",X"75",X"01",X"1C",
		X"00",X"ED",X"B0",X"21",X"92",X"54",X"11",X"9A",X"71",X"01",X"50",X"00",X"ED",X"B0",X"CD",X"1C",
		X"23",X"21",X"84",X"0C",X"22",X"C8",X"72",X"CD",X"8F",X"22",X"CD",X"9C",X"27",X"3E",X"40",X"32",
		X"35",X"70",X"3E",X"08",X"32",X"36",X"70",X"3E",X"01",X"32",X"01",X"A0",X"32",X"02",X"A0",X"3E",
		X"01",X"32",X"03",X"A0",X"CD",X"6A",X"13",X"3A",X"00",X"70",X"FE",X"00",X"28",X"E9",X"FE",X"01",
		X"20",X"1A",X"3A",X"4F",X"70",X"FE",X"01",X"28",X"29",X"CD",X"B5",X"19",X"CD",X"3D",X"1B",X"CD",
		X"9C",X"27",X"CD",X"E1",X"22",X"3E",X"01",X"32",X"4F",X"70",X"18",X"16",X"3A",X"4F",X"70",X"FE",
		X"00",X"28",X"E6",X"3A",X"50",X"70",X"FE",X"01",X"28",X"08",X"CD",X"08",X"23",X"3E",X"01",X"32",
		X"50",X"70",X"3A",X"0F",X"89",X"FE",X"1E",X"28",X"08",X"3A",X"2F",X"89",X"FE",X"1E",X"C2",X"27",
		X"0F",X"3A",X"00",X"70",X"FE",X"00",X"CA",X"27",X"0F",X"3A",X"02",X"70",X"E6",X"04",X"FE",X"04",
		X"28",X"21",X"3A",X"00",X"70",X"FE",X"02",X"DA",X"27",X"0F",X"3A",X"04",X"70",X"E6",X"04",X"FE",
		X"04",X"C2",X"27",X"0F",X"3A",X"00",X"70",X"3D",X"27",X"32",X"00",X"70",X"3E",X"02",X"32",X"0C",
		X"70",X"18",X"05",X"3E",X"01",X"32",X"0C",X"70",X"AF",X"32",X"0B",X"70",X"3A",X"00",X"70",X"3D",
		X"27",X"32",X"00",X"70",X"AF",X"32",X"76",X"72",X"32",X"79",X"72",X"3E",X"01",X"32",X"53",X"70",
		X"CD",X"5A",X"22",X"CD",X"B5",X"19",X"CD",X"6F",X"1A",X"CD",X"8F",X"22",X"CD",X"D4",X"11",X"CD",
		X"3C",X"1C",X"CD",X"89",X"12",X"CD",X"3E",X"23",X"3E",X"00",X"32",X"13",X"70",X"32",X"62",X"70",
		X"32",X"5B",X"70",X"32",X"F7",X"72",X"3E",X"10",X"32",X"35",X"70",X"3A",X"8D",X"72",X"FE",X"00",
		X"28",X"08",X"3A",X"FD",X"70",X"FE",X"03",X"CC",X"7F",X"1D",X"CD",X"B2",X"28",X"CD",X"40",X"22",
		X"CD",X"00",X"24",X"FD",X"21",X"88",X"75",X"11",X"35",X"70",X"DD",X"21",X"BD",X"72",X"CD",X"8A",
		X"23",X"CD",X"C7",X"23",X"FD",X"21",X"98",X"75",X"11",X"85",X"72",X"DD",X"21",X"BE",X"72",X"CD",
		X"8A",X"23",X"CD",X"C7",X"23",X"CD",X"34",X"22",X"3A",X"00",X"B8",X"3A",X"A1",X"72",X"FE",X"01",
		X"CC",X"3C",X"1C",X"CD",X"B0",X"21",X"CD",X"9C",X"27",X"3A",X"56",X"70",X"FE",X"02",X"CC",X"B2",
		X"11",X"3A",X"00",X"B8",X"CD",X"F1",X"1A",X"CD",X"B2",X"2F",X"E5",X"3A",X"20",X"70",X"FE",X"01",
		X"CA",X"07",X"11",X"3A",X"62",X"70",X"FE",X"01",X"CA",X"07",X"11",X"7E",X"CD",X"85",X"1E",X"CA",
		X"92",X"10",X"11",X"E0",X"FF",X"19",X"CD",X"85",X"1E",X"28",X"17",X"E1",X"E5",X"2B",X"CD",X"85",
		X"1E",X"28",X"0F",X"E1",X"E5",X"11",X"DF",X"FF",X"19",X"CD",X"85",X"1E",X"28",X"04",X"E1",X"E5",
		X"18",X"75",X"F5",X"CB",X"0F",X"CB",X"0F",X"E6",X"3F",X"32",X"44",X"70",X"F1",X"D1",X"E5",X"3A",
		X"BC",X"72",X"FE",X"01",X"20",X"61",X"CD",X"8D",X"26",X"AF",X"32",X"BC",X"72",X"3E",X"01",X"32",
		X"20",X"70",X"E5",X"21",X"86",X"0E",X"22",X"06",X"73",X"D5",X"ED",X"5B",X"10",X"73",X"E1",X"E5",
		X"AF",X"ED",X"52",X"D1",X"28",X"06",X"21",X"10",X"00",X"CD",X"6A",X"27",X"E1",X"3A",X"44",X"70",
		X"32",X"84",X"75",X"3E",X"2C",X"32",X"85",X"75",X"3E",X"FE",X"CD",X"35",X"27",X"CD",X"F0",X"26",
		X"22",X"2D",X"70",X"7E",X"E6",X"0F",X"F6",X"20",X"32",X"85",X"75",X"3E",X"00",X"CD",X"35",X"27",
		X"E1",X"E5",X"0E",X"10",X"CD",X"7D",X"21",X"E1",X"3A",X"44",X"70",X"FE",X"29",X"20",X"38",X"E5",
		X"CD",X"49",X"21",X"E1",X"C3",X"37",X"11",X"E1",X"E5",X"3A",X"20",X"70",X"FE",X"00",X"CA",X"19",
		X"11",X"CD",X"75",X"2F",X"20",X"03",X"E1",X"18",X"03",X"E1",X"18",X"1B",X"3A",X"5B",X"70",X"FE",
		X"01",X"28",X"11",X"3A",X"BC",X"72",X"FE",X"01",X"20",X"0D",X"3A",X"00",X"B8",X"AF",X"32",X"BC",
		X"72",X"22",X"10",X"73",X"CD",X"C1",X"1E",X"CD",X"28",X"1F",X"3A",X"00",X"B8",X"3A",X"F7",X"71",
		X"FE",X"00",X"20",X"43",X"3A",X"FD",X"71",X"FE",X"00",X"20",X"3C",X"3A",X"8B",X"72",X"FE",X"01",
		X"CC",X"1B",X"21",X"AF",X"32",X"8B",X"72",X"FD",X"21",X"84",X"72",X"FD",X"7E",X"04",X"FE",X"01",
		X"CC",X"2E",X"2F",X"DD",X"21",X"98",X"75",X"21",X"8A",X"72",X"CD",X"13",X"56",X"FD",X"21",X"84",
		X"72",X"FE",X"01",X"CC",X"2E",X"2F",X"ED",X"5B",X"04",X"73",X"1A",X"FE",X"FF",X"20",X"06",X"21",
		X"7E",X"0E",X"22",X"04",X"73",X"18",X"08",X"3E",X"01",X"32",X"8B",X"72",X"CD",X"3B",X"21",X"CD",
		X"47",X"14",X"FE",X"02",X"CA",X"DF",X"0F",X"FE",X"03",X"20",X"11",X"CD",X"3D",X"1B",X"CD",X"08",
		X"29",X"CD",X"B5",X"19",X"3E",X"01",X"32",X"03",X"A0",X"C3",X"27",X"0F",X"3A",X"00",X"B8",X"C3",
		X"FB",X"0F",X"3E",X"01",X"32",X"5C",X"70",X"CD",X"3D",X"1B",X"CD",X"49",X"12",X"CD",X"39",X"15",
		X"CD",X"89",X"12",X"21",X"D8",X"70",X"06",X"25",X"CD",X"64",X"13",X"3E",X"00",X"32",X"56",X"70",
		X"CD",X"3E",X"23",X"C9",X"21",X"69",X"70",X"AF",X"77",X"23",X"7D",X"FE",X"99",X"20",X"F8",X"7C",
		X"FE",X"71",X"20",X"F3",X"3A",X"07",X"70",X"CB",X"0F",X"E6",X"03",X"C6",X"01",X"32",X"D5",X"70",
		X"3C",X"32",X"6F",X"71",X"AF",X"32",X"4F",X"70",X"32",X"50",X"70",X"AF",X"21",X"26",X"70",X"06",
		X"06",X"77",X"23",X"10",X"FC",X"21",X"D8",X"70",X"CD",X"62",X"13",X"21",X"72",X"71",X"CD",X"62",
		X"13",X"21",X"EB",X"70",X"06",X"14",X"CD",X"64",X"13",X"21",X"85",X"71",X"06",X"12",X"CD",X"64",
		X"13",X"AF",X"32",X"56",X"70",X"32",X"69",X"70",X"32",X"D6",X"70",X"32",X"70",X"71",X"3C",X"32",
		X"FE",X"70",X"32",X"98",X"71",X"3A",X"9E",X"72",X"FE",X"00",X"28",X"06",X"3A",X"F6",X"72",X"32",
		X"FD",X"70",X"CD",X"67",X"12",X"CD",X"49",X"12",X"C9",X"AF",X"32",X"03",X"A0",X"CD",X"9F",X"19",
		X"CD",X"D2",X"19",X"CD",X"8F",X"22",X"3A",X"FD",X"70",X"FE",X"03",X"CC",X"B8",X"2D",X"CD",X"E0",
		X"16",X"3E",X"01",X"32",X"03",X"A0",X"C9",X"CD",X"74",X"12",X"CD",X"39",X"15",X"CD",X"63",X"15",
		X"CD",X"DE",X"20",X"C9",X"3A",X"FD",X"70",X"FE",X"03",X"CA",X"7D",X"12",X"C9",X"CD",X"75",X"2E",
		X"FD",X"21",X"69",X"70",X"E1",X"C9",X"CD",X"6F",X"1A",X"AF",X"32",X"34",X"70",X"3A",X"FD",X"70",
		X"FE",X"03",X"C4",X"28",X"16",X"3A",X"FD",X"70",X"FE",X"03",X"28",X"16",X"21",X"5A",X"55",X"11",
		X"80",X"75",X"01",X"20",X"00",X"ED",X"B0",X"21",X"3A",X"55",X"11",X"80",X"75",X"01",X"20",X"00",
		X"ED",X"B0",X"AF",X"32",X"76",X"72",X"32",X"79",X"72",X"32",X"20",X"70",X"32",X"5D",X"70",X"32",
		X"63",X"70",X"32",X"C3",X"72",X"32",X"FD",X"71",X"3E",X"50",X"CD",X"03",X"00",X"3E",X"02",X"32",
		X"49",X"70",X"32",X"4A",X"70",X"3E",X"01",X"32",X"43",X"70",X"32",X"CA",X"72",X"32",X"5C",X"70",
		X"3E",X"00",X"32",X"FA",X"71",X"CD",X"2D",X"13",X"3A",X"43",X"70",X"FE",X"40",X"CC",X"50",X"13",
		X"FE",X"60",X"CC",X"2D",X"13",X"FE",X"90",X"CC",X"50",X"13",X"FE",X"B0",X"CC",X"2D",X"13",X"FE",
		X"D0",X"20",X"E5",X"CD",X"50",X"13",X"AF",X"32",X"5C",X"70",X"21",X"5F",X"8A",X"11",X"4C",X"58",
		X"CD",X"49",X"19",X"01",X"E0",X"FF",X"00",X"3A",X"FE",X"70",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",
		X"FE",X"00",X"28",X"02",X"77",X"09",X"3A",X"FE",X"70",X"E6",X"0F",X"77",X"C9",X"21",X"5F",X"8A",
		X"11",X"9E",X"57",X"CD",X"49",X"19",X"21",X"BF",X"99",X"3E",X"0F",X"06",X"0A",X"CD",X"60",X"19",
		X"CD",X"9C",X"27",X"AF",X"32",X"BF",X"72",X"32",X"C0",X"72",X"3E",X"20",X"32",X"35",X"70",X"C9",
		X"21",X"5F",X"8A",X"11",X"E0",X"FF",X"06",X"06",X"3E",X"FF",X"77",X"19",X"10",X"FA",X"CD",X"DB",
		X"02",X"C9",X"06",X"09",X"AF",X"77",X"23",X"10",X"FB",X"C9",X"3A",X"00",X"70",X"FE",X"00",X"C0",
		X"3E",X"01",X"32",X"5D",X"70",X"CD",X"67",X"1B",X"CD",X"3D",X"1B",X"3E",X"00",X"32",X"03",X"A0",
		X"CD",X"9E",X"2C",X"CD",X"B5",X"19",X"3E",X"00",X"32",X"5D",X"70",X"3E",X"01",X"32",X"03",X"A0",
		X"3A",X"FD",X"70",X"3C",X"FE",X"07",X"06",X"00",X"28",X"0C",X"FE",X"03",X"06",X"04",X"28",X"06",
		X"32",X"FD",X"70",X"C3",X"6A",X"13",X"78",X"32",X"FD",X"70",X"C3",X"6A",X"13",X"FD",X"21",X"FB",
		X"5E",X"3A",X"FD",X"70",X"FE",X"00",X"C8",X"FD",X"21",X"29",X"5F",X"FE",X"01",X"C8",X"FD",X"21",
		X"CD",X"5E",X"FE",X"02",X"C8",X"FD",X"21",X"85",X"5F",X"FE",X"06",X"C8",X"FD",X"21",X"57",X"5F",
		X"FE",X"04",X"C8",X"FD",X"21",X"B3",X"5F",X"FE",X"05",X"C9",X"CD",X"FB",X"2E",X"E6",X"3F",X"FE",
		X"10",X"D8",X"FD",X"7E",X"00",X"FE",X"00",X"C8",X"2A",X"AF",X"72",X"AF",X"FD",X"77",X"00",X"DD",
		X"77",X"06",X"CD",X"A7",X"1E",X"CD",X"3C",X"1C",X"3E",X"01",X"32",X"3E",X"70",X"C9",X"11",X"05",
		X"09",X"CD",X"FE",X"18",X"7E",X"FE",X"C8",X"20",X"0A",X"3A",X"3E",X"70",X"FE",X"01",X"28",X"07",
		X"3E",X"01",X"C9",X"AF",X"32",X"3E",X"70",X"3E",X"00",X"C9",X"FD",X"21",X"69",X"70",X"CD",X"6D",
		X"15",X"FD",X"7E",X"02",X"E6",X"30",X"B9",X"28",X"09",X"FD",X"23",X"FD",X"23",X"FD",X"23",X"10",
		X"F0",X"C9",X"FD",X"7E",X"02",X"E6",X"CF",X"FD",X"77",X"02",X"CD",X"F0",X"26",X"CD",X"AB",X"2F",
		X"FD",X"75",X"00",X"FD",X"74",X"01",X"C9",X"3A",X"13",X"70",X"FE",X"00",X"C8",X"CD",X"8C",X"0D",
		X"21",X"D2",X"36",X"CD",X"9B",X"0B",X"21",X"D2",X"36",X"CD",X"B5",X"0B",X"21",X"D8",X"36",X"CD",
		X"CF",X"0B",X"CD",X"00",X"24",X"3A",X"34",X"70",X"FE",X"00",X"28",X"08",X"2A",X"AF",X"72",X"0E",
		X"20",X"CD",X"1A",X"14",X"3A",X"20",X"70",X"FE",X"00",X"28",X"08",X"2A",X"AD",X"72",X"0E",X"10",
		X"CD",X"1A",X"14",X"3E",X"3A",X"32",X"80",X"75",X"AF",X"32",X"58",X"70",X"32",X"14",X"70",X"32",
		X"7F",X"72",X"3C",X"32",X"5D",X"70",X"21",X"38",X"5B",X"22",X"59",X"70",X"AF",X"32",X"20",X"70",
		X"32",X"34",X"70",X"CD",X"49",X"1B",X"21",X"9F",X"8A",X"11",X"51",X"58",X"CD",X"54",X"23",X"3A",
		X"0C",X"70",X"FE",X"02",X"28",X"32",X"3A",X"D5",X"70",X"FE",X"00",X"28",X"41",X"3A",X"07",X"70",
		X"E6",X"08",X"FE",X"08",X"28",X"07",X"3A",X"D5",X"70",X"3D",X"32",X"D5",X"70",X"CD",X"5A",X"22",
		X"CD",X"B5",X"19",X"CD",X"3D",X"1B",X"CD",X"8F",X"22",X"CD",X"6F",X"1A",X"CD",X"D2",X"19",X"CD",
		X"8F",X"22",X"CD",X"E0",X"16",X"3E",X"02",X"C9",X"CD",X"16",X"28",X"3A",X"D5",X"70",X"FE",X"00",
		X"20",X"CB",X"CD",X"16",X"28",X"3A",X"D5",X"70",X"FE",X"00",X"28",X"02",X"18",X"BF",X"CD",X"94",
		X"22",X"21",X"6E",X"8A",X"11",X"A1",X"56",X"CD",X"49",X"19",X"3E",X"00",X"32",X"D6",X"70",X"32",
		X"70",X"71",X"3E",X"01",X"32",X"42",X"70",X"AF",X"32",X"53",X"70",X"3A",X"42",X"70",X"FE",X"70",
		X"20",X"F9",X"AF",X"32",X"42",X"70",X"3E",X"01",X"32",X"01",X"A0",X"32",X"02",X"A0",X"3E",X"00",
		X"32",X"03",X"A0",X"CD",X"68",X"19",X"3E",X"03",X"C9",X"FD",X"21",X"69",X"70",X"FD",X"22",X"CB",
		X"72",X"CD",X"74",X"12",X"11",X"16",X"70",X"CD",X"B6",X"15",X"06",X"09",X"DD",X"7E",X"00",X"12",
		X"DD",X"23",X"13",X"10",X"F7",X"CD",X"6D",X"15",X"CD",X"82",X"15",X"FD",X"2A",X"CB",X"72",X"CD",
		X"EA",X"15",X"C9",X"FD",X"21",X"03",X"71",X"FD",X"22",X"CB",X"72",X"18",X"D4",X"06",X"11",X"3A",
		X"FD",X"70",X"FE",X"00",X"C8",X"06",X"18",X"FE",X"01",X"C8",X"06",X"09",X"FE",X"03",X"C8",X"06",
		X"23",X"C9",X"DD",X"21",X"86",X"5C",X"3A",X"FD",X"70",X"FE",X"00",X"C8",X"DD",X"21",X"58",X"5D",
		X"FE",X"01",X"C8",X"DD",X"21",X"AB",X"5B",X"FE",X"02",X"C8",X"DD",X"21",X"EF",X"5C",X"FE",X"04",
		X"C8",X"DD",X"21",X"C1",X"5D",X"FE",X"06",X"C8",X"DD",X"21",X"2A",X"5E",X"FE",X"05",X"C8",X"DD",
		X"21",X"1D",X"5C",X"FE",X"03",X"C9",X"DD",X"21",X"12",X"5B",X"3A",X"FD",X"70",X"FE",X"00",X"C8",
		X"DD",X"21",X"24",X"5B",X"FE",X"01",X"C8",X"DD",X"21",X"00",X"5B",X"FE",X"02",X"C8",X"DD",X"21",
		X"1B",X"5B",X"FE",X"04",X"C8",X"DD",X"21",X"2D",X"5B",X"FE",X"06",X"C8",X"DD",X"21",X"36",X"5B",
		X"FE",X"05",X"C8",X"DD",X"21",X"09",X"5B",X"FE",X"03",X"C9",X"CD",X"FB",X"2E",X"CD",X"FB",X"2E",
		X"11",X"16",X"70",X"E6",X"0F",X"3C",X"FE",X"0A",X"30",X"F0",X"F5",X"83",X"5F",X"1B",X"1A",X"FE",
		X"00",X"28",X"22",X"F1",X"EB",X"35",X"EB",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"FD",X"75",X"00",
		X"FD",X"74",X"01",X"FD",X"77",X"02",X"DD",X"23",X"DD",X"23",X"DD",X"23",X"FD",X"23",X"FD",X"23",
		X"FD",X"23",X"10",X"C6",X"C9",X"F1",X"18",X"C2",X"FD",X"21",X"69",X"70",X"E5",X"21",X"F3",X"36",
		X"22",X"80",X"72",X"E1",X"CD",X"6D",X"15",X"C5",X"FD",X"6E",X"00",X"FD",X"66",X"01",X"CD",X"9D",
		X"2F",X"CD",X"A2",X"2F",X"E5",X"CD",X"05",X"27",X"2A",X"80",X"72",X"CD",X"BD",X"0B",X"AF",X"32",
		X"7C",X"72",X"F3",X"2A",X"80",X"72",X"23",X"23",X"23",X"22",X"80",X"72",X"FB",X"E1",X"CD",X"F0",
		X"26",X"FD",X"7E",X"02",X"E6",X"0F",X"F6",X"20",X"CD",X"35",X"27",X"C1",X"FD",X"23",X"FD",X"23",
		X"FD",X"23",X"3E",X"01",X"32",X"43",X"70",X"E5",X"21",X"68",X"5B",X"22",X"59",X"70",X"3E",X"00",
		X"32",X"58",X"70",X"E1",X"3A",X"D6",X"70",X"FE",X"01",X"28",X"0B",X"3A",X"43",X"70",X"FE",X"07",
		X"20",X"F9",X"AF",X"32",X"43",X"70",X"10",X"9F",X"3E",X"01",X"32",X"D6",X"70",X"C9",X"FD",X"21",
		X"69",X"70",X"CD",X"6D",X"15",X"C5",X"FD",X"6E",X"00",X"FD",X"66",X"01",X"CD",X"9D",X"2F",X"CD",
		X"A2",X"2F",X"E5",X"CD",X"05",X"27",X"E1",X"CD",X"F0",X"26",X"FD",X"7E",X"02",X"E6",X"0F",X"F6",
		X"20",X"CD",X"35",X"27",X"C1",X"FD",X"23",X"FD",X"23",X"FD",X"23",X"3E",X"01",X"32",X"43",X"70",
		X"E5",X"21",X"68",X"5B",X"22",X"59",X"70",X"3E",X"00",X"32",X"58",X"70",X"E1",X"10",X"C6",X"C9",
		X"CD",X"10",X"17",X"3A",X"FD",X"70",X"FE",X"03",X"C8",X"3E",X"0E",X"F5",X"DD",X"46",X"00",X"DD",
		X"4E",X"01",X"C5",X"DD",X"46",X"02",X"DD",X"4E",X"03",X"C5",X"DD",X"7E",X"06",X"DD",X"66",X"04",
		X"DD",X"6E",X"05",X"CD",X"4A",X"17",X"11",X"07",X"00",X"DD",X"19",X"F1",X"3D",X"20",X"DC",X"C9",
		X"DD",X"21",X"7F",X"50",X"3A",X"FD",X"70",X"FE",X"00",X"C8",X"DD",X"21",X"43",X"51",X"FE",X"01",
		X"C8",X"DD",X"21",X"1D",X"50",X"FE",X"02",X"C8",X"DD",X"21",X"E1",X"50",X"FE",X"04",X"C8",X"DD",
		X"21",X"A5",X"51",X"FE",X"06",X"C8",X"DD",X"21",X"07",X"52",X"FE",X"05",X"C8",X"C9",X"ED",X"4B",
		X"A3",X"72",X"E5",X"21",X"88",X"53",X"ED",X"B1",X"E1",X"C9",X"FD",X"E1",X"11",X"20",X"00",X"C1",
		X"2B",X"77",X"10",X"FC",X"41",X"37",X"3F",X"ED",X"52",X"77",X"10",X"F9",X"C1",X"23",X"77",X"10",
		X"FC",X"41",X"19",X"77",X"10",X"FC",X"FD",X"E5",X"C9",X"DD",X"21",X"90",X"75",X"11",X"0E",X"0E",
		X"CD",X"FE",X"18",X"CD",X"FA",X"17",X"C8",X"DD",X"21",X"90",X"75",X"11",X"00",X"0E",X"CD",X"FE",
		X"18",X"CD",X"FA",X"17",X"C9",X"DD",X"21",X"90",X"75",X"11",X"0E",X"00",X"CD",X"FE",X"18",X"CD",
		X"FA",X"17",X"C8",X"DD",X"21",X"90",X"75",X"11",X"00",X"00",X"CD",X"FE",X"18",X"CD",X"FA",X"17",
		X"C9",X"DD",X"21",X"90",X"75",X"11",X"0C",X"00",X"CD",X"FE",X"18",X"CD",X"FA",X"17",X"C8",X"DD",
		X"21",X"90",X"75",X"11",X"0C",X"0E",X"CD",X"FE",X"18",X"CD",X"FA",X"17",X"C9",X"DD",X"21",X"90",
		X"75",X"11",X"00",X"00",X"CD",X"FE",X"18",X"CD",X"FA",X"17",X"C8",X"DD",X"21",X"90",X"75",X"11",
		X"00",X"0E",X"CD",X"FE",X"18",X"CD",X"FA",X"17",X"C9",X"DD",X"21",X"80",X"75",X"11",X"08",X"09",
		X"CD",X"FE",X"18",X"CD",X"FA",X"17",X"C8",X"DD",X"21",X"80",X"75",X"11",X"05",X"09",X"CD",X"FE",
		X"18",X"CD",X"FA",X"17",X"C8",X"AF",X"32",X"12",X"70",X"C9",X"7E",X"E5",X"21",X"27",X"55",X"01",
		X"13",X"00",X"ED",X"B1",X"E1",X"C9",X"3A",X"12",X"70",X"FE",X"00",X"C0",X"CD",X"FB",X"2E",X"E6",
		X"01",X"32",X"49",X"70",X"CD",X"FB",X"2E",X"47",X"10",X"FE",X"CD",X"FB",X"2E",X"E6",X"01",X"32",
		X"4A",X"70",X"3A",X"4B",X"70",X"2F",X"E6",X"01",X"32",X"4B",X"70",X"CD",X"FB",X"2E",X"E6",X"01",
		X"32",X"4C",X"70",X"3A",X"49",X"70",X"47",X"3A",X"4B",X"70",X"B0",X"FE",X"00",X"28",X"C7",X"3E",
		X"01",X"32",X"12",X"70",X"C9",X"3A",X"12",X"70",X"FE",X"00",X"C0",X"CD",X"FB",X"2E",X"E6",X"01",
		X"32",X"49",X"70",X"CD",X"FB",X"2E",X"47",X"10",X"FE",X"CD",X"FB",X"2E",X"E6",X"01",X"32",X"4A",
		X"70",X"CD",X"FB",X"2E",X"E6",X"01",X"32",X"4B",X"70",X"3A",X"4C",X"70",X"2F",X"E6",X"01",X"32",
		X"4C",X"70",X"3A",X"49",X"70",X"47",X"3A",X"4B",X"70",X"B0",X"FE",X"00",X"28",X"C7",X"3E",X"01",
		X"32",X"12",X"70",X"C9",X"DD",X"21",X"E2",X"54",X"11",X"05",X"00",X"7E",X"47",X"DD",X"7E",X"00",
		X"B8",X"28",X"0A",X"DD",X"19",X"DD",X"7E",X"00",X"FE",X"00",X"C8",X"18",X"EE",X"3A",X"12",X"70",
		X"FE",X"00",X"C0",X"3A",X"11",X"70",X"5F",X"16",X"00",X"DD",X"7E",X"00",X"32",X"12",X"70",X"DD",
		X"19",X"DD",X"7E",X"00",X"32",X"11",X"70",X"E5",X"21",X"97",X"5E",X"11",X"03",X"00",X"CD",X"FB",
		X"2E",X"E6",X"0F",X"FE",X"00",X"28",X"F7",X"47",X"19",X"10",X"FD",X"EB",X"1A",X"6F",X"13",X"1A",
		X"67",X"13",X"1A",X"77",X"21",X"97",X"5E",X"11",X"03",X"00",X"CD",X"FB",X"2E",X"E6",X"0F",X"FE",
		X"00",X"28",X"F7",X"47",X"19",X"10",X"FD",X"EB",X"1A",X"6F",X"13",X"1A",X"67",X"13",X"3E",X"10",
		X"77",X"E1",X"C9",X"E5",X"7E",X"21",X"93",X"5E",X"01",X"05",X"00",X"ED",X"B1",X"E1",X"D5",X"CD",
		X"18",X"19",X"D1",X"CD",X"07",X"19",X"C9",X"DD",X"7E",X"03",X"83",X"CB",X"3F",X"CB",X"3F",X"CB",
		X"3F",X"85",X"6F",X"7C",X"CE",X"00",X"67",X"C9",X"DD",X"7E",X"02",X"82",X"FE",X"80",X"38",X"15",
		X"2F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"FE",X"00",X"C8",X"47",X"11",X"20",X"00",X"21",X"00",
		X"88",X"19",X"10",X"FD",X"C9",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"FE",X"00",X"C8",X"47",X"11",
		X"E0",X"FF",X"21",X"E0",X"8B",X"19",X"10",X"FD",X"C9",X"F5",X"3A",X"00",X"A8",X"E6",X"40",X"FE",
		X"40",X"28",X"08",X"E5",X"EB",X"11",X"87",X"02",X"19",X"EB",X"E1",X"F1",X"CD",X"54",X"23",X"C9",
		X"11",X"20",X"00",X"77",X"19",X"10",X"FC",X"C9",X"06",X"08",X"21",X"00",X"98",X"0E",X"00",X"77",
		X"23",X"F5",X"3A",X"00",X"B8",X"F1",X"0D",X"20",X"F6",X"10",X"F2",X"3E",X"0A",X"21",X"40",X"98",
		X"06",X"1C",X"CD",X"60",X"19",X"3E",X"05",X"21",X"41",X"98",X"06",X"1C",X"CD",X"60",X"19",X"3E",
		X"04",X"21",X"7F",X"98",X"06",X"1C",X"CD",X"60",X"19",X"3E",X"00",X"32",X"5F",X"98",X"C9",X"06",
		X"04",X"3E",X"FF",X"21",X"00",X"88",X"0E",X"00",X"77",X"23",X"F5",X"3A",X"00",X"B8",X"F1",X"0D",
		X"20",X"F6",X"10",X"F2",X"C9",X"21",X"01",X"88",X"11",X"20",X"00",X"0E",X"1D",X"23",X"E5",X"06",
		X"20",X"3E",X"FF",X"77",X"19",X"10",X"FC",X"E1",X"0D",X"79",X"FE",X"00",X"20",X"EF",X"CD",X"9C",
		X"27",X"C9",X"CD",X"E1",X"19",X"11",X"00",X"88",X"01",X"00",X"04",X"ED",X"B0",X"CD",X"B0",X"1F",
		X"C9",X"21",X"00",X"38",X"3A",X"FD",X"70",X"FE",X"00",X"C8",X"21",X"00",X"3C",X"FE",X"01",X"C8",
		X"21",X"00",X"40",X"FE",X"02",X"C8",X"21",X"00",X"44",X"FE",X"04",X"C8",X"21",X"00",X"48",X"FE",
		X"06",X"C8",X"21",X"00",X"4C",X"FE",X"05",X"C8",X"FE",X"03",X"CC",X"B8",X"2D",X"E1",X"C9",X"CD",
		X"82",X"15",X"FD",X"21",X"69",X"70",X"CD",X"6D",X"15",X"11",X"20",X"00",X"19",X"7D",X"DD",X"BE",
		X"00",X"20",X"3D",X"7C",X"DD",X"BE",X"01",X"20",X"37",X"7E",X"E6",X"0F",X"DD",X"BE",X"02",X"20",
		X"2F",X"11",X"20",X"00",X"AF",X"ED",X"52",X"5C",X"3A",X"2E",X"70",X"BB",X"20",X"07",X"5D",X"3A",
		X"2D",X"70",X"BB",X"28",X"1B",X"21",X"00",X"01",X"FD",X"7E",X"02",X"E6",X"40",X"FE",X"40",X"28",
		X"0B",X"FD",X"7E",X"02",X"F6",X"40",X"FD",X"77",X"02",X"CD",X"6A",X"27",X"CD",X"9C",X"27",X"C9",
		X"DD",X"23",X"DD",X"23",X"DD",X"23",X"FD",X"23",X"FD",X"23",X"FD",X"23",X"10",X"AF",X"C9",X"3A",
		X"0C",X"70",X"FE",X"01",X"C8",X"3E",X"01",X"32",X"42",X"70",X"CD",X"21",X"1B",X"21",X"75",X"8A",
		X"CD",X"49",X"19",X"3E",X"06",X"08",X"CD",X"9C",X"1A",X"3A",X"42",X"70",X"FE",X"00",X"28",X"02",
		X"18",X"F7",X"21",X"75",X"8A",X"11",X"6C",X"57",X"CD",X"49",X"19",X"C9",X"21",X"94",X"8A",X"06",
		X"08",X"0E",X"01",X"11",X"E0",X"FF",X"3E",X"AE",X"C5",X"CD",X"E5",X"1A",X"3E",X"B4",X"19",X"CD",
		X"E5",X"1A",X"10",X"FA",X"19",X"3E",X"B3",X"CD",X"E5",X"1A",X"41",X"3E",X"B2",X"23",X"CD",X"E5",
		X"1A",X"10",X"FA",X"23",X"3E",X"B1",X"CD",X"E5",X"1A",X"C1",X"11",X"20",X"00",X"19",X"3E",X"B4",
		X"CD",X"E5",X"1A",X"10",X"F8",X"19",X"3E",X"B0",X"CD",X"E5",X"1A",X"41",X"3E",X"AF",X"2B",X"CD",
		X"E5",X"1A",X"10",X"FA",X"C9",X"77",X"E5",X"F5",X"CD",X"F0",X"26",X"F1",X"08",X"77",X"E1",X"08",
		X"C9",X"3A",X"53",X"70",X"FE",X"01",X"C0",X"3A",X"CA",X"72",X"FE",X"20",X"D8",X"FE",X"30",X"30",
		X"03",X"C3",X"13",X"1B",X"3E",X"01",X"32",X"CA",X"72",X"CD",X"21",X"1B",X"11",X"6C",X"57",X"CD",
		X"49",X"19",X"C9",X"CD",X"21",X"1B",X"7E",X"FE",X"FF",X"C0",X"CD",X"49",X"19",X"CD",X"34",X"1B",
		X"C9",X"3A",X"0B",X"70",X"21",X"A0",X"8B",X"11",X"5A",X"57",X"FE",X"01",X"C0",X"11",X"63",X"57",
		X"21",X"20",X"89",X"C9",X"3E",X"0A",X"21",X"40",X"98",X"CD",X"80",X"23",X"C9",X"21",X"5A",X"55",
		X"11",X"80",X"75",X"01",X"1C",X"00",X"ED",X"B0",X"C9",X"06",X"03",X"3E",X"1F",X"3C",X"32",X"81",
		X"75",X"3E",X"01",X"32",X"43",X"70",X"3A",X"43",X"70",X"FE",X"04",X"20",X"F9",X"3A",X"81",X"75",
		X"FE",X"2F",X"20",X"E9",X"10",X"E5",X"C9",X"11",X"AA",X"53",X"21",X"86",X"8A",X"3E",X"0E",X"08",
		X"CD",X"6B",X"23",X"11",X"B5",X"53",X"21",X"87",X"8A",X"3E",X"0E",X"08",X"CD",X"6B",X"23",X"11",
		X"C0",X"53",X"21",X"88",X"8A",X"3E",X"0E",X"08",X"CD",X"6B",X"23",X"11",X"CB",X"53",X"21",X"6B",
		X"8A",X"3E",X"0F",X"08",X"CD",X"6B",X"23",X"3A",X"00",X"A8",X"E6",X"40",X"FE",X"40",X"20",X"0A",
		X"3E",X"BD",X"32",X"8B",X"89",X"3E",X"0F",X"32",X"8B",X"99",X"3E",X"01",X"32",X"43",X"70",X"11",
		X"D4",X"53",X"21",X"4E",X"8B",X"3E",X"2D",X"08",X"CD",X"6B",X"23",X"11",X"EB",X"53",X"21",X"4F",
		X"8B",X"3E",X"2D",X"08",X"CD",X"6B",X"23",X"11",X"02",X"54",X"21",X"50",X"8B",X"3E",X"2D",X"08",
		X"CD",X"6B",X"23",X"11",X"19",X"54",X"21",X"51",X"8B",X"3E",X"2D",X"08",X"CD",X"6B",X"23",X"11",
		X"30",X"54",X"21",X"52",X"8B",X"3E",X"2D",X"08",X"CD",X"6B",X"23",X"11",X"47",X"54",X"21",X"53",
		X"8B",X"3E",X"2D",X"08",X"CD",X"6B",X"23",X"CD",X"8F",X"24",X"3E",X"00",X"32",X"94",X"72",X"3E",
		X"0A",X"32",X"35",X"70",X"3E",X"01",X"32",X"43",X"70",X"3A",X"43",X"70",X"FE",X"30",X"C8",X"3A",
		X"00",X"70",X"FE",X"00",X"C0",X"18",X"F2",X"DD",X"21",X"88",X"75",X"3A",X"11",X"70",X"FE",X"01",
		X"CD",X"69",X"17",X"3A",X"11",X"70",X"FE",X"02",X"CD",X"85",X"17",X"3A",X"11",X"70",X"FE",X"03",
		X"CD",X"A1",X"17",X"3A",X"11",X"70",X"FE",X"04",X"CD",X"BD",X"17",X"C9",X"3E",X"01",X"32",X"5E",
		X"70",X"3A",X"00",X"B8",X"CD",X"5E",X"1C",X"3A",X"00",X"B8",X"CD",X"CD",X"1C",X"3A",X"00",X"B8",
		X"CD",X"7F",X"1D",X"3A",X"00",X"B8",X"AF",X"32",X"5E",X"70",X"32",X"A1",X"72",X"C9",X"CD",X"6D",
		X"15",X"D9",X"21",X"00",X"72",X"11",X"03",X"00",X"CD",X"82",X"15",X"CD",X"6D",X"15",X"FD",X"21",
		X"69",X"70",X"DD",X"7E",X"00",X"FD",X"BE",X"00",X"28",X"0D",X"FD",X"19",X"10",X"F4",X"3E",X"00",
		X"77",X"23",X"77",X"23",X"77",X"18",X"16",X"DD",X"7E",X"01",X"FD",X"BE",X"01",X"20",X"EB",X"FD",
		X"7E",X"00",X"77",X"FD",X"7E",X"01",X"23",X"77",X"FD",X"7E",X"02",X"23",X"77",X"23",X"DD",X"19",
		X"D9",X"05",X"D9",X"20",X"C6",X"C9",X"21",X"51",X"5B",X"3A",X"FD",X"70",X"FE",X"00",X"C8",X"21",
		X"75",X"5B",X"FE",X"01",X"C8",X"21",X"3F",X"5B",X"FE",X"02",X"C8",X"21",X"63",X"5B",X"FE",X"04",
		X"C8",X"21",X"87",X"5B",X"FE",X"06",X"C8",X"21",X"99",X"5B",X"FE",X"05",X"C9",X"CD",X"B6",X"15",
		X"0E",X"01",X"FD",X"21",X"00",X"72",X"CD",X"A6",X"1C",X"DD",X"46",X"00",X"16",X"01",X"FD",X"7E",
		X"02",X"E6",X"0F",X"B9",X"28",X"02",X"16",X"00",X"FD",X"23",X"FD",X"23",X"FD",X"23",X"10",X"EE",
		X"7A",X"FE",X"00",X"C4",X"01",X"1D",X"0C",X"DD",X"23",X"79",X"FE",X"0A",X"C8",X"23",X"23",X"18",
		X"D8",X"E5",X"21",X"D7",X"70",X"7D",X"81",X"6F",X"7E",X"FE",X"01",X"28",X"63",X"3E",X"01",X"77",
		X"E1",X"E5",X"D5",X"EB",X"1A",X"6F",X"13",X"1A",X"67",X"D1",X"E5",X"CD",X"75",X"2F",X"E1",X"20",
		X"0A",X"3E",X"A4",X"CD",X"4D",X"27",X"3E",X"20",X"CD",X"29",X"22",X"E5",X"DD",X"E5",X"21",X"E9",
		X"70",X"DD",X"21",X"E1",X"70",X"41",X"23",X"23",X"DD",X"23",X"10",X"FA",X"DD",X"36",X"00",X"01",
		X"ED",X"53",X"F8",X"71",X"EB",X"DD",X"E1",X"E1",X"E5",X"EB",X"73",X"23",X"72",X"ED",X"5B",X"F8",
		X"71",X"E1",X"E5",X"CD",X"75",X"2F",X"E1",X"20",X"08",X"CD",X"F0",X"26",X"3E",X"20",X"CD",X"35",
		X"27",X"06",X"05",X"3A",X"F7",X"71",X"FE",X"99",X"28",X"08",X"00",X"CD",X"1F",X"00",X"10",X"F3",
		X"E1",X"C9",X"3E",X"01",X"32",X"FD",X"71",X"AF",X"32",X"F7",X"71",X"10",X"E6",X"18",X"F1",X"3A",
		X"FD",X"70",X"FE",X"03",X"20",X"13",X"CD",X"BC",X"2E",X"C0",X"3A",X"F7",X"71",X"FE",X"00",X"20",
		X"34",X"CD",X"1C",X"23",X"CD",X"8C",X"0D",X"18",X"47",X"CD",X"B6",X"15",X"0E",X"01",X"FD",X"21",
		X"00",X"72",X"21",X"22",X"8A",X"DD",X"46",X"00",X"16",X"01",X"FD",X"7E",X"02",X"E6",X"0F",X"B9",
		X"C2",X"6B",X"1E",X"FD",X"23",X"FD",X"23",X"FD",X"23",X"10",X"EF",X"0C",X"DD",X"23",X"CD",X"6E",
		X"1E",X"28",X"02",X"18",X"E0",X"21",X"D0",X"8A",X"11",X"32",X"58",X"CD",X"49",X"19",X"CD",X"8C",
		X"0D",X"CD",X"1C",X"23",X"21",X"83",X"37",X"CD",X"9B",X"0B",X"21",X"DD",X"37",X"CD",X"B5",X"0B",
		X"3E",X"01",X"32",X"A2",X"72",X"AF",X"32",X"D6",X"70",X"3A",X"FE",X"70",X"C6",X"01",X"27",X"32",
		X"FE",X"70",X"3A",X"FD",X"70",X"3C",X"FE",X"07",X"20",X"01",X"AF",X"32",X"FD",X"70",X"21",X"D8",
		X"70",X"CD",X"62",X"13",X"3E",X"02",X"32",X"56",X"70",X"AF",X"32",X"F6",X"71",X"3C",X"32",X"FA",
		X"71",X"32",X"5D",X"70",X"3A",X"F7",X"71",X"FE",X"00",X"28",X"17",X"3D",X"27",X"32",X"F7",X"71",
		X"21",X"00",X"01",X"CD",X"6A",X"27",X"CD",X"9C",X"27",X"3E",X"FF",X"3D",X"FE",X"00",X"20",X"FB",
		X"18",X"E2",X"3A",X"FD",X"71",X"FE",X"00",X"28",X"11",X"AF",X"32",X"FD",X"71",X"21",X"00",X"01",
		X"CD",X"6A",X"27",X"3E",X"99",X"32",X"F7",X"71",X"18",X"CA",X"3E",X"01",X"32",X"43",X"70",X"3A",
		X"43",X"70",X"FE",X"FF",X"28",X"02",X"18",X"F7",X"3E",X"01",X"32",X"43",X"70",X"3A",X"43",X"70",
		X"FE",X"80",X"28",X"02",X"18",X"F7",X"AF",X"32",X"43",X"70",X"C9",X"3E",X"01",X"C9",X"3A",X"FD",
		X"70",X"FE",X"00",X"20",X"04",X"79",X"FE",X"04",X"C9",X"FE",X"01",X"20",X"04",X"79",X"FE",X"07",
		X"C9",X"79",X"FE",X"0A",X"C9",X"E5",X"01",X"0B",X"00",X"2A",X"40",X"70",X"ED",X"B1",X"11",X"0B",
		X"00",X"2A",X"40",X"70",X"19",X"22",X"40",X"70",X"E1",X"C9",X"DD",X"7E",X"04",X"CB",X"07",X"CB",
		X"07",X"E6",X"FC",X"CD",X"4D",X"27",X"C9",X"E5",X"0E",X"20",X"CD",X"1A",X"14",X"E1",X"E5",X"CD",
		X"F0",X"26",X"3A",X"8D",X"75",X"E6",X"0F",X"F6",X"20",X"CD",X"35",X"27",X"E1",X"CD",X"05",X"27",
		X"C9",X"AF",X"32",X"5B",X"70",X"32",X"20",X"70",X"32",X"87",X"75",X"3E",X"2C",X"32",X"81",X"75",
		X"AF",X"32",X"7C",X"72",X"E5",X"21",X"94",X"0E",X"22",X"06",X"73",X"E1",X"E5",X"2A",X"AD",X"72",
		X"DD",X"21",X"80",X"75",X"CD",X"9A",X"1E",X"E1",X"E5",X"2A",X"AD",X"72",X"CD",X"F0",X"26",X"3A",
		X"85",X"75",X"E6",X"0F",X"F6",X"20",X"F5",X"CD",X"35",X"27",X"3A",X"84",X"75",X"FE",X"29",X"20",
		X"09",X"F1",X"E1",X"2A",X"AD",X"72",X"CD",X"F3",X"20",X"C9",X"F1",X"CD",X"0F",X"1A",X"E1",X"2A",
		X"AD",X"72",X"0E",X"10",X"CD",X"1A",X"14",X"3A",X"A0",X"72",X"FE",X"01",X"28",X"04",X"CD",X"3C",
		X"1C",X"C9",X"3E",X"01",X"32",X"A1",X"72",X"C9",X"CD",X"D9",X"17",X"DD",X"21",X"88",X"75",X"FD",
		X"21",X"34",X"70",X"FD",X"7E",X"04",X"FE",X"01",X"CC",X"DA",X"13",X"FD",X"21",X"34",X"70",X"FD",
		X"7E",X"04",X"FE",X"01",X"20",X"04",X"CD",X"2E",X"2F",X"C9",X"DD",X"21",X"88",X"75",X"21",X"3D",
		X"70",X"CD",X"13",X"56",X"FD",X"21",X"34",X"70",X"FE",X"01",X"CC",X"2E",X"2F",X"DD",X"21",X"88",
		X"75",X"CD",X"FE",X"13",X"FE",X"01",X"C0",X"3A",X"34",X"70",X"FE",X"01",X"C8",X"3E",X"01",X"32",
		X"34",X"70",X"E5",X"0E",X"20",X"CD",X"7D",X"21",X"E1",X"E5",X"3E",X"FE",X"CD",X"35",X"27",X"CD",
		X"F0",X"26",X"7E",X"E6",X"0F",X"F6",X"20",X"32",X"8D",X"75",X"E1",X"E5",X"CD",X"F0",X"26",X"3E",
		X"00",X"CD",X"35",X"27",X"E1",X"3E",X"32",X"32",X"8C",X"75",X"C9",X"C4",X"10",X"8C",X"98",X"C4",
		X"1A",X"9E",X"4A",X"9E",X"82",X"98",X"8B",X"86",X"00",X"B0",X"08",X"B6",X"8A",X"9C",X"12",X"9C",
		X"21",X"D1",X"72",X"06",X"24",X"AF",X"77",X"10",X"FD",X"3A",X"FD",X"70",X"01",X"09",X"00",X"21",
		X"83",X"55",X"16",X"01",X"FE",X"00",X"28",X"48",X"01",X"24",X"00",X"21",X"8C",X"55",X"16",X"04",
		X"FE",X"01",X"28",X"3C",X"01",X"24",X"00",X"21",X"B0",X"55",X"16",X"04",X"FE",X"02",X"28",X"30",
		X"01",X"09",X"00",X"21",X"D4",X"55",X"16",X"00",X"FE",X"03",X"28",X"24",X"01",X"12",X"00",X"21",
		X"DD",X"55",X"16",X"02",X"FE",X"06",X"28",X"18",X"01",X"09",X"00",X"21",X"EF",X"55",X"16",X"01",
		X"FE",X"05",X"28",X"0C",X"01",X"1B",X"00",X"21",X"F8",X"55",X"16",X"03",X"FE",X"04",X"28",X"00",
		X"7A",X"32",X"D0",X"72",X"11",X"D1",X"72",X"ED",X"B0",X"C9",X"3A",X"53",X"70",X"FE",X"01",X"28",
		X"06",X"3A",X"9E",X"72",X"FE",X"01",X"C0",X"DD",X"7E",X"04",X"FE",X"03",X"28",X"04",X"DD",X"34",
		X"04",X"C9",X"AF",X"DD",X"77",X"04",X"DD",X"66",X"00",X"DD",X"6E",X"01",X"DD",X"7E",X"02",X"47",
		X"DD",X"7E",X"03",X"80",X"DD",X"77",X"02",X"FE",X"40",X"CC",X"B3",X"20",X"FE",X"4E",X"CC",X"B7",
		X"20",X"E5",X"CD",X"C0",X"20",X"E1",X"C0",X"E5",X"23",X"CD",X"C0",X"20",X"E1",X"C0",X"E5",X"D5",
		X"11",X"20",X"00",X"19",X"D1",X"CD",X"C0",X"20",X"E1",X"C0",X"E5",X"D5",X"11",X"21",X"00",X"19",
		X"D1",X"CD",X"C0",X"20",X"E1",X"C0",X"DD",X"7E",X"02",X"77",X"3C",X"23",X"77",X"D5",X"11",X"20",
		X"00",X"19",X"D1",X"77",X"2B",X"3D",X"77",X"FE",X"44",X"D8",X"DD",X"7E",X"08",X"47",X"3A",X"83",
		X"75",X"B8",X"C0",X"3A",X"82",X"75",X"47",X"DD",X"7E",X"06",X"B8",X"D0",X"DD",X"7E",X"07",X"B8",
		X"D8",X"3E",X"01",X"3A",X"81",X"75",X"FE",X"27",X"C8",X"3E",X"01",X"32",X"13",X"70",X"AF",X"32",
		X"D6",X"72",X"C9",X"AF",X"DD",X"77",X"05",X"DD",X"7E",X"03",X"2F",X"3C",X"DD",X"77",X"03",X"C9",
		X"E5",X"7E",X"21",X"CC",X"20",X"01",X"12",X"00",X"ED",X"B1",X"E1",X"C9",X"40",X"41",X"42",X"43",
		X"44",X"45",X"46",X"47",X"48",X"49",X"4A",X"4B",X"4C",X"4D",X"4E",X"4F",X"FF",X"FE",X"3A",X"FD",
		X"70",X"FE",X"00",X"C0",X"3A",X"6B",X"70",X"08",X"3A",X"9B",X"70",X"32",X"6B",X"70",X"08",X"32",
		X"9B",X"70",X"C9",X"DD",X"E5",X"DD",X"21",X"EB",X"70",X"06",X"09",X"DD",X"7E",X"00",X"FE",X"FF",
		X"28",X"09",X"DD",X"23",X"DD",X"23",X"10",X"F3",X"DD",X"E1",X"C9",X"DD",X"75",X"00",X"DD",X"74",
		X"01",X"AF",X"32",X"63",X"70",X"32",X"C3",X"72",X"DD",X"E1",X"C9",X"06",X"04",X"DD",X"21",X"88",
		X"75",X"DD",X"7E",X"00",X"DD",X"77",X"10",X"DD",X"23",X"10",X"F6",X"3E",X"20",X"32",X"85",X"72",
		X"3E",X"80",X"32",X"86",X"72",X"3E",X"3F",X"32",X"98",X"75",X"C9",X"AF",X"32",X"85",X"72",X"32",
		X"88",X"72",X"32",X"9A",X"75",X"32",X"9B",X"75",X"C9",X"D5",X"DD",X"E5",X"06",X"09",X"DD",X"21",
		X"EB",X"70",X"DD",X"5E",X"00",X"DD",X"56",X"01",X"E5",X"AF",X"ED",X"52",X"E1",X"28",X"0A",X"DD",
		X"23",X"DD",X"23",X"10",X"ED",X"DD",X"E1",X"D1",X"C9",X"3E",X"FF",X"DD",X"77",X"00",X"DD",X"77",
		X"01",X"3E",X"01",X"32",X"63",X"70",X"32",X"C3",X"72",X"DD",X"E1",X"D1",X"C9",X"CD",X"6D",X"15",
		X"FD",X"21",X"69",X"70",X"FD",X"5E",X"00",X"FD",X"56",X"01",X"E5",X"EB",X"CD",X"9D",X"2F",X"CD",
		X"A2",X"2F",X"AF",X"ED",X"52",X"E1",X"28",X"09",X"FD",X"23",X"FD",X"23",X"FD",X"23",X"10",X"E4",
		X"C9",X"FD",X"7E",X"02",X"B1",X"FD",X"77",X"02",X"AF",X"FD",X"77",X"00",X"FD",X"77",X"01",X"C9",
		X"11",X"E2",X"70",X"DD",X"21",X"EB",X"70",X"06",X"09",X"0E",X"A4",X"1A",X"FE",X"B0",X"38",X"3E",
		X"0E",X"A0",X"FE",X"C0",X"38",X"38",X"0E",X"9C",X"FE",X"D0",X"38",X"32",X"DD",X"7E",X"00",X"FE",
		X"FF",X"28",X"46",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"CD",X"21",X"22",X"20",X"13",X"3E",X"FF",
		X"CD",X"35",X"27",X"3E",X"00",X"CD",X"29",X"22",X"3E",X"00",X"DD",X"77",X"00",X"DD",X"77",X"01",
		X"12",X"D5",X"DD",X"E5",X"C5",X"CD",X"9E",X"16",X"C1",X"DD",X"E1",X"D1",X"18",X"1B",X"DD",X"6E",
		X"00",X"DD",X"66",X"01",X"CD",X"21",X"22",X"20",X"10",X"79",X"D5",X"CD",X"4D",X"27",X"E5",X"CD",
		X"F0",X"26",X"3E",X"20",X"CD",X"35",X"27",X"E1",X"D1",X"13",X"DD",X"23",X"DD",X"23",X"10",X"99",
		X"C9",X"E5",X"D5",X"CD",X"6B",X"2F",X"D1",X"E1",X"C9",X"E5",X"F5",X"CD",X"F0",X"26",X"F1",X"CD",
		X"35",X"27",X"E1",X"C9",X"3A",X"C3",X"72",X"FE",X"30",X"D8",X"3E",X"01",X"32",X"5B",X"70",X"C9",
		X"3A",X"62",X"70",X"47",X"3A",X"A6",X"72",X"80",X"47",X"3A",X"63",X"70",X"80",X"06",X"2C",X"21",
		X"81",X"75",X"FE",X"00",X"28",X"02",X"06",X"27",X"70",X"C9",X"AF",X"32",X"43",X"70",X"32",X"5B",
		X"70",X"32",X"34",X"70",X"32",X"BD",X"72",X"32",X"BE",X"72",X"32",X"BF",X"72",X"32",X"C0",X"72",
		X"32",X"62",X"70",X"32",X"63",X"70",X"32",X"BD",X"72",X"32",X"BE",X"72",X"32",X"BF",X"72",X"32",
		X"C0",X"72",X"32",X"8E",X"75",X"32",X"8F",X"75",X"32",X"9E",X"75",X"32",X"9F",X"75",X"C9",X"3E",
		X"00",X"CD",X"68",X"19",X"21",X"A0",X"8B",X"11",X"5A",X"57",X"CD",X"49",X"19",X"3E",X"0A",X"21",
		X"C0",X"9A",X"06",X"08",X"CD",X"60",X"19",X"21",X"20",X"89",X"11",X"63",X"57",X"CD",X"49",X"19",
		X"3E",X"0A",X"21",X"40",X"98",X"06",X"08",X"CD",X"60",X"19",X"21",X"40",X"8A",X"11",X"A4",X"57",
		X"CD",X"49",X"19",X"3E",X"0A",X"21",X"A0",X"99",X"06",X"07",X"CD",X"60",X"19",X"21",X"7F",X"89",
		X"11",X"89",X"56",X"CD",X"54",X"23",X"3E",X"04",X"21",X"7F",X"98",X"06",X"09",X"CD",X"60",X"19",
		X"C9",X"11",X"C3",X"56",X"21",X"AF",X"8B",X"CD",X"49",X"19",X"3E",X"0E",X"21",X"4F",X"98",X"06",
		X"1C",X"CD",X"60",X"19",X"11",X"DF",X"56",X"21",X"11",X"8B",X"CD",X"49",X"19",X"3E",X"0E",X"21",
		X"51",X"98",X"06",X"1C",X"CD",X"60",X"19",X"C9",X"11",X"F2",X"56",X"21",X"11",X"8B",X"CD",X"49",
		X"19",X"3E",X"0E",X"21",X"51",X"98",X"06",X"1C",X"CD",X"60",X"19",X"C9",X"3E",X"0A",X"32",X"7E",
		X"72",X"21",X"D2",X"36",X"22",X"74",X"72",X"21",X"D2",X"36",X"22",X"77",X"72",X"21",X"D2",X"36",
		X"22",X"7A",X"72",X"AF",X"32",X"76",X"72",X"32",X"79",X"72",X"32",X"7C",X"72",X"C9",X"21",X"69",
		X"33",X"CD",X"89",X"0B",X"21",X"00",X"30",X"CD",X"A3",X"0B",X"3E",X"01",X"32",X"7F",X"72",X"AF",
		X"32",X"A2",X"72",X"C9",X"01",X"E0",X"FF",X"1A",X"FE",X"3F",X"C8",X"D6",X"30",X"77",X"E5",X"7C",
		X"C6",X"10",X"67",X"3E",X"03",X"77",X"E1",X"13",X"09",X"18",X"E9",X"01",X"E0",X"FF",X"1A",X"FE",
		X"3F",X"C8",X"77",X"E5",X"7C",X"C6",X"10",X"67",X"08",X"77",X"08",X"E1",X"13",X"09",X"18",X"EB",
		X"11",X"20",X"00",X"06",X"1C",X"77",X"19",X"10",X"FC",X"C9",X"DD",X"7E",X"00",X"FE",X"00",X"C8",
		X"DD",X"7E",X"02",X"FE",X"00",X"C0",X"AF",X"DD",X"77",X"00",X"3E",X"01",X"DD",X"77",X"02",X"E5",
		X"21",X"00",X"10",X"CD",X"6A",X"27",X"E1",X"3E",X"29",X"32",X"94",X"75",X"3E",X"2A",X"32",X"95",
		X"75",X"AF",X"32",X"86",X"75",X"32",X"87",X"75",X"32",X"20",X"70",X"3E",X"FF",X"32",X"A6",X"72",
		X"21",X"00",X"00",X"CD",X"F3",X"20",X"C9",X"CD",X"EF",X"23",X"38",X"11",X"AF",X"DD",X"77",X"00",
		X"DD",X"77",X"02",X"32",X"96",X"75",X"32",X"97",X"75",X"3E",X"10",X"12",X"C9",X"FE",X"00",X"C8",
		X"AF",X"12",X"FD",X"7E",X"02",X"32",X"96",X"75",X"FD",X"7E",X"03",X"32",X"97",X"75",X"C9",X"21",
		X"81",X"53",X"3A",X"FD",X"70",X"85",X"3E",X"00",X"8C",X"DD",X"7E",X"02",X"BE",X"C9",X"3A",X"20",
		X"CD",X"B2",X"2F",X"22",X"B1",X"72",X"CD",X"5A",X"24",X"20",X"03",X"22",X"A9",X"72",X"CD",X"C3",
		X"2F",X"22",X"B1",X"72",X"CD",X"5A",X"24",X"20",X"03",X"22",X"AB",X"72",X"3A",X"20",X"70",X"C5",
		X"47",X"3A",X"34",X"70",X"80",X"C1",X"FE",X"02",X"20",X"21",X"DD",X"21",X"7D",X"24",X"06",X"09",
		X"C5",X"2A",X"A9",X"72",X"DD",X"56",X"01",X"DD",X"5E",X"00",X"19",X"ED",X"5B",X"AB",X"72",X"AF",
		X"ED",X"52",X"28",X"14",X"DD",X"23",X"DD",X"23",X"C1",X"10",X"E5",X"2A",X"A9",X"72",X"22",X"AD",
		X"72",X"2A",X"AB",X"72",X"22",X"AF",X"72",X"C9",X"C1",X"C9",X"DD",X"21",X"7D",X"24",X"06",X"09",
		X"C5",X"2A",X"B1",X"72",X"DD",X"56",X"01",X"DD",X"5E",X"00",X"19",X"E5",X"CD",X"75",X"2F",X"E1",
		X"DD",X"23",X"DD",X"23",X"C1",X"C8",X"10",X"E8",X"3E",X"01",X"FE",X"02",X"C9",X"00",X"00",X"FF",
		X"FF",X"01",X"00",X"E1",X"FF",X"E0",X"FF",X"DF",X"FF",X"1F",X"00",X"20",X"00",X"21",X"00",X"3E",
		X"01",X"32",X"94",X"72",X"3E",X"00",X"32",X"42",X"70",X"32",X"5D",X"70",X"32",X"13",X"70",X"32",
		X"8D",X"72",X"32",X"35",X"70",X"32",X"49",X"70",X"32",X"4A",X"70",X"32",X"4B",X"70",X"32",X"4C",
		X"70",X"32",X"85",X"72",X"32",X"22",X"70",X"CD",X"5A",X"22",X"3A",X"02",X"70",X"06",X"10",X"B0",
		X"32",X"02",X"70",X"11",X"80",X"75",X"21",X"CE",X"2F",X"01",X"1C",X"00",X"ED",X"B0",X"3A",X"82",
		X"75",X"FE",X"40",X"38",X"F9",X"CD",X"85",X"26",X"11",X"DC",X"58",X"21",X"76",X"8A",X"CD",X"54",
		X"23",X"21",X"16",X"99",X"3E",X"0D",X"06",X"0C",X"CD",X"60",X"19",X"3A",X"02",X"70",X"E6",X"07",
		X"32",X"02",X"70",X"3E",X"01",X"32",X"49",X"70",X"32",X"4A",X"70",X"3E",X"00",X"32",X"4B",X"70",
		X"3A",X"92",X"75",X"FE",X"20",X"38",X"F9",X"3E",X"01",X"32",X"4C",X"70",X"3A",X"92",X"75",X"FE",
		X"40",X"38",X"F9",X"CD",X"85",X"26",X"11",X"E5",X"58",X"21",X"78",X"8A",X"CD",X"54",X"23",X"21",
		X"18",X"99",X"06",X"0C",X"3E",X"0D",X"CD",X"60",X"19",X"3E",X"00",X"32",X"49",X"70",X"32",X"4A",
		X"70",X"3E",X"10",X"32",X"35",X"70",X"3E",X"00",X"32",X"86",X"72",X"3A",X"8A",X"75",X"FE",X"40",
		X"38",X"F9",X"CD",X"85",X"26",X"11",X"F2",X"58",X"21",X"7A",X"8A",X"CD",X"54",X"23",X"21",X"1A",
		X"99",X"06",X"0C",X"3E",X"0D",X"CD",X"60",X"19",X"3E",X"00",X"32",X"35",X"70",X"3E",X"10",X"32",
		X"85",X"72",X"3A",X"9A",X"75",X"FE",X"40",X"38",X"F9",X"CD",X"85",X"26",X"11",X"FE",X"58",X"21",
		X"7C",X"8A",X"CD",X"54",X"23",X"21",X"1C",X"99",X"06",X"0C",X"3E",X"0D",X"CD",X"60",X"19",X"3E",
		X"00",X"32",X"85",X"72",X"06",X"01",X"21",X"00",X"90",X"2B",X"E5",X"C5",X"3E",X"B9",X"CD",X"AA",
		X"06",X"C1",X"E1",X"7C",X"FE",X"00",X"20",X"F1",X"CD",X"85",X"26",X"10",X"E9",X"3E",X"01",X"32",
		X"9E",X"72",X"CD",X"B2",X"25",X"AF",X"32",X"9E",X"72",X"3A",X"02",X"70",X"E6",X"07",X"32",X"02",
		X"70",X"C9",X"AF",X"32",X"03",X"A0",X"AF",X"32",X"FD",X"70",X"CD",X"B5",X"19",X"11",X"80",X"75",
		X"21",X"3A",X"55",X"01",X"1C",X"00",X"ED",X"B0",X"CD",X"B0",X"1F",X"CD",X"D4",X"11",X"3E",X"01",
		X"32",X"03",X"A0",X"CD",X"9C",X"27",X"AF",X"32",X"94",X"72",X"CD",X"28",X"16",X"3E",X"10",X"32",
		X"35",X"70",X"3E",X"03",X"32",X"49",X"70",X"3E",X"03",X"32",X"36",X"70",X"3E",X"10",X"32",X"02",
		X"70",X"3E",X"20",X"32",X"36",X"70",X"32",X"22",X"70",X"CD",X"00",X"24",X"CD",X"40",X"22",X"CD",
		X"28",X"1F",X"3A",X"24",X"70",X"FE",X"01",X"20",X"0F",X"CD",X"56",X"26",X"3E",X"00",X"32",X"24",
		X"70",X"3E",X"01",X"32",X"9C",X"72",X"18",X"12",X"DD",X"21",X"80",X"75",X"21",X"9C",X"72",X"FD",
		X"21",X"95",X"72",X"CD",X"13",X"56",X"FE",X"01",X"20",X"00",X"CD",X"85",X"26",X"3A",X"13",X"70",
		X"FE",X"01",X"28",X"06",X"CD",X"B0",X"21",X"18",X"C0",X"C9",X"CD",X"49",X"1B",X"3A",X"F6",X"72",
		X"3C",X"FE",X"03",X"06",X"04",X"28",X"07",X"06",X"00",X"FE",X"07",X"28",X"01",X"47",X"78",X"32",
		X"F6",X"72",X"32",X"FD",X"70",X"C9",X"CD",X"FB",X"2E",X"E6",X"03",X"3C",X"47",X"21",X"7A",X"55",
		X"23",X"10",X"FD",X"3A",X"00",X"B8",X"3A",X"02",X"70",X"E6",X"F8",X"32",X"9D",X"72",X"47",X"E5",
		X"23",X"23",X"23",X"23",X"7E",X"E1",X"B8",X"28",X"DD",X"7E",X"47",X"3A",X"02",X"70",X"E6",X"07",
		X"B0",X"32",X"02",X"70",X"C9",X"3A",X"00",X"70",X"FE",X"00",X"C8",X"F1",X"C9",X"F5",X"DD",X"E5",
		X"D5",X"C5",X"E5",X"7D",X"E6",X"1F",X"6F",X"AF",X"26",X"00",X"CD",X"D5",X"26",X"4F",X"E1",X"E5",
		X"11",X"20",X"00",X"7D",X"E6",X"E0",X"CB",X"1C",X"CB",X"1D",X"CB",X"1C",X"CB",X"1D",X"CB",X"1C",
		X"CB",X"1D",X"CB",X"1C",X"CB",X"1D",X"CB",X"1C",X"CB",X"1D",X"7D",X"E6",X"1F",X"6F",X"AF",X"67",
		X"CD",X"E2",X"26",X"47",X"DD",X"21",X"80",X"75",X"DD",X"71",X"03",X"DD",X"70",X"02",X"E1",X"C1",
		X"D1",X"DD",X"E1",X"F1",X"C9",X"06",X"08",X"7D",X"FE",X"00",X"C8",X"AF",X"5D",X"80",X"1D",X"C8",
		X"18",X"FB",X"06",X"08",X"7D",X"FE",X"00",X"C8",X"3E",X"F0",X"5D",X"90",X"1D",X"C8",X"18",X"FB",
		X"7C",X"C6",X"10",X"67",X"C9",X"7C",X"E6",X"60",X"FE",X"60",X"28",X"07",X"7C",X"3D",X"E6",X"60",
		X"FE",X"60",X"C0",X"F1",X"C9",X"CD",X"F5",X"26",X"3E",X"C8",X"77",X"3E",X"C9",X"E5",X"23",X"77",
		X"11",X"20",X"00",X"19",X"3E",X"CB",X"77",X"2B",X"3E",X"CA",X"77",X"E1",X"C9",X"CD",X"F5",X"26",
		X"3E",X"A4",X"77",X"3E",X"A5",X"E5",X"23",X"77",X"11",X"20",X"00",X"19",X"3E",X"A7",X"77",X"2B",
		X"3E",X"A6",X"77",X"E1",X"C9",X"E5",X"08",X"7C",X"E6",X"80",X"FE",X"80",X"20",X"0D",X"08",X"77",
		X"23",X"77",X"D5",X"11",X"20",X"00",X"19",X"D1",X"77",X"2B",X"77",X"E1",X"C9",X"E5",X"F5",X"7C",
		X"E6",X"80",X"FE",X"80",X"20",X"11",X"F1",X"F5",X"77",X"23",X"3C",X"77",X"D5",X"11",X"1F",X"00",
		X"19",X"D1",X"3C",X"77",X"23",X"3C",X"77",X"F1",X"E1",X"C9",X"3A",X"0B",X"70",X"FE",X"00",X"C2",
		X"95",X"27",X"DD",X"21",X"26",X"70",X"AF",X"7D",X"47",X"DD",X"7E",X"00",X"80",X"27",X"DD",X"77",
		X"00",X"7C",X"47",X"DD",X"7E",X"01",X"88",X"27",X"DD",X"77",X"01",X"DD",X"7E",X"02",X"CE",X"00",
		X"27",X"DD",X"77",X"02",X"C9",X"DD",X"21",X"29",X"70",X"C3",X"76",X"27",X"DD",X"21",X"26",X"70",
		X"21",X"E1",X"8A",X"CD",X"F3",X"27",X"DD",X"21",X"29",X"70",X"21",X"61",X"88",X"CD",X"F3",X"27",
		X"21",X"9F",X"8B",X"11",X"E0",X"FF",X"3A",X"D5",X"70",X"FE",X"00",X"28",X"11",X"08",X"3E",X"67",
		X"77",X"E5",X"CD",X"F0",X"26",X"3E",X"0C",X"77",X"E1",X"19",X"08",X"3D",X"18",X"EB",X"3E",X"FF",
		X"77",X"DD",X"21",X"F7",X"71",X"21",X"01",X"8A",X"06",X"01",X"CD",X"F5",X"27",X"AF",X"32",X"C1",
		X"89",X"32",X"E1",X"89",X"3E",X"FF",X"32",X"41",X"8A",X"3A",X"FD",X"71",X"FE",X"00",X"C8",X"32",
		X"41",X"8A",X"C9",X"06",X"03",X"11",X"20",X"00",X"DD",X"7E",X"00",X"CD",X"04",X"28",X"DD",X"23",
		X"19",X"10",X"F5",X"C9",X"F5",X"E6",X"0F",X"77",X"19",X"F1",X"CB",X"0F",X"CB",X"0F",X"CB",X"0F",
		X"CB",X"0F",X"E6",X"0F",X"77",X"C9",X"DD",X"21",X"69",X"70",X"FD",X"21",X"03",X"71",X"06",X"33",
		X"DD",X"7E",X"00",X"08",X"FD",X"7E",X"00",X"DD",X"77",X"00",X"08",X"FD",X"77",X"00",X"DD",X"7E",
		X"01",X"08",X"FD",X"7E",X"01",X"DD",X"77",X"01",X"08",X"FD",X"77",X"01",X"DD",X"7E",X"02",X"08",
		X"FD",X"7E",X"02",X"DD",X"77",X"02",X"08",X"FD",X"77",X"02",X"DD",X"23",X"DD",X"23",X"DD",X"23",
		X"FD",X"23",X"FD",X"23",X"FD",X"23",X"10",X"C8",X"3A",X"0B",X"70",X"2F",X"E6",X"01",X"32",X"0B",
		X"70",X"06",X"00",X"3A",X"00",X"A8",X"E6",X"80",X"FE",X"80",X"28",X"02",X"06",X"01",X"3A",X"0B",
		X"70",X"A0",X"2F",X"32",X"01",X"A0",X"32",X"02",X"A0",X"C9",X"AF",X"32",X"05",X"A0",X"3E",X"07",
		X"D3",X"08",X"3E",X"38",X"D3",X"09",X"3E",X"0E",X"D3",X"08",X"DB",X"0C",X"2F",X"32",X"F2",X"71",
		X"3E",X"01",X"32",X"05",X"A0",X"C9",X"AF",X"32",X"05",X"A0",X"3E",X"07",X"D3",X"08",X"3E",X"38",
		X"D3",X"09",X"3E",X"0F",X"D3",X"08",X"DB",X"0C",X"2F",X"32",X"F2",X"71",X"3E",X"01",X"32",X"05",
		X"A0",X"C9",X"CD",X"FB",X"2E",X"E6",X"3F",X"47",X"00",X"10",X"FD",X"3E",X"80",X"32",X"36",X"70",
		X"3A",X"FE",X"70",X"FE",X"01",X"20",X"05",X"3E",X"08",X"32",X"36",X"70",X"3A",X"00",X"A8",X"E6",
		X"20",X"FE",X"20",X"3E",X"03",X"28",X"02",X"3E",X"04",X"47",X"3A",X"0B",X"70",X"FE",X"01",X"3A",
		X"28",X"70",X"20",X"03",X"3A",X"2B",X"70",X"B8",X"30",X"05",X"AF",X"32",X"FF",X"70",X"C9",X"3A",
		X"FF",X"70",X"FE",X"00",X"C0",X"3A",X"D5",X"70",X"3C",X"32",X"D5",X"70",X"3E",X"01",X"32",X"FF",
		X"70",X"21",X"6B",X"37",X"CD",X"CF",X"0B",X"C9",X"AF",X"32",X"53",X"70",X"FD",X"21",X"26",X"70",
		X"CD",X"10",X"2A",X"78",X"FE",X"05",X"38",X"0B",X"FD",X"21",X"29",X"70",X"CD",X"10",X"2A",X"78",
		X"FE",X"05",X"D0",X"CD",X"6D",X"2C",X"21",X"83",X"8B",X"01",X"0C",X"18",X"3E",X"03",X"08",X"CD",
		X"A3",X"1A",X"21",X"91",X"8B",X"01",X"0C",X"18",X"3E",X"00",X"08",X"CD",X"A3",X"1A",X"CD",X"4A",
		X"2D",X"CD",X"24",X"2C",X"3A",X"0B",X"70",X"FE",X"01",X"CC",X"16",X"28",X"CD",X"B6",X"2B",X"3E",
		X"01",X"32",X"01",X"A0",X"32",X"02",X"A0",X"FD",X"21",X"26",X"70",X"CD",X"10",X"2A",X"78",X"FE",
		X"05",X"D2",X"97",X"29",X"DD",X"23",X"DD",X"23",X"DD",X"23",X"D5",X"11",X"F0",X"FF",X"DD",X"19",
		X"D1",X"DD",X"E5",X"23",X"23",X"E5",X"CD",X"3C",X"2A",X"3E",X"60",X"32",X"F7",X"71",X"AF",X"32",
		X"FD",X"71",X"E1",X"CD",X"B6",X"2B",X"DD",X"E1",X"3E",X"01",X"32",X"F4",X"71",X"AF",X"32",X"FA",
		X"71",X"CD",X"90",X"2A",X"CD",X"B6",X"2B",X"3A",X"0C",X"70",X"FE",X"01",X"28",X"62",X"3A",X"00",
		X"A8",X"E6",X"80",X"FE",X"80",X"28",X"08",X"3E",X"00",X"32",X"01",X"A0",X"32",X"02",X"A0",X"3A",
		X"02",X"70",X"E6",X"80",X"FE",X"80",X"28",X"F7",X"FD",X"21",X"29",X"70",X"CD",X"10",X"2A",X"78",
		X"FE",X"05",X"30",X"3C",X"CD",X"B6",X"2B",X"DD",X"23",X"DD",X"23",X"DD",X"23",X"D5",X"11",X"F0",
		X"FF",X"DD",X"19",X"D1",X"DD",X"E5",X"23",X"23",X"E5",X"CD",X"3C",X"2A",X"3E",X"60",X"32",X"F7",
		X"71",X"AF",X"32",X"FD",X"71",X"E1",X"CD",X"B6",X"2B",X"DD",X"E1",X"3E",X"00",X"32",X"4A",X"70",
		X"32",X"F4",X"71",X"CD",X"62",X"2B",X"CD",X"62",X"2B",X"CD",X"62",X"2B",X"CD",X"90",X"2A",X"C9",
		X"AF",X"32",X"67",X"72",X"3E",X"01",X"32",X"01",X"A0",X"32",X"02",X"A0",X"32",X"FA",X"71",X"C9",
		X"DD",X"21",X"9A",X"71",X"11",X"10",X"00",X"21",X"0F",X"8A",X"06",X"05",X"FD",X"7E",X"02",X"DD",
		X"BE",X"02",X"D8",X"20",X"10",X"FD",X"7E",X"01",X"DD",X"BE",X"01",X"D8",X"20",X"07",X"FD",X"7E",
		X"00",X"DD",X"BE",X"00",X"D8",X"DD",X"19",X"2B",X"2B",X"10",X"E1",X"C9",X"C5",X"DD",X"21",X"9A",
		X"71",X"78",X"FE",X"04",X"30",X"11",X"C5",X"06",X"10",X"DD",X"7E",X"10",X"DD",X"77",X"00",X"DD",
		X"23",X"10",X"F6",X"C1",X"04",X"18",X"EA",X"C1",X"DD",X"21",X"9A",X"71",X"78",X"FE",X"04",X"30",
		X"05",X"DD",X"19",X"04",X"18",X"F6",X"FD",X"7E",X"00",X"DD",X"77",X"00",X"FD",X"7E",X"01",X"DD",
		X"77",X"01",X"FD",X"7E",X"02",X"DD",X"77",X"02",X"C5",X"06",X"0D",X"DD",X"E5",X"DD",X"23",X"DD",
		X"23",X"DD",X"23",X"3E",X"10",X"DD",X"77",X"00",X"DD",X"23",X"10",X"F9",X"DD",X"E1",X"C1",X"C9",
		X"06",X"11",X"3E",X"00",X"32",X"F2",X"71",X"F3",X"3A",X"F4",X"71",X"FE",X"01",X"20",X"05",X"CD",
		X"7A",X"28",X"18",X"0C",X"3A",X"00",X"A8",X"E6",X"80",X"FE",X"80",X"28",X"F2",X"CD",X"96",X"28",
		X"FB",X"3A",X"F2",X"71",X"E6",X"10",X"FE",X"10",X"CC",X"FB",X"2A",X"3A",X"F2",X"71",X"E6",X"08",
		X"FE",X"08",X"CC",X"0A",X"2B",X"3A",X"F2",X"71",X"E6",X"40",X"FE",X"40",X"CC",X"19",X"2B",X"3A",
		X"F2",X"71",X"E6",X"20",X"FE",X"20",X"CC",X"37",X"2B",X"3A",X"F2",X"71",X"E6",X"80",X"FE",X"80",
		X"C8",X"3A",X"F7",X"71",X"FE",X"00",X"C8",X"CD",X"53",X"2B",X"DD",X"E5",X"E5",X"F5",X"C5",X"D5",
		X"CD",X"9C",X"27",X"D1",X"C1",X"F1",X"E1",X"DD",X"E1",X"18",X"9C",X"78",X"FE",X"2B",X"20",X"02",
		X"06",X"10",X"04",X"CD",X"53",X"2B",X"CD",X"62",X"2B",X"C9",X"78",X"FE",X"10",X"20",X"02",X"06",
		X"2C",X"05",X"CD",X"53",X"2B",X"CD",X"62",X"2B",X"C9",X"7D",X"E6",X"F0",X"FE",X"00",X"20",X"04",
		X"7C",X"FE",X"8A",X"C8",X"06",X"10",X"CD",X"53",X"2B",X"11",X"20",X"00",X"19",X"DD",X"2B",X"46",
		X"CD",X"53",X"2B",X"CD",X"62",X"2B",X"C9",X"7D",X"E6",X"F0",X"FE",X"C0",X"20",X"04",X"7C",X"FE",
		X"89",X"C8",X"11",X"20",X"00",X"AF",X"ED",X"52",X"DD",X"23",X"06",X"11",X"CD",X"53",X"2B",X"CD",
		X"62",X"2B",X"C9",X"78",X"DD",X"77",X"00",X"77",X"E5",X"7C",X"C6",X"10",X"67",X"3E",X"01",X"77",
		X"E1",X"C9",X"C5",X"F5",X"E5",X"06",X"70",X"21",X"00",X"03",X"2B",X"7C",X"FE",X"00",X"20",X"FA",
		X"10",X"F5",X"E1",X"F1",X"C1",X"C9",X"21",X"25",X"8B",X"11",X"4F",X"57",X"CD",X"49",X"19",X"21",
		X"05",X"8A",X"11",X"55",X"57",X"CD",X"49",X"19",X"21",X"85",X"99",X"3E",X"07",X"06",X"0E",X"CD",
		X"60",X"19",X"21",X"E3",X"8A",X"11",X"90",X"56",X"CD",X"49",X"19",X"21",X"03",X"99",X"3E",X"03",
		X"06",X"10",X"CD",X"60",X"19",X"C9",X"77",X"E5",X"F5",X"7C",X"C6",X"10",X"67",X"3E",X"10",X"77",
		X"F1",X"E1",X"23",X"10",X"F1",X"C9",X"DD",X"E5",X"C5",X"E5",X"D5",X"CD",X"76",X"2B",X"11",X"20",
		X"00",X"21",X"8F",X"8A",X"DD",X"21",X"9A",X"71",X"06",X"05",X"C5",X"E5",X"06",X"03",X"DD",X"7E",
		X"00",X"E6",X"0F",X"CD",X"57",X"2B",X"DD",X"7E",X"00",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"11",
		X"20",X"00",X"19",X"CD",X"57",X"2B",X"DD",X"23",X"19",X"10",X"E3",X"E1",X"2B",X"2B",X"C1",X"11",
		X"0D",X"00",X"DD",X"19",X"10",X"D4",X"11",X"20",X"00",X"DD",X"21",X"9A",X"71",X"21",X"0F",X"8A",
		X"06",X"05",X"C5",X"E5",X"DD",X"23",X"DD",X"23",X"DD",X"23",X"06",X"0D",X"DD",X"7E",X"00",X"CD",
		X"57",X"2B",X"DD",X"23",X"ED",X"52",X"10",X"F4",X"E1",X"2B",X"2B",X"C1",X"10",X"E4",X"D1",X"E1",
		X"C1",X"DD",X"E1",X"C9",X"3E",X"01",X"32",X"67",X"72",X"21",X"72",X"8B",X"11",X"1E",X"57",X"CD",
		X"49",X"19",X"21",X"73",X"8B",X"11",X"37",X"57",X"CD",X"49",X"19",X"21",X"7D",X"8B",X"11",X"75",
		X"57",X"CD",X"49",X"19",X"CD",X"76",X"2B",X"C9",X"3E",X"14",X"08",X"CD",X"6B",X"23",X"C9",X"3E",
		X"18",X"08",X"CD",X"59",X"2C",X"CD",X"6B",X"23",X"C9",X"F5",X"3A",X"00",X"A8",X"E6",X"40",X"FE",
		X"40",X"20",X"08",X"E5",X"EB",X"11",X"0A",X"00",X"19",X"EB",X"E1",X"F1",X"C9",X"3E",X"00",X"32",
		X"03",X"A0",X"CD",X"B5",X"19",X"3E",X"07",X"CD",X"68",X"19",X"21",X"41",X"98",X"3E",X"05",X"06",
		X"1E",X"CD",X"60",X"19",X"21",X"40",X"98",X"3E",X"02",X"06",X"1E",X"CD",X"60",X"19",X"21",X"7F",
		X"98",X"3E",X"04",X"06",X"0A",X"CD",X"60",X"19",X"3E",X"01",X"32",X"03",X"A0",X"C9",X"CD",X"6D",
		X"2C",X"AF",X"32",X"03",X"A0",X"21",X"83",X"8B",X"01",X"0D",X"18",X"3E",X"03",X"08",X"CD",X"A3",
		X"1A",X"11",X"AC",X"56",X"21",X"5A",X"8B",X"CD",X"49",X"19",X"11",X"00",X"50",X"21",X"B5",X"8B",
		X"CD",X"54",X"23",X"3E",X"0E",X"21",X"9A",X"98",X"CD",X"80",X"23",X"11",X"A2",X"0E",X"21",X"57",
		X"8B",X"CD",X"54",X"23",X"11",X"A3",X"0E",X"21",X"18",X"8B",X"CD",X"54",X"23",X"3E",X"00",X"21",
		X"57",X"98",X"CD",X"80",X"23",X"3E",X"00",X"21",X"58",X"98",X"CD",X"80",X"23",X"3E",X"03",X"21",
		X"55",X"98",X"CD",X"80",X"23",X"CD",X"B6",X"2B",X"3E",X"01",X"32",X"00",X"A0",X"32",X"42",X"70",
		X"3E",X"0A",X"21",X"40",X"98",X"06",X"1E",X"CD",X"60",X"19",X"3A",X"42",X"70",X"FE",X"00",X"28",
		X"0E",X"3A",X"00",X"70",X"FE",X"00",X"C0",X"3E",X"01",X"32",X"03",X"A0",X"C3",X"0A",X"2D",X"3E",
		X"01",X"32",X"42",X"70",X"3A",X"00",X"70",X"FE",X"00",X"C0",X"3A",X"42",X"70",X"FE",X"FF",X"C8",
		X"18",X"F2",X"3A",X"02",X"70",X"E6",X"80",X"FE",X"80",X"C0",X"3A",X"03",X"70",X"E6",X"80",X"FE",
		X"00",X"C0",X"F5",X"3E",X"01",X"32",X"BC",X"72",X"F1",X"C9",X"21",X"16",X"8A",X"36",X"80",X"23",
		X"36",X"7F",X"23",X"23",X"36",X"7F",X"23",X"36",X"79",X"3E",X"02",X"21",X"16",X"9A",X"77",X"23",
		X"77",X"23",X"23",X"77",X"23",X"77",X"21",X"17",X"9A",X"36",X"0A",X"21",X"19",X"9A",X"36",X"0A",
		X"21",X"75",X"8A",X"11",X"B9",X"57",X"CD",X"49",X"19",X"21",X"F8",X"8A",X"11",X"C1",X"57",X"CD",
		X"49",X"19",X"21",X"9B",X"8A",X"11",X"D3",X"57",X"CD",X"49",X"19",X"21",X"38",X"9A",X"36",X"0A",
		X"21",X"F8",X"99",X"36",X"0A",X"21",X"95",X"99",X"3E",X"02",X"06",X"08",X"CD",X"60",X"19",X"21",
		X"78",X"9A",X"06",X"05",X"CD",X"60",X"19",X"21",X"F8",X"98",X"06",X"07",X"CD",X"60",X"19",X"21",
		X"BB",X"99",X"06",X"09",X"CD",X"60",X"19",X"C9",X"3E",X"01",X"32",X"8D",X"72",X"AF",X"32",X"62",
		X"70",X"CD",X"3D",X"1B",X"21",X"3A",X"55",X"11",X"80",X"75",X"01",X"04",X"00",X"ED",X"B0",X"3E",
		X"58",X"32",X"82",X"75",X"3E",X"C0",X"32",X"83",X"75",X"21",X"73",X"8A",X"11",X"69",X"52",X"3E",
		X"03",X"08",X"CD",X"6B",X"23",X"21",X"B7",X"8A",X"11",X"72",X"52",X"3E",X"03",X"08",X"CD",X"6B",
		X"23",X"21",X"BA",X"8A",X"11",X"7F",X"52",X"3E",X"03",X"08",X"CD",X"6B",X"23",X"3E",X"03",X"08",
		X"06",X"03",X"21",X"74",X"8A",X"CD",X"6C",X"2E",X"06",X"02",X"21",X"B8",X"8A",X"CD",X"6C",X"2E",
		X"21",X"94",X"89",X"06",X"03",X"CD",X"6C",X"2E",X"21",X"58",X"89",X"06",X"02",X"CD",X"6C",X"2E",
		X"21",X"A4",X"8B",X"01",X"0C",X"1A",X"3E",X"00",X"08",X"CD",X"A3",X"1A",X"06",X"09",X"DD",X"21",
		X"1D",X"5C",X"11",X"14",X"5C",X"C5",X"DD",X"66",X"01",X"DD",X"6E",X"00",X"D5",X"11",X"0B",X"00",
		X"ED",X"52",X"D1",X"CD",X"AD",X"2E",X"DD",X"23",X"DD",X"23",X"DD",X"23",X"13",X"C1",X"10",X"E5",
		X"21",X"85",X"8B",X"11",X"E0",X"57",X"CD",X"49",X"19",X"21",X"A6",X"8A",X"11",X"FB",X"57",X"CD",
		X"49",X"19",X"21",X"47",X"8B",X"11",X"06",X"58",X"CD",X"49",X"19",X"C9",X"3E",X"F8",X"CD",X"E5",
		X"1A",X"23",X"10",X"F8",X"C9",X"11",X"14",X"5C",X"06",X"09",X"C5",X"DD",X"21",X"1D",X"5C",X"CD",
		X"FB",X"2E",X"E6",X"0F",X"FE",X"09",X"30",X"F3",X"FE",X"00",X"28",X"0A",X"D5",X"11",X"03",X"00",
		X"47",X"DD",X"19",X"10",X"FC",X"D1",X"DD",X"66",X"01",X"DD",X"6E",X"00",X"E5",X"D5",X"CD",X"75",
		X"2F",X"D1",X"E1",X"20",X"D6",X"CD",X"AD",X"2E",X"13",X"C1",X"10",X"CE",X"C9",X"1A",X"E5",X"CD",
		X"4D",X"27",X"E1",X"CD",X"F0",X"26",X"3E",X"2B",X"CD",X"35",X"27",X"C9",X"3A",X"F7",X"71",X"FE",
		X"00",X"28",X"25",X"06",X"09",X"DD",X"21",X"1D",X"5C",X"11",X"14",X"5C",X"DD",X"66",X"01",X"DD",
		X"6E",X"00",X"7E",X"EB",X"BE",X"EB",X"C0",X"DD",X"23",X"DD",X"23",X"DD",X"23",X"13",X"10",X"EC",
		X"3E",X"70",X"32",X"F7",X"71",X"18",X"0E",X"C9",X"21",X"3E",X"8B",X"11",X"1E",X"58",X"CD",X"49",
		X"19",X"3E",X"02",X"FE",X"02",X"3E",X"00",X"32",X"8D",X"72",X"C9",X"3A",X"93",X"72",X"FE",X"FF",
		X"20",X"05",X"AF",X"32",X"93",X"72",X"C9",X"C5",X"CB",X"07",X"47",X"3E",X"00",X"CB",X"17",X"4F",
		X"78",X"CB",X"0F",X"CB",X"0F",X"CB",X"0F",X"CB",X"0F",X"CB",X"0F",X"E6",X"01",X"A9",X"2F",X"CB",
		X"1F",X"3A",X"00",X"B8",X"3A",X"93",X"72",X"CB",X"17",X"32",X"93",X"72",X"C1",X"C9",X"CD",X"FB",
		X"2E",X"E6",X"03",X"3C",X"47",X"21",X"7A",X"55",X"23",X"10",X"FD",X"FD",X"7E",X"01",X"32",X"90",
		X"72",X"47",X"E5",X"23",X"23",X"23",X"23",X"7E",X"E1",X"B8",X"28",X"12",X"7E",X"FD",X"77",X"01",
		X"AF",X"FD",X"77",X"04",X"32",X"8F",X"72",X"21",X"EA",X"2F",X"CD",X"95",X"0C",X"C9",X"3A",X"8F",
		X"72",X"FE",X"05",X"28",X"E7",X"3C",X"32",X"8F",X"72",X"18",X"C3",X"C5",X"01",X"22",X"00",X"ED",
		X"43",X"A3",X"72",X"18",X"08",X"C5",X"01",X"12",X"00",X"ED",X"43",X"A3",X"72",X"7E",X"CD",X"3E",
		X"17",X"20",X"18",X"23",X"7E",X"CD",X"3E",X"17",X"20",X"11",X"11",X"20",X"00",X"19",X"7E",X"CD",
		X"3E",X"17",X"20",X"07",X"2B",X"7E",X"CD",X"3E",X"17",X"20",X"00",X"C1",X"C9",X"7C",X"D6",X"10",
		X"67",X"C9",X"D5",X"11",X"20",X"00",X"AF",X"ED",X"52",X"D1",X"C9",X"D5",X"11",X"20",X"00",X"19",
		X"D1",X"C9",X"21",X"8C",X"52",X"22",X"40",X"70",X"DD",X"21",X"80",X"75",X"11",X"05",X"09",X"CD",
		X"FE",X"18",X"C9",X"DD",X"21",X"88",X"75",X"11",X"05",X"09",X"CD",X"FE",X"18",X"C9",X"3A",X"2C",
		X"00",X"AC",X"00",X"00",X"00",X"00",X"2F",X"2B",X"00",X"CD",X"00",X"00",X"00",X"00",X"36",X"2A",
		X"00",X"BD",X"00",X"00",X"00",X"00",X"3F",X"2F",X"00",X"DD",X"00",X"1D",X"00",X"00",X"1C",X"00",
		X"00",X"1B",X"00",X"00",X"1A",X"00",X"00",X"19",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"DE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2A",X"24",X"20",X"00",X"00",X"00",X"29",X"25",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"25",X"20",X"1D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"1E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"25",X"22",X"00",X"00",X"00",X"00",X"2A",X"25",X"22",X"00",X"00",X"00",X"00",X"00",
		X"00",X"29",X"24",X"20",X"00",X"00",X"00",X"27",X"24",X"20",X"00",X"00",X"00",X"29",X"25",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"25",X"20",X"1D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"25",X"22",X"1E",X"00",X"00",X"00",X"25",X"20",X"1D",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"1E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"25",X"22",X"00",X"00",X"00",X"00",X"2E",X"25",X"22",X"00",X"00",X"00",X"00",X"00",
		X"00",X"2C",X"27",X"24",X"00",X"00",X"00",X"2A",X"27",X"24",X"00",X"00",X"00",X"29",X"25",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"25",X"20",X"1D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"25",X"22",X"1E",X"00",X"00",X"00",X"25",X"20",X"1D",
		X"19",X"1D",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"19",X"1E",X"22",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1B",X"20",X"24",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"19",X"1E",X"22",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"19",X"1D",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"29",X"2C",X"00",X"00",X"00",X"00",
		X"29",X"2C",X"00",X"00",X"00",X"00",X"29",X"2C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"2A",X"2E",X"00",X"00",X"00",X"00",X"2A",X"2E",X"00",X"00",X"00",X"00",X"2A",X"2E",
		X"00",X"2A",X"2E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2C",X"30",X"00",X"00",X"00",X"00",
		X"2C",X"30",X"00",X"00",X"00",X"00",X"2C",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"2A",X"2E",X"00",X"00",X"00",X"00",X"2A",X"2E",X"00",X"00",X"00",X"00",X"2A",X"2E",
		X"00",X"2A",X"2E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"29",X"2C",X"00",X"00",X"00",X"00",
		X"29",X"2C",X"00",X"00",X"00",X"00",X"29",X"2C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"2A",X"2E",X"00",X"00",X"00",X"00",X"2A",X"2E",X"00",X"00",X"00",X"00",X"2A",X"2E",
		X"00",X"2A",X"2E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2C",X"30",X"00",X"00",X"00",X"00",
		X"2C",X"30",X"00",X"00",X"00",X"00",X"2C",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"2A",X"2E",X"00",X"00",X"00",X"00",X"2A",X"2E",X"00",X"00",X"00",X"00",X"2A",X"2E",
		X"00",X"2A",X"2E",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"29",X"2C",X"00",X"00",X"00",X"00",
		X"29",X"2C",X"05",X"00",X"00",X"00",X"29",X"2C",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",
		X"00",X"06",X"2A",X"2E",X"00",X"00",X"00",X"00",X"2A",X"2E",X"0A",X"00",X"00",X"00",X"2A",X"2E",
		X"00",X"2A",X"2E",X"0D",X"00",X"00",X"00",X"00",X"00",X"08",X"2C",X"30",X"00",X"00",X"00",X"00",
		X"2C",X"30",X"0C",X"00",X"00",X"00",X"2C",X"30",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",
		X"00",X"06",X"2A",X"2E",X"00",X"00",X"00",X"00",X"2A",X"2E",X"0A",X"00",X"00",X"00",X"2A",X"2E",
		X"00",X"2A",X"2E",X"0D",X"00",X"00",X"00",X"00",X"00",X"01",X"29",X"2C",X"01",X"00",X"00",X"00",
		X"29",X"2C",X"05",X"00",X"00",X"00",X"29",X"2C",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",
		X"00",X"06",X"2A",X"2E",X"06",X"00",X"00",X"00",X"2A",X"2E",X"0A",X"00",X"00",X"00",X"2A",X"2E",
		X"00",X"2A",X"2E",X"0D",X"00",X"00",X"00",X"00",X"00",X"08",X"2C",X"30",X"08",X"00",X"00",X"00",
		X"2C",X"30",X"0C",X"00",X"00",X"00",X"2C",X"30",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",
		X"00",X"06",X"2A",X"2E",X"06",X"00",X"00",X"00",X"2A",X"2E",X"0A",X"00",X"00",X"06",X"2A",X"2E",
		X"00",X"2A",X"2E",X"0D",X"00",X"00",X"00",X"00",X"00",X"01",X"29",X"2C",X"00",X"00",X"00",X"00",
		X"29",X"2C",X"05",X"00",X"00",X"00",X"29",X"2C",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",
		X"00",X"06",X"2A",X"2E",X"00",X"00",X"00",X"00",X"2A",X"2E",X"0A",X"00",X"00",X"00",X"2A",X"2E",
		X"00",X"2A",X"2E",X"0D",X"00",X"00",X"00",X"00",X"00",X"08",X"2C",X"30",X"00",X"00",X"00",X"00",
		X"2C",X"30",X"0C",X"00",X"00",X"00",X"2C",X"30",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",
		X"00",X"06",X"2A",X"2E",X"00",X"00",X"00",X"00",X"2A",X"2E",X"0A",X"00",X"00",X"00",X"2A",X"2E",
		X"00",X"2A",X"2E",X"0D",X"00",X"00",X"00",X"00",X"00",X"01",X"29",X"2C",X"01",X"00",X"00",X"00",
		X"29",X"2C",X"05",X"00",X"00",X"00",X"29",X"2C",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",
		X"00",X"06",X"2A",X"2E",X"06",X"00",X"00",X"00",X"2A",X"2E",X"0A",X"00",X"00",X"00",X"2A",X"2E",
		X"00",X"2A",X"2E",X"0D",X"00",X"00",X"00",X"00",X"00",X"08",X"2C",X"30",X"08",X"00",X"00",X"00",
		X"2C",X"30",X"0C",X"00",X"00",X"00",X"2C",X"30",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",
		X"00",X"06",X"2A",X"2E",X"06",X"00",X"00",X"00",X"2A",X"2E",X"0A",X"00",X"00",X"06",X"2A",X"2E",
		X"00",X"2A",X"2E",X"0D",X"00",X"00",X"00",X"00",X"00",X"01",X"29",X"2C",X"00",X"00",X"00",X"00",
		X"29",X"2C",X"05",X"00",X"00",X"00",X"29",X"2C",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",
		X"00",X"06",X"2A",X"2E",X"00",X"00",X"00",X"00",X"2A",X"2E",X"0A",X"00",X"00",X"00",X"2A",X"2E",
		X"00",X"2A",X"2E",X"0D",X"00",X"00",X"00",X"00",X"00",X"08",X"2C",X"30",X"00",X"00",X"00",X"00",
		X"2C",X"30",X"0C",X"00",X"00",X"00",X"2C",X"30",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",
		X"00",X"06",X"2A",X"2E",X"00",X"00",X"00",X"00",X"2A",X"2E",X"0A",X"00",X"00",X"00",X"2A",X"2E",
		X"00",X"2A",X"2E",X"0D",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",
		X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",
		X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",
		X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",
		X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"25",X"00",X"00",X"20",X"00",X"00",X"22",X"00",
		X"00",X"1D",X"00",X"00",X"20",X"00",X"00",X"1D",X"00",X"00",X"1B",X"00",X"00",X"19",X"00",X"00",
		X"00",X"00",X"FF",X"01",X"00",X"00",X"02",X"00",X"00",X"03",X"00",X"00",X"04",X"00",X"00",X"05",
		X"00",X"00",X"06",X"00",X"00",X"07",X"00",X"00",X"08",X"00",X"00",X"09",X"00",X"00",X"0A",X"00",
		X"00",X"0B",X"00",X"00",X"0C",X"00",X"00",X"0D",X"00",X"00",X"0E",X"00",X"00",X"0F",X"00",X"00",
		X"10",X"00",X"00",X"11",X"00",X"00",X"12",X"00",X"00",X"13",X"00",X"00",X"14",X"00",X"00",X"15",
		X"00",X"00",X"16",X"00",X"00",X"17",X"00",X"00",X"18",X"00",X"00",X"19",X"00",X"00",X"1A",X"00",
		X"00",X"1B",X"00",X"00",X"1C",X"00",X"00",X"1D",X"00",X"00",X"1E",X"00",X"00",X"1F",X"00",X"00",
		X"20",X"00",X"00",X"21",X"00",X"00",X"22",X"00",X"00",X"23",X"00",X"00",X"00",X"00",X"FF",X"29",
		X"2C",X"00",X"29",X"2C",X"00",X"00",X"00",X"FF",X"00",X"32",X"FF",X"1B",X"00",X"00",X"00",X"00",
		X"00",X"27",X"00",X"00",X"00",X"00",X"00",X"24",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"14",X"19",X"1D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"16",
		X"19",X"1E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"14",X"19",X"1D",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"16",X"19",X"1E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"14",X"19",X"1D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"16",
		X"19",X"1E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"1B",X"29",X"00",X"00",
		X"00",X"1B",X"20",X"24",X"00",X"00",X"00",X"1D",X"20",X"25",X"00",X"00",X"FF",X"01",X"29",X"00",
		X"00",X"20",X"00",X"00",X"25",X"00",X"01",X"29",X"00",X"06",X"2A",X"00",X"00",X"22",X"00",X"00",
		X"25",X"00",X"00",X"2A",X"00",X"01",X"29",X"00",X"00",X"20",X"00",X"00",X"25",X"00",X"01",X"29",
		X"00",X"06",X"2A",X"00",X"00",X"22",X"00",X"00",X"25",X"00",X"00",X"2A",X"00",X"01",X"29",X"00",
		X"00",X"20",X"00",X"00",X"25",X"00",X"01",X"29",X"00",X"06",X"2A",X"00",X"00",X"22",X"00",X"00",
		X"25",X"00",X"00",X"2A",X"00",X"08",X"29",X"00",X"00",X"00",X"00",X"0C",X"30",X"00",X"00",X"00",
		X"00",X"0D",X"31",X"00",X"00",X"00",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"E3",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",
		X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"E1",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"6B",X"71",X"71",X"71",X"71",X"71",X"71",X"71",X"71",X"6C",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"6F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"6F",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F5",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"EF",
		X"FF",X"FF",X"6F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"6F",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"6F",X"FF",X"FF",X"6B",X"71",X"71",X"71",X"71",X"71",X"6A",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"6F",X"FF",X"FF",X"6F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F7",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F0",
		X"FF",X"FF",X"70",X"71",X"71",X"6A",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F5",X"F8",X"F8",X"F4",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F5",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"F8",X"F8",X"F8",X"F4",X"FF",X"FF",X"EA",X"F8",X"F2",X"FF",X"FF",X"F6",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"F5",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"F8",X"F8",X"F8",X"F2",X"FF",X"FF",X"F3",X"F8",X"F4",X"FF",X"FF",X"F6",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F7",X"F8",X"F8",X"F2",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F5",X"F8",X"F8",X"F8",
		X"F8",X"F8",X"F8",X"F8",X"F8",X"F4",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F5",X"F8",X"F8",X"F4",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F7",X"F8",X"F4",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"F7",X"F8",X"EF",X"FF",X"FF",X"F6",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F7",X"F8",X"F8",X"F8",X"F8",X"F0",X"FF",X"FF",X"F7",X"F8",
		X"F8",X"F8",X"F8",X"F8",X"F8",X"F2",X"FF",X"FF",X"F7",X"F8",X"F8",X"F2",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"E2",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",
		X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"E0",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"E3",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",
		X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"E1",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F5",X"F8",X"F8",X"F4",X"FF",X"FF",X"F5",X"F8",X"F8",X"F4",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F5",X"F8",X"F8",X"F8",X"F8",X"EF",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"F5",X"F8",X"F0",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",
		X"FF",X"FF",X"F5",X"F8",X"F8",X"F8",X"F2",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",
		X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",
		X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"E9",X"FF",X"FF",X"EC",X"FF",X"FF",X"E9",X"FF",X"FF",X"EC",
		X"FF",X"FF",X"F7",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F2",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F5",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F4",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F7",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F2",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"E8",X"FF",X"FF",X"ED",X"FF",X"FF",X"E8",X"FF",X"FF",X"ED",
		X"FF",X"FF",X"F5",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F4",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",
		X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",
		X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",
		X"FF",X"FF",X"F7",X"F8",X"F8",X"F8",X"F4",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"F7",X"F8",X"EF",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F7",X"F8",X"F8",X"F2",X"FF",X"FF",X"F7",X"F8",X"F8",X"F2",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"F8",X"F8",X"F8",X"F8",X"F0",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"E2",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",
		X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"E0",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"E3",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",
		X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"E1",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F5",X"F8",X"F8",X"EF",X"FF",X"FF",X"F5",X"F8",X"F9",X"FF",
		X"FF",X"EB",X"F8",X"F4",X"FF",X"FF",X"EA",X"F8",X"F8",X"F8",X"F8",X"F4",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F7",X"F8",X"F8",X"F0",X"FF",X"FF",X"F7",X"F8",X"F8",X"F8",
		X"F8",X"F8",X"F8",X"F2",X"FF",X"FF",X"F3",X"F8",X"F8",X"F8",X"F8",X"F2",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F5",X"F8",X"F8",X"F4",X"FF",X"FF",X"F5",X"F8",X"F8",X"F8",
		X"F8",X"F8",X"F8",X"F4",X"FF",X"FF",X"F5",X"F8",X"F8",X"F8",X"F8",X"F4",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"EC",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F7",X"F8",X"F4",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F1",X"FF",X"FF",X"F6",X"FF",X"FF",X"F5",X"F8",X"F2",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"F1",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"ED",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F3",X"F8",X"F8",X"F2",X"FF",X"FF",X"F7",X"F8",X"F8",X"F8",
		X"F8",X"F8",X"F8",X"F2",X"FF",X"FF",X"F7",X"F8",X"F8",X"F8",X"F8",X"F0",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F5",X"F8",X"F8",X"F4",X"FF",X"FF",X"F5",X"F8",X"F8",X"F8",
		X"F8",X"F8",X"F8",X"F4",X"FF",X"FF",X"F5",X"F8",X"F8",X"F8",X"F8",X"F4",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"F1",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"F1",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F7",X"F8",X"F8",X"F0",X"FF",X"FF",X"F7",X"F8",X"F8",X"F8",
		X"F9",X"FF",X"FF",X"EE",X"FF",X"FF",X"F3",X"F8",X"F8",X"F8",X"F8",X"F2",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"E2",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",
		X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"E0",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"E3",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",
		X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"E1",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F5",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F4",X"FF",X"FF",
		X"F5",X"F8",X"F8",X"F4",X"F5",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"EF",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",
		X"F6",X"FF",X"FF",X"F6",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EC",X"FF",X"FF",
		X"F6",X"FF",X"FF",X"F6",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F6",X"FF",X"FF",X"F6",X"F7",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F0",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"ED",X"FF",X"FF",
		X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",
		X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F5",X"F8",X"F8",X"F8",X"F8",X"F4",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F7",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F2",X"FF",X"FF",
		X"E9",X"FF",X"FF",X"EC",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E9",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"E8",X"FF",X"FF",X"EB",X"F8",X"F4",X"FF",X"FF",X"F5",X"F8",
		X"F8",X"F8",X"F8",X"F4",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",
		X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"E8",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",
		X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"E9",X"FF",
		X"FF",X"EB",X"F8",X"F2",X"FF",X"FF",X"F7",X"F8",X"F8",X"F8",X"F8",X"F2",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F7",X"F8",X"F8",X"F8",X"F8",X"F2",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"F5",X"F8",X"F8",X"F4",X"FF",X"FF",X"F5",X"F8",X"F8",X"F4",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"EA",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F4",
		X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F1",X"FF",X"FF",X"F6",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",
		X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",
		X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F3",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F2",
		X"FF",X"FF",X"E9",X"FF",X"FF",X"EC",X"FF",X"FF",X"F3",X"F8",X"F8",X"F2",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"E2",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",
		X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"E0",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"E3",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",
		X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"E1",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"6B",X"71",X"71",X"71",X"71",X"71",X"71",X"71",X"71",X"71",X"71",X"6C",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"6F",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F5",X"F8",X"F8",X"F4",X"FF",X"FF",X"E8",X"FF",X"FF",X"ED",
		X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"6F",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",
		X"FF",X"FF",X"F7",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F9",X"FF",X"FF",X"6D",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",
		X"FF",X"FF",X"F5",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F4",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",
		X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",
		X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F7",X"F8",X"F8",X"F2",
		X"FF",X"FF",X"F7",X"F8",X"F8",X"F8",X"F9",X"FF",X"FF",X"EB",X"F8",X"F2",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"EA",X"F8",X"F8",X"F4",
		X"FF",X"FF",X"F5",X"F8",X"F8",X"EF",X"FF",X"FF",X"F5",X"F8",X"F8",X"F4",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"E9",X"FF",X"FF",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",
		X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",
		X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E8",X"FF",X"FF",X"F6",
		X"FF",X"FF",X"F6",X"FF",X"FF",X"ED",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"E8",X"FF",X"FF",X"ED",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",
		X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F7",X"F8",X"F8",X"F2",
		X"FF",X"FF",X"F7",X"F8",X"F8",X"F2",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"F7",X"F8",X"F8",X"F8",X"F8",X"F8",X"F4",
		X"FF",X"FF",X"F5",X"F8",X"F8",X"F4",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",
		X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",
		X"FF",X"FF",X"F6",X"FF",X"FF",X"F1",X"FF",X"FF",X"F6",X"FF",X"FF",X"F1",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F7",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F2",
		X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"70",X"71",X"71",X"72",X"FF",X"FF",X"70",X"71",X"71",X"72",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"E2",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",
		X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"E0",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"E3",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",
		X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"E1",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"6B",X"71",X"71",X"71",X"71",X"71",X"71",X"6C",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"6B",X"71",X"71",X"71",X"71",X"71",X"71",X"6C",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"6F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"6F",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"6F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"F5",X"F8",
		X"F9",X"FF",X"FF",X"ED",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"6F",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"6F",X"FF",X"FF",X"F5",X"F8",X"F8",X"F8",X"F2",X"FF",X"FF",X"F6",X"FF",
		X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"F7",X"F8",X"F8",X"F8",X"F4",X"FF",X"FF",X"6F",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"6F",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",
		X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"6F",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"6F",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"F8",
		X"F8",X"F8",X"F8",X"F2",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"6F",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"6F",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"6F",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"6D",X"FF",X"FF",X"EC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E9",X"FF",X"FF",X"6D",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F5",X"F8",X"F8",X"F8",
		X"F8",X"F4",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F5",X"F8",X"F8",X"EF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",
		X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F5",X"F8",X"F8",X"F4",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",
		X"FF",X"F7",X"F8",X"EF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F1",X"FF",X"FF",X"F6",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"ED",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",
		X"FF",X"F5",X"F8",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F7",X"F8",X"F8",X"F2",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",
		X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F3",X"F8",X"F8",X"F2",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"F8",X"F8",X"F8",
		X"F8",X"F2",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"6E",X"FF",X"FF",X"ED",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E8",X"FF",X"FF",X"6E",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"6F",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"6F",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"6F",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F5",X"F8",
		X"F8",X"F8",X"F8",X"F4",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"6F",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"6F",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",
		X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"6F",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"6F",X"FF",X"FF",X"F7",X"F8",X"F8",X"F8",X"F4",X"FF",X"FF",X"F6",X"FF",
		X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"F5",X"F8",X"F8",X"F8",X"F2",X"FF",X"FF",X"6F",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"6F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"E9",X"FF",
		X"FF",X"EB",X"F8",X"F2",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"6F",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"6F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"6F",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"70",X"71",X"71",X"71",X"71",X"71",X"71",X"6A",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"70",X"71",X"71",X"71",X"71",X"71",X"71",X"6A",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"E2",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",
		X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"E0",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"EA",X"2F",X"42",X"59",X"2F",X"56",X"41",X"4C",X"41",X"44",X"4F",X"4E",X"2F",X"41",X"55",X"54",
		X"4F",X"4D",X"41",X"54",X"49",X"4F",X"4E",X"2F",X"31",X"39",X"38",X"33",X"3F",X"03",X"05",X"04",
		X"05",X"9B",X"4A",X"01",X"07",X"05",X"08",X"05",X"9B",X"54",X"02",X"05",X"05",X"06",X"05",X"9B",
		X"5C",X"03",X"03",X"07",X"04",X"07",X"9A",X"4A",X"04",X"07",X"07",X"08",X"07",X"9A",X"54",X"05",
		X"05",X"07",X"06",X"07",X"9A",X"5C",X"06",X"03",X"03",X"04",X"03",X"99",X"0A",X"07",X"07",X"03",
		X"08",X"03",X"99",X"14",X"08",X"05",X"03",X"06",X"03",X"99",X"1C",X"09",X"02",X"01",X"03",X"01",
		X"99",X"EF",X"05",X"05",X"03",X"06",X"03",X"99",X"1C",X"09",X"05",X"03",X"06",X"03",X"99",X"1C",
		X"09",X"05",X"03",X"06",X"03",X"99",X"1C",X"09",X"05",X"03",X"06",X"03",X"99",X"1C",X"09",X"03",
		X"11",X"04",X"11",X"9B",X"5C",X"02",X"02",X"03",X"03",X"03",X"99",X"D9",X"02",X"09",X"03",X"0A",
		X"03",X"99",X"10",X"03",X"07",X"09",X"08",X"09",X"9B",X"56",X"04",X"06",X"04",X"09",X"04",X"9A",
		X"8F",X"04",X"0D",X"06",X"0E",X"05",X"9A",X"14",X"04",X"03",X"02",X"04",X"02",X"99",X"16",X"04",
		X"09",X"03",X"0A",X"03",X"98",X"DC",X"04",X"05",X"03",X"06",X"03",X"9B",X"4C",X"01",X"03",X"04",
		X"04",X"04",X"9A",X"EA",X"01",X"09",X"03",X"0A",X"03",X"98",X"DC",X"04",X"0B",X"03",X"0D",X"03",
		X"9A",X"36",X"04",X"09",X"03",X"0A",X"03",X"98",X"DC",X"04",X"09",X"03",X"0A",X"03",X"98",X"DC",
		X"04",X"09",X"03",X"0A",X"03",X"9B",X"50",X"03",X"03",X"05",X"04",X"05",X"9B",X"56",X"06",X"03",
		X"05",X"04",X"05",X"9B",X"5C",X"02",X"05",X"05",X"06",X"05",X"9A",X"8C",X"05",X"05",X"03",X"06",
		X"03",X"9A",X"54",X"07",X"05",X"07",X"06",X"07",X"9A",X"5C",X"01",X"07",X"03",X"08",X"03",X"99",
		X"1C",X"09",X"03",X"07",X"04",X"07",X"99",X"94",X"04",X"07",X"07",X"08",X"07",X"99",X"8E",X"08",
		X"07",X"07",X"08",X"07",X"99",X"8E",X"08",X"07",X"07",X"08",X"07",X"99",X"8E",X"08",X"07",X"07",
		X"08",X"07",X"99",X"8E",X"08",X"07",X"07",X"08",X"07",X"99",X"8E",X"08",X"07",X"07",X"08",X"07",
		X"99",X"8E",X"08",X"03",X"07",X"04",X"07",X"99",X"8A",X"01",X"07",X"03",X"08",X"03",X"99",X"9A",
		X"02",X"05",X"03",X"06",X"03",X"99",X"1C",X"02",X"03",X"07",X"04",X"07",X"99",X"90",X"03",X"05",
		X"03",X"06",X"03",X"9B",X"5C",X"04",X"07",X"03",X"08",X"03",X"9A",X"DA",X"04",X"03",X"07",X"04",
		X"07",X"9B",X"4A",X"05",X"03",X"07",X"04",X"07",X"9B",X"50",X"06",X"15",X"01",X"16",X"01",X"9A",
		X"1C",X"07",X"03",X"07",X"04",X"07",X"9B",X"50",X"06",X"03",X"07",X"04",X"07",X"9B",X"50",X"06",
		X"03",X"07",X"04",X"07",X"9B",X"50",X"06",X"03",X"07",X"04",X"07",X"9B",X"50",X"06",X"03",X"07",
		X"04",X"07",X"9B",X"50",X"06",X"06",X"03",X"07",X"03",X"9B",X"50",X"03",X"03",X"07",X"04",X"07",
		X"9B",X"4A",X"03",X"03",X"0B",X"04",X"0B",X"9A",X"0A",X"02",X"03",X"05",X"04",X"05",X"9A",X"90",
		X"05",X"03",X"07",X"04",X"07",X"99",X"90",X"07",X"03",X"05",X"04",X"05",X"9B",X"96",X"01",X"03",
		X"05",X"04",X"05",X"9A",X"96",X"09",X"03",X"0D",X"04",X"0D",X"9B",X"9C",X"04",X"09",X"03",X"0A",
		X"03",X"99",X"9C",X"08",X"0B",X"03",X"0C",X"03",X"98",X"DE",X"06",X"0B",X"03",X"0C",X"03",X"98",
		X"DE",X"06",X"0B",X"03",X"0C",X"03",X"98",X"DE",X"06",X"0B",X"03",X"0C",X"03",X"98",X"DE",X"06",
		X"0B",X"03",X"0C",X"03",X"98",X"DE",X"06",X"04",X"03",X"05",X"03",X"9B",X"8C",X"03",X"03",X"07",
		X"04",X"07",X"9B",X"88",X"03",X"03",X"05",X"04",X"05",X"9A",X"4A",X"02",X"03",X"04",X"04",X"04",
		X"99",X"48",X"05",X"07",X"03",X"08",X"03",X"98",X"CC",X"05",X"05",X"07",X"06",X"07",X"9A",X"72",
		X"01",X"02",X"03",X"03",X"03",X"9A",X"34",X"01",X"05",X"03",X"06",X"03",X"9B",X"54",X"04",X"05",
		X"03",X"06",X"03",X"99",X"14",X"08",X"03",X"05",X"04",X"05",X"9A",X"5C",X"09",X"07",X"03",X"08",
		X"03",X"9B",X"9E",X"06",X"03",X"04",X"04",X"04",X"9B",X"3E",X"06",X"03",X"04",X"04",X"04",X"99",
		X"5E",X"07",X"07",X"03",X"08",X"03",X"98",X"DE",X"07",X"F7",X"F6",X"F6",X"F6",X"F6",X"F6",X"F6",
		X"F5",X"3F",X"F7",X"F6",X"F4",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F2",X"F6",X"F5",X"3F",X"F2",
		X"F6",X"F6",X"F6",X"F6",X"F6",X"F6",X"F6",X"F6",X"F6",X"F6",X"F4",X"3F",X"A4",X"C8",X"54",X"58",
		X"5C",X"60",X"64",X"68",X"6C",X"70",X"74",X"A6",X"CA",X"56",X"5A",X"5E",X"62",X"66",X"6A",X"6E",
		X"72",X"76",X"A5",X"C9",X"55",X"59",X"5D",X"61",X"65",X"69",X"6D",X"71",X"75",X"A7",X"CB",X"57",
		X"5B",X"5F",X"63",X"67",X"6B",X"6F",X"73",X"77",X"13",X"15",X"FF",X"1A",X"15",X"25",X"FF",X"20",
		X"19",X"13",X"1B",X"19",X"1E",X"10",X"15",X"23",X"24",X"FF",X"1C",X"11",X"3F",X"13",X"22",X"15",
		X"11",X"24",X"19",X"1F",X"1E",X"FF",X"1F",X"22",X"19",X"17",X"19",X"1E",X"11",X"1C",X"15",X"FF",
		X"14",X"15",X"3F",X"26",X"11",X"1C",X"11",X"14",X"1F",X"1E",X"FF",X"11",X"25",X"24",X"1F",X"1D",
		X"11",X"24",X"19",X"1F",X"1E",X"3F",X"13",X"1F",X"20",X"29",X"22",X"19",X"17",X"18",X"24",X"FF",
		X"01",X"09",X"08",X"03",X"3F",X"1D",X"15",X"15",X"FF",X"1F",X"00",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"FF",X"1E",X"00",X"1F",X"1F",X"1F",X"1F",X"1F",X"FF",X"1E",X"00",X"1F",X"1F",X"00",X"00",X"B2",
		X"05",X"61",X"05",X"14",X"05",X"CC",X"04",X"86",X"04",X"45",X"04",X"08",X"04",X"CE",X"03",X"97",
		X"03",X"63",X"03",X"34",X"03",X"05",X"03",X"D9",X"02",X"B0",X"02",X"8A",X"02",X"66",X"02",X"43",
		X"02",X"22",X"02",X"04",X"02",X"E7",X"01",X"CB",X"01",X"B2",X"01",X"99",X"01",X"82",X"01",X"6D",
		X"01",X"58",X"01",X"45",X"01",X"33",X"01",X"22",X"01",X"11",X"01",X"02",X"01",X"F4",X"00",X"E6",
		X"00",X"D9",X"00",X"CD",X"00",X"C1",X"00",X"B6",X"00",X"AC",X"00",X"A2",X"00",X"9A",X"00",X"91",
		X"00",X"89",X"00",X"81",X"00",X"7A",X"00",X"73",X"00",X"6C",X"00",X"66",X"00",X"61",X"00",X"5B",
		X"00",X"40",X"38",X"30",X"30",X"28",X"20",X"18",X"FF",X"FE",X"40",X"41",X"42",X"43",X"44",X"45",
		X"46",X"47",X"48",X"49",X"4A",X"4B",X"4C",X"4D",X"4E",X"4F",X"A7",X"A6",X"A5",X"A4",X"A3",X"A2",
		X"A1",X"A0",X"9F",X"9E",X"9D",X"9C",X"9B",X"9A",X"99",X"98",X"DB",X"DA",X"D9",X"D8",X"C1",X"C1",
		X"CA",X"C9",X"C8",X"C1",X"3F",X"D7",X"D6",X"D5",X"D4",X"D0",X"CE",X"CC",X"C7",X"C6",X"C5",X"3F",
		X"C1",X"D3",X"D2",X"D1",X"CF",X"CD",X"CB",X"C4",X"C3",X"C2",X"3F",X"C0",X"BF",X"BE",X"BD",X"BE",
		X"BC",X"BB",X"BE",X"3F",X"00",X"00",X"01",X"02",X"03",X"04",X"05",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"00",X"06",X"07",X"08",X"09",
		X"0A",X"0B",X"00",X"00",X"00",X"00",X"00",X"0C",X"0D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"3F",X"00",X"00",X"50",X"0E",X"0F",X"00",X"10",X"11",X"12",X"00",X"00",X"13",X"14",X"15",
		X"00",X"16",X"17",X"00",X"00",X"00",X"18",X"00",X"3F",X"00",X"19",X"1A",X"1B",X"1C",X"1D",X"1E",
		X"1F",X"20",X"21",X"22",X"23",X"24",X"25",X"26",X"27",X"28",X"29",X"2A",X"2B",X"4F",X"00",X"3F",
		X"00",X"2C",X"2D",X"2E",X"2F",X"30",X"31",X"32",X"33",X"34",X"35",X"36",X"37",X"38",X"39",X"3A",
		X"3B",X"3C",X"3D",X"3E",X"00",X"00",X"3F",X"00",X"51",X"40",X"00",X"00",X"41",X"42",X"43",X"44",
		X"45",X"46",X"47",X"48",X"49",X"4A",X"4B",X"4C",X"4D",X"4E",X"00",X"00",X"00",X"3F",X"13",X"15",
		X"10",X"1A",X"15",X"25",X"10",X"1C",X"15",X"10",X"12",X"11",X"17",X"1E",X"11",X"22",X"14",X"10",
		X"11",X"10",X"15",X"24",X"15",X"10",X"13",X"22",X"15",X"15",X"3F",X"20",X"11",X"22",X"10",X"26",
		X"11",X"1C",X"11",X"14",X"1F",X"1E",X"10",X"11",X"25",X"24",X"1F",X"1D",X"11",X"24",X"19",X"1F",
		X"1E",X"3F",X"00",X"42",X"01",X"13",X"14",X"17",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"00",X"51",X"01",X"17",X"20",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"00",X"60",X"01",X"26",X"17",X"15",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"00",X"79",X"01",X"16",X"1D",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"00",X"89",X"01",X"26",X"2B",X"11",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"04",X"00",X"04",X"01",X"00",X"04",X"02",X"04",X"01",X"03",X"04",X"04",X"01",X"02",
		X"03",X"04",X"03",X"01",X"04",X"02",X"04",X"03",X"00",X"00",X"02",X"04",X"02",X"03",X"04",X"01",
		X"04",X"04",X"00",X"02",X"00",X"04",X"00",X"03",X"00",X"01",X"FD",X"02",X"01",X"04",X"03",X"FC",
		X"02",X"01",X"04",X"03",X"FB",X"02",X"01",X"04",X"03",X"FA",X"02",X"01",X"04",X"03",X"00",X"FA",
		X"FD",X"FC",X"FB",X"F5",X"F3",X"F0",X"EF",X"FA",X"FD",X"FC",X"FB",X"FA",X"FA",X"FA",X"FA",X"72",
		X"71",X"70",X"6F",X"6E",X"6D",X"6C",X"6B",X"6A",X"69",X"69",X"3A",X"2C",X"6F",X"E0",X"00",X"00",
		X"00",X"00",X"2F",X"2B",X"70",X"20",X"00",X"00",X"00",X"00",X"36",X"2A",X"98",X"E0",X"00",X"00",
		X"00",X"00",X"2F",X"2F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"40",X"10",X"08",X"40",
		X"20",X"08",X"10",X"8A",X"DC",X"42",X"02",X"00",X"00",X"33",X"4B",X"E0",X"8B",X"0A",X"42",X"02",
		X"00",X"00",X"23",X"3B",X"50",X"8A",X"8A",X"42",X"02",X"00",X"10",X"43",X"5B",X"50",X"89",X"4A",
		X"42",X"02",X"00",X"30",X"93",X"AB",X"50",X"88",X"CA",X"42",X"02",X"00",X"40",X"B3",X"CB",X"50",
		X"8A",X"0A",X"42",X"02",X"00",X"00",X"63",X"7B",X"50",X"89",X"8A",X"42",X"02",X"00",X"10",X"83",
		X"9B",X"50",X"8A",X"FC",X"42",X"02",X"00",X"20",X"2B",X"43",X"E0",X"88",X"DC",X"42",X"02",X"00",
		X"30",X"B3",X"CB",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"89",X"4A",X"42",
		X"02",X"00",X"00",X"93",X"AB",X"50",X"88",X"CA",X"42",X"02",X"00",X"10",X"B3",X"CB",X"50",X"89",
		X"FC",X"42",X"02",X"00",X"00",X"6B",X"83",X"E0",X"89",X"04",X"42",X"02",X"00",X"00",X"A3",X"BB",
		X"20",X"8B",X"10",X"42",X"02",X"00",X"10",X"23",X"3B",X"80",X"89",X"DC",X"42",X"02",X"00",X"30",
		X"73",X"8B",X"E0",X"11",X"05",X"00",X"CD",X"AD",X"13",X"06",X"17",X"DD",X"7E",X"02",X"3D",X"FD",
		X"BE",X"00",X"28",X"12",X"3C",X"FD",X"BE",X"00",X"28",X"0C",X"3C",X"FD",X"BE",X"00",X"28",X"06",
		X"3C",X"FD",X"BE",X"00",X"20",X"1B",X"DD",X"7E",X"03",X"3D",X"FD",X"BE",X"01",X"28",X"1B",X"3C",
		X"FD",X"BE",X"01",X"28",X"15",X"3C",X"FD",X"BE",X"01",X"28",X"0F",X"3C",X"FD",X"BE",X"01",X"28",
		X"09",X"FD",X"23",X"FD",X"23",X"10",X"C4",X"AF",X"77",X"C9",X"3E",X"01",X"7E",X"FE",X"01",X"3E",
		X"00",X"C8",X"3E",X"01",X"77",X"C9",X"CD",X"75",X"56",X"C9",X"78",X"77",X"E5",X"7C",X"C6",X"08",
		X"67",X"FF",X"6A",X"7A",X"0F",X"8D",X"6B",X"7F",X"FE",X"45",X"0F",X"54",X"BE",X"55",X"1F",X"6C",
		X"50",X"4C",X"41",X"59",X"45",X"52",X"2F",X"31",X"3F",X"43",X"52",X"45",X"44",X"49",X"54",X"3F",
		X"2F",X"2F",X"2F",X"48",X"49",X"47",X"48",X"2F",X"53",X"43",X"4F",X"52",X"45",X"2F",X"2F",X"2F",
		X"3F",X"47",X"41",X"4D",X"45",X"2F",X"4F",X"56",X"45",X"52",X"2F",X"3F",X"2F",X"2F",X"2F",X"2F",
		X"2F",X"49",X"4E",X"53",X"45",X"52",X"54",X"2F",X"43",X"4F",X"49",X"4E",X"53",X"2F",X"2F",X"2F",
		X"2F",X"2F",X"3F",X"2F",X"2F",X"2F",X"2F",X"2F",X"50",X"55",X"53",X"48",X"2F",X"53",X"54",X"41",
		X"52",X"54",X"2F",X"42",X"55",X"54",X"54",X"4F",X"4E",X"2F",X"2F",X"2F",X"2F",X"2F",X"3F",X"2F",
		X"4F",X"4E",X"45",X"2F",X"50",X"4C",X"41",X"59",X"45",X"52",X"2F",X"4F",X"4E",X"4C",X"59",X"2F",
		X"2F",X"3F",X"4F",X"4E",X"45",X"2F",X"4F",X"52",X"2F",X"54",X"57",X"4F",X"2F",X"50",X"4C",X"41",
		X"59",X"45",X"52",X"53",X"3F",X"42",X"4F",X"4E",X"55",X"53",X"3F",X"56",X"41",X"4C",X"41",X"44",
		X"4F",X"4E",X"2F",X"41",X"55",X"54",X"4F",X"4D",X"41",X"54",X"49",X"4F",X"4E",X"3F",X"2F",X"2F",
		X"2F",X"2F",X"2F",X"2F",X"4D",X"4F",X"56",X"45",X"2F",X"4A",X"4F",X"59",X"53",X"54",X"49",X"43",
		X"4B",X"2F",X"2F",X"2F",X"2F",X"2F",X"3F",X"2F",X"2F",X"54",X"4F",X"2F",X"44",X"49",X"53",X"50",
		X"4C",X"41",X"59",X"2F",X"59",X"4F",X"55",X"52",X"2F",X"4E",X"41",X"4D",X"45",X"2F",X"3F",X"53",
		X"43",X"4F",X"52",X"45",X"3F",X"4E",X"41",X"4D",X"45",X"3F",X"50",X"4C",X"41",X"59",X"45",X"52",
		X"2F",X"31",X"3F",X"50",X"4C",X"41",X"59",X"45",X"52",X"2F",X"32",X"3F",X"2F",X"2F",X"2F",X"2F",
		X"2F",X"2F",X"2F",X"2F",X"3F",X"2F",X"2F",X"45",X"4E",X"44",X"2F",X"42",X"59",X"2F",X"41",X"43",
		X"54",X"49",X"4F",X"4E",X"2F",X"42",X"55",X"54",X"54",X"4F",X"4E",X"3F",X"2F",X"2F",X"3F",X"43",
		X"4F",X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"2F",X"31",X"39",X"38",X"33",X"3F",X"52",X"45",
		X"41",X"44",X"59",X"3F",X"42",X"4F",X"4E",X"55",X"53",X"3F",X"43",X"4F",X"4E",X"47",X"52",X"41",
		X"54",X"55",X"4C",X"41",X"54",X"49",X"4F",X"4E",X"3F",X"2F",X"A8",X"DD",X"DC",X"DB",X"DA",X"2F",
		X"3F",X"B5",X"B4",X"B3",X"B2",X"B1",X"AE",X"AD",X"2F",X"AC",X"AB",X"CD",X"CC",X"CB",X"CA",X"C9",
		X"C8",X"2F",X"3F",X"2F",X"2F",X"BE",X"BD",X"BC",X"BB",X"BA",X"2F",X"2F",X"3F",X"2F",X"2F",X"2F",
		X"43",X"4F",X"4D",X"50",X"4C",X"45",X"54",X"45",X"2F",X"50",X"55",X"5A",X"5A",X"4C",X"45",X"2F",
		X"4C",X"49",X"4B",X"45",X"2F",X"54",X"48",X"49",X"53",X"2F",X"3F",X"2F",X"2F",X"42",X"45",X"46",
		X"4F",X"52",X"45",X"2F",X"2F",X"3F",X"2F",X"2F",X"2F",X"42",X"4F",X"4E",X"55",X"53",X"2F",X"47",
		X"45",X"54",X"53",X"2F",X"54",X"4F",X"2F",X"5A",X"45",X"52",X"4F",X"2F",X"2F",X"3F",X"2F",X"2F",
		X"2F",X"53",X"4F",X"52",X"52",X"59",X"2F",X"4E",X"4F",X"2F",X"42",X"4F",X"4E",X"55",X"53",X"2F",
		X"2F",X"3F",X"43",X"4F",X"4E",X"47",X"52",X"41",X"54",X"55",X"4C",X"41",X"54",X"49",X"4F",X"4E",
		X"53",X"3F",X"46",X"52",X"45",X"45",X"2F",X"50",X"4C",X"41",X"59",X"3F",X"41",X"43",X"54",X"3F",
		X"3F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"3F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",
		X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",
		X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",
		X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",
		X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",
		X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",
		X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",
		X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",
		X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"5E",X"50",X"49",X"43",
		X"4B",X"45",X"52",X"5D",X"3F",X"5E",X"54",X"52",X"41",X"4E",X"53",X"50",X"4F",X"53",X"45",X"52",
		X"5D",X"3F",X"5E",X"44",X"49",X"53",X"54",X"55",X"52",X"42",X"45",X"52",X"5D",X"3F",X"5E",X"4B",
		X"49",X"4C",X"4C",X"45",X"52",X"5D",X"3F",X"4A",X"4F",X"55",X"45",X"55",X"52",X"2F",X"31",X"3F",
		X"43",X"52",X"45",X"44",X"49",X"54",X"3F",X"4D",X"45",X"49",X"4C",X"4C",X"45",X"55",X"52",X"53",
		X"2F",X"53",X"43",X"4F",X"52",X"45",X"53",X"3F",X"4A",X"45",X"55",X"2F",X"46",X"49",X"4E",X"49",
		X"2F",X"2F",X"3F",X"49",X"4E",X"54",X"52",X"4F",X"44",X"55",X"49",X"53",X"45",X"5A",X"2F",X"56",
		X"4F",X"53",X"2F",X"50",X"49",X"45",X"43",X"45",X"53",X"3F",X"41",X"50",X"50",X"55",X"59",X"45",
		X"5A",X"2F",X"53",X"55",X"52",X"2F",X"4C",X"45",X"2F",X"42",X"4F",X"55",X"54",X"4F",X"4E",X"2F",
		X"53",X"54",X"41",X"52",X"54",X"3F",X"31",X"2F",X"4A",X"4F",X"55",X"45",X"55",X"52",X"2F",X"53",
		X"45",X"55",X"4C",X"45",X"4D",X"45",X"4E",X"54",X"3F",X"2F",X"2F",X"31",X"2F",X"30",X"55",X"2F",
		X"32",X"2F",X"4A",X"4F",X"55",X"45",X"55",X"52",X"53",X"2F",X"2F",X"3F",X"42",X"4F",X"4E",X"55",
		X"53",X"3F",X"56",X"41",X"4C",X"41",X"44",X"4F",X"4E",X"2F",X"41",X"55",X"54",X"4F",X"4D",X"41",
		X"54",X"49",X"4F",X"4E",X"3F",X"55",X"54",X"49",X"4C",X"49",X"53",X"45",X"5A",X"2F",X"4C",X"45",
		X"2F",X"4D",X"41",X"4E",X"49",X"50",X"55",X"4C",X"41",X"54",X"45",X"55",X"52",X"3F",X"50",X"4F",
		X"55",X"52",X"2F",X"49",X"4E",X"53",X"43",X"52",X"49",X"52",X"45",X"2F",X"56",X"4F",X"54",X"52",
		X"45",X"2F",X"4E",X"4F",X"4D",X"3F",X"53",X"43",X"4F",X"52",X"45",X"3F",X"4E",X"4F",X"4D",X"2F",
		X"3F",X"4A",X"4F",X"55",X"45",X"55",X"52",X"2F",X"31",X"3F",X"4A",X"4F",X"55",X"45",X"55",X"52",
		X"2F",X"32",X"3F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"3F",X"2F",X"2F",X"2F",X"41",
		X"43",X"54",X"49",X"4F",X"4E",X"2F",X"50",X"4F",X"55",X"52",X"2F",X"46",X"49",X"4E",X"49",X"52",
		X"3F",X"2F",X"2F",X"2F",X"2F",X"3F",X"43",X"4F",X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"2F",
		X"31",X"39",X"38",X"33",X"3F",X"2F",X"50",X"52",X"45",X"54",X"3F",X"42",X"4F",X"4E",X"55",X"53",
		X"3F",X"2F",X"46",X"45",X"4C",X"49",X"43",X"49",X"54",X"41",X"54",X"49",X"4F",X"4E",X"53",X"2F",
		X"D9",X"D8",X"D7",X"D6",X"D5",X"D4",X"D3",X"3F",X"2F",X"B9",X"B8",X"B7",X"B6",X"AE",X"AD",X"2F",
		X"AC",X"AB",X"D2",X"D1",X"D0",X"CF",X"CE",X"2F",X"2F",X"3F",X"C7",X"C6",X"C5",X"C4",X"C3",X"C2",
		X"C1",X"C0",X"BF",X"3F",X"2F",X"2F",X"2F",X"2F",X"2F",X"43",X"4F",X"4D",X"50",X"4C",X"45",X"54",
		X"45",X"5A",X"2F",X"4C",X"45",X"2F",X"50",X"55",X"5A",X"5A",X"4C",X"45",X"2F",X"2F",X"2F",X"2F",
		X"2F",X"3F",X"41",X"56",X"41",X"4E",X"54",X"2F",X"51",X"55",X"45",X"2F",X"3F",X"4C",X"45",X"2F",
		X"42",X"4F",X"4E",X"55",X"53",X"2F",X"4E",X"45",X"2F",X"53",X"4F",X"49",X"54",X"2F",X"41",X"2F",
		X"5A",X"45",X"52",X"4F",X"3F",X"44",X"45",X"53",X"4F",X"4C",X"45",X"2F",X"50",X"41",X"53",X"2F",
		X"44",X"45",X"2F",X"42",X"4F",X"4E",X"55",X"53",X"3F",X"46",X"45",X"4C",X"49",X"43",X"49",X"54",
		X"41",X"54",X"49",X"4F",X"4E",X"53",X"3F",X"2F",X"2F",X"46",X"52",X"45",X"45",X"2F",X"50",X"4C",
		X"41",X"59",X"3F",X"41",X"43",X"54",X"45",X"3F",X"80",X"4A",X"F0",X"80",X"4A",X"F7",X"80",X"4B",
		X"47",X"40",X"4B",X"53",X"40",X"FF",X"FF",X"FF",X"58",X"93",X"02",X"A8",X"91",X"01",X"12",X"91",
		X"01",X"98",X"90",X"01",X"2E",X"93",X"01",X"36",X"93",X"01",X"C8",X"91",X"02",X"4C",X"92",X"02",
		X"02",X"06",X"04",X"03",X"08",X"06",X"01",X"03",X"02",X"09",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"04",X"09",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"02",X"04",X"03",X"04",
		X"02",X"02",X"09",X"03",X"03",X"06",X"03",X"06",X"03",X"03",X"00",X"00",X"00",X"02",X"05",X"06",
		X"06",X"02",X"05",X"03",X"04",X"02",X"07",X"02",X"05",X"02",X"05",X"05",X"05",X"02",X"02",X"09",
		X"8B",X"51",X"8B",X"15",X"8B",X"05",X"8A",X"D3",X"89",X"1B",X"8A",X"C9",X"88",X"8F",X"88",X"D5",
		X"88",X"0B",X"8B",X"95",X"89",X"CF",X"88",X"05",X"89",X"95",X"89",X"95",X"89",X"95",X"89",X"95",
		X"89",X"95",X"89",X"D5",X"89",X"17",X"8B",X"05",X"8B",X"91",X"89",X"C7",X"89",X"53",X"8B",X"4F",
		X"8A",X"0D",X"89",X"DB",X"88",X"87",X"89",X"DB",X"88",X"8D",X"89",X"1B",X"8B",X"47",X"8A",X"4D",
		X"8A",X"4D",X"8A",X"4D",X"8A",X"4D",X"8A",X"55",X"8B",X"07",X"8A",X"47",X"8A",X"5B",X"8B",X"0B",
		X"8A",X"DB",X"88",X"8D",X"88",X"97",X"89",X"15",X"8A",X"F3",X"89",X"C9",X"89",X"85",X"8A",X"4F",
		X"8B",X"45",X"89",X"9B",X"8A",X"5B",X"89",X"91",X"88",X"17",X"8A",X"27",X"9B",X"01",X"E7",X"9A",
		X"01",X"2D",X"9B",X"02",X"ED",X"9A",X"02",X"EF",X"9A",X"02",X"31",X"9B",X"02",X"2F",X"9B",X"02",
		X"F1",X"9A",X"02",X"37",X"9B",X"03",X"F7",X"9A",X"03",X"F9",X"9A",X"03",X"39",X"9B",X"03",X"A7",
		X"99",X"04",X"27",X"9A",X"04",X"E7",X"99",X"04",X"2D",X"9A",X"05",X"31",X"9A",X"05",X"AD",X"99",
		X"05",X"AF",X"99",X"05",X"EF",X"99",X"05",X"B1",X"99",X"05",X"2F",X"9A",X"05",X"F1",X"99",X"05",
		X"B7",X"99",X"06",X"37",X"9A",X"06",X"39",X"9A",X"06",X"F7",X"99",X"06",X"B9",X"99",X"06",X"F9",
		X"99",X"06",X"E7",X"98",X"07",X"ED",X"98",X"08",X"EF",X"98",X"08",X"F1",X"98",X"08",X"F7",X"98",
		X"09",X"F9",X"98",X"09",X"54",X"60",X"6C",X"58",X"64",X"70",X"5C",X"68",X"74",X"34",X"8A",X"01",
		X"36",X"8A",X"01",X"38",X"8A",X"02",X"F4",X"89",X"02",X"F6",X"89",X"02",X"F8",X"89",X"02",X"B4",
		X"89",X"02",X"B6",X"89",X"02",X"B8",X"89",X"03",X"DB",X"89",X"03",X"DB",X"89",X"03",X"DB",X"89",
		X"03",X"DB",X"89",X"04",X"DB",X"89",X"04",X"DB",X"89",X"04",X"DB",X"89",X"05",X"DB",X"89",X"05",
		X"DB",X"89",X"05",X"DB",X"89",X"05",X"DB",X"89",X"05",X"DB",X"89",X"05",X"DB",X"89",X"05",X"DB",
		X"89",X"05",X"DB",X"89",X"06",X"DB",X"89",X"06",X"DB",X"89",X"06",X"DB",X"89",X"06",X"DB",X"89",
		X"06",X"DB",X"89",X"06",X"DB",X"89",X"07",X"DB",X"89",X"08",X"DB",X"89",X"08",X"DB",X"89",X"08",
		X"DB",X"89",X"09",X"DB",X"89",X"09",X"27",X"9B",X"01",X"E7",X"9A",X"01",X"A7",X"9A",X"01",X"29",
		X"9B",X"01",X"39",X"9B",X"02",X"F9",X"9A",X"02",X"B9",X"9A",X"02",X"79",X"9A",X"02",X"39",X"9A",
		X"02",X"F9",X"99",X"02",X"B9",X"99",X"02",X"79",X"99",X"02",X"B7",X"99",X"02",X"E7",X"98",X"03",
		X"E9",X"98",X"03",X"EB",X"98",X"03",X"ED",X"98",X"03",X"ED",X"98",X"03",X"ED",X"98",X"03",X"ED",
		X"98",X"03",X"ED",X"98",X"03",X"ED",X"98",X"03",X"ED",X"98",X"03",X"ED",X"98",X"03",X"ED",X"98",
		X"03",X"ED",X"98",X"03",X"ED",X"98",X"03",X"ED",X"98",X"03",X"ED",X"98",X"03",X"ED",X"98",X"03",
		X"ED",X"98",X"03",X"ED",X"98",X"03",X"ED",X"98",X"03",X"ED",X"98",X"03",X"D9",X"98",X"03",X"37",
		X"9A",X"01",X"39",X"9A",X"01",X"F7",X"99",X"01",X"F9",X"99",X"01",X"B7",X"99",X"01",X"B9",X"99",
		X"01",X"39",X"9B",X"02",X"F9",X"9A",X"02",X"27",X"9B",X"03",X"29",X"9B",X"03",X"2B",X"9B",X"03",
		X"2D",X"9B",X"03",X"71",X"99",X"04",X"31",X"99",X"04",X"F1",X"98",X"04",X"67",X"9A",X"05",X"69",
		X"9A",X"05",X"27",X"9A",X"05",X"29",X"9A",X"05",X"33",X"9B",X"06",X"F3",X"9A",X"06",X"2F",X"9A",
		X"07",X"31",X"9A",X"07",X"67",X"99",X"08",X"69",X"99",X"08",X"6B",X"99",X"08",X"27",X"99",X"08",
		X"29",X"99",X"08",X"2B",X"99",X"08",X"E7",X"98",X"08",X"E9",X"98",X"08",X"EB",X"98",X"08",X"F5",
		X"98",X"09",X"F7",X"98",X"09",X"F9",X"98",X"09",X"E7",X"98",X"01",X"27",X"99",X"01",X"67",X"99",
		X"01",X"73",X"99",X"02",X"75",X"99",X"02",X"77",X"99",X"02",X"37",X"99",X"02",X"F7",X"98",X"02",
		X"F9",X"98",X"02",X"ED",X"98",X"03",X"2D",X"99",X"03",X"6D",X"99",X"03",X"B3",X"9A",X"04",X"B5",
		X"9A",X"04",X"B7",X"9A",X"04",X"F7",X"9A",X"04",X"37",X"9B",X"04",X"39",X"9B",X"04",X"27",X"9B",
		X"05",X"E7",X"9A",X"05",X"A7",X"9A",X"05",X"2D",X"9B",X"06",X"ED",X"9A",X"06",X"AD",X"9A",X"06",
		X"AD",X"9A",X"06",X"AD",X"9A",X"06",X"AD",X"9A",X"06",X"AD",X"9A",X"06",X"AD",X"9A",X"06",X"AD",
		X"9A",X"06",X"AD",X"9A",X"06",X"AD",X"9A",X"06",X"AD",X"9A",X"06",X"AD",X"9A",X"06",X"AD",X"9A",
		X"06",X"73",X"9B",X"01",X"33",X"9B",X"01",X"E7",X"99",X"02",X"A7",X"99",X"02",X"67",X"99",X"02",
		X"27",X"99",X"02",X"E7",X"98",X"02",X"27",X"9B",X"03",X"29",X"9B",X"03",X"2B",X"9B",X"03",X"2D",
		X"9B",X"03",X"E7",X"9A",X"03",X"A7",X"9A",X"03",X"79",X"9B",X"04",X"39",X"9B",X"04",X"F9",X"9A",
		X"04",X"B9",X"9A",X"04",X"79",X"9A",X"04",X"39",X"9A",X"04",X"6D",X"9A",X"05",X"2D",X"9A",X"05",
		X"B3",X"98",X"06",X"B5",X"98",X"06",X"B7",X"98",X"06",X"B9",X"98",X"06",X"BB",X"98",X"06",X"6D",
		X"99",X"07",X"2D",X"99",X"07",X"ED",X"98",X"07",X"73",X"99",X"08",X"75",X"99",X"08",X"77",X"99",
		X"08",X"79",X"99",X"08",X"73",X"9A",X"09",X"33",X"9A",X"09",X"4F",X"9A",X"01",X"4D",X"9A",X"01",
		X"0D",X"9A",X"01",X"0F",X"9A",X"01",X"11",X"9A",X"01",X"CD",X"99",X"01",X"CF",X"99",X"01",X"27",
		X"9A",X"02",X"E7",X"99",X"02",X"65",X"9B",X"03",X"67",X"9B",X"03",X"69",X"9B",X"03",X"25",X"9B",
		X"03",X"E5",X"9A",X"03",X"2F",X"9B",X"04",X"31",X"9B",X"04",X"25",X"99",X"05",X"E5",X"98",X"05",
		X"A5",X"98",X"05",X"A7",X"98",X"05",X"A9",X"98",X"05",X"77",X"9B",X"06",X"79",X"9B",X"06",X"7B",
		X"9B",X"06",X"3B",X"9B",X"06",X"FB",X"9A",X"06",X"B7",X"98",X"07",X"B9",X"98",X"07",X"BB",X"98",
		X"07",X"FB",X"98",X"07",X"3B",X"99",X"07",X"EF",X"98",X"08",X"F1",X"98",X"08",X"39",X"9A",X"09",
		X"F9",X"99",X"09",X"FE",X"F5",X"F0",X"EF",X"00",X"00",X"00",X"43",X"89",X"FC",X"63",X"89",X"FD",
		X"83",X"8A",X"FC",X"A3",X"8A",X"FD",X"6C",X"88",X"FC",X"6D",X"88",X"F8",X"76",X"88",X"FC",X"77",
		X"88",X"F8",X"5D",X"89",X"F8",X"7D",X"89",X"F3",X"9D",X"8A",X"F8",X"BD",X"8A",X"F3",X"8C",X"8B",
		X"FD",X"8D",X"8B",X"F3",X"96",X"8B",X"FD",X"97",X"8B",X"F3",X"97",X"8B",X"F3",X"58",X"20",X"70",
		X"20",X"A8",X"20",X"18",X"50",X"30",X"50",X"58",X"50",X"A8",X"50",X"C0",X"50",X"D8",X"50",X"D8",
		X"78",X"18",X"88",X"18",X"A0",X"30",X"A0",X"58",X"A0",X"A8",X"A0",X"D8",X"A0",X"C0",X"A0",X"58",
		X"E0",X"70",X"E0",X"A8",X"E0",X"80",X"A0",X"80",X"88",X"C0",X"78",X"58",X"20",X"A8",X"20",X"30",
		X"60",X"18",X"60",X"A8",X"80",X"C0",X"80",X"18",X"B0",X"90",X"A0",X"A8",X"A0",X"B8",X"E0",X"90",
		X"C8",X"B8",X"E0",X"B8",X"E0",X"B8",X"E0",X"B8",X"E0",X"B8",X"E0",X"B8",X"E0",X"B8",X"E0",X"B8",
		X"E0",X"B8",X"E0",X"B8",X"E0",X"B8",X"E0",X"B8",X"E0",X"68",X"20",X"88",X"20",X"68",X"38",X"88",
		X"38",X"68",X"50",X"88",X"50",X"68",X"68",X"88",X"68",X"68",X"80",X"88",X"80",X"68",X"D0",X"88",
		X"D0",X"68",X"E0",X"88",X"E0",X"30",X"E0",X"C0",X"E0",X"18",X"50",X"18",X"80",X"18",X"A0",X"D8",
		X"50",X"D8",X"80",X"D8",X"A0",X"D8",X"A0",X"30",X"20",X"48",X"20",X"88",X"20",X"88",X"38",X"30",
		X"50",X"48",X"60",X"58",X"60",X"88",X"60",X"B0",X"70",X"18",X"80",X"58",X"78",X"88",X"88",X"80",
		X"A0",X"18",X"98",X"30",X"B0",X"C0",X"E0",X"58",X"E0",X"A8",X"E0",X"18",X"B0",X"D8",X"70",X"B0",
		X"58",X"80",X"B8",X"D8",X"70",X"68",X"20",X"68",X"38",X"D8",X"50",X"88",X"50",X"70",X"50",X"88",
		X"68",X"30",X"80",X"48",X"80",X"88",X"80",X"B8",X"80",X"48",X"98",X"48",X"B0",X"70",X"B0",X"88",
		X"B0",X"A0",X"B0",X"B8",X"D8",X"E0",X"88",X"E0",X"88",X"E0",X"88",X"E0",X"88",X"E0",X"88",X"E0",
		X"88",X"E0",X"88",X"58",X"28",X"98",X"28",X"58",X"40",X"58",X"50",X"80",X"50",X"98",X"50",X"98",
		X"40",X"D0",X"60",X"D8",X"88",X"D0",X"A0",X"78",X"78",X"78",X"A0",X"20",X"60",X"18",X"78",X"20",
		X"A0",X"58",X"D8",X"98",X"D8",X"70",X"B0",X"58",X"C0",X"98",X"B0",X"98",X"B0",X"98",X"B0",X"98",
		X"B0",X"0F",X"02",X"37",X"1F",X"00",X"00",X"FF",X"04",X"00",X"0F",X"1F",X"37",X"1F",X"00",X"00",
		X"FF",X"00",X"00",X"38",X"1F",X"1F",X"1F",X"FF",X"2E",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"01");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
