library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity burger_time_prog is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of burger_time_prog is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"4C",X"3C",X"CF",X"4C",X"0F",X"C0",X"85",X"F5",X"EA",X"4C",X"03",X"B0",X"85",X"F5",X"EA",X"78",
		X"D8",X"A2",X"FF",X"9A",X"AD",X"03",X"40",X"29",X"10",X"F0",X"EE",X"A9",X"00",X"85",X"01",X"85",
		X"F9",X"8D",X"00",X"40",X"20",X"32",X"C3",X"20",X"1D",X"C3",X"A9",X"01",X"85",X"01",X"A9",X"00",
		X"85",X"1A",X"20",X"0D",X"C7",X"85",X"F7",X"EA",X"A9",X"FE",X"8D",X"05",X"50",X"A9",X"00",X"8D",
		X"02",X"40",X"85",X"1B",X"85",X"20",X"A9",X"00",X"85",X"1C",X"20",X"16",X"C4",X"A2",X"FF",X"20",
		X"2C",X"CA",X"20",X"D9",X"C3",X"A2",X"FF",X"20",X"2C",X"CA",X"20",X"78",X"C4",X"A2",X"3F",X"20",
		X"2C",X"CA",X"20",X"61",X"C5",X"85",X"F5",X"EA",X"20",X"0D",X"C7",X"20",X"48",X"C7",X"A9",X"01",
		X"85",X"1C",X"85",X"F5",X"EA",X"20",X"67",X"C7",X"85",X"F5",X"EA",X"AD",X"03",X"40",X"10",X"FB",
		X"58",X"EA",X"EA",X"EA",X"EA",X"78",X"20",X"45",X"D0",X"20",X"6E",X"D0",X"E6",X"13",X"A5",X"13",
		X"29",X"3F",X"D0",X"03",X"85",X"F5",X"EA",X"E6",X"14",X"D0",X"03",X"E6",X"15",X"EA",X"E6",X"16",
		X"AD",X"00",X"40",X"6D",X"01",X"40",X"65",X"16",X"85",X"16",X"85",X"F5",X"EA",X"AD",X"03",X"40",
		X"30",X"FB",X"20",X"E6",X"C8",X"20",X"7B",X"D1",X"20",X"96",X"D7",X"20",X"98",X"D8",X"A5",X"1B",
		X"F0",X"0C",X"20",X"28",X"DB",X"20",X"BB",X"DB",X"20",X"77",X"DC",X"85",X"F5",X"EA",X"20",X"65",
		X"DD",X"20",X"8D",X"EA",X"20",X"DF",X"E6",X"20",X"41",X"E1",X"20",X"90",X"E1",X"20",X"35",X"E8",
		X"20",X"60",X"E7",X"20",X"6C",X"E8",X"A6",X"1F",X"B5",X"2B",X"D0",X"2D",X"A5",X"13",X"29",X"3F",
		X"D0",X"19",X"A2",X"FC",X"A0",X"C0",X"20",X"BC",X"C9",X"4C",X"19",X"C1",X"3A",X"10",X"00",X"00",
		X"00",X"FF",X"3A",X"10",X"51",X"52",X"53",X"FF",X"85",X"F6",X"EA",X"C9",X"0F",X"D0",X"0A",X"A2",
		X"02",X"A0",X"C1",X"20",X"BC",X"C9",X"85",X"F6",X"EA",X"A5",X"C6",X"D0",X"0D",X"A5",X"C5",X"F0",
		X"03",X"4C",X"75",X"C0",X"4C",X"7B",X"C0",X"85",X"F7",X"EA",X"A9",X"00",X"85",X"C6",X"C9",X"1B",
		X"D0",X"0B",X"A2",X"3F",X"20",X"2C",X"CA",X"4C",X"38",X"C0",X"85",X"F7",X"6E",X"20",X"A3",X"C8",
		X"20",X"E3",X"CB",X"A5",X"21",X"D0",X"17",X"A5",X"29",X"30",X"0D",X"A9",X"01",X"85",X"20",X"08",
		X"52",X"C2",X"4C",X"75",X"C0",X"85",X"F5",X"6E",X"4C",X"F1",X"C1",X"85",X"F7",X"6E",X"A6",X"1F",
		X"D0",X"4D",X"A5",X"29",X"25",X"2A",X"30",X"41",X"A5",X"2A",X"10",X"0D",X"20",X"6D",X"C2",X"A9",
		X"01",X"85",X"20",X"4C",X"75",X"C0",X"85",X"F7",X"EA",X"A5",X"29",X"10",X"09",X"20",X"95",X"C2",
		X"20",X"A3",X"C8",X"85",X"F7",X"6E",X"20",X"03",X"C3",X"A9",X"01",X"85",X"1F",X"C1",X"20",X"CD",
		X"03",X"40",X"29",X"40",X"F0",X"0D",X"A9",X"00",X"8D",X"05",X"50",X"A9",X"01",X"8D",X"02",X"40",
		X"85",X"F7",X"EA",X"20",X"81",X"C2",X"4C",X"75",X"C0",X"4C",X"F1",X"C1",X"85",X"F7",X"6E",X"A5",
		X"2A",X"25",X"29",X"30",X"3C",X"A5",X"29",X"10",X"0D",X"A9",X"01",X"85",X"20",X"08",X"81",X"C2",
		X"4C",X"75",X"C0",X"85",X"F7",X"6E",X"A5",X"2A",X"10",X"09",X"20",X"AD",X"C2",X"20",X"A3",X"C8",
		X"85",X"F7",X"EA",X"20",X"03",X"C3",X"A9",X"00",X"85",X"1F",X"A9",X"01",X"85",X"20",X"4D",X"FE",
		X"8D",X"05",X"50",X"A9",X"00",X"8D",X"02",X"40",X"20",X"6D",X"C2",X"4C",X"75",X"C0",X"85",X"F7",
		X"EA",X"20",X"C5",X"C2",X"20",X"A3",X"C8",X"A9",X"FE",X"8D",X"05",X"50",X"4D",X"00",X"8D",X"02",
		X"40",X"A9",X"00",X"85",X"CB",X"A5",X"2D",X"85",X"CC",X"A5",X"2E",X"85",X"CD",X"A5",X"2F",X"85",
		X"CE",X"20",X"F3",X"EF",X"20",X"A3",X"C8",X"AD",X"03",X"40",X"29",X"40",X"F0",X"0D",X"A9",X"00",
		X"8D",X"05",X"50",X"A9",X"01",X"8D",X"02",X"40",X"85",X"F7",X"EA",X"A9",X"01",X"85",X"CB",X"A5",
		X"30",X"85",X"CC",X"A5",X"31",X"85",X"CD",X"A5",X"32",X"85",X"CE",X"20",X"F3",X"EF",X"A2",X"00",
		X"86",X"1B",X"A5",X"1D",X"05",X"1E",X"F0",X"05",X"E6",X"1A",X"85",X"F7",X"EA",X"4C",X"38",X"C0",
		X"85",X"F7",X"EA",X"A2",X"E8",X"A0",X"C2",X"20",X"BC",X"C9",X"85",X"F5",X"EA",X"A9",X"03",X"20",
		X"5D",X"EA",X"85",X"F5",X"EA",X"A2",X"1F",X"20",X"2C",X"CA",X"60",X"85",X"F7",X"EA",X"A2",X"D2",
		X"A0",X"C2",X"20",X"BC",X"C9",X"A2",X"E8",X"A0",X"C2",X"20",X"BC",X"C9",X"4C",X"5D",X"C2",X"85",
		X"F7",X"EA",X"A2",X"DD",X"A0",X"C2",X"20",X"BC",X"C9",X"A2",X"E8",X"A0",X"C2",X"20",X"BC",X"C9",
		X"4C",X"5D",X"C2",X"85",X"F7",X"EA",X"E6",X"C8",X"A2",X"D2",X"A0",X"C2",X"20",X"BC",X"C9",X"E6",
		X"C8",X"A2",X"F5",X"A0",X"C2",X"20",X"BC",X"C9",X"4C",X"65",X"C2",X"85",X"F7",X"EA",X"E6",X"C8",
		X"A2",X"DD",X"A0",X"C2",X"20",X"BC",X"C9",X"E6",X"C8",X"A2",X"F5",X"A0",X"C2",X"20",X"BC",X"C9",
		X"4C",X"65",X"C2",X"85",X"F7",X"EA",X"E6",X"C8",X"A2",X"F5",X"A0",X"C2",X"20",X"BC",X"C9",X"4C",
		X"65",X"C2",X"CD",X"11",X"1A",X"16",X"0B",X"23",X"0F",X"1C",X"00",X"02",X"FF",X"CD",X"11",X"1A",
		X"16",X"0B",X"23",X"0F",X"1C",X"00",X"03",X"FF",X"0C",X"12",X"11",X"0B",X"17",X"0F",X"00",X"1C",
		X"0F",X"0B",X"0E",X"23",X"FF",X"0C",X"12",X"11",X"0B",X"17",X"0F",X"00",X"19",X"20",X"0F",X"1C",
		X"FF",X"85",X"F7",X"EA",X"A0",X"00",X"85",X"F7",X"EA",X"B9",X"00",X"02",X"AA",X"B9",X"00",X"03",
		X"99",X"00",X"02",X"8A",X"99",X"00",X"03",X"64",X"D0",X"EF",X"60",X"85",X"F6",X"6E",X"A9",X"00",
		X"8D",X"05",X"50",X"85",X"25",X"C5",X"03",X"40",X"A9",X"80",X"85",X"27",X"C5",X"00",X"40",X"28",
		X"85",X"F6",X"EA",X"85",X"F6",X"6E",X"A9",X"00",X"85",X"03",X"A9",X"10",X"85",X"04",X"4A",X"10",
		X"85",X"F6",X"EA",X"A0",X"00",X"85",X"F6",X"6E",X"A9",X"00",X"91",X"03",X"64",X"D0",X"F9",X"E6",
		X"04",X"CA",X"D0",X"EF",X"85",X"F6",X"6E",X"95",X"01",X"E8",X"E0",X"E1",X"D0",X"F9",X"A2",X"00",
		X"85",X"F6",X"EA",X"9D",X"00",X"02",X"D5",X"00",X"03",X"E8",X"D0",X"F7",X"A9",X"02",X"85",X"35",
		X"A9",X"80",X"85",X"34",X"4D",X"00",X"85",X"33",X"A2",X"23",X"85",X"F6",X"6E",X"BD",X"B3",X"C3",
		X"95",X"36",X"CA",X"10",X"F8",X"85",X"F6",X"6E",X"A0",X"00",X"85",X"F6",X"6E",X"A2",X"00",X"85",
		X"F6",X"EA",X"BD",X"A3",X"C3",X"99",X"00",X"0C",X"C8",X"E8",X"E0",X"10",X"D0",X"F4",X"C0",X"20",
		X"D0",X"EB",X"60",X"FF",X"00",X"D0",X"C0",X"F8",X"C7",X"E1",X"D4",X"FF",X"52",X"07",X"3F",X"00",
		X"F8",X"C0",X"38",X"00",X"80",X"02",X"00",X"01",X"01",X"00",X"94",X"00",X"50",X"65",X"00",X"50",
		X"48",X"00",X"FF",X"FF",X"FF",X"15",X"0F",X"18",X"12",X"CD",X"13",X"11",X"19",X"18",X"12",X"CD",
		X"15",X"15",X"CD",X"12",X"FF",X"FF",X"FF",X"85",X"F5",X"EA",X"20",X"A3",X"C8",X"20",X"E3",X"CB",
		X"A2",X"0F",X"A0",X"CE",X"20",X"BC",X"C9",X"A2",X"29",X"A0",X"CE",X"20",X"BC",X"C9",X"A2",X"BE",
		X"A0",X"CE",X"20",X"BC",X"C9",X"A6",X"5B",X"E8",X"8E",X"D5",X"12",X"A5",X"5A",X"29",X"F0",X"4A",
		X"4A",X"4A",X"4A",X"AA",X"E8",X"8E",X"D6",X"12",X"A2",X"01",X"8E",X"D7",X"12",X"8E",X"D8",X"12",
		X"8E",X"D9",X"12",X"60",X"85",X"F5",X"EA",X"20",X"A3",X"C8",X"20",X"E3",X"CB",X"A2",X"0F",X"A0",
		X"CE",X"20",X"BC",X"C9",X"A2",X"EF",X"A0",X"CE",X"20",X"BC",X"C9",X"A9",X"C9",X"85",X"03",X"A9",
		X"11",X"85",X"04",X"A2",X"12",X"85",X"F5",X"EA",X"A0",X"00",X"B5",X"36",X"91",X"03",X"C8",X"B5",
		X"37",X"91",X"03",X"C8",X"B5",X"38",X"91",X"03",X"18",X"A5",X"03",X"69",X"40",X"85",X"03",X"A5",
		X"04",X"69",X"00",X"85",X"04",X"E8",X"E8",X"E8",X"E0",X"21",X"90",X"DC",X"A2",X"03",X"20",X"4E",
		X"C9",X"A2",X"04",X"20",X"4E",X"C9",X"A2",X"05",X"20",X"4E",X"C9",X"A2",X"06",X"20",X"4E",X"C9",
		X"A2",X"07",X"20",X"4E",X"C9",X"60",X"85",X"F5",X"EA",X"A9",X"FF",X"85",X"19",X"85",X"F5",X"EA",
		X"A9",X"01",X"85",X"1C",X"20",X"48",X"C7",X"20",X"67",X"C7",X"A0",X"01",X"84",X"68",X"C8",X"84",
		X"69",X"C8",X"84",X"6A",X"A9",X"90",X"8D",X"02",X"18",X"A9",X"4D",X"8D",X"03",X"18",X"A9",X"60",
		X"8D",X"06",X"18",X"A9",X"3D",X"8D",X"07",X"18",X"A9",X"30",X"8D",X"0A",X"18",X"A9",X"3D",X"8D",
		X"0B",X"18",X"A9",X"40",X"85",X"A9",X"85",X"AA",X"85",X"AB",X"85",X"B0",X"A9",X"04",X"85",X"A8",
		X"85",X"BA",X"A9",X"18",X"8D",X"1E",X"18",X"A9",X"1D",X"8D",X"1F",X"18",X"20",X"65",X"DD",X"85",
		X"F5",X"EA",X"A2",X"01",X"20",X"2C",X"CA",X"E6",X"13",X"A2",X"07",X"20",X"C3",X"D3",X"F0",X"04",
		X"60",X"85",X"F5",X"EA",X"A2",X"07",X"20",X"69",X"D2",X"20",X"98",X"D8",X"20",X"8D",X"EA",X"20",
		X"90",X"E1",X"A5",X"19",X"D0",X"06",X"4C",X"D2",X"C4",X"85",X"F5",X"EA",X"A2",X"0F",X"A0",X"C5",
		X"20",X"BC",X"C9",X"A2",X"FF",X"20",X"2C",X"CA",X"A9",X"00",X"85",X"19",X"A4",X"80",X"C4",X"86",
		X"11",X"3B",X"40",X"60",X"36",X"3D",X"42",X"00",X"32",X"3D",X"35",X"61",X"62",X"FE",X"86",X"15",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"CE",X"10",X"3B",
		X"40",X"60",X"3E",X"37",X"31",X"39",X"3A",X"33",X"61",X"62",X"FE",X"CE",X"14",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"56",X"11",X"3B",X"40",X"60",X"33",X"35",
		X"35",X"61",X"62",X"FE",X"56",X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"85",
		X"F5",X"EA",X"20",X"48",X"C7",X"20",X"67",X"C7",X"A0",X"01",X"84",X"68",X"C0",X"69",X"64",X"84",
		X"6A",X"84",X"6B",X"C8",X"84",X"6C",X"C0",X"6D",X"A9",X"1D",X"8D",X"03",X"18",X"C5",X"07",X"18",
		X"8D",X"0B",X"18",X"8D",X"0F",X"18",X"C5",X"13",X"18",X"8D",X"17",X"18",X"C5",X"1F",X"18",X"4D",
		X"40",X"85",X"A9",X"85",X"AA",X"C1",X"AB",X"C1",X"AC",X"85",X"AD",X"85",X"AE",X"4D",X"89",X"8D",
		X"02",X"18",X"A9",X"59",X"8D",X"06",X"18",X"4D",X"60",X"8D",X"0A",X"18",X"4D",X"90",X"8D",X"0E",
		X"18",X"A9",X"97",X"8D",X"12",X"18",X"4D",X"30",X"8D",X"16",X"18",X"A9",X"18",X"8D",X"1E",X"18",
		X"A9",X"01",X"85",X"13",X"C1",X"14",X"08",X"65",X"DD",X"85",X"F5",X"EA",X"A2",X"01",X"20",X"2C",
		X"CA",X"E6",X"13",X"D0",X"03",X"E6",X"14",X"6E",X"A2",X"07",X"20",X"C3",X"D3",X"F0",X"1B",X"A5",
		X"14",X"C9",X"04",X"90",X"3C",X"A2",X"30",X"A0",X"C6",X"20",X"BC",X"C9",X"A2",X"FF",X"20",X"2C",
		X"CA",X"A2",X"40",X"20",X"2C",X"CA",X"60",X"85",X"F5",X"EA",X"A5",X"6E",X"10",X"23",X"A2",X"07",
		X"20",X"69",X"D2",X"AD",X"1E",X"18",X"C9",X"22",X"F0",X"0B",X"C9",X"4A",X"F0",X"07",X"C9",X"82",
		X"D0",X"0F",X"85",X"F5",X"EA",X"20",X"AD",X"D1",X"EE",X"1E",X"18",X"EE",X"1E",X"18",X"85",X"F5",
		X"EA",X"20",X"96",X"D7",X"20",X"98",X"D8",X"20",X"DF",X"E6",X"20",X"90",X"E1",X"4C",X"CC",X"C5",
		X"C7",X"10",X"32",X"3D",X"3C",X"64",X"42",X"00",X"45",X"2F",X"41",X"42",X"33",X"00",X"3E",X"33",
		X"3E",X"3E",X"33",X"40",X"41",X"FE",X"C7",X"14",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"04",X"11",X"47",X"3D",
		X"43",X"00",X"41",X"42",X"2F",X"40",X"42",X"00",X"45",X"37",X"42",X"36",X"00",X"3D",X"3C",X"3A",
		X"47",X"00",X"34",X"37",X"44",X"33",X"FE",X"04",X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FE",X"42",X"11",X"33",X"2F",X"40",X"3C",X"00",X"33",X"46",X"42",X"40",X"2F",X"00",X"3E",
		X"33",X"3E",X"3E",X"33",X"40",X"41",X"00",X"63",X"00",X"30",X"3D",X"3C",X"43",X"41",X"33",X"41",
		X"FE",X"42",X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",
		X"83",X"11",X"31",X"3A",X"2F",X"37",X"3B",X"00",X"31",X"3D",X"3C",X"33",X"41",X"4A",X"31",X"3D",
		X"34",X"34",X"33",X"33",X"41",X"00",X"63",X"00",X"34",X"40",X"37",X"33",X"41",X"FE",X"83",X"15",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"85",X"F5",X"6E",X"AD",X"04",
		X"40",X"49",X"FF",X"A8",X"A2",X"02",X"29",X"01",X"F0",X"05",X"A2",X"04",X"85",X"F5",X"6E",X"86",
		X"29",X"86",X"2A",X"98",X"4A",X"29",X"03",X"AA",X"BD",X"3E",X"C7",X"85",X"5A",X"C1",X"5C",X"C1",
		X"5E",X"BD",X"42",X"C7",X"85",X"5B",X"C1",X"5D",X"85",X"5F",X"20",X"C3",X"EB",X"60",X"00",X"50",
		X"00",X"00",X"01",X"01",X"02",X"03",X"85",X"F7",X"EA",X"A9",X"01",X"85",X"61",X"C1",X"62",X"4D",
		X"04",X"20",X"5D",X"EA",X"A9",X"00",X"85",X"65",X"85",X"66",X"85",X"1F",X"08",X"0F",X"CC",X"20",
		X"03",X"C3",X"C6",X"61",X"28",X"85",X"F5",X"6E",X"20",X"A3",X"C8",X"A5",X"20",X"D0",X"2C",X"A9",
		X"04",X"20",X"5D",X"EA",X"AD",X"04",X"40",X"29",X"10",X"D0",X"12",X"A5",X"1B",X"F0",X"0E",X"A6",
		X"1F",X"B5",X"2B",X"18",X"F8",X"69",X"01",X"95",X"2B",X"D8",X"85",X"F6",X"6E",X"A6",X"1F",X"F6",
		X"61",X"A9",X"00",X"95",X"65",X"08",X"0F",X"CC",X"85",X"F5",X"EA",X"A9",X"00",X"85",X"20",X"08",
		X"64",X"CC",X"A6",X"1F",X"B4",X"61",X"88",X"85",X"F5",X"EA",X"C0",X"06",X"90",X"0B",X"98",X"38",
		X"E9",X"06",X"A8",X"4C",X"AA",X"C7",X"85",X"F5",X"EA",X"84",X"63",X"B4",X"61",X"88",X"C0",X"06",
		X"90",X"05",X"A0",X"05",X"85",X"F5",X"6E",X"84",X"64",X"A4",X"63",X"B9",X"EF",X"CD",X"8D",X"1C",
		X"18",X"B9",X"F7",X"CD",X"8D",X"1D",X"18",X"5D",X"FF",X"CD",X"8D",X"1E",X"18",X"5D",X"07",X"CE",
		X"8D",X"1F",X"18",X"A2",X"07",X"A9",X"FF",X"85",X"F5",X"EA",X"95",X"68",X"66",X"10",X"FB",X"A2",
		X"07",X"A9",X"01",X"85",X"F5",X"6E",X"95",X"99",X"CA",X"10",X"FB",X"A2",X"07",X"A9",X"04",X"85",
		X"F5",X"EA",X"95",X"A1",X"CA",X"10",X"FB",X"A2",X"07",X"A9",X"00",X"85",X"F5",X"EA",X"95",X"A9",
		X"CA",X"10",X"FB",X"85",X"6F",X"A9",X"03",X"85",X"A8",X"A9",X"00",X"85",X"C5",X"85",X"C4",X"20",
		X"89",X"DA",X"20",X"C6",X"C8",X"A5",X"21",X"F0",X"0B",X"A5",X"1F",X"49",X"01",X"AA",X"20",X"4E",
		X"C9",X"85",X"F5",X"EA",X"A6",X"1F",X"20",X"4E",X"C9",X"A2",X"02",X"20",X"4E",X"C9",X"20",X"54",
		X"CA",X"20",X"94",X"CA",X"A6",X"1F",X"20",X"C4",X"CA",X"20",X"1E",X"CB",X"A9",X"3E",X"85",X"13",
		X"A5",X"1B",X"F0",X"04",X"60",X"85",X"F5",X"EA",X"A9",X"01",X"85",X"68",X"A9",X"02",X"85",X"69",
		X"A9",X"03",X"85",X"6A",X"A9",X"90",X"8D",X"02",X"18",X"A9",X"4D",X"8D",X"03",X"18",X"A9",X"60",
		X"8D",X"06",X"18",X"A9",X"3D",X"8D",X"07",X"18",X"A9",X"30",X"8D",X"0A",X"18",X"A9",X"3D",X"8D",
		X"0B",X"18",X"A9",X"80",X"85",X"A9",X"85",X"AA",X"85",X"AB",X"A9",X"40",X"85",X"B0",X"A9",X"18",
		X"8D",X"1E",X"18",X"A9",X"1D",X"8D",X"1F",X"18",X"A9",X"FF",X"85",X"A1",X"85",X"A2",X"85",X"A3",
		X"60",X"85",X"F6",X"EA",X"A0",X"00",X"84",X"03",X"A9",X"10",X"85",X"04",X"85",X"F6",X"EA",X"A9",
		X"00",X"91",X"03",X"C8",X"D0",X"F9",X"E6",X"04",X"A5",X"04",X"C9",X"18",X"D0",X"F1",X"A2",X"01",
		X"20",X"2C",X"CA",X"60",X"85",X"F5",X"EA",X"A2",X"35",X"A0",X"C9",X"20",X"BC",X"C9",X"A2",X"29",
		X"A0",X"C9",X"20",X"BC",X"C9",X"A5",X"21",X"F0",X"0A",X"A2",X"40",X"A0",X"C9",X"20",X"BC",X"C9",
		X"85",X"F5",X"EA",X"60",X"85",X"F5",X"EA",X"A5",X"21",X"F0",X"3D",X"A5",X"13",X"29",X"3F",X"D0",
		X"1A",X"A5",X"1F",X"D0",X"0B",X"A2",X"2F",X"A0",X"C9",X"20",X"BC",X"C9",X"60",X"85",X"F5",X"EA",
		X"A2",X"46",X"A0",X"C9",X"20",X"BC",X"C9",X"60",X"85",X"F5",X"EA",X"C9",X"0F",X"D0",X"19",X"A5",
		X"1F",X"D0",X"0B",X"A2",X"29",X"A0",X"C9",X"20",X"BC",X"C9",X"60",X"85",X"F5",X"6E",X"A2",X"40",
		X"A0",X"C9",X"20",X"BC",X"C9",X"85",X"F5",X"6E",X"60",X"24",X"10",X"26",X"43",X"3E",X"FF",X"24",
		X"10",X"00",X"00",X"00",X"FF",X"29",X"10",X"36",X"37",X"49",X"41",X"31",X"3D",X"40",X"33",X"FF",
		X"34",X"10",X"27",X"43",X"3E",X"FF",X"34",X"10",X"00",X"00",X"00",X"FF",X"85",X"F5",X"6E",X"86",
		X"03",X"8A",X"0A",X"A8",X"18",X"65",X"03",X"AA",X"85",X"F5",X"EA",X"B9",X"A0",X"C9",X"85",X"03",
		X"B9",X"A1",X"C9",X"85",X"04",X"48",X"05",X"85",X"F5",X"EA",X"B5",X"2D",X"29",X"0F",X"85",X"05",
		X"E6",X"05",X"A5",X"05",X"91",X"03",X"44",X"B5",X"2D",X"4A",X"4A",X"4A",X"4A",X"85",X"05",X"EA",
		X"05",X"A5",X"05",X"91",X"03",X"6C",X"88",X"10",X"E1",X"C8",X"85",X"F5",X"6E",X"B1",X"03",X"C9",
		X"01",X"D0",X"0C",X"A9",X"00",X"91",X"03",X"64",X"C0",X"05",X"D0",X"F1",X"85",X"F5",X"6E",X"60",
		X"42",X"10",X"52",X"10",X"4A",X"10",X"CD",X"11",X"0D",X"12",X"4D",X"12",X"8D",X"12",X"CD",X"12",
		X"92",X"12",X"D2",X"12",X"12",X"13",X"52",X"13",X"92",X"13",X"85",X"F6",X"6E",X"86",X"03",X"C0",
		X"04",X"85",X"F6",X"EA",X"A0",X"00",X"84",X"08",X"B1",X"03",X"85",X"05",X"64",X"B1",X"03",X"85",
		X"06",X"85",X"F6",X"EA",X"C8",X"B1",X"03",X"C9",X"FF",X"F0",X"4A",X"C9",X"FE",X"F0",X"1D",X"C9",
		X"FD",X"F0",X"2C",X"84",X"07",X"C8",X"08",X"91",X"05",X"E6",X"08",X"A4",X"07",X"A5",X"C8",X"F0",
		X"E3",X"A2",X"0A",X"20",X"2C",X"CA",X"4C",X"D4",X"C9",X"85",X"F6",X"EA",X"C8",X"18",X"98",X"65",
		X"03",X"85",X"03",X"A5",X"04",X"69",X"00",X"85",X"04",X"4C",X"C4",X"C9",X"85",X"F6",X"EA",X"18",
		X"A5",X"05",X"69",X"20",X"85",X"05",X"A5",X"06",X"69",X"00",X"85",X"06",X"A9",X"00",X"85",X"08",
		X"F0",X"B2",X"85",X"F6",X"EA",X"A9",X"00",X"85",X"C8",X"60",X"85",X"F6",X"EA",X"AD",X"03",X"40",
		X"10",X"FB",X"58",X"EA",X"EA",X"EA",X"EA",X"78",X"20",X"45",X"D0",X"A5",X"1A",X"F0",X"0A",X"8A",
		X"48",X"20",X"6E",X"D0",X"68",X"AA",X"85",X"F6",X"EA",X"AD",X"03",X"40",X"30",X"FB",X"CA",X"D0",
		X"DC",X"60",X"85",X"F5",X"EA",X"A6",X"1F",X"38",X"A9",X"5C",X"F5",X"29",X"85",X"F3",X"A9",X"18",
		X"85",X"F4",X"B5",X"29",X"C9",X"09",X"B0",X"16",X"A0",X"10",X"A9",X"00",X"99",X"4C",X"18",X"88",
		X"D0",X"FA",X"B4",X"29",X"F0",X"07",X"A9",X"C8",X"91",X"F3",X"88",X"D0",X"FB",X"60",X"A0",X"09",
		X"A9",X"53",X"85",X"F3",X"4C",X"76",X"CA",X"F6",X"EA",X"91",X"F3",X"88",X"D0",X"FB",X"85",X"F7",
		X"EA",X"60",X"85",X"F5",X"EA",X"98",X"48",X"A0",X"51",X"8C",X"3A",X"10",X"C8",X"8C",X"3B",X"10",
		X"C8",X"8C",X"3C",X"10",X"A6",X"1F",X"B5",X"2B",X"4A",X"4A",X"4A",X"4A",X"A8",X"F0",X"04",X"C8",
		X"85",X"F5",X"EA",X"8C",X"5B",X"10",X"B5",X"2B",X"29",X"0F",X"A8",X"C8",X"8C",X"5C",X"10",X"68",
		X"A8",X"60",X"85",X"F5",X"EA",X"B5",X"61",X"85",X"03",X"AD",X"1A",X"CB",X"85",X"04",X"AD",X"1B",
		X"CB",X"85",X"05",X"A9",X"04",X"85",X"06",X"A0",X"80",X"85",X"F5",X"EA",X"A6",X"03",X"E0",X"0A",
		X"90",X"0D",X"A5",X"03",X"E9",X"0A",X"85",X"03",X"A9",X"C6",X"D0",X"1F",X"85",X"F5",X"EA",X"E0",
		X"05",X"90",X"0D",X"A5",X"03",X"E9",X"05",X"85",X"03",X"A9",X"C5",X"D0",X"0E",X"85",X"F5",X"EA",
		X"E0",X"01",X"90",X"15",X"C6",X"03",X"4D",X"C4",X"85",X"F5",X"EA",X"91",X"04",X"54",X"38",X"E9",
		X"20",X"A8",X"C6",X"06",X"10",X"C6",X"85",X"F5",X"EA",X"60",X"1D",X"13",X"85",X"F5",X"6E",X"20",
		X"E3",X"CB",X"A5",X"63",X"0A",X"A8",X"B9",X"D7",X"CD",X"85",X"03",X"B9",X"D8",X"CD",X"85",X"04",
		X"A9",X"10",X"85",X"05",X"4D",X"04",X"85",X"06",X"A2",X"68",X"A0",X"00",X"85",X"F5",X"6E",X"B1",
		X"03",X"29",X"F0",X"11",X"05",X"91",X"05",X"EA",X"05",X"B1",X"03",X"0A",X"0A",X"0A",X"0A",X"11",
		X"05",X"91",X"05",X"E6",X"05",X"EA",X"03",X"70",X"05",X"E6",X"04",X"85",X"F5",X"6E",X"CA",X"A5",
		X"05",X"29",X"07",X"D0",X"DA",X"18",X"A5",X"05",X"69",X"7F",X"85",X"05",X"C9",X"06",X"69",X"00",
		X"85",X"06",X"85",X"F5",X"6E",X"B1",X"03",X"29",X"F0",X"11",X"05",X"91",X"05",X"E2",X"05",X"59",
		X"03",X"0A",X"0A",X"0A",X"0A",X"11",X"05",X"91",X"05",X"C6",X"05",X"E6",X"03",X"70",X"05",X"E6",
		X"04",X"85",X"F5",X"EA",X"CA",X"A5",X"05",X"29",X"07",X"C9",X"07",X"D0",X"D8",X"38",X"A5",X"05",
		X"E9",X"77",X"85",X"05",X"C9",X"06",X"E9",X"00",X"85",X"06",X"E0",X"00",X"D0",X"91",X"A5",X"63",
		X"29",X"0F",X"85",X"F3",X"46",X"48",X"CD",X"03",X"40",X"29",X"40",X"F0",X"07",X"A5",X"1F",X"D0",
		X"13",X"85",X"F5",X"EA",X"A6",X"F3",X"BD",X"D9",X"CB",X"09",X"10",X"8D",X"04",X"40",X"2C",X"AA",
		X"60",X"85",X"F5",X"EA",X"A5",X"F3",X"4C",X"C9",X"CB",X"03",X"00",X"01",X"02",X"07",X"04",X"05",
		X"06",X"85",X"F5",X"EA",X"A0",X"00",X"A9",X"04",X"85",X"04",X"A9",X"00",X"85",X"03",X"C1",X"F5",
		X"EA",X"B1",X"03",X"29",X"0F",X"91",X"03",X"64",X"D0",X"F7",X"E6",X"04",X"CA",X"04",X"E0",X"08",
		X"D0",X"EF",X"A9",X"00",X"8D",X"04",X"40",X"A2",X"01",X"20",X"2C",X"CA",X"60",X"85",X"F5",X"EA",
		X"A6",X"1F",X"B4",X"61",X"88",X"85",X"F5",X"EA",X"C0",X"06",X"90",X"0B",X"98",X"38",X"E9",X"06",
		X"A8",X"4C",X"18",X"CC",X"85",X"F5",X"EA",X"98",X"0A",X"A8",X"B9",X"E3",X"CD",X"85",X"03",X"B9",
		X"E4",X"CD",X"85",X"04",X"A0",X"00",X"A2",X"00",X"85",X"F5",X"EA",X"B1",X"03",X"C9",X"FF",X"F0",
		X"18",X"9D",X"02",X"02",X"C8",X"E8",X"8A",X"29",X"03",X"C9",X"03",X"D0",X"EE",X"E8",X"A9",X"00",
		X"9D",X"02",X"02",X"4C",X"3B",X"CC",X"85",X"F5",X"EA",X"A9",X"00",X"9D",X"02",X"02",X"E8",X"D0",
		X"F8",X"60",X"85",X"F7",X"EA",X"A9",X"02",X"85",X"0B",X"A9",X"02",X"85",X"0C",X"A9",X"00",X"85",
		X"0D",X"85",X"F7",X"EA",X"A4",X"0D",X"B1",X"0B",X"F0",X"1C",X"85",X"03",X"C8",X"B1",X"0B",X"85",
		X"04",X"C8",X"B1",X"0B",X"85",X"05",X"20",X"99",X"CC",X"A5",X"0D",X"18",X"69",X"04",X"85",X"0D",
		X"4C",X"74",X"CC",X"85",X"F7",X"EA",X"60",X"85",X"F5",X"EA",X"A9",X"00",X"85",X"0E",X"F0",X"12",
		X"85",X"F5",X"EA",X"A9",X"00",X"85",X"0E",X"A5",X"05",X"29",X"F8",X"D0",X"05",X"E6",X"0E",X"85",
		X"F5",X"EA",X"98",X"48",X"A5",X"03",X"29",X"0F",X"0A",X"AA",X"BD",X"B7",X"CD",X"85",X"07",X"A5",
		X"05",X"29",X"07",X"0A",X"0A",X"18",X"65",X"07",X"85",X"07",X"BD",X"B8",X"CD",X"85",X"08",X"A5",
		X"04",X"49",X"FF",X"85",X"04",X"46",X"04",X"46",X"04",X"46",X"04",X"A9",X"00",X"85",X"06",X"A5",
		X"05",X"29",X"F8",X"85",X"05",X"06",X"05",X"26",X"06",X"06",X"05",X"26",X"06",X"18",X"A5",X"05",
		X"65",X"04",X"85",X"05",X"A5",X"06",X"69",X"10",X"85",X"06",X"A5",X"03",X"29",X"0F",X"C9",X"0F",
		X"F0",X"35",X"A0",X"00",X"A5",X"07",X"AA",X"20",X"95",X"CD",X"A4",X"0E",X"D0",X"0C",X"A0",X"20",
		X"18",X"69",X"1D",X"AA",X"20",X"95",X"CD",X"85",X"F5",X"EA",X"18",X"A5",X"06",X"69",X"04",X"85",
		X"06",X"A0",X"00",X"A5",X"08",X"20",X"AA",X"CD",X"A4",X"0E",X"D0",X"64",X"A0",X"20",X"20",X"AA",
		X"CD",X"4C",X"90",X"CD",X"85",X"F5",X"6E",X"38",X"A5",X"05",X"E9",X"21",X"85",X"05",X"C9",X"06",
		X"E9",X"00",X"85",X"06",X"48",X"00",X"A5",X"07",X"91",X"05",X"AA",X"E8",X"E8",X"8A",X"A0",X"05",
		X"91",X"05",X"E6",X"07",X"C9",X"07",X"A0",X"21",X"91",X"05",X"C8",X"91",X"05",X"64",X"91",X"05",
		X"C8",X"91",X"05",X"18",X"A5",X"06",X"69",X"04",X"85",X"06",X"A0",X"21",X"A9",X"00",X"91",X"05",
		X"C8",X"91",X"05",X"C8",X"91",X"05",X"64",X"91",X"05",X"38",X"A5",X"06",X"E9",X"04",X"85",X"06",
		X"18",X"A5",X"05",X"69",X"21",X"85",X"05",X"C9",X"06",X"69",X"00",X"85",X"06",X"C1",X"F5",X"6E",
		X"68",X"A8",X"60",X"85",X"F7",X"6E",X"91",X"05",X"C8",X"E8",X"8A",X"91",X"05",X"64",X"E8",X"8A",
		X"91",X"05",X"C8",X"E8",X"8A",X"91",X"05",X"28",X"85",X"F7",X"EA",X"91",X"05",X"64",X"91",X"05",
		X"C8",X"91",X"05",X"C8",X"91",X"05",X"28",X"00",X"00",X"00",X"02",X"40",X"02",X"80",X"02",X"C0",
		X"02",X"00",X"03",X"40",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"C9",X"00",X"81",X"ED",X"51",X"EE",X"B9",X"EE",X"21",X"EF",X"E9",
		X"ED",X"89",X"EF",X"D7",X"EB",X"4B",X"EC",X"88",X"EC",X"D1",X"EC",X"14",X"EC",X"3E",X"ED",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"47",X"47",X"47",X"47",X"47",X"47",X"47",X"47",X"78",
		X"78",X"78",X"78",X"48",X"78",X"78",X"78",X"AD",X"BD",X"CD",X"8D",X"CD",X"AD",X"AD",X"AD",X"AA",
		X"10",X"30",X"43",X"40",X"35",X"33",X"40",X"00",X"42",X"37",X"3B",X"33",X"FE",X"EB",X"10",X"4D",
		X"4E",X"4F",X"50",X"00",X"26",X"2E",X"2D",X"27",X"FF",X"2C",X"11",X"CC",X"1D",X"0D",X"19",X"1C",
		X"0F",X"CC",X"FE",X"65",X"11",X"00",X"01",X"02",X"03",X"00",X"00",X"40",X"41",X"42",X"43",X"00",
		X"00",X"80",X"81",X"82",X"83",X"FE",X"65",X"15",X"02",X"02",X"02",X"02",X"00",X"00",X"03",X"03",
		X"03",X"03",X"00",X"00",X"02",X"02",X"02",X"02",X"FE",X"A5",X"11",X"C0",X"C1",X"C2",X"C3",X"00",
		X"00",X"00",X"01",X"02",X"03",X"00",X"00",X"40",X"41",X"42",X"43",X"FE",X"A5",X"15",X"02",X"02",
		X"02",X"02",X"00",X"00",X"03",X"03",X"03",X"03",X"00",X"00",X"02",X"02",X"02",X"02",X"FE",X"E5",
		X"11",X"BC",X"BD",X"00",X"00",X"C0",X"C1",X"00",X"00",X"B8",X"B9",X"FE",X"05",X"12",X"BE",X"BF",
		X"00",X"00",X"C2",X"C3",X"00",X"00",X"BA",X"BB",X"FE",X"25",X"12",X"DC",X"DD",X"00",X"00",X"E0",
		X"E1",X"00",X"00",X"B4",X"B5",X"FE",X"96",X"11",X"06",X"01",X"00",X"1A",X"1E",X"1D",X"FE",X"10",
		X"12",X"CC",X"0C",X"19",X"18",X"1F",X"1D",X"00",X"02",X"00",X"51",X"52",X"53",X"FF",X"C3",X"12",
		X"0C",X"19",X"18",X"1F",X"1D",X"00",X"00",X"00",X"10",X"19",X"1C",X"00",X"0F",X"20",X"0F",X"1C",
		X"23",X"00",X"00",X"00",X"00",X"00",X"00",X"1A",X"1E",X"1D",X"FE",X"A8",X"12",X"1C",X"1D",X"FE",
		X"C8",X"12",X"1E",X"1F",X"FE",X"A8",X"16",X"01",X"01",X"FE",X"C8",X"16",X"01",X"01",X"FF",X"67",
		X"11",X"0C",X"0F",X"1D",X"1E",X"00",X"10",X"13",X"20",X"0F",X"00",X"1A",X"16",X"0B",X"23",X"0F",
		X"1C",X"1D",X"FE",X"C7",X"11",X"02",X"FE",X"D4",X"11",X"1A",X"1E",X"1D",X"FE",X"07",X"12",X"03",
		X"FE",X"14",X"12",X"1A",X"1E",X"1D",X"FE",X"47",X"12",X"04",X"FE",X"54",X"12",X"1A",X"1E",X"1D",
		X"FE",X"87",X"12",X"05",X"FE",X"94",X"12",X"1A",X"1E",X"1D",X"FE",X"C7",X"12",X"06",X"FE",X"D4",
		X"12",X"1A",X"1E",X"1D",X"FF",X"68",X"4C",X"00",X"B0",X"85",X"F5",X"EA",X"48",X"CD",X"03",X"40",
		X"29",X"10",X"F0",X"F1",X"8A",X"48",X"54",X"48",X"EA",X"D8",X"A5",X"01",X"F0",X"40",X"AD",X"04",
		X"40",X"49",X"FF",X"29",X"E0",X"85",X"02",X"26",X"4A",X"4A",X"4A",X"4A",X"A8",X"20",X"34",X"D0",
		X"AD",X"02",X"40",X"29",X"C0",X"F0",X"27",X"85",X"26",X"20",X"34",X"D0",X"AD",X"02",X"40",X"25",
		X"26",X"F0",X"1B",X"20",X"34",X"D0",X"AD",X"02",X"40",X"25",X"26",X"F0",X"11",X"20",X"34",X"D0",
		X"AD",X"02",X"40",X"25",X"26",X"F0",X"07",X"A9",X"01",X"85",X"F9",X"85",X"F6",X"6E",X"8D",X"00",
		X"40",X"68",X"A8",X"68",X"AA",X"68",X"40",X"85",X"F6",X"EA",X"E6",X"1E",X"4D",X"1B",X"8D",X"03",
		X"40",X"A5",X"02",X"C9",X"80",X"F0",X"31",X"A2",X"00",X"AD",X"03",X"40",X"49",X"FF",X"29",X"0F",
		X"06",X"26",X"90",X"05",X"4A",X"4A",X"85",X"F5",X"EA",X"29",X"03",X"F0",X"46",X"E8",X"C9",X"01",
		X"F0",X"41",X"E8",X"C9",X"02",X"F0",X"31",X"E8",X"85",X"F5",X"EA",X"A5",X"1E",X"C9",X"02",X"B0",
		X"1F",X"85",X"F5",X"EA",X"60",X"85",X"F5",X"6E",X"A2",X"05",X"A5",X"26",X"C9",X"80",X"F0",X"23",
		X"E8",X"C9",X"40",X"F0",X"1E",X"E8",X"C9",X"C0",X"F0",X"19",X"4C",X"D4",X"CF",X"85",X"F5",X"6E",
		X"C6",X"1E",X"4C",X"03",X"D0",X"85",X"F5",X"6E",X"A5",X"02",X"C9",X"60",X"D0",X"05",X"A2",X"04",
		X"85",X"F5",X"EA",X"A5",X"1D",X"F8",X"18",X"7D",X"5C",X"D0",X"D9",X"64",X"D0",X"90",X"06",X"B9",
		X"64",X"D0",X"85",X"F5",X"EA",X"85",X"1D",X"D8",X"C6",X"1E",X"A5",X"1B",X"D0",X"11",X"8D",X"00",
		X"40",X"A9",X"01",X"85",X"1A",X"A2",X"FF",X"9A",X"EA",X"4C",X"38",X"C0",X"85",X"F6",X"EA",X"4C",
		X"D4",X"CF",X"85",X"F5",X"EA",X"A2",X"E7",X"85",X"F5",X"EA",X"A5",X"FF",X"A5",X"FF",X"EA",X"CA",
		X"D0",X"F8",X"60",X"85",X"F6",X"EA",X"A5",X"F9",X"F0",X"11",X"AD",X"02",X"40",X"29",X"C0",X"D0",
		X"0A",X"A9",X"00",X"85",X"F9",X"20",X"99",X"CF",X"85",X"F6",X"EA",X"60",X"01",X"02",X"03",X"01",
		X"06",X"08",X"03",X"01",X"09",X"09",X"09",X"09",X"09",X"09",X"09",X"09",X"85",X"F5",X"EA",X"A5",
		X"1A",X"F0",X"1E",X"A5",X"1C",X"D0",X"09",X"20",X"11",X"D1",X"20",X"3F",X"D1",X"85",X"F5",X"EA",
		X"AD",X"02",X"40",X"29",X"01",X"F0",X"0E",X"AD",X"02",X"40",X"29",X"02",X"F0",X"32",X"85",X"F5",
		X"EA",X"60",X"85",X"F5",X"EA",X"20",X"6E",X"D1",X"A9",X"00",X"85",X"21",X"85",X"20",X"85",X"1C",
		X"A9",X"01",X"85",X"1B",X"A9",X"00",X"85",X"1A",X"20",X"A3",X"C8",X"20",X"E3",X"CB",X"A2",X"E8",
		X"A0",X"C2",X"20",X"BC",X"C9",X"A2",X"1F",X"20",X"2C",X"CA",X"4C",X"FD",X"D0",X"85",X"F5",X"EA",
		X"A5",X"1D",X"C9",X"02",X"B0",X"03",X"4C",X"91",X"D0",X"20",X"6E",X"D1",X"20",X"6E",X"D1",X"A9",
		X"01",X"85",X"21",X"A9",X"00",X"85",X"20",X"85",X"1C",X"A9",X"01",X"85",X"1B",X"A9",X"00",X"85",
		X"1A",X"20",X"A3",X"C8",X"20",X"E3",X"CB",X"A2",X"D2",X"A0",X"C2",X"20",X"BC",X"C9",X"A2",X"E8",
		X"A0",X"C2",X"20",X"BC",X"C9",X"A2",X"1F",X"20",X"2C",X"CA",X"85",X"F5",X"EA",X"A2",X"05",X"A9",
		X"00",X"85",X"F5",X"EA",X"95",X"2D",X"66",X"10",X"FB",X"A2",X"FF",X"9A",X"4C",X"68",X"C0",X"85",
		X"F5",X"EA",X"AD",X"67",X"13",X"CD",X"55",X"D1",X"F0",X"3A",X"A0",X"00",X"85",X"F5",X"6E",X"B9",
		X"55",X"D1",X"99",X"67",X"13",X"64",X"C0",X"11",X"D0",X"F5",X"85",X"F5",X"6E",X"A0",X"00",X"85",
		X"F5",X"EA",X"B9",X"66",X"D1",X"99",X"AB",X"13",X"C8",X"C0",X"06",X"D0",X"F5",X"85",X"F5",X"6E",
		X"A5",X"1D",X"4A",X"4A",X"4A",X"4A",X"AA",X"E8",X"A5",X"1D",X"29",X"0F",X"AA",X"E8",X"8E",X"B3",
		X"13",X"85",X"F5",X"EA",X"60",X"1A",X"1F",X"1D",X"12",X"00",X"1D",X"1E",X"0B",X"1C",X"1E",X"00",
		X"0C",X"1F",X"1E",X"1E",X"19",X"18",X"0D",X"1C",X"0F",X"0E",X"13",X"1E",X"85",X"F5",X"6E",X"F8",
		X"38",X"A5",X"1D",X"E9",X"01",X"85",X"1D",X"74",X"60",X"85",X"F5",X"EA",X"A5",X"6F",X"10",X"04",
		X"85",X"F5",X"EA",X"60",X"A5",X"1B",X"D0",X"03",X"4C",X"36",X"D2",X"A6",X"1F",X"A4",X"1F",X"AD",
		X"03",X"40",X"29",X"40",X"D0",X"02",X"A0",X"00",X"B9",X"00",X"40",X"49",X"FF",X"29",X"10",X"F0",
		X"40",X"A5",X"B9",X"D0",X"43",X"B5",X"2B",X"F0",X"2D",X"85",X"B9",X"85",X"F5",X"6E",X"A9",X"00",
		X"85",X"6E",X"A9",X"05",X"85",X"A0",X"C9",X"BA",X"AA",X"18",X"BD",X"4D",X"D2",X"6D",X"1E",X"18",
		X"8D",X"1A",X"18",X"18",X"BD",X"4E",X"D2",X"6D",X"1F",X"18",X"8D",X"1B",X"18",X"4D",X"0D",X"20",
		X"5D",X"EA",X"60",X"85",X"F5",X"6E",X"A9",X"0E",X"20",X"5D",X"EA",X"4C",X"E8",X"D1",X"85",X"F5",
		X"EA",X"A9",X"00",X"85",X"B9",X"C1",X"F5",X"6E",X"B9",X"00",X"40",X"49",X"FF",X"29",X"0F",X"A8",
		X"B9",X"57",X"D2",X"A8",X"C5",X"BB",X"F0",X"09",X"0A",X"0A",X"0A",X"0A",X"85",X"B0",X"C1",X"F5",
		X"EA",X"84",X"BB",X"98",X"F0",X"05",X"84",X"BA",X"85",X"F5",X"EA",X"A5",X"BB",X"F0",X"0A",X"A2",
		X"07",X"20",X"C3",X"D3",X"D0",X"1C",X"85",X"F5",X"EA",X"A2",X"07",X"20",X"69",X"D2",X"A5",X"B0",
		X"29",X"F0",X"F0",X"0E",X"A0",X"06",X"C9",X"60",X"B0",X"01",X"C8",X"98",X"20",X"5D",X"EA",X"85",
		X"F5",X"EA",X"60",X"85",X"F5",X"EA",X"A2",X"07",X"20",X"C3",X"D3",X"F0",X"0A",X"A9",X"47",X"8D",
		X"1D",X"18",X"E6",X"C6",X"85",X"F5",X"EA",X"A2",X"07",X"20",X"69",X"D2",X"60",X"00",X"10",X"F0",
		X"00",X"10",X"00",X"00",X"F0",X"00",X"10",X"00",X"02",X"04",X"00",X"06",X"00",X"00",X"00",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"85",X"F5",X"EA",X"B5",X"68",X"10",X"01",X"60",X"A5",
		X"13",X"35",X"91",X"D0",X"01",X"60",X"D6",X"99",X"F0",X"01",X"60",X"B5",X"A1",X"95",X"99",X"B5",
		X"A9",X"29",X"0F",X"85",X"03",X"B5",X"A9",X"4A",X"4A",X"4A",X"F0",X"0B",X"18",X"65",X"03",X"85",
		X"03",X"4C",X"AC",X"D2",X"85",X"F5",X"EA",X"E0",X"07",X"D0",X"11",X"A0",X"00",X"A5",X"BA",X"C9",
		X"06",X"D0",X"04",X"C8",X"85",X"F5",X"EA",X"84",X"03",X"85",X"F5",X"EA",X"8A",X"0A",X"0A",X"85",
		X"09",X"B5",X"68",X"29",X"07",X"0A",X"A8",X"B9",X"4B",X"D3",X"85",X"05",X"B9",X"4C",X"D3",X"85",
		X"06",X"A4",X"03",X"B1",X"05",X"C9",X"FF",X"F0",X"4B",X"A4",X"09",X"99",X"01",X"18",X"B5",X"A9",
		X"4A",X"4A",X"4A",X"4A",X"29",X"02",X"09",X"01",X"99",X"00",X"18",X"B5",X"A9",X"29",X"F0",X"F0",
		X"69",X"F6",X"A9",X"B5",X"A9",X"29",X"F3",X"95",X"A9",X"86",X"08",X"A4",X"09",X"4A",X"4A",X"4A",
		X"4A",X"AA",X"18",X"BD",X"B7",X"D3",X"79",X"02",X"18",X"99",X"02",X"18",X"18",X"BD",X"B8",X"D3",
		X"79",X"03",X"18",X"C9",X"1D",X"B0",X"02",X"A9",X"1D",X"99",X"03",X"18",X"CA",X"08",X"4C",X"4A",
		X"D3",X"85",X"F5",X"EA",X"A4",X"09",X"B5",X"A9",X"30",X"0D",X"B9",X"03",X"18",X"85",X"0B",X"EA",
		X"0B",X"4C",X"31",X"D3",X"85",X"F5",X"6E",X"B9",X"03",X"18",X"85",X"0B",X"E2",X"0B",X"C1",X"F5",
		X"EA",X"A5",X"0B",X"99",X"03",X"18",X"C1",X"F5",X"EA",X"B5",X"A9",X"29",X"F0",X"F0",X"0B",X"F6",
		X"A9",X"B5",X"A9",X"29",X"F3",X"95",X"A9",X"C1",X"F5",X"EA",X"60",X"5B",X"D3",X"6F",X"D3",X"83",
		X"D3",X"97",X"D3",X"AE",X"D3",X"B1",X"D3",X"B4",X"D3",X"B7",X"D3",X"47",X"48",X"47",X"48",X"40",
		X"41",X"42",X"41",X"40",X"41",X"42",X"41",X"45",X"FF",X"46",X"FF",X"43",X"FF",X"44",X"FF",X"00",
		X"00",X"00",X"00",X"58",X"59",X"58",X"59",X"58",X"59",X"58",X"59",X"5C",X"FF",X"5D",X"FF",X"5A",
		X"FF",X"5B",X"FF",X"00",X"00",X"00",X"00",X"64",X"65",X"64",X"65",X"64",X"65",X"64",X"65",X"68",
		X"FF",X"69",X"FF",X"66",X"FF",X"67",X"FF",X"00",X"00",X"00",X"00",X"70",X"71",X"70",X"71",X"70",
		X"71",X"70",X"71",X"74",X"FF",X"75",X"FF",X"72",X"FF",X"73",X"FF",X"85",X"F5",X"6E",X"85",X"F5",
		X"EA",X"85",X"F5",X"EA",X"85",X"F5",X"6E",X"00",X"00",X"FE",X"00",X"02",X"00",X"00",X"FD",X"00",
		X"03",X"85",X"F5",X"EA",X"B5",X"A9",X"4A",X"4A",X"4A",X"4A",X"A8",X"B9",X"E8",X"D3",X"85",X"05",
		X"B9",X"E9",X"D3",X"85",X"06",X"46",X"0A",X"0A",X"A8",X"B9",X"02",X"18",X"85",X"03",X"5D",X"03",
		X"18",X"85",X"04",X"E6",X"67",X"AC",X"05",X"00",X"F5",X"D3",X"FD",X"D3",X"2E",X"D4",X"5F",X"D4",
		X"AD",X"D4",X"85",X"F5",X"6E",X"A9",X"00",X"85",X"67",X"60",X"85",X"F5",X"6E",X"A5",X"03",X"C9",
		X"16",X"B0",X"0A",X"A9",X"17",X"99",X"02",X"18",X"D0",X"20",X"85",X"F5",X"EA",X"20",X"00",X"D5",
		X"D0",X"18",X"20",X"88",X"D5",X"D0",X"13",X"A5",X"04",X"38",X"E9",X"01",X"29",X"F0",X"09",X"0D",
		X"99",X"03",X"18",X"A9",X"00",X"85",X"67",X"85",X"F5",X"EA",X"60",X"85",X"F5",X"EA",X"A5",X"03",
		X"C9",X"D8",X"90",X"0A",X"A9",X"D8",X"99",X"02",X"18",X"D0",X"20",X"85",X"F5",X"EA",X"20",X"00",
		X"D5",X"D0",X"18",X"20",X"AB",X"D5",X"D0",X"13",X"A5",X"04",X"38",X"E9",X"01",X"29",X"F0",X"09",
		X"0D",X"99",X"03",X"18",X"A9",X"00",X"85",X"67",X"85",X"F5",X"EA",X"60",X"85",X"F5",X"EA",X"A5",
		X"04",X"C9",X"1D",X"B0",X"0A",X"A9",X"1D",X"99",X"03",X"18",X"D0",X"34",X"85",X"F5",X"EA",X"20",
		X"23",X"D5",X"D0",X"2C",X"20",X"1E",X"D6",X"D0",X"27",X"8A",X"48",X"A5",X"08",X"29",X"F8",X"48",
		X"AD",X"03",X"40",X"29",X"40",X"F0",X"1D",X"68",X"A6",X"1F",X"85",X"F5",X"EA",X"18",X"7D",X"FA",
		X"D4",X"99",X"02",X"18",X"68",X"AA",X"85",X"F5",X"EA",X"A9",X"00",X"85",X"67",X"85",X"F5",X"EA",
		X"60",X"85",X"F5",X"EA",X"68",X"A2",X"00",X"4C",X"8D",X"D4",X"85",X"F5",X"EA",X"A5",X"04",X"C9",
		X"DD",X"90",X"0A",X"A9",X"DD",X"99",X"03",X"18",X"D0",X"36",X"85",X"F5",X"EA",X"A5",X"03",X"20",
		X"23",X"D5",X"D0",X"2C",X"20",X"41",X"D6",X"D0",X"27",X"8A",X"48",X"A5",X"08",X"29",X"F8",X"48",
		X"AD",X"03",X"40",X"29",X"40",X"F0",X"1D",X"68",X"A6",X"1F",X"85",X"F5",X"EA",X"18",X"7D",X"FA",
		X"D4",X"99",X"02",X"18",X"68",X"AA",X"85",X"F5",X"EA",X"A9",X"00",X"85",X"67",X"85",X"F5",X"EA",
		X"60",X"85",X"F5",X"EA",X"68",X"A2",X"00",X"4C",X"DD",X"D4",X"FF",X"01",X"FE",X"02",X"85",X"F5",
		X"EA",X"A5",X"04",X"29",X"0F",X"F0",X"19",X"C9",X"0F",X"F0",X"15",X"C9",X"0E",X"F0",X"11",X"C9",
		X"0D",X"F0",X"0D",X"C9",X"0C",X"F0",X"09",X"C9",X"0B",X"F0",X"05",X"C9",X"0A",X"85",X"F5",X"6E",
		X"60",X"85",X"F5",X"EA",X"A5",X"03",X"85",X"08",X"AD",X"03",X"40",X"29",X"40",X"F0",X"0B",X"A5",
		X"1F",X"F0",X"07",X"C6",X"08",X"E2",X"08",X"C1",X"F5",X"EA",X"E6",X"08",X"EA",X"08",X"EA",X"08",
		X"A5",X"08",X"29",X"0F",X"C9",X"06",X"90",X"28",X"C9",X"08",X"90",X"39",X"C9",X"0E",X"B0",X"33",
		X"85",X"F5",X"EA",X"A5",X"08",X"29",X"F0",X"C9",X"10",X"F0",X"2A",X"C9",X"40",X"F0",X"26",X"C9",
		X"70",X"F0",X"22",X"C9",X"A0",X"F0",X"1E",X"C9",X"D0",X"F0",X"1A",X"D0",X"18",X"85",X"F5",X"6E",
		X"A5",X"08",X"29",X"F0",X"C9",X"30",X"F0",X"0D",X"C9",X"60",X"F0",X"09",X"C9",X"90",X"F0",X"05",
		X"C9",X"C0",X"85",X"F5",X"6E",X"60",X"85",X"F5",X"EA",X"A5",X"03",X"38",X"E9",X"08",X"4A",X"4A",
		X"4A",X"4A",X"85",X"12",X"4D",X"0F",X"38",X"E5",X"12",X"85",X"12",X"A5",X"04",X"18",X"69",X"07",
		X"29",X"F0",X"18",X"65",X"12",X"AA",X"4C",X"CC",X"D5",X"85",X"F5",X"EA",X"A5",X"03",X"18",X"69",
		X"19",X"4A",X"4A",X"4A",X"4A",X"85",X"12",X"4D",X"0F",X"38",X"E5",X"12",X"85",X"12",X"C9",X"04",
		X"18",X"69",X"07",X"29",X"F0",X"18",X"65",X"12",X"AA",X"85",X"F5",X"EA",X"BD",X"8E",X"D6",X"AA",
		X"BD",X"00",X"04",X"4A",X"4A",X"4A",X"4A",X"C9",X"00",X"F0",X"3E",X"C9",X"05",X"F0",X"3A",X"C9",
		X"06",X"F0",X"36",X"C9",X"07",X"F0",X"32",X"A5",X"03",X"18",X"69",X"05",X"4A",X"4A",X"4A",X"4A",
		X"85",X"12",X"A9",X"0F",X"38",X"E5",X"12",X"85",X"12",X"A5",X"04",X"18",X"69",X"10",X"29",X"F0",
		X"18",X"65",X"12",X"AA",X"BD",X"8E",X"D6",X"AA",X"BD",X"00",X"04",X"4A",X"4A",X"4A",X"4A",X"C9",
		X"07",X"F0",X"06",X"A9",X"00",X"60",X"85",X"F5",X"EA",X"A9",X"FF",X"60",X"85",X"F5",X"EA",X"A5",
		X"03",X"18",X"69",X"07",X"4A",X"4A",X"4A",X"4A",X"85",X"12",X"A9",X"0F",X"38",X"E5",X"12",X"85",
		X"12",X"A5",X"04",X"18",X"69",X"11",X"29",X"F0",X"18",X"65",X"12",X"AA",X"4C",X"62",X"D6",X"85",
		X"F5",X"EA",X"A5",X"03",X"18",X"69",X"07",X"4A",X"4A",X"4A",X"4A",X"85",X"12",X"A9",X"0F",X"38",
		X"E5",X"12",X"85",X"12",X"A5",X"04",X"18",X"69",X"14",X"29",X"F0",X"18",X"65",X"12",X"AA",X"85",
		X"F5",X"EA",X"BD",X"8E",X"D6",X"AA",X"BD",X"00",X"04",X"4A",X"4A",X"4A",X"4A",X"C9",X"00",X"F0",
		X"1A",X"C9",X"01",X"F0",X"16",X"C9",X"02",X"F0",X"12",X"C9",X"09",X"F0",X"0E",X"C9",X"0A",X"F0",
		X"0A",X"C9",X"0B",X"F0",X"06",X"A9",X"00",X"60",X"85",X"F5",X"EA",X"A9",X"FF",X"60",X"00",X"01",
		X"02",X"03",X"04",X"05",X"06",X"07",X"87",X"86",X"85",X"84",X"83",X"82",X"81",X"80",X"08",X"09",
		X"0A",X"0B",X"0C",X"0D",X"0E",X"0F",X"8F",X"8E",X"8D",X"8C",X"8B",X"8A",X"89",X"88",X"10",X"11",
		X"12",X"13",X"14",X"15",X"16",X"17",X"97",X"96",X"95",X"94",X"93",X"92",X"91",X"90",X"18",X"19",
		X"1A",X"1B",X"1C",X"1D",X"1E",X"1F",X"9F",X"9E",X"9D",X"9C",X"9B",X"9A",X"99",X"98",X"20",X"21",
		X"22",X"23",X"24",X"25",X"26",X"27",X"A7",X"A6",X"A5",X"A4",X"A3",X"A2",X"A1",X"A0",X"28",X"29",
		X"2A",X"2B",X"2C",X"2D",X"2E",X"2F",X"AF",X"AE",X"AD",X"AC",X"AB",X"AA",X"A9",X"A8",X"30",X"31",
		X"32",X"33",X"34",X"35",X"36",X"37",X"B7",X"B6",X"B5",X"B4",X"B3",X"B2",X"B1",X"B0",X"38",X"39",
		X"3A",X"3B",X"3C",X"3D",X"3E",X"3F",X"BF",X"BE",X"BD",X"BC",X"BB",X"BA",X"B9",X"B8",X"40",X"41",
		X"42",X"43",X"44",X"45",X"46",X"47",X"C7",X"C6",X"C5",X"C4",X"C3",X"C2",X"C1",X"C0",X"48",X"49",
		X"4A",X"4B",X"4C",X"4D",X"4E",X"4F",X"CF",X"CE",X"CD",X"CC",X"CB",X"CA",X"C9",X"C8",X"50",X"51",
		X"52",X"53",X"54",X"55",X"56",X"57",X"D7",X"D6",X"D5",X"D4",X"D3",X"D2",X"D1",X"D0",X"58",X"59",
		X"5A",X"5B",X"5C",X"5D",X"5E",X"5F",X"DF",X"DE",X"DD",X"DC",X"DB",X"DA",X"D9",X"D8",X"60",X"61",
		X"62",X"63",X"64",X"65",X"66",X"67",X"E7",X"E6",X"E5",X"E4",X"E3",X"E2",X"E1",X"E0",X"68",X"69",
		X"6A",X"6B",X"6C",X"6D",X"6E",X"6F",X"EF",X"EE",X"ED",X"EC",X"EB",X"EA",X"E9",X"E8",X"70",X"71",
		X"72",X"73",X"74",X"75",X"76",X"77",X"F7",X"F6",X"F5",X"F4",X"F3",X"F2",X"F1",X"F0",X"78",X"79",
		X"7A",X"7B",X"7C",X"7D",X"7E",X"7F",X"FF",X"FE",X"FD",X"FC",X"FB",X"FA",X"F9",X"F8",X"85",X"F6",
		X"EA",X"4C",X"38",X"D8",X"85",X"F5",X"6E",X"A5",X"6E",X"C9",X"FF",X"D0",X"03",X"4C",X"63",X"D8",
		X"20",X"72",X"E6",X"E6",X"6E",X"C9",X"6E",X"C9",X"01",X"F0",X"1A",X"C9",X"09",X"F0",X"4B",X"C9",
		X"11",X"F0",X"66",X"C9",X"19",X"F0",X"DA",X"C9",X"22",X"F0",X"04",X"60",X"85",X"F6",X"6E",X"4C",
		X"57",X"D8",X"85",X"F5",X"6E",X"A5",X"BA",X"4A",X"A8",X"B9",X"64",X"D8",X"8D",X"1C",X"18",X"5D",
		X"6E",X"D8",X"8D",X"1D",X"18",X"5D",X"69",X"D8",X"8D",X"18",X"18",X"B9",X"82",X"D8",X"8D",X"19",
		X"18",X"A6",X"1F",X"B5",X"2B",X"38",X"F8",X"E9",X"01",X"95",X"2B",X"D8",X"A5",X"1B",X"F0",X"06",
		X"20",X"94",X"CA",X"85",X"F6",X"6E",X"60",X"85",X"F5",X"EA",X"A5",X"BA",X"4A",X"A8",X"AD",X"1D",
		X"18",X"D9",X"6E",X"D8",X"D0",X"09",X"B9",X"73",X"D8",X"8D",X"1D",X"18",X"85",X"F6",X"EA",X"B9",
		X"87",X"D8",X"8D",X"19",X"18",X"60",X"85",X"F5",X"EA",X"A5",X"BA",X"4A",X"A8",X"AD",X"1D",X"18",
		X"D9",X"73",X"D8",X"D0",X"09",X"B9",X"78",X"D8",X"8D",X"1D",X"18",X"85",X"F6",X"EA",X"B9",X"8C",
		X"D8",X"8D",X"19",X"18",X"60",X"85",X"F5",X"EA",X"A5",X"BA",X"4A",X"A8",X"AD",X"1D",X"18",X"D9",
		X"78",X"D8",X"D0",X"09",X"B9",X"7D",X"D8",X"8D",X"1D",X"18",X"85",X"F6",X"EA",X"B9",X"91",X"D8",
		X"8D",X"19",X"18",X"60",X"85",X"F5",X"EA",X"A9",X"FF",X"85",X"6E",X"A9",X"00",X"8D",X"18",X"18",
		X"85",X"F5",X"EA",X"60",X"03",X"03",X"01",X"01",X"01",X"03",X"03",X"01",X"01",X"05",X"49",X"49",
		X"49",X"4B",X"4A",X"41",X"41",X"41",X"48",X"47",X"49",X"49",X"49",X"4B",X"4A",X"41",X"41",X"41",
		X"48",X"47",X"20",X"20",X"20",X"24",X"24",X"21",X"21",X"21",X"25",X"25",X"22",X"22",X"22",X"26",
		X"26",X"23",X"23",X"23",X"27",X"27",X"85",X"F5",X"EA",X"A5",X"BA",X"C9",X"06",X"F0",X"50",X"C9",
		X"08",X"F0",X"4C",X"AD",X"1E",X"18",X"49",X"FF",X"38",X"E9",X"28",X"4A",X"4A",X"4A",X"85",X"03",
		X"A9",X"00",X"85",X"04",X"AD",X"1F",X"18",X"29",X"F8",X"18",X"69",X"10",X"0A",X"26",X"04",X"0A",
		X"26",X"04",X"18",X"65",X"03",X"85",X"05",X"85",X"03",X"A5",X"04",X"69",X"10",X"85",X"04",X"18",
		X"69",X"04",X"85",X"06",X"A0",X"24",X"B1",X"05",X"29",X"03",X"F0",X"13",X"A0",X"04",X"B1",X"05",
		X"29",X"03",X"F0",X"0B",X"B1",X"03",X"29",X"1F",X"C9",X"04",X"90",X"06",X"85",X"F5",X"EA",X"4C",
		X"55",X"DA",X"85",X"F5",X"EA",X"A9",X"08",X"20",X"5D",X"EA",X"20",X"6A",X"DA",X"A5",X"BA",X"C9",
		X"02",X"F0",X"15",X"C8",X"85",X"F5",X"6E",X"20",X"58",X"DA",X"F0",X"1F",X"C8",X"C0",X"08",X"D0",
		X"F6",X"A0",X"04",X"D0",X"5F",X"85",X"F5",X"6E",X"88",X"85",X"F5",X"EA",X"20",X"58",X"DA",X"F0",
		X"2E",X"88",X"D0",X"F8",X"A0",X"01",X"D0",X"4C",X"85",X"F5",X"EA",X"8A",X"D0",X"0D",X"85",X"F5",
		X"EA",X"C8",X"B1",X"05",X"29",X"03",X"D0",X"F9",X"85",X"F5",X"EA",X"A2",X"04",X"85",X"F5",X"6E",
		X"88",X"B1",X"03",X"29",X"1C",X"F0",X"A8",X"CA",X"D0",X"F6",X"F0",X"28",X"85",X"F5",X"6E",X"8A",
		X"D0",X"0D",X"85",X"F5",X"6E",X"88",X"B1",X"05",X"29",X"03",X"D0",X"F9",X"85",X"F5",X"6E",X"A2",
		X"04",X"85",X"F5",X"EA",X"C8",X"B1",X"03",X"29",X"1C",X"F0",X"84",X"CA",X"D0",X"F6",X"88",X"88",
		X"88",X"85",X"F5",X"EA",X"A9",X"09",X"20",X"5D",X"EA",X"98",X"18",X"65",X"03",X"85",X"07",X"C9",
		X"04",X"69",X"00",X"29",X"03",X"85",X"08",X"C9",X"07",X"29",X"1F",X"0A",X"0A",X"0A",X"85",X"09",
		X"46",X"08",X"66",X"07",X"A2",X"08",X"AA",X"07",X"A5",X"07",X"29",X"F8",X"85",X"07",X"4A",X"00",
		X"85",X"F5",X"EA",X"BD",X"02",X"02",X"F0",X"1E",X"BD",X"03",X"02",X"49",X"FF",X"29",X"F8",X"C5",
		X"09",X"D0",X"0C",X"BD",X"04",X"02",X"29",X"F8",X"C5",X"07",X"F0",X"10",X"85",X"F5",X"6E",X"E8",
		X"E8",X"E8",X"E8",X"4C",X"A3",X"D9",X"4C",X"31",X"DA",X"85",X"F5",X"EA",X"BD",X"02",X"02",X"C9",
		X"0F",X"B0",X"EC",X"29",X"0F",X"09",X"10",X"9D",X"02",X"02",X"BD",X"04",X"02",X"29",X"FC",X"09",
		X"04",X"9D",X"04",X"02",X"4D",X"01",X"9D",X"05",X"02",X"A0",X"00",X"84",X"0A",X"C1",X"F5",X"6E",
		X"A4",X"0A",X"B9",X"68",X"00",X"29",X"A0",X"D0",X"2D",X"98",X"0A",X"0A",X"A8",X"B9",X"02",X"18",
		X"18",X"69",X"08",X"DD",X"03",X"02",X"B0",X"1E",X"18",X"69",X"20",X"DD",X"03",X"02",X"90",X"16",
		X"B9",X"03",X"18",X"29",X"F8",X"18",X"69",X"10",X"85",X"0B",X"BD",X"04",X"02",X"29",X"F8",X"C5",
		X"0B",X"F0",X"13",X"85",X"F5",X"EA",X"E6",X"0A",X"A4",X"0A",X"C0",X"06",X"D0",X"C2",X"85",X"F5",
		X"EA",X"F0",X"22",X"85",X"F5",X"EA",X"A4",X"0A",X"B9",X"68",X"00",X"29",X"0F",X"09",X"40",X"99",
		X"68",X"00",X"96",X"B1",X"FE",X"05",X"02",X"FE",X"05",X"02",X"A9",X"12",X"20",X"5D",X"EA",X"4C",
		X"26",X"DA",X"85",X"F5",X"EA",X"60",X"85",X"F5",X"EA",X"A2",X"FF",X"B1",X"05",X"29",X"03",X"F0",
		X"25",X"E8",X"B1",X"03",X"29",X"1C",X"F0",X"1E",X"85",X"F5",X"EA",X"84",X"12",X"18",X"B1",X"03",
		X"69",X"04",X"91",X"03",X"18",X"98",X"69",X"20",X"A8",X"B1",X"03",X"69",X"04",X"91",X"03",X"A4",
		X"12",X"A9",X"FF",X"85",X"F5",X"EA",X"60",X"85",X"F5",X"EA",X"A0",X"00",X"AD",X"04",X"40",X"29",
		X"08",X"D0",X"05",X"A0",X"06",X"85",X"F5",X"EA",X"18",X"98",X"65",X"64",X"AA",X"BD",X"02",X"DB",
		X"85",X"BC",X"BD",X"0E",X"DB",X"85",X"BD",X"BD",X"1A",X"DB",X"85",X"BE",X"A9",X"00",X"85",X"C2",
		X"85",X"C3",X"85",X"BF",X"85",X"C0",X"85",X"C1",X"85",X"90",X"A6",X"1F",X"B5",X"61",X"4A",X"4A",
		X"85",X"03",X"C9",X"08",X"90",X"02",X"A9",X"07",X"AA",X"BD",X"F0",X"DA",X"A0",X"05",X"85",X"F5",
		X"EA",X"99",X"91",X"00",X"88",X"10",X"FA",X"BD",X"F9",X"DA",X"A0",X"05",X"85",X"F5",X"EA",X"99",
		X"A1",X"00",X"88",X"10",X"FA",X"AD",X"F4",X"DA",X"85",X"98",X"AD",X"FD",X"DA",X"85",X"A8",X"60",
		X"0F",X"03",X"07",X"0F",X"03",X"07",X"0F",X"03",X"07",X"04",X"03",X"03",X"03",X"02",X"02",X"02",
		X"01",X"01",X"03",X"03",X"02",X"04",X"00",X"02",X"05",X"05",X"02",X"04",X"00",X"02",X"00",X"00",
		X"03",X"02",X"02",X"02",X"00",X"00",X"03",X"02",X"02",X"02",X"01",X"01",X"01",X"00",X"04",X"02",
		X"01",X"01",X"01",X"00",X"04",X"02",X"85",X"F5",X"EA",X"A5",X"6F",X"30",X"6E",X"A5",X"13",X"29",
		X"1F",X"D0",X"68",X"E6",X"C2",X"CA",X"C2",X"E0",X"03",X"D0",X"02",X"A2",X"00",X"86",X"C2",X"D9",
		X"BC",X"D5",X"BF",X"F0",X"56",X"A0",X"00",X"85",X"F5",X"EA",X"B9",X"68",X"00",X"C9",X"FF",X"F0",
		X"0B",X"C8",X"C0",X"06",X"D0",X"F4",X"4C",X"9B",X"DB",X"85",X"F5",X"EA",X"F6",X"BF",X"6C",X"8A",
		X"09",X"20",X"99",X"68",X"00",X"C0",X"0A",X"4D",X"01",X"99",X"99",X"00",X"EA",X"C3",X"C9",X"C3",
		X"29",X"03",X"85",X"C3",X"0D",X"01",X"AA",X"BD",X"9C",X"DB",X"99",X"A9",X"00",X"54",X"0A",X"0A",
		X"A8",X"BD",X"9E",X"DB",X"99",X"02",X"18",X"C9",X"63",X"0A",X"0A",X"18",X"65",X"C3",X"AA",X"BD",
		X"A1",X"DB",X"99",X"03",X"18",X"08",X"EB",X"DC",X"85",X"F5",X"EA",X"60",X"20",X"40",X"F0",X"00",
		X"1D",X"1D",X"AD",X"AD",X"1D",X"1D",X"5D",X"5D",X"1D",X"1D",X"8D",X"AD",X"1D",X"1D",X"8D",X"8D",
		X"1D",X"1D",X"CD",X"CD",X"1D",X"2D",X"9D",X"8D",X"80",X"85",X"F5",X"EA",X"A5",X"6F",X"30",X"1C",
		X"A2",X"00",X"85",X"F5",X"6E",X"B5",X"68",X"29",X"D0",X"D0",X"09",X"B5",X"68",X"29",X"20",X"D0",
		X"0F",X"85",X"F5",X"EA",X"E8",X"E0",X"06",X"D0",X"EC",X"85",X"F5",X"EA",X"60",X"85",X"F5",X"6E",
		X"86",X"70",X"B5",X"A9",X"85",X"71",X"46",X"0A",X"0A",X"A8",X"B9",X"02",X"18",X"85",X"03",X"5D",
		X"03",X"18",X"85",X"04",X"C9",X"03",X"C9",X"D9",X"B0",X"54",X"C9",X"18",X"90",X"60",X"20",X"B6",
		X"E0",X"D0",X"42",X"C9",X"10",X"F0",X"13",X"C9",X"40",X"F0",X"0F",X"C9",X"70",X"F0",X"0B",X"C9",
		X"A0",X"F0",X"07",X"C9",X"D0",X"D0",X"2E",X"85",X"F5",X"EA",X"20",X"9D",X"E0",X"D0",X"0D",X"20",
		X"7B",X"E0",X"F0",X"13",X"20",X"8C",X"E0",X"F0",X"0E",X"85",X"F5",X"EA",X"20",X"59",X"E0",X"F0",
		X"06",X"4C",X"6B",X"DC",X"85",X"F5",X"EA",X"A6",X"70",X"B5",X"68",X"29",X"0F",X"95",X"68",X"4C",
		X"6B",X"DC",X"85",X"F5",X"EA",X"A5",X"03",X"C9",X"80",X"B0",X"13",X"85",X"F5",X"EA",X"A6",X"70",
		X"B5",X"A9",X"29",X"0F",X"09",X"20",X"95",X"A9",X"4C",X"6B",X"DC",X"85",X"F5",X"EA",X"A6",X"70",
		X"B5",X"A9",X"29",X"0F",X"09",X"40",X"95",X"A9",X"85",X"F5",X"EA",X"A6",X"70",X"20",X"69",X"D2",
		X"A6",X"70",X"4C",X"D4",X"DB",X"85",X"F5",X"EA",X"A5",X"13",X"29",X"3F",X"D0",X"6A",X"E6",X"90",
		X"A5",X"90",X"C9",X"14",X"90",X"2E",X"A9",X"00",X"85",X"90",X"A2",X"05",X"85",X"F5",X"EA",X"B5",
		X"91",X"29",X"10",X"F0",X"11",X"B5",X"A1",X"C9",X"02",X"F0",X"13",X"D6",X"A1",X"A9",X"03",X"95",
		X"91",X"D0",X"0B",X"85",X"F5",X"EA",X"38",X"B5",X"91",X"36",X"91",X"85",X"F5",X"EA",X"CA",X"10",
		X"DE",X"85",X"F5",X"EA",X"A0",X"05",X"A2",X"14",X"85",X"F5",X"EA",X"B9",X"68",X"00",X"30",X"09",
		X"B5",X"73",X"F0",X"11",X"D6",X"73",X"85",X"F5",X"EA",X"88",X"CA",X"CA",X"CA",X"CA",X"10",X"EB",
		X"30",X"16",X"85",X"F5",X"EA",X"8A",X"48",X"98",X"48",X"84",X"0A",X"20",X"EB",X"DC",X"68",X"A8",
		X"68",X"AA",X"4C",X"C9",X"DC",X"85",X"F5",X"EA",X"60",X"85",X"F5",X"EA",X"A4",X"0A",X"B9",X"68",
		X"00",X"29",X"03",X"0A",X"A8",X"B9",X"2A",X"DD",X"85",X"03",X"B9",X"2B",X"DD",X"85",X"04",X"B9",
		X"30",X"DD",X"85",X"05",X"5D",X"31",X"DD",X"85",X"06",X"A5",X"0A",X"0A",X"0A",X"AA",X"B4",X"75",
		X"B1",X"03",X"95",X"72",X"59",X"05",X"95",X"73",X"A9",X"00",X"95",X"74",X"FA",X"75",X"D8",X"75",
		X"B1",X"03",X"10",X"07",X"A9",X"00",X"95",X"75",X"85",X"F5",X"EA",X"60",X"38",X"DD",X"4D",X"DD",
		X"5A",X"DD",X"43",X"DD",X"54",X"DD",X"5F",X"DD",X"04",X"03",X"04",X"05",X"04",X"04",X"05",X"04",
		X"04",X"04",X"FF",X"03",X"03",X"07",X"05",X"03",X"03",X"05",X"03",X"03",X"03",X"03",X"03",X"04",
		X"03",X"03",X"04",X"FF",X"03",X"03",X"07",X"09",X"0D",X"03",X"05",X"05",X"04",X"05",X"FF",X"09",
		X"17",X"09",X"13",X"85",X"F5",X"6E",X"A5",X"6F",X"30",X"19",X"A2",X"05",X"86",X"70",X"C1",X"F5",
		X"EA",X"A6",X"70",X"B5",X"68",X"29",X"F0",X"F0",X"0E",X"85",X"F5",X"EA",X"C6",X"70",X"10",X"F1",
		X"85",X"F5",X"EA",X"60",X"85",X"F5",X"6E",X"8A",X"0A",X"0A",X"A8",X"B9",X"02",X"18",X"85",X"03",
		X"B9",X"03",X"18",X"85",X"04",X"D9",X"8A",X"F0",X"0B",X"D6",X"8A",X"85",X"F5",X"6E",X"4C",X"BB",
		X"DE",X"85",X"F5",X"EA",X"20",X"9D",X"E0",X"D0",X"F5",X"20",X"B6",X"E0",X"D0",X"F0",X"AD",X"1E",
		X"18",X"85",X"17",X"AD",X"1F",X"18",X"85",X"18",X"A5",X"70",X"0A",X"0A",X"AA",X"B4",X"72",X"F0",
		X"11",X"88",X"F0",X"14",X"88",X"F0",X"17",X"88",X"F0",X"1A",X"88",X"F0",X"20",X"D0",X"44",X"85",
		X"F5",X"EA",X"4C",X"ED",X"DD",X"85",X"F5",X"6E",X"4C",X"13",X"DE",X"85",X"F5",X"6E",X"4C",X"ED",
		X"DD",X"85",X"F5",X"EA",X"A5",X"17",X"69",X"08",X"85",X"17",X"85",X"F5",X"6E",X"A6",X"70",X"B5",
		X"A9",X"85",X"71",X"29",X"F0",X"C9",X"20",X"85",X"F5",X"EA",X"F0",X"23",X"C9",X"40",X"85",X"F5",
		X"EA",X"F0",X"31",X"C9",X"60",X"85",X"F5",X"EA",X"F0",X"3F",X"85",X"F5",X"EA",X"4C",X"5E",X"DE",
		X"85",X"F5",X"EA",X"A5",X"18",X"69",X"08",X"85",X"18",X"4C",X"ED",X"DD",X"85",X"F5",X"EA",X"A5",
		X"18",X"29",X"F8",X"85",X"05",X"A5",X"04",X"29",X"F8",X"C5",X"05",X"B0",X"46",X"F0",X"4A",X"90",
		X"4E",X"85",X"F5",X"EA",X"A5",X"18",X"29",X"F8",X"85",X"05",X"A5",X"04",X"29",X"F8",X"C5",X"05",
		X"B0",X"43",X"F0",X"47",X"90",X"4B",X"85",X"F5",X"EA",X"A5",X"17",X"29",X"F8",X"85",X"05",X"A5",
		X"03",X"29",X"F8",X"C5",X"05",X"90",X"4C",X"F0",X"44",X"B0",X"3C",X"85",X"F5",X"EA",X"A5",X"17",
		X"29",X"F8",X"85",X"05",X"A5",X"03",X"29",X"F8",X"C5",X"05",X"90",X"49",X"F0",X"41",X"B0",X"39",
		X"85",X"F5",X"EA",X"4C",X"E7",X"DE",X"85",X"F5",X"EA",X"4C",X"01",X"DF",X"85",X"F5",X"EA",X"4C",
		X"1B",X"DF",X"85",X"F5",X"EA",X"4C",X"35",X"DF",X"85",X"F5",X"EA",X"4C",X"55",X"DF",X"85",X"F5",
		X"EA",X"4C",X"6F",X"DF",X"85",X"F5",X"EA",X"4C",X"89",X"DF",X"85",X"F5",X"EA",X"4C",X"A3",X"DF",
		X"85",X"F5",X"EA",X"4C",X"BD",X"DF",X"85",X"F5",X"EA",X"4C",X"D7",X"DF",X"85",X"F5",X"EA",X"4C",
		X"F1",X"DF",X"85",X"F5",X"EA",X"4C",X"0B",X"E0",X"85",X"F5",X"EA",X"A6",X"70",X"20",X"C3",X"D3",
		X"D0",X"0B",X"A6",X"70",X"20",X"69",X"D2",X"4C",X"7C",X"DD",X"85",X"F5",X"EA",X"A6",X"70",X"B5",
		X"A9",X"85",X"71",X"29",X"F0",X"C9",X"20",X"F0",X"28",X"C9",X"40",X"F0",X"AE",X"C9",X"60",X"F0",
		X"BC",X"4C",X"F1",X"DF",X"85",X"F5",X"EA",X"20",X"59",X"E0",X"F0",X"63",X"20",X"7B",X"E0",X"F0",
		X"5E",X"20",X"8C",X"E0",X"F0",X"59",X"20",X"6A",X"E0",X"F0",X"54",X"4C",X"3D",X"E0",X"85",X"F5",
		X"EA",X"20",X"7B",X"E0",X"F0",X"49",X"20",X"59",X"E0",X"F0",X"44",X"20",X"6A",X"E0",X"F0",X"3F",
		X"20",X"8C",X"E0",X"F0",X"3A",X"4C",X"3D",X"E0",X"85",X"F5",X"EA",X"20",X"6A",X"E0",X"F0",X"2F",
		X"20",X"7B",X"E0",X"F0",X"2A",X"20",X"8C",X"E0",X"F0",X"25",X"20",X"59",X"E0",X"F0",X"20",X"4C",
		X"3D",X"E0",X"85",X"F5",X"6E",X"20",X"59",X"E0",X"F0",X"15",X"20",X"8C",X"E0",X"F0",X"10",X"20",
		X"6A",X"E0",X"F0",X"0B",X"20",X"7B",X"E0",X"F0",X"06",X"4C",X"3D",X"E0",X"85",X"F5",X"6E",X"4C",
		X"25",X"E0",X"85",X"F5",X"6E",X"20",X"8C",X"E0",X"F0",X"F5",X"20",X"6A",X"E0",X"F0",X"F0",X"20",
		X"59",X"E0",X"F0",X"EB",X"20",X"7B",X"E0",X"F0",X"E6",X"4C",X"3D",X"E0",X"85",X"F5",X"6E",X"20",
		X"6A",X"E0",X"F0",X"DB",X"20",X"8C",X"E0",X"F0",X"D6",X"20",X"59",X"E0",X"F0",X"D1",X"20",X"7B",
		X"E0",X"F0",X"CC",X"4C",X"3D",X"E0",X"85",X"F5",X"EA",X"20",X"7B",X"E0",X"F0",X"C1",X"20",X"59",
		X"E0",X"F0",X"BC",X"20",X"8C",X"E0",X"F0",X"B7",X"20",X"6A",X"E0",X"F0",X"B2",X"4C",X"3D",X"E0",
		X"85",X"F5",X"EA",X"20",X"59",X"E0",X"F0",X"7D",X"20",X"7B",X"E0",X"F0",X"78",X"20",X"8C",X"E0",
		X"F0",X"73",X"20",X"6A",X"E0",X"F0",X"6E",X"4C",X"3D",X"E0",X"85",X"F5",X"6E",X"20",X"8C",X"E0",
		X"F0",X"63",X"20",X"59",X"E0",X"F0",X"5E",X"20",X"7B",X"E0",X"F0",X"59",X"20",X"6A",X"E0",X"F0",
		X"54",X"4C",X"3D",X"E0",X"85",X"F5",X"6E",X"20",X"7B",X"E0",X"F0",X"49",X"20",X"6A",X"E0",X"F0",
		X"44",X"20",X"8C",X"E0",X"F0",X"3F",X"20",X"59",X"E0",X"F0",X"3A",X"4C",X"3D",X"E0",X"85",X"F5",
		X"EA",X"20",X"6A",X"E0",X"F0",X"2F",X"20",X"8C",X"E0",X"F0",X"2A",X"20",X"7B",X"E0",X"F0",X"25",
		X"20",X"59",X"E0",X"F0",X"20",X"4C",X"3D",X"E0",X"85",X"F5",X"EA",X"20",X"8C",X"E0",X"F0",X"15",
		X"20",X"6A",X"E0",X"F0",X"10",X"20",X"7B",X"E0",X"F0",X"0B",X"20",X"59",X"E0",X"F0",X"06",X"4C",
		X"3D",X"E0",X"85",X"F5",X"EA",X"A6",X"70",X"A9",X"00",X"95",X"74",X"A9",X"10",X"95",X"8A",X"85",
		X"F5",X"EA",X"A6",X"70",X"20",X"69",X"D2",X"4C",X"7B",X"DD",X"85",X"F5",X"EA",X"A6",X"70",X"B5",
		X"68",X"29",X"03",X"AA",X"D6",X"BE",X"A6",X"70",X"0A",X"0A",X"A8",X"A9",X"00",X"99",X"00",X"18",
		X"A9",X"FF",X"95",X"68",X"4C",X"7C",X"DD",X"85",X"F5",X"EA",X"A6",X"70",X"A5",X"71",X"29",X"0F",
		X"09",X"60",X"95",X"A9",X"20",X"C3",X"D3",X"60",X"85",X"F5",X"EA",X"A6",X"70",X"A5",X"71",X"29",
		X"0F",X"09",X"80",X"95",X"A9",X"20",X"C3",X"D3",X"60",X"85",X"F5",X"EA",X"A6",X"70",X"A5",X"71",
		X"29",X"0F",X"09",X"20",X"95",X"A9",X"20",X"C3",X"D3",X"60",X"85",X"F5",X"EA",X"A6",X"70",X"A5",
		X"71",X"29",X"0F",X"09",X"40",X"95",X"A9",X"20",X"C3",X"D3",X"60",X"85",X"F5",X"EA",X"A5",X"04",
		X"29",X"0F",X"C9",X"0F",X"F0",X"0D",X"C9",X"0E",X"F0",X"09",X"C9",X"0D",X"F0",X"05",X"C9",X"0C",
		X"85",X"F5",X"EA",X"60",X"85",X"F5",X"EA",X"A5",X"03",X"85",X"08",X"E6",X"08",X"E6",X"08",X"A5",
		X"08",X"29",X"0C",X"F0",X"1E",X"C9",X"08",X"D0",X"2F",X"A5",X"08",X"29",X"F0",X"C9",X"10",X"F0",
		X"27",X"C9",X"40",X"F0",X"23",X"C9",X"70",X"F0",X"1F",X"C9",X"A0",X"F0",X"1B",X"C9",X"D0",X"60",
		X"85",X"F5",X"EA",X"A5",X"08",X"29",X"F0",X"C9",X"30",X"F0",X"0D",X"C9",X"60",X"F0",X"09",X"C9",
		X"90",X"F0",X"05",X"C9",X"C0",X"85",X"F5",X"EA",X"60",X"85",X"F5",X"EA",X"86",X"11",X"84",X"12",
		X"A4",X"64",X"B9",X"88",X"E1",X"85",X"C4",X"C8",X"63",X"98",X"0A",X"AA",X"BD",X"76",X"E1",X"85",
		X"03",X"BD",X"77",X"E1",X"85",X"04",X"5D",X"82",X"E1",X"AA",X"A0",X"00",X"91",X"03",X"6C",X"8A",
		X"C8",X"91",X"03",X"A0",X"20",X"E8",X"8A",X"91",X"03",X"E8",X"8A",X"C8",X"91",X"03",X"4D",X"00",
		X"85",X"60",X"A4",X"12",X"A6",X"11",X"A9",X"0B",X"20",X"5D",X"EA",X"85",X"F5",X"6E",X"60",X"85",
		X"F5",X"EA",X"A5",X"C4",X"F0",X"2F",X"20",X"F2",X"E8",X"A5",X"13",X"29",X"3F",X"D0",X"26",X"C6",
		X"C4",X"D0",X"22",X"A5",X"63",X"0A",X"AA",X"BD",X"76",X"E1",X"85",X"03",X"DD",X"77",X"E1",X"85",
		X"04",X"A9",X"00",X"A8",X"91",X"03",X"64",X"91",X"03",X"A0",X"20",X"91",X"03",X"64",X"91",X"03",
		X"85",X"60",X"85",X"F5",X"6E",X"60",X"4F",X"11",X"CF",X"11",X"CF",X"11",X"8F",X"10",X"15",X"11",
		X"8F",X"11",X"BC",X"C0",X"B8",X"BC",X"C0",X"B8",X"07",X"06",X"05",X"05",X"05",X"05",X"85",X"F5",
		X"EA",X"A9",X"00",X"8D",X"00",X"02",X"C1",X"F5",X"EA",X"AC",X"00",X"02",X"B9",X"02",X"02",X"D0",
		X"04",X"60",X"85",X"F5",X"6E",X"29",X"0F",X"85",X"03",X"B9",X"03",X"02",X"85",X"04",X"5D",X"04",
		X"02",X"85",X"05",X"B9",X"02",X"02",X"29",X"F0",X"4A",X"4A",X"4A",X"AA",X"BD",X"C9",X"E1",X"85",
		X"06",X"BD",X"CA",X"E1",X"85",X"07",X"AC",X"06",X"00",X"00",X"E2",X"18",X"E2",X"36",X"E2",X"78",
		X"E2",X"B0",X"E2",X"E8",X"E2",X"00",X"E4",X"EC",X"E1",X"EF",X"E1",X"F2",X"E1",X"20",X"E3",X"58",
		X"E3",X"90",X"E3",X"C8",X"E3",X"57",X"E4",X"03",X"E2",X"85",X"F5",X"EA",X"85",X"F5",X"6E",X"85",
		X"F5",X"EA",X"00",X"B9",X"02",X"02",X"29",X"0F",X"09",X"10",X"99",X"02",X"02",X"C1",X"F5",X"6E",
		X"85",X"F5",X"EA",X"20",X"BE",X"E5",X"EE",X"00",X"02",X"EE",X"00",X"02",X"EE",X"00",X"02",X"EE",
		X"00",X"02",X"4C",X"99",X"E1",X"85",X"F5",X"EA",X"20",X"16",X"E5",X"D0",X"13",X"20",X"6E",X"E5",
		X"D0",X"0E",X"20",X"A2",X"CC",X"98",X"AA",X"FE",X"04",X"02",X"20",X"6B",X"EB",X"85",X"F5",X"EA",
		X"4C",X"03",X"E2",X"85",X"F5",X"EA",X"B9",X"05",X"02",X"29",X"10",X"D0",X"1E",X"38",X"A5",X"05",
		X"E9",X"08",X"85",X"05",X"99",X"04",X"02",X"20",X"A9",X"E4",X"B9",X"05",X"02",X"09",X"10",X"99",
		X"05",X"02",X"85",X"F5",X"EA",X"4C",X"03",X"E2",X"85",X"F5",X"EA",X"A5",X"13",X"29",X"03",X"D0",
		X"F4",X"B9",X"05",X"02",X"29",X"0F",X"99",X"05",X"02",X"B9",X"02",X"02",X"29",X"0F",X"09",X"30",
		X"99",X"02",X"02",X"D0",X"E0",X"85",X"F5",X"EA",X"B9",X"05",X"02",X"29",X"10",X"D0",X"14",X"20",
		X"B2",X"E4",X"B9",X"05",X"02",X"09",X"10",X"99",X"05",X"02",X"85",X"F5",X"EA",X"4C",X"03",X"E2",
		X"85",X"F5",X"EA",X"A5",X"13",X"29",X"03",X"D0",X"F4",X"B9",X"05",X"02",X"29",X"0F",X"99",X"05",
		X"02",X"B9",X"02",X"02",X"29",X"0F",X"09",X"40",X"99",X"02",X"02",X"D0",X"E0",X"85",X"F5",X"EA",
		X"B9",X"05",X"02",X"29",X"10",X"D0",X"14",X"20",X"BB",X"E4",X"B9",X"05",X"02",X"09",X"10",X"99",
		X"05",X"02",X"85",X"F5",X"EA",X"4C",X"03",X"E2",X"85",X"F5",X"EA",X"A5",X"13",X"29",X"03",X"D0",
		X"F4",X"B9",X"05",X"02",X"29",X"0F",X"99",X"05",X"02",X"B9",X"02",X"02",X"09",X"50",X"29",X"5F",
		X"99",X"02",X"02",X"D0",X"E0",X"85",X"F5",X"EA",X"B9",X"05",X"02",X"29",X"10",X"D0",X"14",X"20",
		X"C4",X"E4",X"B9",X"05",X"02",X"09",X"10",X"99",X"05",X"02",X"85",X"F5",X"EA",X"4C",X"03",X"E2",
		X"85",X"F5",X"EA",X"A5",X"13",X"29",X"03",X"D0",X"F4",X"B9",X"05",X"02",X"29",X"0F",X"99",X"05",
		X"02",X"B9",X"02",X"02",X"09",X"60",X"29",X"6F",X"99",X"02",X"02",X"D0",X"E0",X"85",X"F5",X"6E",
		X"B9",X"05",X"02",X"29",X"10",X"D0",X"14",X"20",X"A9",X"E4",X"B9",X"05",X"02",X"09",X"10",X"99",
		X"05",X"02",X"85",X"F5",X"6E",X"4C",X"03",X"E2",X"85",X"F5",X"EA",X"A5",X"13",X"29",X"03",X"D0",
		X"F4",X"B9",X"05",X"02",X"29",X"0F",X"99",X"05",X"02",X"B9",X"02",X"02",X"29",X"0F",X"09",X"B0",
		X"99",X"02",X"02",X"D0",X"E0",X"85",X"F5",X"6E",X"B9",X"05",X"02",X"29",X"10",X"D0",X"14",X"20",
		X"B2",X"E4",X"B9",X"05",X"02",X"09",X"10",X"99",X"05",X"02",X"85",X"F5",X"6E",X"4C",X"03",X"E2",
		X"85",X"F5",X"EA",X"A5",X"13",X"29",X"03",X"D0",X"F4",X"B9",X"05",X"02",X"29",X"0F",X"99",X"05",
		X"02",X"B9",X"02",X"02",X"09",X"C0",X"29",X"CF",X"99",X"02",X"02",X"D0",X"E0",X"85",X"F5",X"6E",
		X"B9",X"05",X"02",X"29",X"10",X"D0",X"14",X"20",X"BB",X"E4",X"B9",X"05",X"02",X"09",X"10",X"99",
		X"05",X"02",X"85",X"F5",X"6E",X"4C",X"03",X"E2",X"85",X"F5",X"EA",X"A5",X"13",X"29",X"03",X"D0",
		X"F4",X"B9",X"05",X"02",X"29",X"0F",X"99",X"05",X"02",X"B9",X"02",X"02",X"09",X"D0",X"29",X"DF",
		X"99",X"02",X"02",X"D0",X"E0",X"85",X"F5",X"6E",X"B9",X"05",X"02",X"29",X"10",X"D0",X"14",X"20",
		X"C4",X"E4",X"B9",X"05",X"02",X"09",X"10",X"99",X"05",X"02",X"85",X"F5",X"6E",X"4C",X"03",X"E2",
		X"85",X"F5",X"EA",X"A5",X"13",X"29",X"03",X"D0",X"F4",X"B9",X"05",X"02",X"29",X"0F",X"99",X"05",
		X"02",X"B9",X"02",X"02",X"09",X"E0",X"29",X"EF",X"99",X"02",X"02",X"D0",X"E0",X"85",X"F5",X"6E",
		X"20",X"A2",X"CC",X"98",X"AA",X"FE",X"04",X"02",X"BD",X"04",X"02",X"29",X"07",X"D0",X"42",X"B9",
		X"02",X"02",X"29",X"0F",X"09",X"10",X"99",X"02",X"02",X"B9",X"05",X"02",X"29",X"0F",X"99",X"05",
		X"02",X"B9",X"06",X"02",X"29",X"0F",X"C9",X"0F",X"F0",X"0C",X"B9",X"06",X"02",X"29",X"F0",X"C9",
		X"F0",X"D0",X"1E",X"85",X"F5",X"EA",X"A9",X"00",X"99",X"05",X"02",X"B9",X"02",X"02",X"09",X"F0",
		X"99",X"02",X"02",X"A9",X"00",X"20",X"8C",X"E9",X"20",X"FA",X"E5",X"20",X"C8",X"E7",X"85",X"F5",
		X"EA",X"4C",X"03",X"E2",X"85",X"F5",X"EA",X"20",X"A2",X"CC",X"98",X"AA",X"BD",X"05",X"02",X"29",
		X"0F",X"9D",X"05",X"02",X"F0",X"08",X"DE",X"05",X"02",X"D0",X"19",X"85",X"F5",X"EA",X"B9",X"02",
		X"02",X"29",X"0F",X"99",X"02",X"02",X"A9",X"00",X"20",X"8C",X"E9",X"20",X"FA",X"E5",X"4C",X"03",
		X"E2",X"85",X"F5",X"EA",X"B9",X"02",X"02",X"29",X"0F",X"09",X"10",X"99",X"02",X"02",X"B9",X"04",
		X"02",X"69",X"02",X"99",X"04",X"02",X"4C",X"03",X"E2",X"00",X"01",X"01",X"05",X"02",X"04",X"03",
		X"00",X"01",X"01",X"05",X"02",X"04",X"03",X"85",X"F5",X"EA",X"A9",X"00",X"85",X"11",X"F0",X"1C",
		X"85",X"F5",X"EA",X"A9",X"01",X"85",X"11",X"F0",X"13",X"85",X"F5",X"EA",X"A9",X"02",X"85",X"11",
		X"F0",X"0A",X"85",X"F5",X"EA",X"A9",X"03",X"85",X"11",X"85",X"F5",X"EA",X"98",X"48",X"A6",X"11",
		X"A5",X"05",X"18",X"7D",X"0C",X"E5",X"85",X"05",X"20",X"99",X"CC",X"A0",X"01",X"A6",X"11",X"A5",
		X"06",X"29",X"FB",X"85",X"06",X"B1",X"05",X"18",X"7D",X"10",X"E5",X"91",X"05",X"C8",X"B1",X"05",
		X"18",X"7D",X"10",X"E5",X"91",X"05",X"A0",X"21",X"B1",X"05",X"18",X"7D",X"10",X"E5",X"91",X"05",
		X"C8",X"B1",X"05",X"18",X"7D",X"10",X"E5",X"91",X"05",X"68",X"A8",X"60",X"04",X"03",X"02",X"01",
		X"04",X"FC",X"04",X"FC",X"85",X"F5",X"6E",X"A5",X"05",X"29",X"07",X"D0",X"4C",X"B9",X"07",X"02",
		X"C5",X"04",X"D0",X"45",X"B9",X"08",X"02",X"38",X"E5",X"05",X"C9",X"09",X"B0",X"3B",X"B9",X"02",
		X"02",X"29",X"0F",X"09",X"20",X"99",X"02",X"02",X"B9",X"06",X"02",X"29",X"F0",X"C9",X"F0",X"F0",
		X"1D",X"B9",X"06",X"02",X"29",X"0F",X"C9",X"0F",X"F0",X"14",X"B9",X"06",X"02",X"09",X"10",X"99",
		X"06",X"02",X"B9",X"08",X"02",X"18",X"69",X"04",X"99",X"08",X"02",X"85",X"F5",X"6E",X"A9",X"0A",
		X"20",X"5D",X"EA",X"A9",X"FF",X"60",X"85",X"F5",X"EA",X"A9",X"00",X"60",X"85",X"F5",X"6E",X"A5",
		X"05",X"29",X"0F",X"C9",X"08",X"D0",X"2D",X"A5",X"04",X"4A",X"4A",X"4A",X"4A",X"85",X"12",X"4D",
		X"10",X"38",X"E5",X"12",X"85",X"12",X"C9",X"05",X"29",X"F0",X"18",X"65",X"12",X"AA",X"BD",X"8E",
		X"D6",X"AA",X"BD",X"00",X"04",X"4A",X"4A",X"4A",X"4A",X"C9",X"09",X"F0",X"0D",X"C9",X"08",X"F0",
		X"09",X"85",X"F5",X"EA",X"A9",X"00",X"60",X"85",X"F5",X"EA",X"B9",X"02",X"02",X"29",X"0F",X"09",
		X"A0",X"99",X"02",X"02",X"4D",X"0A",X"20",X"5D",X"EA",X"A9",X"FF",X"60",X"85",X"F5",X"6E",X"A2",
		X"00",X"85",X"F5",X"EA",X"B5",X"68",X"29",X"E0",X"C9",X"40",X"F0",X"0C",X"85",X"F5",X"6E",X"E8",
		X"E0",X"06",X"D0",X"F0",X"60",X"85",X"F5",X"6E",X"B5",X"B1",X"85",X"0D",X"E0",X"0D",X"D0",X"EF",
		X"84",X"0E",X"38",X"B9",X"04",X"02",X"E9",X"0C",X"85",X"0F",X"8A",X"0A",X"0A",X"A8",X"A5",X"0F",
		X"99",X"03",X"18",X"A4",X"0E",X"4C",X"CF",X"E5",X"85",X"F5",X"EA",X"A2",X"00",X"86",X"C9",X"C1",
		X"F5",X"EA",X"B5",X"68",X"30",X"07",X"29",X"40",X"D0",X"2F",X"85",X"F5",X"EA",X"E8",X"E0",X"06",
		X"D0",X"F0",X"A6",X"C9",X"F0",X"1F",X"BD",X"63",X"E6",X"20",X"8C",X"E9",X"98",X"48",X"A6",X"CA",
		X"BC",X"4F",X"EB",X"A6",X"C9",X"BD",X"69",X"E6",X"99",X"01",X"18",X"A9",X"01",X"99",X"00",X"18",
		X"68",X"A8",X"85",X"F5",X"EA",X"60",X"85",X"F5",X"EA",X"B5",X"B1",X"85",X"0D",X"C4",X"0D",X"D0",
		X"CC",X"E6",X"C9",X"86",X"CA",X"B5",X"68",X"29",X"0F",X"09",X"20",X"95",X"68",X"84",X"0E",X"29",
		X"03",X"A8",X"B9",X"4C",X"E7",X"BC",X"4F",X"EB",X"99",X"01",X"18",X"A4",X"0E",X"A9",X"7F",X"95",
		X"99",X"4C",X"0D",X"E6",X"04",X"05",X"07",X"08",X"09",X"0A",X"37",X"38",X"39",X"3A",X"3B",X"3C",
		X"85",X"F5",X"EA",X"AD",X"1A",X"18",X"85",X"03",X"AD",X"1B",X"18",X"85",X"04",X"A2",X"00",X"85",
		X"F5",X"EA",X"B5",X"68",X"10",X"0C",X"85",X"F5",X"EA",X"E8",X"E0",X"06",X"D0",X"F4",X"60",X"85",
		X"F5",X"EA",X"8A",X"0A",X"0A",X"A8",X"B9",X"02",X"18",X"18",X"69",X"0C",X"C5",X"03",X"90",X"E9",
		X"E9",X"18",X"C5",X"03",X"B0",X"E3",X"B9",X"03",X"18",X"18",X"69",X"0C",X"C5",X"04",X"90",X"D9",
		X"E9",X"18",X"C5",X"04",X"B0",X"D3",X"B5",X"68",X"09",X"10",X"95",X"68",X"A4",X"1F",X"B9",X"61",
		X"00",X"C9",X"08",X"90",X"02",X"A9",X"08",X"A8",X"B9",X"D4",X"E6",X"95",X"99",X"A9",X"0F",X"20",
		X"5D",X"EA",X"4C",X"89",X"E6",X"D1",X"C1",X"B1",X"A1",X"91",X"81",X"71",X"61",X"85",X"F5",X"EA",
		X"A2",X"00",X"85",X"F5",X"EA",X"B5",X"68",X"30",X"07",X"29",X"10",X"D0",X"0C",X"85",X"F5",X"EA",
		X"E8",X"E0",X"06",X"D0",X"F0",X"60",X"85",X"F5",X"EA",X"B5",X"99",X"C9",X"01",X"F0",X"39",X"D6",
		X"99",X"B5",X"99",X"29",X"0F",X"D0",X"E9",X"B5",X"99",X"29",X"10",X"F0",X"0F",X"B5",X"68",X"29",
		X"03",X"A8",X"B9",X"4C",X"E7",X"85",X"03",X"70",X"10",X"85",X"F5",X"EA",X"B5",X"68",X"29",X"03",
		X"A8",X"B9",X"53",X"E7",X"85",X"03",X"C1",X"F5",X"EA",X"8A",X"0A",X"0A",X"A8",X"A5",X"03",X"99",
		X"01",X"18",X"4C",X"F0",X"E6",X"85",X"F5",X"6E",X"B5",X"68",X"29",X"EF",X"95",X"68",X"0D",X"03",
		X"A8",X"B9",X"5A",X"E7",X"85",X"03",X"A4",X"29",X"E7",X"85",X"F5",X"EA",X"00",X"62",X"6E",X"7A",
		X"85",X"F5",X"EA",X"00",X"63",X"6F",X"7B",X"85",X"F5",X"EA",X"00",X"5A",X"66",X"72",X"85",X"F5",
		X"EA",X"A5",X"6F",X"30",X"1E",X"AD",X"1E",X"18",X"85",X"03",X"AD",X"1F",X"18",X"85",X"04",X"4A",
		X"00",X"85",X"F5",X"EA",X"B5",X"68",X"10",X"0F",X"85",X"F5",X"EA",X"E8",X"E0",X"06",X"D0",X"F4",
		X"85",X"F5",X"EA",X"60",X"85",X"F5",X"6E",X"29",X"70",X"D0",X"F0",X"8A",X"0A",X"0A",X"A8",X"B9",
		X"02",X"18",X"18",X"69",X"08",X"C5",X"03",X"90",X"E2",X"E9",X"10",X"C5",X"03",X"B0",X"DC",X"B9",
		X"03",X"18",X"18",X"69",X"04",X"C5",X"04",X"90",X"D2",X"E9",X"0D",X"C5",X"04",X"B0",X"CC",X"A9",
		X"10",X"20",X"5D",X"EA",X"A5",X"6F",X"09",X"F0",X"85",X"6F",X"A9",X"FF",X"85",X"A0",X"4D",X"00",
		X"20",X"5D",X"EA",X"4C",X"7B",X"E7",X"85",X"F5",X"EA",X"A6",X"1F",X"F6",X"65",X"C8",X"63",X"B5",
		X"65",X"85",X"05",X"D9",X"15",X"E8",X"D0",X"03",X"20",X"FB",X"E0",X"A5",X"05",X"D9",X"1B",X"E8",
		X"D0",X"03",X"20",X"FB",X"E0",X"A5",X"05",X"D9",X"21",X"E8",X"D0",X"03",X"20",X"FB",X"E0",X"A5",
		X"05",X"D9",X"27",X"E8",X"D0",X"03",X"20",X"FB",X"E0",X"A5",X"05",X"D9",X"2D",X"E8",X"90",X"14",
		X"A5",X"6F",X"29",X"0F",X"09",X"80",X"85",X"6F",X"A9",X"FF",X"85",X"A0",X"A9",X"05",X"20",X"5D",
		X"EA",X"85",X"F5",X"EA",X"60",X"04",X"05",X"04",X"06",X"03",X"03",X"08",X"07",X"08",X"10",X"06",
		X"07",X"0C",X"0D",X"0E",X"16",X"09",X"0C",X"FF",X"FF",X"0E",X"1C",X"FF",X"0E",X"10",X"10",X"12",
		X"20",X"10",X"12",X"85",X"F5",X"EA",X"A5",X"6F",X"29",X"F0",X"C9",X"80",X"D0",X"2B",X"A5",X"A0",
		X"F0",X"22",X"C6",X"A0",X"A5",X"A0",X"29",X"0F",X"D0",X"1F",X"A5",X"A0",X"29",X"10",X"F0",X"07",
		X"A9",X"47",X"D0",X"08",X"85",X"F5",X"EA",X"A9",X"4C",X"85",X"F5",X"EA",X"8D",X"1D",X"18",X"D0",
		X"08",X"85",X"F5",X"EA",X"E6",X"C5",X"85",X"F5",X"EA",X"60",X"85",X"F5",X"EA",X"A5",X"C6",X"30",
		X"46",X"A5",X"6F",X"29",X"F0",X"C9",X"F0",X"F0",X"04",X"60",X"85",X"F5",X"EA",X"A2",X"1B",X"A5",
		X"A0",X"85",X"F5",X"EA",X"DD",X"B8",X"E8",X"F0",X"09",X"CA",X"10",X"F8",X"C6",X"A0",X"60",X"85",
		X"F5",X"EA",X"BD",X"D4",X"E8",X"8D",X"1D",X"18",X"C6",X"A0",X"8A",X"D0",X"0E",X"A6",X"1F",X"D6",
		X"29",X"A9",X"FF",X"85",X"C6",X"4C",X"B7",X"E8",X"85",X"F5",X"EA",X"E0",X"18",X"D0",X"08",X"A9",
		X"10",X"20",X"5D",X"EA",X"85",X"F5",X"EA",X"60",X"01",X"08",X"10",X"18",X"20",X"28",X"30",X"38",
		X"40",X"48",X"50",X"58",X"60",X"68",X"78",X"80",X"88",X"90",X"98",X"A0",X"A8",X"B0",X"B8",X"C0",
		X"C8",X"D0",X"F8",X"FE",X"52",X"51",X"52",X"51",X"52",X"51",X"52",X"51",X"52",X"51",X"52",X"51",
		X"52",X"51",X"52",X"51",X"52",X"51",X"52",X"51",X"52",X"51",X"52",X"51",X"50",X"4F",X"4E",X"4D",
		X"85",X"F5",X"EA",X"A5",X"60",X"D0",X"7A",X"A6",X"63",X"BD",X"72",X"E9",X"85",X"03",X"BD",X"78",
		X"E9",X"85",X"04",X"AD",X"1E",X"18",X"18",X"69",X"08",X"C5",X"03",X"90",X"64",X"E9",X"10",X"C5",
		X"03",X"B0",X"5E",X"AD",X"1F",X"18",X"18",X"69",X"08",X"C5",X"04",X"90",X"54",X"E9",X"10",X"C5",
		X"04",X"B0",X"4E",X"8A",X"0A",X"A8",X"B9",X"76",X"E1",X"85",X"03",X"B9",X"77",X"E1",X"85",X"04",
		X"BC",X"81",X"E9",X"B9",X"7E",X"E9",X"85",X"05",X"A0",X"00",X"91",X"03",X"64",X"E6",X"05",X"C9",
		X"05",X"91",X"03",X"A9",X"00",X"A0",X"20",X"91",X"03",X"C8",X"91",X"03",X"4D",X"02",X"85",X"C4",
		X"E6",X"60",X"BC",X"81",X"E9",X"B9",X"87",X"E9",X"20",X"8C",X"E9",X"A6",X"1F",X"B5",X"2B",X"18",
		X"F8",X"69",X"01",X"95",X"2B",X"74",X"20",X"94",X"CA",X"A9",X"11",X"20",X"5D",X"EA",X"85",X"F5",
		X"EA",X"60",X"78",X"78",X"78",X"78",X"48",X"78",X"50",X"70",X"70",X"20",X"40",X"60",X"AC",X"B0",
		X"B4",X"00",X"01",X"02",X"00",X"01",X"02",X"04",X"05",X"06",X"85",X"F5",X"6E",X"85",X"04",X"46",
		X"48",X"98",X"48",X"A5",X"1B",X"D0",X"06",X"4C",X"33",X"EA",X"85",X"F5",X"6E",X"A6",X"1F",X"BC",
		X"59",X"EA",X"A6",X"04",X"18",X"F8",X"B9",X"2D",X"00",X"7D",X"38",X"EA",X"99",X"2D",X"00",X"5D",
		X"2E",X"00",X"7D",X"43",X"EA",X"99",X"2E",X"00",X"B9",X"2F",X"00",X"7D",X"4E",X"EA",X"99",X"2F",
		X"00",X"D8",X"A6",X"1F",X"20",X"4E",X"C9",X"A6",X"1F",X"BC",X"59",X"EA",X"A5",X"35",X"D9",X"2F",
		X"00",X"90",X"15",X"D0",X"2A",X"A5",X"34",X"D9",X"2E",X"00",X"90",X"0C",X"D0",X"21",X"A5",X"33",
		X"D9",X"2D",X"00",X"B0",X"1A",X"85",X"F5",X"6E",X"B9",X"2D",X"00",X"85",X"33",X"5D",X"2E",X"00",
		X"85",X"34",X"B9",X"2F",X"00",X"85",X"35",X"4A",X"02",X"20",X"4E",X"C9",X"85",X"F5",X"6E",X"A6",
		X"1F",X"BC",X"59",X"EA",X"8A",X"0A",X"AA",X"B9",X"2F",X"00",X"D5",X"5D",X"90",X"25",X"B9",X"2E",
		X"00",X"D5",X"5C",X"90",X"1E",X"18",X"F8",X"B5",X"5C",X"65",X"5A",X"95",X"5C",X"B5",X"5D",X"65",
		X"5B",X"95",X"5D",X"D8",X"A6",X"1F",X"F6",X"29",X"20",X"54",X"CA",X"A9",X"02",X"20",X"5D",X"EA",
		X"85",X"F5",X"EA",X"68",X"A8",X"68",X"AA",X"60",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"02",X"03",X"05",X"10",X"15",X"20",X"40",X"80",X"60",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"03",X"85",X"F5",X"EA",X"86",X"C7",
		X"A6",X"1B",X"F0",X"0A",X"AA",X"BD",X"71",X"EA",X"8D",X"03",X"40",X"85",X"F5",X"EA",X"A6",X"C7",
		X"60",X"00",X"1B",X"1C",X"04",X"01",X"02",X"20",X"21",X"11",X"12",X"13",X"14",X"15",X"16",X"17",
		X"18",X"19",X"1A",X"1D",X"13",X"14",X"15",X"16",X"17",X"05",X"03",X"85",X"F5",X"EA",X"A2",X"05",
		X"85",X"F5",X"EA",X"B5",X"68",X"29",X"F0",X"C9",X"80",X"F0",X"0D",X"85",X"F5",X"EA",X"CA",X"10",
		X"F2",X"85",X"F5",X"EA",X"60",X"85",X"F5",X"EA",X"B5",X"99",X"C9",X"01",X"F0",X"48",X"D6",X"99",
		X"B5",X"99",X"C9",X"40",X"F0",X"43",X"C9",X"38",X"F0",X"53",X"C9",X"30",X"F0",X"63",X"C9",X"28",
		X"F0",X"23",X"C9",X"20",X"D0",X"D8",X"B5",X"68",X"29",X"03",X"A8",X"B9",X"65",X"EB",X"20",X"8C",
		X"E9",X"B9",X"62",X"EB",X"BC",X"4F",X"EB",X"99",X"01",X"18",X"A9",X"01",X"99",X"00",X"18",X"4C",
		X"9E",X"EA",X"85",X"F5",X"EA",X"B5",X"68",X"29",X"03",X"A8",X"B9",X"5F",X"EB",X"BC",X"4F",X"EB",
		X"99",X"01",X"18",X"4C",X"9E",X"EA",X"4C",X"35",X"EB",X"B5",X"68",X"29",X"03",X"A8",X"B9",X"56",
		X"EB",X"BC",X"4F",X"EB",X"99",X"01",X"18",X"A4",X"9E",X"EA",X"85",X"F5",X"6E",X"B5",X"68",X"29",
		X"03",X"A8",X"B9",X"59",X"EB",X"BC",X"4F",X"EB",X"99",X"01",X"18",X"4C",X"9E",X"EA",X"85",X"F5",
		X"EA",X"B5",X"68",X"29",X"03",X"A8",X"B9",X"5C",X"EB",X"BC",X"4F",X"EB",X"99",X"01",X"18",X"A4",
		X"9E",X"EA",X"85",X"F5",X"6E",X"86",X"03",X"D9",X"68",X"29",X"03",X"AA",X"D6",X"BE",X"CA",X"03",
		X"A9",X"FF",X"95",X"68",X"DC",X"4F",X"EB",X"A9",X"00",X"99",X"00",X"18",X"A4",X"9E",X"EA",X"00",
		X"04",X"08",X"0C",X"10",X"14",X"18",X"1C",X"5E",X"6A",X"76",X"5F",X"6B",X"77",X"60",X"6C",X"78",
		X"61",X"6D",X"79",X"34",X"35",X"36",X"01",X"02",X"03",X"85",X"F5",X"EA",X"A2",X"05",X"85",X"F5",
		X"EA",X"B5",X"68",X"10",X"0A",X"85",X"F5",X"6E",X"CA",X"10",X"F6",X"60",X"85",X"F5",X"6E",X"BC",
		X"4F",X"EB",X"B9",X"02",X"18",X"85",X"03",X"5D",X"03",X"18",X"85",X"04",X"CC",X"00",X"02",X"B9",
		X"03",X"02",X"E9",X"08",X"C5",X"03",X"90",X"E0",X"E9",X"20",X"C5",X"03",X"B0",X"DA",X"B9",X"04",
		X"02",X"E9",X"05",X"C5",X"04",X"B0",X"D1",X"69",X"0C",X"C5",X"04",X"90",X"CB",X"B5",X"68",X"29",
		X"0F",X"09",X"80",X"95",X"68",X"4D",X"42",X"95",X"99",X"A9",X"0C",X"20",X"5E",X"EA",X"4C",X"78",
		X"EB",X"85",X"F6",X"EA",X"A9",X"05",X"85",X"2B",X"85",X"2C",X"AD",X"04",X"40",X"29",X"10",X"D0",
		X"05",X"C6",X"2B",X"85",X"F6",X"6E",X"60",X"01",X"D7",X"48",X"06",X"D7",X"68",X"04",X"D7",X"98",
		X"02",X"D7",X"B8",X"0F",X"D7",X"E8",X"01",X"A7",X"28",X"06",X"A7",X"78",X"04",X"A7",X"98",X"02",
		X"A7",X"B8",X"0F",X"A7",X"E8",X"01",X"77",X"28",X"06",X"77",X"48",X"04",X"77",X"78",X"02",X"77",
		X"B8",X"0F",X"77",X"E8",X"01",X"47",X"28",X"06",X"47",X"48",X"04",X"47",X"68",X"02",X"47",X"88",
		X"0F",X"47",X"E8",X"FF",X"01",X"A7",X"28",X"05",X"A7",X"38",X"06",X"A7",X"48",X"04",X"A7",X"58",
		X"06",X"A7",X"68",X"04",X"A7",X"78",X"05",X"A7",X"88",X"02",X"A7",X"98",X"0F",X"A7",X"E8",X"01",
		X"77",X"28",X"05",X"77",X"38",X"04",X"77",X"48",X"06",X"77",X"58",X"04",X"77",X"68",X"05",X"77",
		X"78",X"06",X"77",X"88",X"02",X"77",X"98",X"0F",X"77",X"E8",X"FF",X"01",X"D7",X"28",X"06",X"D7",
		X"38",X"03",X"D7",X"48",X"02",X"D7",X"68",X"0F",X"D7",X"B8",X"01",X"A7",X"28",X"03",X"A7",X"38",
		X"06",X"A7",X"58",X"02",X"A7",X"A8",X"0F",X"A7",X"E8",X"01",X"77",X"28",X"03",X"77",X"78",X"06",
		X"77",X"98",X"02",X"77",X"A8",X"0F",X"77",X"E8",X"01",X"47",X"28",X"06",X"47",X"48",X"03",X"47",
		X"58",X"02",X"47",X"68",X"0F",X"47",X"B8",X"FF",X"01",X"D7",X"28",X"04",X"D7",X"48",X"02",X"D7",
		X"58",X"0F",X"D7",X"88",X"01",X"D7",X"98",X"05",X"D7",X"A8",X"02",X"D7",X"B8",X"0F",X"D7",X"E8",
		X"01",X"A7",X"28",X"05",X"A7",X"38",X"02",X"A7",X"58",X"0F",X"A7",X"B8",X"01",X"77",X"28",X"04",
		X"77",X"38",X"02",X"77",X"58",X"0F",X"77",X"B8",X"01",X"47",X"28",X"05",X"47",X"48",X"02",X"47",
		X"58",X"0F",X"47",X"88",X"01",X"47",X"98",X"04",X"47",X"A8",X"02",X"47",X"B8",X"0F",X"47",X"E8",
		X"FF",X"01",X"D7",X"28",X"03",X"D7",X"38",X"05",X"D7",X"48",X"06",X"D7",X"58",X"04",X"D7",X"68",
		X"06",X"D7",X"78",X"05",X"D7",X"88",X"02",X"D7",X"98",X"0F",X"D7",X"E8",X"01",X"A7",X"28",X"06",
		X"A7",X"38",X"05",X"A7",X"48",X"04",X"A7",X"58",X"05",X"A7",X"68",X"03",X"A7",X"78",X"06",X"A7",
		X"88",X"02",X"A7",X"98",X"0F",X"A7",X"E8",X"01",X"77",X"28",X"05",X"77",X"38",X"06",X"77",X"48",
		X"05",X"77",X"58",X"04",X"77",X"68",X"03",X"77",X"78",X"06",X"77",X"88",X"02",X"77",X"98",X"0F",
		X"77",X"E8",X"01",X"47",X"28",X"03",X"47",X"38",X"06",X"47",X"48",X"04",X"47",X"58",X"05",X"47",
		X"68",X"06",X"47",X"78",X"05",X"47",X"88",X"02",X"47",X"98",X"0F",X"47",X"E8",X"FF",X"01",X"D7",
		X"38",X"03",X"D7",X"58",X"04",X"D7",X"78",X"02",X"D7",X"B8",X"0F",X"D7",X"E8",X"01",X"A7",X"28",
		X"03",X"A7",X"48",X"04",X"A7",X"68",X"03",X"A7",X"88",X"02",X"A7",X"A8",X"0F",X"A7",X"E8",X"01",
		X"77",X"38",X"03",X"77",X"58",X"03",X"77",X"78",X"04",X"77",X"98",X"02",X"77",X"B8",X"0F",X"77",
		X"E8",X"01",X"47",X"28",X"04",X"47",X"48",X"03",X"47",X"68",X"02",X"47",X"88",X"0F",X"47",X"E8",
		X"FF",X"01",X"B9",X"AB",X"9A",X"A9",X"BA",X"9B",X"10",X"05",X"60",X"56",X"75",X"50",X"65",X"06",
		X"50",X"03",X"D9",X"C4",X"73",X"C9",X"DC",X"9D",X"30",X"00",X"07",X"3D",X"8C",X"37",X"65",X"06",
		X"50",X"01",X"B8",X"C4",X"05",X"57",X"4C",X"9D",X"30",X"05",X"67",X"3D",X"9C",X"C8",X"D3",X"70",
		X"00",X"05",X"67",X"56",X"05",X"50",X"4C",X"8B",X"10",X"03",X"D8",X"CD",X"9C",X"C9",X"D3",X"76",
		X"50",X"05",X"60",X"56",X"05",X"50",X"65",X"76",X"50",X"03",X"D9",X"CD",X"9C",X"C9",X"DC",X"8D",
		X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"B9",X"AB",X"9A",X"A9",X"BA",X"9B",
		X"10",X"03",X"D9",X"AB",X"9A",X"A9",X"BA",X"8D",X"30",X"01",X"B9",X"AB",X"9C",X"C9",X"D3",X"76",
		X"50",X"03",X"D9",X"AB",X"9A",X"A9",X"B1",X"76",X"50",X"03",X"D9",X"AB",X"9A",X"A9",X"DC",X"8D",
		X"30",X"03",X"D9",X"CD",X"9A",X"A9",X"B1",X"76",X"50",X"03",X"D9",X"AB",X"9A",X"A9",X"D3",X"76",
		X"50",X"03",X"D9",X"AB",X"9A",X"A9",X"D3",X"76",X"50",X"05",X"60",X"00",X"00",X"00",X"2A",X"8D",
		X"30",X"05",X"60",X"00",X"00",X"00",X"65",X"06",X"50",X"05",X"60",X"00",X"00",X"00",X"65",X"06",
		X"50",X"03",X"40",X"00",X"00",X"00",X"4C",X"9D",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"B9",X"AB",X"9A",X"A9",X"BA",X"9B",X"10",X"03",X"D8",X"CD",X"8C",X"37",X"65",X"76",
		X"50",X"03",X"D8",X"C4",X"73",X"C8",X"DC",X"8D",X"30",X"05",X"67",X"3D",X"8C",X"37",X"4C",X"8D",
		X"30",X"03",X"D8",X"CD",X"8C",X"C8",X"DC",X"8D",X"30",X"00",X"00",X"00",X"73",X"C8",X"B1",X"00",
		X"00",X"00",X"00",X"1B",X"8C",X"37",X"00",X"00",X"00",X"00",X"00",X"00",X"73",X"C8",X"B1",X"00",
		X"00",X"00",X"00",X"1B",X"8C",X"C8",X"B1",X"00",X"00",X"00",X"00",X"00",X"05",X"50",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"B9",X"AB",X"9A",X"A9",X"BA",X"9B",
		X"10",X"03",X"D9",X"CD",X"8A",X"A8",X"BA",X"9D",X"30",X"03",X"D9",X"CD",X"9C",X"30",X"4C",X"9D",
		X"30",X"03",X"D9",X"AB",X"8C",X"C9",X"DC",X"9D",X"30",X"00",X"00",X"34",X"73",X"C8",X"B1",X"00",
		X"00",X"00",X"00",X"3D",X"8C",X"C9",X"D3",X"00",X"00",X"00",X"00",X"34",X"00",X"00",X"65",X"00",
		X"00",X"01",X"B9",X"C4",X"00",X"00",X"4C",X"9B",X"10",X"03",X"D8",X"C4",X"00",X"00",X"4C",X"9D",
		X"30",X"03",X"D8",X"C4",X"00",X"00",X"4C",X"8D",X"30",X"00",X"00",X"3D",X"9A",X"A9",X"D3",X"00",
		X"00",X"00",X"00",X"3D",X"8A",X"A8",X"D3",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"B9",X"AB",X"9A",X"A9",X"BA",X"9B",X"10",X"03",X"D9",X"CD",X"9C",X"C9",X"DC",X"9D",
		X"30",X"01",X"B8",X"AB",X"8A",X"A8",X"BA",X"8B",X"10",X"03",X"D9",X"CD",X"9C",X"C9",X"DC",X"9D",
		X"30",X"01",X"B8",X"AB",X"8C",X"C8",X"BA",X"8B",X"10",X"03",X"D9",X"CD",X"9C",X"C9",X"DC",X"9D",
		X"30",X"03",X"D8",X"AB",X"8A",X"A8",X"BA",X"8D",X"30",X"03",X"D9",X"CD",X"9C",X"C9",X"DC",X"9D",
		X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1B",X"9A",X"10",X"2A",X"9B",
		X"10",X"01",X"B9",X"C4",X"71",X"A9",X"D3",X"00",X"00",X"00",X"00",X"3D",X"8A",X"17",X"2A",X"9B",
		X"10",X"01",X"B9",X"C4",X"73",X"C8",X"D3",X"00",X"00",X"00",X"00",X"1B",X"8C",X"30",X"4C",X"9B",
		X"10",X"01",X"B9",X"C4",X"03",X"C9",X"D3",X"00",X"00",X"00",X"00",X"3D",X"9A",X"17",X"2A",X"9B",
		X"10",X"01",X"B9",X"C4",X"73",X"C8",X"D3",X"00",X"00",X"00",X"00",X"1B",X"8A",X"17",X"4C",X"9B",
		X"10",X"01",X"B9",X"C4",X"03",X"C8",X"D3",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"85",X"F5",X"EA",X"A9",X"00",X"85",X"F3",X"85",X"F5",X"EA",X"A9",X"00",X"85",X"ED",X"4D",
		X"36",X"85",X"E4",X"A9",X"00",X"85",X"E5",X"85",X"F5",X"EA",X"A0",X"02",X"85",X"F5",X"EA",X"B1",
		X"E4",X"99",X"E7",X"00",X"88",X"10",X"F8",X"A5",X"E7",X"C9",X"FF",X"D0",X"04",X"60",X"85",X"F5",
		X"EA",X"A5",X"E4",X"18",X"69",X"03",X"85",X"E4",X"A5",X"E5",X"69",X"00",X"85",X"E5",X"E6",X"ED",
		X"F8",X"A5",X"E7",X"38",X"E5",X"CC",X"A5",X"E8",X"E5",X"CD",X"A5",X"E9",X"E5",X"CE",X"D8",X"B0",
		X"C9",X"A6",X"ED",X"BD",X"7E",X"F0",X"18",X"69",X"36",X"85",X"D8",X"A9",X"00",X"85",X"D9",X"A9",
		X"02",X"85",X"DA",X"20",X"8C",X"F0",X"A2",X"02",X"85",X"F5",X"EA",X"A9",X"00",X"95",X"CC",X"CA",
		X"10",X"F9",X"A6",X"ED",X"BD",X"84",X"F0",X"18",X"69",X"36",X"85",X"D8",X"A9",X"00",X"85",X"D9",
		X"A9",X"02",X"85",X"DA",X"20",X"8C",X"F0",X"20",X"D1",X"F0",X"20",X"E3",X"CB",X"60",X"00",X"00",
		X"03",X"06",X"09",X"0C",X"00",X"12",X"15",X"18",X"1B",X"1E",X"85",X"F5",X"EA",X"A4",X"DA",X"85",
		X"F5",X"EA",X"B1",X"D8",X"99",X"EA",X"00",X"88",X"10",X"F8",X"A5",X"EA",X"C9",X"FF",X"D0",X"04",
		X"60",X"85",X"F5",X"EA",X"A4",X"DA",X"85",X"F5",X"EA",X"B9",X"CC",X"00",X"91",X"D8",X"88",X"10",
		X"F8",X"A6",X"DA",X"85",X"F5",X"EA",X"B5",X"EA",X"95",X"CC",X"CA",X"10",X"F9",X"A6",X"DA",X"E8",
		X"8A",X"18",X"65",X"D8",X"85",X"D8",X"A5",X"D9",X"69",X"00",X"85",X"D9",X"4C",X"8D",X"F0",X"85",
		X"F5",X"EA",X"20",X"A3",X"C8",X"20",X"DC",X"F1",X"20",X"F8",X"F2",X"A9",X"05",X"85",X"DC",X"85",
		X"F5",X"EA",X"A5",X"DC",X"18",X"69",X"03",X"85",X"DD",X"0A",X"18",X"65",X"DD",X"AA",X"A5",X"DC",
		X"0A",X"18",X"69",X"10",X"A8",X"20",X"5A",X"C9",X"C6",X"DC",X"10",X"E6",X"A9",X"04",X"85",X"DC",
		X"20",X"B6",X"F1",X"A9",X"00",X"85",X"DE",X"4D",X"07",X"85",X"DF",X"A9",X"06",X"85",X"E0",X"4D",
		X"00",X"85",X"E1",X"85",X"E2",X"C1",X"E3",X"C1",X"F5",X"EA",X"20",X"B8",X"F2",X"20",X"D1",X"F2",
		X"A5",X"E2",X"29",X"0F",X"C9",X"0F",X"D0",X"0C",X"20",X"B8",X"F2",X"A9",X"00",X"8D",X"03",X"40",
		X"60",X"85",X"F5",X"EA",X"A5",X"E2",X"10",X"15",X"A5",X"E3",X"30",X"11",X"A9",X"FF",X"85",X"DE",
		X"A5",X"E3",X"09",X"80",X"85",X"E3",X"4D",X"00",X"85",X"DF",X"85",X"F5",X"6E",X"A5",X"DE",X"05",
		X"DF",X"D0",X"12",X"A5",X"E2",X"10",X"07",X"09",X"0F",X"85",X"E2",X"85",X"F5",X"6E",X"09",X"80",
		X"85",X"E2",X"85",X"F5",X"6E",X"20",X"2F",X"F3",X"20",X"7C",X"F3",X"20",X"E9",X"F3",X"20",X"2F",
		X"F4",X"20",X"9C",X"F5",X"A5",X"E2",X"29",X"20",X"F0",X"1D",X"20",X"DC",X"F1",X"20",X"B6",X"F1",
		X"20",X"F8",X"F2",X"A5",X"E2",X"49",X"20",X"AA",X"A5",X"E3",X"29",X"40",X"D0",X"04",X"E8",X"85",
		X"F5",X"EA",X"86",X"E2",X"C1",X"F5",X"6E",X"20",X"3E",X"F6",X"A5",X"E3",X"29",X"BF",X"85",X"E3",
		X"A5",X"E2",X"29",X"0F",X"C9",X"03",X"90",X"09",X"A5",X"E3",X"09",X"20",X"85",X"E3",X"C1",X"F5",
		X"EA",X"4C",X"1A",X"F1",X"85",X"F5",X"6E",X"A9",X"B4",X"8D",X"02",X"18",X"4D",X"40",X"8D",X"03",
		X"18",X"A9",X"47",X"8D",X"01",X"18",X"4D",X"01",X"8D",X"00",X"18",X"A9",X"00",X"8D",X"04",X"18",
		X"85",X"EE",X"85",X"EF",X"4D",X"17",X"8D",X"05",X"18",X"60",X"85",X"F5",X"6E",X"A9",X"08",X"85",
		X"DD",X"85",X"F5",X"EA",X"A5",X"DD",X"0A",X"AA",X"BD",X"12",X"F2",X"85",X"D8",X"DD",X"24",X"F2",
		X"85",X"DA",X"E8",X"BD",X"12",X"F2",X"85",X"D9",X"BD",X"24",X"F2",X"85",X"DB",X"CA",X"DD",X"BD",
		X"36",X"F2",X"A8",X"85",X"F5",X"EA",X"B1",X"D8",X"91",X"DA",X"88",X"10",X"F9",X"C6",X"DD",X"10",
		X"D3",X"60",X"3F",X"F2",X"52",X"F2",X"65",X"F2",X"78",X"F2",X"83",X"F2",X"92",X"F2",X"9B",X"F2",
		X"A4",X"F2",X"AD",X"F2",X"A8",X"10",X"08",X"11",X"68",X"11",X"C8",X"11",X"4B",X"12",X"D4",X"18",
		X"14",X"1B",X"34",X"1B",X"54",X"1B",X"12",X"12",X"12",X"0A",X"0E",X"08",X"08",X"08",X"08",X"0B",
		X"00",X"0C",X"00",X"0D",X"00",X"0E",X"00",X"0F",X"00",X"10",X"00",X"11",X"00",X"12",X"00",X"13",
		X"00",X"14",X"15",X"00",X"16",X"00",X"17",X"00",X"18",X"00",X"19",X"00",X"1A",X"00",X"1B",X"00",
		X"1C",X"00",X"1D",X"00",X"1E",X"1F",X"00",X"20",X"00",X"21",X"00",X"22",X"00",X"23",X"00",X"24",
		X"00",X"CC",X"00",X"CD",X"00",X"CE",X"00",X"CF",X"1D",X"1A",X"0B",X"00",X"1C",X"1F",X"0C",X"00",
		X"0F",X"18",X"0E",X"3C",X"2F",X"3B",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"41",X"31",X"3D",
		X"40",X"33",X"26",X"00",X"27",X"00",X"28",X"00",X"29",X"00",X"2A",X"3E",X"00",X"3E",X"00",X"3E",
		X"00",X"3E",X"00",X"3E",X"42",X"00",X"42",X"00",X"42",X"00",X"42",X"00",X"42",X"41",X"00",X"41",
		X"00",X"41",X"00",X"41",X"00",X"41",X"85",X"F5",X"EA",X"AD",X"03",X"40",X"10",X"FB",X"85",X"F5",
		X"EA",X"AD",X"03",X"40",X"30",X"FB",X"58",X"EA",X"EA",X"EA",X"78",X"20",X"45",X"D0",X"60",X"85",
		X"F5",X"EA",X"A5",X"DE",X"38",X"E9",X"01",X"85",X"DE",X"A5",X"DF",X"E9",X"00",X"85",X"DF",X"C6",
		X"E0",X"10",X"07",X"A9",X"04",X"85",X"E0",X"85",X"F5",X"EA",X"C6",X"E1",X"10",X"07",X"A9",X"00",
		X"85",X"E1",X"85",X"F5",X"EA",X"60",X"85",X"F5",X"EA",X"A9",X"8B",X"85",X"D8",X"A9",X"12",X"85",
		X"D9",X"A2",X"00",X"85",X"F5",X"6E",X"A0",X"00",X"85",X"F5",X"EA",X"B5",X"48",X"91",X"D8",X"6C",
		X"E0",X"0F",X"D0",X"04",X"60",X"85",X"F5",X"6E",X"C8",X"C0",X"03",X"D0",X"EE",X"A5",X"D8",X"18",
		X"69",X"40",X"85",X"D8",X"C9",X"D9",X"69",X"00",X"85",X"D9",X"4C",X"06",X"F3",X"85",X"F5",X"6E",
		X"A5",X"E0",X"D0",X"45",X"A5",X"E2",X"29",X"10",X"4A",X"4A",X"4A",X"4A",X"18",X"69",X"43",X"8D",
		X"01",X"18",X"A5",X"E2",X"10",X"2A",X"C6",X"DC",X"F0",X"07",X"A9",X"47",X"D0",X"1C",X"85",X"F5",
		X"EA",X"E6",X"F3",X"A5",X"F3",X"C9",X"01",X"D0",X"08",X"A9",X"1E",X"8D",X"03",X"40",X"C1",X"F5",
		X"EA",X"A9",X"03",X"85",X"DC",X"4D",X"4C",X"85",X"F5",X"EA",X"8D",X"01",X"18",X"C1",X"F5",X"6E",
		X"A5",X"E2",X"49",X"10",X"85",X"E2",X"C1",X"F5",X"EA",X"60",X"85",X"F5",X"6E",X"AD",X"02",X"40",
		X"49",X"FF",X"29",X"03",X"F0",X"08",X"BA",X"E8",X"E8",X"9A",X"60",X"85",X"F5",X"6E",X"A5",X"E0",
		X"D0",X"42",X"A5",X"E2",X"29",X"E0",X"D0",X"3C",X"A6",X"CB",X"AD",X"03",X"40",X"29",X"40",X"D0",
		X"05",X"A2",X"00",X"85",X"F5",X"6E",X"BD",X"00",X"40",X"49",X"FF",X"29",X"0F",X"AA",X"BD",X"D5",
		X"F3",X"C5",X"EF",X"F0",X"1F",X"85",X"EF",X"14",X"65",X"EE",X"10",X"05",X"A9",X"00",X"85",X"F5",
		X"EA",X"C9",X"24",X"90",X"05",X"A9",X"23",X"85",X"F5",X"EA",X"85",X"EE",X"4D",X"15",X"8D",X"03",
		X"40",X"85",X"F5",X"EA",X"60",X"00",X"01",X"FF",X"00",X"F6",X"00",X"00",X"00",X"0A",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"85",X"F5",X"EA",X"A5",X"E2",X"29",X"E0",X"D0",X"32",
		X"A2",X"78",X"A5",X"EE",X"C9",X"1E",X"B0",X"11",X"A2",X"60",X"C9",X"14",X"B0",X"0B",X"A2",X"48",
		X"C9",X"0A",X"B0",X"05",X"A2",X"30",X"85",X"F5",X"EA",X"8E",X"03",X"18",X"A5",X"EE",X"38",X"85",
		X"F5",X"EA",X"E9",X"0A",X"B0",X"FC",X"69",X"0A",X"AA",X"BD",X"23",X"F4",X"8D",X"02",X"18",X"85",
		X"F5",X"EA",X"60",X"B4",X"A4",X"94",X"84",X"74",X"64",X"54",X"44",X"34",X"24",X"85",X"F5",X"EA",
		X"A5",X"E1",X"D0",X"4F",X"A5",X"E2",X"29",X"E0",X"D0",X"49",X"A6",X"CB",X"AD",X"03",X"40",X"29",
		X"40",X"D0",X"05",X"A2",X"00",X"85",X"F5",X"EA",X"BD",X"00",X"40",X"49",X"FF",X"29",X"10",X"F0",
		X"32",X"A5",X"E2",X"29",X"03",X"C9",X"03",X"F0",X"06",X"A9",X"11",X"8D",X"03",X"40",X"EA",X"A5",
		X"EE",X"C9",X"1E",X"90",X"22",X"38",X"E9",X"1E",X"0A",X"AA",X"BD",X"EB",X"F4",X"85",X"D8",X"BD",
		X"EC",X"F4",X"85",X"D9",X"A9",X"3F",X"85",X"E1",X"A9",X"17",X"8D",X"03",X"40",X"6C",X"D8",X"00",
		X"85",X"F5",X"EA",X"60",X"85",X"F5",X"EA",X"A5",X"E3",X"29",X"20",X"D0",X"F6",X"A9",X"60",X"85",
		X"D9",X"A6",X"EE",X"E0",X"1A",X"90",X"15",X"E0",X"1E",X"B0",X"11",X"8A",X"E9",X"18",X"AA",X"A9",
		X"50",X"85",X"D8",X"A9",X"66",X"85",X"D9",X"D0",X"0A",X"85",X"F5",X"EA",X"A9",X"50",X"85",X"D8",
		X"85",X"F5",X"EA",X"A5",X"D8",X"18",X"69",X"08",X"85",X"D8",X"A5",X"D9",X"69",X"00",X"85",X"D9",
		X"CA",X"10",X"F0",X"85",X"F5",X"EA",X"A9",X"E0",X"85",X"DA",X"A9",X"62",X"85",X"DB",X"20",X"4B",
		X"F5",X"20",X"35",X"F5",X"A9",X"01",X"8D",X"04",X"18",X"20",X"71",X"F5",X"A9",X"00",X"A8",X"91",
		X"D8",X"A5",X"E2",X"09",X"40",X"85",X"E2",X"85",X"F5",X"EA",X"60",X"FA",X"F4",X"FA",X"F4",X"16",
		X"F5",X"16",X"F5",X"0C",X"F5",X"0C",X"F5",X"85",X"F5",X"EA",X"A5",X"E3",X"29",X"20",X"D0",X"EA",
		X"A9",X"F5",X"85",X"EE",X"CA",X"ED",X"4C",X"09",X"F6",X"85",X"F5",X"EA",X"A5",X"E2",X"09",X"80",
		X"85",X"E2",X"60",X"85",X"F5",X"6E",X"A5",X"E2",X"29",X"0F",X"F0",X"16",X"C6",X"E2",X"4D",X"F5",
		X"85",X"EE",X"A6",X"ED",X"20",X"08",X"F6",X"A5",X"E3",X"09",X"40",X"29",X"DF",X"85",X"E3",X"C1",
		X"F5",X"EA",X"60",X"85",X"F5",X"6E",X"AD",X"02",X"18",X"38",X"E9",X"04",X"8D",X"06",X"18",X"CD",
		X"03",X"18",X"38",X"E9",X"08",X"8D",X"07",X"18",X"60",X"85",X"F5",X"EA",X"A2",X"02",X"85",X"F5",
		X"EA",X"A0",X"07",X"85",X"F5",X"6E",X"B1",X"D8",X"91",X"DA",X"88",X"10",X"F9",X"A5",X"D9",X"18",
		X"69",X"20",X"85",X"D9",X"C9",X"DB",X"18",X"69",X"20",X"85",X"DB",X"CA",X"10",X"E3",X"60",X"85",
		X"F5",X"EA",X"AD",X"07",X"18",X"85",X"D9",X"CD",X"06",X"18",X"49",X"FF",X"85",X"D8",X"A2",X"D9",
		X"46",X"D9",X"46",X"D9",X"A2",X"D9",X"AA",X"D8",X"46",X"D9",X"66",X"D8",X"A2",X"D9",X"AA",X"D8",
		X"A5",X"D9",X"18",X"69",X"10",X"85",X"D9",X"E2",X"D8",X"60",X"85",X"F5",X"6E",X"A5",X"E2",X"29",
		X"E0",X"C9",X"40",X"F0",X"04",X"60",X"85",X"F5",X"EA",X"A9",X"9B",X"85",X"D8",X"C9",X"E2",X"29",
		X"0F",X"F0",X"11",X"AA",X"85",X"F5",X"6E",X"A5",X"D8",X"38",X"E9",X"08",X"85",X"D8",X"66",X"D0",
		X"F6",X"85",X"F5",X"EA",X"A6",X"ED",X"BD",X"00",X"F6",X"85",X"D9",X"A5",X"D8",X"CD",X"02",X"18",
		X"F0",X"10",X"90",X"08",X"EE",X"02",X"18",X"70",X"09",X"85",X"F5",X"EA",X"CE",X"02",X"18",X"C1",
		X"F5",X"EA",X"A5",X"D9",X"CD",X"03",X"18",X"F0",X"0D",X"EE",X"03",X"18",X"C1",X"F5",X"6E",X"20",
		X"35",X"F5",X"60",X"85",X"F5",X"6E",X"A5",X"D8",X"CD",X"02",X"18",X"F0",X"0C",X"4C",X"EF",X"F5",
		X"00",X"A8",X"B8",X"C8",X"D8",X"E8",X"85",X"F5",X"EA",X"A5",X"E2",X"09",X"20",X"29",X"BF",X"85",
		X"E2",X"BD",X"84",X"F0",X"18",X"69",X"36",X"85",X"D8",X"A9",X"00",X"85",X"D9",X"A5",X"E2",X"29",
		X"0F",X"A8",X"A5",X"EE",X"C9",X"1A",X"90",X"0B",X"C9",X"1E",X"B0",X"07",X"69",X"B2",X"30",X"09",
		X"85",X"F5",X"EA",X"18",X"69",X"0B",X"85",X"F5",X"EA",X"91",X"D8",X"60",X"85",X"F5",X"EA",X"A5",
		X"E2",X"10",X"18",X"A9",X"D0",X"8D",X"02",X"18",X"A6",X"ED",X"BD",X"00",X"F6",X"38",X"E9",X"0C",
		X"8D",X"03",X"18",X"A9",X"00",X"8D",X"04",X"18",X"85",X"F5",X"EA",X"60",X"45",X"09",X"41",X"54",
		X"32",X"30",X"37",X"30",X"09",X"2F",X"20",X"4B",X"4F",X"52",X"45",X"4B",X"41",X"52",X"41",X"20",
		X"44",X"49",X"53",X"50",X"2E",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"0D",X"0A",X"09",X"4A",X"4D",X"50",X"09",X"41",X"54",X"32",X"30",X"33",X"30",X"0D",
		X"0A",X"0D",X"0A",X"09",X"53",X"54",X"41",X"09",X"44",X"55",X"4D",X"59",X"50",X"0D",X"0A",X"09",
		X"4E",X"4F",X"50",X"0D",X"0A",X"41",X"54",X"32",X"30",X"37",X"30",X"09",X"4C",X"44",X"58",X"09",
		X"23",X"3E",X"54",X"45",X"4B",X"4E",X"41",X"4D",X"20",X"20",X"20",X"20",X"2F",X"20",X"54",X"45",
		X"4B",X"49",X"20",X"4E",X"41",X"4D",X"45",X"20",X"44",X"49",X"53",X"50",X"4C",X"41",X"59",X"2E",
		X"20",X"53",X"54",X"4F",X"50",X"20",X"4D",X"4F",X"54",X"49",X"4F",X"4E",X"0D",X"0A",X"09",X"4C",
		X"44",X"59",X"09",X"23",X"3C",X"54",X"45",X"4B",X"4E",X"41",X"4D",X"0D",X"0A",X"09",X"4A",X"53",
		X"52",X"09",X"43",X"48",X"52",X"4F",X"55",X"54",X"2D",X"31",X"09",X"2F",X"20",X"44",X"49",X"53",
		X"50",X"4C",X"41",X"59",X"20",X"4F",X"55",X"54",X"0D",X"0A",X"09",X"09",X"09",X"2F",X"20",X"4D",
		X"52",X"2E",X"48",X"4F",X"54",X"20",X"44",X"4F",X"47",X"2C",X"4D",X"52",X"2E",X"50",X"49",X"43",
		X"4B",X"4C",X"45",X"2C",X"4D",X"52",X"2E",X"45",X"47",X"47",X"0D",X"0A",X"09",X"4C",X"44",X"58",
		X"09",X"23",X"30",X"46",X"46",X"0D",X"0A",X"09",X"4A",X"53",X"52",X"09",X"57",X"41",X"49",X"54",
		X"45",X"2D",X"31",X"09",X"20",X"20",X"20",X"20",X"20",X"20",X"0D",X"0A",X"09",X"4C",X"44",X"41",
		X"09",X"23",X"30",X"30",X"0D",X"0A",X"09",X"53",X"54",X"41",X"09",X"46",X"4C",X"47",X"46",X"4C",
		X"47",X"09",X"20",X"20",X"20",X"2F",X"20",X"4E",X"41",X"4D",X"45",X"20",X"44",X"49",X"53",X"50",
		X"2E",X"20",X"45",X"4E",X"44",X"0D",X"0A",X"09",X"4A",X"4D",X"50",X"09",X"41",X"54",X"32",X"30",
		X"30",X"30",X"0D",X"0A",X"0D",X"0A",X"54",X"45",X"4B",X"4E",X"41",X"4D",X"09",X"45",X"51",X"55",
		X"09",X"2E",X"0D",X"0A",X"09",X"44",X"46",X"41",X"09",X"31",X"31",X"38",X"36",X"09",X"09",X"2F",
		X"20",X"4D",X"52",X"2E",X"48",X"4F",X"54",X"44",X"4F",X"47",X"0D",X"0A",X"09",X"44",X"46",X"43",
		X"09",X"33",X"42",X"2C",X"34",X"30",X"2C",X"36",X"30",X"2C",X"33",X"36",X"2C",X"33",X"44",X"2C",
		X"34",X"32",X"2C",X"30",X"30",X"2C",X"33",X"32",X"0D",X"0A",X"09",X"44",X"46",X"43",X"09",X"33",
		X"44",X"2C",X"33",X"35",X"2C",X"36",X"31",X"2C",X"36",X"32",X"2C",X"30",X"46",X"45",X"0D",X"0A",
		X"09",X"44",X"46",X"41",X"09",X"31",X"35",X"38",X"36",X"0D",X"0A",X"09",X"44",X"46",X"43",X"09",
		X"30",X"30",X"2C",X"30",X"30",X"2C",X"30",X"30",X"2C",X"30",X"30",X"2C",X"30",X"30",X"2C",X"30",
		X"30",X"2C",X"30",X"30",X"2C",X"30",X"30",X"0D",X"0A",X"09",X"44",X"46",X"43",X"09",X"30",X"30",
		X"2C",X"30",X"30",X"2C",X"30",X"30",X"2C",X"30",X"30",X"2C",X"30",X"46",X"45",X"0D",X"0A",X"0D",
		X"0A",X"09",X"44",X"46",X"41",X"09",X"31",X"30",X"43",X"45",X"09",X"09",X"2F",X"20",X"4D",X"52",
		X"2E",X"50",X"49",X"43",X"4B",X"4C",X"45",X"0D",X"0A",X"09",X"44",X"46",X"43",X"09",X"33",X"42",
		X"2C",X"34",X"30",X"2C",X"36",X"30",X"2C",X"33",X"45",X"2C",X"33",X"37",X"2C",X"33",X"31",X"2C",
		X"33",X"39",X"2C",X"33",X"41",X"0D",X"0A",X"09",X"44",X"46",X"43",X"09",X"33",X"33",X"2C",X"36",
		X"31",X"2C",X"36",X"32",X"2C",X"30",X"46",X"45",X"0D",X"0A",X"09",X"44",X"46",X"41",X"09",X"31",
		X"34",X"43",X"45",X"0D",X"0A",X"09",X"44",X"46",X"43",X"09",X"30",X"30",X"2C",X"30",X"30",X"2C",
		X"30",X"30",X"2C",X"30",X"30",X"2C",X"30",X"30",X"2C",X"30",X"30",X"2C",X"30",X"30",X"2C",X"30",
		X"30",X"0D",X"0A",X"09",X"44",X"46",X"43",X"09",X"30",X"30",X"2C",X"30",X"30",X"2C",X"30",X"30",
		X"2C",X"30",X"46",X"45",X"0D",X"0A",X"0D",X"0A",X"09",X"44",X"46",X"41",X"09",X"31",X"31",X"35",
		X"36",X"09",X"09",X"2F",X"20",X"4D",X"52",X"2E",X"45",X"47",X"47",X"0D",X"0A",X"09",X"44",X"46",
		X"43",X"09",X"33",X"42",X"2C",X"34",X"30",X"2C",X"36",X"30",X"2C",X"33",X"33",X"2C",X"33",X"35",
		X"2C",X"33",X"35",X"2C",X"36",X"31",X"2C",X"36",X"32",X"2C",X"30",X"46",X"45",X"0D",X"0A",X"09",
		X"44",X"46",X"41",X"09",X"31",X"35",X"35",X"36",X"0D",X"0A",X"09",X"44",X"46",X"43",X"09",X"30",
		X"30",X"2C",X"30",X"30",X"2C",X"30",X"30",X"2C",X"30",X"30",X"2C",X"30",X"30",X"2C",X"30",X"30",
		X"2C",X"30",X"30",X"2C",X"30",X"30",X"2C",X"30",X"46",X"46",X"0D",X"0A",X"0D",X"0A",X"2F",X"0D",
		X"0A",X"2F",X"2A",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",
		X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",
		X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",
		X"2D",X"2A",X"0D",X"0A",X"2F",X"2A",X"09",X"50",X"45",X"50",X"50",X"45",X"52",X"20",X"26",X"20",
		X"54",X"45",X"4B",X"49",X"20",X"4C",X"41",X"4B",X"4B",X"41",X"20",X"41",X"54",X"52",X"41",X"43",
		X"54",X"49",X"4F",X"4E",X"09",X"09",X"2A",X"0D",X"0A",X"2F",X"2A",X"2D",X"2D",X"2D",X"2D",X"2D",
		X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",
		X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",
		X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"2A",X"0D",X"0A",X"2F",X"0D",X"0A",X"09",
		X"53",X"54",X"41",X"09",X"44",X"55",X"4D",X"59",X"50",X"09",X"2F",X"20",X"44",X"55",X"4D",X"4D",
		X"59",X"20",X"57",X"52",X"49",X"54",X"45",X"0D",X"0A",X"09",X"4E",X"4F",X"50",X"09",X"09",X"2F",
		X"20",X"44",X"55",X"4D",X"4D",X"59",X"20",X"4E",X"4F",X"50",X"0D",X"0A",X"41",X"54",X"52",X"43",
		X"54",X"33",X"09",X"45",X"51",X"55",X"09",X"2E",X"0D",X"0A",X"09",X"4A",X"53",X"52",X"09",X"47",
		X"41",X"4D",X"49",X"4E",X"4C",X"2D",X"31",X"0D",X"0A",X"09",X"4A",X"53",X"52",X"09",X"52",X"4E",
		X"44",X"49",X"4E",X"4C",X"2D",X"31",X"0D",X"0A",X"2F",X"0D",X"0A",X"09",X"4C",X"44",X"59",X"09",
		X"23",X"30",X"31",X"0D",X"0A",X"09",X"53",X"54",X"59",X"09",X"4C",X"49",X"56",X"45",X"2B",X"30",
		X"0D",X"0A",X"09",X"53",X"54",X"59",X"09",X"4C",X"49",X"56",X"45",X"2B",X"31",X"0D",X"0A",X"09",
		X"49",X"4E",X"59",X"0D",X"0A",X"09",X"53",X"54",X"59",X"09",X"4C",X"49",X"56",X"45",X"2B",X"32",
		X"0D",X"0A",X"09",X"53",X"54",X"59",X"09",X"4C",X"49",X"56",X"45",X"2B",X"33",X"0D",X"0A",X"09",
		X"49",X"4E",X"59",X"0D",X"0A",X"09",X"53",X"54",X"59",X"09",X"4C",X"49",X"56",X"45",X"2B",X"34",
		X"0D",X"0A",X"09",X"53",X"54",X"59",X"09",X"4C",X"49",X"56",X"45",X"2B",X"35",X"0D",X"0A",X"2F",
		X"0D",X"0A",X"09",X"4C",X"44",X"41",X"09",X"23",X"31",X"44",X"0D",X"0A",X"09",X"53",X"54",X"41",
		X"09",X"30",X"31",X"38",X"30",X"33",X"0D",X"0A",X"09",X"53",X"54",X"41",X"09",X"30",X"31",X"38",
		X"30",X"37",X"0D",X"0A",X"09",X"53",X"54",X"41",X"09",X"30",X"31",X"38",X"30",X"42",X"0D",X"0A",
		X"09",X"53",X"54",X"41",X"09",X"30",X"31",X"38",X"30",X"46",X"0D",X"0A",X"09",X"53",X"54",X"41",
		X"09",X"30",X"31",X"38",X"31",X"33",X"0D",X"0A",X"09",X"53",X"54",X"41",X"09",X"30",X"31",X"38",
		X"31",X"37",X"0D",X"0A",X"09",X"53",X"54",X"41",X"09",X"30",X"31",X"38",X"31",X"46",X"0D",X"0A",
		X"2F",X"0D",X"0A",X"09",X"4C",X"44",X"41",X"09",X"23",X"34",X"30",X"0D",X"0A",X"09",X"53",X"54",
		X"41",X"09",X"44",X"49",X"52",X"45",X"43",X"54",X"2B",X"30",X"0D",X"0A",X"09",X"53",X"54",X"41",
		X"09",X"44",X"49",X"52",X"45",X"43",X"54",X"2B",X"31",X"0D",X"0A",X"09",X"53",X"54",X"41",X"09",
		X"44",X"49",X"52",X"45",X"43",X"54",X"2B",X"32",X"0D",X"0A",X"09",X"53",X"54",X"41",X"09",X"44",
		X"49",X"52",X"45",X"43",X"54",X"2B",X"33",X"0D",X"0A",X"09",X"53",X"54",X"41",X"09",X"44",X"49",
		X"52",X"45",X"43",X"54",X"2B",X"34",X"0D",X"0A",X"09",X"53",X"54",X"41",X"09",X"44",X"49",X"52",
		X"45",X"43",X"54",X"2B",X"35",X"0D",X"0A",X"2F",X"0D",X"0A",X"09",X"4C",X"44",X"41",X"09",X"23",
		X"38",X"39",X"0D",X"0A",X"09",X"53",X"54",X"41",X"09",X"30",X"31",X"38",X"30",X"32",X"0D",X"0A",
		X"09",X"4C",X"44",X"41",X"09",X"23",X"35",X"39",X"0D",X"0A",X"09",X"53",X"54",X"41",X"09",X"30",
		X"31",X"38",X"30",X"36",X"0D",X"0A",X"09",X"4C",X"44",X"41",X"09",X"23",X"36",X"30",X"0D",X"0A",
		X"09",X"53",X"54",X"41",X"09",X"30",X"31",X"38",X"30",X"41",X"0D",X"0A",X"09",X"4C",X"44",X"41",
		X"09",X"23",X"39",X"30",X"0D",X"0A",X"09",X"53",X"54",X"41",X"09",X"30",X"31",X"38",X"30",X"45",
		X"0D",X"0A",X"09",X"4C",X"44",X"41",X"09",X"23",X"39",X"37",X"0D",X"0A",X"09",X"53",X"54",X"41",
		X"09",X"30",X"31",X"38",X"31",X"32",X"0D",X"0A",X"09",X"4C",X"44",X"41",X"09",X"23",X"33",X"30",
		X"0D",X"0A",X"09",X"53",X"54",X"41",X"09",X"30",X"31",X"38",X"31",X"36",X"0D",X"0A",X"09",X"4C",
		X"44",X"41",X"09",X"23",X"31",X"38",X"0D",X"0A",X"09",X"53",X"54",X"41",X"09",X"30",X"31",X"38",
		X"31",X"45",X"0D",X"0A",X"2F",X"09",X"0D",X"0A",X"09",X"4C",X"44",X"41",X"09",X"23",X"30",X"31",
		X"0D",X"0A",X"09",X"53",X"54",X"41",X"09",X"54",X"49",X"4D",X"45",X"52",X"31",X"0D",X"0A",X"09",
		X"53",X"54",X"41",X"09",X"54",X"49",X"4D",X"45",X"52",X"32",X"0D",X"0A",X"2F",X"0D",X"0A",X"09",
		X"4A",X"53",X"52",X"09",X"54",X"45",X"4B",X"4D",X"4F",X"56",X"2D",X"31",X"09",X"2F",X"20",X"54",
		X"45",X"4B",X"49",X"20",X"44",X"49",X"53",X"50",X"4C",X"41",X"59",X"0D",X"0A",X"2F",X"0D",X"0A",
		X"09",X"53",X"54",X"41",X"09",X"44",X"55",X"4D",X"59",X"50",X"09",X"2F",X"20",X"44",X"55",X"4D",
		X"4D",X"59",X"20",X"57",X"52",X"49",X"54",X"45",X"0D",X"0A",X"09",X"4E",X"4F",X"50",X"09",X"09",
		X"2F",X"20",X"44",X"55",X"4D",X"4D",X"59",X"20",X"4E",X"4F",X"50",X"0D",X"0A",X"41",X"54",X"33",
		X"30",X"33",X"30",X"09",X"45",X"51",X"55",X"09",X"2E",X"0D",X"0A",X"09",X"4C",X"44",X"58",X"09",
		X"23",X"30",X"31",X"0D",X"0A",X"09",X"4A",X"53",X"52",X"09",X"57",X"41",X"49",X"54",X"45",X"2D",
		X"31",X"0D",X"0A",X"09",X"49",X"4E",X"43",X"09",X"54",X"49",X"4D",X"45",X"52",X"31",X"0D",X"0A",
		X"09",X"42",X"4E",X"45",X"09",X"2E",X"2B",X"35",X"0D",X"0A",X"09",X"49",X"4E",X"43",X"09",X"54",
		X"49",X"4D",X"45",X"52",X"32",X"0D",X"0A",X"09",X"4E",X"4F",X"50",X"0D",X"0A",X"2F",X"0D",X"0A",
		X"09",X"4C",X"44",X"58",X"09",X"23",X"30",X"37",X"0D",X"0A",X"09",X"4A",X"53",X"52",X"09",X"4C",
		X"49",X"4D",X"49",X"54",X"2D",X"31",X"0D",X"0A",X"09",X"42",X"45",X"51",X"09",X"41",X"54",X"33",
		X"30",X"34",X"30",X"0D",X"0A",X"09",X"4C",X"44",X"41",X"09",X"54",X"49",X"4D",X"45",X"52",X"32",
		X"0D",X"0A",X"09",X"43",X"4D",X"50",X"09",X"23",X"30",X"34",X"0D",X"0A",X"09",X"42",X"43",X"43",
		X"09",X"41",X"54",X"33",X"30",X"36",X"30",X"0D",X"0A",X"09",X"0D",X"0A",X"09",X"4C",X"44",X"58",
		X"09",X"23",X"3E",X"50",X"45",X"50",X"4D",X"53",X"47",X"0D",X"0A",X"09",X"4C",X"44",X"59",X"09",
		X"23",X"3C",X"50",X"45",X"50",X"4D",X"53",X"47",X"0D",X"0A",X"09",X"4A",X"53",X"52",X"09",X"43",
		X"48",X"52",X"4F",X"55",X"54",X"2D",X"31",X"20",X"20",X"20",X"2F",X"20",X"50",X"45",X"50",X"50",
		X"45",X"52",X"20",X"53",X"45",X"54",X"53",X"55",X"4D",X"45",X"49",X"20",X"44",X"49",X"53",X"50",
		X"4C",X"41",X"59",X"0D",X"0A",X"09",X"4C",X"44",X"58",X"09",X"23",X"30",X"46",X"46",X"0D",X"0A",
		X"09",X"4A",X"53",X"52",X"09",X"57",X"41",X"49",X"54",X"45",X"2D",X"31",X"0D",X"0A",X"09",X"4C",
		X"44",X"58",X"09",X"23",X"30",X"34",X"30",X"0D",X"0A",X"09",X"4A",X"53",X"52",X"09",X"57",X"41",
		X"49",X"54",X"45",X"2D",X"31",X"0D",X"0A",X"09",X"52",X"54",X"53",X"0D",X"0A",X"0D",X"0A",X"09",
		X"53",X"54",X"41",X"09",X"44",X"55",X"4D",X"59",X"50",X"09",X"2F",X"20",X"44",X"55",X"4D",X"4D",
		X"59",X"20",X"57",X"52",X"49",X"54",X"45",X"0D",X"0A",X"09",X"4E",X"4F",X"50",X"09",X"09",X"2F",
		X"20",X"44",X"55",X"4D",X"4D",X"59",X"20",X"4E",X"4F",X"50",X"0D",X"0A",X"41",X"54",X"33",X"30",
		X"34",X"30",X"09",X"4C",X"44",X"41",X"09",X"4C",X"49",X"56",X"45",X"2B",X"36",X"0D",X"0A",X"09",
		X"42",X"50",X"4C",X"09",X"41",X"54",X"33",X"30",X"36",X"30",X"0D",X"0A",X"20",X"20",X"20",X"20",
		X"20",X"20",X"09",X"4C",X"44",X"58",X"09",X"23",X"30",X"37",X"0D",X"0A",X"09",X"4A",X"53",X"52",
		X"09",X"53",X"50",X"52",X"4D",X"4F",X"56",X"2D",X"31",X"0D",X"0A",X"2F",X"0D",X"0A",X"09",X"4C",
		X"44",X"41",X"09",X"30",X"31",X"38",X"31",X"45",X"0D",X"0A",X"09",X"43",X"4D",X"50",X"09",X"23",
		X"32",X"32",X"0D",X"0A",X"09",X"42",X"45",X"51",X"09",X"41",X"54",X"33",X"30",X"35",X"30",X"09",
		X"2F",X"20",X"50",X"45",X"50",X"50",X"45",X"52",X"20",X"4F",X"4E",X"0D",X"0A",X"09",X"43",X"4D",
		X"50",X"09",X"23",X"34",X"41",X"0D",X"0A",X"09",X"42",X"45",X"51",X"09",X"41",X"54",X"33",X"30",
		X"35",X"30",X"0D",X"0A",X"09",X"43",X"4D",X"50",X"09",X"23",X"38",X"32",X"0D",X"0A",X"09",X"42",
		X"4E",X"45",X"09",X"41",X"54",X"33",X"30",X"36",X"30",X"0D",X"0A",X"09",X"53",X"54",X"41",X"09",
		X"44",X"55",X"4D",X"59",X"50",X"09",X"2F",X"20",X"44",X"55",X"4D",X"4D",X"59",X"20",X"57",X"52",
		X"49",X"54",X"45",X"0D",X"0A",X"09",X"4E",X"4F",X"50",X"09",X"09",X"2F",X"20",X"44",X"55",X"4D",
		X"4D",X"59",X"20",X"4E",X"4F",X"50",X"0D",X"0A",X"41",X"54",X"33",X"30",X"35",X"30",X"09",X"4A",
		X"53",X"52",X"09",X"43",X"4F",X"4B",X"50",X"50",X"53",X"2D",X"31",X"09",X"2F",X"20",X"50",X"45",
		X"50",X"50",X"45",X"52",X"20",X"53",X"45",X"54",X"0D",X"0A",X"09",X"49",X"4E",X"43",X"09",X"30",
		X"31",X"38",X"31",X"45",X"0D",X"0A",X"09",X"49",X"4E",X"43",X"09",X"30",X"31",X"38",X"31",X"45",
		X"0D",X"0A",X"09",X"53",X"54",X"41",X"09",X"44",X"55",X"4D",X"59",X"50",X"09",X"2F",X"20",X"44",
		X"55",X"4D",X"4D",X"59",X"20",X"57",X"52",X"49",X"54",X"45",X"0D",X"0A",X"09",X"4E",X"4F",X"50",
		X"09",X"09",X"2F",X"20",X"44",X"55",X"4D",X"4D",X"59",X"20",X"4E",X"4F",X"50",X"0D",X"0A",X"41",
		X"54",X"33",X"30",X"36",X"30",X"09",X"4A",X"53",X"52",X"09",X"43",X"4F",X"4B",X"50",X"45",X"50",
		X"2D",X"31",X"0D",X"0A",X"09",X"4A",X"53",X"52",X"09",X"4B",X"41",X"54",X"41",X"4D",X"4B",X"2D",
		X"31",X"0D",X"0A",X"09",X"4A",X"53",X"52",X"09",X"50",X"50",X"54",X"4B",X"50",X"54",X"2D",X"31",
		X"0D",X"0A",X"09",X"4A",X"53",X"52",X"09",X"4C",X"41",X"4B",X"4D",X"4F",X"56",X"2D",X"31",X"0D",
		X"0A",X"09",X"4A",X"4D",X"50",X"09",X"41",X"54",X"33",X"30",X"33",X"30",X"0D",X"0A",X"0D",X"0A",
		X"2F",X"50",X"45",X"50",X"50",X"45",X"52",X"20",X"4D",X"45",X"53",X"53",X"41",X"47",X"45",X"20",
		X"54",X"41",X"42",X"4C",X"45",X"0D",X"0A",X"2F",X"09",X"4D",X"45",X"53",X"53",X"41",X"47",X"45",
		X"20",X"20",X"3A",X"20",X"20",X"44",X"4F",X"4E",X"27",X"54",X"20",X"57",X"41",X"53",X"54",X"45",
		X"20",X"50",X"45",X"50",X"50",X"45",X"52",X"53",X"0D",X"0A",X"09",X"09",X"2F",X"20",X"20",X"20",
		X"59",X"4F",X"55",X"20",X"53",X"54",X"41",X"52",X"54",X"20",X"57",X"49",X"54",X"48",X"20",X"4F",
		X"4E",X"4C",X"59",X"20",X"46",X"49",X"56",X"45",X"0D",X"0A",X"09",X"09",X"2F",X"20",X"20",X"20",
		X"45",X"41",X"52",X"4E",X"20",X"45",X"58",X"54",X"52",X"41",X"20",X"50",X"45",X"50",X"50",X"45",
		X"52",X"53",X"20",X"26",X"20",X"42",X"4F",X"4E",X"55",X"53",X"45",X"53",X"0D",X"0A",X"09",X"09",
		X"2F",X"20",X"20",X"20",X"43",X"4C",X"41",X"49",X"4D",X"20",X"43",X"4F",X"4E",X"45",X"53",X"2C",
		X"43",X"4F",X"46",X"46",X"45",X"45",X"53",X"20",X"26",X"20",X"46",X"52",X"49",X"45",X"53",X"0D",
		X"0A",X"0D",X"0A",X"50",X"45",X"50",X"4D",X"53",X"47",X"09",X"45",X"51",X"55",X"09",X"2E",X"09",
		X"2F",X"20",X"44",X"4F",X"4E",X"27",X"54",X"2E",X"2E",X"2E",X"2E",X"2E",X"0D",X"0A",X"09",X"44",
		X"46",X"41",X"09",X"30",X"31",X"30",X"43",X"37",X"0D",X"0A",X"09",X"44",X"46",X"43",X"09",X"33",
		X"32",X"2C",X"33",X"44",X"2C",X"33",X"43",X"2C",X"36",X"34",X"2C",X"34",X"32",X"2C",X"30",X"30",
		X"2C",X"34",X"35",X"2C",X"32",X"46",X"0D",X"0A",X"09",X"44",X"00",X"C0",X"03",X"C0",X"00",X"C0");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
