library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity mw02 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of mw02 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"3D",X"32",X"51",X"20",X"F2",X"18",X"08",X"E6",X"0F",X"32",X"51",X"20",X"F3",X"2A",X"3B",X"20",
		X"2B",X"22",X"3B",X"20",X"FB",X"C3",X"18",X"08",X"CD",X"79",X"0A",X"E6",X"F0",X"CA",X"4E",X"08",
		X"21",X"51",X"20",X"35",X"EE",X"10",X"CA",X"2E",X"08",X"EE",X"30",X"CA",X"3E",X"08",X"2A",X"49",
		X"20",X"7C",X"FE",X"28",X"DA",X"4E",X"08",X"25",X"22",X"49",X"20",X"C3",X"4E",X"08",X"2A",X"49",
		X"20",X"7C",X"FE",X"E0",X"D2",X"4E",X"08",X"24",X"22",X"49",X"20",X"C3",X"4E",X"08",X"AF",X"32",
		X"4F",X"20",X"CD",X"1C",X"0A",X"DF",X"01",X"3A",X"52",X"20",X"A7",X"CA",X"AF",X"07",X"01",X"00",
		X"10",X"21",X"E8",X"20",X"7E",X"A7",X"CA",X"6C",X"08",X"F2",X"78",X"08",X"23",X"23",X"23",X"23",
		X"0C",X"05",X"C2",X"64",X"08",X"C3",X"AF",X"07",X"E5",X"C5",X"57",X"79",X"21",X"68",X"20",X"87",
		X"87",X"87",X"CD",X"2D",X"02",X"7E",X"FE",X"28",X"D2",X"A1",X"08",X"23",X"5E",X"3A",X"4A",X"20",
		X"C6",X"02",X"47",X"C6",X"0A",X"BB",X"DA",X"A1",X"08",X"23",X"23",X"7B",X"86",X"B8",X"D2",X"A6",
		X"08",X"C1",X"E1",X"C3",X"6C",X"08",X"7A",X"FE",X"40",X"CA",X"98",X"09",X"E6",X"F0",X"87",X"B1",
		X"3C",X"32",X"2C",X"20",X"3E",X"3F",X"32",X"0A",X"20",X"7A",X"FE",X"40",X"C1",X"E1",X"36",X"00",
		X"11",X"24",X"FA",X"FA",X"D1",X"08",X"FE",X"70",X"11",X"E0",X"FC",X"DA",X"D1",X"08",X"11",X"30",
		X"F8",X"2A",X"3B",X"20",X"19",X"7C",X"A7",X"FA",X"4A",X"09",X"3E",X"04",X"EF",X"0A",X"3E",X"20",
		X"EF",X"0B",X"DF",X"03",X"AF",X"32",X"66",X"20",X"D5",X"CD",X"50",X"0A",X"2A",X"49",X"20",X"3A",
		X"51",X"20",X"3D",X"32",X"51",X"20",X"0F",X"DA",X"FF",X"08",X"25",X"25",X"C3",X"01",X"09",X"24",
		X"24",X"22",X"49",X"20",X"CD",X"1C",X"0A",X"D1",X"2A",X"3B",X"20",X"2B",X"2B",X"2B",X"2B",X"2B",
		X"2B",X"00",X"00",X"22",X"3B",X"20",X"13",X"13",X"13",X"13",X"13",X"13",X"00",X"00",X"7A",X"A7",
		X"FA",X"E2",X"08",X"06",X"01",X"3E",X"04",X"F7",X"0A",X"3E",X"20",X"F7",X"0B",X"3E",X"01",X"32",
		X"30",X"20",X"AF",X"32",X"0A",X"20",X"78",X"E6",X"02",X"C2",X"43",X"09",X"3A",X"48",X"20",X"A7",
		X"F2",X"AF",X"07",X"78",X"32",X"2A",X"20",X"CD",X"C0",X"01",X"22",X"3B",X"20",X"3E",X"04",X"EF",
		X"0A",X"3E",X"20",X"EF",X"0B",X"2A",X"49",X"20",X"11",X"FE",X"FD",X"19",X"22",X"49",X"20",X"21",
		X"05",X"17",X"22",X"4B",X"20",X"21",X"54",X"1C",X"22",X"4D",X"20",X"CD",X"1C",X"0A",X"3E",X"64",
		X"32",X"51",X"20",X"21",X"51",X"20",X"35",X"CA",X"7F",X"09",X"DF",X"01",X"C3",X"73",X"09",X"06",
		X"03",X"C3",X"25",X"09",X"06",X"83",X"C3",X"25",X"09",X"3E",X"7F",X"32",X"0A",X"20",X"AF",X"32",
		X"2E",X"20",X"11",X"18",X"FC",X"C3",X"D1",X"08",X"C1",X"E1",X"CD",X"FC",X"09",X"DF",X"01",X"CD",
		X"50",X"0A",X"21",X"18",X"8A",X"22",X"49",X"20",X"CD",X"1C",X"0A",X"DF",X"01",X"3E",X"02",X"32",
		X"2D",X"20",X"3E",X"10",X"EF",X"0A",X"11",X"DC",X"05",X"DB",X"02",X"E6",X"08",X"CA",X"C3",X"09",
		X"11",X"E8",X"03",X"2A",X"3B",X"20",X"23",X"23",X"23",X"23",X"23",X"23",X"22",X"3B",X"20",X"E5",
		X"D5",X"CD",X"1C",X"0A",X"D1",X"E1",X"DF",X"02",X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",X"7A",X"A7",
		X"F2",X"C3",X"09",X"3E",X"10",X"F7",X"0A",X"3E",X"80",X"32",X"2D",X"20",X"3C",X"32",X"30",X"20",
		X"DF",X"01",X"3A",X"2D",X"20",X"A7",X"C2",X"F0",X"09",X"C3",X"AF",X"07",X"21",X"8F",X"19",X"11",
		X"AD",X"1B",X"3A",X"FC",X"1F",X"86",X"23",X"47",X"7D",X"AB",X"C2",X"12",X"0A",X"7C",X"AA",X"CA",
		X"16",X"0A",X"78",X"C3",X"05",X"0A",X"78",X"A7",X"C8",X"C3",X"30",X"0A",X"2A",X"49",X"20",X"CD",
		X"70",X"15",X"EB",X"2A",X"4B",X"20",X"E5",X"2A",X"4D",X"20",X"C1",X"EB",X"AF",X"32",X"52",X"20",
		X"E5",X"C5",X"1A",X"A6",X"CA",X"3A",X"0A",X"32",X"52",X"20",X"1A",X"B6",X"77",X"13",X"23",X"0D",
		X"C2",X"32",X"0A",X"C1",X"05",X"E1",X"C8",X"D5",X"11",X"20",X"00",X"19",X"D1",X"C3",X"30",X"0A",
		X"2A",X"49",X"20",X"CD",X"70",X"15",X"EB",X"2A",X"4B",X"20",X"E5",X"2A",X"4D",X"20",X"C1",X"EB",
		X"E5",X"C5",X"00",X"1A",X"AE",X"77",X"23",X"13",X"0D",X"C2",X"62",X"0A",X"C1",X"E1",X"05",X"C8",
		X"D5",X"11",X"20",X"00",X"19",X"D1",X"C3",X"60",X"0A",X"3A",X"48",X"20",X"A7",X"CA",X"9A",X"0A",
		X"F2",X"91",X"0A",X"0F",X"DA",X"91",X"0A",X"DB",X"00",X"07",X"07",X"47",X"DB",X"02",X"C3",X"96",
		X"0A",X"DB",X"00",X"47",X"DB",X"01",X"0F",X"E6",X"38",X"C9",X"3A",X"5B",X"20",X"C6",X"10",X"07",
		X"E6",X"38",X"C9",X"AF",X"32",X"5C",X"20",X"32",X"64",X"20",X"3E",X"64",X"32",X"66",X"20",X"3E",
		X"20",X"32",X"65",X"20",X"3E",X"01",X"32",X"5F",X"20",X"3A",X"2C",X"20",X"A7",X"C2",X"8D",X"0C",
		X"3A",X"E8",X"20",X"FE",X"40",X"CA",X"9F",X"0C",X"3E",X"0F",X"F7",X"0C",X"3A",X"58",X"20",X"A7",
		X"CA",X"FA",X"0A",X"21",X"66",X"20",X"35",X"C2",X"DF",X"0A",X"36",X"64",X"C3",X"14",X"0B",X"CD",
		X"DC",X"0C",X"DF",X"01",X"C3",X"B9",X"0A",X"CD",X"79",X"0A",X"E6",X"08",X"C2",X"3E",X"0B",X"3A",
		X"5C",X"20",X"E6",X"01",X"32",X"5C",X"20",X"C3",X"3E",X"0B",X"CD",X"79",X"0A",X"E6",X"08",X"C2",
		X"0D",X"0B",X"3A",X"5C",X"20",X"E6",X"01",X"32",X"5C",X"20",X"C3",X"DF",X"0A",X"3A",X"5C",X"20",
		X"A7",X"C2",X"DF",X"0A",X"3A",X"0A",X"20",X"E6",X"FF",X"C2",X"DF",X"0A",X"3E",X"03",X"32",X"5C",
		X"20",X"3E",X"02",X"EF",X"0A",X"3E",X"08",X"32",X"67",X"20",X"F3",X"2A",X"3B",X"20",X"2B",X"2B",
		X"22",X"3B",X"20",X"FB",X"2A",X"49",X"20",X"11",X"10",X"07",X"19",X"C3",X"66",X"0B",X"CD",X"DC",
		X"0C",X"DF",X"01",X"11",X"05",X"0D",X"06",X"01",X"2A",X"5D",X"20",X"CD",X"DD",X"15",X"21",X"67",
		X"20",X"35",X"C2",X"59",X"0B",X"3E",X"02",X"F7",X"0A",X"2A",X"5D",X"20",X"2C",X"2C",X"2C",X"2C",
		X"7D",X"FE",X"D8",X"D2",X"D7",X"0B",X"22",X"5D",X"20",X"11",X"05",X"0D",X"06",X"01",X"CD",X"A0",
		X"15",X"DF",X"01",X"79",X"A7",X"CA",X"E7",X"0A",X"01",X"00",X"10",X"21",X"E8",X"20",X"7E",X"A7",
		X"CA",X"86",X"0B",X"F2",X"94",X"0B",X"23",X"23",X"23",X"23",X"0C",X"05",X"C2",X"7E",X"0B",X"DF",
		X"01",X"C3",X"E7",X"0A",X"FE",X"40",X"CA",X"E7",X"0A",X"E5",X"C5",X"57",X"79",X"21",X"68",X"20",
		X"87",X"87",X"87",X"CD",X"2D",X"02",X"D5",X"EB",X"2A",X"5D",X"20",X"EB",X"1C",X"1C",X"1C",X"7B",
		X"4E",X"B9",X"DA",X"D1",X"0B",X"23",X"7A",X"46",X"B8",X"DA",X"D1",X"0B",X"23",X"23",X"23",X"7E",
		X"87",X"87",X"87",X"81",X"BB",X"DA",X"D1",X"0B",X"23",X"7E",X"E6",X"1F",X"80",X"BA",X"D2",X"E2",
		X"0B",X"D1",X"C1",X"E1",X"C3",X"86",X"0B",X"3A",X"5C",X"20",X"E6",X"FE",X"32",X"5C",X"20",X"C3",
		X"E2",X"0A",X"D1",X"C1",X"E1",X"7A",X"FE",X"40",X"06",X"00",X"D2",X"F8",X"0B",X"3A",X"3D",X"20",
		X"E6",X"07",X"47",X"3A",X"3F",X"20",X"80",X"47",X"7A",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"57",
		X"59",X"21",X"08",X"0D",X"CD",X"2D",X"02",X"80",X"4F",X"06",X"00",X"2A",X"41",X"20",X"09",X"22",
		X"41",X"20",X"3A",X"64",X"20",X"A7",X"CA",X"26",X"0C",X"D5",X"2A",X"63",X"20",X"44",X"4D",X"2A",
		X"5F",X"20",X"CD",X"7F",X"15",X"D1",X"7B",X"21",X"E8",X"20",X"87",X"87",X"CD",X"2D",X"02",X"36",
		X"00",X"7A",X"FE",X"04",X"D2",X"81",X"0C",X"3E",X"08",X"EF",X"0A",X"7B",X"87",X"87",X"87",X"21",
		X"68",X"20",X"CD",X"2D",X"02",X"D6",X"02",X"4F",X"23",X"7E",X"D6",X"02",X"47",X"C5",X"7A",X"87",
		X"87",X"21",X"10",X"0D",X"CD",X"2D",X"02",X"5F",X"23",X"56",X"23",X"4E",X"23",X"46",X"21",X"64",
		X"20",X"70",X"2B",X"71",X"2B",X"72",X"2B",X"73",X"E1",X"22",X"5F",X"20",X"3A",X"5C",X"20",X"E6",
		X"FE",X"32",X"5C",X"20",X"DF",X"01",X"CD",X"25",X"15",X"3E",X"32",X"32",X"65",X"20",X"C3",X"E2",
		X"0A",X"FE",X"05",X"C2",X"3B",X"0C",X"3E",X"17",X"E7",X"0B",X"C3",X"3B",X"0C",X"3D",X"57",X"E6",
		X"1F",X"4F",X"7A",X"1F",X"57",X"AF",X"32",X"2C",X"20",X"32",X"66",X"20",X"C3",X"E5",X"0B",X"21",
		X"65",X"20",X"35",X"F2",X"D0",X"0C",X"36",X"20",X"3A",X"64",X"20",X"3C",X"FE",X"04",X"C2",X"B3",
		X"0C",X"3E",X"00",X"32",X"64",X"20",X"3E",X"0F",X"F7",X"0C",X"3A",X"2D",X"20",X"E6",X"02",X"C2",
		X"D0",X"0C",X"21",X"D8",X"0C",X"3A",X"64",X"20",X"3D",X"E6",X"03",X"CD",X"2D",X"02",X"EF",X"0C",
		X"CD",X"DC",X"0C",X"DF",X"01",X"C3",X"B9",X"0A",X"01",X"04",X"02",X"08",X"3A",X"64",X"20",X"A7",
		X"C8",X"21",X"65",X"20",X"35",X"C0",X"2B",X"46",X"36",X"00",X"2B",X"4E",X"2B",X"2B",X"2B",X"7E",
		X"2B",X"6E",X"67",X"CD",X"7F",X"15",X"3E",X"08",X"F7",X"0A",X"3A",X"35",X"20",X"FE",X"17",X"C0",
		X"3E",X"1F",X"E7",X"0B",X"C9",X"0F",X"00",X"00",X"10",X"20",X"30",X"40",X"05",X"06",X"00",X"80",
		X"19",X"1C",X"02",X"13",X"19",X"1C",X"02",X"13",X"19",X"1C",X"02",X"13",X"19",X"1C",X"02",X"13",
		X"3F",X"1C",X"01",X"0C",X"3F",X"1C",X"01",X"0C",X"4A",X"1C",X"02",X"07",X"02",X"4F",X"05",X"28",
		X"21",X"2D",X"20",X"7E",X"A7",X"36",X"00",X"C2",X"5C",X"0E",X"3A",X"48",X"20",X"A7",X"C4",X"37",
		X"0F",X"21",X"E8",X"20",X"06",X"40",X"CD",X"40",X"00",X"CD",X"4F",X"0D",X"C3",X"66",X"0D",X"3E",
		X"DF",X"F7",X"0A",X"F7",X"0B",X"F7",X"0C",X"3A",X"40",X"20",X"E6",X"07",X"C8",X"FE",X"06",X"F0",
		X"3E",X"15",X"C3",X"DA",X"0F",X"0A",X"DF",X"01",X"3A",X"40",X"20",X"87",X"87",X"21",X"7F",X"0D",
		X"CD",X"2D",X"02",X"5F",X"23",X"56",X"23",X"7E",X"23",X"66",X"6F",X"E9",X"06",X"06",X"08",X"49",
		X"0D",X"49",X"0D",X"03",X"0F",X"58",X"0E",X"19",X"0F",X"58",X"0E",X"20",X"0F",X"58",X"0E",X"0C",
		X"0F",X"58",X"0E",X"30",X"0F",X"58",X"0E",X"FA",X"0E",X"58",X"0E",X"FD",X"0E",X"58",X"0E",X"00",
		X"0F",X"6C",X"0E",X"CF",X"0E",X"58",X"0E",X"D8",X"0E",X"58",X"0E",X"DF",X"0E",X"58",X"0E",X"EA",
		X"0E",X"58",X"0E",X"F3",X"0E",X"58",X"0E",X"FA",X"0E",X"58",X"0E",X"FD",X"0E",X"58",X"0E",X"00",
		X"0F",X"6C",X"0E",X"03",X"0F",X"58",X"0E",X"0C",X"0F",X"58",X"0E",X"10",X"0F",X"58",X"0E",X"19",
		X"0F",X"58",X"0E",X"20",X"0F",X"58",X"0E",X"FA",X"0E",X"58",X"0E",X"FD",X"0E",X"58",X"0E",X"00",
		X"0F",X"6C",X"0E",X"29",X"0F",X"58",X"0E",X"20",X"0F",X"58",X"0E",X"EA",X"0E",X"58",X"0E",X"03",
		X"0F",X"58",X"0E",X"0C",X"0F",X"58",X"0E",X"FA",X"0E",X"58",X"0E",X"FD",X"0E",X"58",X"0E",X"00",
		X"0F",X"6C",X"0E",X"7E",X"3C",X"C8",X"3D",X"23",X"32",X"2A",X"21",X"7E",X"23",X"E5",X"CD",X"43",
		X"0F",X"E1",X"C3",X"03",X"0E",X"AF",X"32",X"29",X"21",X"3D",X"32",X"2A",X"21",X"3E",X"06",X"C3",
		X"26",X"0E",X"0D",X"CD",X"2D",X"02",X"32",X"28",X"21",X"CD",X"ED",X"0F",X"3A",X"2A",X"21",X"FE",
		X"10",X"F0",X"21",X"28",X"21",X"35",X"C2",X"29",X"0E",X"DF",X"01",X"C3",X"1D",X"0E",X"DF",X"01",
		X"3A",X"29",X"21",X"A7",X"C0",X"3A",X"40",X"20",X"3C",X"32",X"40",X"20",X"FE",X"21",X"DA",X"56",
		X"0E",X"3E",X"01",X"32",X"40",X"20",X"AF",X"C9",X"EB",X"CD",X"03",X"0E",X"CD",X"15",X"0E",X"CD",
		X"3E",X"0E",X"C2",X"5C",X"0E",X"AF",X"32",X"2D",X"20",X"C3",X"49",X"0D",X"EB",X"3E",X"80",X"32",
		X"2B",X"21",X"CD",X"03",X"0E",X"CD",X"15",X"0E",X"3A",X"2D",X"20",X"E6",X"02",X"C2",X"90",X"0E",
		X"21",X"2B",X"21",X"35",X"CA",X"BD",X"0E",X"CD",X"3E",X"0E",X"C2",X"75",X"0E",X"C3",X"49",X"0D",
		X"DF",X"01",X"CD",X"15",X"0E",X"21",X"26",X"32",X"06",X"08",X"3E",X"AA",X"CD",X"41",X"00",X"DF",
		X"01",X"CD",X"15",X"0E",X"21",X"26",X"32",X"06",X"08",X"3E",X"55",X"CD",X"41",X"00",X"3A",X"2D",
		X"20",X"A7",X"F2",X"90",X"0E",X"21",X"26",X"32",X"06",X"08",X"CD",X"40",X"00",X"21",X"E9",X"20",
		X"06",X"08",X"36",X"00",X"23",X"23",X"23",X"23",X"05",X"C2",X"C2",X"0E",X"C3",X"5C",X"0E",X"00",
		X"00",X"01",X"01",X"02",X"02",X"03",X"03",X"FF",X"00",X"04",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"05",X"01",X"06",X"02",X"07",X"03",X"08",X"04",X"09",X"FF",X"00",X"0B",X"01",X"0C",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"00",X"0D",X"01",X"0E",X"02",X"0F",X"FF",X"00",X"0A",X"FF",X"00",X"13",X"FF",
		X"00",X"12",X"FF",X"00",X"10",X"01",X"11",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"18",X"FF",X"FF",
		X"00",X"16",X"01",X"17",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"19",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"14",X"01",X"15",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"1A",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"1B",X"FF",X"FF",X"FF",X"FF",X"FF",X"21",X"DB",X"17",X"11",X"8F",X"19",X"3A",X"FD",X"1F",
		X"C3",X"05",X"0A",X"87",X"21",X"00",X"40",X"CD",X"2D",X"02",X"5F",X"23",X"56",X"3A",X"2A",X"21",
		X"21",X"68",X"20",X"87",X"87",X"87",X"CD",X"2D",X"02",X"06",X"06",X"3A",X"40",X"20",X"EE",X"07",
		X"4F",X"E6",X"07",X"C2",X"77",X"0F",X"79",X"D6",X"08",X"F2",X"6E",X"0F",X"3E",X"18",X"4F",X"05",
		X"1A",X"91",X"91",X"00",X"77",X"13",X"23",X"CD",X"34",X"16",X"21",X"E8",X"20",X"3A",X"2A",X"21",
		X"87",X"87",X"CD",X"2D",X"02",X"1A",X"13",X"77",X"47",X"78",X"FE",X"38",X"C2",X"96",X"0F",X"3E",
		X"01",X"EF",X"0A",X"C3",X"E3",X"0F",X"78",X"FE",X"33",X"C2",X"A3",X"0F",X"3E",X"01",X"E7",X"0B",
		X"C3",X"12",X"4D",X"78",X"FE",X"70",X"C2",X"BC",X"0F",X"3E",X"10",X"EF",X"0C",X"D5",X"E5",X"21",
		X"AD",X"1B",X"11",X"E0",X"1F",X"3E",X"A3",X"C3",X"EB",X"4F",X"19",X"4D",X"78",X"FE",X"50",X"C2",
		X"CD",X"0F",X"3E",X"01",X"EF",X"0A",X"3E",X"1F",X"E7",X"0B",X"C3",X"E3",X"0F",X"78",X"FE",X"3F",
		X"C2",X"E5",X"0F",X"3E",X"1F",X"E7",X"0B",X"C3",X"12",X"4D",X"E7",X"0B",X"3E",X"01",X"EF",X"0A",
		X"C9",X"4F",X"4F",X"DF",X"01",X"23",X"36",X"00",X"23",X"73",X"23",X"72",X"C9",X"3A",X"2A",X"21",
		X"3C",X"32",X"2A",X"21",X"FE",X"10",X"F0",X"21",X"E8",X"20",X"87",X"87",X"F3",X"CD",X"2D",X"02");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
