library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity prom_ic40 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of prom_ic40 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7C",X"12",X"12",X"12",X"12",X"7C",X"00",
		X"00",X"34",X"4A",X"4A",X"4A",X"4A",X"7E",X"00",X"00",X"24",X"42",X"42",X"42",X"42",X"3C",X"00",
		X"00",X"3C",X"42",X"42",X"42",X"42",X"7E",X"00",X"00",X"42",X"4A",X"4A",X"4A",X"4A",X"7E",X"00",
		X"00",X"02",X"0A",X"0A",X"0A",X"0A",X"7E",X"00",X"00",X"34",X"52",X"52",X"42",X"42",X"3C",X"00",
		X"00",X"7E",X"08",X"08",X"08",X"08",X"7E",X"00",X"00",X"42",X"42",X"7E",X"42",X"42",X"00",X"00",
		X"00",X"02",X"3E",X"42",X"42",X"40",X"20",X"00",X"00",X"42",X"24",X"18",X"08",X"7E",X"00",X"00",
		X"00",X"40",X"40",X"40",X"40",X"40",X"7E",X"00",X"00",X"7E",X"04",X"08",X"08",X"04",X"7E",X"00",
		X"00",X"7E",X"20",X"10",X"08",X"04",X"7E",X"00",X"00",X"3C",X"42",X"42",X"42",X"42",X"3C",X"00",
		X"00",X"04",X"0A",X"0A",X"0A",X"0A",X"7E",X"00",X"80",X"7C",X"62",X"42",X"42",X"42",X"3C",X"00",
		X"00",X"44",X"2A",X"1A",X"0A",X"0A",X"7E",X"00",X"00",X"24",X"52",X"4A",X"4A",X"4A",X"24",X"00",
		X"00",X"02",X"02",X"7E",X"02",X"02",X"00",X"00",X"00",X"3E",X"40",X"40",X"40",X"40",X"3E",X"00",
		X"00",X"1E",X"20",X"40",X"40",X"20",X"1E",X"00",X"00",X"3E",X"40",X"3C",X"20",X"40",X"3E",X"00",
		X"00",X"42",X"24",X"18",X"18",X"24",X"42",X"00",X"00",X"02",X"04",X"78",X"04",X"02",X"00",X"00",
		X"00",X"42",X"46",X"4A",X"52",X"62",X"42",X"00",X"00",X"00",X"00",X"42",X"42",X"7E",X"00",X"00",
		X"00",X"3C",X"42",X"66",X"66",X"5A",X"3C",X"00",X"00",X"00",X"7E",X"42",X"42",X"00",X"00",X"00",
		X"00",X"08",X"04",X"7E",X"04",X"08",X"00",X"00",X"00",X"40",X"40",X"40",X"40",X"40",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",
		X"00",X"00",X"06",X"00",X"06",X"00",X"00",X"00",X"00",X"24",X"7E",X"24",X"24",X"7E",X"24",X"00",
		X"00",X"24",X"52",X"FF",X"4A",X"24",X"00",X"00",X"00",X"00",X"06",X"09",X"09",X"06",X"00",X"00",
		X"00",X"50",X"24",X"5A",X"5A",X"24",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"42",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"42",X"00",X"00",X"00",
		X"00",X"24",X"18",X"7E",X"18",X"24",X"00",X"00",X"00",X"08",X"08",X"3E",X"08",X"08",X"00",X"00",
		X"00",X"00",X"00",X"70",X"10",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"08",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"60",X"60",X"00",X"00",X"00",X"02",X"04",X"08",X"10",X"20",X"40",X"00",
		X"00",X"3C",X"46",X"4A",X"52",X"62",X"3C",X"00",X"00",X"40",X"40",X"7E",X"42",X"44",X"00",X"00",
		X"00",X"44",X"4A",X"4A",X"52",X"52",X"64",X"00",X"00",X"34",X"4A",X"4A",X"4A",X"42",X"42",X"00",
		X"00",X"10",X"7E",X"12",X"14",X"18",X"10",X"00",X"00",X"32",X"4A",X"4A",X"4A",X"4A",X"2E",X"00",
		X"00",X"30",X"4A",X"4A",X"4A",X"4A",X"3C",X"00",X"00",X"02",X"06",X"0A",X"72",X"02",X"02",X"00",
		X"00",X"34",X"4A",X"4A",X"4A",X"4A",X"34",X"00",X"00",X"3C",X"52",X"52",X"52",X"52",X"0C",X"00",
		X"00",X"00",X"00",X"24",X"24",X"00",X"00",X"00",X"00",X"00",X"00",X"64",X"24",X"00",X"00",X"00",
		X"00",X"00",X"00",X"22",X"14",X"08",X"00",X"00",X"00",X"24",X"24",X"24",X"24",X"24",X"24",X"00",
		X"00",X"00",X"08",X"14",X"22",X"00",X"00",X"00",X"00",X"04",X"0A",X"0A",X"52",X"02",X"04",X"00",
		X"40",X"40",X"50",X"58",X"5C",X"5C",X"5E",X"1E",X"00",X"C0",X"F4",X"E8",X"D4",X"AC",X"5E",X"3E",
		X"00",X"7F",X"00",X"FC",X"F8",X"F0",X"C0",X"00",X"3E",X"5E",X"AC",X"D4",X"E8",X"F4",X"C0",X"00",
		X"1E",X"5E",X"5C",X"5C",X"58",X"50",X"40",X"40",X"7C",X"7A",X"35",X"2B",X"17",X"2F",X"03",X"00",
		X"00",X"FE",X"00",X"3F",X"1F",X"0F",X"03",X"00",X"00",X"03",X"2F",X"17",X"2B",X"35",X"7A",X"7C",
		X"FE",X"FE",X"FC",X"FC",X"F8",X"F0",X"C0",X"00",X"7F",X"7F",X"3F",X"3F",X"1F",X"0F",X"03",X"00",
		X"00",X"C0",X"F0",X"F8",X"FC",X"FC",X"FE",X"FE",X"00",X"03",X"0F",X"1F",X"3F",X"3F",X"7F",X"7F",
		X"3C",X"7E",X"FE",X"FE",X"FE",X"FE",X"7E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"40",X"40",X"50",X"58",X"5C",X"5C",X"5E",X"1E",X"00",X"C0",X"F4",X"E8",X"D4",X"AC",X"5E",X"3E",
		X"00",X"7F",X"00",X"FC",X"F8",X"F0",X"C0",X"00",X"3E",X"5E",X"AC",X"D4",X"E8",X"F4",X"C0",X"00",
		X"1E",X"5E",X"5C",X"5C",X"58",X"50",X"40",X"40",X"7C",X"7A",X"35",X"2B",X"17",X"2F",X"03",X"00",
		X"00",X"FE",X"00",X"3F",X"1F",X"0F",X"03",X"00",X"00",X"03",X"2F",X"17",X"2B",X"35",X"7A",X"7C",
		X"FE",X"FE",X"FC",X"FC",X"F8",X"F0",X"C0",X"00",X"7F",X"7F",X"3F",X"3F",X"1F",X"0F",X"03",X"00",
		X"00",X"C0",X"F0",X"F8",X"FC",X"FC",X"FE",X"FE",X"00",X"03",X"0F",X"1F",X"3F",X"3F",X"7F",X"7F",
		X"00",X"24",X"18",X"7E",X"18",X"24",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3C",X"7E",X"FF",X"FF",X"FF",X"FF",X"7E",X"3C",X"3C",X"7E",X"FF",X"FF",X"FF",X"FF",X"7E",X"3C",
		X"10",X"F8",X"F0",X"38",X"10",X"F0",X"40",X"00",X"09",X"1B",X"09",X"1B",X"0D",X"0F",X"19",X"30",
		X"00",X"00",X"00",X"00",X"04",X"4C",X"E8",X"38",X"00",X"00",X"00",X"00",X"00",X"07",X"0D",X"1B",
		X"40",X"E0",X"C0",X"60",X"40",X"C0",X"00",X"00",X"26",X"6F",X"27",X"6C",X"36",X"3F",X"65",X"C0",
		X"00",X"00",X"00",X"00",X"10",X"30",X"A0",X"60",X"00",X"00",X"00",X"00",X"00",X"1D",X"37",X"6C",
		X"FE",X"64",X"C6",X"7A",X"D3",X"01",X"00",X"00",X"06",X"02",X"06",X"03",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"50",X"FC",X"64",X"C6",X"7C",X"00",X"00",X"0C",X"06",X"03",X"03",X"06",X"02",
		X"C6",X"7C",X"FE",X"4C",X"C6",X"7C",X"D6",X"03",X"06",X"02",X"06",X"02",X"06",X"03",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"50",X"FC",X"4C",X"00",X"00",X"00",X"00",X"08",X"08",X"0D",X"07",
		X"10",X"F0",X"48",X"04",X"00",X"00",X"00",X"00",X"0D",X"07",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"E0",X"90",X"10",X"F8",X"F0",X"98",X"20",X"17",X"0D",X"1B",X"09",X"1B",X"09",X"1B",
		X"4C",X"FC",X"57",X"01",X"00",X"00",X"00",X"00",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"D0",X"78",X"C4",X"4C",X"FE",X"7C",X"C6",X"0C",X"05",X"07",X"06",X"02",X"06",X"02",X"02",
		X"E0",X"C0",X"40",X"80",X"80",X"00",X"00",X"00",X"6F",X"24",X"2C",X"77",X"5D",X"C0",X"00",X"00",
		X"00",X"00",X"10",X"30",X"E0",X"C0",X"60",X"C0",X"00",X"00",X"00",X"05",X"1F",X"34",X"6C",X"27",
		X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"2C",X"77",X"DD",X"80",X"00",X"00",X"00",X"00",
		X"30",X"20",X"E0",X"40",X"60",X"C0",X"E0",X"40",X"00",X"05",X"1F",X"36",X"6C",X"27",X"6F",X"26",
		X"00",X"00",X"00",X"C0",X"00",X"00",X"08",X"04",X"00",X"02",X"00",X"02",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"20",X"10",X"00",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"10",X"01",X"08",X"00",X"0A",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"00",X"0A",
		X"80",X"10",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"08",X"00",X"00",
		X"00",X"00",X"01",X"07",X"00",X"10",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"00",X"80",X"10",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"0C",
		X"00",X"00",X"00",X"00",X"03",X"06",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"30",X"00",X"00",X"00",X"00",
		X"04",X"04",X"08",X"60",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"02",X"00",X"02",X"00",X"02",
		X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0C",X"08",X"08",X"00",X"00",X"00",X"00",
		X"01",X"0F",X"00",X"88",X"10",X"80",X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"00",X"40",X"70",X"00",X"00",X"08",X"01",X"08",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"F0",X"10",X"00",X"01",X"08",X"00",
		X"20",X"20",X"30",X"10",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"70",X"00",X"01",X"0A",X"00",X"08",X"01",
		X"00",X"00",X"00",X"C0",X"00",X"00",X"08",X"04",X"00",X"02",X"00",X"02",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"20",X"10",X"00",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"10",X"01",X"08",X"00",X"0A",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"00",X"0A",
		X"80",X"10",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"08",X"00",X"00",
		X"00",X"00",X"01",X"07",X"00",X"10",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"00",X"80",X"10",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"0C",
		X"00",X"00",X"00",X"00",X"03",X"06",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"30",X"00",X"00",X"00",X"00",
		X"04",X"04",X"08",X"60",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"02",X"00",X"02",X"00",X"02",
		X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0C",X"08",X"08",X"00",X"00",X"00",X"00",
		X"01",X"0F",X"00",X"88",X"10",X"80",X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"00",X"40",X"70",X"00",X"00",X"08",X"01",X"08",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"F0",X"10",X"00",X"01",X"08",X"00",
		X"20",X"20",X"30",X"10",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"70",X"00",X"01",X"0A",X"00",X"08",X"01",
		X"10",X"F8",X"F0",X"F8",X"10",X"F0",X"40",X"00",X"09",X"19",X"09",X"19",X"0D",X"0F",X"19",X"30",
		X"00",X"00",X"00",X"00",X"04",X"4C",X"E8",X"F8",X"00",X"00",X"00",X"00",X"00",X"07",X"0D",X"19",
		X"40",X"E0",X"C0",X"60",X"40",X"C0",X"00",X"00",X"27",X"67",X"27",X"66",X"37",X"3F",X"65",X"C0",
		X"00",X"00",X"00",X"00",X"10",X"30",X"A0",X"60",X"00",X"00",X"00",X"00",X"00",X"1D",X"37",X"66",
		X"7E",X"74",X"66",X"7A",X"D3",X"01",X"00",X"00",X"06",X"02",X"06",X"03",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"50",X"FC",X"74",X"66",X"7C",X"00",X"00",X"0C",X"06",X"03",X"03",X"06",X"02",
		X"4E",X"7C",X"7E",X"5C",X"4E",X"7C",X"D6",X"03",X"06",X"02",X"06",X"02",X"06",X"03",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"50",X"FC",X"5C",X"00",X"00",X"00",X"00",X"08",X"08",X"0D",X"07",
		X"10",X"F0",X"48",X"04",X"00",X"00",X"00",X"00",X"0D",X"07",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"E0",X"F0",X"10",X"F8",X"F0",X"F8",X"20",X"17",X"0D",X"19",X"09",X"19",X"09",X"19",
		X"5C",X"FC",X"57",X"01",X"00",X"00",X"00",X"00",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"D0",X"78",X"4C",X"5C",X"7E",X"7C",X"4E",X"0C",X"05",X"07",X"06",X"02",X"06",X"02",X"02",
		X"E0",X"C0",X"C0",X"80",X"80",X"00",X"00",X"00",X"67",X"25",X"24",X"77",X"5D",X"C0",X"00",X"00",
		X"00",X"00",X"10",X"30",X"E0",X"C0",X"E0",X"C0",X"00",X"00",X"00",X"05",X"1F",X"35",X"64",X"27",
		X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"26",X"77",X"DD",X"80",X"00",X"00",X"00",X"00",
		X"30",X"20",X"E0",X"40",X"60",X"C0",X"E0",X"40",X"00",X"05",X"1F",X"37",X"66",X"27",X"67",X"27",
		X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",
		X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",
		X"18",X"18",X"18",X"F8",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F8",X"18",X"18",X"18",
		X"18",X"18",X"18",X"1F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"1F",X"18",X"18",X"18",
		X"18",X"18",X"18",X"F8",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F8",X"18",X"18",X"18",
		X"18",X"18",X"18",X"1F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"1F",X"18",X"18",X"18",
		X"00",X"3C",X"42",X"66",X"66",X"5A",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"3C",X"42",X"42",X"42",X"42",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"81",X"BD",X"A5",X"A5",X"BD",X"81",X"FF",X"00",X"7E",X"42",X"5A",X"5A",X"42",X"7E",X"00",
		X"DB",X"ED",X"F6",X"7B",X"BD",X"DE",X"6F",X"B7",X"08",X"14",X"22",X"41",X"80",X"41",X"22",X"14");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
