`define BUILD_DATE "190421"
`define BUILD_TIME "114651"
