library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity rom_cpu3 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of rom_cpu3 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"18",X"D3",X"DC",X"01",X"B5",X"B3",X"06",X"D9",X"76",X"A8",X"61",X"D9",X"22",X"01",X"F4",X"00",
		X"7D",X"1C",X"D9",X"24",X"00",X"D9",X"05",X"01",X"D9",X"66",X"CB",X"A4",X"2B",X"3D",X"00",X"00",
		X"76",X"A9",X"60",X"D1",X"DC",X"D9",X"3E",X"EE",X"D9",X"F8",X"00",X"D9",X"F8",X"01",X"D9",X"C0",
		X"D9",X"C0",X"89",X"D7",X"B5",X"EE",X"B3",X"03",X"D9",X"FA",X"00",X"A4",X"3B",X"33",X"E2",X"1F",
		X"00",X"E2",X"C0",X"E2",X"C1",X"00",X"E2",X"C0",X"5C",X"D9",X"C0",X"D9",X"C0",X"D9",X"C0",X"D9",
		X"C0",X"89",X"E5",X"B5",X"B3",X"0C",X"D9",X"76",X"9C",X"61",X"D9",X"22",X"01",X"F4",X"00",X"7D",
		X"16",X"D9",X"24",X"00",X"D9",X"05",X"01",X"D9",X"66",X"CB",X"A4",X"2B",X"3D",X"DC",X"D9",X"3E",
		X"EE",X"D9",X"F8",X"00",X"D9",X"F8",X"01",X"D9",X"C0",X"D9",X"C0",X"89",X"DD",X"B5",X"4B",X"B4",
		X"61",X"6D",X"0F",X"9B",X"A4",X"40",X"76",X"21",X"60",X"19",X"4A",X"19",X"03",X"B3",X"04",X"76",
		X"2B",X"60",X"15",X"05",X"00",X"3D",X"1C",X"9D",X"40",X"19",X"03",X"19",X"4A",X"40",X"89",X"F5",
		X"EE",X"DE",X"B4",X"61",X"A4",X"F8",X"40",X"A4",X"B0",X"3C",X"6D",X"0F",X"7D",X"1D",X"A4",X"5C",
		X"2E",X"A4",X"CC",X"40",X"B3",X"04",X"76",X"2B",X"60",X"7A",X"C2",X"40",X"26",X"15",X"05",X"00",
		X"40",X"D3",X"19",X"FA",X"7D",X"03",X"A4",X"BA",X"42",X"89",X"F1",X"B5",X"4B",X"C3",X"61",X"72",
		X"19",X"8B",X"19",X"8B",X"19",X"8B",X"19",X"8B",X"57",X"19",X"AE",X"ED",X"10",X"19",X"80",X"ED",
		X"08",X"19",X"F6",X"7D",X"12",X"25",X"CC",X"1A",X"06",X"25",X"80",X"1A",X"02",X"25",X"33",X"76",
		X"B5",X"61",X"03",X"F8",X"EA",X"01",X"7C",X"B5",X"A4",X"26",X"1F",X"76",X"A6",X"0E",X"F4",X"33",
		X"E7",X"05",X"41",X"25",X"32",X"57",X"CE",X"00",X"40",X"69",X"76",X"D8",X"0E",X"4B",X"02",X"90",
		X"19",X"04",X"ED",X"03",X"76",X"E8",X"0E",X"4B",X"B7",X"61",X"19",X"02",X"19",X"02",X"19",X"02",
		X"19",X"02",X"6B",X"F4",X"10",X"2C",X"02",X"25",X"0F",X"57",X"40",X"22",X"DE",X"C3",X"61",X"B5",
		X"19",X"72",X"ED",X"1B",X"19",X"04",X"ED",X"2A",X"19",X"48",X"ED",X"39",X"25",X"02",X"6B",X"57",
		X"A4",X"0A",X"3C",X"22",X"F4",X"35",X"7D",X"3F",X"F4",X"37",X"7D",X"3B",X"7A",X"85",X"41",X"1D",
		X"6E",X"01",X"48",X"A4",X"0A",X"3C",X"22",X"F4",X"3D",X"7D",X"2C",X"F4",X"3F",X"7D",X"28",X"7A",
		X"85",X"41",X"6A",X"6E",X"07",X"57",X"A4",X"0A",X"3C",X"22",X"F4",X"35",X"7D",X"19",X"F4",X"37",
		X"7D",X"15",X"7A",X"85",X"41",X"25",X"08",X"EC",X"48",X"A4",X"0A",X"3C",X"22",X"F4",X"3F",X"7D",
		X"06",X"F4",X"3D",X"7D",X"02",X"0A",X"B5",X"A8",X"B5",X"19",X"72",X"ED",X"2C",X"19",X"04",X"ED",
		X"4B",X"19",X"48",X"ED",X"6A",X"25",X"02",X"6B",X"72",X"57",X"A4",X"0A",X"3C",X"22",X"F4",X"4A",
		X"9B",X"22",X"42",X"F4",X"45",X"7D",X"7B",X"65",X"5A",X"02",X"57",X"A4",X"0A",X"3C",X"22",X"F4",
		X"41",X"7D",X"6F",X"F4",X"46",X"7D",X"6B",X"1A",X"67",X"1D",X"6E",X"01",X"72",X"48",X"A4",X"0A",
		X"3C",X"22",X"F4",X"45",X"7D",X"5C",X"F4",X"46",X"7D",X"58",X"65",X"6E",X"02",X"48",X"A4",X"0A",
		X"3C",X"22",X"F4",X"4A",X"7D",X"4C",X"F4",X"41",X"7D",X"48",X"1A",X"44",X"6A",X"6E",X"81",X"72",
		X"57",X"A4",X"0A",X"3C",X"22",X"F4",X"49",X"7D",X"39",X"F4",X"43",X"7D",X"35",X"65",X"6E",X"06",
		X"57",X"A4",X"0A",X"3C",X"22",X"F4",X"41",X"7D",X"29",X"F4",X"46",X"7D",X"25",X"1A",X"21",X"25",
		X"02",X"EC",X"72",X"48",X"A4",X"0A",X"3C",X"22",X"F4",X"44",X"7D",X"16",X"F4",X"47",X"7D",X"12",
		X"65",X"5A",X"06",X"48",X"A4",X"0A",X"3C",X"22",X"F4",X"4A",X"7D",X"06",X"F4",X"41",X"7D",X"02",
		X"0A",X"B5",X"A8",X"B5",X"D9",X"22",X"00",X"F4",X"02",X"2C",X"0A",X"7D",X"0C",X"F4",X"04",X"7D",
		X"0C",X"D9",X"D1",X"02",X"B5",X"D9",X"9E",X"01",X"B5",X"D9",X"9E",X"02",X"B5",X"D9",X"D1",X"01",
		X"B5",X"D9",X"76",X"BE",X"61",X"D9",X"0D",X"00",X"D9",X"69",X"01",X"B3",X"01",X"3D",X"EA",X"0A",
		X"19",X"ED",X"19",X"5B",X"7D",X"F7",X"EE",X"7A",X"4B",X"42",X"DE",X"C8",X"61",X"CB",X"80",X"A4",
		X"11",X"39",X"DC",X"4B",X"C8",X"61",X"2C",X"E8",X"DE",X"C8",X"61",X"CB",X"65",X"D9",X"0D",X"00",
		X"D9",X"69",X"01",X"A4",X"30",X"41",X"DC",X"4B",X"C8",X"61",X"2C",X"D4",X"80",X"B5",X"32",X"1D",
		X"6D",X"0F",X"F4",X"08",X"ED",X"32",X"6A",X"6D",X"0F",X"F4",X"06",X"ED",X"2B",X"32",X"6D",X"05",
		X"ED",X"08",X"8D",X"1D",X"A4",X"7A",X"37",X"7A",X"9F",X"42",X"90",X"6A",X"A4",X"DA",X"36",X"19",
		X"4B",X"19",X"9D",X"E7",X"AA",X"42",X"C8",X"7A",X"9F",X"42",X"A4",X"03",X"37",X"7D",X"07",X"2C",
		X"07",X"19",X"30",X"7A",X"A6",X"42",X"A8",X"B5",X"0A",X"B5",X"66",X"26",X"CB",X"A4",X"F0",X"43",
		X"F7",X"03",X"00",X"76",X"BA",X"61",X"15",X"BD",X"61",X"B6",X"B2",X"EE",X"DE",X"C1",X"61",X"DE",
		X"C2",X"61",X"76",X"BD",X"61",X"22",X"C0",X"0D",X"C0",X"69",X"A4",X"7E",X"42",X"1C",X"3A",X"43",
		X"A4",X"E6",X"42",X"7A",X"BA",X"43",X"D9",X"76",X"BE",X"61",X"3E",X"DC",X"CB",X"66",X"25",X"04",
		X"49",X"04",X"B3",X"00",X"76",X"C4",X"61",X"D6",X"0D",X"A4",X"11",X"39",X"2C",X"13",X"26",X"1D",
		X"76",X"BE",X"61",X"0D",X"C0",X"69",X"A4",X"30",X"41",X"D3",X"2C",X"05",X"76",X"BD",X"61",X"91",
		X"B5",X"4B",X"C1",X"61",X"C4",X"DE",X"C1",X"61",X"76",X"BD",X"61",X"22",X"72",X"8C",X"7D",X"09",
		X"65",X"C0",X"0D",X"C0",X"69",X"A4",X"30",X"41",X"DF",X"4B",X"BD",X"61",X"72",X"4B",X"C1",X"61",
		X"B2",X"DE",X"C1",X"61",X"A4",X"41",X"42",X"7A",X"0C",X"43",X"76",X"BD",X"61",X"22",X"C0",X"0D",
		X"C0",X"69",X"A4",X"89",X"41",X"EA",X"12",X"4B",X"BD",X"61",X"72",X"19",X"02",X"19",X"02",X"19",
		X"ED",X"19",X"ED",X"B2",X"6D",X"0F",X"DE",X"BD",X"61",X"76",X"BD",X"61",X"22",X"C0",X"0D",X"C0",
		X"69",X"F4",X"02",X"7D",X"0D",X"2C",X"12",X"F4",X"04",X"7D",X"0B",X"6A",X"6E",X"04",X"57",X"7A",
		X"7B",X"43",X"38",X"7A",X"7B",X"43",X"78",X"78",X"78",X"78",X"78",X"A4",X"0A",X"3C",X"22",X"F4",
		X"63",X"F3",X"BA",X"43",X"A4",X"E5",X"3F",X"A4",X"2B",X"3D",X"66",X"76",X"01",X"60",X"19",X"F4",
		X"76",X"5F",X"60",X"19",X"11",X"3E",X"DC",X"CB",X"76",X"B4",X"61",X"25",X"04",X"49",X"7D",X"0B",
		X"F4",X"02",X"7D",X"0C",X"2C",X"0F",X"19",X"BF",X"7A",X"CE",X"43",X"19",X"5A",X"7A",X"CE",X"43",
		X"19",X"6E",X"7A",X"CE",X"43",X"19",X"54",X"7A",X"CE",X"43",X"D9",X"76",X"BD",X"61",X"A4",X"24",
		X"42",X"76",X"C2",X"61",X"D1",X"22",X"DC",X"D3",X"26",X"CB",X"4C",X"F3",X"D2",X"42",X"DC",X"D3",
		X"3E",X"66",X"26",X"CB",X"4B",X"BD",X"61",X"19",X"99",X"19",X"99",X"19",X"99",X"19",X"99",X"19",
		X"9C",X"F8",X"4B",X"BE",X"61",X"C0",X"F8",X"4B",X"BF",X"61",X"C0",X"F8",X"DC",X"D3",X"3E",X"B5",
		X"15",X"BA",X"61",X"22",X"19",X"02",X"19",X"02",X"19",X"02",X"19",X"02",X"18",X"C7",X"C0",X"22",
		X"18",X"C7",X"C0",X"22",X"18",X"B5",X"15",X"05",X"00",X"B3",X"04",X"76",X"2B",X"60",X"66",X"CB",
		X"19",X"3C",X"F3",X"E5",X"5F",X"40",X"89",X"F8",X"DC",X"3E",X"19",X"FA",X"7D",X"23",X"40",X"89",
		X"F9",X"76",X"5F",X"60",X"19",X"86",X"F9",X"D9",X"76",X"21",X"60",X"D9",X"71",X"00",X"82",X"D9",
		X"71",X"01",X"58",X"D9",X"71",X"02",X"86",X"A4",X"7F",X"1F",X"D9",X"F8",X"03",X"D9",X"A3",X"04",
		X"B5",X"66",X"CB",X"B3",X"04",X"76",X"2B",X"60",X"19",X"FA",X"7D",X"1B",X"66",X"D9",X"3E",X"25",
		X"58",X"D9",X"21",X"01",X"ED",X"11",X"25",X"86",X"D9",X"21",X"02",X"2C",X"0A",X"25",X"94",X"D9",
		X"21",X"02",X"EA",X"03",X"DC",X"3E",X"B5",X"40",X"89",X"DE",X"DC",X"65",X"6E",X"04",X"B6",X"CF",
		X"04",X"A4",X"61",X"30",X"3E",X"19",X"4A",X"19",X"5A",X"B5",X"DC",X"3E",X"B5",X"4B",X"5F",X"60",
		X"19",X"57",X"9B",X"9A",X"44",X"B6",X"27",X"D3",X"61",X"B6",X"41",X"D5",X"61",X"AB",X"62",X"4B",
		X"D7",X"61",X"F4",X"00",X"9B",X"CA",X"44",X"7A",X"42",X"45",X"A4",X"C4",X"45",X"F7",X"CF",X"62",
		X"15",X"FF",X"62",X"25",X"FF",X"D8",X"18",X"76",X"26",X"60",X"19",X"FA",X"31",X"C0",X"26",X"CB",
		X"0D",X"C0",X"69",X"25",X"35",X"4C",X"E7",X"BC",X"44",X"DC",X"D3",X"B5",X"A4",X"DC",X"45",X"DC",
		X"D3",X"9A",X"D8",X"AB",X"62",X"EB",X"22",X"FE",X"0F",X"F8",X"3F",X"F4",X"FF",X"9B",X"3C",X"45",
		X"EB",X"19",X"22",X"7D",X"12",X"66",X"26",X"15",X"F0",X"FF",X"40",X"D3",X"22",X"6D",X"0F",X"ED",
		X"05",X"19",X"54",X"38",X"92",X"18",X"3E",X"19",X"86",X"7D",X"0D",X"66",X"E1",X"22",X"6D",X"0F",
		X"ED",X"05",X"19",X"5A",X"38",X"92",X"18",X"3E",X"19",X"24",X"7D",X"12",X"66",X"26",X"15",X"10",
		X"00",X"40",X"D3",X"22",X"6D",X"0F",X"ED",X"05",X"19",X"BF",X"38",X"92",X"18",X"3E",X"19",X"05",
		X"7D",X"0D",X"66",X"A7",X"22",X"6D",X"0F",X"ED",X"05",X"19",X"6E",X"38",X"92",X"18",X"3E",X"77",
		X"66",X"76",X"01",X"90",X"19",X"22",X"3E",X"9B",X"CA",X"44",X"76",X"5F",X"60",X"19",X"BF",X"B6",
		X"8D",X"D3",X"61",X"B6",X"2F",X"D5",X"61",X"EE",X"DE",X"D7",X"61",X"B5",X"7B",X"F4",X"FF",X"9B",
		X"BE",X"45",X"7B",X"F4",X"FF",X"9B",X"B8",X"45",X"EB",X"19",X"22",X"7D",X"12",X"66",X"26",X"15",
		X"F0",X"FF",X"40",X"D3",X"22",X"6D",X"0F",X"ED",X"05",X"19",X"54",X"9A",X"92",X"D8",X"3E",X"19",
		X"86",X"7D",X"0D",X"66",X"E1",X"22",X"6D",X"0F",X"ED",X"05",X"19",X"5A",X"9A",X"92",X"D8",X"3E",
		X"19",X"24",X"7D",X"12",X"66",X"26",X"15",X"10",X"00",X"40",X"D3",X"22",X"6D",X"0F",X"ED",X"05",
		X"19",X"BF",X"9A",X"92",X"D8",X"3E",X"19",X"05",X"7D",X"0D",X"66",X"A7",X"22",X"6D",X"0F",X"ED",
		X"05",X"19",X"6E",X"9A",X"92",X"D8",X"3E",X"7C",X"66",X"76",X"01",X"90",X"19",X"22",X"3E",X"9B",
		X"42",X"45",X"76",X"5F",X"60",X"19",X"BF",X"B6",X"8D",X"D3",X"61",X"B6",X"2F",X"D5",X"61",X"19",
		X"FB",X"DE",X"D7",X"61",X"B5",X"7A",X"42",X"45",X"3F",X"F4",X"FF",X"F3",X"CA",X"44",X"76",X"5F",
		X"60",X"19",X"12",X"B5",X"15",X"10",X"00",X"76",X"00",X"62",X"66",X"B3",X"0B",X"22",X"6D",X"F0",
		X"F8",X"C0",X"89",X"F9",X"3E",X"40",X"25",X"B0",X"3A",X"ED",X"EF",X"B5",X"19",X"4B",X"19",X"4B",
		X"19",X"4B",X"19",X"4B",X"6A",X"6E",X"30",X"19",X"02",X"19",X"02",X"19",X"02",X"19",X"02",X"04",
		X"25",X"0A",X"82",X"19",X"99",X"19",X"99",X"19",X"99",X"19",X"99",X"C4",X"B5",X"D9",X"76",X"A2",
		X"0D",X"76",X"A0",X"62",X"B3",X"0B",X"15",X"F0",X"FF",X"66",X"CB",X"B3",X"05",X"D9",X"22",X"00",
		X"04",X"6D",X"0F",X"19",X"99",X"19",X"99",X"19",X"99",X"19",X"99",X"F8",X"40",X"C2",X"6D",X"F0",
		X"F8",X"40",X"D9",X"C0",X"89",X"E7",X"D9",X"22",X"00",X"19",X"99",X"19",X"99",X"19",X"99",X"19",
		X"99",X"F8",X"DC",X"3E",X"D9",X"C0",X"C0",X"89",X"D0",X"B5",X"7A",X"42",X"56",X"22",X"DE",X"C8",
		X"61",X"F4",X"36",X"AB",X"62",X"A5",X"F7",X"F0",X"FF",X"7D",X"1A",X"4B",X"C8",X"61",X"F4",X"3E",
		X"F9",X"19",X"F4",X"19",X"CD",X"0C",X"19",X"F4",X"19",X"11",X"D6",X"19",X"55",X"19",X"11",X"C0",
		X"19",X"55",X"19",X"CD",X"B5",X"19",X"6D",X"19",X"21",X"0C",X"19",X"FE",X"19",X"21",X"D6",X"19",
		X"FE",X"19",X"AA",X"C0",X"19",X"6D",X"19",X"AA",X"B5",X"FF",X"FF",X"7A",X"3D",X"46",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"A4",X"26",X"1F",X"F4",X"1E",X"2C",X"02",X"25",
		X"1E",X"76",X"88",X"47",X"DE",X"C8",X"61",X"5E",X"1E",X"EB",X"25",X"00",X"C9",X"E9",X"22",X"76",
		X"A6",X"47",X"1E",X"EB",X"25",X"00",X"C9",X"E9",X"22",X"72",X"97",X"4B",X"B8",X"61",X"04",X"65",
		X"B3",X"00",X"BA",X"2C",X"03",X"14",X"1A",X"FA",X"CB",X"C2",X"06",X"89",X"FD",X"DC",X"19",X"02",
		X"89",X"FC",X"72",X"01",X"33",X"ED",X"3C",X"4B",X"B6",X"61",X"F4",X"3B",X"ED",X"35",X"76",X"D2",
		X"61",X"22",X"D1",X"6D",X"03",X"76",X"CE",X"61",X"1E",X"EB",X"25",X"00",X"C9",X"E9",X"22",X"F4",
		X"00",X"ED",X"20",X"66",X"76",X"AE",X"47",X"4B",X"02",X"90",X"19",X"72",X"ED",X"03",X"76",X"CD",
		X"47",X"4B",X"B7",X"61",X"19",X"02",X"19",X"02",X"19",X"02",X"1E",X"EB",X"25",X"00",X"C9",X"E9",
		X"22",X"3E",X"F8",X"E2",X"76",X"C4",X"61",X"15",X"05",X"00",X"D9",X"76",X"2C",X"60",X"76",X"CE",
		X"61",X"B3",X"04",X"22",X"F4",X"00",X"7D",X"18",X"26",X"D9",X"0D",X"00",X"D9",X"69",X"01",X"A4",
		X"DC",X"45",X"57",X"CE",X"62",X"7B",X"6D",X"0F",X"D3",X"F4",X"0F",X"7D",X"03",X"E2",X"F8",X"00",
		X"E2",X"C0",X"D9",X"40",X"C0",X"89",X"DC",X"B5",X"00",X"02",X"03",X"04",X"01",X"02",X"03",X"02",
		X"03",X"04",X"03",X"04",X"05",X"05",X"06",X"06",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",
		X"07",X"07",X"07",X"07",X"07",X"07",X"05",X"05",X"05",X"04",X"03",X"02",X"01",X"01",X"03",X"03",
		X"04",X"04",X"05",X"05",X"06",X"06",X"07",X"07",X"08",X"08",X"09",X"09",X"0A",X"0A",X"0B",X"0B",
		X"0C",X"0C",X"0D",X"0D",X"0E",X"0E",X"0F",X"0F",X"10",X"10",X"11",X"11",X"12",X"0A",X"0B",X"0C",
		X"0D",X"0E",X"0F",X"10",X"11",X"12",X"13",X"14",X"15",X"16",X"17",X"18",X"19",X"1A",X"1B",X"1C",
		X"1D",X"1E",X"1F",X"20",X"21",X"22",X"23",X"24",X"25",X"26",X"27",X"28",X"F5",X"E5",X"D5",X"C5",
		X"DD",X"E5",X"06",X"0C",X"21",X"9D",X"D0",X"11",X"20",X"00",X"3E",X"FF",X"77",X"23",X"77",X"19",
		X"77",X"2B",X"77",X"19",X"10",X"F6",X"06",X"0C",X"21",X"9D",X"D4",X"3E",X"01",X"77",X"23",X"77",
		X"19",X"77",X"2B",X"77",X"19",X"10",X"F6",X"06",X"16",X"21",X"9E",X"D0",X"DD",X"21",X"08",X"49",
		X"DD",X"7E",X"00",X"77",X"19",X"DD",X"23",X"10",X"F7",X"06",X"13",X"21",X"9D",X"D0",X"DD",X"21",
		X"1E",X"49",X"DD",X"7E",X"00",X"77",X"19",X"DD",X"23",X"10",X"F7",X"DD",X"E1",X"C1",X"D1",X"E1",
		X"F1",X"C9",X"CD",X"EC",X"47",X"E5",X"D5",X"C5",X"F5",X"E5",X"D5",X"C5",X"F5",X"11",X"DE",X"D0",
		X"06",X"05",X"21",X"01",X"00",X"39",X"3E",X"00",X"ED",X"6F",X"CD",X"B2",X"48",X"ED",X"6F",X"CD",
		X"C0",X"48",X"23",X"10",X"F1",X"F1",X"C1",X"D1",X"E1",X"F1",X"C1",X"D1",X"E1",X"C5",X"D5",X"E5",
		X"DD",X"E5",X"FD",X"E5",X"C5",X"D5",X"E5",X"DD",X"E5",X"FD",X"E5",X"11",X"5D",X"D3",X"06",X"03",
		X"21",X"00",X"00",X"39",X"3E",X"00",X"ED",X"67",X"CD",X"CE",X"48",X"ED",X"67",X"CD",X"CE",X"48",
		X"23",X"ED",X"67",X"CD",X"CE",X"48",X"ED",X"67",X"CD",X"DE",X"48",X"23",X"10",X"E6",X"FD",X"E1",
		X"DD",X"E1",X"E1",X"D1",X"C1",X"FD",X"E1",X"DD",X"E1",X"E1",X"D1",X"C1",X"C9",X"76",X"CD",X"D5",
		X"22",X"C9",X"E5",X"F5",X"6B",X"62",X"77",X"11",X"20",X"00",X"19",X"5D",X"54",X"F1",X"E1",X"C9",
		X"E5",X"F5",X"6B",X"62",X"77",X"11",X"80",X"00",X"19",X"5D",X"54",X"F1",X"E1",X"C9",X"E5",X"F5",
		X"6B",X"62",X"77",X"11",X"20",X"00",X"A7",X"ED",X"52",X"5D",X"54",X"F1",X"E1",X"C9",X"E5",X"F5",
		X"6B",X"62",X"77",X"11",X"A0",X"00",X"A7",X"ED",X"52",X"5D",X"54",X"F1",X"E1",X"C9",X"21",X"00",
		X"60",X"7E",X"CD",X"42",X"48",X"DD",X"21",X"00",X"90",X"DD",X"CB",X"00",X"76",X"20",X"FA",X"DD",
		X"CB",X"00",X"76",X"28",X"FA",X"23",X"18",X"E9",X"0A",X"2A",X"FF",X"FF",X"FF",X"0C",X"2A",X"FF",
		X"FF",X"FF",X"0B",X"2A",X"FF",X"FF",X"FF",X"0E",X"2A",X"FF",X"FF",X"FF",X"0D",X"2A",X"11",X"15",
		X"2A",X"FF",X"FF",X"FF",X"FF",X"FF",X"12",X"21",X"2A",X"FF",X"FF",X"FF",X"FF",X"FF",X"12",X"22",
		X"2A",X"71",X"19",X"40",X"71",X"FF",X"40",X"7A",X"EB",X"1D",X"71",X"19",X"40",X"71",X"FF",X"40",
		X"7A",X"FE",X"1D",X"26",X"EE",X"DE",X"E0",X"61",X"7A",X"6E",X"37",X"4B",X"26",X"60",X"19",X"02",
		X"19",X"02",X"19",X"02",X"7A",X"77",X"36",X"DE",X"5F",X"60",X"DE",X"E3",X"61",X"7A",X"DC",X"02",
		X"76",X"5E",X"60",X"9E",X"9E",X"76",X"E2",X"61",X"D1",X"7A",X"E1",X"03",X"DE",X"65",X"60",X"76",
		X"E3",X"61",X"22",X"F4",X"00",X"9B",X"86",X"49",X"4B",X"5F",X"60",X"19",X"04",X"9B",X"81",X"49",
		X"9E",X"9E",X"EE",X"DE",X"E2",X"61",X"7A",X"E5",X"03",X"D9",X"76",X"2B",X"60",X"76",X"2B",X"62",
		X"15",X"05",X"00",X"B3",X"04",X"EE",X"D9",X"19",X"00",X"4E",X"ED",X"03",X"F8",X"1A",X"1F",X"21",
		X"7D",X"1C",X"D9",X"19",X"00",X"8E",X"D9",X"19",X"00",X"C6",X"97",X"D9",X"22",X"03",X"F4",X"48",
		X"7D",X"04",X"D9",X"71",X"03",X"30",X"01",X"66",X"76",X"01",X"60",X"19",X"54",X"3E",X"C0",X"D9",
		X"40",X"89",X"D3",X"25",X"00",X"DE",X"0D",X"62",X"D9",X"76",X"2B",X"60",X"76",X"2B",X"62",X"15",
		X"05",X"00",X"B3",X"04",X"66",X"26",X"CB",X"A4",X"64",X"4A",X"DC",X"D3",X"3E",X"C0",X"D9",X"40",
		X"89",X"F2",X"A4",X"C7",X"1F",X"A4",X"8F",X"17",X"A4",X"5A",X"2D",X"A4",X"01",X"4A",X"76",X"2B",
		X"62",X"B3",X"04",X"EE",X"21",X"ED",X"D1",X"C0",X"89",X"FA",X"4B",X"0E",X"62",X"5F",X"ED",X"E2",
		X"B5",X"76",X"0D",X"62",X"EE",X"21",X"31",X"19",X"3C",X"7D",X"09",X"C0",X"71",X"09",X"0C",X"19",
		X"03",X"19",X"54",X"B5",X"C0",X"22",X"5F",X"ED",X"18",X"0C",X"F8",X"76",X"00",X"D0",X"15",X"20",
		X"00",X"B3",X"04",X"CB",X"66",X"B3",X"08",X"F8",X"C0",X"89",X"FC",X"3E",X"40",X"DC",X"89",X"F3",
		X"B5",X"76",X"0D",X"62",X"4B",X"0E",X"62",X"6D",X"0F",X"72",X"B6",X"CF",X"04",X"4B",X"00",X"D0",
		X"33",X"ED",X"04",X"19",X"AC",X"1A",X"05",X"67",X"ED",X"02",X"19",X"6E",X"F4",X"00",X"ED",X"08",
		X"66",X"76",X"0E",X"62",X"9E",X"3E",X"7D",X"C3",X"19",X"0D",X"ED",X"04",X"6E",X"01",X"1A",X"BB",
		X"5A",X"01",X"1A",X"B7",X"22",X"5F",X"31",X"6D",X"0F",X"F4",X"01",X"7D",X"0D",X"F4",X"02",X"7D",
		X"28",X"F4",X"03",X"7D",X"38",X"F4",X"04",X"7D",X"58",X"B5",X"D9",X"22",X"01",X"5A",X"02",X"D9",
		X"F8",X"01",X"F4",X"B0",X"2C",X"06",X"22",X"6D",X"F0",X"FE",X"02",X"F8",X"D9",X"22",X"02",X"5A",
		X"02",X"D9",X"F8",X"02",X"F4",X"E6",X"EA",X"49",X"B5",X"D9",X"22",X"01",X"6E",X"02",X"D9",X"F8",
		X"01",X"F4",X"06",X"EA",X"E7",X"22",X"6D",X"F0",X"FE",X"01",X"F8",X"1A",X"DF",X"D9",X"22",X"01",
		X"6E",X"02",X"D9",X"F8",X"01",X"F4",X"06",X"EA",X"02",X"71",X"04",X"D9",X"22",X"02",X"6E",X"02",
		X"D9",X"F8",X"02",X"F4",X"32",X"DF",X"22",X"F4",X"04",X"25",X"02",X"ED",X"02",X"25",X"01",X"F8",
		X"B5",X"D9",X"22",X"01",X"5A",X"02",X"D9",X"F8",X"01",X"F4",X"B0",X"2C",X"DE",X"71",X"03",X"1A",
		X"DA",X"D9",X"22",X"03",X"F4",X"48",X"7D",X"1C",X"19",X"05",X"ED",X"18",X"4B",X"3C",X"62",X"5F",
		X"7D",X"0F",X"4B",X"3B",X"62",X"72",X"25",X"08",X"5A",X"10",X"89",X"FC",X"D9",X"21",X"01",X"EA",
		X"10",X"19",X"6D",X"B5",X"D9",X"22",X"02",X"F4",X"F0",X"84",X"D9",X"71",X"00",X"00",X"71",X"00",
		X"B5",X"66",X"76",X"00",X"60",X"19",X"BF",X"4B",X"3D",X"62",X"5C",X"72",X"76",X"7D",X"D0",X"15",
		X"40",X"00",X"40",X"89",X"FD",X"25",X"A4",X"15",X"20",X"00",X"A4",X"F6",X"26",X"25",X"02",X"26",
		X"15",X"00",X"04",X"40",X"D3",X"A4",X"56",X"4B",X"4B",X"3C",X"62",X"5E",X"DE",X"3C",X"62",X"4B",
		X"3D",X"62",X"5C",X"DE",X"3D",X"62",X"4B",X"0D",X"62",X"19",X"FB",X"DE",X"0D",X"62",X"3E",X"D9",
		X"71",X"00",X"00",X"71",X"00",X"B5",X"97",X"66",X"66",X"F8",X"40",X"F8",X"3E",X"0C",X"F8",X"40",
		X"F8",X"3E",X"01",X"B5",X"76",X"A6",X"D0",X"F7",X"16",X"16",X"A4",X"52",X"5D",X"76",X"22",X"60",
		X"B3",X"1E",X"71",X"00",X"C0",X"89",X"FB",X"4B",X"3D",X"62",X"5F",X"ED",X"11",X"76",X"54",X"4C",
		X"A4",X"36",X"5D",X"76",X"01",X"60",X"19",X"BF",X"A4",X"9E",X"4B",X"7A",X"37",X"4C",X"76",X"44",
		X"4C",X"A4",X"36",X"5D",X"B3",X"03",X"76",X"5C",X"62",X"71",X"00",X"C0",X"89",X"FB",X"D9",X"66",
		X"B3",X"4F",X"CB",X"A4",X"C7",X"1F",X"A4",X"8F",X"17",X"A4",X"5A",X"2D",X"DC",X"89",X"F3",X"D9",
		X"3E",X"4B",X"3D",X"62",X"5F",X"31",X"76",X"7D",X"D0",X"15",X"40",X"00",X"72",X"40",X"89",X"FD",
		X"66",X"66",X"15",X"20",X"00",X"71",X"E7",X"40",X"71",X"FF",X"3E",X"0C",X"71",X"E6",X"40",X"71",
		X"E5",X"3E",X"26",X"15",X"00",X"04",X"40",X"D3",X"25",X"02",X"A4",X"56",X"4B",X"76",X"00",X"60",
		X"19",X"F4",X"B3",X"00",X"D4",X"05",X"CE",X"00",X"D9",X"66",X"D9",X"76",X"5C",X"62",X"D9",X"22",
		X"02",X"EC",X"99",X"D9",X"F8",X"02",X"D9",X"22",X"01",X"C3",X"99",X"D9",X"F8",X"01",X"D9",X"22",
		X"00",X"56",X"99",X"D9",X"F8",X"00",X"76",X"91",X"D1",X"A4",X"06",X"1E",X"D9",X"3E",X"76",X"3D",
		X"62",X"9E",X"ED",X"8A",X"A4",X"9E",X"4B",X"76",X"01",X"60",X"19",X"54",X"76",X"5F",X"60",X"19",
		X"05",X"ED",X"14",X"D9",X"66",X"D9",X"76",X"5C",X"62",X"D9",X"3C",X"00",X"D9",X"FA",X"01",X"D9",
		X"0D",X"02",X"A4",X"72",X"3C",X"D9",X"3E",X"A4",X"9E",X"4B",X"76",X"A6",X"D0",X"F7",X"16",X"16",
		X"A4",X"52",X"5D",X"B5",X"53",X"D1",X"03",X"0C",X"0B",X"18",X"17",X"1E",X"1C",X"FF",X"19",X"18",
		X"12",X"17",X"1D",X"1C",X"93",X"D1",X"01",X"08",X"17",X"18",X"FF",X"0B",X"18",X"17",X"1E",X"1C",
		X"A4",X"91",X"4C",X"A4",X"C2",X"4C",X"A4",X"FE",X"4C",X"A4",X"DE",X"4C",X"A4",X"62",X"4D",X"1A",
		X"09",X"A4",X"91",X"4C",X"0A",X"7D",X"0B",X"A4",X"FE",X"4C",X"15",X"1C",X"60",X"A4",X"98",X"4D",
		X"1A",X"09",X"A4",X"32",X"4D",X"15",X"1C",X"60",X"A4",X"A0",X"4D",X"B3",X"01",X"A4",X"A9",X"4D",
		X"B5",X"76",X"01",X"90",X"19",X"22",X"F9",X"1A",X"F8",X"A4",X"91",X"4C",X"A4",X"D0",X"4C",X"A4",
		X"42",X"4D",X"A4",X"52",X"4D",X"B3",X"05",X"CB",X"EE",X"A4",X"87",X"4D",X"B3",X"20",X"A4",X"A9",
		X"4D",X"25",X"01",X"A4",X"87",X"4D",X"B3",X"20",X"A4",X"A9",X"4D",X"DC",X"89",X"E9",X"A4",X"FB",
		X"5B",X"B5",X"76",X"AC",X"D4",X"25",X"05",X"DE",X"6B",X"62",X"25",X"0E",X"D4",X"16",X"1A",X"1A",
		X"76",X"31",X"D5",X"25",X"0B",X"DE",X"6B",X"62",X"25",X"0E",X"D4",X"0E",X"1A",X"0C",X"76",X"82",
		X"D5",X"25",X"03",X"DE",X"6B",X"62",X"25",X"00",X"D4",X"07",X"15",X"20",X"00",X"66",X"97",X"4B",
		X"6B",X"62",X"72",X"01",X"F8",X"C0",X"89",X"FC",X"3E",X"40",X"9A",X"ED",X"F0",X"B5",X"76",X"AC",
		X"D0",X"D9",X"76",X"38",X"4E",X"25",X"05",X"DE",X"6B",X"62",X"D4",X"01",X"A4",X"70",X"4D",X"D9",
		X"76",X"CA",X"4D",X"D4",X"07",X"A4",X"70",X"4D",X"D9",X"76",X"3D",X"4E",X"D4",X"04",X"A4",X"70",
		X"4D",X"D9",X"76",X"0B",X"4E",X"D4",X"09",X"A4",X"70",X"4D",X"D9",X"76",X"38",X"4E",X"D4",X"01",
		X"1A",X"3E",X"76",X"AC",X"D0",X"D9",X"76",X"CA",X"4D",X"25",X"05",X"DE",X"6B",X"62",X"D4",X"16",
		X"1A",X"2E",X"76",X"AC",X"D0",X"25",X"05",X"DE",X"6B",X"62",X"D9",X"76",X"79",X"4E",X"D4",X"16",
		X"1A",X"1E",X"76",X"31",X"D1",X"D9",X"76",X"E7",X"4E",X"25",X"0B",X"DE",X"6B",X"62",X"D4",X"0E",
		X"1A",X"0E",X"76",X"82",X"D1",X"D9",X"76",X"DB",X"4F",X"25",X"03",X"DE",X"6B",X"62",X"D4",X"07",
		X"15",X"20",X"00",X"66",X"4B",X"6B",X"62",X"72",X"D9",X"22",X"00",X"F8",X"D9",X"C0",X"C0",X"89",
		X"F7",X"3E",X"40",X"9A",X"ED",X"ED",X"B5",X"15",X"1C",X"60",X"F7",X"2D",X"00",X"0A",X"76",X"AE",
		X"4F",X"ED",X"13",X"76",X"81",X"4F",X"1A",X"0E",X"76",X"51",X"4E",X"F7",X"14",X"00",X"1A",X"06",
		X"76",X"65",X"4E",X"F7",X"14",X"00",X"B6",X"B2",X"B5",X"4B",X"5E",X"60",X"0A",X"ED",X"0B",X"CB",
		X"A4",X"C7",X"1F",X"A4",X"8F",X"17",X"DC",X"89",X"F0",X"B5",X"F4",X"02",X"4B",X"00",X"90",X"8B",
		X"2C",X"03",X"6D",X"60",X"F9",X"6D",X"20",X"F9",X"1A",X"E5",X"00",X"00",X"58",X"57",X"00",X"56",
		X"55",X"54",X"53",X"00",X"52",X"51",X"50",X"4F",X"00",X"4E",X"4D",X"4C",X"4B",X"00",X"4A",X"49",
		X"48",X"47",X"46",X"45",X"44",X"43",X"42",X"41",X"40",X"3F",X"3E",X"3D",X"3C",X"3B",X"3A",X"39",
		X"38",X"37",X"36",X"35",X"34",X"33",X"32",X"31",X"30",X"00",X"00",X"2F",X"2E",X"00",X"00",X"00",
		X"2D",X"2C",X"2B",X"00",X"00",X"2A",X"29",X"28",X"27",X"26",X"25",X"24",X"23",X"22",X"21",X"20",
		X"1F",X"1E",X"1D",X"1C",X"1B",X"1A",X"19",X"18",X"17",X"16",X"15",X"14",X"00",X"13",X"12",X"11",
		X"10",X"0F",X"0E",X"00",X"0D",X"0C",X"0B",X"0A",X"00",X"09",X"08",X"07",X"00",X"00",X"06",X"05",
		X"04",X"03",X"00",X"00",X"00",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"6A",X"69",X"68",
		X"67",X"66",X"65",X"64",X"63",X"62",X"61",X"60",X"5F",X"00",X"00",X"5E",X"5D",X"5C",X"5B",X"5A",
		X"59",X"81",X"4C",X"74",X"78",X"03",X"11",X"5C",X"74",X"84",X"03",X"41",X"10",X"66",X"90",X"00",
		X"11",X"98",X"66",X"90",X"00",X"81",X"4C",X"74",X"60",X"03",X"11",X"5C",X"74",X"6C",X"03",X"41",
		X"08",X"66",X"90",X"00",X"11",X"A0",X"66",X"90",X"00",X"00",X"BE",X"BD",X"00",X"00",X"BC",X"BB",
		X"BA",X"00",X"00",X"B9",X"B8",X"B7",X"00",X"00",X"B6",X"B5",X"B4",X"B3",X"00",X"B2",X"B1",X"B0",
		X"AF",X"AE",X"AD",X"AC",X"AB",X"AA",X"A9",X"A8",X"A7",X"A6",X"A5",X"A4",X"A3",X"A2",X"A1",X"A0",
		X"9F",X"9E",X"9D",X"9C",X"9B",X"9A",X"00",X"99",X"98",X"97",X"90",X"96",X"95",X"94",X"90",X"90",
		X"00",X"93",X"92",X"91",X"90",X"8F",X"8E",X"00",X"00",X"8D",X"8C",X"8B",X"8A",X"00",X"89",X"88",
		X"87",X"86",X"85",X"84",X"83",X"82",X"81",X"80",X"7F",X"7E",X"7D",X"7C",X"7B",X"7A",X"79",X"78",
		X"77",X"76",X"00",X"75",X"74",X"73",X"72",X"00",X"71",X"70",X"6F",X"00",X"00",X"6E",X"6D",X"00",
		X"00",X"00",X"6C",X"6B",X"00",X"00",X"00",X"00",X"00",X"00",X"EF",X"EE",X"ED",X"EC",X"EB",X"00",
		X"00",X"00",X"00",X"EA",X"E9",X"E8",X"90",X"90",X"90",X"E7",X"E6",X"00",X"00",X"E5",X"E4",X"90",
		X"E3",X"90",X"90",X"90",X"E2",X"E1",X"E0",X"00",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",
		X"90",X"DF",X"00",X"DE",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"DD",X"DC",X"90",X"90",
		X"90",X"90",X"90",X"00",X"90",X"90",X"90",X"90",X"DB",X"90",X"90",X"90",X"90",X"90",X"00",X"90",
		X"90",X"90",X"DA",X"D9",X"90",X"90",X"90",X"90",X"90",X"00",X"90",X"90",X"90",X"D8",X"D7",X"D6",
		X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"D5",X"D4",X"90",X"90",X"90",X"90",X"90",
		X"90",X"90",X"90",X"D3",X"D2",X"D1",X"90",X"D0",X"90",X"90",X"90",X"90",X"90",X"90",X"CF",X"00",
		X"00",X"CE",X"CD",X"CC",X"CB",X"90",X"90",X"CA",X"C9",X"C8",X"00",X"00",X"00",X"C7",X"C6",X"C5",
		X"C4",X"C3",X"C2",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C1",X"C0",X"BF",X"00",X"00",X"00",
		X"00",X"81",X"44",X"9A",X"90",X"13",X"81",X"44",X"AA",X"94",X"13",X"81",X"44",X"BA",X"98",X"13",
		X"81",X"54",X"9A",X"9C",X"13",X"81",X"54",X"AA",X"A0",X"13",X"81",X"54",X"BA",X"A4",X"13",X"81",
		X"64",X"9A",X"A8",X"13",X"81",X"64",X"AA",X"AC",X"13",X"81",X"64",X"BA",X"B0",X"13",X"81",X"44",
		X"9A",X"B4",X"13",X"81",X"44",X"AA",X"B8",X"13",X"81",X"44",X"BA",X"BC",X"13",X"81",X"54",X"9A",
		X"C0",X"13",X"81",X"54",X"AA",X"C4",X"13",X"81",X"54",X"BA",X"C8",X"13",X"81",X"64",X"9A",X"CC",
		X"13",X"81",X"64",X"AA",X"D0",X"13",X"81",X"64",X"BA",X"D4",X"13",X"A9",X"FF",X"FF",X"AA",X"B6",
		X"B1",X"AB",X"B7",X"B2",X"AC",X"B8",X"B3",X"AD",X"B9",X"B4",X"AE",X"BA",X"B5",X"AF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"4B",X"02",X"90",X"6D",X"20",X"9B",X"0E",X"52",X"4B",X"65",X"60",X"0A",X"9B",X"0E",X"52",X"7A",
		X"13",X"52",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"76",X"30",X"68",X"B3",X"10",X"F8",X"C0",X"89",X"FC",X"B5",X"CB",X"A4",
		X"C7",X"1F",X"A4",X"8F",X"17",X"DC",X"89",X"F6",X"B5",X"6D",X"02",X"7D",X"0C",X"1A",X"39",X"A4",
		X"A4",X"50",X"2C",X"05",X"1A",X"42",X"A4",X"F6",X"50",X"A4",X"3E",X"25",X"A4",X"93",X"4C",X"A4",
		X"B1",X"5B",X"B5",X"A4",X"8F",X"17",X"76",X"80",X"D0",X"F7",X"18",X"20",X"A4",X"52",X"5D",X"B5",
		X"15",X"68",X"60",X"4B",X"65",X"60",X"0A",X"7D",X"03",X"15",X"6B",X"60",X"A4",X"A4",X"50",X"34",
		X"F6",X"50",X"4B",X"5F",X"60",X"7A",X"39",X"50",X"15",X"6B",X"60",X"4B",X"65",X"60",X"0A",X"7D",
		X"03",X"15",X"68",X"60",X"7A",X"3F",X"50",X"84",X"4B",X"65",X"60",X"0A",X"7D",X"02",X"25",X"FF",
		X"8B",X"DE",X"65",X"60",X"72",X"4B",X"02",X"90",X"6D",X"20",X"7D",X"04",X"65",X"DE",X"00",X"A0",
		X"7A",X"46",X"50",X"B5",X"76",X"73",X"60",X"F7",X"00",X"09",X"CB",X"26",X"66",X"A4",X"2C",X"5D",
		X"EA",X"0C",X"3E",X"F7",X"03",X"00",X"D6",X"D3",X"DC",X"77",X"89",X"EE",X"A8",X"B5",X"3E",X"D3",
		X"DC",X"D9",X"76",X"00",X"68",X"D9",X"71",X"00",X"5C",X"D9",X"71",X"01",X"20",X"D9",X"71",X"02",
		X"03",X"4B",X"02",X"90",X"6D",X"04",X"ED",X"04",X"D9",X"71",X"02",X"03",X"D9",X"71",X"03",X"00",
		X"D9",X"08",X"04",X"51",X"15",X"05",X"68",X"F7",X"03",X"00",X"B6",X"B2",X"51",X"B3",X"0A",X"71",
		X"FF",X"C0",X"89",X"FB",X"0A",X"B5",X"E2",X"76",X"12",X"68",X"E2",X"71",X"00",X"82",X"E2",X"71",
		X"01",X"58",X"E2",X"71",X"02",X"36",X"76",X"85",X"D0",X"F7",X"18",X"1A",X"A4",X"52",X"5D",X"76",
		X"4E",X"54",X"A4",X"36",X"5D",X"76",X"59",X"54",X"A4",X"36",X"5D",X"76",X"65",X"54",X"A4",X"36",
		X"5D",X"D9",X"22",X"04",X"72",X"B7",X"17",X"57",X"CE",X"00",X"76",X"6F",X"54",X"40",X"51",X"26",
		X"76",X"DE",X"D1",X"F7",X"00",X"03",X"A4",X"3F",X"5D",X"D3",X"76",X"DD",X"D0",X"F7",X"02",X"03",
		X"A4",X"3F",X"5D",X"A4",X"6D",X"5D",X"A4",X"BC",X"5D",X"F7",X"0A",X"05",X"76",X"E7",X"D0",X"15",
		X"20",X"00",X"CB",X"66",X"71",X"31",X"40",X"71",X"31",X"40",X"71",X"33",X"40",X"40",X"89",X"F4",
		X"3E",X"C0",X"C0",X"DC",X"9A",X"ED",X"EB",X"25",X"0A",X"B3",X"03",X"76",X"98",X"D1",X"A4",X"15",
		X"54",X"F7",X"04",X"05",X"76",X"16",X"D1",X"CB",X"66",X"A4",X"15",X"54",X"3E",X"0C",X"0C",X"DC",
		X"9A",X"ED",X"F4",X"B3",X"03",X"A4",X"15",X"54",X"25",X"01",X"B3",X"02",X"A4",X"15",X"54",X"B3",
		X"05",X"76",X"0C",X"D1",X"A4",X"15",X"54",X"B3",X"02",X"76",X"0A",X"D1",X"A4",X"15",X"54",X"25",
		X"27",X"B3",X"01",X"A4",X"15",X"54",X"25",X"28",X"B3",X"01",X"A4",X"15",X"54",X"25",X"24",X"B3",
		X"01",X"A4",X"15",X"54",X"25",X"2D",X"B3",X"01",X"76",X"88",X"D1",X"A4",X"15",X"54",X"25",X"29",
		X"B3",X"01",X"76",X"88",X"D2",X"A4",X"15",X"54",X"76",X"F8",X"D0",X"A4",X"28",X"54",X"76",X"F8",
		X"D2",X"A4",X"28",X"54",X"76",X"E8",X"D0",X"A4",X"28",X"54",X"A4",X"3C",X"54",X"A4",X"47",X"5E",
		X"A4",X"9C",X"5E",X"D9",X"66",X"E2",X"66",X"A4",X"C7",X"1F",X"A4",X"8F",X"17",X"E2",X"3E",X"D9",
		X"3E",X"D9",X"9E",X"01",X"ED",X"12",X"D9",X"71",X"01",X"20",X"00",X"00",X"00",X"76",X"00",X"60",
		X"19",X"6D",X"D9",X"9E",X"00",X"9B",X"29",X"53",X"7A",X"00",X"50",X"00",X"00",X"00",X"4B",X"00",
		X"90",X"1A",X"03",X"4B",X"01",X"90",X"8B",X"6D",X"0F",X"7D",X"C5",X"3D",X"2C",X"68",X"3D",X"2C",
		X"44",X"3D",X"2C",X"21",X"E2",X"71",X"00",X"82",X"E2",X"22",X"02",X"F4",X"D6",X"1C",X"E0",X"51",
		X"E2",X"FA",X"01",X"76",X"BD",X"53",X"A4",X"9F",X"53",X"1C",X"E0",X"51",X"E2",X"08",X"01",X"E2",
		X"D1",X"02",X"7A",X"E0",X"51",X"E2",X"71",X"00",X"42",X"E2",X"22",X"01",X"F4",X"A8",X"1C",X"E0",
		X"51",X"E2",X"FA",X"02",X"76",X"B1",X"53",X"A4",X"9F",X"53",X"1C",X"E0",X"51",X"E2",X"08",X"02",
		X"E2",X"D1",X"01",X"1A",X"3F",X"E2",X"71",X"00",X"22",X"E2",X"22",X"02",X"F4",X"37",X"E7",X"E0",
		X"51",X"E2",X"FA",X"01",X"76",X"BD",X"53",X"A4",X"9F",X"53",X"1C",X"E0",X"51",X"E2",X"08",X"01",
		X"E2",X"9E",X"02",X"7A",X"E0",X"51",X"E2",X"71",X"00",X"12",X"E2",X"22",X"01",X"F4",X"09",X"E7",
		X"E0",X"51",X"E2",X"FA",X"02",X"76",X"B1",X"53",X"A4",X"9F",X"53",X"1C",X"E0",X"51",X"E2",X"08",
		X"02",X"E2",X"9E",X"01",X"65",X"6E",X"02",X"E7",X"E0",X"51",X"F4",X"09",X"1C",X"E0",X"51",X"72",
		X"B7",X"B7",X"17",X"48",X"E2",X"FA",X"01",X"76",X"C4",X"53",X"A4",X"9F",X"53",X"0A",X"F3",X"E0",
		X"51",X"65",X"5E",X"EC",X"57",X"CE",X"00",X"76",X"94",X"54",X"40",X"22",X"0A",X"ED",X"07",X"76",
		X"00",X"60",X"19",X"F4",X"1A",X"53",X"F4",X"80",X"ED",X"1F",X"76",X"01",X"60",X"19",X"54",X"D9",
		X"22",X"03",X"0A",X"9B",X"E0",X"51",X"D9",X"9E",X"03",X"76",X"10",X"68",X"15",X"11",X"68",X"F7",
		X"09",X"00",X"B6",X"33",X"51",X"71",X"FF",X"1A",X"21",X"72",X"76",X"00",X"60",X"19",X"5A",X"D9",
		X"22",X"03",X"D9",X"21",X"02",X"1C",X"E0",X"51",X"D9",X"D1",X"03",X"CB",X"76",X"09",X"68",X"15",
		X"08",X"68",X"F7",X"09",X"00",X"B6",X"B2",X"51",X"DC",X"A3",X"F7",X"00",X"0A",X"15",X"08",X"68",
		X"76",X"5D",X"D1",X"A4",X"3F",X"5D",X"7A",X"E0",X"51",X"76",X"08",X"68",X"B3",X"0A",X"25",X"FF",
		X"21",X"ED",X"0E",X"C0",X"89",X"FA",X"76",X"8E",X"54",X"15",X"0C",X"68",X"F7",X"06",X"00",X"B6",
		X"B2",X"15",X"8D",X"60",X"D9",X"22",X"04",X"6E",X"08",X"EA",X"0D",X"B6",X"CF",X"72",X"B7",X"17",
		X"04",X"B3",X"00",X"76",X"8A",X"60",X"B6",X"33",X"76",X"07",X"68",X"F7",X"03",X"00",X"B6",X"33",
		X"15",X"C6",X"D3",X"D9",X"22",X"04",X"6E",X"08",X"EA",X"0F",X"B6",X"CF",X"B7",X"B7",X"B7",X"00",
		X"00",X"04",X"B3",X"00",X"76",X"BE",X"D3",X"B6",X"33",X"76",X"11",X"68",X"F7",X"06",X"00",X"B6",
		X"33",X"25",X"FF",X"18",X"9D",X"18",X"EE",X"DE",X"26",X"60",X"A4",X"C7",X"1F",X"A4",X"8F",X"17",
		X"76",X"80",X"D0",X"F7",X"18",X"20",X"A4",X"52",X"5D",X"B5",X"00",X"00",X"00",X"00",X"B5",X"3C",
		X"C0",X"22",X"82",X"EA",X"02",X"B6",X"CF",X"F4",X"07",X"2C",X"04",X"C0",X"89",X"F3",X"B5",X"FA",
		X"B5",X"0B",X"36",X"46",X"56",X"66",X"76",X"86",X"96",X"A6",X"B6",X"C6",X"D6",X"06",X"08",X"28",
		X"48",X"68",X"88",X"A8",X"05",X"1B",X"3B",X"5B",X"7B",X"9B",X"D9",X"22",X"00",X"F4",X"0C",X"2C",
		X"2C",X"F4",X"23",X"2C",X"1F",X"F4",X"3A",X"2C",X"14",X"F4",X"51",X"2C",X"09",X"6E",X"5C",X"B6",
		X"CF",X"15",X"1C",X"D6",X"1A",X"1E",X"6E",X"3A",X"15",X"65",X"D7",X"1A",X"21",X"6E",X"23",X"15",
		X"85",X"D4",X"1A",X"10",X"6E",X"22",X"B6",X"CF",X"15",X"86",X"D4",X"1A",X"11",X"6E",X"0B",X"B6",
		X"CF",X"15",X"BC",X"D4",X"EB",X"AB",X"00",X"4F",X"4F",X"4F",X"4F",X"4F",X"1A",X"03",X"EB",X"AB",
		X"00",X"40",X"71",X"05",X"B5",X"15",X"00",X"04",X"CB",X"66",X"F8",X"40",X"71",X"00",X"3E",X"F7",
		X"80",X"00",X"D6",X"DC",X"5C",X"89",X"F1",X"B5",X"F7",X"20",X"00",X"15",X"00",X"04",X"66",X"71",
		X"2B",X"40",X"71",X"01",X"3E",X"D6",X"71",X"2C",X"40",X"71",X"01",X"B5",X"25",X"57",X"DE",X"E8",
		X"D2",X"5C",X"DE",X"08",X"D3",X"25",X"02",X"DE",X"E8",X"D6",X"DE",X"08",X"D7",X"B5",X"DE",X"D0",
		X"00",X"07",X"22",X"18",X"1E",X"FF",X"10",X"0E",X"1D",X"5E",X"D2",X"00",X"08",X"11",X"12",X"FF",
		X"1C",X"0C",X"18",X"1B",X"0E",X"DD",X"D2",X"00",X"06",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1D",
		X"18",X"19",X"02",X"17",X"0D",X"03",X"1B",X"0D",X"04",X"1D",X"11",X"05",X"1D",X"11",X"06",X"1D",
		X"11",X"07",X"1D",X"11",X"08",X"1D",X"11",X"09",X"1D",X"11",X"FF",X"FF",X"FF",X"FF",X"16",X"1B",
		X"2D",X"20",X"11",X"18",X"80",X"0C",X"0B",X"0A",X"80",X"11",X"10",X"0F",X"0E",X"0D",X"16",X"15",
		X"14",X"13",X"12",X"1B",X"1A",X"19",X"18",X"17",X"20",X"1F",X"1E",X"1D",X"1C",X"02",X"01",X"23",
		X"22",X"21",X"07",X"06",X"05",X"04",X"03",X"24",X"28",X"27",X"09",X"08",X"00",X"29",X"FF",X"2D",
		X"80",X"97",X"CB",X"26",X"66",X"76",X"0B",X"62",X"71",X"00",X"C0",X"71",X"00",X"C0",X"71",X"00",
		X"C0",X"71",X"00",X"76",X"D1",X"57",X"3C",X"C0",X"22",X"CB",X"66",X"A4",X"00",X"55",X"3E",X"DC",
		X"23",X"ED",X"F4",X"76",X"D1",X"57",X"3C",X"A4",X"22",X"55",X"04",X"C0",X"22",X"CB",X"26",X"66",
		X"76",X"F9",X"D4",X"A4",X"23",X"56",X"08",X"3E",X"D3",X"DC",X"23",X"ED",X"EA",X"7A",X"A1",X"55",
		X"97",X"66",X"76",X"1F",X"62",X"B6",X"57",X"03",X"F8",X"76",X"2F",X"62",X"19",X"72",X"7D",X"03",
		X"22",X"8B",X"F8",X"22",X"19",X"72",X"7D",X"05",X"3E",X"01",X"7A",X"52",X"55",X"3E",X"01",X"7A",
		X"78",X"55",X"CB",X"B6",X"57",X"3D",X"1E",X"3D",X"6D",X"03",X"7D",X"F7",X"72",X"4B",X"1F",X"62",
		X"17",X"DE",X"1F",X"62",X"6D",X"03",X"F4",X"03",X"ED",X"04",X"25",X"03",X"1A",X"12",X"F4",X"02",
		X"ED",X"04",X"25",X"02",X"1A",X"0A",X"F4",X"01",X"ED",X"04",X"25",X"01",X"1A",X"02",X"25",X"00",
		X"DC",X"B5",X"76",X"FB",X"D0",X"A4",X"23",X"56",X"00",X"00",X"00",X"22",X"00",X"F4",X"33",X"ED",
		X"04",X"25",X"3B",X"1A",X"02",X"25",X"3C",X"F8",X"0C",X"71",X"3D",X"0C",X"71",X"3E",X"0C",X"71",
		X"3F",X"15",X"E1",X"FF",X"40",X"71",X"40",X"B5",X"76",X"B9",X"D0",X"A4",X"23",X"56",X"00",X"00",
		X"00",X"00",X"00",X"22",X"00",X"F4",X"33",X"ED",X"04",X"25",X"34",X"1A",X"02",X"25",X"38",X"F8",
		X"15",X"20",X"00",X"40",X"71",X"35",X"40",X"71",X"36",X"C0",X"71",X"39",X"0C",X"40",X"71",X"37",
		X"B5",X"76",X"D1",X"57",X"A4",X"D2",X"55",X"B6",X"57",X"72",X"45",X"A2",X"61",X"A4",X"C1",X"55",
		X"45",X"A4",X"61",X"A4",X"C1",X"55",X"45",X"A6",X"61",X"A4",X"C1",X"55",X"3E",X"D3",X"DC",X"01",
		X"B5",X"25",X"03",X"15",X"00",X"04",X"40",X"F8",X"C0",X"F8",X"15",X"E0",X"FF",X"40",X"F8",X"0C",
		X"F8",X"B5",X"3C",X"C0",X"22",X"97",X"CB",X"66",X"76",X"F9",X"D0",X"A4",X"23",X"56",X"22",X"F4",
		X"36",X"7D",X"06",X"F4",X"3E",X"7D",X"1D",X"1A",X"33",X"15",X"00",X"04",X"40",X"15",X"E0",X"FF",
		X"3C",X"C0",X"A3",X"C0",X"A3",X"0C",X"0C",X"40",X"A3",X"40",X"A3",X"15",X"20",X"00",X"40",X"40",
		X"40",X"A3",X"1A",X"18",X"15",X"00",X"04",X"40",X"15",X"C0",X"FF",X"3C",X"40",X"A3",X"15",X"20",
		X"00",X"40",X"A3",X"40",X"C0",X"A3",X"C0",X"A3",X"0C",X"0C",X"0C",X"A3",X"3E",X"DC",X"01",X"23",
		X"ED",X"B1",X"B5",X"72",X"3D",X"3D",X"3D",X"3D",X"6D",X"0F",X"F4",X"01",X"7D",X"05",X"0C",X"0C",
		X"5E",X"1A",X"F7",X"15",X"40",X"00",X"65",X"6D",X"0F",X"F4",X"01",X"7D",X"04",X"40",X"5E",X"1A",
		X"F8",X"B5",X"97",X"B3",X"0A",X"D4",X"0A",X"65",X"06",X"06",X"06",X"06",X"C8",X"CB",X"97",X"76",
		X"F9",X"D0",X"A4",X"23",X"56",X"01",X"72",X"22",X"76",X"00",X"62",X"A5",X"F7",X"F0",X"FF",X"F4",
		X"36",X"7D",X"0D",X"F4",X"3E",X"7D",X"16",X"DC",X"9A",X"ED",X"DC",X"23",X"ED",X"D7",X"01",X"B5",
		X"19",X"21",X"0C",X"19",X"21",X"D6",X"19",X"AA",X"C0",X"19",X"AA",X"1A",X"EA",X"19",X"CD",X"0C",
		X"19",X"11",X"D6",X"19",X"11",X"C0",X"19",X"CD",X"1A",X"DD",X"97",X"66",X"19",X"7C",X"19",X"38",
		X"25",X"0F",X"E5",X"8B",X"5A",X"0E",X"72",X"19",X"7C",X"19",X"38",X"25",X"F0",X"E5",X"6E",X"20",
		X"B2",X"06",X"06",X"06",X"06",X"72",X"3E",X"01",X"B5",X"C2",X"F4",X"00",X"7D",X"0D",X"65",X"6D",
		X"0F",X"F4",X"01",X"ED",X"03",X"25",X"01",X"B5",X"25",X"03",X"B5",X"65",X"3D",X"3D",X"3D",X"3D",
		X"6D",X"0F",X"F4",X"01",X"ED",X"03",X"25",X"01",X"B5",X"25",X"03",X"B5",X"97",X"CB",X"26",X"66",
		X"76",X"D1",X"57",X"A4",X"DB",X"56",X"3E",X"D3",X"DC",X"01",X"B5",X"3C",X"C0",X"22",X"97",X"CB",
		X"66",X"76",X"F9",X"D0",X"A4",X"23",X"56",X"22",X"F4",X"36",X"7D",X"06",X"F4",X"3E",X"7D",X"32",
		X"1A",X"29",X"15",X"C0",X"03",X"40",X"22",X"6D",X"0F",X"72",X"15",X"40",X"00",X"40",X"22",X"6D",
		X"0F",X"33",X"7D",X"17",X"A4",X"48",X"57",X"15",X"20",X"00",X"40",X"A3",X"15",X"E0",X"FF",X"40",
		X"A3",X"C0",X"A3",X"C0",X"A3",X"0C",X"0C",X"40",X"A3",X"40",X"A3",X"3E",X"DC",X"01",X"23",X"ED",
		X"BB",X"B5",X"15",X"02",X"04",X"40",X"22",X"6D",X"0F",X"72",X"0C",X"0C",X"22",X"6D",X"0F",X"33",
		X"7D",X"E9",X"A4",X"48",X"57",X"15",X"E0",X"FF",X"0C",X"A3",X"C0",X"A3",X"C0",X"A3",X"C0",X"A3",
		X"0C",X"0C",X"40",X"A3",X"40",X"A3",X"1A",X"D3",X"25",X"AA",X"DE",X"0F",X"62",X"66",X"26",X"CB",
		X"97",X"F2",X"00",X"A4",X"2C",X"3C",X"01",X"DC",X"D3",X"3E",X"A4",X"26",X"1F",X"F4",X"02",X"EA",
		X"03",X"B3",X"03",X"B5",X"65",X"F4",X"00",X"ED",X"03",X"B3",X"01",X"B5",X"F4",X"01",X"ED",X"03",
		X"B3",X"03",X"B5",X"F4",X"02",X"ED",X"03",X"B3",X"03",X"B5",X"F4",X"03",X"ED",X"03",X"B3",X"00",
		X"B5",X"B3",X"02",X"B5",X"66",X"26",X"CB",X"97",X"76",X"D1",X"57",X"C0",X"22",X"76",X"F9",X"D4",
		X"A4",X"23",X"56",X"22",X"6D",X"0F",X"72",X"D4",X"00",X"CB",X"76",X"D1",X"57",X"A4",X"B3",X"57",
		X"DC",X"C2",X"F4",X"00",X"ED",X"07",X"01",X"DC",X"D3",X"3E",X"A8",X"02",X"B5",X"01",X"DC",X"D3",
		X"3E",X"A8",X"B5",X"3C",X"C0",X"22",X"66",X"CB",X"76",X"F9",X"D4",X"A4",X"23",X"56",X"22",X"DC",
		X"3E",X"D9",X"3E",X"D3",X"6D",X"0F",X"DD",X"7D",X"01",X"7C",X"26",X"D9",X"66",X"23",X"ED",X"E4",
		X"B5",X"1F",X"11",X"41",X"71",X"A1",X"22",X"52",X"33",X"63",X"93",X"14",X"44",X"74",X"A4",X"25",
		X"85",X"36",X"66",X"96",X"17",X"47",X"77",X"A7",X"28",X"58",X"88",X"69",X"99",X"1A",X"4A",X"7A",
		X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"66",X"26",X"CB",X"97",X"DE",X"3F",X"62",X"76",X"2B",X"60",X"B3",X"04",X"22",
		X"B6",X"8D",X"AE",X"62",X"6D",X"03",X"F4",X"00",X"ED",X"0D",X"C0",X"C0",X"C0",X"C0",X"C0",X"7A",
		X"44",X"58",X"00",X"00",X"00",X"00",X"00",X"19",X"22",X"7D",X"04",X"19",X"21",X"19",X"55",X"C0",
		X"22",X"5A",X"00",X"6D",X"F0",X"5A",X"08",X"F8",X"C0",X"22",X"5A",X"02",X"6D",X"F0",X"5A",X"06",
		X"F8",X"A4",X"94",X"58",X"23",X"ED",X"C8",X"76",X"01",X"90",X"19",X"22",X"ED",X"FC",X"19",X"22",
		X"7D",X"FC",X"A4",X"C7",X"1F",X"CE",X"08",X"26",X"A4",X"C7",X"1F",X"A4",X"8F",X"17",X"A4",X"C7",
		X"1F",X"A4",X"8F",X"17",X"A4",X"C7",X"1F",X"A4",X"8F",X"17",X"76",X"D1",X"57",X"FA",X"C0",X"66",
		X"3C",X"65",X"76",X"F9",X"D4",X"CB",X"A4",X"23",X"56",X"22",X"6D",X"0F",X"72",X"4B",X"3F",X"62",
		X"33",X"ED",X"03",X"A4",X"40",X"59",X"DC",X"3E",X"9A",X"ED",X"E3",X"D3",X"2A",X"ED",X"C8",X"01",
		X"DC",X"D3",X"3E",X"B5",X"66",X"26",X"CB",X"97",X"69",X"0C",X"0D",X"1D",X"19",X"02",X"19",X"02",
		X"19",X"02",X"19",X"02",X"6D",X"0F",X"5A",X"01",X"48",X"6A",X"8B",X"5A",X"F0",X"6D",X"F0",X"EC",
		X"48",X"76",X"F9",X"D0",X"A4",X"23",X"56",X"22",X"F4",X"36",X"ED",X"03",X"A4",X"03",X"59",X"F4",
		X"3E",X"ED",X"03",X"A4",X"03",X"59",X"C0",X"C0",X"22",X"F4",X"36",X"ED",X"03",X"A4",X"09",X"59",
		X"F4",X"3E",X"ED",X"03",X"A4",X"09",X"59",X"15",X"C0",X"FF",X"40",X"22",X"F4",X"36",X"ED",X"03",
		X"A4",X"0F",X"59",X"F4",X"3E",X"ED",X"03",X"A4",X"0F",X"59",X"0C",X"0C",X"22",X"F4",X"36",X"ED",
		X"03",X"A4",X"15",X"59",X"F4",X"3E",X"ED",X"03",X"A4",X"15",X"59",X"01",X"DC",X"D3",X"3E",X"C0",
		X"C0",X"C0",X"B5",X"66",X"CB",X"D4",X"03",X"1A",X"10",X"66",X"CB",X"D4",X"04",X"1A",X"0A",X"66",
		X"CB",X"D4",X"01",X"1A",X"04",X"66",X"CB",X"D4",X"02",X"15",X"00",X"04",X"40",X"22",X"6D",X"0F",
		X"72",X"4B",X"3F",X"62",X"33",X"ED",X"16",X"C2",X"B6",X"27",X"AE",X"62",X"76",X"2F",X"62",X"15",
		X"FF",X"FF",X"04",X"65",X"F4",X"00",X"7D",X"04",X"40",X"5E",X"ED",X"FC",X"08",X"DC",X"3E",X"B5",
		X"4B",X"3F",X"62",X"48",X"F7",X"00",X"FC",X"D6",X"22",X"F4",X"36",X"ED",X"03",X"7A",X"88",X"59",
		X"F4",X"48",X"ED",X"03",X"7A",X"C0",X"59",X"F4",X"3E",X"ED",X"03",X"7A",X"14",X"5A",X"7A",X"56",
		X"5A",X"F7",X"C0",X"FF",X"F2",X"FF",X"66",X"D6",X"07",X"F7",X"1F",X"00",X"D6",X"07",X"C0",X"07",
		X"C0",X"07",X"F7",X"1E",X"00",X"D6",X"07",X"C0",X"07",X"C0",X"07",X"C0",X"07",X"F7",X"1D",X"00",
		X"D6",X"07",X"C0",X"07",X"C0",X"07",X"3E",X"B5",X"A4",X"61",X"59",X"71",X"48",X"F7",X"00",X"04",
		X"66",X"D6",X"91",X"3E",X"66",X"C0",X"71",X"47",X"D6",X"91",X"3E",X"66",X"CB",X"F7",X"21",X"00",
		X"D6",X"71",X"46",X"DC",X"D6",X"91",X"3E",X"66",X"CB",X"F7",X"E0",X"FF",X"D6",X"DC",X"71",X"49",
		X"D6",X"91",X"3E",X"66",X"CB",X"F7",X"DF",X"FF",X"D6",X"71",X"4A",X"DC",X"D6",X"91",X"3E",X"B5",
		X"A4",X"61",X"59",X"F7",X"00",X"04",X"66",X"71",X"3E",X"D6",X"91",X"3E",X"66",X"C0",X"71",X"3D",
		X"D6",X"91",X"3E",X"66",X"C0",X"C0",X"92",X"6D",X"1F",X"F4",X"1A",X"2C",X"04",X"71",X"3C",X"1A",
		X"02",X"71",X"3B",X"D6",X"91",X"3E",X"66",X"0C",X"71",X"3F",X"D6",X"91",X"3E",X"66",X"CB",X"F7",
		X"E0",X"FF",X"D6",X"DC",X"71",X"40",X"D6",X"91",X"3E",X"E0",X"F4",X"D0",X"ED",X"08",X"92",X"6D",
		X"E0",X"F4",X"E0",X"ED",X"01",X"B5",X"66",X"CB",X"F7",X"C0",X"FF",X"D6",X"71",X"33",X"DC",X"D6",
		X"71",X"00",X"3E",X"B5",X"A4",X"61",X"59",X"F7",X"00",X"04",X"66",X"71",X"42",X"D6",X"91",X"3E",
		X"66",X"0C",X"71",X"44",X"D6",X"91",X"3E",X"66",X"CB",X"F7",X"E0",X"FF",X"D6",X"DC",X"71",X"40",
		X"D6",X"91",X"3E",X"66",X"CB",X"F7",X"E1",X"FF",X"D6",X"DC",X"71",X"41",X"D6",X"91",X"3E",X"66",
		X"CB",X"F7",X"20",X"00",X"D6",X"DC",X"71",X"43",X"D6",X"91",X"3E",X"66",X"CB",X"F7",X"1F",X"00",
		X"D6",X"DC",X"D6",X"91",X"3E",X"B5",X"A4",X"61",X"59",X"F7",X"00",X"04",X"66",X"71",X"36",X"D6",
		X"91",X"3E",X"66",X"C0",X"71",X"39",X"D6",X"91",X"3E",X"66",X"CB",X"F7",X"20",X"00",X"D6",X"DC",
		X"71",X"37",X"D6",X"91",X"3E",X"66",X"CB",X"F7",X"E0",X"FF",X"D6",X"DC",X"71",X"35",X"D6",X"91",
		X"3E",X"66",X"CB",X"F7",X"C0",X"FF",X"D6",X"DC",X"E0",X"F4",X"D0",X"ED",X"0B",X"92",X"6D",X"E0",
		X"F4",X"A0",X"ED",X"04",X"71",X"38",X"1A",X"02",X"71",X"34",X"D6",X"91",X"3E",X"92",X"6D",X"1F",
		X"F4",X"19",X"EA",X"09",X"66",X"C0",X"C0",X"71",X"33",X"D6",X"71",X"00",X"3E",X"B5",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"EE",X"DE",X"65",X"60",X"76",X"0F",X"5C",X"15",X"1C",X"60",X"F7",X"32",X"00",X"00",
		X"00",X"76",X"56",X"5C",X"A4",X"36",X"5D",X"4B",X"03",X"90",X"6D",X"0F",X"97",X"76",X"27",X"D1",
		X"A4",X"41",X"5C",X"01",X"72",X"25",X"06",X"DE",X"27",X"D5",X"DE",X"27",X"D6",X"4B",X"03",X"90",
		X"6D",X"F0",X"BC",X"BC",X"BC",X"BC",X"33",X"31",X"76",X"25",X"D1",X"A4",X"41",X"5C",X"25",X"06",
		X"DE",X"25",X"D5",X"DE",X"25",X"D6",X"76",X"1B",X"5D",X"A4",X"36",X"5D",X"51",X"A4",X"36",X"5D",
		X"B5",X"97",X"CB",X"B3",X"1F",X"A4",X"2E",X"50",X"DC",X"01",X"B5",X"76",X"1C",X"60",X"71",X"00",
		X"15",X"1D",X"60",X"F7",X"31",X"00",X"B6",X"B2",X"A4",X"C7",X"1F",X"7A",X"53",X"50",X"B5",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"66",X"B7",X"57",X"CE",X"00",X"76",X"65",X"5C",X"40",X"69",X"C0",X"0D",X"3E",X"B3",X"0F",
		X"D4",X"02",X"A4",X"3F",X"5D",X"B5",X"69",X"D1",X"00",X"0B",X"12",X"17",X"1C",X"0E",X"1B",X"1D",
		X"FF",X"0C",X"18",X"12",X"17",X"85",X"5C",X"85",X"5C",X"85",X"5C",X"85",X"5C",X"85",X"5C",X"85",
		X"5C",X"0C",X"5D",X"FD",X"5C",X"EE",X"5C",X"DF",X"5C",X"D0",X"5C",X"C1",X"5C",X"B2",X"5C",X"A3",
		X"5C",X"94",X"5C",X"85",X"5C",X"01",X"FF",X"0C",X"18",X"12",X"17",X"FF",X"FF",X"01",X"FF",X"19",
		X"15",X"0A",X"22",X"FF",X"01",X"FF",X"0C",X"18",X"12",X"17",X"FF",X"FF",X"02",X"FF",X"19",X"15",
		X"0A",X"22",X"1C",X"01",X"FF",X"0C",X"18",X"12",X"17",X"FF",X"FF",X"03",X"FF",X"19",X"15",X"0A",
		X"22",X"1C",X"01",X"FF",X"0C",X"18",X"12",X"17",X"FF",X"FF",X"04",X"FF",X"19",X"15",X"0A",X"22",
		X"1C",X"01",X"FF",X"0C",X"18",X"12",X"17",X"FF",X"FF",X"05",X"FF",X"19",X"15",X"0A",X"22",X"1C",
		X"02",X"FF",X"0C",X"18",X"12",X"17",X"1C",X"FF",X"01",X"FF",X"19",X"15",X"0A",X"22",X"FF",X"02",
		X"FF",X"0C",X"18",X"12",X"17",X"1C",X"FF",X"03",X"FF",X"19",X"15",X"0A",X"22",X"1C",X"03",X"FF",
		X"0C",X"18",X"12",X"17",X"1C",X"FF",X"01",X"FF",X"19",X"15",X"0A",X"22",X"FF",X"03",X"FF",X"0C",
		X"18",X"12",X"17",X"1C",X"FF",X"02",X"FF",X"19",X"15",X"0A",X"22",X"1C",X"04",X"FF",X"0C",X"18",
		X"12",X"17",X"1C",X"FF",X"01",X"FF",X"19",X"15",X"0A",X"22",X"FF",X"E8",X"D0",X"01",X"05",X"1B",
		X"12",X"10",X"11",X"1D",X"E6",X"D0",X"01",X"04",X"15",X"0E",X"0F",X"1D",X"B3",X"03",X"7B",X"21",
		X"F9",X"C7",X"C0",X"89",X"F9",X"B5",X"69",X"C0",X"0D",X"C0",X"FA",X"C0",X"3C",X"C0",X"51",X"26",
		X"66",X"7B",X"F8",X"15",X"00",X"04",X"40",X"08",X"3E",X"15",X"20",X"00",X"40",X"D3",X"C7",X"89",
		X"EE",X"B5",X"26",X"15",X"00",X"04",X"CB",X"66",X"66",X"71",X"FF",X"40",X"71",X"00",X"3E",X"C0",
		X"89",X"F6",X"3E",X"F7",X"20",X"00",X"D6",X"DC",X"9A",X"ED",X"EB",X"D3",X"B5",X"15",X"BD",X"D2",
		X"76",X"05",X"68",X"EE",X"B3",X"06",X"B6",X"EB",X"7D",X"09",X"FE",X"80",X"97",X"6D",X"0F",X"5A",
		X"00",X"18",X"01",X"66",X"76",X"20",X"00",X"40",X"51",X"3E",X"19",X"81",X"7D",X"05",X"B6",X"EB",
		X"C0",X"1A",X"06",X"19",X"AE",X"ED",X"02",X"FE",X"80",X"89",X"DB",X"B5",X"F7",X"18",X"18",X"76",
		X"85",X"D0",X"A4",X"52",X"5D",X"76",X"1C",X"60",X"15",X"05",X"00",X"71",X"00",X"40",X"71",X"00",
		X"40",X"B3",X"07",X"40",X"71",X"00",X"89",X"FB",X"A4",X"BC",X"5D",X"B5",X"7A",X"EB",X"5D",X"91",
		X"C0",X"07",X"C0",X"66",X"26",X"15",X"FE",X"03",X"40",X"F8",X"C0",X"F8",X"D3",X"3E",X"89",X"EF",
		X"B5",X"91",X"CB",X"F7",X"20",X"00",X"D6",X"07",X"D6",X"DC",X"66",X"26",X"15",X"C0",X"03",X"40",
		X"F8",X"15",X"20",X"00",X"40",X"F8",X"D3",X"3E",X"89",X"E7",X"B5",X"15",X"E5",X"E5",X"25",X"02",
		X"B3",X"0B",X"76",X"BC",X"D0",X"A4",X"D1",X"5D",X"15",X"52",X"52",X"25",X"02",X"B3",X"0C",X"76",
		X"85",X"D0",X"A4",X"D1",X"5D",X"15",X"4C",X"4C",X"25",X"02",X"B3",X"0C",X"76",X"86",X"D0",X"A4",
		X"BF",X"5D",X"15",X"50",X"50",X"B3",X"0C",X"76",X"66",X"D3",X"A4",X"BF",X"5D",X"15",X"54",X"54",
		X"76",X"9E",X"D0",X"25",X"02",X"B3",X"0C",X"A4",X"D1",X"5D",X"25",X"4D",X"DE",X"85",X"D0",X"25",
		X"51",X"DE",X"65",X"D3",X"25",X"4B",X"DE",X"9E",X"D0",X"25",X"4E",X"76",X"7E",X"D3",X"F8",X"25",
		X"4F",X"0C",X"F8",X"0C",X"F8",X"B5",X"FF",X"D9",X"66",X"E2",X"66",X"A4",X"D1",X"1D",X"A4",X"8B",
		X"1E",X"B3",X"06",X"25",X"05",X"76",X"A1",X"D5",X"A4",X"7D",X"1E",X"A4",X"E0",X"1E",X"A4",X"26",
		X"28",X"B3",X"05",X"25",X"01",X"76",X"E1",X"D4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"D9",X"76",X"1C",X"60",X"D9",X"71",X"00",X"82",X"D9",X"71",X"01",X"08",
		X"D9",X"71",X"02",X"0F",X"A4",X"7F",X"1F",X"D9",X"F8",X"03",X"D9",X"A3",X"04",X"A4",X"C7",X"1F",
		X"A4",X"8F",X"17",X"D9",X"71",X"00",X"81",X"E2",X"3E",X"D9",X"3E",X"B5",X"15",X"26",X"60",X"76",
		X"12",X"68",X"F7",X"03",X"00",X"B6",X"B2",X"51",X"71",X"00",X"C0",X"71",X"00",X"B5",X"15",X"3F",
		X"60",X"1A",X"EC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"40",X"71",X"0D",
		X"40",X"7A",X"FA",X"1E",X"71",X"1C",X"40",X"71",X"0C",X"40",X"71",X"18",X"40",X"71",X"1B",X"40",
		X"71",X"0E",X"40",X"04",X"B3",X"01",X"B5",X"A4",X"0D",X"30",X"A4",X"41",X"5F",X"A4",X"06",X"44",
		X"B5",X"76",X"0C",X"62",X"19",X"0D",X"31",X"D9",X"66",X"76",X"01",X"60",X"19",X"5A",X"B3",X"48",
		X"CB",X"A4",X"C7",X"1F",X"A4",X"8F",X"17",X"A4",X"5A",X"2D",X"A4",X"6C",X"5F",X"DC",X"89",X"F0",
		X"EE",X"DE",X"49",X"60",X"76",X"26",X"60",X"19",X"54",X"D9",X"3E",X"B5",X"3E",X"DC",X"CB",X"66",
		X"65",X"F4",X"01",X"ED",X"2C",X"76",X"0C",X"62",X"71",X"00",X"0C",X"22",X"DE",X"C3",X"61",X"D9",
		X"76",X"2B",X"60",X"15",X"05",X"00",X"B3",X"04",X"D9",X"19",X"00",X"4E",X"7D",X"0E",X"D9",X"19",
		X"04",X"66",X"7D",X"08",X"D9",X"19",X"00",X"86",X"D9",X"19",X"00",X"8E",X"D9",X"40",X"89",X"E8",
		X"B5",X"BC",X"84",X"BC",X"84",X"BC",X"84",X"6D",X"0F",X"31",X"72",X"25",X"68",X"5A",X"04",X"89",
		X"FC",X"D4",X"1C",X"D9",X"66",X"D9",X"76",X"2B",X"60",X"15",X"05",X"00",X"B3",X"04",X"D9",X"19",
		X"00",X"4E",X"7D",X"18",X"97",X"25",X"48",X"D9",X"21",X"03",X"7D",X"06",X"D9",X"19",X"04",X"66",
		X"7D",X"09",X"01",X"D9",X"F8",X"03",X"D9",X"08",X"04",X"1A",X"01",X"01",X"D9",X"40",X"89",X"DE",
		X"D9",X"3E",X"B5",X"FF",X"FF",X"EE",X"DE",X"21",X"60",X"7A",X"7A",X"44",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
