library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity Qbert_snd2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of Qbert_snd2 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"4C",X"CC",X"77",X"60",X"95",X"00",X"9E",X"00",X"A7",X"00",X"B1",X"00",X"BC",X"00",X"C7",X"00",
		X"D3",X"00",X"DF",X"00",X"ED",X"00",X"FB",X"00",X"0B",X"01",X"1A",X"01",X"2B",X"01",X"44",X"24",
		X"44",X"23",X"24",X"14",X"24",X"64",X"44",X"64",X"42",X"34",X"44",X"74",X"44",X"74",X"B3",X"B3",
		X"00",X"A5",X"20",X"38",X"E9",X"01",X"0A",X"0A",X"A8",X"A2",X"00",X"B9",X"8A",X"78",X"95",X"00",
		X"C8",X"E8",X"E0",X"04",X"D0",X"F5",X"A9",X"00",X"85",X"06",X"85",X"04",X"85",X"05",X"A9",X"FF",
		X"85",X"07",X"18",X"A5",X"06",X"65",X"02",X"85",X"06",X"A5",X"00",X"69",X"00",X"85",X"00",X"A5",
		X"03",X"69",X"00",X"85",X"03",X"A5",X"00",X"C5",X"01",X"B0",X"1C",X"18",X"A5",X"04",X"65",X"00",
		X"85",X"04",X"A5",X"05",X"65",X"03",X"85",X"05",X"29",X"0F",X"A8",X"B9",X"88",X"71",X"25",X"07",
		X"4A",X"8D",X"00",X"90",X"4C",X"52",X"78",X"4C",X"35",X"70",X"0A",X"60",X"0F",X"00",X"3F",X"7F",
		X"10",X"00",X"7F",X"C0",X"0E",X"00",X"C0",X"FF",X"0C",X"00",X"00",X"7F",X"17",X"01",X"7F",X"FF",
		X"1C",X"01",X"00",X"D0",X"37",X"02",X"00",X"FF",X"4F",X"03",X"A9",X"41",X"85",X"00",X"85",X"01",
		X"A9",X"78",X"85",X"2B",X"A9",X"F0",X"85",X"2A",X"A9",X"FF",X"8D",X"00",X"B0",X"A0",X"00",X"84",
		X"29",X"B1",X"2A",X"49",X"FF",X"8D",X"00",X"A0",X"38",X"A5",X"00",X"E9",X"02",X"85",X"00",X"A5",
		X"01",X"E9",X"00",X"85",X"01",X"B0",X"F1",X"E6",X"2A",X"D0",X"02",X"E6",X"2B",X"A9",X"CD",X"8D",
		X"00",X"B0",X"A0",X"00",X"84",X"29",X"B1",X"2A",X"49",X"FF",X"8D",X"00",X"A0",X"4C",X"35",X"70",
		X"0E",X"15",X"09",X"22",X"3F",X"0E",X"15",X"02",X"29",X"3F",X"A9",X"3F",X"49",X"FF",X"8D",X"00",
		X"A0",X"A9",X"03",X"85",X"03",X"A9",X"20",X"85",X"02",X"A9",X"00",X"85",X"00",X"85",X"01",X"85",
		X"06",X"A9",X"FF",X"85",X"05",X"85",X"04",X"A2",X"01",X"38",X"A5",X"04",X"E9",X"14",X"85",X"04",
		X"A5",X"05",X"E9",X"00",X"85",X"05",X"29",X"7F",X"F0",X"19",X"18",X"A5",X"00",X"65",X"02",X"85",
		X"00",X"A5",X"01",X"65",X"03",X"85",X"01",X"A8",X"B9",X"00",X"7E",X"25",X"05",X"8D",X"00",X"90",
		X"4C",X"19",X"79",X"A5",X"06",X"D0",X"12",X"46",X"03",X"66",X"02",X"66",X"07",X"C6",X"05",X"CA",
		X"D0",X"C7",X"A9",X"01",X"85",X"06",X"4C",X"19",X"79",X"06",X"07",X"26",X"02",X"26",X"03",X"C6",
		X"05",X"E8",X"E0",X"07",X"D0",X"B3",X"4C",X"35",X"70",X"A2",X"00",X"20",X"A5",X"79",X"A9",X"00",
		X"85",X"05",X"85",X"06",X"38",X"A5",X"07",X"E5",X"03",X"85",X"07",X"A5",X"01",X"E5",X"02",X"85",
		X"01",X"A5",X"00",X"E9",X"00",X"85",X"00",X"C5",X"04",X"F0",X"17",X"18",X"A5",X"05",X"65",X"01",
		X"85",X"05",X"A5",X"06",X"65",X"00",X"85",X"06",X"A8",X"B9",X"00",X"7E",X"8D",X"00",X"90",X"4C",
		X"74",X"79",X"4C",X"35",X"70",X"A9",X"00",X"E0",X"00",X"F0",X"07",X"18",X"69",X"05",X"CA",X"4C",
		X"A9",X"79",X"AA",X"A0",X"00",X"BD",X"C2",X"79",X"99",X"00",X"00",X"E8",X"C8",X"C0",X"05",X"D0",
		X"F4",X"60",X"0E",X"AE",X"00",X"F5",X"0D",X"F8",X"06",X"F9",X"0C",X"E0",X"FA",X"1F",X"FB",X"08",
		X"4C",X"47",X"52",X"5B",X"67",X"4C",X"47",X"54",X"60",X"67",X"43",X"47",X"52",X"5B",X"67",X"23",
		X"56",X"66",X"23",X"54",X"64",X"23",X"52",X"62",X"23",X"51",X"61",X"23",X"52",X"62",X"43",X"42",
		X"50",X"56",X"64",X"23",X"49",X"59",X"23",X"4B",X"5B",X"23",X"52",X"62",X"23",X"50",X"60",X"23",
		X"49",X"59",X"23",X"47",X"57",X"13",X"7C",X"23",X"47",X"57",X"4A",X"37",X"52",X"5B",X"67",X"FF",
		X"A9",X"00",X"85",X"24",X"A9",X"7F",X"85",X"25",X"20",X"48",X"7A",X"4C",X"35",X"70",X"A9",X"59",
		X"85",X"24",X"A9",X"7F",X"85",X"25",X"20",X"48",X"7A",X"4C",X"35",X"70",X"A9",X"B0",X"85",X"24",
		X"A9",X"7F",X"85",X"25",X"20",X"48",X"7A",X"4C",X"35",X"70",X"A9",X"C7",X"85",X"24",X"A9",X"79",
		X"85",X"25",X"20",X"48",X"7A",X"4C",X"35",X"70",X"A9",X"00",X"85",X"13",X"A9",X"02",X"85",X"1A",
		X"A9",X"01",X"85",X"18",X"A9",X"03",X"85",X"19",X"20",X"8D",X"7B",X"20",X"BD",X"7A",X"58",X"C9",
		X"FF",X"F0",X"59",X"29",X"F0",X"C9",X"F0",X"D0",X"45",X"A5",X"15",X"29",X"0F",X"C9",X"07",X"B0",
		X"02",X"85",X"12",X"C9",X"08",X"D0",X"08",X"20",X"BD",X"7A",X"85",X"1A",X"4C",X"A8",X"7A",X"C9",
		X"09",X"D0",X"0D",X"20",X"BD",X"7A",X"85",X"19",X"20",X"BD",X"7A",X"85",X"18",X"4C",X"A8",X"7A",
		X"C9",X"0A",X"D0",X"08",X"20",X"BD",X"7A",X"85",X"1D",X"4C",X"A8",X"7A",X"C9",X"0B",X"D0",X"08",
		X"20",X"BD",X"7A",X"85",X"1E",X"4C",X"A8",X"7A",X"20",X"BD",X"7A",X"4C",X"5F",X"7A",X"A5",X"15",
		X"20",X"37",X"7B",X"20",X"CA",X"7A",X"20",X"BD",X"7A",X"4C",X"5F",X"7A",X"60",X"84",X"1F",X"A4",
		X"13",X"B1",X"24",X"85",X"15",X"E6",X"13",X"A4",X"1F",X"60",X"A2",X"06",X"18",X"B5",X"08",X"75",
		X"00",X"95",X"08",X"B5",X"09",X"75",X"01",X"95",X"09",X"A8",X"B9",X"00",X"7E",X"C5",X"1C",X"B0",
		X"04",X"A9",X"00",X"90",X"03",X"18",X"90",X"00",X"18",X"65",X"16",X"85",X"16",X"A5",X"17",X"69",
		X"00",X"85",X"17",X"CA",X"CA",X"10",X"D5",X"A5",X"16",X"46",X"17",X"6A",X"46",X"17",X"6A",X"8D",
		X"00",X"90",X"A9",X"00",X"85",X"16",X"85",X"17",X"18",X"A5",X"1B",X"65",X"1E",X"85",X"1B",X"A5",
		X"1C",X"69",X"00",X"85",X"1C",X"38",X"A5",X"10",X"E5",X"18",X"85",X"10",X"A5",X"11",X"E5",X"19",
		X"85",X"11",X"90",X"05",X"48",X"68",X"18",X"90",X"A1",X"A5",X"14",X"C5",X"1A",X"D0",X"03",X"20",
		X"8D",X"7B",X"C6",X"14",X"D0",X"94",X"60",X"48",X"29",X"0F",X"AA",X"BD",X"B5",X"7B",X"85",X"14",
		X"68",X"4A",X"4A",X"4A",X"4A",X"A8",X"20",X"8D",X"7B",X"20",X"BD",X"7A",X"48",X"29",X"0F",X"0A",
		X"AA",X"BD",X"9B",X"7B",X"85",X"16",X"E8",X"BD",X"9B",X"7B",X"85",X"17",X"68",X"4A",X"4A",X"4A",
		X"4A",X"85",X"12",X"38",X"A9",X"07",X"E5",X"12",X"F0",X"08",X"AA",X"46",X"17",X"66",X"16",X"CA",
		X"D0",X"F9",X"98",X"38",X"E9",X"01",X"0A",X"AA",X"A5",X"16",X"95",X"00",X"E8",X"A5",X"17",X"95",
		X"00",X"88",X"D0",X"C5",X"A9",X"00",X"85",X"1B",X"A5",X"1D",X"85",X"1C",X"60",X"A2",X"07",X"A9",
		X"00",X"95",X"00",X"A9",X"40",X"95",X"08",X"CA",X"10",X"F5",X"60",X"FB",X"4A",X"6D",X"4F",X"28",
		X"54",X"28",X"59",X"75",X"5E",X"13",X"64",X"07",X"6A",X"54",X"70",X"03",X"77",X"16",X"7E",X"95",
		X"85",X"86",X"8D",X"00",X"00",X"60",X"30",X"18",X"0C",X"06",X"20",X"10",X"08",X"04",X"02",X"90",
		X"48",X"24",X"12",X"09",X"78",X"31",X"78",X"31",X"78",X"31",X"78",X"31",X"78",X"31",X"78",X"31",
		X"78",X"31",X"78",X"31",X"71",X"14",X"71",X"14",X"71",X"14",X"71",X"98",X"73",X"F4",X"73",X"A6",
		X"74",X"4A",X"70",X"35",X"72",X"AA",X"72",X"AA",X"72",X"AA",X"72",X"AA",X"72",X"AA",X"72",X"D5",
		X"73",X"09",X"75",X"4F",X"74",X"B6",X"75",X"EA",X"76",X"BA",X"71",X"E9",X"70",X"35",X"70",X"35",
		X"70",X"35",X"70",X"35",X"78",X"FA",X"76",X"EE",X"75",X"63",X"78",X"AA",X"79",X"69",X"7A",X"10",
		X"7A",X"1E",X"7A",X"2C",X"7A",X"3A",X"70",X"35",X"70",X"00",X"70",X"35",X"70",X"35",X"70",X"35",
		X"70",X"35",X"74",X"E2",X"76",X"0B",X"70",X"35",X"70",X"35",X"00",X"03",X"03",X"03",X"03",X"03",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"05",X"03",X"04",X"03",X"03",X"03",X"03",X"03",X"03",
		X"05",X"05",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"0F",X"03",X"03",X"03",X"03",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"A9",X"00",X"85",X"00",X"85",
		X"01",X"A8",X"A9",X"02",X"85",X"02",X"A9",X"04",X"85",X"06",X"85",X"05",X"A9",X"00",X"85",X"03",
		X"85",X"04",X"18",X"A5",X"03",X"65",X"05",X"85",X"03",X"A5",X"04",X"65",X"06",X"85",X"04",X"A8",
		X"B9",X"00",X"7E",X"8D",X"00",X"90",X"18",X"A5",X"00",X"69",X"02",X"85",X"00",X"A5",X"01",X"69",
		X"00",X"85",X"01",X"90",X"DD",X"C6",X"02",X"D0",X"D9",X"4C",X"35",X"70",X"20",X"7A",X"CA",X"54",
		X"55",X"42",X"44",X"41",X"43",X"7A",X"CC",X"54",X"55",X"53",X"51",X"31",X"20",X"7A",X"E5",X"54",
		X"55",X"53",X"51",X"32",X"20",X"7A",X"E8",X"54",X"55",X"53",X"51",X"20",X"20",X"7A",X"E8",X"54",
		X"55",X"45",X"51",X"31",X"20",X"7B",X"29",X"54",X"55",X"4E",X"59",X"45",X"54",X"7B",X"32",X"54",
		X"55",X"4E",X"4F",X"54",X"45",X"7B",X"37",X"54",X"55",X"56",X"46",X"31",X"20",X"7B",X"49",X"54",
		X"55",X"44",X"49",X"56",X"20",X"7B",X"6B",X"54",X"55",X"46",X"52",X"4F",X"20",X"7B",X"72",X"54",
		X"55",X"43",X"4C",X"52",X"20",X"7B",X"8D",X"54",X"55",X"43",X"4C",X"52",X"31",X"7B",X"8F",X"4E",
		X"4F",X"54",X"56",X"41",X"4C",X"7B",X"9B",X"54",X"55",X"4E",X"44",X"55",X"52",X"7B",X"B5",X"4A",
		X"4D",X"50",X"54",X"42",X"4C",X"7B",X"C4",X"50",X"52",X"49",X"4F",X"54",X"20",X"7C",X"2A",X"53",
		X"54",X"52",X"20",X"20",X"20",X"7C",X"5B",X"53",X"54",X"52",X"54",X"54",X"20",X"00",X"00",X"53",
		X"54",X"52",X"42",X"43",X"20",X"00",X"02",X"53",X"54",X"52",X"57",X"50",X"20",X"00",X"03",X"53",
		X"54",X"52",X"50",X"49",X"20",X"00",X"05",X"53",X"54",X"52",X"4C",X"55",X"50",X"7C",X"72",X"CB",
		X"2B",X"4B",X"9B",X"DB",X"8B",X"29",X"5B",X"CB",X"0B",X"4B",X"0B",X"DB",X"8B",X"CB",X"BB",X"7B",
		X"2B",X"0B",X"4B",X"BB",X"0B",X"0B",X"0B",X"9B",X"0B",X"1B",X"8B",X"BB",X"0B",X"8B",X"8B",X"CB",
		X"0B",X"0B",X"8B",X"9B",X"1B",X"5B",X"0B",X"8B",X"8B",X"1B",X"8B",X"7B",X"0B",X"2B",X"8B",X"4B",
		X"1B",X"CB",X"8B",X"CB",X"9B",X"8B",X"8B",X"AB",X"0B",X"0B",X"CB",X"FB",X"0B",X"CB",X"1B",X"AB",
		X"0B",X"1B",X"0B",X"EB",X"0B",X"9B",X"1B",X"6B",X"0B",X"9B",X"CB",X"DB",X"0B",X"6B",X"2B",X"EB",
		X"0B",X"CB",X"BB",X"9B",X"8B",X"DB",X"9B",X"9B",X"9B",X"1B",X"8B",X"BB",X"0B",X"CB",X"DB",X"CB",
		X"0B",X"AB",X"4B",X"1B",X"0B",X"0B",X"1B",X"EB",X"0B",X"8B",X"3B",X"4B",X"1B",X"CB",X"AB",X"FB",
		X"0B",X"AB",X"0B",X"6B",X"8B",X"9B",X"9B",X"BB",X"8B",X"6B",X"5B",X"7B",X"0B",X"9B",X"1B",X"FB",
		X"0B",X"8B",X"0B",X"9B",X"1B",X"0B",X"0B",X"4B",X"4B",X"2B",X"BB",X"5B",X"0B",X"CB",X"0B",X"FB",
		X"2B",X"9B",X"0B",X"FB",X"0B",X"8B",X"4B",X"6B",X"9B",X"2B",X"8B",X"DB",X"0B",X"DB",X"CB",X"AB",
		X"8B",X"5B",X"0B",X"6B",X"0B",X"CB",X"1B",X"BB",X"4B",X"1B",X"0B",X"BB",X"4B",X"8B",X"2B",X"BB",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FD",X"FD",X"FD",X"FC",X"FB",X"FB",X"FA",X"F9",X"F8",X"F7",X"F6",
		X"F5",X"F4",X"F2",X"F1",X"F0",X"EE",X"ED",X"EB",X"E9",X"E7",X"E6",X"E4",X"E2",X"E0",X"DE",X"DC",
		X"D9",X"D7",X"D5",X"D3",X"D0",X"CE",X"CB",X"C9",X"C6",X"C4",X"C1",X"BE",X"BC",X"B9",X"B6",X"B3",
		X"B0",X"AE",X"AB",X"A8",X"A5",X"A2",X"9F",X"9C",X"99",X"96",X"93",X"8F",X"8C",X"89",X"86",X"83",
		X"80",X"7D",X"7A",X"77",X"73",X"70",X"6D",X"6A",X"67",X"64",X"61",X"5E",X"5B",X"58",X"55",X"52",
		X"4F",X"4C",X"4A",X"47",X"44",X"41",X"3F",X"3C",X"39",X"37",X"34",X"32",X"2F",X"2D",X"2B",X"28",
		X"26",X"24",X"22",X"20",X"1E",X"1C",X"1A",X"18",X"16",X"15",X"13",X"11",X"10",X"0E",X"0D",X"0C",
		X"0A",X"09",X"08",X"07",X"06",X"05",X"05",X"04",X"03",X"03",X"02",X"02",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"02",X"02",X"02",X"03",X"04",X"04",X"05",X"06",X"07",X"08",X"09",
		X"0A",X"0B",X"0D",X"0E",X"0F",X"11",X"12",X"14",X"16",X"18",X"19",X"1B",X"1D",X"1F",X"21",X"23",
		X"26",X"28",X"2A",X"2C",X"2F",X"31",X"34",X"36",X"39",X"3B",X"3E",X"41",X"43",X"46",X"49",X"4C",
		X"4F",X"51",X"54",X"57",X"5A",X"5D",X"60",X"63",X"66",X"69",X"6C",X"70",X"73",X"76",X"79",X"7C",
		X"7F",X"82",X"85",X"88",X"8C",X"8F",X"92",X"95",X"98",X"9B",X"9E",X"A1",X"A4",X"A7",X"AA",X"AD",
		X"B0",X"B3",X"B5",X"B8",X"BB",X"BE",X"C0",X"C3",X"C6",X"C8",X"CB",X"CD",X"D0",X"D2",X"D4",X"D7",
		X"D9",X"DB",X"DD",X"DF",X"E1",X"E3",X"E5",X"E7",X"E9",X"EA",X"EC",X"EE",X"EF",X"F1",X"F2",X"F3",
		X"F5",X"F6",X"F7",X"F8",X"F9",X"FA",X"FA",X"FB",X"FC",X"FC",X"FD",X"FD",X"FE",X"FE",X"FE",X"FE",
		X"F8",X"00",X"F9",X"13",X"7F",X"FA",X"00",X"FB",X"00",X"22",X"44",X"54",X"22",X"40",X"50",X"22",
		X"44",X"54",X"22",X"47",X"57",X"22",X"50",X"60",X"22",X"44",X"54",X"22",X"47",X"57",X"22",X"50",
		X"60",X"42",X"45",X"55",X"58",X"62",X"42",X"45",X"55",X"58",X"62",X"42",X"45",X"55",X"58",X"60",
		X"42",X"45",X"55",X"58",X"62",X"46",X"40",X"57",X"60",X"64",X"46",X"40",X"54",X"57",X"60",X"46",
		X"40",X"57",X"60",X"64",X"46",X"40",X"60",X"64",X"67",X"46",X"40",X"57",X"60",X"64",X"46",X"40",
		X"60",X"64",X"67",X"42",X"40",X"64",X"67",X"70",X"FF",X"F8",X"00",X"F9",X"1C",X"20",X"FA",X"1F",
		X"FB",X"00",X"12",X"49",X"22",X"49",X"54",X"22",X"49",X"59",X"22",X"49",X"60",X"22",X"49",X"5B",
		X"22",X"49",X"54",X"22",X"48",X"5B",X"22",X"48",X"62",X"22",X"49",X"60",X"12",X"44",X"22",X"49",
		X"64",X"12",X"50",X"22",X"4B",X"58",X"12",X"44",X"22",X"4B",X"64",X"12",X"52",X"22",X"50",X"59",
		X"12",X"54",X"22",X"49",X"59",X"12",X"60",X"22",X"48",X"5B",X"12",X"54",X"22",X"44",X"5B",X"12",
		X"62",X"22",X"49",X"60",X"12",X"44",X"22",X"49",X"59",X"12",X"50",X"32",X"49",X"59",X"69",X"FF",
		X"F8",X"0A",X"F9",X"14",X"D0",X"FA",X"00",X"FB",X"00",X"32",X"40",X"50",X"60",X"22",X"47",X"67",
		X"22",X"47",X"62",X"42",X"47",X"52",X"5B",X"64",X"32",X"40",X"50",X"60",X"22",X"47",X"67",X"22",
		X"47",X"62",X"42",X"47",X"52",X"5B",X"64",X"31",X"40",X"50",X"60",X"11",X"7C",X"41",X"50",X"54",
		X"67",X"70",X"12",X"7C",X"42",X"40",X"47",X"54",X"60",X"4A",X"40",X"47",X"54",X"60",X"FF",X"2B",
		X"7B",X"3B",X"DB",X"4B",X"FB",X"7B",X"6B",X"0B",X"6B",X"6B",X"20",X"72",X"03",X"70",X"89",X"70");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
