library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity mpa_33k is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of mpa_33k is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"DD",X"34",X"00",X"DD",X"7E",X"0C",X"E6",X"7F",X"C8",X"CD",X"28",X"1F",X"DD",X"7E",X"00",X"FE",
		X"25",X"CA",X"83",X"1F",X"FE",X"24",X"CA",X"AA",X"1E",X"C9",X"CD",X"63",X"1C",X"CD",X"DB",X"20",
		X"22",X"D6",X"E0",X"7C",X"D6",X"08",X"FE",X"F0",X"D2",X"52",X"08",X"ED",X"5B",X"DC",X"E0",X"2A",
		X"DA",X"E0",X"19",X"22",X"DA",X"E0",X"7C",X"FE",X"30",X"DA",X"52",X"08",X"7A",X"A7",X"FA",X"78",
		X"1F",X"21",X"00",X"00",X"A7",X"ED",X"52",X"22",X"DC",X"E0",X"C3",X"78",X"1F",X"3A",X"03",X"E3",
		X"16",X"00",X"C6",X"10",X"DD",X"96",X"03",X"30",X"03",X"ED",X"44",X"15",X"1F",X"1F",X"1F",X"E6",
		X"1E",X"4F",X"06",X"00",X"21",X"24",X"2D",X"09",X"FE",X"12",X"38",X"01",X"04",X"7E",X"CB",X"7A",
		X"28",X"06",X"2F",X"5F",X"78",X"2F",X"47",X"7B",X"DD",X"77",X"04",X"DD",X"70",X"05",X"23",X"5E",
		X"16",X"00",X"79",X"FE",X"0A",X"30",X"01",X"14",X"DD",X"72",X"09",X"DD",X"73",X"08",X"DD",X"36",
		X"00",X"29",X"2A",X"1A",X"E3",X"DD",X"75",X"0B",X"DD",X"74",X"0F",X"C9",X"CD",X"63",X"1C",X"CD",
		X"FB",X"20",X"22",X"D6",X"E0",X"7C",X"2A",X"DC",X"E0",X"C3",X"F1",X"1C",X"DD",X"35",X"0A",X"C2",
		X"B8",X"08",X"DD",X"36",X"0A",X"06",X"DD",X"7E",X"0D",X"FE",X"39",X"D2",X"52",X"08",X"DD",X"34",
		X"0D",X"C3",X"B8",X"08",X"DD",X"35",X"0A",X"C2",X"B8",X"08",X"DD",X"7E",X"07",X"FE",X"80",X"D2",
		X"52",X"08",X"06",X"80",X"DD",X"36",X"00",X"00",X"C3",X"69",X"08",X"DD",X"E5",X"E1",X"11",X"D4",
		X"E0",X"01",X"0A",X"00",X"ED",X"B0",X"ED",X"5B",X"D6",X"E0",X"2A",X"D8",X"E0",X"19",X"C9",X"DD",
		X"E5",X"D1",X"21",X"D4",X"E0",X"01",X"0A",X"00",X"ED",X"B0",X"C9",X"CD",X"DB",X"20",X"EB",X"DD",
		X"6E",X"0B",X"DD",X"66",X"0F",X"ED",X"4B",X"1A",X"E3",X"ED",X"42",X"19",X"C9",X"21",X"51",X"E0",
		X"3A",X"00",X"E3",X"3D",X"28",X"11",X"7E",X"A7",X"F0",X"21",X"11",X"E5",X"3E",X"01",X"86",X"27",
		X"77",X"23",X"7E",X"CE",X"00",X"27",X"77",X"3E",X"37",X"32",X"51",X"E0",X"11",X"90",X"80",X"FD",
		X"21",X"90",X"84",X"0E",X"02",X"CD",X"E7",X"03",X"3A",X"12",X"E5",X"CD",X"BD",X"03",X"3A",X"11",
		X"E5",X"C3",X"AE",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"06",X"01",X"03",X"34",X"07",X"49",X"08",X"63",X"0F",X"73",X"07",X"80",X"19",X"92",X"0F",
		X"A0",X"06",X"A1",X"03",X"A2",X"2A",X"E0",X"32",X"FF",X"28",X"0F",X"0F",X"3F",X"30",X"40",X"06",
		X"41",X"03",X"42",X"2A",X"4C",X"0F",X"92",X"0F",X"9F",X"28",X"A5",X"07",X"B8",X"0F",X"CD",X"0F",
		X"E0",X"06",X"E1",X"03",X"00",X"19",X"01",X"08",X"14",X"07",X"20",X"33",X"4F",X"0F",X"7F",X"30",
		X"80",X"06",X"81",X"03",X"82",X"22",X"9C",X"1C",X"B6",X"1C",X"C0",X"2A",X"D9",X"1C",X"DF",X"20",
		X"03",X"0F",X"08",X"28",X"16",X"07",X"20",X"06",X"21",X"03",X"3C",X"22",X"52",X"1C",X"60",X"32",
		X"6E",X"1C",X"7F",X"20",X"A6",X"08",X"B7",X"0F",X"BF",X"30",X"C0",X"06",X"C1",X"03",X"C4",X"08",
		X"D3",X"0A",X"E6",X"0E",X"F6",X"0F",X"0C",X"10",X"1C",X"0F",X"2D",X"0E",X"39",X"07",X"4A",X"0F",
		X"5B",X"0F",X"60",X"06",X"61",X"03",X"6E",X"19",X"6F",X"09",X"82",X"0F",X"8F",X"09",X"A0",X"2B",
		X"A2",X"0F",X"B1",X"0F",X"FF",X"28",X"00",X"06",X"01",X"03",X"02",X"22",X"14",X"1C",X"28",X"1C",
		X"40",X"2A",X"54",X"1C",X"5F",X"20",X"9F",X"28",X"A0",X"06",X"A1",X"03",X"A2",X"23",X"A6",X"1C",
		X"D3",X"1C",X"E9",X"0F",X"F7",X"0A",X"FF",X"20",X"07",X"10",X"17",X"0E",X"29",X"10",X"35",X"0A",
		X"40",X"06",X"41",X"02",X"42",X"1A",X"60",X"03",X"6F",X"12",X"78",X"12",X"88",X"12",X"92",X"12",
		X"A3",X"12",X"A4",X"12",X"B1",X"12",X"C2",X"12",X"CD",X"12",X"CE",X"12",X"D9",X"12",X"E0",X"06",
		X"E1",X"03",X"EB",X"12",X"FA",X"12",X"06",X"12",X"07",X"12",X"14",X"12",X"23",X"12",X"2C",X"12",
		X"37",X"12",X"42",X"12",X"56",X"12",X"57",X"12",X"65",X"12",X"6E",X"12",X"7A",X"12",X"80",X"06",
		X"81",X"03",X"85",X"12",X"86",X"12",X"91",X"12",X"92",X"12",X"A3",X"12",X"A4",X"12",X"AE",X"12",
		X"B8",X"12",X"B9",X"12",X"CA",X"12",X"CB",X"12",X"D7",X"12",X"E3",X"12",X"F3",X"12",X"00",X"19",
		X"20",X"06",X"21",X"03",X"22",X"2C",X"60",X"33",X"9F",X"28",X"BF",X"30",X"C0",X"06",X"C1",X"03",
		X"C2",X"24",X"D5",X"1C",X"EA",X"1C",X"00",X"33",X"05",X"1C",X"18",X"1C",X"31",X"1C",X"3F",X"20",
		X"48",X"30",X"60",X"06",X"61",X"03",X"7B",X"24",X"87",X"1C",X"99",X"1C",X"A0",X"2B",X"AE",X"1C",
		X"C5",X"1C",X"D7",X"1C",X"DF",X"20",X"E0",X"28",X"00",X"06",X"01",X"04",X"13",X"14",X"1E",X"16",
		X"2D",X"16",X"2F",X"16",X"3A",X"15",X"4C",X"16",X"4E",X"16",X"58",X"16",X"66",X"16",X"68",X"16",
		X"72",X"02",X"73",X"14",X"7E",X"16",X"80",X"19",X"A0",X"86",X"A1",X"03",X"A2",X"34",X"C7",X"0F",
		X"EC",X"10",X"0F",X"0A",X"1F",X"30",X"2A",X"10",X"40",X"86",X"41",X"02",X"42",X"19",X"60",X"32",
		X"61",X"05",X"80",X"2A",X"BF",X"30",X"C0",X"02",X"DF",X"28",X"E0",X"06",X"E1",X"03",X"E2",X"2B",
		X"00",X"23",X"01",X"03",X"2A",X"1C",X"3F",X"28",X"45",X"1C",X"57",X"1C",X"6C",X"1C",X"6D",X"20",
		X"80",X"06",X"81",X"02",X"A0",X"03",X"A8",X"10",X"B4",X"0A",X"C5",X"07",X"DC",X"0F",X"E3",X"09",
		X"F2",X"07",X"0A",X"10",X"0D",X"09",X"1C",X"08",X"20",X"06",X"21",X"03",X"2C",X"0F",X"2F",X"0F",
		X"32",X"0A",X"45",X"13",X"54",X"13",X"66",X"13",X"77",X"0A",X"8A",X"13",X"98",X"13",X"A7",X"13",
		X"B4",X"13",X"C0",X"06",X"C1",X"03",X"C5",X"09",X"D4",X"0A",X"E0",X"02",X"E7",X"0A",X"F5",X"09",
		X"00",X"04",X"1C",X"16",X"2A",X"15",X"2C",X"15",X"35",X"16",X"3D",X"14",X"40",X"02",X"48",X"14",
		X"4A",X"14",X"60",X"86",X"61",X"02",X"62",X"19",X"80",X"03",X"81",X"2C",X"A0",X"33",X"DF",X"28",
		X"FF",X"30",X"00",X"86",X"01",X"03",X"02",X"2C",X"40",X"23",X"57",X"1C",X"5F",X"28",X"6C",X"1C",
		X"83",X"1C",X"9A",X"1C",X"A0",X"86",X"A1",X"03",X"A2",X"23",X"AE",X"1C",X"C5",X"1C",X"D5",X"1C",
		X"E0",X"33",X"E8",X"1C",X"F5",X"0F",X"FF",X"20",X"0A",X"09",X"1C",X"0A",X"28",X"30",X"32",X"10",
		X"40",X"06",X"42",X"02",X"5B",X"2B",X"60",X"03",X"80",X"33",X"9F",X"28",X"D0",X"30",X"E0",X"06",
		X"E1",X"03",X"E2",X"1B",X"20",X"17",X"60",X"18",X"80",X"06",X"81",X"03",X"C6",X"13",X"D2",X"0F",
		X"DD",X"0F",X"EE",X"0E",X"FC",X"0A",X"01",X"13",X"0D",X"09",X"20",X"06",X"21",X"03",X"22",X"13",
		X"2B",X"13",X"39",X"13",X"49",X"13",X"4C",X"0A",X"5C",X"0F",X"6A",X"0F",X"79",X"13",X"84",X"13",
		X"86",X"0A",X"95",X"0F",X"A4",X"13",X"B3",X"13",X"B5",X"09",X"C0",X"06",X"C1",X"02",X"C2",X"19",
		X"E0",X"03",X"E1",X"2C",X"EA",X"07",X"F9",X"09",X"07",X"0A",X"19",X"0F",X"2A",X"0F",X"39",X"09",
		X"48",X"28",X"54",X"0F",X"60",X"06",X"61",X"03",X"7B",X"23",X"84",X"1C",X"92",X"1C",X"A0",X"23",
		X"A3",X"1C",X"B3",X"1C",X"C3",X"1C",X"DC",X"1C",X"EF",X"1C",X"FF",X"20",X"00",X"06",X"01",X"03",
		X"07",X"10",X"0A",X"0A",X"1A",X"0F",X"2C",X"09",X"32",X"0F",X"41",X"07",X"4F",X"08",X"5C",X"0F",
		X"63",X"09",X"70",X"07",X"7D",X"0E",X"80",X"19",X"A0",X"06",X"A1",X"03",X"A2",X"24",X"AF",X"1C",
		X"BC",X"1C",X"C0",X"2C",X"CA",X"1C",X"D9",X"1C",X"E8",X"1C",X"F6",X"1C",X"FF",X"28",X"05",X"0A",
		X"10",X"1C",X"11",X"20",X"25",X"0C",X"32",X"0F",X"35",X"0C",X"40",X"06",X"41",X"03",X"42",X"19",
		X"60",X"33",X"80",X"2B",X"83",X"0A",X"92",X"07",X"BF",X"30",X"C6",X"0F",X"C9",X"0A",X"D9",X"09",
		X"DF",X"28",X"E0",X"06",X"E1",X"03",X"E2",X"24",X"EA",X"1C",X"04",X"0A",X"14",X"0F",X"1C",X"1C",
		X"24",X"20",X"34",X"09",X"45",X"0F",X"49",X"0F",X"4B",X"0C",X"58",X"0C",X"67",X"0C",X"75",X"0C",
		X"7A",X"0F",X"80",X"06",X"81",X"02",X"90",X"04",X"AD",X"16",X"B7",X"15",X"BE",X"14",X"C5",X"16",
		X"C7",X"16",X"D4",X"14",X"DB",X"15",X"E6",X"14",X"E8",X"14",X"E9",X"16",X"F0",X"14",X"F1",X"16",
		X"F2",X"14",X"02",X"15",X"04",X"15",X"0E",X"16",X"0F",X"02",X"10",X"14",X"13",X"16",X"17",X"14",
		X"19",X"14",X"20",X"86",X"21",X"03",X"22",X"19",X"40",X"2C",X"41",X"33",X"42",X"03",X"BE",X"28",
		X"BF",X"30",X"C0",X"86",X"C1",X"03",X"C2",X"1A",X"E8",X"12",X"F2",X"12",X"F4",X"12",X"FD",X"12",
		X"08",X"12",X"13",X"12",X"22",X"12",X"23",X"12",X"2E",X"12",X"36",X"12",X"42",X"12",X"4E",X"12",
		X"57",X"12",X"60",X"86",X"61",X"03",X"65",X"12",X"67",X"12",X"72",X"12",X"7A",X"12",X"83",X"12",
		X"8F",X"12",X"97",X"12",X"A2",X"12",X"AB",X"12",X"B7",X"12",X"C2",X"12",X"D0",X"12",X"D8",X"12",
		X"E4",X"12",X"00",X"86",X"01",X"03",X"20",X"25",X"25",X"09",X"33",X"1C",X"40",X"2C",X"48",X"10",
		X"54",X"1C",X"65",X"0F",X"6F",X"1C",X"7F",X"20",X"80",X"02",X"88",X"28",X"A0",X"86",X"A1",X"05",
		X"BB",X"35",X"C0",X"2C",X"DF",X"02",X"FF",X"30",X"0A",X"10",X"19",X"0A",X"1F",X"28",X"20",X"03",
		X"29",X"0F",X"2C",X"0A",X"32",X"0F",X"3A",X"0F",X"40",X"06",X"41",X"02",X"47",X"0F",X"4A",X"0A",
		X"50",X"0F",X"60",X"03",X"65",X"07",X"79",X"08",X"80",X"17",X"8A",X"0A",X"A0",X"18",X"C8",X"09",
		X"E0",X"06",X"E1",X"03",X"EF",X"10",X"F4",X"0F",X"F7",X"0A",X"06",X"0F",X"11",X"10",X"14",X"09",
		X"1A",X"1A",X"3A",X"12",X"42",X"12",X"44",X"12",X"4E",X"12",X"57",X"12",X"59",X"12",X"63",X"12",
		X"6B",X"12",X"80",X"06",X"81",X"02",X"8F",X"13",X"92",X"0A",X"A0",X"03",X"A5",X"10",X"A8",X"07",
		X"B2",X"0F",X"B5",X"0F",X"C5",X"13",X"D4",X"09",X"E4",X"0F",X"E6",X"0C",X"F4",X"0C",X"04",X"10",
		X"06",X"0C",X"13",X"0C",X"20",X"06",X"21",X"03",X"22",X"10",X"23",X"19",X"28",X"10",X"2A",X"0A",
		X"3B",X"10",X"40",X"25",X"41",X"33",X"4A",X"1C",X"55",X"1C",X"65",X"1C",X"74",X"1C",X"82",X"0F",
		X"88",X"1C",X"95",X"0F",X"A5",X"1C",X"A8",X"30",X"B1",X"1C",X"B2",X"20",X"BE",X"0F",X"C0",X"06",
		X"C1",X"02",X"C2",X"1B",X"CA",X"10",X"E0",X"03",X"E6",X"0A",X"F0",X"17",X"03",X"08",X"12",X"18",
		X"13",X"09",X"40",X"1A",X"4A",X"0A",X"60",X"06",X"61",X"03",X"74",X"12",X"85",X"12",X"87",X"12",
		X"92",X"12",X"94",X"12",X"A9",X"12",X"AA",X"12",X"B4",X"10",X"BD",X"12",X"C3",X"12",X"CC",X"0F",
		X"D5",X"12",X"D7",X"12",X"E5",X"12",X"E7",X"12",X"F4",X"12",X"00",X"06",X"01",X"02",X"02",X"25",
		X"03",X"2C",X"0A",X"1C",X"17",X"1C",X"20",X"03",X"27",X"10",X"37",X"1C",X"48",X"1C",X"59",X"1C",
		X"6A",X"0A",X"79",X"1C",X"80",X"28",X"8D",X"0F",X"90",X"1C",X"91",X"20",X"A0",X"06",X"A1",X"03",
		X"AD",X"0C",X"B2",X"0F",X"BB",X"0C",X"CB",X"0C",X"D8",X"0F",X"E5",X"0F",X"E7",X"10",X"F1",X"0F",
		X"F9",X"0F",X"08",X"0C",X"0D",X"0F",X"16",X"0C",X"20",X"19",X"25",X"0F",X"28",X"09",X"36",X"10",
		X"40",X"06",X"41",X"02",X"42",X"25",X"4A",X"1C",X"5A",X"0F",X"60",X"03",X"61",X"2C",X"65",X"10",
		X"79",X"1C",X"88",X"1C",X"94",X"1C",X"A2",X"1C",X"AE",X"1C",X"BB",X"1C",X"BF",X"20",X"CA",X"0F",
		X"D0",X"28",X"DC",X"10",X"E0",X"06",X"E1",X"03",X"E8",X"0F",X"EA",X"10",X"EC",X"0A",X"F9",X"0F",
		X"08",X"13",X"0A",X"07",X"17",X"0F",X"1A",X"0A",X"2A",X"0C",X"37",X"10",X"3C",X"0C",X"43",X"02",
		X"80",X"06",X"00",X"06",X"20",X"03",X"28",X"10",X"34",X"0A",X"47",X"0C",X"55",X"0C",X"5A",X"0F",
		X"63",X"09",X"72",X"07",X"85",X"13",X"94",X"13",X"A0",X"06",X"A1",X"04",X"B3",X"14",X"BF",X"16",
		X"CD",X"16",X"DA",X"15",X"EC",X"16",X"EE",X"16",X"F8",X"16",X"F9",X"03",X"00",X"2B",X"20",X"23",
		X"40",X"86",X"4A",X"1C",X"50",X"28",X"65",X"1C",X"77",X"1C",X"7E",X"05",X"7F",X"20",X"80",X"33",
		X"C8",X"03",X"CF",X"30",X"E0",X"06",X"00",X"17",X"20",X"18",X"6A",X"0A",X"73",X"07",X"01",X"02",
		X"20",X"01",X"34",X"C0",X"3A",X"C2",X"48",X"20",X"54",X"C2",X"59",X"20",X"64",X"C2",X"69",X"E2",
		X"6D",X"C2",X"76",X"22",X"82",X"20",X"90",X"C0",X"96",X"C0",X"9C",X"C0",X"A2",X"C0",X"BE",X"C1",
		X"CB",X"C0",X"D8",X"20",X"E6",X"C2",X"F4",X"22",X"00",X"C2",X"05",X"FF",X"4D",X"00",X"4E",X"02",
		X"5E",X"22",X"77",X"22",X"8A",X"22",X"8B",X"FF",X"D8",X"00",X"E0",X"02",X"45",X"22",X"55",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"21",X"46",X"E0",X"35",X"FB",X"78",X"32",X"13",X"E5",X"FE",X"05",X"CA",X"D2",X"27",X"A7",X"C2",
		X"5E",X"28",X"CD",X"FA",X"29",X"3E",X"1E",X"CD",X"75",X"0D",X"21",X"0F",X"E5",X"36",X"00",X"23",
		X"34",X"CD",X"48",X"29",X"CD",X"E8",X"05",X"21",X"24",X"2C",X"CD",X"00",X"03",X"CD",X"BA",X"28",
		X"21",X"0C",X"2C",X"CD",X"00",X"03",X"3A",X"13",X"E5",X"17",X"17",X"17",X"17",X"26",X"00",X"E6",
		X"F0",X"6F",X"20",X"01",X"24",X"22",X"98",X"E0",X"CD",X"71",X"29",X"2A",X"96",X"E0",X"56",X"2B",
		X"5E",X"2A",X"11",X"E5",X"A7",X"ED",X"52",X"30",X"0E",X"19",X"EB",X"2A",X"96",X"E0",X"72",X"2B",
		X"73",X"21",X"39",X"2C",X"CD",X"4E",X"03",X"2A",X"94",X"E0",X"ED",X"5B",X"11",X"E5",X"7D",X"D6",
		X"01",X"27",X"6F",X"30",X"01",X"25",X"22",X"94",X"E0",X"A7",X"ED",X"52",X"38",X"50",X"CD",X"68",
		X"29",X"2A",X"98",X"E0",X"7D",X"C6",X"01",X"27",X"6F",X"30",X"01",X"24",X"22",X"98",X"E0",X"CD",
		X"71",X"29",X"3E",X"10",X"CD",X"75",X"0D",X"3E",X"0C",X"CD",X"EA",X"05",X"18",X"C9",X"3E",X"1D",
		X"CD",X"75",X"0D",X"CD",X"D6",X"29",X"CD",X"12",X"0D",X"CD",X"48",X"29",X"3E",X"30",X"CD",X"EA",
		X"05",X"CD",X"BA",X"28",X"38",X"0D",X"21",X"E4",X"2B",X"CD",X"4E",X"03",X"3A",X"F9",X"E0",X"3C",
		X"C3",X"F9",X"27",X"21",X"F9",X"2B",X"CD",X"4E",X"03",X"CD",X"E8",X"05",X"18",X"0E",X"CD",X"E8",
		X"05",X"11",X"01",X"E5",X"21",X"98",X"E0",X"06",X"02",X"CD",X"36",X"06",X"21",X"00",X"00",X"22",
		X"11",X"E5",X"21",X"13",X"E5",X"7E",X"A7",X"C2",X"B7",X"0B",X"36",X"05",X"21",X"A2",X"23",X"22",
		X"16",X"E5",X"3E",X"1A",X"32",X"0E",X"E5",X"C3",X"B7",X"0B",X"CD",X"E8",X"05",X"CD",X"5A",X"29",
		X"3A",X"10",X"E5",X"D6",X"02",X"28",X"07",X"3E",X"0A",X"FA",X"CE",X"28",X"3E",X"05",X"5F",X"3A",
		X"13",X"E5",X"01",X"80",X"00",X"FE",X"08",X"30",X"09",X"01",X"00",X"01",X"FE",X"03",X"30",X"02",
		X"0E",X"20",X"ED",X"43",X"94",X"E0",X"83",X"87",X"5F",X"FE",X"0A",X"20",X"09",X"3A",X"10",X"E5",
		X"FE",X"03",X"28",X"02",X"1E",X"14",X"16",X"00",X"21",X"0C",X"E0",X"19",X"7E",X"23",X"22",X"96",
		X"E0",X"B6",X"20",X"03",X"70",X"2B",X"71",X"21",X"79",X"2B",X"CD",X"4E",X"03",X"CD",X"81",X"29",
		X"A7",X"20",X"02",X"3E",X"1A",X"C6",X"40",X"1B",X"1B",X"12",X"21",X"94",X"2B",X"CD",X"4E",X"03",
		X"21",X"12",X"E5",X"13",X"CD",X"9A",X"03",X"21",X"B0",X"2B",X"CD",X"4E",X"03",X"CD",X"68",X"29",
		X"21",X"CC",X"2B",X"CD",X"4E",X"03",X"2A",X"96",X"E0",X"13",X"CD",X"9A",X"03",X"2A",X"94",X"E0",
		X"ED",X"5B",X"11",X"E5",X"A7",X"ED",X"52",X"C9",X"21",X"00",X"E1",X"01",X"A4",X"00",X"CD",X"FA",
		X"05",X"01",X"20",X"02",X"21",X"E0",X"80",X"C3",X"FA",X"05",X"21",X"00",X"E1",X"01",X"C6",X"00",
		X"CD",X"FA",X"05",X"01",X"20",X"03",X"18",X"EC",X"11",X"D9",X"81",X"21",X"95",X"E0",X"C3",X"9A",
		X"03",X"21",X"99",X"E0",X"11",X"97",X"82",X"CD",X"93",X"03",X"EB",X"36",X"30",X"23",X"36",X"30",
		X"C9",X"3A",X"0E",X"E5",X"FE",X"1A",X"D8",X"D6",X"1A",X"C9",X"21",X"CC",X"80",X"11",X"CC",X"84",
		X"01",X"02",X"10",X"CD",X"E7",X"03",X"79",X"36",X"21",X"12",X"23",X"13",X"10",X"F9",X"21",X"CC",
		X"80",X"06",X"05",X"34",X"23",X"23",X"23",X"10",X"FA",X"36",X"1B",X"CD",X"81",X"29",X"21",X"CC",
		X"80",X"06",X"05",X"FE",X"05",X"38",X"0C",X"16",X"03",X"36",X"29",X"23",X"15",X"20",X"FA",X"D6",
		X"05",X"10",X"F0",X"57",X"87",X"87",X"82",X"5F",X"FE",X"08",X"38",X"10",X"28",X"01",X"3D",X"36",
		X"29",X"23",X"D6",X"08",X"18",X"F2",X"2A",X"F4",X"E0",X"3A",X"F6",X"E0",X"3C",X"57",X"C6",X"21",
		X"CB",X"66",X"28",X"07",X"D6",X"06",X"FE",X"20",X"20",X"01",X"3D",X"77",X"7A",X"FE",X"08",X"38",
		X"02",X"AF",X"2C",X"32",X"F6",X"E0",X"22",X"F4",X"E0",X"C9",X"21",X"CC",X"80",X"06",X"0F",X"36",
		X"29",X"23",X"10",X"FB",X"36",X"1F",X"3E",X"5A",X"32",X"52",X"80",X"C9",X"00",X"00",X"00",X"20",
		X"00",X"00",X"50",X"00",X"00",X"80",X"00",X"00",X"00",X"01",X"00",X"00",X"02",X"00",X"00",X"03",
		X"00",X"00",X"05",X"00",X"00",X"08",X"00",X"00",X"10",X"00",X"08",X"81",X"08",X"54",X"4F",X"20",
		X"43",X"4F",X"55",X"4E",X"54",X"49",X"4E",X"55",X"45",X"20",X"47",X"41",X"4D",X"45",X"22",X"2D",
		X"82",X"08",X"54",X"49",X"4D",X"45",X"21",X"46",X"81",X"08",X"42",X"45",X"47",X"49",X"4E",X"4E",
		X"45",X"52",X"20",X"43",X"4F",X"55",X"52",X"53",X"45",X"20",X"47",X"4F",X"20",X"5B",X"21",X"46",
		X"81",X"00",X"43",X"48",X"41",X"4D",X"50",X"49",X"4F",X"4E",X"20",X"43",X"4F",X"55",X"52",X"53",
		X"45",X"20",X"31",X"20",X"47",X"4F",X"20",X"5B",X"21",X"4C",X"82",X"00",X"46",X"52",X"45",X"45",
		X"20",X"50",X"4C",X"41",X"59",X"21",X"EA",X"81",X"00",X"4F",X"4E",X"4C",X"59",X"20",X"31",X"20",
		X"50",X"4C",X"41",X"59",X"45",X"52",X"21",X"EA",X"81",X"00",X"31",X"20",X"4F",X"52",X"20",X"32",
		X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"53",X"21",X"06",X"82",X"00",X"50",X"49",X"43",X"54",
		X"55",X"52",X"45",X"20",X"4E",X"55",X"4D",X"42",X"45",X"52",X"20",X"53",X"45",X"54",X"22",X"4A",
		X"82",X"00",X"4E",X"45",X"58",X"54",X"20",X"31",X"50",X"20",X"42",X"55",X"54",X"54",X"4F",X"4E",
		X"21",X"6A",X"81",X"00",X"20",X"50",X"55",X"53",X"48",X"20",X"42",X"55",X"54",X"54",X"4F",X"4E",
		X"20",X"21",X"D4",X"83",X"00",X"43",X"52",X"45",X"44",X"49",X"54",X"20",X"21",X"88",X"81",X"00",
		X"47",X"41",X"4D",X"45",X"20",X"4F",X"56",X"45",X"52",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",
		X"20",X"21",X"0C",X"82",X"00",X"47",X"41",X"4D",X"45",X"20",X"4F",X"56",X"45",X"52",X"21",X"2B",
		X"80",X"02",X"04",X"25",X"0F",X"14",X"05",X"22",X"41",X"80",X"01",X"0C",X"0D",X"25",X"06",X"00",
		X"22",X"49",X"80",X"09",X"3F",X"22",X"4B",X"80",X"02",X"06",X"50",X"4F",X"49",X"4E",X"54",X"25",
		X"04",X"00",X"12",X"25",X"05",X"00",X"07",X"22",X"6B",X"80",X"02",X"06",X"25",X"09",X"00",X"12",
		X"25",X"05",X"00",X"07",X"22",X"8B",X"80",X"02",X"06",X"0E",X"0F",X"10",X"11",X"25",X"05",X"00",
		X"12",X"25",X"05",X"00",X"07",X"22",X"AB",X"80",X"02",X"08",X"16",X"15",X"15",X"17",X"15",X"15",
		X"18",X"15",X"15",X"19",X"15",X"15",X"1A",X"15",X"15",X"09",X"22",X"81",X"80",X"01",X"31",X"50",
		X"3F",X"21",X"A1",X"80",X"01",X"32",X"50",X"3F",X"21",X"25",X"81",X"01",X"54",X"49",X"4D",X"45",
		X"20",X"54",X"4F",X"20",X"52",X"45",X"41",X"43",X"48",X"20",X"50",X"4F",X"49",X"4E",X"54",X"20",
		X"5E",X"00",X"5E",X"21",X"84",X"81",X"00",X"59",X"4F",X"55",X"52",X"20",X"54",X"49",X"4D",X"45",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"22",X"97",X"81",X"01",X"5D",X"21",
		X"C4",X"81",X"00",X"54",X"48",X"45",X"20",X"41",X"56",X"45",X"52",X"41",X"47",X"45",X"20",X"54",
		X"49",X"4D",X"45",X"20",X"20",X"20",X"22",X"D7",X"81",X"01",X"5D",X"21",X"04",X"82",X"01",X"54",
		X"4F",X"50",X"20",X"52",X"45",X"43",X"4F",X"52",X"44",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"5D",X"21",X"85",X"82",X"00",X"47",X"4F",X"4F",X"44",X"20",X"42",X"4F",X"4E",X"55",
		X"53",X"20",X"50",X"4F",X"49",X"4E",X"54",X"53",X"21",X"67",X"82",X"00",X"53",X"4F",X"52",X"52",
		X"59",X"20",X"4E",X"4F",X"20",X"42",X"4F",X"4E",X"55",X"53",X"5B",X"21",X"65",X"82",X"01",X"53",
		X"50",X"45",X"43",X"49",X"41",X"4C",X"20",X"42",X"4F",X"4E",X"55",X"53",X"20",X"50",X"4F",X"49",
		X"4E",X"54",X"53",X"21",X"25",X"81",X"00",X"43",X"4F",X"4E",X"47",X"52",X"41",X"54",X"55",X"4C",
		X"41",X"54",X"49",X"4F",X"4E",X"53",X"20",X"5B",X"21",X"E5",X"82",X"01",X"59",X"4F",X"55",X"20",
		X"48",X"41",X"56",X"45",X"20",X"42",X"52",X"4F",X"4B",X"45",X"4E",X"20",X"41",X"20",X"52",X"45",
		X"43",X"4F",X"52",X"44",X"20",X"5B",X"21",X"6A",X"81",X"00",X"49",X"4E",X"53",X"45",X"52",X"54",
		X"20",X"43",X"4F",X"49",X"4E",X"20",X"21",X"C7",X"81",X"00",X"31",X"20",X"50",X"4C",X"41",X"59",
		X"45",X"52",X"20",X"20",X"20",X"31",X"20",X"43",X"4F",X"49",X"4E",X"20",X"21",X"C5",X"81",X"00",
		X"41",X"20",X"5F",X"20",X"31",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"20",X"20",X"20",X"31",
		X"20",X"43",X"4F",X"49",X"4E",X"20",X"21",X"C8",X"82",X"00",X"5C",X"31",X"39",X"38",X"32",X"20",
		X"49",X"52",X"45",X"4D",X"20",X"43",X"4F",X"52",X"50",X"2F",X"21",X"76",X"80",X"02",X"3A",X"3B",
		X"3C",X"3D",X"3E",X"21",X"F0",X"F0",X"ED",X"F0",X"F0",X"FB",X"FB",X"FB",X"F0",X"E8",X"F0",X"F0",
		X"F0",X"EE",X"F0",X"F0",X"F0",X"F0",X"E0",X"F0",X"F0",X"FB",X"FB",X"FB",X"F0",X"F0",X"F0",X"F2",
		X"F2",X"F0",X"F0",X"F0",X"E9",X"F2",X"EF",X"E3",X"D2",X"FC",X"FD",X"FE",X"E0",X"D4",X"D3",X"EB",
		X"FF",X"D5",X"F1",X"E5",X"E2",X"D0",X"D6",X"E6",X"D7",X"F0",X"E1",X"D8",X"F9",X"FB",X"F0",X"F2",
		X"D9",X"EC",X"FC",X"D1",X"34",X"32",X"32",X"43",X"34",X"23",X"32",X"11",X"23",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"12",X"12",X"12",X"24",X"77",X"21",X"10",X"56",X"21",X"10",X"34",X"21",
		X"23",X"23",X"21",X"31",X"22",X"21",X"11",X"00",X"77",X"77",X"66",X"65",X"55",X"44",X"43",X"33",
		X"43",X"33",X"21",X"31",X"00",X"9A",X"51",X"98",X"8D",X"5F",X"B6",X"30",X"D2",X"06",X"E3",X"E3",
		X"EF",X"C7",X"F7",X"B0",X"FC",X"9E",X"00",X"8E",X"03",X"82",X"06",X"77",X"07",X"6E",X"08",X"66",
		X"09",X"5F",X"0A",X"59",X"03",X"48",X"81",X"B0",X"B1",X"B2",X"B3",X"B4",X"02",X"B5",X"B6",X"B7",
		X"B8",X"02",X"B9",X"BA",X"BB",X"BC",X"BD",X"02",X"BE",X"BF",X"C0",X"C1",X"C2",X"02",X"C3",X"C4",
		X"C5",X"C6",X"BD",X"02",X"03",X"6D",X"81",X"C7",X"C8",X"C9",X"CA",X"02",X"CB",X"BF",X"CC",X"02",
		X"CD",X"BC",X"CE",X"CF",X"02",X"D0",X"D1",X"D2",X"CA",X"02",X"D3",X"D4",X"D5",X"C2",X"02",X"D6",
		X"D7",X"BC",X"BD",X"02",X"D8",X"C0",X"C1",X"C2",X"02",X"D9",X"BC",X"C5",X"DA",X"02",X"DB",X"C1",
		X"DC",X"02",X"03",X"06",X"82",X"B0",X"B1",X"B2",X"B3",X"B4",X"02",X"DD",X"DE",X"DF",X"B8",X"02",
		X"E0",X"E1",X"E2",X"02",X"E3",X"E4",X"E5",X"02",X"00",X"E6",X"B2",X"E7",X"E8",X"02",X"00",X"E9",
		X"EA",X"EB",X"EC",X"02",X"00",X"ED",X"EE",X"EF",X"B4",X"02",X"00",X"F0",X"F1",X"F2",X"02",X"F3",
		X"F4",X"F5",X"BF",X"02",X"F7",X"F8",X"F9",X"B0",X"FA",X"02",X"00",X"B2",X"B3",X"FB",X"FC",X"02",
		X"00",X"FD",X"B8",X"02",X"00",X"FE",X"BC",X"CE",X"CF",X"02",X"00",X"D0",X"D1",X"D2",X"CA",X"02",
		X"00",X"D3",X"D4",X"D5",X"C2",X"02",X"00",X"D6",X"D7",X"BC",X"BD",X"02",X"C5",X"BF",X"C0",X"FF",
		X"EC",X"02",X"C3",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"19",X"2F",X"08",X"02",X"18",X"2F",X"08",X"02",X"15",X"38",X"0D",X"04",X"15",X"38",X"0D",X"04",
		X"15",X"42",X"10",X"04",X"15",X"33",X"10",X"00",X"01",X"00",X"0E",X"04",X"09",X"00",X"24",X"04",
		X"0D",X"00",X"24",X"04",X"11",X"01",X"08",X"06",X"17",X"01",X"08",X"06",X"1D",X"01",X"08",X"06",
		X"23",X"01",X"0A",X"02",X"25",X"01",X"0A",X"02",X"27",X"01",X"0C",X"01",X"28",X"01",X"1C",X"01",
		X"29",X"01",X"1C",X"01",X"2A",X"01",X"1C",X"01",X"2B",X"01",X"1C",X"01",X"2C",X"01",X"1C",X"01",
		X"2D",X"04",X"00",X"01",X"2E",X"04",X"00",X"01",X"2F",X"04",X"00",X"01",X"30",X"04",X"00",X"01",
		X"31",X"04",X"00",X"01",X"31",X"84",X"00",X"01",X"31",X"C4",X"00",X"01",X"31",X"44",X"00",X"01",
		X"32",X"04",X"00",X"01",X"33",X"04",X"00",X"01",X"34",X"04",X"00",X"01",X"33",X"C4",X"00",X"01",
		X"34",X"C4",X"00",X"01",X"36",X"04",X"00",X"01",X"36",X"84",X"00",X"01",X"37",X"04",X"00",X"01",
		X"36",X"C4",X"00",X"01",X"36",X"44",X"00",X"01",X"37",X"C4",X"00",X"01",X"38",X"09",X"00",X"01",
		X"39",X"00",X"00",X"01",X"3A",X"09",X"02",X"02",X"05",X"00",X"2C",X"01",X"3D",X"0A",X"28",X"01",
		X"3E",X"01",X"00",X"01",X"3F",X"01",X"00",X"01",X"40",X"01",X"00",X"01",X"41",X"01",X"00",X"01",
		X"42",X"07",X"1A",X"80",X"45",X"07",X"1A",X"80",X"46",X"07",X"1A",X"80",X"47",X"07",X"1A",X"80",
		X"47",X"47",X"1A",X"80",X"46",X"47",X"1A",X"80",X"45",X"47",X"1A",X"80",X"43",X"07",X"1A",X"01",
		X"44",X"07",X"1A",X"01",X"43",X"87",X"1A",X"01",X"44",X"47",X"1A",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"48",X"01",X"1A",X"80",X"49",X"01",X"1A",X"80",X"4A",X"01",X"1A",X"80",
		X"35",X"0A",X"2A",X"80",X"4B",X"01",X"1A",X"80",X"4C",X"01",X"1A",X"80",X"4D",X"01",X"1A",X"80",
		X"4E",X"01",X"00",X"C0",X"4F",X"01",X"10",X"C0",X"53",X"01",X"10",X"C0",X"57",X"01",X"10",X"C0",
		X"5B",X"01",X"12",X"C0",X"61",X"03",X"1E",X"C0",X"62",X"03",X"1E",X"C0",X"63",X"03",X"1E",X"C0",
		X"64",X"03",X"14",X"C0",X"68",X"03",X"14",X"C0",X"6C",X"03",X"16",X"C0",X"6E",X"03",X"16",X"C0",
		X"78",X"08",X"22",X"02",X"70",X"02",X"04",X"04",X"73",X"02",X"06",X"04",X"74",X"02",X"18",X"04",
		X"75",X"02",X"20",X"04",X"7A",X"01",X"1A",X"80",X"4B",X"41",X"1A",X"80",X"4C",X"41",X"1A",X"80",
		X"7B",X"09",X"26",X"02",X"07",X"00",X"2C",X"01",X"7D",X"0E",X"2E",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A3");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
