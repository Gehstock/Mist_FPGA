library IEEE;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

entity rom_crt is
	port (
		clk: in std_logic;
		addr: in std_logic_vector(12 downto 0);
		data: out std_logic_vector(7 downto 0)
	);
end entity;

architecture Behavioral of rom_crt is
	type romDef is array(0 to 8191) of std_logic_vector(7 downto 0);
	constant romData: romDef := (
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"08", x"08", x"08", x"08", x"08", x"00", x"08", x"00",
x"14", x"14", x"00", x"00", x"00", x"00", x"00", x"00",
x"28", x"28", x"7C", x"28", x"7C", x"28", x"28", x"00",
x"10", x"78", x"14", x"38", x"50", x"3C", x"10", x"00",
x"46", x"26", x"10", x"08", x"64", x"62", x"00", x"00",
x"08", x"14", x"14", x"0C", x"52", x"22", x"5C", x"00",
x"20", x"10", x"08", x"00", x"00", x"00", x"00", x"00",
x"20", x"10", x"08", x"08", x"08", x"10", x"20", x"00",
x"04", x"08", x"10", x"10", x"10", x"08", x"04", x"00",
x"00", x"10", x"54", x"38", x"54", x"10", x"00", x"00",
x"00", x"10", x"10", x"7C", x"10", x"10", x"00", x"00",
x"00", x"00", x"00", x"00", x"18", x"18", x"04", x"00",
x"00", x"00", x"00", x"7C", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"18", x"18", x"00", x"00",
x"00", x"40", x"20", x"10", x"08", x"04", x"00", x"00",
x"38", x"44", x"64", x"54", x"4C", x"44", x"38", x"00",
x"10", x"18", x"10", x"10", x"10", x"10", x"38", x"00",
x"38", x"44", x"40", x"20", x"18", x"04", x"7C", x"00",
x"7C", x"20", x"10", x"20", x"40", x"44", x"38", x"00",
x"20", x"30", x"28", x"24", x"7C", x"20", x"20", x"00",
x"7C", x"04", x"3C", x"40", x"40", x"44", x"38", x"00",
x"30", x"08", x"04", x"3C", x"44", x"44", x"38", x"00",
x"7C", x"40", x"20", x"10", x"08", x"08", x"08", x"00",
x"38", x"44", x"44", x"38", x"44", x"44", x"38", x"00",
x"38", x"44", x"44", x"78", x"40", x"20", x"18", x"00",
x"00", x"18", x"18", x"00", x"18", x"18", x"00", x"00",
x"00", x"18", x"18", x"00", x"18", x"18", x"04", x"00",
x"20", x"10", x"08", x"04", x"08", x"10", x"20", x"00",
x"00", x"00", x"7C", x"00", x"7C", x"00", x"00", x"00",
x"04", x"08", x"10", x"20", x"10", x"08", x"04", x"00",
x"1C", x"22", x"20", x"18", x"08", x"00", x"08", x"00",
x"38", x"44", x"74", x"54", x"74", x"04", x"78", x"00",
x"38", x"44", x"44", x"7C", x"44", x"44", x"44", x"00",
x"3C", x"48", x"48", x"38", x"48", x"48", x"3C", x"00",
x"38", x"44", x"04", x"04", x"04", x"44", x"38", x"00",
x"3C", x"48", x"48", x"48", x"48", x"48", x"3C", x"00",
x"7C", x"04", x"04", x"1C", x"04", x"04", x"7C", x"00",
x"7C", x"04", x"04", x"1C", x"04", x"04", x"04", x"00",
x"38", x"44", x"04", x"04", x"74", x"44", x"78", x"00",
x"44", x"44", x"44", x"7C", x"44", x"44", x"44", x"00",
x"38", x"10", x"10", x"10", x"10", x"10", x"38", x"00",
x"70", x"20", x"20", x"20", x"20", x"24", x"18", x"00",
x"44", x"24", x"14", x"0C", x"14", x"24", x"44", x"00",
x"04", x"04", x"04", x"04", x"04", x"04", x"7C", x"00",
x"44", x"6C", x"54", x"54", x"44", x"44", x"44", x"00",
x"44", x"44", x"4C", x"54", x"64", x"44", x"44", x"00",
x"38", x"44", x"44", x"44", x"44", x"44", x"38", x"00",
x"3C", x"44", x"44", x"3C", x"04", x"04", x"04", x"00",
x"38", x"44", x"44", x"44", x"54", x"24", x"58", x"00",
x"3C", x"44", x"44", x"3C", x"14", x"24", x"44", x"00",
x"38", x"44", x"08", x"10", x"20", x"44", x"38", x"00",
x"7C", x"10", x"10", x"10", x"10", x"10", x"10", x"00",
x"44", x"44", x"44", x"44", x"44", x"44", x"38", x"00",
x"44", x"44", x"44", x"44", x"44", x"28", x"10", x"00",
x"44", x"44", x"44", x"54", x"54", x"54", x"28", x"00",
x"44", x"44", x"28", x"10", x"28", x"44", x"44", x"00",
x"44", x"44", x"44", x"28", x"10", x"10", x"10", x"00",
x"7C", x"40", x"20", x"10", x"08", x"04", x"7C", x"00",
x"28", x"38", x"44", x"04", x"04", x"44", x"38", x"00",
x"20", x"38", x"44", x"04", x"04", x"44", x"38", x"00",
x"3C", x"48", x"48", x"5C", x"48", x"48", x"3C", x"00",
x"28", x"38", x"44", x"08", x"30", x"44", x"38", x"00",
x"28", x"7C", x"40", x"20", x"10", x"08", x"7C", x"00",
x"10", x"28", x"44", x"00", x"00", x"00", x"00", x"00",
x"00", x"18", x"20", x"38", x"24", x"38", x"00", x"00",
x"04", x"04", x"1C", x"24", x"24", x"1C", x"00", x"00",
x"00", x"38", x"04", x"04", x"04", x"38", x"00", x"00",
x"20", x"20", x"38", x"24", x"24", x"38", x"00", x"00",
x"00", x"18", x"24", x"1C", x"04", x"18", x"00", x"00",
x"10", x"28", x"08", x"1C", x"08", x"08", x"08", x"00",
x"00", x"38", x"24", x"24", x"38", x"20", x"18", x"00",
x"04", x"04", x"1C", x"24", x"24", x"24", x"00", x"00",
x"10", x"00", x"18", x"10", x"10", x"38", x"00", x"00",
x"10", x"00", x"18", x"10", x"10", x"14", x"08", x"00",
x"04", x"04", x"14", x"0C", x"14", x"24", x"00", x"00",
x"18", x"10", x"10", x"10", x"10", x"38", x"00", x"00",
x"00", x"2C", x"54", x"54", x"54", x"54", x"00", x"00",
x"00", x"1C", x"24", x"24", x"24", x"24", x"00", x"00",
x"00", x"18", x"24", x"24", x"24", x"18", x"00", x"00",
x"00", x"1C", x"24", x"24", x"1C", x"04", x"04", x"00",
x"00", x"1C", x"12", x"12", x"1C", x"10", x"78", x"00",
x"00", x"34", x"0C", x"04", x"04", x"04", x"00", x"00",
x"00", x"38", x"04", x"18", x"20", x"1C", x"00", x"00",
x"10", x"38", x"10", x"10", x"10", x"20", x"00", x"00",
x"00", x"24", x"24", x"24", x"24", x"38", x"00", x"00",
x"00", x"44", x"44", x"44", x"28", x"10", x"00", x"00",
x"00", x"44", x"44", x"54", x"54", x"28", x"00", x"00",
x"00", x"44", x"28", x"10", x"28", x"44", x"00", x"00",
x"00", x"24", x"24", x"24", x"38", x"20", x"18", x"00",
x"00", x"3C", x"20", x"10", x"08", x"3C", x"00", x"00",
x"38", x"00", x"38", x"04", x"04", x"38", x"00", x"00",
x"20", x"00", x"38", x"04", x"04", x"38", x"00", x"00",
x"20", x"70", x"20", x"38", x"24", x"38", x"00", x"00",
x"28", x"38", x"04", x"18", x"20", x"1C", x"00", x"00",
x"38", x"00", x"3C", x"10", x"08", x"3C", x"00", x"00",
x"09", x"0A", x"0B", x"1F", x"14", x"13", x"12", x"11",
x"36", x"74", x"7A", x"72", x"37", x"75", x"69", x"6F",
x"31", x"77", x"71", x"65", x"6D", x"6B", x"6A", x"6C",
x"79", x"73", x"61", x"64", x"6E", x"67", x"68", x"66",
x"3A", x"7F", x"7C", x"7B", x"3B", x"7E", x"7D", x"70",
x"00", x"0D", x"00", x"20", x"34", x"35", x"39", x"38",
x"33", x"32", x"2E", x"2C", x"63", x"78", x"76", x"62",
x"60", x"2F", x"30", x"2D", x"87", x"FC", x"87", x"FA",
x"87", x"F6", x"87", x"EE", x"87", x"DE", x"87", x"BE",
x"87", x"7E", x"86", x"FE", x"85", x"FE", x"83", x"FE",
x"85", x"FC", x"8A", x"48", x"98", x"48", x"A5", x"FC",
x"A8", x"2A", x"2A", x"2A", x"2A", x"29", x"03", x"AA",
x"BD", x"00", x"02", x"D0", x"05", x"BD", x"04", x"02",
x"F0", x"24", x"85", x"F1", x"98", x"0A", x"0A", x"0A",
x"85", x"F0", x"A0", x"07", x"B1", x"F0", x"84", x"FA",
x"A4", x"E9", x"20", x"C1", x"EE", x"EA", x"EA", x"EA",
x"91", x"E6", x"A5", x"E6", x"38", x"E9", x"20", x"85",
x"E6", x"A4", x"FA", x"88", x"10", x"E6", x"68", x"A8",
x"68", x"AA", x"A5", x"FC", x"60", x"A6", x"EA", x"86",
x"E8", x"A4", x"EC", x"84", x"E9", x"A9", x"E0", x"85",
x"E6", x"A5", x"E8", x"4C", x"9E", x"EE", x"EA", x"EA",
x"EA", x"60", x"A6", x"EB", x"18", x"90", x"05", x"20",
x"95", x"E3", x"A4", x"EC", x"20", x"AD", x"E4", x"C4",
x"ED", x"C8", x"90", x"F8", x"E4", x"EB", x"B0", x"15",
x"E8", x"E6", x"E7", x"90", x"ED", x"C6", x"E9", x"C4",
x"EC", x"D0", x"0D", x"A4", x"ED", x"84", x"E9", x"E4",
x"EA", x"F0", x"05", x"C6", x"E8", x"20", x"9D", x"E3",
x"68", x"A8", x"68", x"AA", x"A5", x"FC", x"60", x"85",
x"FC", x"8A", x"48", x"98", x"48", x"A5", x"FC", x"A6",
x"E8", x"A4", x"E9", x"C9", x"20", x"B0", x"39", x"2C",
x"08", x"02", x"30", x"34", x"C9", x"05", x"F0", x"B2",
x"C9", x"0C", x"F0", x"B3", x"C9", x"06", x"F0", x"B4",
x"C9", x"08", x"F0", x"C1", x"C9", x"0B", x"F0", x"C7",
x"C9", x"09", x"F0", x"1F", x"C9", x"0A", x"F0", x"25",
x"C9", x"0D", x"F0", x"6A", x"C9", x"04", x"D0", x"06",
x"20", x"95", x"E3", x"4C", x"D8", x"E3", x"C9", x"07",
x"D0", x"B6", x"20", x"F4", x"E4", x"4C", x"D8", x"E3",
x"20", x"50", x"E3", x"E6", x"E9", x"C4", x"ED", x"90",
x"A7", x"A4", x"EC", x"84", x"E9", x"E6", x"E8", x"E4",
x"EB", x"90", x"9A", x"C6", x"E8", x"A5", x"EA", x"20",
x"A3", x"E3", x"A5", x"E6", x"18", x"90", x"13", x"E6",
x"E7", x"A4", x"EC", x"B1", x"E6", x"91", x"EE", x"C4",
x"ED", x"C8", x"90", x"F7", x"A5", x"E6", x"E9", x"20",
x"85", x"E6", x"85", x"EE", x"B0", x"EB", x"A5", x"E7",
x"85", x"EF", x"38", x"E9", x"60", x"C5", x"EB", x"90",
x"DE", x"2C", x"43", x"02", x"10", x"03", x"20", x"4E",
x"F0", x"4C", x"B2", x"E3", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"4C", x"9F",
x"E4", x"F0", x"1C", x"A0", x"09", x"88", x"F0", x"17",
x"A2", x"FF", x"20", x"E3", x"E4", x"20", x"0F", x"E6",
x"D0", x"F3", x"A4", x"E9", x"20", x"C2", x"E4", x"20",
x"0F", x"E6", x"F0", x"FB", x"20", x"C2", x"E4", x"A6",
x"E8", x"AD", x"09", x"02", x"D0", x"8B", x"A4", x"EC",
x"84", x"E9", x"4C", x"D8", x"E3", x"86", x"FB", x"A2",
x"08", x"A9", x"00", x"91", x"E6", x"A5", x"E6", x"38",
x"E9", x"20", x"85", x"E6", x"CA", x"D0", x"F2", x"A6",
x"FB", x"60", x"86", x"FB", x"A2", x"08", x"B1", x"E6",
x"49", x"FF", x"91", x"E6", x"A5", x"E6", x"38", x"E9",
x"20", x"85", x"E6", x"CA", x"D0", x"F0", x"A6", x"FB",
x"60", x"48", x"98", x"A0", x"BB", x"88", x"D0", x"FD",
x"A8", x"68", x"60", x"20", x"D9", x"E4", x"CA", x"D0",
x"FA", x"60", x"8E", x"00", x"88", x"20", x"D9", x"E4",
x"CA", x"D0", x"F7", x"60", x"48", x"8A", x"A2", x"70",
x"20", x"EA", x"E4", x"AA", x"68", x"60", x"FF", x"FF",
x"8A", x"48", x"98", x"48", x"20", x"42", x"F0", x"8D",
x"42", x"02", x"20", x"42", x"F0", x"49", x"FF", x"91",
x"E6", x"A0", x"00", x"88", x"F0", x"F4", x"20", x"B0",
x"E5", x"90", x"3E", x"85", x"FC", x"F0", x"3A", x"A2",
x"0A", x"20", x"E3", x"E4", x"20", x"B0", x"E5", x"90",
x"30", x"C5", x"FC", x"D0", x"2C", x"A4", x"E9", x"AD",
x"42", x"02", x"91", x"E6", x"AD", x"0C", x"02", x"D0",
x"06", x"38", x"6E", x"0C", x"02", x"90", x"23", x"2C",
x"0C", x"02", x"10", x"0E", x"A9", x"40", x"8D", x"0C",
x"02", x"A0", x"30", x"20", x"3F", x"F0", x"90", x"09",
x"B0", x"10", x"A0", x"08", x"20", x"3F", x"F0", x"B0",
x"09", x"A9", x"00", x"8D", x"0C", x"02", x"4C", x"13",
x"E5", x"EA", x"AD", x"FB", x"87", x"29", x"20", x"0A",
x"85", x"FA", x"AD", x"FD", x"87", x"29", x"20", x"05",
x"FA", x"0A", x"85", x"FA", x"A5", x"FC", x"C9", x"21",
x"90", x"2D", x"C9", x"60", x"B0", x"0F", x"2C", x"0E",
x"02", x"10", x"02", x"EA", x"EA", x"A4", x"FA", x"30",
x"1E", x"49", x"10", x"D0", x"1A", x"F0", x"05", x"2C",
x"0D", x"02", x"10", x"04", x"A4", x"FA", x"30", x"02",
x"49", x"20", x"EA", x"EA", x"EA", x"EA", x"EA", x"EA",
x"EA", x"24", x"FA", x"70", x"02", x"29", x"1F", x"85",
x"FC", x"68", x"A8", x"68", x"AA", x"A5", x"FC", x"60",
x"8A", x"48", x"98", x"48", x"A2", x"14", x"CA", x"CA",
x"30", x"2D", x"BD", x"3C", x"E3", x"85", x"F1", x"BD",
x"3D", x"E3", x"85", x"F0", x"20", x"F9", x"E5", x"90",
x"ED", x"C0", x"00", x"D0", x"21", x"0A", x"B0", x"09",
x"C8", x"0A", x"B0", x"05", x"C8", x"0A", x"B0", x"01",
x"C8", x"8A", x"0A", x"84", x"FA", x"18", x"65", x"FA",
x"AA", x"BD", x"00", x"E3", x"85", x"FA", x"38", x"68",
x"A8", x"68", x"AA", x"A5", x"FA", x"60", x"29", x"10",
x"D0", x"01", x"88", x"8A", x"18", x"69", x"28", x"D0",
x"E2", x"38", x"A0", x"00", x"B1", x"F0", x"09", x"0F",
x"49", x"FF", x"D0", x"0A", x"C8", x"B1", x"F0", x"09",
x"CF", x"49", x"FF", x"D0", x"01", x"18", x"60", x"AD",
x"00", x"80", x"09", x"0F", x"49", x"FF", x"D0", x"07",
x"AD", x"01", x"80", x"09", x"CF", x"49", x"FF", x"60",
x"4C", x"2D", x"F0", x"C9", x"57", x"D0", x"03", x"4C",
x"03", x"C0", x"C9", x"43", x"D0", x"03", x"4C", x"00",
x"C0", x"60", x"E8", x"BD", x"80", x"02", x"C9", x"20",
x"F0", x"F8", x"60", x"85", x"F3", x"84", x"F2", x"98",
x"48", x"A0", x"00", x"B1", x"F2", x"C9", x"04", x"F0",
x"0B", x"20", x"F1", x"FF", x"E6", x"F2", x"D0", x"F3",
x"E6", x"F3", x"D0", x"EF", x"68", x"A8", x"60", x"A2",
x"00", x"8A", x"F0", x"01", x"CA", x"20", x"EE", x"FF",
x"9D", x"80", x"02", x"C9", x"0D", x"F0", x"1B", x"C9",
x"08", x"F0", x"EE", x"C9", x"18", x"F0", x"0D", x"C9",
x"20", x"90", x"EA", x"E8", x"10", x"E7", x"20", x"F4",
x"E4", x"38", x"B0", x"E0", x"A9", x"0D", x"A2", x"00",
x"F0", x"DE", x"60", x"FF", x"0D", x"0A", x"00", x"00",
x"00", x"00", x"2A", x"04", x"E0", x"2F", x"00", x"00",
x"00", x"00", x"E0", x"60", x"00", x"00", x"00", x"1F",
x"00", x"1F", x"E0", x"20", x"00", x"00", x"00", x"00",
x"00", x"E0", x"E1", x"E2", x"00", x"00", x"00", x"00",
x"FF", x"00", x"00", x"00", x"00", x"FF", x"FD", x"53",
x"FF", x"FF", x"1C", x"E7", x"62", x"E7", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"20", x"E6", x"FD", x"E8", x"06", x"E9", x"0E", x"E9",
x"D0", x"EA", x"09", x"EB", x"48", x"EB", x"6A", x"EB",
x"AB", x"EB", x"80", x"EC", x"D0", x"EE", x"57", x"EF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"42", x"4A", x"55", x"45", x"43", x"51", x"46", x"4D",
x"41", x"58", x"48", x"23", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"20", x"00", x"E5", x"C9",
x"11", x"D0", x"0B", x"AD", x"0D", x"02", x"49", x"FF",
x"8D", x"0D", x"02", x"6C", x"16", x"02", x"C9", x"12",
x"D0", x"0B", x"AD", x"10", x"02", x"49", x"FF", x"8D",
x"10", x"02", x"6C", x"16", x"02", x"C9", x"13", x"D0",
x"0B", x"AD", x"0E", x"02", x"49", x"FF", x"8D", x"0E",
x"02", x"6C", x"16", x"02", x"4C", x"45", x"F0", x"EA",
x"2C", x"0F", x"02", x"30", x"03", x"20", x"F1", x"FF",
x"60", x"48", x"8A", x"2C", x"00", x"80", x"10", x"FB",
x"30", x"0A", x"20", x"DF", x"E3", x"2C", x"10", x"02",
x"10", x"EE", x"30", x"ED", x"48", x"98", x"48", x"BA",
x"BD", x"03", x"01", x"A2", x"09", x"18", x"2A", x"6A",
x"B0", x"05", x"8D", x"00", x"98", x"90", x"07", x"29",
x"FF", x"30", x"03", x"8D", x"00", x"90", x"AC", x"13",
x"02", x"20", x"B8", x"E7", x"CA", x"30", x"06", x"D0",
x"E6", x"09", x"01", x"D0", x"E2", x"68", x"A8", x"68",
x"AA", x"68", x"60", x"FF", x"FF", x"FF", x"FF", x"A0",
x"00", x"8C", x"00", x"98", x"8C", x"00", x"90", x"2C",
x"FF", x"87", x"10", x"03", x"C8", x"D0", x"F8", x"88",
x"84", x"F4", x"60", x"AE", x"2A", x"0A", x"04", x"EA",
x"EA", x"EA", x"EA", x"EA", x"EA", x"EA", x"88", x"D0",
x"F6", x"60", x"FF", x"48", x"10", x"05", x"38", x"90",
x"02", x"49", x"80", x"0A", x"D0", x"F9", x"68", x"60",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"48", x"A9", x"20", x"20",
x"F1", x"FF", x"68", x"60", x"A2", x"03", x"20", x"DC",
x"E7", x"CA", x"D0", x"FA", x"60", x"C9", x"0A", x"90",
x"02", x"69", x"06", x"69", x"30", x"60", x"A9", x"0D",
x"20", x"F1", x"FF", x"A9", x"0A", x"4C", x"F1", x"FF",
x"20", x"DC", x"E7", x"48", x"4A", x"4A", x"4A", x"4A",
x"20", x"ED", x"E7", x"20", x"F1", x"FF", x"68", x"29",
x"0F", x"20", x"ED", x"E7", x"4C", x"F1", x"FF", x"20",
x"DC", x"E7", x"A5", x"FF", x"20", x"03", x"E8", x"A5",
x"FE", x"4C", x"03", x"E8", x"20", x"33", x"E6", x"BD",
x"80", x"02", x"E8", x"C9", x"30", x"90", x"0F", x"E9",
x"30", x"C9", x"0A", x"90", x"0A", x"C9", x"11", x"90",
x"05", x"E9", x"07", x"C9", x"10", x"60", x"38", x"60",
x"20", x"27", x"E8", x"90", x"06", x"60", x"20", x"24",
x"E8", x"B0", x"0F", x"0A", x"0A", x"0A", x"0A", x"85",
x"FC", x"20", x"27", x"E8", x"B0", x"04", x"05", x"FC",
x"85", x"FC", x"60", x"20", x"46", x"E8", x"B0", x"07",
x"85", x"F7", x"20", x"40", x"E8", x"85", x"F6", x"60",
x"20", x"7D", x"E8", x"B0", x"1D", x"20", x"92", x"E8",
x"B0", x"18", x"4C", x"5B", x"E8", x"20", x"7D", x"E8",
x"B0", x"10", x"4C", x"5B", x"E8", x"20", x"5B", x"E8",
x"B0", x"08", x"A5", x"F6", x"85", x"FE", x"A5", x"F7",
x"85", x"FF", x"60", x"E6", x"FE", x"D0", x"02", x"E6",
x"FF", x"60", x"20", x"5B", x"E8", x"B0", x"08", x"A5",
x"F6", x"85", x"F4", x"A5", x"F7", x"85", x"F5", x"60",
x"E6", x"F4", x"D0", x"02", x"E6", x"F5", x"60", x"18",
x"A5", x"FE", x"65", x"F6", x"85", x"FE", x"A5", x"FF",
x"65", x"F7", x"85", x"FF", x"60", x"38", x"A5", x"FE",
x"E5", x"F4", x"85", x"FE", x"A5", x"FF", x"E5", x"F5",
x"85", x"FF", x"60", x"38", x"A5", x"F6", x"E5", x"F4",
x"A5", x"F7", x"E5", x"F5", x"60", x"38", x"A5", x"FE",
x"E5", x"F4", x"A5", x"FF", x"E5", x"F5", x"60", x"18",
x"A5", x"F6", x"E9", x"00", x"85", x"F6", x"A5", x"F7",
x"E9", x"00", x"85", x"F7", x"60", x"18", x"A5", x"FE",
x"E9", x"00", x"85", x"FE", x"A5", x"FF", x"E9", x"00",
x"85", x"FF", x"60", x"38", x"A5", x"FE", x"E5", x"F6",
x"A5", x"FF", x"E5", x"F7", x"60", x"20", x"5B", x"E8",
x"B0", x"2C", x"68", x"68", x"90", x"05", x"20", x"5B",
x"E8", x"B0", x"23", x"6C", x"F6", x"00", x"20", x"75",
x"E8", x"B0", x"1B", x"A0", x"00", x"20", x"F6", x"E7",
x"20", x"17", x"E8", x"A2", x"09", x"CA", x"F0", x"F5",
x"B1", x"FE", x"20", x"00", x"E8", x"20", x"F3", x"E8",
x"20", x"8B", x"E8", x"90", x"F0", x"18", x"60", x"FF",
x"00", x"90", x"6D", x"65", x"69", x"7D", x"79", x"61",
x"71", x"75", x"D0", x"2D", x"25", x"29", x"3D", x"39",
x"21", x"31", x"35", x"30", x"0A", x"0E", x"06", x"1E",
x"16", x"08", x"90", x"08", x"B0", x"88", x"F0", x"48",
x"2C", x"24", x"C8", x"30", x"C8", x"D0", x"28", x"10",
x"28", x"00", x"A8", x"50", x"A8", x"70", x"D8", x"18",
x"D8", x"D8", x"D8", x"58", x"D8", x"B8", x"D8", x"CD",
x"C5", x"C9", x"DD", x"D9", x"C1", x"D1", x"D5", x"38",
x"EC", x"E4", x"E0", x"38", x"CC", x"C4", x"C0", x"84",
x"CE", x"C6", x"DE", x"D6", x"84", x"CA", x"84", x"88",
x"D4", x"4D", x"45", x"49", x"5D", x"59", x"41", x"51",
x"55", x"D2", x"EE", x"E6", x"FE", x"F6", x"D2", x"E8",
x"D2", x"C8", x"CA", x"4C", x"6C", x"2A", x"20", x"86",
x"AD", x"A5", x"A9", x"BD", x"B9", x"A1", x"B1", x"B5",
x"86", x"AE", x"A6", x"A2", x"BE", x"B6", x"86", x"AC",
x"A4", x"A0", x"BC", x"B4", x"26", x"4A", x"4E", x"46",
x"5E", x"56", x"CE", x"EA", x"3E", x"0D", x"05", x"09",
x"1D", x"19", x"01", x"11", x"15", x"41", x"48", x"41",
x"08", x"C1", x"68", x"C1", x"28", x"C9", x"2A", x"2E",
x"26", x"3E", x"36", x"C9", x"6A", x"6E", x"66", x"7E",
x"76", x"A9", x"40", x"A9", x"60", x"19", x"ED", x"E5",
x"E9", x"FD", x"F9", x"E1", x"F1", x"F5", x"99", x"38",
x"99", x"F8", x"99", x"78", x"B9", x"8D", x"85", x"9D",
x"99", x"81", x"91", x"95", x"B9", x"8E", x"86", x"96",
x"B9", x"8C", x"84", x"94", x"05", x"AA", x"05", x"A8",
x"25", x"BA", x"65", x"8A", x"65", x"9A", x"65", x"98",
x"00", x"60", x"82", x"81", x"C1", x"8A", x"86", x"99",
x"95", x"89", x"11", x"82", x"81", x"C1", x"8A", x"86",
x"99", x"95", x"89", x"1B", x"80", x"82", x"81", x"8A",
x"89", x"63", x"A1", x"67", x"A1", x"46", x"A1", x"16",
x"82", x"81", x"4A", x"A1", x"51", x"A1", x"18", x"A1",
x"69", x"80", x"61", x"A1", x"65", x"A1", x"60", x"80",
x"10", x"80", x"48", x"80", x"34", x"80", x"06", x"82",
x"81", x"C1", x"8A", x"86", x"99", x"95", x"89", x"0C",
x"82", x"81", x"C1", x"4C", x"82", x"81", x"C1", x"62",
x"82", x"81", x"8A", x"89", x"0E", x"80", x"4E", x"80",
x"27", x"82", x"81", x"C1", x"8A", x"86", x"99", x"95",
x"89", x"61", x"82", x"81", x"8A", x"89", x"0D", x"80",
x"4D", x"80", x"06", x"82", x"92", x"27", x"82", x"40",
x"82", x"81", x"C1", x"8A", x"86", x"99", x"95", x"89",
x"0C", x"82", x"81", x"C1", x"86", x"85", x"4C", x"82",
x"81", x"C1", x"8A", x"89", x"27", x"80", x"82", x"81",
x"8A", x"89", x"07", x"80", x"41", x"82", x"81", x"C1",
x"8A", x"86", x"99", x"95", x"89", x"40", x"80", x"04",
x"80", x"40", x"80", x"04", x"80", x"1B", x"80", x"82",
x"81", x"8A", x"89", x"27", x"80", x"82", x"81", x"8A",
x"89", x"48", x"80", x"64", x"80", x"61", x"82", x"81",
x"C1", x"8A", x"86", x"99", x"95", x"89", x"62", x"80",
x"12", x"80", x"4A", x"80", x"40", x"82", x"81", x"8A",
x"86", x"99", x"95", x"89", x"0C", x"82", x"81", x"85",
x"4C", x"82", x"81", x"89", x"0E", x"80", x"4E", x"80",
x"0F", x"80", x"40", x"80", x"64", x"80", x"42", x"80",
x"20", x"75", x"E8", x"B0", x"33", x"A2", x"00", x"86",
x"F4", x"86", x"F5", x"A0", x"00", x"8A", x"71", x"FE",
x"AA", x"90", x"06", x"E6", x"F4", x"D0", x"02", x"E6",
x"F5", x"20", x"F3", x"E8", x"20", x"8B", x"E8", x"90",
x"EC", x"20", x"F6", x"E7", x"A9", x"3D", x"20", x"F1",
x"FF", x"A5", x"F5", x"20", x"00", x"E8", x"A5", x"F4",
x"20", x"00", x"E8", x"8A", x"20", x"00", x"E8", x"18",
x"60", x"20", x"68", x"E8", x"B0", x"25", x"20", x"C3",
x"E8", x"90", x"33", x"A0", x"00", x"20", x"CD", x"E8",
x"90", x"1A", x"20", x"B5", x"E8", x"20", x"A7", x"E8",
x"B0", x"11", x"B1", x"F6", x"91", x"FE", x"20", x"D7",
x"E8", x"90", x"08", x"20", x"E5", x"E8", x"20", x"C3",
x"E8", x"B0", x"EF", x"60", x"B1", x"F4", x"91", x"FE",
x"20", x"A0", x"E8", x"F0", x"F6", x"20", x"8B", x"E8",
x"20", x"C3", x"E8", x"B0", x"EF", x"60", x"38", x"60",
x"20", x"75", x"E8", x"B0", x"1C", x"A0", x"00", x"20",
x"46", x"E8", x"90", x"09", x"C9", x"27", x"D0", x"EE",
x"BD", x"80", x"02", x"AA", x"8A", x"91", x"FE", x"AA",
x"20", x"F3", x"E8", x"20", x"8B", x"E8", x"90", x"F4",
x"18", x"60", x"20", x"7D", x"E8", x"A0", x"00", x"F0",
x"0D", x"BD", x"80", x"02", x"91", x"FE", x"D1", x"FE",
x"38", x"D0", x"2F", x"20", x"8B", x"E8", x"20", x"F6",
x"E7", x"20", x"17", x"E8", x"B1", x"FE", x"20", x"00",
x"E8", x"20", x"DC", x"E7", x"20", x"57", x"E6", x"A2",
x"00", x"20", x"46", x"E8", x"90", x"DE", x"C9", x"0D",
x"F0", x"E1", x"C9", x"27", x"F0", x"D3", x"C9", x"2D",
x"18", x"D0", x"07", x"20", x"E5", x"E8", x"18", x"90",
x"D5", x"18", x"60", x"20", x"7D", x"E8", x"20", x"F6",
x"E7", x"20", x"17", x"E8", x"20", x"57", x"E6", x"A2",
x"00", x"20", x"33", x"E6", x"20", x"C2", x"EB", x"90",
x"ED", x"60", x"A9", x"FD", x"85", x"FC", x"A0", x"04",
x"BD", x"80", x"02", x"E8", x"0A", x"0A", x"0A", x"0A",
x"66", x"F5", x"66", x"F4", x"88", x"10", x"F8", x"E6",
x"FC", x"30", x"EB", x"F0", x"F2", x"20", x"33", x"E6",
x"A9", x"80", x"D0", x"02", x"05", x"F8", x"85", x"F8",
x"20", x"40", x"E8", x"90", x"18", x"C9", x"23", x"D0",
x"04", x"A9", x"40", x"D0", x"EF", x"C9", x"28", x"D0",
x"04", x"A9", x"10", x"D0", x"E7", x"C9", x"27", x"D0",
x"30", x"BD", x"80", x"02", x"E8", x"85", x"E4", x"E6",
x"F8", x"20", x"40", x"E8", x"B0", x"07", x"85", x"E5",
x"E6", x"F8", x"20", x"40", x"E8", x"C9", x"21", x"D0",
x"08", x"A9", x"08", x"05", x"F8", x"85", x"F8", x"D0",
x"10", x"C9", x"22", x"D0", x"04", x"A9", x"04", x"D0",
x"F2", x"C9", x"2C", x"F0", x"E5", x"C9", x"29", x"F0",
x"E1", x"A2", x"D0", x"CA", x"F0", x"43", x"BD", x"00",
x"EA", x"30", x"F8", x"C5", x"F5", x"D0", x"F4", x"BD",
x"30", x"E9", x"C5", x"F4", x"D0", x"ED", x"E8", x"BD",
x"00", x"EA", x"10", x"2D", x"C5", x"F8", x"F0", x"10",
x"29", x"20", x"F0", x"F2", x"A5", x"E5", x"38", x"E9",
x"02", x"38", x"E5", x"FE", x"85", x"E4", x"A9", x"01",
x"29", x"03", x"48", x"A0", x"00", x"BD", x"30", x"E9",
x"91", x"FE", x"68", x"AA", x"18", x"20", x"8B", x"E8",
x"CA", x"30", x"07", x"B5", x"E4", x"91", x"FE", x"90",
x"F4", x"38", x"60", x"FF", x"FF", x"FF", x"FF", x"FF",
x"20", x"75", x"E8", x"90", x"14", x"A2", x"0C", x"8A",
x"48", x"20", x"F6", x"E7", x"20", x"A9", x"EC", x"20",
x"8B", x"E8", x"68", x"AA", x"CA", x"D0", x"F0", x"18",
x"60", x"20", x"F6", x"E7", x"20", x"A9", x"EC", x"20",
x"F3", x"E8", x"20", x"8B", x"E8", x"90", x"F2", x"18",
x"60", x"20", x"17", x"E8", x"A0", x"00", x"B1", x"FE",
x"A0", x"80", x"84", x"F8", x"A2", x"D0", x"CA", x"F0",
x"0D", x"DD", x"30", x"E9", x"D0", x"F8", x"BC", x"00",
x"EA", x"10", x"F3", x"84", x"F8", x"CA", x"BD", x"00",
x"EA", x"30", x"FA", x"85", x"F5", x"BD", x"30", x"E9",
x"85", x"F4", x"98", x"29", x"03", x"AA", x"A0", x"FF",
x"C8", x"B1", x"FE", x"20", x"00", x"E8", x"CA", x"10",
x"F7", x"C8", x"20", x"E4", x"E7", x"C0", x"04", x"D0",
x"F8", x"88", x"A2", x"05", x"A9", x"02", x"46", x"F5",
x"66", x"F4", x"2A", x"CA", x"D0", x"F8", x"20", x"F1",
x"FF", x"88", x"D0", x"EE", x"20", x"DC", x"E7", x"A5",
x"F8", x"0A", x"F0", x"A3", x"10", x"04", x"A9", x"23",
x"D0", x"08", x"29", x"20", x"F0", x"02", x"A9", x"08",
x"09", x"20", x"20", x"F1", x"FF", x"A5", x"F8", x"C9",
x"A1", x"D0", x"1D", x"20", x"8B", x"E8", x"B1", x"FE",
x"A8", x"38", x"65", x"FE", x"48", x"A6", x"FF", x"98",
x"10", x"03", x"B0", x"04", x"CA", x"90", x"01", x"E8",
x"8A", x"20", x"03", x"E8", x"68", x"4C", x"03", x"E8",
x"29", x"03", x"A8", x"B1", x"FE", x"20", x"03", x"E8",
x"20", x"8B", x"E8", x"88", x"88", x"F0", x"F4", x"A2",
x"58", x"A5", x"F8", x"29", x"1C", x"F0", x"22", x"0A",
x"0A", x"0A", x"0A", x"F0", x"0B", x"B0", x"04", x"10",
x"0E", x"30", x"0D", x"10", x"07", x"20", x"68", x"ED",
x"A9", x"29", x"D0", x"0A", x"20", x"60", x"ED", x"E8",
x"A9", x"2C", x"20", x"F1", x"FF", x"8A", x"4C", x"F1",
x"FF", x"18", x"60", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"A5", x"7B", x"85", x"FE", x"A5", x"7C", x"85", x"FF",
x"A9", x"00", x"85", x"F4", x"A9", x"04", x"85", x"F5",
x"20", x"B5", x"E8", x"E6", x"FE", x"E6", x"FF", x"A9",
x"60", x"A2", x"00", x"A0", x"14", x"20", x"B7", x"E7",
x"8D", x"00", x"88", x"CA", x"D0", x"F5", x"A8", x"88",
x"98", x"D0", x"F0", x"A0", x"08", x"20", x"DC", x"ED",
x"A5", x"FE", x"20", x"D8", x"ED", x"A5", x"FF", x"20",
x"D8", x"ED", x"20", x"D7", x"ED", x"20", x"D7", x"ED",
x"B1", x"F4", x"A2", x"07", x"A0", x"07", x"20", x"DC",
x"ED", x"E6", x"F4", x"D0", x"02", x"E6", x"F5", x"C6",
x"FE", x"D0", x"EA", x"C6", x"FF", x"D0", x"E9", x"60",
x"A2", x"07", x"A0", x"09", x"20", x"B7", x"E7", x"6A",
x"B0", x"05", x"8D", x"00", x"88", x"90", x"0D", x"A0",
x"0A", x"20", x"B7", x"E7", x"8D", x"00", x"88", x"A0",
x"09", x"20", x"B7", x"E7", x"A0", x"0A", x"20", x"B7",
x"E7", x"8D", x"00", x"88", x"CA", x"10", x"DB", x"60",
x"E8", x"F0", x"05", x"2C", x"FF", x"87", x"70", x"F8",
x"60", x"E8", x"F0", x"05", x"2C", x"FF", x"87", x"50",
x"F8", x"60", x"A0", x"08", x"20", x"1C", x"EE", x"6A",
x"88", x"D0", x"F9", x"60", x"A2", x"00", x"2C", x"FF",
x"87", x"50", x"08", x"20", x"00", x"EE", x"20", x"09",
x"EE", x"70", x"06", x"20", x"09", x"EE", x"20", x"00",
x"EE", x"E0", x"33", x"60", x"A2", x"00", x"2C", x"FF",
x"87", x"50", x"06", x"20", x"00", x"EE", x"E0", x"19",
x"60", x"20", x"09", x"EE", x"E0", x"19", x"60", x"20",
x"34", x"EE", x"90", x"FB", x"E0", x"33", x"B0", x"F7",
x"A0", x"0A", x"20", x"34", x"EE", x"90", x"F0", x"88",
x"D0", x"F8", x"20", x"34", x"EE", x"B0", x"FB", x"20",
x"34", x"EE", x"B0", x"E3", x"60", x"A0", x"FF", x"A9",
x"03", x"84", x"7B", x"85", x"7C", x"20", x"47", x"EE",
x"20", x"12", x"EE", x"85", x"FE", x"20", x"12", x"EE",
x"85", x"FF", x"20", x"12", x"EE", x"E6", x"7B", x"D0",
x"02", x"E6", x"7C", x"91", x"7B", x"C6", x"FE", x"D0",
x"F1", x"C6", x"FF", x"D0", x"ED", x"60", x"C9", x"10",
x"90", x"07", x"29", x"0F", x"09", x"70", x"85", x"E1",
x"60", x"09", x"60", x"85", x"E1", x"60", x"C9", x"10",
x"B0", x"07", x"29", x"0F", x"09", x"60", x"85", x"E7",
x"60", x"29", x"0F", x"09", x"70", x"85", x"E7", x"60",
x"A2", x"23", x"BD", x"9C", x"E6", x"9D", x"00", x"02",
x"CA", x"10", x"F7", x"A9", x"00", x"8D", x"43", x"02",
x"60", x"2C", x"0E", x"02", x"10", x"03", x"49", x"FF",
x"60", x"24", x"FC", x"30", x"F9", x"60", x"FF", x"FF",
x"20", x"75", x"E8", x"90", x"03", x"20", x"49", x"EF",
x"A0", x"00", x"20", x"F6", x"E7", x"20", x"17", x"E8",
x"A2", x"FF", x"E8", x"E0", x"05", x"B0", x"0E", x"B1",
x"FE", x"20", x"00", x"E8", x"20", x"F3", x"E8", x"20",
x"8B", x"E8", x"90", x"EE", x"E8", x"A5", x"FE", x"48",
x"86", x"FE", x"38", x"E5", x"FE", x"85", x"FE", x"A5",
x"FF", x"48", x"E9", x"00", x"85", x"FF", x"20", x"40",
x"EF", x"E8", x"E0", x"06", x"90", x"F8", x"CA", x"F0",
x"1B", x"B1", x"FE", x"C9", x"20", x"90", x"04", x"C9",
x"80", x"90", x"02", x"A9", x"2E", x"20", x"F1", x"FF",
x"20", x"F3", x"E8", x"20", x"8B", x"E8", x"90", x"E6",
x"68", x"68", x"18", x"60", x"20", x"B0", x"E5", x"C9",
x"71", x"F0", x"F5", x"C9", x"0D", x"F0", x"F5", x"68",
x"85", x"FF", x"68", x"85", x"FE", x"4C", x"DA", x"EE",
x"20", x"DC", x"E7", x"20", x"DC", x"E7", x"4C", x"DC",
x"E7", x"A5", x"FE", x"18", x"69", x"04", x"85", x"F6",
x"A5", x"FF", x"69", x"00", x"85", x"F7", x"60", x"20",
x"7D", x"E8", x"B0", x"FA", x"90", x"58", x"20", x"0C",
x"DB", x"18", x"60", x"20", x"9D", x"F9", x"D0", x"6A",
x"C9", x"01", x"F0", x"0E", x"A8", x"D0", x"53", x"20",
x"85", x"EF", x"D0", x"1E", x"20", x"3D", x"A7", x"4C",
x"C5", x"00", x"20", x"85", x"EF", x"D0", x"13", x"20",
x"B6", x"A4", x"4C", x"C5", x"00", x"AD", x"00", x"A4",
x"C9", x"A9", x"D0", x"05", x"AD", x"02", x"A4", x"C9",
x"8D", x"60", x"A9", x"EF", x"A0", x"9C", x"20", x"3B",
x"E6", x"4C", x"03", x"C0", x"0D", x"0A", x"0A", x"20",
x"43", x"52", x"54", x"20", x"4E", x"4F", x"54", x"20",
x"49", x"4D", x"50", x"4C", x"45", x"4D", x"45", x"4E",
x"54", x"45", x"44", x"0D", x"0A", x"04", x"20", x"F6",
x"E7", x"A5", x"FF", x"A6", x"FE", x"20", x"0C", x"DB",
x"18", x"60", x"C9", x"02", x"D0", x"0C", x"20", x"85",
x"EF", x"D0", x"C7", x"18", x"20", x"B6", x"A4", x"4C",
x"C5", x"00", x"A2", x"02", x"4C", x"59", x"C2", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"4C", x"6D", x"FA", x"4C", x"67", x"F0", x"4C", x"FF",
x"FF", x"4C", x"FF", x"FF", x"4C", x"A0", x"F3", x"4C",
x"87", x"F5", x"4C", x"73", x"F3", x"4C", x"0F", x"F5",
x"4C", x"D2", x"F5", x"4C", x"17", x"F4", x"4C", x"F6",
x"F0", x"4C", x"93", x"F8", x"4C", x"EE", x"FF", x"4C",
x"43", x"F4", x"4C", x"09", x"F3", x"4C", x"A1", x"F0",
x"4C", x"ED", x"F0", x"4C", x"90", x"F8", x"4C", x"B0",
x"F8", x"4C", x"57", x"F9", x"4C", x"82", x"F9", x"4C",
x"72", x"F1", x"4C", x"87", x"F1", x"4C", x"C4", x"F1",
x"4C", x"D6", x"FB", x"4C", x"D9", x"FB", x"4C", x"1F",
x"FC", x"20", x"C5", x"CC", x"20", x"C5", x"00", x"4C",
x"DC", x"D4", x"20", x"54", x"F0", x"86", x"E2", x"20",
x"51", x"F0", x"86", x"E3", x"4C", x"C5", x"00", x"20",
x"54", x"F0", x"86", x"E4", x"20", x"51", x"F0", x"86",
x"E5", x"20", x"8B", x"FE", x"20", x"C5", x"00", x"F0",
x"6D", x"20", x"51", x"F0", x"86", x"E4", x"4C", x"6C",
x"F0", x"20", x"5A", x"F0", x"20", x"69", x"FE", x"4C",
x"C5", x"00", x"20", x"5A", x"F0", x"20", x"51", x"F0",
x"86", x"F8", x"20", x"06", x"FF", x"4C", x"C5", x"00",
x"20", x"54", x"F0", x"8E", x"0A", x"02", x"4C", x"C5",
x"00", x"A9", x"00", x"8D", x"5A", x"02", x"20", x"ED",
x"F0", x"20", x"33", x"E6", x"C9", x"57", x"D0", x"03",
x"4C", x"03", x"C0", x"C9", x"43", x"D0", x"2F", x"A9",
x"14", x"8D", x"4F", x"02", x"A9", x"54", x"8D", x"66",
x"02", x"A9", x"FD", x"8D", x"5F", x"02", x"8D", x"61",
x"02", x"8D", x"63", x"02", x"8D", x"65", x"02", x"A9",
x"8F", x"8D", x"5E", x"02", x"A9", x"9D", x"8D", x"60",
x"02", x"A9", x"A1", x"8D", x"62", x"02", x"A9", x"AB",
x"8D", x"64", x"02", x"4C", x"00", x"C0", x"60", x"A9",
x"20", x"8D", x"40", x"02", x"60", x"20", x"E7", x"F0",
x"A9", x"20", x"8D", x"41", x"02", x"60", x"20", x"00",
x"C9", x"A5", x"81", x"85", x"14", x"A5", x"82", x"85",
x"15", x"20", x"36", x"C4", x"A0", x"02", x"B1", x"A7",
x"AA", x"C8", x"B1", x"A7", x"84", x"91", x"20", x"0C",
x"DB", x"A9", x"20", x"A4", x"91", x"29", x"7F", x"20",
x"51", x"F1", x"C8", x"B1", x"A7", x"D0", x"03", x"4C",
x"00", x"C9", x"10", x"F3", x"C9", x"C6", x"90", x"09",
x"20", x"85", x"F8", x"38", x"E9", x"C5", x"4C", x"37",
x"F1", x"20", x"7A", x"F8", x"38", x"E9", x"7F", x"AA",
x"84", x"91", x"A0", x"FF", x"CA", x"F0", x"07", x"C8",
x"B1", x"FE", x"10", x"FB", x"30", x"F6", x"C8", x"B1",
x"FE", x"30", x"C8", x"20", x"6C", x"C9", x"4C", x"46",
x"F1", x"20", x"6C", x"C9", x"98", x"38", x"65", x"A7",
x"85", x"A7", x"90", x"02", x"E6", x"A8", x"A0", x"FF",
x"84", x"91", x"C5", x"C6", x"D0", x"0B", x"A5", x"A8",
x"C5", x"C7", x"D0", x"05", x"A9", x"BF", x"20", x"6C",
x"C9", x"60", x"A2", x"0A", x"20", x"E3", x"E4", x"20",
x"B0", x"E5", x"90", x"09", x"F0", x"07", x"85", x"FC",
x"88", x"D0", x"EF", x"38", x"60", x"18", x"60", x"A4",
x"E9", x"B1", x"E6", x"60", x"8A", x"48", x"A2", x"00",
x"F0", x"04", x"8A", x"48", x"A2", x"05", x"A0", x"00",
x"B9", x"E6", x"00", x"9D", x"44", x"02", x"E8", x"C8",
x"C0", x"04", x"D0", x"F4", x"A8", x"68", x"AA", x"60",
x"8A", x"48", x"A2", x"00", x"F0", x"04", x"8A", x"48",
x"A2", x"05", x"A0", x"00", x"BD", x"44", x"02", x"99",
x"E6", x"00", x"E8", x"C8", x"C0", x"04", x"D0", x"F4",
x"A8", x"68", x"AA", x"60", x"C9", x"08", x"D0", x"1D",
x"2C", x"43", x"02", x"10", x"25", x"20", x"92", x"F1",
x"20", x"A8", x"F1", x"20", x"C2", x"E4", x"20", x"F2",
x"F1", x"20", x"8C", x"F1", x"20", x"C2", x"E4", x"20",
x"AE", x"F1", x"A9", x"08", x"60", x"C9", x"1F", x"D0",
x"18", x"2C", x"43", x"02", x"10", x"04", x"A9", x"08",
x"D0", x"25", x"A9", x"08", x"20", x"50", x"E7", x"A9",
x"20", x"20", x"50", x"E7", x"A9", x"08", x"4C", x"50",
x"E7", x"C9", x"0A", x"D0", x"18", x"2C", x"43", x"02",
x"30", x"0D", x"48", x"A9", x"FF", x"8D", x"43", x"02",
x"20", x"8C", x"F1", x"20", x"C2", x"E4", x"68", x"20",
x"50", x"E7", x"6C", x"16", x"02", x"C9", x"09", x"F0",
x"E4", x"C9", x"0B", x"F0", x"E0", x"C9", x"0D", x"D0",
x"15", x"2C", x"43", x"02", x"10", x"0D", x"48", x"20",
x"A8", x"F1", x"20", x"C2", x"E4", x"A9", x"00", x"8D",
x"43", x"02", x"68", x"4C", x"50", x"E7", x"C9", x"14",
x"F0", x"23", x"C9", x"20", x"90", x"F5", x"48", x"2C",
x"43", x"02", x"10", x"EE", x"20", x"92", x"F1", x"20",
x"A8", x"F1", x"20", x"C2", x"E4", x"68", x"48", x"20",
x"50", x"E7", x"20", x"8C", x"F1", x"20", x"C2", x"E4",
x"20", x"AE", x"F1", x"68", x"60", x"2C", x"43", x"02",
x"30", x"03", x"6C", x"16", x"02", x"20", x"92", x"F1",
x"20", x"A8", x"F1", x"20", x"C2", x"E4", x"20", x"8D",
x"F2", x"20", x"8C", x"F1", x"20", x"C2", x"E4", x"20",
x"AE", x"F1", x"A9", x"09", x"20", x"50", x"E7", x"AD",
x"48", x"02", x"F0", x"DE", x"60", x"8A", x"48", x"98",
x"48", x"AD", x"49", x"02", x"18", x"6D", x"4C", x"02",
x"69", x"20", x"85", x"F0", x"85", x"FC", x"AD", x"4A",
x"02", x"85", x"F1", x"A2", x"00", x"A9", x"20", x"8D",
x"48", x"02", x"E8", x"A9", x"20", x"8D", x"5D", x"02",
x"BD", x"00", x"02", x"85", x"FE", x"BD", x"04", x"02",
x"85", x"FF", x"A0", x"00", x"84", x"FA", x"A0", x"00",
x"B1", x"F0", x"A4", x"FA", x"D1", x"FE", x"F0", x"1E",
x"EE", x"48", x"02", x"2C", x"48", x"02", x"30", x"32",
x"A5", x"FC", x"85", x"F0", x"A5", x"FE", x"CE", x"5D",
x"02", x"F0", x"CF", x"18", x"69", x"08", x"85", x"FE",
x"90", x"D8", x"E6", x"FF", x"D0", x"D4", x"C8", x"84",
x"FA", x"C0", x"07", x"F0", x"0A", x"A5", x"F0", x"18",
x"69", x"20", x"85", x"F0", x"4C", x"BE", x"F2", x"AD",
x"48", x"02", x"20", x"50", x"E7", x"68", x"A8", x"68",
x"AA", x"60", x"A9", x"00", x"8D", x"48", x"02", x"F0",
x"F4", x"24", x"10", x"30", x"12", x"48", x"C9", x"20",
x"90", x"0C", x"A5", x"11", x"C5", x"12", x"D0", x"04",
x"A9", x"00", x"85", x"11", x"E6", x"11", x"68", x"29",
x"FF", x"60", x"A9", x"20", x"A2", x"09", x"9D", x"50",
x"02", x"CA", x"10", x"FA", x"20", x"C5", x"00", x"D0",
x"03", x"4C", x"92", x"FA", x"20", x"71", x"F6", x"CA",
x"F0", x"0A", x"B1", x"6A", x"99", x"50", x"02", x"C8",
x"C0", x"0A", x"D0", x"F3", x"4C", x"C5", x"00", x"86",
x"FA", x"A2", x"03", x"A9", x"1B", x"9D", x"80", x"02",
x"CA", x"10", x"FA", x"A9", x"42", x"8D", x"84", x"02",
x"A2", x"05", x"BD", x"4B", x"02", x"9D", x"80", x"02",
x"E8", x"E0", x"0F", x"D0", x"F5", x"AD", x"4E", x"02",
x"8D", x"8F", x"02", x"A9", x"10", x"8D", x"4D", x"02",
x"A6", x"FA", x"60", x"8A", x"48", x"AD", x"66", x"02",
x"8D", x"41", x"02", x"20", x"C5", x"00", x"20", x"22",
x"F3", x"BA", x"9D", x"04", x"01", x"A9", x"00", x"8D",
x"4E", x"02", x"20", x"47", x"F3", x"AD", x"41", x"02",
x"C9", x"44", x"D0", x"09", x"38", x"20", x"E1", x"F3",
x"90", x"03", x"4C", x"60", x"FD", x"68", x"AA", x"60",
x"85", x"FC", x"48", x"8A", x"48", x"98", x"48", x"20",
x"40", x"C6", x"A5", x"FC", x"AE", x"4D", x"02", x"9D",
x"80", x"02", x"EE", x"4D", x"02", x"D0", x"11", x"20",
x"D1", x"F3", x"EE", x"4E", x"02", x"AD", x"4E", x"02",
x"8D", x"8F", x"02", x"A9", x"10", x"8D", x"4D", x"02",
x"68", x"A8", x"68", x"AA", x"20", x"C5", x"00", x"68",
x"60", x"AD", x"41", x"02", x"C9", x"44", x"D0", x"0C",
x"20", x"E0", x"F3", x"90", x"F3", x"4C", x"60", x"FD",
x"18", x"6C", x"5E", x"02", x"AD", x"4F", x"02", x"A2",
x"00", x"A0", x"14", x"20", x"B7", x"E7", x"8D", x"00",
x"88", x"CA", x"D0", x"F5", x"A8", x"88", x"98", x"D0",
x"F0", x"A0", x"08", x"20", x"DC", x"ED", x"EA", x"EA",
x"EA", x"20", x"D7", x"ED", x"AE", x"4D", x"02", x"BD",
x"80", x"02", x"A2", x"07", x"A0", x"06", x"20", x"DC",
x"ED", x"EE", x"4D", x"02", x"D0", x"E8", x"60", x"8A",
x"48", x"AE", x"4D", x"02", x"A9", x"20", x"9D", x"80",
x"02", x"E8", x"D0", x"FA", x"8E", x"4D", x"02", x"20",
x"D1", x"F3", x"AD", x"41", x"02", x"C9", x"44", x"D0",
x"0B", x"20", x"39", x"F4", x"90", x"06", x"4C", x"60",
x"FD", x"6C", x"60", x"02", x"20", x"ED", x"F0", x"68",
x"AA", x"18", x"60", x"48", x"AD", x"40", x"02", x"20",
x"D8", x"C6", x"F0", x"04", x"68", x"4C", x"F1", x"FF",
x"68", x"60", x"8A", x"48", x"A2", x"00", x"BD", x"50",
x"02", x"20", x"F1", x"FF", x"E8", x"E0", x"0A", x"D0",
x"F5", x"68", x"AA", x"A9", x"22", x"4C", x"F1", x"FF",
x"8A", x"48", x"AD", x"40", x"02", x"C9", x"44", x"F0",
x"43", x"A2", x"00", x"BD", x"85", x"02", x"20", x"F1",
x"FF", x"E8", x"E0", x"0A", x"D0", x"F5", x"A9", x"22",
x"20", x"F1", x"FF", x"A9", x"20", x"20", x"F1", x"FF",
x"AD", x"84", x"02", x"20", x"F1", x"FF", x"AE", x"8F",
x"02", x"AD", x"40", x"02", x"48", x"20", x"E7", x"F0",
x"A9", x"00", x"20", x"0C", x"DB", x"68", x"8D", x"40",
x"02", x"AD", x"84", x"02", x"C9", x"4F", x"D0", x"0C",
x"AD", x"91", x"02", x"20", x"00", x"E8", x"AD", x"90",
x"02", x"20", x"03", x"E8", x"68", x"AA", x"60", x"A2",
x"05", x"BD", x"4B", x"02", x"C9", x"20", x"F0", x"0A",
x"DD", x"80", x"02", x"D0", x"10", x"E8", x"E0", x"0F",
x"D0", x"EF", x"08", x"AD", x"8F", x"02", x"D0", x"03",
x"28", x"18", x"60", x"28", x"38", x"60", x"AD", x"40",
x"02", x"C9", x"44", x"F0", x"F8", x"B9", x"24", x"F6",
x"F0", x"F3", x"20", x"F1", x"FF", x"C8", x"D0", x"F5",
x"AD", x"40", x"02", x"C9", x"44", x"D0", x"08", x"20",
x"F8", x"F4", x"90", x"03", x"4C", x"60", x"FD", x"60",
x"38", x"6C", x"62", x"02", x"AD", x"40", x"02", x"C9",
x"44", x"D0", x"09", x"18", x"20", x"F9", x"F4", x"90",
x"EE", x"4C", x"60", x"FD", x"4C", x"F1", x"F5", x"AD",
x"66", x"02", x"8D", x"40", x"02", x"8A", x"48", x"98",
x"48", x"20", x"C5", x"00", x"20", x"22", x"F3", x"20",
x"E8", x"F4", x"A9", x"42", x"48", x"A0", x"00", x"AD",
x"40", x"02", x"C9", x"44", x"F0", x"06", x"20", x"D6",
x"F4", x"20", x"52", x"F4", x"20", x"FC", x"F4", x"20",
x"B7", x"F4", x"F0", x"0B", x"A0", x"1C", x"20", x"D6",
x"F4", x"20", x"68", x"F4", x"4C", x"34", x"F5", x"90",
x"1E", x"A0", x"1C", x"20", x"D6", x"F4", x"20", x"68",
x"F4", x"68", x"48", x"CD", x"84", x"02", x"D0", x"DC",
x"A0", x"2A", x"20", x"D6", x"F4", x"20", x"EE", x"FF",
x"C9", x"0D", x"F0", x"D0", x"4C", x"58", x"C6", x"68",
x"48", x"CD", x"84", x"02", x"D0", x"CE", x"68", x"A0",
x"0E", x"20", x"D6", x"F4", x"20", x"68", x"F4", x"A9",
x"10", x"8D", x"4D", x"02", x"A9", x"01", x"8D", x"4E",
x"02", x"68", x"A8", x"68", x"AA", x"18", x"60", x"8A",
x"48", x"98", x"48", x"AE", x"4D", x"02", x"F0", x"10",
x"BD", x"80", x"02", x"EE", x"4D", x"02", x"85", x"FA",
x"68", x"A8", x"68", x"AA", x"A5", x"FA", x"18", x"60",
x"20", x"FC", x"F4", x"A0", x"1C", x"20", x"D6", x"F4",
x"20", x"68", x"F4", x"20", x"B7", x"F4", x"F0", x"0F",
x"A0", x"39", x"20", x"D6", x"F4", x"20", x"DE", x"F5",
x"20", x"ED", x"F0", x"A9", x"1A", x"D0", x"D7", x"AD",
x"8F", x"02", x"CD", x"4E", x"02", x"D0", x"E9", x"EE",
x"4E", x"02", x"A9", x"10", x"8D", x"4D", x"02", x"4C",
x"8B", x"F5", x"20", x"DE", x"F5", x"20", x"ED", x"F0",
x"20", x"00", x"C9", x"4C", x"00", x"C9", x"AD", x"40",
x"02", x"C9", x"44", x"D0", x"08", x"20", x"EE", x"F5",
x"90", x"03", x"4C", x"60", x"FD", x"60", x"6C", x"64",
x"02", x"20", x"40", x"C6", x"A9", x"04", x"8D", x"4D",
x"02", x"A0", x"20", x"20", x"1C", x"EE", x"90", x"F1",
x"88", x"D0", x"F8", x"20", x"47", x"EE", x"A9", x"04",
x"85", x"FA", x"20", x"12", x"EE", x"C9", x"1B", x"D0",
x"E0", x"C6", x"FA", x"D0", x"F5", x"20", x"12", x"EE",
x"AE", x"4D", x"02", x"9D", x"80", x"02", x"EE", x"4D",
x"02", x"D0", x"F2", x"60", x"0D", x"0A", x"53", x"45",
x"41", x"52", x"43", x"48", x"49", x"4E", x"47", x"20",
x"22", x"00", x"0D", x"0A", x"4C", x"4F", x"41", x"44",
x"49", x"4E", x"47", x"20", x"20", x"20", x"22", x"00",
x"0D", x"0A", x"20", x"20", x"20", x"20", x"20", x"20",
x"20", x"20", x"20", x"20", x"22", x"00", x"0D", x"0A",
x"0A", x"52", x"45", x"57", x"49", x"4E", x"44", x"20",
x"54", x"41", x"50", x"45", x"00", x"0D", x"0A", x"0A",
x"4C", x"4F", x"41", x"44", x"49", x"4E", x"47", x"20",
x"45", x"52", x"52", x"4F", x"52", x"0D", x"0A", x"0A",
x"00", x"20", x"7F", x"CB", x"20", x"70", x"CB", x"20",
x"E4", x"D3", x"AA", x"A0", x"00", x"E8", x"60", x"20",
x"71", x"F6", x"CA", x"F0", x"08", x"B1", x"6A", x"99",
x"80", x"02", x"C8", x"D0", x"F5", x"A9", x"00", x"99",
x"80", x"02", x"20", x"C5", x"00", x"20", x"51", x"F0",
x"8E", x"5B", x"02", x"20", x"51", x"F0", x"8A", x"29",
x"03", x"6A", x"6A", x"6A", x"8D", x"5C", x"02", x"A2",
x"00", x"AD", x"0A", x"02", x"48", x"BD", x"80", x"02",
x"F0", x"08", x"20", x"C6", x"F6", x"B0", x"0A", x"E8",
x"D0", x"F3", x"68", x"8D", x"0A", x"02", x"4C", x"C5",
x"00", x"A2", x"08", x"4C", x"59", x"C2", x"29", x"7F",
x"85", x"FC", x"C9", x"20", x"B0", x"02", x"38", x"60",
x"8A", x"48", x"98", x"48", x"A5", x"FC", x"A8", x"2A",
x"2A", x"2A", x"2A", x"29", x"03", x"AA", x"BD", x"00",
x"02", x"D0", x"03", x"BD", x"04", x"02", x"85", x"FF",
x"98", x"0A", x"0A", x"0A", x"85", x"FE", x"A5", x"E2",
x"8D", x"50", x"02", x"A5", x"E3", x"8D", x"51", x"02",
x"A0", x"07", x"AD", x"5B", x"02", x"8D", x"52", x"02",
x"2C", x"5C", x"02", x"50", x"08", x"A5", x"E3", x"8D",
x"53", x"02", x"4C", x"12", x"F7", x"A5", x"E2", x"8D",
x"53", x"02", x"B1", x"FE", x"A2", x"08", x"48", x"6A",
x"90", x"06", x"20", x"75", x"F7", x"4C", x"23", x"F7",
x"20", x"79", x"F7", x"68", x"6A", x"CA", x"D0", x"EE",
x"AD", x"53", x"02", x"2C", x"5C", x"02", x"50", x"10",
x"08", x"85", x"E3", x"28", x"10", x"05", x"E6", x"E2",
x"4C", x"4D", x"F7", x"C6", x"E2", x"4C", x"4D", x"F7",
x"08", x"85", x"E2", x"28", x"10", x"05", x"C6", x"E3",
x"4C", x"4D", x"F7", x"E6", x"E3", x"CE", x"52", x"02",
x"D0", x"C0", x"88", x"10", x"A5", x"AD", x"50", x"02",
x"85", x"E2", x"AD", x"51", x"02", x"85", x"E3", x"AE",
x"5B", x"02", x"F0", x"0B", x"A0", x"08", x"20", x"91",
x"F7", x"88", x"D0", x"FA", x"CA", x"D0", x"F5", x"68",
x"A8", x"68", x"AA", x"18", x"60", x"A9", x"00", x"F0",
x"02", x"A9", x"01", x"8D", x"0A", x"02", x"8A", x"48",
x"AE", x"5B", x"02", x"F0", x"09", x"20", x"69", x"FE",
x"20", x"91", x"F7", x"CA", x"D0", x"F7", x"68", x"AA",
x"60", x"2C", x"5C", x"02", x"30", x"05", x"70", x"0B",
x"E6", x"E2", x"60", x"70", x"03", x"C6", x"E2", x"60",
x"C6", x"E3", x"60", x"E6", x"E3", x"60", x"4D", x"4F",
x"44", x"C5", x"4D", x"4F", x"56", x"C5", x"45", x"58",
x"49", x"D4", x"4C", x"4E", x"CB", x"4C", x"45", x"54",
x"54", x"45", x"D2", x"44", x"4D", x"45", x"CD", x"4C",
x"4D", x"45", x"CD", x"49", x"4E", x"4B", x"45", x"D9",
x"4F", x"50", x"45", x"4E", x"D7", x"57", x"52", x"49",
x"54", x"C5", x"43", x"4C", x"4F", x"53", x"45", x"D7",
x"4F", x"50", x"45", x"4E", x"C7", x"43", x"4C", x"4F",
x"53", x"45", x"C7", x"53", x"4F", x"55", x"4E", x"C4",
x"43", x"4C", x"D3", x"56", x"44", x"D5", x"52", x"41",
x"54", x"C5", x"43", x"55", x"D2", x"54", x"47", x"41",
x"D0", x"53", x"43", x"52", x"45", x"45", x"4E", x"A4",
x"44", x"4F", x"D4", x"43", x"52", x"D4", x"49", x"4E",
x"D6", x"53", x"4D", x"4F", x"56", x"C5", x"43", x"49",
x"D2", x"50", x"4C", x"4F", x"D4", x"50", x"54", x"D2",
x"44", x"4F", x"53", x"C9", x"44", x"4F", x"D3", x"43",
x"4F", x"4D", x"CD", x"41", x"54", x"45", x"4F", x"C6",
x"54", x"41", x"50", x"C5", x"44", x"49", x"53", x"CB",
x"43", x"48", x"41", x"D2", x"00", x"00", x"97", x"F0",
x"59", x"F0", x"FB", x"FD", x"8D", x"F9", x"7E", x"F6",
x"AE", x"F9", x"01", x"FA", x"A7", x"F9", x"4F", x"FA",
x"70", x"FA", x"C5", x"FA", x"DD", x"FA", x"01", x"FB",
x"09", x"FB", x"33", x"FB", x"42", x"FB", x"81", x"FB",
x"A2", x"FB", x"BC", x"FB", x"EA", x"FB", x"02", x"FC",
x"62", x"EF", x"2F", x"FC", x"3F", x"FC", x"89", x"F0",
x"80", x"F0", x"70", x"FB", x"C5", x"FB", x"CD", x"FB",
x"67", x"FD", x"C5", x"FD", x"53", x"FD", x"5B", x"FD",
x"D5", x"FD", x"48", x"A9", x"90", x"85", x"FE", x"A9",
x"C0", x"85", x"FF", x"68", x"60", x"48", x"A9", x"A6",
x"85", x"FE", x"A9", x"F7", x"85", x"FF", x"68", x"60",
x"D0", x"01", x"60", x"E9", x"80", x"B0", x"03", x"4C",
x"05", x"C6", x"C9", x"46", x"B0", x"03", x"4C", x"07",
x"C6", x"E9", x"46", x"0A", x"A8", x"B9", x"37", x"F8",
x"48", x"B9", x"36", x"F8", x"48", x"4C", x"BF", x"00",
x"20", x"7A", x"F8", x"A9", x"00", x"8D", x"5B", x"02",
x"20", x"C5", x"F8", x"20", x"85", x"F8", x"A9", x"80",
x"8D", x"5B", x"02", x"E6", x"C6", x"A6", x"C6", x"A0",
x"04", x"84", x"0C", x"B5", x"00", x"30", x"41", x"C9",
x"20", x"F0", x"3D", x"85", x"07", x"C9", x"22", x"F0",
x"5B", x"24", x"0C", x"70", x"33", x"C9", x"3F", x"D0",
x"04", x"A9", x"97", x"D0", x"2B", x"C9", x"30", x"90",
x"04", x"C9", x"3C", x"90", x"23", x"84", x"B9", x"A0",
x"00", x"84", x"08", x"88", x"86", x"C6", x"CA", x"C8",
x"E8", x"B5", x"00", x"38", x"F1", x"FE", x"F0", x"F7",
x"C9", x"80", x"D0", x"37", x"05", x"08", x"2C", x"5B",
x"02", x"10", x"03", x"18", x"69", x"46", x"A4", x"B9",
x"E8", x"C8", x"99", x"11", x"00", x"B9", x"11", x"00",
x"F0", x"32", x"38", x"E9", x"3A", x"F0", x"04", x"C9",
x"49", x"D0", x"02", x"85", x"0C", x"38", x"E9", x"54",
x"D0", x"A1", x"85", x"07", x"B5", x"00", x"F0", x"E0",
x"C5", x"07", x"F0", x"DC", x"C8", x"99", x"11", x"00",
x"E8", x"D0", x"F1", x"A6", x"C6", x"E6", x"08", x"B1",
x"FE", x"10", x"11", x"C8", x"B1", x"FE", x"D0", x"B1",
x"B5", x"00", x"10", x"C2", x"99", x"13", x"00", x"A9",
x"15", x"85", x"C6", x"60", x"C8", x"D0", x"E8", x"38",
x"E9", x"7F", x"C9", x"47", x"B0", x"03", x"4C", x"41",
x"C5", x"E9", x"46", x"AA", x"84", x"91", x"A0", x"FF",
x"CA", x"F0", x"08", x"C8", x"B9", x"A6", x"F7", x"10",
x"FA", x"30", x"F5", x"C8", x"B9", x"A6", x"F7", x"10",
x"03", x"4C", x"0C", x"C5", x"20", x"6C", x"C9", x"4C",
x"73", x"F9", x"C9", x"60", x"F0", x"07", x"C9", x"80",
x"90", x"02", x"18", x"60", x"38", x"60", x"20", x"9D",
x"F9", x"20", x"97", x"F9", x"4C", x"C5", x"00", x"6C",
x"14", x"00", x"20", x"C5", x"CC", x"20", x"6B", x"CB",
x"20", x"36", x"D5", x"A5", x"14", x"A4", x"15", x"60",
x"A9", x"00", x"85", x"FA", x"4C", x"AD", x"C9", x"48",
x"A9", x"54", x"8D", x"41", x"02", x"68", x"20", x"22",
x"F3", x"20", x"47", x"F3", x"A9", x"4F", x"8D", x"84",
x"02", x"20", x"9A", x"F9", x"85", x"F4", x"8D", x"90",
x"02", x"84", x"F5", x"8C", x"91", x"02", x"20", x"9A",
x"F9", x"85", x"FE", x"8D", x"92", x"02", x"84", x"FF",
x"8C", x"93", x"02", x"A9", x"00", x"8D", x"8F", x"02",
x"A2", x"14", x"A9", x"20", x"9D", x"80", x"02", x"E8",
x"D0", x"FA", x"8E", x"4D", x"02", x"20", x"E4", x"F3",
x"AD", x"4F", x"02", x"E6", x"FE", x"E6", x"FF", x"20",
x"99", x"ED", x"A9", x"20", x"8D", x"41", x"02", x"4C",
x"C5", x"00", x"48", x"A9", x"54", x"8D", x"40", x"02",
x"68", x"20", x"22", x"F3", x"A0", x"4F", x"20", x"49",
x"FA", x"A5", x"7B", x"48", x"A5", x"7C", x"48", x"AD",
x"90", x"02", x"38", x"E9", x"01", x"85", x"7B", x"AD",
x"91", x"02", x"E9", x"00", x"85", x"7C", x"20", x"C5",
x"00", x"F0", x"0D", x"20", x"9A", x"F9", x"38", x"E9",
x"01", x"85", x"7B", x"98", x"E9", x"00", x"85", x"7C",
x"20", x"6D", x"EE", x"A9", x"20", x"8D", x"40", x"02",
x"68", x"85", x"7C", x"68", x"85", x"7B", x"4C", x"C5",
x"00", x"8A", x"48", x"98", x"48", x"4C", x"24", x"F5",
x"20", x"22", x"F3", x"A9", x"00", x"8D", x"4E", x"02",
x"A9", x"80", x"8D", x"5A", x"02", x"20", x"47", x"F3",
x"A9", x"44", x"8D", x"84", x"02", x"A9", x"54", x"8D",
x"41", x"02", x"4C", x"C5", x"00", x"A9", x"00", x"F0",
x"06", x"C9", x"23", x"D0", x"0F", x"A9", x"80", x"A0",
x"00", x"20", x"42", x"B0", x"A2", x"1C", x"20", x"06",
x"B0", x"B0", x"0F", x"60", x"AD", x"41", x"02", x"C9",
x"54", x"D0", x"07", x"2C", x"5A", x"02", x"70", x"02",
x"30", x"08", x"20", x"ED", x"F0", x"A2", x"02", x"4C",
x"59", x"C2", x"20", x"C5", x"00", x"D0", x"03", x"4C",
x"00", x"C9", x"20", x"7F", x"CB", x"24", x"0A", x"30",
x"06", x"20", x"1C", x"DB", x"20", x"C5", x"D1", x"20",
x"4D", x"C9", x"20", x"C5", x"00", x"F0", x"E8", x"C9",
x"2C", x"D0", x"D7", x"20", x"A0", x"F3", x"20", x"BF",
x"00", x"D0", x"DF", x"4C", x"00", x"C9", x"2C", x"5A",
x"02", x"10", x"C7", x"A9", x"1A", x"20", x"A0", x"F3",
x"20", x"A0", x"F3", x"A9", x"00", x"8D", x"5A", x"02",
x"20", x"17", x"F4", x"4C", x"C5", x"00", x"20", x"22",
x"F3", x"A9", x"54", x"8D", x"40", x"02", x"A0", x"44",
x"20", x"49", x"FA", x"A9", x"40", x"8D", x"5A", x"02",
x"4C", x"C5", x"00", x"2C", x"5A", x"02", x"50", x"9A",
x"30", x"98", x"20", x"87", x"F5", x"C9", x"1A", x"F0",
x"01", x"60", x"A9", x"00", x"8D", x"5A", x"02", x"4C",
x"D2", x"F5", x"20", x"54", x"F0", x"8E", x"5B", x"02",
x"20", x"51", x"F0", x"8E", x"5C", x"02", x"AE", x"5B",
x"02", x"A0", x"00", x"F0", x"0B", x"AD", x"00", x"88",
x"88", x"D0", x"05", x"CE", x"5C", x"02", x"F0", x"09",
x"CA", x"D0", x"F5", x"AE", x"5B", x"02", x"4C", x"1D",
x"FB", x"4C", x"C5", x"00", x"A9", x"0C", x"20", x"F1",
x"FF", x"A9", x"00", x"85", x"11", x"20", x"9D", x"E3",
x"4C", x"C5", x"00", x"20", x"C5", x"00", x"F0", x"17",
x"20", x"54", x"F0", x"86", x"EC", x"20", x"51", x"F0",
x"86", x"ED", x"20", x"51", x"F0", x"86", x"EA", x"20",
x"51", x"F0", x"86", x"EB", x"4C", x"C5", x"00", x"20",
x"64", x"FB", x"D0", x"D0", x"A9", x"00", x"85", x"EC",
x"85", x"EA", x"A9", x"1F", x"85", x"ED", x"85", x"EB",
x"60", x"20", x"54", x"F0", x"8A", x"C9", x"02", x"B0",
x"10", x"18", x"6A", x"6A", x"8D", x"10", x"02", x"4C",
x"C5", x"00", x"20", x"54", x"F0", x"E0", x"04", x"90",
x"05", x"A2", x"08", x"4C", x"59", x"C2", x"BD", x"97",
x"FB", x"8D", x"13", x"02", x"4C", x"C5", x"00", x"A7",
x"53", x"2A", x"15", x"00", x"01", x"03", x"07", x"0F",
x"1F", x"3F", x"7F", x"20", x"54", x"F0", x"8A", x"29",
x"1F", x"85", x"11", x"85", x"E9", x"20", x"51", x"F0",
x"8A", x"29", x"1F", x"85", x"E8", x"18", x"69", x"0F",
x"85", x"E7", x"4C", x"3D", x"FB", x"20", x"54", x"F0",
x"8E", x"4F", x"02", x"4C", x"C5", x"00", x"20", x"00",
x"B0", x"90", x"08", x"4C", x"60", x"FD", x"20", x"12",
x"B0", x"B0", x"F8", x"4C", x"C5", x"00", x"4C", x"F6",
x"E7", x"20", x"C5", x"00", x"C9", x"D9", x"F0", x"0B",
x"C9", x"DA", x"F0", x"1F", x"C9", x"DB", x"F0", x"31",
x"4C", x"7F", x"CB", x"20", x"92", x"F1", x"20", x"8D",
x"F2", x"A9", x"01", x"20", x"BB", x"D1", x"A0", x"00",
x"AD", x"48", x"02", x"91", x"AA", x"20", x"08", x"D2",
x"4C", x"BF", x"00", x"20", x"5A", x"FE", x"E8", x"B1",
x"E0", x"2A", x"6A", x"CA", x"D0", x"FC", x"29", x"01",
x"A8", x"A9", x"00", x"20", x"D1", x"D0", x"4C", x"BF",
x"00", x"20", x"9F", x"E7", x"4C", x"11", x"FC", x"20",
x"8C", x"F1", x"20", x"AE", x"F1", x"C6", x"E8", x"20",
x"9D", x"E3", x"20", x"92", x"F1", x"4C", x"A8", x"F1",
x"20", x"54", x"F0", x"8A", x"D0", x"06", x"8D", x"0E",
x"02", x"4C", x"C5", x"00", x"A9", x"FF", x"D0", x"F6",
x"20", x"54", x"F0", x"8A", x"29", x"03", x"18", x"6A",
x"6A", x"6A", x"8D", x"5B", x"02", x"20", x"9A", x"F9",
x"20", x"5A", x"FE", x"18", x"98", x"65", x"E0", x"85",
x"E0", x"8E", x"50", x"02", x"A2", x"00", x"A0", x"00",
x"B1", x"14", x"9D", x"A0", x"02", x"E8", x"C8", x"B1",
x"14", x"9D", x"A0", x"02", x"C8", x"E8", x"A9", x"00",
x"9D", x"A0", x"02", x"E8", x"C0", x"20", x"D0", x"E8",
x"A2", x"00", x"AC", x"50", x"02", x"F0", x"14", x"18",
x"7E", x"A0", x"02", x"7E", x"A1", x"02", x"7E", x"A2",
x"02", x"88", x"D0", x"F3", x"E8", x"E8", x"E8", x"E0",
x"30", x"D0", x"E7", x"A2", x"2F", x"A0", x"08", x"A9",
x"00", x"8D", x"51", x"02", x"18", x"BD", x"A0", x"02",
x"6A", x"2E", x"51", x"02", x"88", x"D0", x"F9", x"AD",
x"51", x"02", x"9D", x"A0", x"02", x"CA", x"10", x"E5",
x"AE", x"50", x"02", x"AD", x"5B", x"02", x"C9", x"40",
x"F0", x"04", x"C9", x"80", x"D0", x"5B", x"BD", x"9B",
x"FB", x"8D", x"51", x"02", x"49", x"FF", x"8D", x"52",
x"02", x"A2", x"00", x"A0", x"00", x"B1", x"E0", x"2D",
x"51", x"02", x"1D", x"A0", x"02", x"2C", x"5B", x"02",
x"10", x"02", x"31", x"E0", x"91", x"E0", x"C8", x"BD",
x"A1", x"02", x"2C", x"5B", x"02", x"10", x"05", x"B1",
x"E0", x"3D", x"A1", x"02", x"91", x"E0", x"C8", x"B1",
x"E0", x"2D", x"52", x"02", x"1D", x"A2", x"02", x"2C",
x"5B", x"02", x"10", x"02", x"31", x"E0", x"91", x"E0",
x"20", x"08", x"FD", x"D0", x"C6", x"4C", x"C5", x"00",
x"18", x"A5", x"E0", x"69", x"20", x"85", x"E0", x"90",
x"02", x"E6", x"E1", x"E8", x"E8", x"E8", x"E0", x"30",
x"60", x"A2", x"00", x"A0", x"00", x"B1", x"E0", x"2C",
x"5B", x"02", x"50", x"05", x"1D", x"A0", x"02", x"70",
x"03", x"5D", x"A0", x"02", x"91", x"E0", x"C8", x"B1",
x"E0", x"50", x"05", x"1D", x"A1", x"02", x"70", x"03",
x"5D", x"A1", x"02", x"91", x"E0", x"C8", x"B1", x"E0",
x"50", x"05", x"1D", x"A2", x"02", x"70", x"03", x"5D",
x"A2", x"02", x"91", x"E0", x"20", x"08", x"FD", x"D0",
x"CA", x"4C", x"C5", x"00", x"A9", x"54", x"8D", x"66",
x"02", x"4C", x"C5", x"00", x"A9", x"44", x"D0", x"F6",
x"A9", x"FF", x"8D", x"00", x"5F", x"4C", x"92", x"FA",
x"20", x"71", x"F6", x"CA", x"F0", x"0A", x"B1", x"6A",
x"99", x"22", x"5F", x"C8", x"C0", x"50", x"D0", x"F3",
x"A9", x"00", x"99", x"22", x"5F", x"A2", x"0A", x"20",
x"06", x"B0", x"B0", x"DC", x"CE", x"21", x"5F", x"20",
x"48", x"B0", x"B0", x"D4", x"4C", x"C5", x"00", x"90",
x"08", x"A2", x"16", x"20", x"06", x"B0", x"B0", x"C8",
x"60", x"A2", x"17", x"D0", x"F6", x"A2", x"19", x"D0",
x"F2", x"90", x"04", x"A2", x"1A", x"D0", x"EC", x"A2",
x"1B", x"D0", x"E8", x"AD", x"5C", x"5E", x"AC", x"5D",
x"5E", x"20", x"42", x"B0", x"20", x"0C", x"B0", x"B0",
x"A7", x"A9", x"00", x"8D", x"5C", x"5E", x"8D", x"5D",
x"5E", x"20", x"ED", x"F0", x"18", x"60", x"20", x"DA",
x"C7", x"AD", x"1A", x"5F", x"29", x"01", x"D0", x"03",
x"4C", x"C5", x"00", x"4C", x"17", x"C7", x"20", x"54",
x"F0", x"E0", x"03", x"90", x"03", x"4C", x"C1", x"F6",
x"8A", x"48", x"20", x"51", x"F0", x"68", x"A8", x"E0",
x"00", x"F0", x"0B", x"E0", x"04", x"90", x"EE", x"8A",
x"99", x"05", x"02", x"4C", x"C5", x"00", x"18", x"98",
x"69", x"E0", x"D0", x"F4", x"A2", x"FF", x"9A", x"20",
x"64", x"FB", x"4C", x"A3", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"A5", x"E3", x"49", x"FF", x"AA",
x"4A", x"4A", x"4A", x"20", x"8E", x"EE", x"EA", x"8A",
x"0A", x"0A", x"0A", x"0A", x"0A", x"85", x"E0", x"60",
x"FF", x"FF", x"FF", x"A5", x"E2", x"4A", x"4A", x"4A",
x"A8", x"60", x"01", x"02", x"04", x"08", x"10", x"20",
x"40", x"80", x"20", x"33", x"FE", x"20", x"4B", x"FE",
x"A5", x"E2", x"29", x"07", x"AA", x"BD", x"52", x"FE",
x"60", x"8A", x"48", x"98", x"48", x"20", x"5A", x"FE",
x"18", x"AE", x"0A", x"02", x"30", x"06", x"D0", x"08",
x"11", x"E0", x"90", x"08", x"51", x"E0", x"90", x"04",
x"49", x"FF", x"31", x"E0", x"91", x"E0", x"68", x"A8",
x"68", x"AA", x"60", x"8A", x"48", x"98", x"48", x"A2",
x"01", x"A5", x"E4", x"38", x"E5", x"E2", x"B0", x"06",
x"A2", x"FF", x"49", x"FF", x"69", x"01", x"85", x"F4",
x"85", x"F8", x"4A", x"69", x"00", x"85", x"F7", x"A0",
x"01", x"A5", x"E5", x"38", x"E5", x"E3", x"B0", x"06",
x"A0", x"FF", x"49", x"FF", x"69", x"01", x"85", x"F6",
x"C5", x"F4", x"B0", x"02", x"85", x"F8", x"4A", x"69",
x"00", x"85", x"F5", x"18", x"90", x"2C", x"A5", x"F5",
x"38", x"E5", x"F8", x"85", x"F5", x"90", x"03", x"D0",
x"0B", x"18", x"65", x"F6", x"85", x"F5", x"8A", x"18",
x"65", x"E2", x"85", x"E2", x"A5", x"F7", x"38", x"E5",
x"F8", x"85", x"F7", x"90", x"03", x"D0", x"0B", x"18",
x"65", x"F4", x"85", x"F7", x"98", x"18", x"65", x"E3",
x"85", x"E3", x"20", x"69", x"FE", x"A5", x"E2", x"C5",
x"E4", x"D0", x"CB", x"A5", x"E3", x"C5", x"E5", x"D0",
x"C5", x"68", x"A8", x"68", x"AA", x"60", x"8A", x"48",
x"98", x"48", x"A5", x"E2", x"85", x"E4", x"A5", x"E3",
x"85", x"E5", x"A9", x"00", x"85", x"F6", x"85", x"F7",
x"A9", x"7F", x"85", x"F4", x"A5", x"F8", x"85", x"F5",
x"A2", x"04", x"A0", x"24", x"A5", x"F7", x"0A", x"90",
x"03", x"E6", x"F5", x"18", x"E5", x"F4", x"49", x"FF",
x"85", x"F4", x"90", x"02", x"C6", x"F5", x"A5", x"F5",
x"0A", x"90", x"03", x"C6", x"F7", x"18", x"65", x"F6",
x"85", x"F6", x"90", x"02", x"E6", x"F7", x"A5", x"F5",
x"18", x"65", x"E4", x"85", x"E2", x"EA", x"EA", x"EA",
x"EA", x"A5", x"F7", x"18", x"65", x"E5", x"EA", x"EA",
x"EA", x"EA", x"85", x"E3", x"20", x"69", x"FE", x"88",
x"D0", x"C2", x"CA", x"D0", x"BF", x"A5", x"E4", x"85",
x"E2", x"A5", x"E5", x"85", x"E3", x"68", x"A8", x"68",
x"AA", x"60", x"48", x"8A", x"48", x"98", x"48", x"D8",
x"BA", x"BD", x"04", x"01", x"29", x"10", x"D0", x"06",
x"6C", x"1E", x"02", x"6C", x"20", x"02", x"6C", x"22",
x"02", x"78", x"D8", x"A2", x"FF", x"9A", x"A2", x"0F",
x"BD", x"8C", x"E6", x"95", x"E0", x"CA", x"10", x"F8",
x"20", x"B0", x"EE", x"A9", x"0C", x"20", x"F1", x"FF",
x"EA", x"EA", x"EA", x"A0", x"84", x"A9", x"E6", x"20",
x"3B", x"E6", x"20", x"57", x"E6", x"A2", x"00", x"20",
x"33", x"E6", x"E8", x"C9", x"0D", x"F0", x"EC", x"A0",
x"FF", x"C8", x"B9", x"00", x"E7", x"C9", x"FF", x"F0",
x"17", x"DD", x"7F", x"02", x"D0", x"F3", x"98", x"0A",
x"A8", x"B9", x"C8", x"E6", x"85", x"F6", x"B9", x"C9",
x"E6", x"85", x"F7", x"20", x"0B", x"E9", x"90", x"CB",
x"20", x"F4", x"E4", x"20", x"F6", x"E7", x"A9", x"3F",
x"20", x"F1", x"FF", x"38", x"B0", x"BD", x"FF", x"FF",
x"6C", x"FE", x"00", x"6C", x"14", x"02", x"6C", x"16",
x"02", x"6C", x"18", x"02", x"6C", x"1A", x"02", x"6C",
x"1C", x"02", x"83", x"FF", x"89", x"FF", x"72", x"FF"
	);
begin
	process(clk)
	begin
		if rising_edge(clk) then
			data <= romData(conv_integer(addr));
		end if;
	end process;
end architecture;

