library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity guzzler_big_sprite_tile_bit1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of guzzler_big_sprite_tile_bit1 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"1F",X"3F",X"3F",X"3F",X"3F",X"1F",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"FC",X"FC",X"FC",X"FC",X"F8",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0D",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"60",X"E0",X"F0",X"F0",X"F8",X"FC",X"FE",X"0F",
		X"C0",X"80",X"80",X"80",X"80",X"80",X"C0",X"40",X"0C",X"FF",X"FC",X"F8",X"F0",X"E0",X"C0",X"40",
		X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",
		X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",
		X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"3F",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",
		X"60",X"40",X"C0",X"80",X"80",X"80",X"C0",X"60",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"1F",X"30",
		X"0C",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",
		X"0C",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",
		X"C0",X"70",X"1C",X"07",X"01",X"00",X"00",X"00",X"06",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"1F",X"30",X"20",X"30",X"18",X"0C",X"F8",X"8F",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"1F",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"E0",X"3C",X"0F",X"0C",X"0F",X"FF",X"FF",X"1F",X"03",X"00",X"00",X"00",
		X"CE",X"8C",X"08",X"08",X"08",X"0C",X"0C",X"0E",X"08",X"FC",X"FE",X"FF",X"7F",X"7F",X"7F",X"4F",
		X"0E",X"0F",X"0C",X"0C",X"0F",X"0E",X"0C",X"08",X"08",X"0C",X"0F",X"0E",X"0C",X"08",X"08",X"0C",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"0D",X"0F",X"0E",X"0C",X"0C",X"08",X"08",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"00",X"81",X"FF",X"0E",X"0C",X"0C",X"08",X"08",
		X"FC",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"0C",X"0C",X"0E",X"0F",X"0D",X"0C",X"8C",
		X"0F",X"FE",X"FC",X"FC",X"F8",X"F8",X"F8",X"08",X"0F",X"0E",X"0C",X"08",X"08",X"08",X"08",X"0D",
		X"0C",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"0C",X"0C",X"0C",X"0F",X"0E",X"0C",X"08",X"08",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"3F",X"83",X"FF",X"FF",X"FF",X"FF",X"3F",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"FF",X"F8",X"C0",X"00",
		X"00",X"FE",X"03",X"00",X"F0",X"1F",X"01",X"00",X"01",X"01",X"FD",X"07",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"F9",X"0F",X"03",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"F8",X"0E",X"03",X"01",X"00",X"00",X"00",
		X"07",X"80",X"F8",X"0F",X"00",X"00",X"00",X"00",X"18",X"0C",X"07",X"01",X"00",X"C0",X"70",X"1C",
		X"01",X"00",X"00",X"1F",X"3F",X"3F",X"3F",X"30",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"80",X"E0",X"F8",X"0C",X"3F",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"0D",X"FF",X"FF",X"FF",X"FF",X"FE",X"F8",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FC",X"8E",X"0F",X"00",X"00",X"00",X"FF",X"80",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"0D",X"0C",X"0C",X"FC",X"1F",X"0F",X"0D",X"0C",X"FC",X"1F",X"00",X"00",X"00",
		X"1C",X"0C",X"06",X"03",X"F0",X"98",X"0C",X"0E",X"0F",X"0D",X"0C",X"0C",X"8C",X"CC",X"6C",X"3C",
		X"1C",X"0C",X"06",X"03",X"F0",X"98",X"0C",X"0E",X"00",X"00",X"00",X"00",X"80",X"FC",X"6F",X"3C",
		X"80",X"F8",X"0F",X"CC",X"7F",X"00",X"00",X"00",X"08",X"08",X"18",X"F0",X"00",X"00",X"01",X"00",
		X"E0",X"3F",X"0F",X"07",X"C3",X"F1",X"F9",X"08",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"3F",X"7F",X"7F",X"7F",X"7F",X"7F",X"3C",X"FC",X"06",X"03",X"01",X"01",X"01",X"01",X"03",
		X"00",X"00",X"00",X"00",X"00",X"07",X"7C",X"C0",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"C0",X"40",X"40",X"C0",X"80",X"00",X"80",X"C0",X"40",X"C0",X"F8",X"0F",X"00",
		X"20",X"20",X"60",X"C0",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"60",X"2F",X"38",X"30",X"20",
		X"20",X"20",X"60",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"18",X"F0",X"20",
		X"31",X"10",X"F0",X"30",X"E0",X"00",X"00",X"00",X"78",X"00",X"00",X"00",X"00",X"00",X"F8",X"6F",
		X"00",X"FF",X"E3",X"F0",X"F8",X"F8",X"F8",X"F8",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"06",X"0C",X"1C",X"FC",X"8C",X"0C",X"0C",X"3C",X"0F",X"07",X"03",X"01",X"01",X"01",X"01",
		X"03",X"01",X"01",X"01",X"F3",X"9E",X"CC",X"6C",X"01",X"03",X"03",X"07",X"FF",X"1F",X"0F",X"06",
		X"1C",X"0C",X"06",X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"03",X"02",X"02",X"06",X"8C",X"FC",
		X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"03",X"02",X"FA",X"0E",X"06",X"02",
		X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"03",X"02",X"06",X"FC",X"04",X"06",X"02",
		X"FC",X"3C",X"0C",X"06",X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"03",X"06",X"0C",
		X"06",X"FF",X"FF",X"7F",X"1F",X"07",X"03",X"01",X"FC",X"06",X"03",X"01",X"01",X"01",X"01",X"03",
		X"4C",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0C",X"7E",X"3C",X"1C",X"0C",X"1C",X"3C",X"7E",X"0C",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"20",X"30",X"10",X"18",X"0C",X"06",X"03",
		X"C0",X"80",X"80",X"80",X"80",X"80",X"C0",X"40",X"00",X"07",X"0C",X"18",X"30",X"60",X"40",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"60",X"40",X"C0",X"80",X"80",X"80",X"C0",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"70",X"1C",X"07",X"01",X"00",X"00",X"00",X"06",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"1F",X"30",X"20",X"30",X"18",X"0C",X"F8",X"8F",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"E0",X"3C",X"07",X"00",X"03",X"80",X"F0",X"1E",X"03",X"00",X"00",X"00",
		X"C6",X"8C",X"08",X"08",X"08",X"0C",X"04",X"06",X"08",X"0C",X"86",X"C3",X"41",X"40",X"41",X"43",
		X"06",X"03",X"00",X"00",X"03",X"06",X"0C",X"08",X"08",X"0C",X"07",X"06",X"0C",X"08",X"08",X"0C",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"0F",X"0F",X"07",X"06",X"04",X"0C",X"08",X"08",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"81",X"FF",X"07",X"07",X"0F",X"0F",X"0F",
		X"F8",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"07",X"07",X"03",X"01",X"00",X"80",
		X"07",X"07",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"03",X"06",X"0C",X"08",X"08",X"08",X"08",X"0D",
		X"0C",X"04",X"06",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"03",X"06",X"0C",X"08",X"08",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"3F",X"83",X"FE",X"00",X"00",X"E0",X"3E",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"FF",X"78",X"C0",X"00",
		X"00",X"FE",X"03",X"00",X"F0",X"1F",X"01",X"00",X"01",X"01",X"FD",X"07",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"FF",X"FF",X"0F",X"03",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"F8",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"07",X"80",X"F8",X"0F",X"00",X"00",X"00",X"00",X"F8",X"FC",X"FF",X"FF",X"FF",X"FF",X"7F",X"1F",
		X"FF",X"FF",X"FF",X"FF",X"F1",X"E0",X"E0",X"F0",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"80",X"E0",X"38",X"0C",X"3F",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"01",X"00",X"00",X"01",X"03",X"0E",X"F8",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FC",X"86",X"03",X"00",X"00",X"00",X"FF",X"80",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"01",X"00",X"00",X"F0",X"1F",X"03",X"01",X"00",X"F0",X"1F",X"00",X"00",X"00",
		X"18",X"0C",X"06",X"03",X"F0",X"98",X"0C",X"06",X"03",X"01",X"00",X"00",X"80",X"C0",X"60",X"30",
		X"F8",X"FC",X"FE",X"FF",X"FF",X"9F",X"0F",X"07",X"00",X"00",X"00",X"00",X"80",X"FC",X"E7",X"F0",
		X"FF",X"FF",X"0F",X"C0",X"7F",X"00",X"00",X"00",X"0F",X"0F",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"E0",X"FF",X"FC",X"FE",X"FF",X"7F",X"1F",X"0F",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"3C",X"60",X"40",X"40",X"40",X"60",X"30",X"FC",X"06",X"03",X"01",X"01",X"01",X"01",X"03",
		X"00",X"00",X"00",X"00",X"00",X"07",X"7C",X"C0",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"C0",X"40",X"40",X"C0",X"80",X"00",X"80",X"C0",X"40",X"C0",X"F8",X"0F",X"00",
		X"20",X"20",X"60",X"C0",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"7F",X"3F",X"38",X"30",X"20",
		X"3F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"0F",X"1F",X"FF",X"3F",
		X"F1",X"F0",X"F0",X"30",X"E0",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",
		X"00",X"FF",X"7F",X"3F",X"1F",X"0F",X"8F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"06",X"0C",X"18",X"F0",X"80",X"00",X"00",X"38",X"0C",X"06",X"03",X"01",X"01",X"01",X"01",
		X"03",X"01",X"01",X"01",X"F3",X"9E",X"C0",X"60",X"01",X"03",X"02",X"06",X"FC",X"18",X"0C",X"06",
		X"18",X"0C",X"06",X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"03",X"02",X"02",X"06",X"8C",X"F8",
		X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"FF",X"FF",X"FF",X"FE",X"FE",X"0E",X"06",X"02",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"03",X"02",X"06",X"FC",X"FC",X"FE",X"FE",
		X"F8",X"38",X"0C",X"06",X"03",X"01",X"01",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",
		X"06",X"FC",X"C0",X"F0",X"FC",X"FE",X"FF",X"FF",X"FC",X"06",X"03",X"01",X"01",X"01",X"01",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"7B",X"7B",X"31",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"01",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"70",X"78",X"18",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"06",X"0F",X"0F",X"06",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"F0",
		X"00",X"00",X"00",X"18",X"3C",X"3C",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"78",X"78",X"30",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"1E",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DE",
		X"FE",X"FF",X"F9",X"79",X"3E",X"00",X"F8",X"FC",X"00",X"00",X"01",X"03",X"03",X"03",X"01",X"7C",
		X"32",X"1C",X"00",X"1F",X"0F",X"07",X"00",X"00",X"FE",X"E6",X"E6",X"FC",X"00",X"3E",X"7F",X"73",
		X"70",X"00",X"07",X"00",X"78",X"00",X"7C",X"FE",X"01",X"01",X"0F",X"1F",X"3F",X"7F",X"7C",X"78",
		X"03",X"00",X"3E",X"3F",X"3F",X"1F",X"0F",X"07",X"00",X"0F",X"1F",X"3F",X"3C",X"1C",X"0F",X"00",
		X"00",X"0F",X"1F",X"3F",X"3C",X"1C",X"0F",X"00",X"07",X"0F",X"1F",X"3F",X"3F",X"3E",X"00",X"1E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1E",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1E",X"3E",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1E",
		X"7C",X"3C",X"3C",X"3C",X"3C",X"3E",X"FE",X"FE",X"00",X"00",X"C0",X"E0",X"F0",X"F0",X"F8",X"F8",
		X"00",X"00",X"00",X"F8",X"F0",X"FC",X"FC",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"80",X"E0",X"E0",X"C0",X"80",X"C0",X"00",X"00",
		X"C0",X"00",X"30",X"70",X"FC",X"FC",X"F0",X"30",X"00",X"00",X"80",X"C0",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"80",X"C0",X"C0",X"80",X"00",X"00",X"30",X"F0",X"FC",X"FC",X"70",X"30",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"1E",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",
		X"07",X"07",X"07",X"07",X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"03",X"07",
		X"07",X"07",X"07",X"07",X"0F",X"03",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"07",
		X"07",X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"07",X"0F",X"07",X"07",X"07",
		X"03",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"07",X"07",X"07",X"07",X"07",X"07",
		X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"03",
		X"00",X"00",X"60",X"F0",X"F0",X"60",X"00",X"00",X"00",X"01",X"03",X"07",X"07",X"03",X"01",X"00",
		X"00",X"01",X"03",X"07",X"07",X"03",X"01",X"00",X"00",X"00",X"60",X"F0",X"F0",X"60",X"00",X"00",
		X"30",X"78",X"78",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"07",X"03",X"00",X"00",X"00",X"00",
		X"70",X"78",X"78",X"30",X"00",X"00",X"00",X"00",X"3E",X"3F",X"7C",X"5D",X"CE",X"87",X"C0",X"40",
		X"5F",X"7F",X"3F",X"3F",X"3E",X"3D",X"1D",X"3D",X"03",X"07",X"1F",X"33",X"60",X"C7",X"8F",X"DF",
		X"3C",X"3C",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"03",X"00",X"00",X"03",X"03",X"18",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7C",X"07",X"07",X"07",X"03",X"01",X"00",X"00",X"01",X"F0",X"F8",X"CD",X"CC",X"F8",X"F0",X"00",
		X"00",X"F0",X"F8",X"CC",X"CD",X"F8",X"F0",X"01",X"00",X"00",X"01",X"03",X"07",X"07",X"07",X"F0",
		X"61",X"61",X"03",X"07",X"07",X"03",X"03",X"01",X"30",X"01",X"30",X"09",X"0C",X"1C",X"01",X"61",
		X"7E",X"7E",X"7E",X"0C",X"0C",X"04",X"04",X"18",X"00",X"80",X"80",X"00",X"00",X"00",X"1C",X"3E",
		X"61",X"61",X"03",X"07",X"07",X"03",X"03",X"01",X"3E",X"FF",X"3E",X"CF",X"CE",X"1C",X"F9",X"61",
		X"FF",X"FF",X"FF",X"0F",X"EF",X"E7",X"E7",X"DF",X"00",X"80",X"80",X"1F",X"FF",X"FF",X"FF",X"FF",
		X"F1",X"EA",X"F4",X"DF",X"60",X"1F",X"00",X"00",X"01",X"07",X"07",X"98",X"81",X"81",X"01",X"7F",
		X"F8",X"18",X"31",X"71",X"31",X"20",X"C0",X"0C",X"01",X"03",X"03",X"01",X"00",X"00",X"70",X"F8",
		X"7C",X"FC",X"FC",X"F8",X"F0",X"E0",X"00",X"00",X"02",X"00",X"06",X"80",X"28",X"F8",X"7C",X"7C",
		X"7C",X"7C",X"F8",X"28",X"80",X"06",X"00",X"02",X"00",X"00",X"E0",X"F0",X"F8",X"FC",X"FC",X"7C",
		X"55",X"95",X"D4",X"F4",X"F0",X"F3",X"E7",X"C7",X"1E",X"9E",X"1E",X"9F",X"1F",X"FF",X"56",X"34",
		X"00",X"70",X"FC",X"FE",X"FE",X"7E",X"3E",X"1E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"95",X"D5",X"F4",X"F0",X"F3",X"E7",X"C7",X"3F",X"9F",X"1F",X"9F",X"1F",X"FF",X"57",X"35",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"41",X"C3",X"43",X"80",X"00",X"83",X"0F",X"0F",X"3C",X"78",X"F8",X"F0",X"F0",X"F0",X"B0",X"80",
		X"00",X"F0",X"FC",X"FE",X"FE",X"FE",X"7E",X"FC",X"80",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"07",X"07",X"07",X"07",X"06",X"0C",
		X"0C",X"06",X"07",X"07",X"07",X"07",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"C0",X"0C",X"3C",X"F8",X"F0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"3F",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"FC",X"FC",X"FC",X"F8",X"F0",X"C0",X"00",X"FE",X"FC",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",
		X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"00",X"00",X"00",X"C0",X"F0",X"F8",X"FC",X"FC",
		X"FE",X"F0",X"80",X"1C",X"FC",X"F8",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"1F",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3C",X"3C",X"18",X"00",X"00",X"00",X"00",X"00",X"73",X"EB",X"AB",X"A8",X"90",X"CB",X"67",X"3B",
		X"3F",X"3C",X"3B",X"17",X"36",X"75",X"7B",X"7F",X"03",X"06",X"04",X"05",X"07",X"0F",X"1F",X"3F",
		X"00",X"06",X"0F",X"0F",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3C",X"3C",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",
		X"00",X"30",X"78",X"78",X"30",X"00",X"00",X"00",X"1F",X"07",X"03",X"03",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"06",X"06",X"0F",X"1F",X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"01",X"01",X"18",X"3C",X"3C",X"18",
		X"60",X"30",X"19",X"0B",X"E7",X"3F",X"07",X"77",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E8",X"F5",X"F2",X"DF",X"60",X"1F",X"00",X"00",X"F1",X"E7",X"E7",X"F8",X"C1",X"C1",X"C1",X"FF",
		X"FF",X"1F",X"BF",X"7F",X"3F",X"38",X"F8",X"FC",X"FD",X"03",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7E",X"7F",X"3F",X"1F",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"01",X"01",X"35",X"3E",X"7E",
		X"7E",X"3E",X"35",X"01",X"01",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"1F",X"3F",X"7F",X"7E",
		X"3B",X"3B",X"11",X"00",X"00",X"00",X"00",X"00",X"80",X"A0",X"A0",X"80",X"80",X"88",X"7B",X"3B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"81",X"FE",X"FE",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"7D",X"7C",X"3C",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"F1",X"7D",
		X"00",X"00",X"80",X"80",X"C0",X"C0",X"80",X"00",X"FF",X"FF",X"3F",X"00",X"00",X"00",X"00",X"00",
		X"4F",X"DF",X"4F",X"87",X"01",X"83",X"0F",X"0F",X"3F",X"7F",X"FF",X"F3",X"F3",X"F3",X"B7",X"87",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"80",X"C0",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"3B",X"FC",X"FC",X"FC",X"F8",X"F0",X"00",X"00",X"78",X"E4",X"E6",X"FE",X"FE",X"FC",X"78",
		X"78",X"FC",X"FE",X"FE",X"E6",X"E4",X"78",X"00",X"00",X"00",X"F0",X"F8",X"FC",X"FC",X"38",X"07",
		X"F0",X"F0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"7F",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"F8",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F8",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"8F",X"8F",X"81",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FC",X"FC",X"FC",X"FC",X"F8",X"E0",X"00",X"FE",X"FC",X"FC",X"FC",X"FC",X"FE",X"FF",X"FF",
		X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"C0",X"F0",X"F8",X"FC",
		X"03",X"83",X"03",X"03",X"03",X"03",X"00",X"00",X"00",X"80",X"80",X"10",X"00",X"00",X"03",X"03",
		X"03",X"03",X"00",X"00",X"10",X"80",X"80",X"00",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"83",
		X"3E",X"7F",X"7F",X"0E",X"0E",X"0F",X"0F",X"06",X"18",X"3C",X"7C",X"7C",X"7C",X"3E",X"3E",X"1E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"3E",X"7F",X"7F",X"0E",X"1C",X"3C",X"3C",X"18",X"18",X"3C",X"7C",X"7C",X"7C",X"3E",X"3E",X"1E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"FC",X"FC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0C",X"1E",X"1E",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"3C",X"3C",X"18",X"00",X"00",X"00",X"00",
		X"33",X"7B",X"7B",X"31",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"01",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"70",X"78",X"18",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"18",X"3C",X"3C",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"78",X"78",X"30",X"00",X"00",
		X"F0",X"F0",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"60",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"06",X"0F",X"0F",X"06",X"00",X"00",X"00",X"00",
		X"06",X"00",X"01",X"03",X"03",X"01",X"00",X"00",X"1B",X"3E",X"F9",X"79",X"7E",X"3F",X"7F",X"36",
		X"1F",X"7F",X"79",X"39",X"3F",X"26",X"00",X"10",X"07",X"0F",X"0F",X"1F",X"1F",X"19",X"01",X"0B",
		X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"1E",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DE",
		X"F2",X"F3",X"FF",X"7F",X"3E",X"00",X"F8",X"E4",X"00",X"00",X"01",X"03",X"03",X"03",X"01",X"7C",
		X"03",X"00",X"3E",X"3F",X"3F",X"1F",X"0F",X"07",X"00",X"0F",X"1C",X"3C",X"3F",X"1F",X"0F",X"00",
		X"00",X"0F",X"1C",X"3C",X"3F",X"1F",X"0F",X"00",X"07",X"0F",X"1F",X"3F",X"3F",X"3E",X"00",X"1E",
		X"38",X"7C",X"7E",X"7F",X"7F",X"3F",X"1D",X"00",X"FF",X"7E",X"00",X"80",X"F0",X"00",X"03",X"00",
		X"F3",X"7F",X"3E",X"00",X"F2",X"F3",X"FF",X"FF",X"00",X"0F",X"1F",X"3F",X"3F",X"00",X"7E",X"F3",
		X"1F",X"3E",X"FC",X"FC",X"F8",X"E0",X"00",X"00",X"00",X"00",X"80",X"80",X"0A",X"1F",X"BF",X"1F",
		X"E0",X"80",X"80",X"01",X"B0",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"E0",X"F0",X"F0",X"E0",
		X"1E",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1E",X"3E",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1E",
		X"7C",X"3C",X"3C",X"3C",X"3C",X"3E",X"FE",X"FE",X"00",X"00",X"C0",X"E0",X"F0",X"F0",X"F8",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"F0",X"E0",X"F8",X"E0",X"78",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"FE",X"FE",X"F2",X"F8",X"00",X"F0",X"00",
		X"03",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"07",X"07",X"07",X"07",X"07",X"07",
		X"07",X"07",X"07",X"87",X"07",X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"03",
		X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"1E",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",
		X"07",X"07",X"07",X"07",X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"03",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"07",X"07",X"07",X"0F",X"07",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"07",
		X"07",X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"07",X"0F",X"07",X"07",X"07");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
