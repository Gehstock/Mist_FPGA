library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity CHEWINGGUM_ROM_PGM_0 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of CHEWINGGUM_ROM_PGM_0 is
	type rom is array(0 to  10239) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"C3",X"4A",X"00",X"BA",X"CA",X"69",X"B5",X"6E",X"C3",X"00",X"06",X"54",X"16",X"2A",X"6E",X"3A",
		X"C3",X"40",X"04",X"C2",X"AE",X"F5",X"09",X"C9",X"6A",X"BF",X"64",X"A5",X"7F",X"61",X"35",X"2A",
		X"0E",X"F6",X"78",X"BA",X"6E",X"1A",X"B2",X"4F",X"11",X"11",X"00",X"FF",X"19",X"FF",X"19",X"FF",
		X"19",X"FF",X"C9",X"BF",X"6A",X"15",X"98",X"E6",X"7E",X"2C",X"4E",X"77",X"06",X"07",X"2C",X"7E",
		X"71",X"2C",X"4E",X"77",X"10",X"F8",X"C9",X"BF",X"EA",X"AF",X"3E",X"FF",X"32",X"00",X"78",X"AF",
		X"21",X"00",X"58",X"77",X"2C",X"C2",X"53",X"00",X"2E",X"09",X"06",X"06",X"70",X"2E",X"0B",X"70",
		X"2E",X"39",X"70",X"2E",X"3D",X"00",X"2E",X"35",X"36",X"05",X"06",X"01",X"2E",X"0F",X"3E",X"33",
		X"70",X"2C",X"2C",X"BD",X"C2",X"70",X"00",X"21",X"00",X"50",X"3E",X"1C",X"06",X"04",X"77",X"2C",
		X"C2",X"7E",X"00",X"24",X"10",X"F8",X"11",X"20",X"00",X"21",X"04",X"51",X"06",X"10",X"3E",X"E0",
		X"77",X"3C",X"19",X"10",X"FB",X"21",X"05",X"51",X"06",X"10",X"77",X"3C",X"19",X"10",X"FB",X"21",
		X"DA",X"50",X"36",X"16",X"19",X"36",X"0E",X"19",X"36",X"10",X"19",X"36",X"0A",X"19",X"36",X"17",
		X"19",X"36",X"16",X"19",X"19",X"19",X"36",X"17",X"19",X"36",X"0E",X"19",X"36",X"0B",X"19",X"19",
		X"19",X"36",X"16",X"19",X"36",X"0D",X"19",X"36",X"0D",X"19",X"36",X"13",X"21",X"9C",X"51",X"36",
		X"1B",X"21",X"3C",X"52",X"36",X"1A",X"21",X"9E",X"51",X"36",X"17",X"19",X"36",X"0F",X"19",X"36",
		X"0D",X"19",X"36",X"0E",X"19",X"36",X"15",X"19",X"36",X"0C",X"31",X"00",X"44",X"21",X"A7",X"50",
		X"06",X"16",X"3E",X"D1",X"77",X"19",X"10",X"FC",X"21",X"B8",X"50",X"3E",X"D6",X"06",X"16",X"77",
		X"19",X"10",X"FC",X"21",X"88",X"50",X"11",X"B0",X"00",X"06",X"10",X"3E",X"D4",X"CD",X"44",X"01",
		X"19",X"06",X"10",X"CD",X"44",X"01",X"19",X"06",X"10",X"CD",X"44",X"01",X"19",X"06",X"10",X"CD",
		X"44",X"01",X"21",X"28",X"51",X"3E",X"D3",X"06",X"10",X"CD",X"44",X"01",X"19",X"06",X"10",X"CD",
		X"44",X"01",X"19",X"06",X"10",X"CD",X"44",X"01",X"19",X"06",X"10",X"CD",X"44",X"01",X"C3",X"50",
		X"01",X"FF",X"FF",X"FF",X"77",X"2C",X"10",X"FC",X"C9",X"C3",X"BA",X"CA",X"AF",X"F0",X"7A",X"6B",
		X"21",X"87",X"50",X"3E",X"D2",X"11",X"C0",X"00",X"77",X"19",X"77",X"19",X"77",X"19",X"77",X"21",
		X"98",X"50",X"3E",X"D7",X"77",X"19",X"77",X"19",X"77",X"19",X"77",X"21",X"27",X"51",X"3E",X"D0",
		X"77",X"19",X"77",X"19",X"77",X"19",X"77",X"21",X"38",X"51",X"3E",X"D5",X"77",X"19",X"77",X"19",
		X"77",X"19",X"77",X"21",X"6F",X"50",X"36",X"D8",X"2C",X"36",X"D9",X"21",X"8F",X"53",X"36",X"D8",
		X"2C",X"36",X"D9",X"21",X"8F",X"50",X"3E",X"DC",X"06",X"DD",X"77",X"2C",X"70",X"19",X"70",X"2D",
		X"77",X"19",X"77",X"2C",X"70",X"19",X"70",X"2D",X"77",X"C3",X"B0",X"01",X"FF",X"EA",X"26",X"5A",
		X"11",X"1D",X"00",X"3E",X"20",X"06",X"04",X"21",X"B2",X"50",X"CD",X"30",X"02",X"3E",X"20",X"06",
		X"04",X"21",X"72",X"51",X"CD",X"30",X"02",X"3E",X"20",X"06",X"04",X"21",X"F2",X"52",X"CD",X"30",
		X"02",X"3E",X"30",X"06",X"04",X"21",X"32",X"52",X"CD",X"30",X"02",X"3E",X"90",X"06",X"04",X"21",
		X"AE",X"50",X"CD",X"30",X"02",X"3E",X"90",X"06",X"04",X"21",X"6E",X"51",X"CD",X"30",X"02",X"3E",
		X"90",X"06",X"04",X"21",X"EE",X"52",X"CD",X"30",X"02",X"3E",X"60",X"06",X"04",X"21",X"AA",X"50",
		X"CD",X"30",X"02",X"3E",X"60",X"06",X"04",X"21",X"6A",X"51",X"CD",X"30",X"02",X"3E",X"60",X"06",
		X"04",X"21",X"EA",X"52",X"CD",X"30",X"02",X"3E",X"B0",X"06",X"04",X"21",X"2E",X"52",X"CD",X"30",
		X"02",X"3E",X"80",X"06",X"04",X"21",X"2A",X"52",X"CD",X"30",X"02",X"C3",X"40",X"02",X"FF",X"FF",
		X"77",X"3C",X"2C",X"77",X"3C",X"2C",X"77",X"3C",X"2C",X"77",X"3C",X"19",X"10",X"F2",X"C9",X"FF",
		X"11",X"1F",X"00",X"3E",X"A2",X"06",X"03",X"21",X"A8",X"50",X"CD",X"90",X"02",X"3E",X"B2",X"21",
		X"68",X"51",X"CD",X"90",X"02",X"3E",X"A2",X"21",X"28",X"52",X"CD",X"90",X"02",X"3E",X"A2",X"21",
		X"E8",X"52",X"CD",X"90",X"02",X"3E",X"B0",X"21",X"B6",X"50",X"CD",X"90",X"02",X"3E",X"B0",X"21",
		X"76",X"51",X"CD",X"90",X"02",X"3E",X"90",X"21",X"36",X"52",X"CD",X"90",X"02",X"3E",X"B0",X"21",
		X"F6",X"52",X"CD",X"90",X"02",X"3A",X"00",X"78",X"00",X"00",X"00",X"C3",X"B0",X"02",X"FF",X"FF",
		X"77",X"2C",X"3C",X"77",X"19",X"80",X"77",X"2C",X"3C",X"77",X"19",X"80",X"77",X"2C",X"3C",X"77",
		X"19",X"80",X"77",X"2C",X"3C",X"77",X"C9",X"7B",X"B6",X"E5",X"12",X"32",X"80",X"01",X"23",X"45",
		X"11",X"C0",X"00",X"21",X"2F",X"51",X"3E",X"DA",X"06",X"DB",X"77",X"2C",X"70",X"19",X"70",X"2D",
		X"77",X"19",X"77",X"2C",X"70",X"19",X"70",X"2D",X"77",X"AF",X"32",X"FE",X"50",X"32",X"1E",X"51",
		X"32",X"3E",X"51",X"32",X"5E",X"51",X"3A",X"00",X"78",X"AF",X"C3",X"00",X"03",X"01",X"23",X"45",
		X"67",X"89",X"AB",X"CD",X"EF",X"A6",X"3B",X"2D",X"66",X"BB",X"94",X"0A",X"D6",X"C7",X"C2",X"A5",
		X"BE",X"F6",X"37",X"B9",X"AE",X"68",X"2B",X"54",X"7B",X"F3",X"05",X"16",X"82",X"BE",X"69",X"BF",
		X"21",X"00",X"40",X"06",X"30",X"77",X"2C",X"10",X"FC",X"21",X"20",X"40",X"3E",X"16",X"77",X"2C",
		X"77",X"CD",X"00",X"08",X"C3",X"2B",X"03",X"32",X"20",X"40",X"21",X"00",X"70",X"46",X"3E",X"02",
		X"A0",X"C2",X"26",X"03",X"3E",X"17",X"C6",X"14",X"32",X"21",X"40",X"3E",X"01",X"32",X"02",X"60",
		X"21",X"3E",X"53",X"3E",X"1C",X"77",X"2E",X"5E",X"77",X"2E",X"7E",X"77",X"2E",X"9E",X"77",X"AF",
		X"32",X"FC",X"50",X"32",X"1C",X"51",X"32",X"3C",X"51",X"32",X"5C",X"51",X"32",X"DC",X"51",X"32",
		X"FC",X"51",X"32",X"7C",X"52",X"32",X"9C",X"52",X"32",X"BC",X"52",X"CF",X"3A",X"5E",X"51",X"FE",
		X"00",X"C2",X"80",X"03",X"3A",X"3E",X"51",X"FE",X"00",X"C2",X"80",X"03",X"3A",X"1E",X"51",X"FE",
		X"00",X"C2",X"80",X"03",X"3A",X"FE",X"50",X"FE",X"00",X"C2",X"80",X"03",X"C3",X"5B",X"03",X"FF",
		X"CF",X"3A",X"00",X"60",X"06",X"08",X"A0",X"C3",X"E4",X"06",X"21",X"20",X"40",X"46",X"21",X"10",
		X"40",X"4E",X"0C",X"3E",X"16",X"B9",X"CC",X"A0",X"03",X"71",X"C3",X"AF",X"03",X"FF",X"FF",X"FF",
		X"0E",X"00",X"11",X"11",X"40",X"1A",X"3C",X"B8",X"CC",X"AD",X"03",X"12",X"C9",X"AF",X"C9",X"D7",
		X"CF",X"21",X"00",X"60",X"46",X"3E",X"08",X"A0",X"CA",X"8A",X"03",X"CD",X"00",X"05",X"CF",X"21",
		X"00",X"60",X"46",X"3E",X"08",X"A0",X"C2",X"BB",X"03",X"CF",X"3A",X"00",X"60",X"06",X"10",X"A0",
		X"C3",X"D0",X"07",X"CF",X"21",X"21",X"40",X"46",X"21",X"13",X"40",X"0C",X"3E",X"16",X"B9",X"CC",
		X"E6",X"03",X"71",X"C3",X"F5",X"03",X"0E",X"00",X"11",X"12",X"40",X"1A",X"3C",X"B8",X"CC",X"F3",
		X"03",X"12",X"C9",X"AF",X"C9",X"21",X"00",X"60",X"46",X"3E",X"10",X"A0",X"C2",X"00",X"07",X"00",
		X"21",X"00",X"60",X"46",X"3E",X"08",X"A0",X"C2",X"BB",X"03",X"21",X"00",X"60",X"46",X"3E",X"06",
		X"A0",X"CA",X"D3",X"03",X"CF",X"CD",X"90",X"05",X"21",X"00",X"60",X"46",X"3E",X"06",X"A0",X"C2",
		X"14",X"04",X"21",X"FC",X"51",X"46",X"AF",X"B8",X"C2",X"D3",X"03",X"21",X"DC",X"51",X"46",X"B8",
		X"C2",X"D3",X"03",X"C3",X"5B",X"03",X"BA",X"CA",X"72",X"BF",X"64",X"29",X"1A",X"0A",X"BA",X"27",
		X"3A",X"00",X"60",X"E6",X"40",X"C8",X"11",X"20",X"00",X"06",X"03",X"21",X"1E",X"51",X"7E",X"B7",
		X"20",X"19",X"19",X"10",X"F9",X"3A",X"FE",X"50",X"C3",X"C5",X"04",X"47",X"AF",X"32",X"FE",X"50",
		X"21",X"02",X"60",X"CD",X"A1",X"04",X"10",X"FB",X"C3",X"C8",X"07",X"06",X"03",X"21",X"1E",X"51",
		X"35",X"F2",X"7A",X"04",X"3E",X"09",X"77",X"19",X"10",X"F6",X"21",X"3E",X"53",X"7E",X"FE",X"1C",
		X"20",X"07",X"06",X"04",X"AF",X"77",X"19",X"10",X"FB",X"21",X"5E",X"53",X"06",X"03",X"7E",X"3C",
		X"27",X"E6",X"0F",X"77",X"20",X"03",X"19",X"10",X"F5",X"21",X"01",X"60",X"CD",X"B3",X"04",X"18",
		X"9F",X"3E",X"01",X"21",X"00",X"60",X"77",X"CD",X"E6",X"04",X"AF",X"21",X"00",X"60",X"77",X"CD",
		X"E6",X"04",X"C9",X"3E",X"01",X"21",X"01",X"60",X"77",X"CD",X"E6",X"04",X"AF",X"21",X"01",X"60",
		X"77",X"CD",X"E6",X"04",X"C9",X"FE",X"00",X"CA",X"C8",X"07",X"32",X"3E",X"53",X"C3",X"5B",X"04",
		X"00",X"00",X"00",X"00",X"3E",X"00",X"32",X"01",X"60",X"CD",X"E6",X"04",X"3A",X"00",X"60",X"E6",
		X"40",X"C8",X"C3",X"46",X"04",X"FF",X"1E",X"0F",X"16",X"FF",X"CF",X"15",X"C2",X"EA",X"04",X"1D",
		X"C2",X"EA",X"04",X"C9",X"3A",X"26",X"15",X"00",X"6B",X"A9",X"2A",X"8E",X"BF",X"CF",X"2A",X"45",
		X"3A",X"5E",X"51",X"FE",X"00",X"C2",X"1E",X"05",X"3A",X"3E",X"51",X"FE",X"00",X"C2",X"1E",X"05",
		X"3A",X"1E",X"51",X"FE",X"00",X"C2",X"1E",X"05",X"3A",X"FE",X"50",X"FE",X"00",X"C8",X"CD",X"00",
		X"09",X"00",X"00",X"C8",X"3A",X"DC",X"51",X"3C",X"32",X"DC",X"51",X"FE",X"0A",X"C2",X"3C",X"05",
		X"3E",X"00",X"32",X"DC",X"51",X"3A",X"FC",X"51",X"3C",X"32",X"FC",X"51",X"3A",X"FE",X"50",X"3D",
		X"32",X"FE",X"50",X"00",X"00",X"00",X"00",X"FE",X"FF",X"C2",X"7A",X"05",X"3E",X"09",X"32",X"FE",
		X"50",X"3A",X"1E",X"51",X"3D",X"32",X"1E",X"51",X"FE",X"FF",X"C2",X"7A",X"05",X"3E",X"09",X"32",
		X"1E",X"51",X"3A",X"3E",X"51",X"3D",X"32",X"3E",X"51",X"FE",X"FF",X"C2",X"7A",X"05",X"3E",X"09",
		X"32",X"3E",X"51",X"3A",X"5E",X"51",X"3D",X"32",X"5E",X"51",X"CD",X"EC",X"07",X"1E",X"1F",X"16",
		X"FF",X"CF",X"15",X"C2",X"81",X"05",X"1D",X"C2",X"81",X"05",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3A",X"FC",X"51",X"FE",X"00",X"C2",X"9E",X"05",X"3A",X"DC",X"51",X"FE",X"00",X"C8",X"3A",X"DC",
		X"51",X"3D",X"32",X"DC",X"51",X"FE",X"FF",X"C2",X"B6",X"05",X"3E",X"09",X"32",X"DC",X"51",X"3A",
		X"FC",X"51",X"3D",X"32",X"FC",X"51",X"3A",X"FE",X"50",X"3C",X"32",X"FE",X"50",X"FE",X"0A",X"C2",
		X"F0",X"05",X"3E",X"00",X"32",X"FE",X"50",X"3A",X"1E",X"51",X"3C",X"32",X"1E",X"51",X"FE",X"0A",
		X"C2",X"F0",X"05",X"3E",X"00",X"32",X"1E",X"51",X"3A",X"3E",X"51",X"3C",X"32",X"3E",X"51",X"FE",
		X"0A",X"C2",X"F0",X"05",X"3E",X"00",X"32",X"3E",X"51",X"3A",X"5E",X"51",X"3C",X"32",X"5E",X"51",
		X"1E",X"1F",X"16",X"FF",X"CF",X"15",X"C2",X"F4",X"05",X"1D",X"C2",X"F4",X"05",X"C9",X"FF",X"FF",
		X"3A",X"00",X"78",X"3A",X"00",X"60",X"E6",X"01",X"CA",X"7D",X"06",X"1E",X"0F",X"06",X"FF",X"3A",
		X"00",X"78",X"10",X"FB",X"1D",X"C2",X"0F",X"06",X"3A",X"00",X"60",X"E6",X"01",X"CA",X"7D",X"06",
		X"3A",X"FE",X"50",X"3C",X"32",X"FE",X"50",X"FE",X"0A",X"C2",X"5A",X"06",X"3E",X"00",X"32",X"FE",
		X"50",X"3A",X"1E",X"51",X"3C",X"32",X"1E",X"51",X"FE",X"0A",X"C2",X"5A",X"06",X"3E",X"00",X"32",
		X"1E",X"51",X"3A",X"3E",X"51",X"3C",X"32",X"3E",X"51",X"FE",X"0A",X"C2",X"5A",X"06",X"3E",X"00",
		X"32",X"3E",X"51",X"3A",X"5E",X"51",X"3C",X"32",X"5E",X"51",X"3E",X"01",X"32",X"03",X"60",X"3A",
		X"00",X"78",X"3A",X"00",X"60",X"E6",X"01",X"C2",X"5F",X"06",X"1E",X"0F",X"06",X"FF",X"3A",X"00",
		X"78",X"10",X"FB",X"1D",X"C2",X"6E",X"06",X"3E",X"00",X"32",X"03",X"60",X"C9",X"3A",X"00",X"60",
		X"E6",X"80",X"C8",X"1E",X"0F",X"06",X"FF",X"3A",X"00",X"78",X"10",X"FB",X"1D",X"C2",X"87",X"06",
		X"3A",X"00",X"60",X"E6",X"80",X"C8",X"00",X"00",X"3A",X"1E",X"51",X"3C",X"32",X"1E",X"51",X"FE",
		X"0A",X"C2",X"C1",X"06",X"3E",X"00",X"32",X"1E",X"51",X"3A",X"3E",X"51",X"3C",X"32",X"3E",X"51",
		X"FE",X"0A",X"C2",X"C1",X"06",X"3E",X"00",X"32",X"3E",X"51",X"3A",X"5E",X"51",X"3C",X"32",X"5E",
		X"51",X"3E",X"00",X"32",X"00",X"60",X"3A",X"00",X"78",X"3A",X"00",X"60",X"E6",X"80",X"C2",X"C6",
		X"06",X"1E",X"0F",X"06",X"FF",X"3A",X"00",X"78",X"10",X"FB",X"1D",X"C2",X"D5",X"06",X"3E",X"00",
		X"32",X"00",X"60",X"C9",X"C2",X"80",X"03",X"1E",X"0F",X"06",X"FF",X"3A",X"00",X"78",X"10",X"FB",
		X"1D",X"C2",X"EB",X"06",X"3A",X"00",X"60",X"06",X"08",X"A0",X"C2",X"80",X"03",X"C3",X"8A",X"03",
		X"CD",X"19",X"08",X"00",X"00",X"00",X"3A",X"09",X"40",X"32",X"31",X"40",X"3A",X"0A",X"40",X"32",
		X"32",X"40",X"3A",X"0B",X"40",X"32",X"33",X"40",X"78",X"32",X"3A",X"40",X"CD",X"60",X"21",X"CD",
		X"2A",X"23",X"20",X"F8",X"CD",X"78",X"23",X"CD",X"60",X"21",X"3A",X"30",X"40",X"21",X"10",X"40",
		X"46",X"B8",X"C2",X"27",X"07",X"CD",X"81",X"23",X"CD",X"60",X"22",X"3A",X"11",X"40",X"FE",X"16",
		X"DA",X"45",X"07",X"D6",X"16",X"47",X"3A",X"31",X"40",X"FE",X"16",X"DA",X"50",X"07",X"D6",X"16",
		X"B8",X"C2",X"38",X"07",X"CD",X"8A",X"23",X"CD",X"D0",X"22",X"3A",X"12",X"40",X"FE",X"16",X"DA",
		X"64",X"07",X"D6",X"16",X"47",X"3A",X"32",X"40",X"FE",X"16",X"DA",X"6F",X"07",X"D6",X"16",X"B8",
		X"C2",X"57",X"07",X"CD",X"F7",X"26",X"CD",X"30",X"23",X"3A",X"33",X"40",X"21",X"13",X"40",X"46",
		X"B8",X"C2",X"76",X"07",X"CD",X"80",X"23",X"3A",X"30",X"40",X"C6",X"30",X"6F",X"26",X"20",X"7E",
		X"32",X"40",X"40",X"3A",X"31",X"40",X"C6",X"30",X"6F",X"26",X"21",X"7E",X"32",X"41",X"40",X"3A",
		X"32",X"40",X"C6",X"30",X"6F",X"26",X"22",X"7E",X"32",X"42",X"40",X"3A",X"33",X"40",X"C6",X"30",
		X"6F",X"26",X"20",X"7E",X"32",X"43",X"40",X"00",X"00",X"00",X"C3",X"90",X"23",X"FF",X"FF",X"FF",
		X"3A",X"3A",X"40",X"3D",X"32",X"3A",X"40",X"C9",X"F1",X"C3",X"5B",X"03",X"FF",X"FF",X"FF",X"FF",
		X"C2",X"C9",X"03",X"1E",X"0F",X"06",X"FF",X"3A",X"00",X"78",X"10",X"FB",X"1D",X"C2",X"D7",X"07",
		X"3A",X"00",X"60",X"06",X"10",X"A0",X"C2",X"C9",X"03",X"C3",X"D3",X"03",X"3E",X"3F",X"32",X"00",
		X"78",X"16",X"FF",X"CF",X"1D",X"C2",X"F3",X"07",X"3E",X"FF",X"32",X"00",X"78",X"C9",X"FF",X"FF",
		X"21",X"00",X"70",X"46",X"3E",X"03",X"A0",X"32",X"22",X"40",X"32",X"24",X"40",X"3E",X"0C",X"A0",
		X"1F",X"1F",X"32",X"23",X"40",X"32",X"25",X"40",X"C9",X"3A",X"08",X"40",X"32",X"30",X"40",X"3A",
		X"10",X"40",X"C6",X"30",X"16",X"20",X"5F",X"1A",X"32",X"00",X"40",X"3A",X"11",X"40",X"C6",X"30",
		X"16",X"21",X"5F",X"1A",X"32",X"01",X"40",X"3A",X"12",X"40",X"C6",X"30",X"16",X"22",X"5F",X"1A",
		X"32",X"02",X"40",X"3A",X"13",X"40",X"C6",X"30",X"16",X"20",X"5F",X"1A",X"32",X"03",X"40",X"00",
		X"3A",X"00",X"40",X"21",X"01",X"40",X"46",X"B8",X"20",X"35",X"3A",X"02",X"40",X"B8",X"20",X"69",
		X"21",X"03",X"40",X"46",X"B8",X"20",X"37",X"3A",X"22",X"40",X"E6",X"03",X"C8",X"3A",X"24",X"40",
		X"E6",X"03",X"20",X"07",X"3A",X"22",X"40",X"32",X"24",X"40",X"C9",X"3D",X"32",X"24",X"40",X"3A",
		X"11",X"40",X"3C",X"FE",X"16",X"20",X"04",X"3A",X"11",X"40",X"3D",X"32",X"11",X"40",X"C9",X"21",
		X"02",X"40",X"46",X"3A",X"00",X"40",X"B8",X"20",X"28",X"3A",X"03",X"40",X"B8",X"C0",X"3A",X"23",
		X"40",X"E6",X"03",X"C8",X"3A",X"25",X"40",X"E6",X"03",X"28",X"3E",X"3D",X"32",X"25",X"40",X"00",
		X"00",X"3A",X"12",X"40",X"3C",X"FE",X"16",X"20",X"04",X"3A",X"12",X"40",X"3D",X"32",X"12",X"40",
		X"C9",X"3A",X"01",X"40",X"B8",X"C0",X"C3",X"99",X"08",X"21",X"01",X"40",X"46",X"3A",X"03",X"40",
		X"B8",X"C0",X"3A",X"23",X"40",X"E6",X"03",X"C8",X"3A",X"25",X"40",X"00",X"E6",X"03",X"28",X"09",
		X"3D",X"32",X"25",X"40",X"00",X"00",X"C3",X"7F",X"08",X"3A",X"23",X"40",X"32",X"25",X"40",X"C9",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3A",X"00",X"68",X"E6",X"80",X"20",X"0D",X"3A",X"00",X"68",X"E6",X"40",X"20",X"0C",X"3A",X"FC",
		X"51",X"FE",X"02",X"C9",X"3A",X"FC",X"51",X"FE",X"01",X"C9",X"3A",X"DC",X"51",X"FE",X"06",X"C9",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C3",X"4A",X"00",X"BA",X"CA",X"69",X"B5",X"6E",X"C3",X"00",X"06",X"54",X"16",X"2A",X"6E",X"3A",
		X"C3",X"40",X"04",X"C2",X"AE",X"F5",X"09",X"C9",X"6A",X"BF",X"64",X"A5",X"7F",X"61",X"35",X"2A",
		X"0E",X"F6",X"78",X"BA",X"6E",X"1A",X"B2",X"4F",X"11",X"11",X"00",X"FF",X"19",X"FF",X"19",X"FF",
		X"19",X"FF",X"C9",X"BF",X"6A",X"15",X"98",X"E6",X"7E",X"2C",X"4E",X"77",X"06",X"07",X"2C",X"7E",
		X"71",X"2C",X"4E",X"77",X"10",X"F8",X"C9",X"BF",X"EA",X"AF",X"3E",X"FF",X"32",X"00",X"78",X"AF",
		X"21",X"00",X"58",X"77",X"2C",X"C2",X"53",X"00",X"2E",X"09",X"06",X"06",X"70",X"2E",X"0B",X"70",
		X"2E",X"39",X"70",X"2E",X"3D",X"00",X"2E",X"35",X"36",X"05",X"06",X"01",X"2E",X"0F",X"3E",X"33",
		X"70",X"2C",X"2C",X"BD",X"C2",X"70",X"00",X"21",X"00",X"50",X"3E",X"1C",X"06",X"04",X"77",X"2C",
		X"C2",X"7E",X"00",X"24",X"10",X"F8",X"11",X"20",X"00",X"21",X"04",X"51",X"06",X"10",X"3E",X"E0",
		X"77",X"3C",X"19",X"10",X"FB",X"21",X"05",X"51",X"06",X"10",X"77",X"3C",X"19",X"10",X"FB",X"21",
		X"DA",X"50",X"36",X"16",X"19",X"36",X"0E",X"19",X"36",X"10",X"19",X"36",X"0A",X"19",X"36",X"17",
		X"19",X"36",X"16",X"19",X"19",X"19",X"36",X"17",X"19",X"36",X"0E",X"19",X"36",X"0B",X"19",X"19",
		X"19",X"36",X"16",X"19",X"36",X"0D",X"19",X"36",X"0D",X"19",X"36",X"13",X"21",X"9C",X"51",X"36",
		X"1B",X"21",X"3C",X"52",X"36",X"1A",X"21",X"9E",X"51",X"36",X"17",X"19",X"36",X"0F",X"19",X"36",
		X"0D",X"19",X"36",X"0E",X"19",X"36",X"15",X"19",X"36",X"0C",X"31",X"00",X"44",X"21",X"A7",X"50",
		X"06",X"16",X"3E",X"D1",X"77",X"19",X"10",X"FC",X"21",X"B8",X"50",X"3E",X"D6",X"06",X"16",X"77",
		X"19",X"10",X"FC",X"21",X"88",X"50",X"11",X"B0",X"00",X"06",X"10",X"3E",X"D4",X"CD",X"44",X"01",
		X"19",X"06",X"10",X"CD",X"44",X"01",X"19",X"06",X"10",X"CD",X"44",X"01",X"19",X"06",X"10",X"CD",
		X"44",X"01",X"21",X"28",X"51",X"3E",X"D3",X"06",X"10",X"CD",X"44",X"01",X"19",X"06",X"10",X"CD",
		X"44",X"01",X"19",X"06",X"10",X"CD",X"44",X"01",X"19",X"06",X"10",X"CD",X"44",X"01",X"C3",X"50",
		X"01",X"FF",X"FF",X"FF",X"77",X"2C",X"10",X"FC",X"C9",X"C3",X"BA",X"CA",X"AF",X"F0",X"7A",X"6B",
		X"21",X"87",X"50",X"3E",X"D2",X"11",X"C0",X"00",X"77",X"19",X"77",X"19",X"77",X"19",X"77",X"21",
		X"98",X"50",X"3E",X"D7",X"77",X"19",X"77",X"19",X"77",X"19",X"77",X"21",X"27",X"51",X"3E",X"D0",
		X"77",X"19",X"77",X"19",X"77",X"19",X"77",X"21",X"38",X"51",X"3E",X"D5",X"77",X"19",X"77",X"19",
		X"77",X"19",X"77",X"21",X"6F",X"50",X"36",X"D8",X"2C",X"36",X"D9",X"21",X"8F",X"53",X"36",X"D8",
		X"2C",X"36",X"D9",X"21",X"8F",X"50",X"3E",X"DC",X"06",X"DD",X"77",X"2C",X"70",X"19",X"70",X"2D",
		X"77",X"19",X"77",X"2C",X"70",X"19",X"70",X"2D",X"77",X"C3",X"B0",X"01",X"FF",X"EA",X"26",X"5A",
		X"11",X"1D",X"00",X"3E",X"20",X"06",X"04",X"21",X"B2",X"50",X"CD",X"30",X"02",X"3E",X"20",X"06",
		X"04",X"21",X"72",X"51",X"CD",X"30",X"02",X"3E",X"20",X"06",X"04",X"21",X"F2",X"52",X"CD",X"30",
		X"02",X"3E",X"30",X"06",X"04",X"21",X"32",X"52",X"CD",X"30",X"02",X"3E",X"90",X"06",X"04",X"21",
		X"AE",X"50",X"CD",X"30",X"02",X"3E",X"90",X"06",X"04",X"21",X"6E",X"51",X"CD",X"30",X"02",X"3E",
		X"90",X"06",X"04",X"21",X"EE",X"52",X"CD",X"30",X"02",X"3E",X"60",X"06",X"04",X"21",X"AA",X"50",
		X"CD",X"30",X"02",X"3E",X"60",X"06",X"04",X"21",X"6A",X"51",X"CD",X"30",X"02",X"3E",X"60",X"06",
		X"04",X"21",X"EA",X"52",X"CD",X"30",X"02",X"3E",X"B0",X"06",X"04",X"21",X"2E",X"52",X"CD",X"30",
		X"02",X"3E",X"80",X"06",X"04",X"21",X"2A",X"52",X"CD",X"30",X"02",X"C3",X"40",X"02",X"FF",X"FF",
		X"77",X"3C",X"2C",X"77",X"3C",X"2C",X"77",X"3C",X"2C",X"77",X"3C",X"19",X"10",X"F2",X"C9",X"FF",
		X"11",X"1F",X"00",X"3E",X"A2",X"06",X"03",X"21",X"A8",X"50",X"CD",X"90",X"02",X"3E",X"B2",X"21",
		X"68",X"51",X"CD",X"90",X"02",X"3E",X"A2",X"21",X"28",X"52",X"CD",X"90",X"02",X"3E",X"A2",X"21",
		X"E8",X"52",X"CD",X"90",X"02",X"3E",X"B0",X"21",X"B6",X"50",X"CD",X"90",X"02",X"3E",X"B0",X"21",
		X"76",X"51",X"CD",X"90",X"02",X"3E",X"90",X"21",X"36",X"52",X"CD",X"90",X"02",X"3E",X"B0",X"21",
		X"F6",X"52",X"CD",X"90",X"02",X"3A",X"00",X"78",X"00",X"00",X"00",X"C3",X"B0",X"02",X"FF",X"FF",
		X"77",X"2C",X"3C",X"77",X"19",X"80",X"77",X"2C",X"3C",X"77",X"19",X"80",X"77",X"2C",X"3C",X"77",
		X"19",X"80",X"77",X"2C",X"3C",X"77",X"C9",X"7B",X"B6",X"E5",X"12",X"32",X"80",X"01",X"23",X"45",
		X"11",X"C0",X"00",X"21",X"2F",X"51",X"3E",X"DA",X"06",X"DB",X"77",X"2C",X"70",X"19",X"70",X"2D",
		X"77",X"19",X"77",X"2C",X"70",X"19",X"70",X"2D",X"77",X"AF",X"32",X"FE",X"50",X"32",X"1E",X"51",
		X"32",X"3E",X"51",X"32",X"5E",X"51",X"3A",X"00",X"78",X"AF",X"C3",X"00",X"03",X"01",X"23",X"45",
		X"67",X"89",X"AB",X"CD",X"EF",X"A6",X"3B",X"2D",X"66",X"BB",X"94",X"0A",X"D6",X"C7",X"C2",X"A5",
		X"BE",X"F6",X"37",X"B9",X"AE",X"68",X"2B",X"54",X"7B",X"F3",X"05",X"16",X"82",X"BE",X"69",X"BF",
		X"21",X"00",X"40",X"06",X"30",X"77",X"2C",X"10",X"FC",X"21",X"20",X"40",X"3E",X"16",X"77",X"2C",
		X"77",X"CD",X"00",X"08",X"C3",X"2B",X"03",X"32",X"20",X"40",X"21",X"00",X"70",X"46",X"3E",X"02",
		X"A0",X"C2",X"26",X"03",X"3E",X"17",X"C6",X"14",X"32",X"21",X"40",X"3E",X"01",X"32",X"02",X"60",
		X"21",X"3E",X"53",X"3E",X"1C",X"77",X"2E",X"5E",X"77",X"2E",X"7E",X"77",X"2E",X"9E",X"77",X"AF",
		X"32",X"FC",X"50",X"32",X"1C",X"51",X"32",X"3C",X"51",X"32",X"5C",X"51",X"32",X"DC",X"51",X"32",
		X"FC",X"51",X"32",X"7C",X"52",X"32",X"9C",X"52",X"32",X"BC",X"52",X"CF",X"3A",X"5E",X"51",X"FE",
		X"00",X"C2",X"80",X"03",X"3A",X"3E",X"51",X"FE",X"00",X"C2",X"80",X"03",X"3A",X"1E",X"51",X"FE",
		X"00",X"C2",X"80",X"03",X"3A",X"FE",X"50",X"FE",X"00",X"C2",X"80",X"03",X"C3",X"5B",X"03",X"FF",
		X"CF",X"3A",X"00",X"60",X"06",X"08",X"A0",X"C3",X"E4",X"06",X"21",X"20",X"40",X"46",X"21",X"10",
		X"40",X"4E",X"0C",X"3E",X"16",X"B9",X"CC",X"A0",X"03",X"71",X"C3",X"AF",X"03",X"FF",X"FF",X"FF",
		X"0E",X"00",X"11",X"11",X"40",X"1A",X"3C",X"B8",X"CC",X"AD",X"03",X"12",X"C9",X"AF",X"C9",X"D7",
		X"CF",X"21",X"00",X"60",X"46",X"3E",X"08",X"A0",X"CA",X"8A",X"03",X"CD",X"00",X"05",X"CF",X"21",
		X"00",X"60",X"46",X"3E",X"08",X"A0",X"C2",X"BB",X"03",X"CF",X"3A",X"00",X"60",X"06",X"10",X"A0",
		X"C3",X"D0",X"07",X"CF",X"21",X"21",X"40",X"46",X"21",X"13",X"40",X"0C",X"3E",X"16",X"B9",X"CC",
		X"E6",X"03",X"71",X"C3",X"F5",X"03",X"0E",X"00",X"11",X"12",X"40",X"1A",X"3C",X"B8",X"CC",X"F3",
		X"03",X"12",X"C9",X"AF",X"C9",X"21",X"00",X"60",X"46",X"3E",X"10",X"A0",X"C2",X"00",X"07",X"00",
		X"21",X"00",X"60",X"46",X"3E",X"08",X"A0",X"C2",X"BB",X"03",X"21",X"00",X"60",X"46",X"3E",X"06",
		X"A0",X"CA",X"D3",X"03",X"CF",X"CD",X"90",X"05",X"21",X"00",X"60",X"46",X"3E",X"06",X"A0",X"C2",
		X"14",X"04",X"21",X"FC",X"51",X"46",X"AF",X"B8",X"C2",X"D3",X"03",X"21",X"DC",X"51",X"46",X"B8",
		X"C2",X"D3",X"03",X"C3",X"5B",X"03",X"BA",X"CA",X"72",X"BF",X"64",X"29",X"1A",X"0A",X"BA",X"27",
		X"3A",X"00",X"60",X"E6",X"40",X"C8",X"11",X"20",X"00",X"06",X"03",X"21",X"1E",X"51",X"7E",X"B7",
		X"20",X"19",X"19",X"10",X"F9",X"3A",X"FE",X"50",X"C3",X"C5",X"04",X"47",X"AF",X"32",X"FE",X"50",
		X"21",X"02",X"60",X"CD",X"A1",X"04",X"10",X"FB",X"C3",X"C8",X"07",X"06",X"03",X"21",X"1E",X"51",
		X"35",X"F2",X"7A",X"04",X"3E",X"09",X"77",X"19",X"10",X"F6",X"21",X"3E",X"53",X"7E",X"FE",X"1C",
		X"20",X"07",X"06",X"04",X"AF",X"77",X"19",X"10",X"FB",X"21",X"5E",X"53",X"06",X"03",X"7E",X"3C",
		X"27",X"E6",X"0F",X"77",X"20",X"03",X"19",X"10",X"F5",X"21",X"01",X"60",X"CD",X"B3",X"04",X"18",
		X"9F",X"3E",X"01",X"21",X"00",X"60",X"77",X"CD",X"E6",X"04",X"AF",X"21",X"00",X"60",X"77",X"CD",
		X"E6",X"04",X"C9",X"3E",X"01",X"21",X"01",X"60",X"77",X"CD",X"E6",X"04",X"AF",X"21",X"01",X"60",
		X"77",X"CD",X"E6",X"04",X"C9",X"FE",X"00",X"CA",X"C8",X"07",X"32",X"3E",X"53",X"C3",X"5B",X"04",
		X"00",X"00",X"00",X"00",X"3E",X"00",X"32",X"01",X"60",X"CD",X"E6",X"04",X"3A",X"00",X"60",X"E6",
		X"40",X"C8",X"C3",X"46",X"04",X"FF",X"1E",X"0F",X"16",X"FF",X"CF",X"15",X"C2",X"EA",X"04",X"1D",
		X"C2",X"EA",X"04",X"C9",X"3A",X"26",X"15",X"00",X"6B",X"A9",X"2A",X"8E",X"BF",X"CF",X"2A",X"45",
		X"3A",X"5E",X"51",X"FE",X"00",X"C2",X"1E",X"05",X"3A",X"3E",X"51",X"FE",X"00",X"C2",X"1E",X"05",
		X"3A",X"1E",X"51",X"FE",X"00",X"C2",X"1E",X"05",X"3A",X"FE",X"50",X"FE",X"00",X"C8",X"CD",X"00",
		X"09",X"00",X"00",X"C8",X"3A",X"DC",X"51",X"3C",X"32",X"DC",X"51",X"FE",X"0A",X"C2",X"3C",X"05",
		X"3E",X"00",X"32",X"DC",X"51",X"3A",X"FC",X"51",X"3C",X"32",X"FC",X"51",X"3A",X"FE",X"50",X"3D",
		X"32",X"FE",X"50",X"00",X"00",X"00",X"00",X"FE",X"FF",X"C2",X"7A",X"05",X"3E",X"09",X"32",X"FE",
		X"50",X"3A",X"1E",X"51",X"3D",X"32",X"1E",X"51",X"FE",X"FF",X"C2",X"7A",X"05",X"3E",X"09",X"32",
		X"1E",X"51",X"3A",X"3E",X"51",X"3D",X"32",X"3E",X"51",X"FE",X"FF",X"C2",X"7A",X"05",X"3E",X"09",
		X"32",X"3E",X"51",X"3A",X"5E",X"51",X"3D",X"32",X"5E",X"51",X"CD",X"EC",X"07",X"1E",X"1F",X"16",
		X"FF",X"CF",X"15",X"C2",X"81",X"05",X"1D",X"C2",X"81",X"05",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3A",X"FC",X"51",X"FE",X"00",X"C2",X"9E",X"05",X"3A",X"DC",X"51",X"FE",X"00",X"C8",X"3A",X"DC",
		X"51",X"3D",X"32",X"DC",X"51",X"FE",X"FF",X"C2",X"B6",X"05",X"3E",X"09",X"32",X"DC",X"51",X"3A",
		X"FC",X"51",X"3D",X"32",X"FC",X"51",X"3A",X"FE",X"50",X"3C",X"32",X"FE",X"50",X"FE",X"0A",X"C2",
		X"F0",X"05",X"3E",X"00",X"32",X"FE",X"50",X"3A",X"1E",X"51",X"3C",X"32",X"1E",X"51",X"FE",X"0A",
		X"C2",X"F0",X"05",X"3E",X"00",X"32",X"1E",X"51",X"3A",X"3E",X"51",X"3C",X"32",X"3E",X"51",X"FE",
		X"0A",X"C2",X"F0",X"05",X"3E",X"00",X"32",X"3E",X"51",X"3A",X"5E",X"51",X"3C",X"32",X"5E",X"51",
		X"1E",X"1F",X"16",X"FF",X"CF",X"15",X"C2",X"F4",X"05",X"1D",X"C2",X"F4",X"05",X"C9",X"FF",X"FF",
		X"3A",X"00",X"78",X"3A",X"00",X"60",X"E6",X"01",X"CA",X"7D",X"06",X"1E",X"0F",X"06",X"FF",X"3A",
		X"00",X"78",X"10",X"FB",X"1D",X"C2",X"0F",X"06",X"3A",X"00",X"60",X"E6",X"01",X"CA",X"7D",X"06",
		X"3A",X"FE",X"50",X"3C",X"32",X"FE",X"50",X"FE",X"0A",X"C2",X"5A",X"06",X"3E",X"00",X"32",X"FE",
		X"50",X"3A",X"1E",X"51",X"3C",X"32",X"1E",X"51",X"FE",X"0A",X"C2",X"5A",X"06",X"3E",X"00",X"32",
		X"1E",X"51",X"3A",X"3E",X"51",X"3C",X"32",X"3E",X"51",X"FE",X"0A",X"C2",X"5A",X"06",X"3E",X"00",
		X"32",X"3E",X"51",X"3A",X"5E",X"51",X"3C",X"32",X"5E",X"51",X"3E",X"01",X"32",X"03",X"60",X"3A",
		X"00",X"78",X"3A",X"00",X"60",X"E6",X"01",X"C2",X"5F",X"06",X"1E",X"0F",X"06",X"FF",X"3A",X"00",
		X"78",X"10",X"FB",X"1D",X"C2",X"6E",X"06",X"3E",X"00",X"32",X"03",X"60",X"C9",X"3A",X"00",X"60",
		X"E6",X"80",X"C8",X"1E",X"0F",X"06",X"FF",X"3A",X"00",X"78",X"10",X"FB",X"1D",X"C2",X"87",X"06",
		X"3A",X"00",X"60",X"E6",X"80",X"C8",X"00",X"00",X"3A",X"1E",X"51",X"3C",X"32",X"1E",X"51",X"FE",
		X"0A",X"C2",X"C1",X"06",X"3E",X"00",X"32",X"1E",X"51",X"3A",X"3E",X"51",X"3C",X"32",X"3E",X"51",
		X"FE",X"0A",X"C2",X"C1",X"06",X"3E",X"00",X"32",X"3E",X"51",X"3A",X"5E",X"51",X"3C",X"32",X"5E",
		X"51",X"3E",X"00",X"32",X"00",X"60",X"3A",X"00",X"78",X"3A",X"00",X"60",X"E6",X"80",X"C2",X"C6",
		X"06",X"1E",X"0F",X"06",X"FF",X"3A",X"00",X"78",X"10",X"FB",X"1D",X"C2",X"D5",X"06",X"3E",X"00",
		X"32",X"00",X"60",X"C9",X"C2",X"80",X"03",X"1E",X"0F",X"06",X"FF",X"3A",X"00",X"78",X"10",X"FB",
		X"1D",X"C2",X"EB",X"06",X"3A",X"00",X"60",X"06",X"08",X"A0",X"C2",X"80",X"03",X"C3",X"8A",X"03",
		X"CD",X"19",X"08",X"00",X"00",X"00",X"3A",X"09",X"40",X"32",X"31",X"40",X"3A",X"0A",X"40",X"32",
		X"32",X"40",X"3A",X"0B",X"40",X"32",X"33",X"40",X"78",X"32",X"3A",X"40",X"CD",X"60",X"21",X"CD",
		X"2A",X"23",X"20",X"F8",X"CD",X"78",X"23",X"CD",X"60",X"21",X"3A",X"30",X"40",X"21",X"10",X"40",
		X"46",X"B8",X"C2",X"27",X"07",X"CD",X"81",X"23",X"CD",X"60",X"22",X"3A",X"11",X"40",X"FE",X"16",
		X"DA",X"45",X"07",X"D6",X"16",X"47",X"3A",X"31",X"40",X"FE",X"16",X"DA",X"50",X"07",X"D6",X"16",
		X"B8",X"C2",X"38",X"07",X"CD",X"8A",X"23",X"CD",X"D0",X"22",X"3A",X"12",X"40",X"FE",X"16",X"DA",
		X"64",X"07",X"D6",X"16",X"47",X"3A",X"32",X"40",X"FE",X"16",X"DA",X"6F",X"07",X"D6",X"16",X"B8",
		X"C2",X"57",X"07",X"CD",X"F7",X"26",X"CD",X"30",X"23",X"3A",X"33",X"40",X"21",X"13",X"40",X"46",
		X"B8",X"C2",X"76",X"07",X"CD",X"80",X"23",X"3A",X"30",X"40",X"C6",X"30",X"6F",X"26",X"20",X"7E",
		X"32",X"40",X"40",X"3A",X"31",X"40",X"C6",X"30",X"6F",X"26",X"21",X"7E",X"32",X"41",X"40",X"3A",
		X"32",X"40",X"C6",X"30",X"6F",X"26",X"22",X"7E",X"32",X"42",X"40",X"3A",X"33",X"40",X"C6",X"30",
		X"6F",X"26",X"20",X"7E",X"32",X"43",X"40",X"00",X"00",X"00",X"C3",X"90",X"23",X"FF",X"FF",X"FF",
		X"3A",X"3A",X"40",X"3D",X"32",X"3A",X"40",X"C9",X"F1",X"C3",X"5B",X"03",X"FF",X"FF",X"FF",X"FF",
		X"C2",X"C9",X"03",X"1E",X"0F",X"06",X"FF",X"3A",X"00",X"78",X"10",X"FB",X"1D",X"C2",X"D7",X"07",
		X"3A",X"00",X"60",X"06",X"10",X"A0",X"C2",X"C9",X"03",X"C3",X"D3",X"03",X"3E",X"3F",X"32",X"00",
		X"78",X"16",X"FF",X"CF",X"1D",X"C2",X"F3",X"07",X"3E",X"FF",X"32",X"00",X"78",X"C9",X"FF",X"FF",
		X"21",X"00",X"70",X"46",X"3E",X"03",X"A0",X"32",X"22",X"40",X"32",X"24",X"40",X"3E",X"0C",X"A0",
		X"1F",X"1F",X"32",X"23",X"40",X"32",X"25",X"40",X"C9",X"3A",X"08",X"40",X"32",X"30",X"40",X"3A",
		X"10",X"40",X"C6",X"30",X"16",X"20",X"5F",X"1A",X"32",X"00",X"40",X"3A",X"11",X"40",X"C6",X"30",
		X"16",X"21",X"5F",X"1A",X"32",X"01",X"40",X"3A",X"12",X"40",X"C6",X"30",X"16",X"22",X"5F",X"1A",
		X"32",X"02",X"40",X"3A",X"13",X"40",X"C6",X"30",X"16",X"20",X"5F",X"1A",X"32",X"03",X"40",X"00",
		X"3A",X"00",X"40",X"21",X"01",X"40",X"46",X"B8",X"20",X"35",X"3A",X"02",X"40",X"B8",X"20",X"69",
		X"21",X"03",X"40",X"46",X"B8",X"20",X"37",X"3A",X"22",X"40",X"E6",X"03",X"C8",X"3A",X"24",X"40",
		X"E6",X"03",X"20",X"07",X"3A",X"22",X"40",X"32",X"24",X"40",X"C9",X"3D",X"32",X"24",X"40",X"3A",
		X"11",X"40",X"3C",X"FE",X"16",X"20",X"04",X"3A",X"11",X"40",X"3D",X"32",X"11",X"40",X"C9",X"21",
		X"02",X"40",X"46",X"3A",X"00",X"40",X"B8",X"20",X"28",X"3A",X"03",X"40",X"B8",X"C0",X"3A",X"23",
		X"40",X"E6",X"03",X"C8",X"3A",X"25",X"40",X"E6",X"03",X"28",X"3E",X"3D",X"32",X"25",X"40",X"00",
		X"00",X"3A",X"12",X"40",X"3C",X"FE",X"16",X"20",X"04",X"3A",X"12",X"40",X"3D",X"32",X"12",X"40",
		X"C9",X"3A",X"01",X"40",X"B8",X"C0",X"C3",X"99",X"08",X"21",X"01",X"40",X"46",X"3A",X"03",X"40",
		X"B8",X"C0",X"3A",X"23",X"40",X"E6",X"03",X"C8",X"3A",X"25",X"40",X"00",X"E6",X"03",X"28",X"09",
		X"3D",X"32",X"25",X"40",X"00",X"00",X"C3",X"7F",X"08",X"3A",X"23",X"40",X"32",X"25",X"40",X"C9",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3A",X"00",X"68",X"E6",X"80",X"20",X"0D",X"3A",X"00",X"68",X"E6",X"40",X"20",X"0C",X"3A",X"FC",
		X"51",X"FE",X"02",X"C9",X"3A",X"FC",X"51",X"FE",X"01",X"C9",X"3A",X"DC",X"51",X"FE",X"06",X"C9",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"A0",X"40",X"A0",X"50",X"90",X"80",X"A0",X"70",X"A0",X"30",X"90",X"60",X"A0",X"80",X"A0",X"50",
		X"A0",X"70",X"B0",X"20",X"90",X"60",X"FF",X"9E",X"7B",X"62",X"4A",X"BF",X"15",X"04",X"26",X"51",
		X"7A",X"9E",X"11",X"00",X"C2",X"A5",X"05",X"BF",X"CF",X"76",X"5A",X"3A",X"26",X"55",X"BA",X"EF",
		X"10",X"04",X"08",X"20",X"08",X"06",X"10",X"18",X"08",X"02",X"08",X"40",X"10",X"04",X"08",X"18",
		X"08",X"06",X"08",X"02",X"01",X"60",X"FF",X"BB",X"CF",X"6A",X"59",X"52",X"41",X"05",X"27",X"B6",
		X"21",X"E8",X"52",X"EF",X"3A",X"30",X"40",X"6F",X"26",X"20",X"46",X"3A",X"38",X"40",X"80",X"21",
		X"E8",X"52",X"11",X"20",X"00",X"77",X"19",X"C6",X"04",X"77",X"19",X"C6",X"04",X"77",X"19",X"C6",
		X"04",X"77",X"21",X"28",X"52",X"EF",X"3A",X"31",X"40",X"6F",X"26",X"21",X"46",X"3A",X"38",X"40",
		X"80",X"21",X"28",X"52",X"11",X"20",X"00",X"77",X"19",X"C6",X"04",X"77",X"19",X"C6",X"04",X"77",
		X"19",X"C6",X"04",X"77",X"21",X"68",X"51",X"EF",X"3A",X"32",X"40",X"6F",X"26",X"22",X"46",X"3A",
		X"38",X"40",X"80",X"21",X"68",X"51",X"11",X"20",X"00",X"77",X"19",X"C6",X"04",X"77",X"19",X"C6",
		X"04",X"77",X"19",X"C6",X"04",X"77",X"21",X"A8",X"50",X"EF",X"3A",X"33",X"40",X"6F",X"26",X"20",
		X"46",X"3A",X"38",X"40",X"80",X"21",X"A8",X"50",X"11",X"20",X"00",X"77",X"19",X"C6",X"04",X"77",
		X"19",X"C6",X"04",X"77",X"19",X"C6",X"04",X"77",X"C9",X"CA",X"30",X"03",X"3A",X"00",X"78",X"3A",
		X"00",X"60",X"E6",X"01",X"CA",X"F8",X"27",X"CF",X"3A",X"00",X"60",X"E6",X"18",X"CA",X"30",X"03",
		X"E6",X"08",X"CA",X"E7",X"20",X"CD",X"E0",X"26",X"00",X"00",X"00",X"00",X"C3",X"C8",X"23",X"FF",
		X"A0",X"50",X"B0",X"80",X"90",X"40",X"B0",X"80",X"A0",X"80",X"B0",X"70",X"B0",X"20",X"80",X"60",
		X"B0",X"80",X"90",X"30",X"B0",X"80",X"90",X"50",X"B0",X"80",X"90",X"40",X"B0",X"80",X"A0",X"80",
		X"B0",X"70",X"B0",X"20",X"80",X"60",X"B0",X"80",X"90",X"30",X"B0",X"80",X"FF",X"FF",X"FF",X"FF",
		X"01",X"18",X"08",X"06",X"01",X"18",X"10",X"20",X"01",X"18",X"08",X"18",X"01",X"02",X"01",X"60",
		X"18",X"04",X"01",X"18",X"10",X"40",X"FF",X"9A",X"26",X"56",X"94",X"11",X"37",X"21",X"05",X"04",
		X"98",X"DC",X"BE",X"A6",X"96",X"25",X"7B",X"FE",X"6A",X"5B",X"46",X"2B",X"D9",X"36",X"75",X"42",
		X"3E",X"01",X"32",X"38",X"40",X"CD",X"50",X"20",X"CD",X"D0",X"21",X"AF",X"32",X"38",X"40",X"CD",
		X"50",X"20",X"CD",X"D0",X"21",X"3A",X"30",X"40",X"3C",X"FE",X"16",X"C2",X"80",X"21",X"3E",X"00",
		X"32",X"30",X"40",X"3A",X"31",X"40",X"3C",X"FE",X"16",X"C2",X"8E",X"21",X"3E",X"00",X"32",X"31",
		X"40",X"00",X"00",X"00",X"00",X"3A",X"32",X"40",X"3C",X"FE",X"16",X"C2",X"A0",X"21",X"3E",X"00",
		X"32",X"32",X"40",X"00",X"00",X"00",X"00",X"3A",X"33",X"40",X"3C",X"FE",X"16",X"C2",X"B2",X"21",
		X"3E",X"00",X"32",X"33",X"40",X"3E",X"03",X"32",X"38",X"40",X"CD",X"50",X"20",X"CD",X"D0",X"21",
		X"3E",X"02",X"32",X"38",X"40",X"CD",X"50",X"20",X"CD",X"D0",X"21",X"C9",X"FF",X"FF",X"FF",X"FF",
		X"3E",X"01",X"32",X"00",X"78",X"1E",X"FF",X"CF",X"1D",X"C2",X"D7",X"21",X"3E",X"FF",X"32",X"00",
		X"78",X"C9",X"CF",X"32",X"65",X"04",X"3A",X"7B",X"5A",X"E8",X"61",X"45",X"BF",X"20",X"10",X"41",
		X"8C",X"E7",X"21",X"7B",X"55",X"41",X"6B",X"E9",X"8A",X"55",X"21",X"7B",X"FE",X"44",X"00",X"6A",
		X"B0",X"90",X"80",X"30",X"B0",X"90",X"A0",X"50",X"B0",X"90",X"80",X"40",X"B0",X"90",X"A0",X"90",
		X"B0",X"70",X"B0",X"20",X"90",X"60",X"B0",X"90",X"80",X"30",X"B0",X"90",X"A0",X"50",X"B0",X"90",
		X"80",X"40",X"B0",X"90",X"A0",X"90",X"B0",X"70",X"B0",X"20",X"90",X"60",X"FF",X"FF",X"FF",X"FF",
		X"10",X"04",X"01",X"10",X"18",X"40",X"01",X"10",X"08",X"06",X"01",X"10",X"18",X"20",X"01",X"10",
		X"08",X"10",X"01",X"02",X"01",X"60",X"FF",X"CF",X"3A",X"54",X"00",X"7B",X"65",X"41",X"7B",X"AA",
		X"9F",X"BA",X"CA",X"25",X"06",X"49",X"81",X"BA",X"3B",X"5A",X"11",X"2B",X"20",X"DE",X"4A",X"89",
		X"3E",X"01",X"32",X"38",X"40",X"CD",X"72",X"20",X"CD",X"D0",X"21",X"AF",X"32",X"38",X"40",X"CD",
		X"72",X"20",X"CD",X"D0",X"21",X"3A",X"31",X"40",X"3C",X"FE",X"16",X"C2",X"80",X"22",X"3E",X"00",
		X"32",X"31",X"40",X"00",X"00",X"00",X"00",X"3A",X"32",X"40",X"3C",X"FE",X"16",X"C2",X"92",X"22",
		X"3E",X"00",X"32",X"32",X"40",X"00",X"00",X"00",X"00",X"3A",X"33",X"40",X"3C",X"FE",X"16",X"C2",
		X"A4",X"22",X"3E",X"00",X"32",X"33",X"40",X"3E",X"03",X"32",X"38",X"40",X"CD",X"72",X"20",X"CD",
		X"D0",X"21",X"3E",X"02",X"32",X"38",X"40",X"CD",X"72",X"20",X"CD",X"D0",X"21",X"C9",X"FF",X"FF",
		X"1E",X"FF",X"CF",X"1D",X"C2",X"C2",X"22",X"C9",X"3A",X"00",X"60",X"2F",X"E6",X"20",X"18",X"58",
		X"3E",X"01",X"32",X"38",X"40",X"CD",X"94",X"20",X"CD",X"D0",X"21",X"AF",X"32",X"38",X"40",X"CD",
		X"94",X"20",X"CD",X"D0",X"21",X"3A",X"32",X"40",X"3C",X"FE",X"16",X"C2",X"F0",X"22",X"3E",X"00",
		X"32",X"32",X"40",X"00",X"00",X"00",X"00",X"3A",X"33",X"40",X"3C",X"FE",X"16",X"C2",X"02",X"23",
		X"3E",X"00",X"32",X"33",X"40",X"3E",X"03",X"32",X"38",X"40",X"CD",X"94",X"20",X"CD",X"D0",X"21",
		X"3E",X"02",X"32",X"38",X"40",X"CD",X"94",X"20",X"CD",X"D0",X"21",X"C9",X"FF",X"FF",X"FF",X"FF",
		X"1E",X"FF",X"CF",X"1D",X"C2",X"22",X"23",X"C9",X"28",X"40",X"CD",X"C0",X"07",X"C0",X"18",X"3A",
		X"3E",X"01",X"32",X"38",X"40",X"CD",X"B6",X"20",X"CD",X"D0",X"21",X"AF",X"32",X"38",X"40",X"CD",
		X"B6",X"20",X"CD",X"D0",X"21",X"3A",X"33",X"40",X"3C",X"FE",X"16",X"C2",X"50",X"23",X"3E",X"00",
		X"32",X"33",X"40",X"3E",X"03",X"32",X"38",X"40",X"CD",X"B6",X"20",X"CD",X"D0",X"21",X"3E",X"02",
		X"32",X"38",X"40",X"CD",X"B6",X"20",X"CD",X"D0",X"21",X"C9",X"3E",X"10",X"32",X"3A",X"40",X"C9",
		X"1E",X"FF",X"CF",X"1D",X"C2",X"72",X"23",X"C9",X"CD",X"60",X"21",X"CD",X"C8",X"22",X"20",X"F8",
		X"C9",X"CD",X"60",X"22",X"CD",X"C8",X"22",X"20",X"F8",X"C9",X"CD",X"D0",X"22",X"C3",X"98",X"27",
		X"3A",X"30",X"40",X"32",X"08",X"40",X"3A",X"31",X"40",X"32",X"09",X"40",X"3A",X"32",X"40",X"32",
		X"0A",X"40",X"3A",X"33",X"40",X"32",X"0B",X"40",X"C3",X"00",X"24",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3E",X"1F",X"32",X"00",X"78",X"16",X"0F",X"1E",X"FF",X"CF",X"1D",X"C2",X"B9",X"23",X"15",X"C2",
		X"B9",X"23",X"3E",X"FF",X"32",X"00",X"78",X"C9",X"3A",X"00",X"60",X"E6",X"08",X"CA",X"30",X"03",
		X"3A",X"00",X"78",X"3A",X"00",X"60",X"E6",X"01",X"CA",X"C8",X"23",X"CF",X"CD",X"00",X"05",X"CF",
		X"3A",X"00",X"60",X"E6",X"08",X"C2",X"DC",X"23",X"3E",X"0F",X"32",X"11",X"40",X"3E",X"15",X"32",
		X"12",X"40",X"32",X"13",X"40",X"CF",X"3A",X"00",X"60",X"E6",X"10",X"C3",X"F0",X"26",X"FF",X"FF",
		X"3A",X"00",X"78",X"3A",X"FC",X"51",X"FE",X"1C",X"20",X"01",X"AF",X"4F",X"1E",X"0A",X"CD",X"00",
		X"27",X"3A",X"DC",X"51",X"83",X"32",X"88",X"40",X"CD",X"00",X"25",X"32",X"8A",X"40",X"A7",X"CA",
		X"D0",X"24",X"4F",X"3A",X"00",X"78",X"06",X"00",X"11",X"64",X"0A",X"79",X"93",X"28",X"02",X"38",
		X"04",X"4F",X"04",X"18",X"F6",X"78",X"A7",X"28",X"00",X"32",X"BC",X"52",X"06",X"00",X"3A",X"00",
		X"78",X"79",X"92",X"28",X"02",X"38",X"04",X"4F",X"04",X"18",X"F3",X"78",X"A7",X"20",X"07",X"3A",
		X"BC",X"52",X"FE",X"1C",X"28",X"04",X"78",X"32",X"9C",X"52",X"79",X"32",X"7C",X"52",X"3A",X"00",
		X"78",X"3A",X"88",X"40",X"4F",X"3A",X"8A",X"40",X"5F",X"CD",X"00",X"27",X"ED",X"53",X"8C",X"40",
		X"C3",X"B0",X"27",X"3A",X"00",X"78",X"21",X"5E",X"51",X"11",X"20",X"22",X"06",X"04",X"7E",X"FE",
		X"09",X"20",X"0C",X"05",X"CA",X"8F",X"24",X"3A",X"00",X"78",X"AF",X"ED",X"52",X"18",X"EF",X"2A",
		X"8C",X"40",X"11",X"01",X"00",X"3A",X"00",X"78",X"AF",X"ED",X"52",X"22",X"8C",X"40",X"CD",X"18",
		X"27",X"21",X"FE",X"50",X"11",X"20",X"00",X"3A",X"00",X"78",X"7E",X"FE",X"09",X"20",X"05",X"36",
		X"00",X"19",X"18",X"F3",X"FE",X"1C",X"20",X"01",X"AF",X"3C",X"77",X"3A",X"00",X"78",X"CD",X"B0",
		X"23",X"CD",X"F8",X"24",X"2A",X"8C",X"40",X"AF",X"BD",X"C2",X"73",X"24",X"BC",X"C2",X"73",X"24",
		X"0E",X"FF",X"CD",X"F8",X"24",X"0D",X"20",X"FA",X"21",X"DC",X"51",X"11",X"20",X"00",X"AF",X"77",
		X"19",X"77",X"21",X"7C",X"52",X"06",X"03",X"77",X"19",X"10",X"FC",X"3A",X"00",X"78",X"C3",X"C8",
		X"27",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"06",X"FF",X"3A",X"00",X"78",X"10",X"FB",X"C9",
		X"21",X"40",X"40",X"06",X"04",X"3A",X"00",X"78",X"7E",X"A7",X"C8",X"E6",X"80",X"20",X"05",X"23",
		X"10",X"F6",X"18",X"02",X"AF",X"C9",X"2B",X"56",X"2B",X"4E",X"2B",X"46",X"2B",X"5E",X"3A",X"00",
		X"78",X"78",X"B9",X"C2",X"BA",X"25",X"7B",X"BA",X"C2",X"78",X"25",X"B8",X"CA",X"51",X"25",X"E6",
		X"9F",X"20",X"08",X"78",X"E6",X"9F",X"20",X"03",X"3E",X"14",X"C9",X"3A",X"00",X"78",X"7B",X"FE",
		X"01",X"28",X"0B",X"E6",X"F9",X"28",X"07",X"78",X"E6",X"F9",X"28",X"02",X"AF",X"C9",X"3E",X"02",
		X"C9",X"3A",X"00",X"78",X"7B",X"21",X"63",X"25",X"01",X"0B",X"00",X"ED",X"B1",X"21",X"6D",X"25",
		X"09",X"7E",X"C9",X"01",X"02",X"04",X"06",X"08",X"10",X"18",X"20",X"40",X"60",X"00",X"FA",X"FA",
		X"FA",X"32",X"14",X"14",X"C8",X"C8",X"C8",X"14",X"3A",X"00",X"78",X"7B",X"B8",X"28",X"05",X"78",
		X"BA",X"C2",X"9E",X"25",X"78",X"21",X"63",X"25",X"01",X"0B",X"00",X"ED",X"B1",X"21",X"93",X"25",
		X"09",X"7E",X"C9",X"00",X"C8",X"64",X"32",X"14",X"0E",X"0A",X"14",X"14",X"14",X"0A",X"E6",X"9F",
		X"20",X"0D",X"7B",X"E6",X"9F",X"28",X"05",X"7A",X"E6",X"9F",X"20",X"03",X"3E",X"14",X"C9",X"3E",
		X"01",X"BB",X"28",X"04",X"BA",X"C2",X"47",X"25",X"3C",X"C9",X"3A",X"00",X"78",X"78",X"E6",X"9F",
		X"20",X"03",X"79",X"E6",X"9F",X"C2",X"EC",X"25",X"7B",X"E6",X"9F",X"20",X"03",X"3E",X"14",X"C9",
		X"7A",X"E6",X"9F",X"28",X"F8",X"3E",X"01",X"BB",X"28",X"03",X"BA",X"20",X"02",X"3C",X"C9",X"7B",
		X"BA",X"20",X"07",X"E6",X"F9",X"20",X"03",X"3E",X"02",X"C9",X"AF",X"C9",X"3A",X"00",X"78",X"7B",
		X"B8",X"20",X"0B",X"FE",X"01",X"20",X"03",X"3E",X"05",X"C9",X"E6",X"F9",X"28",X"0E",X"7A",X"B9",
		X"C2",X"14",X"26",X"FE",X"01",X"28",X"F0",X"E6",X"F9",X"C2",X"14",X"26",X"7B",X"BA",X"C2",X"20",
		X"26",X"3E",X"14",X"C9",X"3A",X"00",X"78",X"7B",X"BA",X"C2",X"2A",X"26",X"E6",X"F9",X"20",X"03",
		X"3E",X"02",X"C9",X"7B",X"FE",X"01",X"28",X"F8",X"AF",X"C9",X"3A",X"00",X"78",X"7B",X"B9",X"20",
		X"07",X"E6",X"F9",X"20",X"03",X"3E",X"02",X"C9",X"7B",X"FE",X"01",X"28",X"F8",X"7A",X"B8",X"20",
		X"04",X"E6",X"F9",X"28",X"F0",X"7A",X"FE",X"01",X"28",X"EB",X"AF",X"C9",X"16",X"0B",X"06",X"0A",
		X"8A",X"37",X"FE",X"76",X"5A",X"9E",X"DA",X"45",X"22",X"00",X"7B",X"FF",X"6B",X"9E",X"6A",X"58",
		X"DC",X"C2",X"0F",X"1A",X"3A",X"5B",X"71",X"6A",X"8E",X"B7",X"22",X"33",X"7B",X"00",X"11",X"22",
		X"33",X"44",X"55",X"66",X"77",X"88",X"99",X"AA",X"BB",X"CC",X"DD",X"EE",X"FF",X"01",X"23",X"45",
		X"67",X"89",X"AB",X"CD",X"EF",X"01",X"12",X"23",X"34",X"45",X"56",X"67",X"78",X"89",X"9A",X"AB",
		X"BC",X"CD",X"DE",X"EF",X"F0",X"00",X"01",X"02",X"03",X"04",X"05",X"06",X"07",X"08",X"09",X"0A",
		X"0B",X"0C",X"0D",X"0E",X"0F",X"F0",X"F1",X"F2",X"F3",X"F4",X"F5",X"F6",X"F7",X"F8",X"F9",X"FA",
		X"FB",X"FC",X"FD",X"FE",X"FF",X"05",X"AF",X"16",X"B2",X"73",X"49",X"E8",X"DC",X"21",X"65",X"A9",
		X"20",X"37",X"B8",X"3A",X"26",X"54",X"32",X"05",X"48",X"CF",X"76",X"9A",X"B5",X"48",X"05",X"CD",
		X"BF",X"62",X"40",X"B9",X"FA",X"96",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"1E",X"1F",X"16",X"FF",X"CF",X"1D",X"C2",X"E4",X"26",X"15",X"C2",X"E4",X"26",X"C9",X"FF",X"FF",
		X"CA",X"F5",X"23",X"C3",X"00",X"07",X"FF",X"CD",X"30",X"23",X"CD",X"C8",X"22",X"20",X"F8",X"C9",
		X"3A",X"00",X"78",X"AF",X"57",X"06",X"08",X"CB",X"1B",X"30",X"03",X"7A",X"81",X"57",X"CB",X"3A",
		X"10",X"F5",X"CB",X"1B",X"3A",X"00",X"78",X"C9",X"21",X"FC",X"50",X"11",X"20",X"00",X"06",X"04",
		X"00",X"00",X"19",X"10",X"FB",X"2A",X"8C",X"40",X"11",X"E8",X"03",X"06",X"00",X"22",X"8E",X"40",
		X"3A",X"00",X"78",X"AF",X"ED",X"52",X"28",X"02",X"38",X"03",X"04",X"18",X"F0",X"78",X"A7",X"28",
		X"00",X"D6",X"0A",X"F2",X"A0",X"27",X"78",X"32",X"5C",X"51",X"2A",X"8E",X"40",X"11",X"64",X"00",
		X"06",X"00",X"22",X"8E",X"40",X"3A",X"00",X"78",X"AF",X"ED",X"52",X"28",X"02",X"38",X"03",X"04",
		X"18",X"F0",X"78",X"A7",X"20",X"07",X"3A",X"5C",X"51",X"FE",X"1C",X"28",X"04",X"78",X"32",X"3C",
		X"51",X"3A",X"00",X"78",X"3A",X"8E",X"40",X"1E",X"0A",X"06",X"00",X"4F",X"93",X"28",X"02",X"38",
		X"03",X"04",X"18",X"F7",X"78",X"A7",X"20",X"07",X"3A",X"3C",X"51",X"FE",X"1C",X"28",X"04",X"78",
		X"32",X"1C",X"51",X"79",X"32",X"FC",X"50",X"C9",X"CD",X"C8",X"22",X"C2",X"8A",X"23",X"C9",X"FF",
		X"21",X"0F",X"27",X"22",X"8C",X"40",X"C3",X"18",X"27",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"CD",X"18",X"27",X"11",X"FF",X"FF",X"CF",X"1D",X"C2",X"B6",X"27",X"15",X"C2",X"B6",X"27",X"3A",
		X"FC",X"50",X"32",X"3A",X"40",X"C3",X"73",X"24",X"3A",X"3A",X"40",X"FE",X"00",X"CA",X"30",X"03",
		X"3A",X"00",X"60",X"E6",X"04",X"CA",X"30",X"03",X"3A",X"00",X"78",X"3A",X"00",X"60",X"E6",X"01",
		X"CA",X"D0",X"27",X"CF",X"3A",X"00",X"60",X"E6",X"14",X"CA",X"30",X"03",X"E6",X"10",X"CA",X"E3",
		X"27",X"CD",X"E0",X"26",X"00",X"00",X"00",X"00",X"3A",X"00",X"60",X"E6",X"10",X"C3",X"D9",X"20");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
