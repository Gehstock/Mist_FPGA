library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity kick_sp_bits_4 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of kick_sp_bits_4 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"EE",X"EE",X"E0",X"EE",X"EE",X"00",X"E0",X"00",X"0E",X"00",X"E0",X"00",X"0E",X"00",X"E0",
		X"00",X"0E",X"00",X"E0",X"00",X"0E",X"00",X"E0",X"00",X"0E",X"00",X"E0",X"00",X"0E",X"E0",X"00",
		X"0E",X"0E",X"0E",X"00",X"E0",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"E0",X"0E",X"00",X"00",
		X"EE",X"0E",X"0E",X"00",X"EE",X"0E",X"EE",X"00",X"0E",X"0E",X"E0",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"0E",X"0E",X"E0",X"00",X"EE",X"0E",X"EE",X"00",X"EE",X"0E",X"0E",X"00",
		X"E0",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"E0",X"0E",X"00",X"00",X"0E",X"0E",X"0E",X"00",
		X"00",X"0E",X"E0",X"00",X"00",X"0E",X"00",X"E0",X"00",X"0E",X"00",X"E0",X"00",X"0E",X"00",X"E0",
		X"00",X"0E",X"00",X"E0",X"00",X"0E",X"00",X"E0",X"EE",X"EE",X"00",X"E0",X"EE",X"EE",X"00",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"0E",X"0E",X"E0",X"00",X"EE",X"0E",X"EE",X"00",X"EE",X"0E",X"0E",X"00",
		X"E0",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"E0",X"0E",X"00",X"00",X"DD",X"0E",X"0E",X"00",
		X"DD",X"0E",X"E0",X"00",X"DD",X"0E",X"00",X"E0",X"DD",X"0E",X"00",X"E0",X"DD",X"0E",X"00",X"E0",
		X"D0",X"0E",X"00",X"E0",X"D0",X"0E",X"00",X"E0",X"D2",X"EE",X"00",X"E0",X"D2",X"EE",X"EE",X"E0",
		X"44",X"4F",X"77",X"77",X"44",X"4F",X"77",X"77",X"44",X"4F",X"77",X"77",X"44",X"4F",X"77",X"77",
		X"44",X"4F",X"77",X"77",X"44",X"4F",X"77",X"77",X"44",X"4F",X"77",X"77",X"44",X"40",X"77",X"00",
		X"40",X"40",X"77",X"00",X"00",X"40",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"3F",X"77",X"22",X"43",X"3F",X"77",X"22",X"43",X"3F",X"77",X"22",X"44",X"3F",X"77",X"22",
		X"44",X"3F",X"77",X"22",X"44",X"3F",X"77",X"00",X"44",X"3F",X"77",X"00",X"44",X"00",X"70",X"00",
		X"44",X"00",X"BB",X"00",X"44",X"00",X"B0",X"00",X"44",X"45",X"00",X"00",X"44",X"4F",X"00",X"00",
		X"44",X"55",X"BB",X"00",X"44",X"55",X"BB",X"00",X"44",X"4F",X"00",X"00",X"44",X"05",X"00",X"00",
		X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"3B",X"77",X"77",X"33",X"3B",X"77",X"77",X"43",X"3B",X"77",X"77",X"43",X"BB",X"77",X"77",
		X"44",X"BB",X"77",X"22",X"44",X"FB",X"77",X"00",X"44",X"5B",X"77",X"00",X"44",X"F0",X"77",X"00",
		X"44",X"50",X"70",X"00",X"44",X"00",X"70",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",
		X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"B0",X"00",X"00",X"4B",X"B0",
		X"00",X"00",X"4B",X"BB",X"00",X"00",X"4B",X"BB",X"00",X"00",X"4B",X"BB",X"00",X"00",X"4B",X"BB",
		X"00",X"00",X"4B",X"BB",X"00",X"00",X"4B",X"00",X"00",X"00",X"4B",X"00",X"00",X"00",X"40",X"00",
		X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"BB",X"00",X"00",X"40",X"BB",X"00",X"00",X"40",X"7B",
		X"00",X"00",X"4B",X"BB",X"00",X"00",X"4B",X"BB",X"00",X"00",X"4B",X"BB",X"00",X"00",X"4B",X"AB",
		X"00",X"00",X"4B",X"A0",X"00",X"00",X"4B",X"A0",X"00",X"00",X"4B",X"A0",X"00",X"00",X"4B",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",
		X"00",X"00",X"4B",X"00",X"00",X"00",X"4B",X"A0",X"00",X"00",X"4B",X"AB",X"00",X"00",X"4B",X"BB",
		X"00",X"00",X"4A",X"BB",X"00",X"00",X"4A",X"BB",X"00",X"00",X"4A",X"00",X"00",X"00",X"4A",X"00",
		X"00",X"00",X"4A",X"00",X"00",X"00",X"4A",X"00",X"00",X"00",X"4A",X"00",X"00",X"00",X"AA",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",
		X"00",X"00",X"11",X"10",X"00",X"00",X"11",X"10",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",
		X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",
		X"00",X"00",X"77",X"11",X"00",X"3F",X"77",X"11",X"00",X"3F",X"77",X"77",X"00",X"3F",X"77",X"77",
		X"50",X"3F",X"77",X"77",X"55",X"3F",X"77",X"77",X"33",X"3F",X"77",X"77",X"33",X"3F",X"77",X"77",
		X"00",X"00",X"DD",X"00",X"00",X"0D",X"DD",X"00",X"00",X"DD",X"DD",X"07",X"00",X"DD",X"DD",X"00",
		X"00",X"DD",X"DD",X"00",X"00",X"DD",X"77",X"00",X"00",X"0D",X"77",X"00",X"00",X"00",X"77",X"00",
		X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",
		X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",
		X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",
		X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"B0",X"B0",X"77",X"00",X"BB",X"00",X"77",X"70",
		X"2B",X"00",X"77",X"77",X"0B",X"00",X"77",X"77",X"BB",X"00",X"77",X"77",X"BB",X"00",X"77",X"77",
		X"BB",X"00",X"77",X"77",X"25",X"00",X"77",X"77",X"25",X"00",X"77",X"77",X"25",X"00",X"77",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"EE",X"EE",X"E0",X"EE",X"EE",X"00",X"E0",X"00",X"0E",X"00",X"E0",X"00",X"0E",X"00",X"E0",
		X"00",X"0E",X"00",X"E0",X"00",X"0E",X"00",X"E0",X"00",X"0E",X"00",X"E0",X"00",X"0E",X"E0",X"00",
		X"0E",X"0E",X"0E",X"00",X"E0",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"E0",X"0E",X"00",X"00",
		X"EE",X"0E",X"0E",X"00",X"EE",X"0E",X"EE",X"00",X"0E",X"0E",X"E0",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DE",X"EE",X"22",X"E0",X"DD",X"EE",X"22",X"E0",X"DD",X"0E",X"00",X"E0",X"77",X"5E",X"00",X"E0",
		X"00",X"0E",X"00",X"E0",X"00",X"0E",X"00",X"E0",X"00",X"0E",X"E0",X"E0",X"00",X"0E",X"0E",X"00",
		X"0E",X"0E",X"00",X"00",X"E0",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"E0",X"0E",X"00",X"00",
		X"EE",X"0E",X"0E",X"00",X"EE",X"0E",X"EE",X"00",X"00",X"0E",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"EE",X"EE",X"E0",X"7E",X"88",X"00",X"E0",X"00",X"88",X"00",X"E0",X"00",X"80",X"00",X"E0",
		X"00",X"22",X"00",X"E0",X"00",X"22",X"00",X"E0",X"0E",X"22",X"00",X"E0",X"E0",X"22",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"0E",X"00",
		X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",
		X"EE",X"00",X"0E",X"00",X"EE",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",
		X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"70",X"BB",X"00",X"77",X"70",
		X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",
		X"50",X"00",X"77",X"77",X"55",X"3F",X"77",X"77",X"33",X"3F",X"77",X"77",X"33",X"3F",X"77",X"77",
		X"33",X"4F",X"77",X"77",X"33",X"4F",X"77",X"77",X"33",X"44",X"77",X"27",X"34",X"44",X"77",X"27",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"B0",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"05",X"00",X"11",X"00",X"04",X"00",X"11",
		X"00",X"44",X"00",X"11",X"00",X"44",X"00",X"11",X"00",X"44",X"77",X"11",X"00",X"44",X"77",X"11",
		X"50",X"44",X"77",X"11",X"55",X"B3",X"77",X"11",X"33",X"B3",X"77",X"00",X"33",X"B3",X"77",X"00",
		X"33",X"F5",X"77",X"77",X"33",X"F5",X"77",X"77",X"33",X"F5",X"77",X"77",X"33",X"44",X"77",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0B",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"01",X"00",
		X"BB",X"00",X"11",X"00",X"BB",X"00",X"11",X"00",X"BB",X"00",X"11",X"00",X"BB",X"00",X"11",X"00",
		X"BB",X"00",X"11",X"00",X"BB",X"00",X"11",X"10",X"05",X"00",X"11",X"11",X"00",X"00",X"11",X"11",
		X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"40",X"71",X"11",X"00",X"44",X"77",X"11",
		X"50",X"44",X"77",X"11",X"55",X"3F",X"77",X"77",X"33",X"3F",X"77",X"77",X"33",X"3F",X"77",X"77",
		X"33",X"3F",X"77",X"77",X"33",X"3F",X"77",X"77",X"33",X"3F",X"77",X"77",X"33",X"3F",X"77",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"B0",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"40",X"00",X"77",
		X"00",X"40",X"00",X"77",X"00",X"40",X"00",X"77",X"00",X"40",X"00",X"77",X"00",X"40",X"00",X"77",
		X"00",X"40",X"00",X"77",X"00",X"40",X"00",X"77",X"00",X"40",X"00",X"77",X"00",X"30",X"77",X"77",
		X"50",X"3F",X"77",X"77",X"55",X"3F",X"77",X"77",X"33",X"3F",X"77",X"77",X"33",X"3F",X"77",X"77",
		X"33",X"3F",X"77",X"77",X"33",X"3F",X"77",X"22",X"33",X"3F",X"77",X"22",X"33",X"3F",X"77",X"27",
		X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"0D",X"DD",X"DD",X"00",X"0D",X"DD",X"DD",
		X"00",X"DD",X"DD",X"D0",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",
		X"00",X"DD",X"D0",X"00",X"00",X"0D",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"07",
		X"00",X"00",X"BB",X"77",X"00",X"00",X"B0",X"77",X"00",X"00",X"B0",X"77",X"00",X"05",X"00",X"77",
		X"00",X"0F",X"00",X"77",X"00",X"44",X"00",X"77",X"00",X"44",X"00",X"77",X"00",X"44",X"00",X"77",
		X"00",X"44",X"00",X"77",X"04",X"44",X"00",X"77",X"44",X"40",X"00",X"70",X"44",X"00",X"07",X"70",
		X"44",X"00",X"77",X"70",X"44",X"00",X"77",X"00",X"44",X"00",X"77",X"00",X"44",X"00",X"77",X"00",
		X"44",X"33",X"77",X"00",X"33",X"33",X"77",X"00",X"53",X"33",X"77",X"0E",X"55",X"33",X"77",X"EE",
		X"55",X"33",X"77",X"EE",X"53",X"33",X"77",X"EE",X"33",X"33",X"77",X"00",X"44",X"33",X"77",X"10",
		X"44",X"33",X"77",X"10",X"44",X"00",X"71",X"11",X"44",X"00",X"11",X"11",X"44",X"00",X"11",X"11",
		X"44",X"00",X"01",X"11",X"44",X"40",X"00",X"11",X"04",X"44",X"00",X"11",X"00",X"44",X"00",X"11",
		X"00",X"44",X"00",X"11",X"00",X"44",X"00",X"11",X"00",X"44",X"00",X"11",X"05",X"40",X"00",X"11",
		X"BB",X"40",X"00",X"11",X"BB",X"00",X"00",X"11",X"BB",X"00",X"11",X"11",X"BB",X"00",X"11",X"10",
		X"B0",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"10",X"DD",
		X"00",X"00",X"00",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"0D",X"DD",X"DD",X"00",X"0D",X"DD",X"DD",
		X"00",X"0D",X"DD",X"DD",X"00",X"0D",X"DD",X"DD",X"00",X"0D",X"DD",X"DD",X"00",X"0D",X"00",X"DD",
		X"77",X"55",X"20",X"E0",X"77",X"FF",X"20",X"E0",X"77",X"55",X"E0",X"E0",X"77",X"00",X"0E",X"E0",
		X"EE",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",
		X"0E",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"E0",X"00",
		X"EE",X"00",X"EE",X"00",X"EE",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"5F",X"DD",X"00",X"E0",X"35",X"DD",X"00",X"E0",X"30",X"DE",X"00",X"E0",X"00",X"2E",X"00",X"E0",
		X"00",X"2E",X"00",X"E0",X"00",X"2E",X"EE",X"E0",X"00",X"20",X"00",X"E0",X"00",X"00",X"00",X"00",
		X"0E",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",
		X"EE",X"00",X"EE",X"00",X"EE",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"EE",X"00",X"EE",X"00",X"EE",X"00",
		X"E0",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"88",X"00",X"00",
		X"00",X"88",X"00",X"00",X"00",X"88",X"00",X"00",X"E0",X"88",X"00",X"00",X"7E",X"08",X"00",X"00",
		X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"E0",X"77",X"0E",X"EE",X"E0",X"77",X"0E",X"00",X"E0",
		X"75",X"0D",X"00",X"E0",X"75",X"DD",X"00",X"E0",X"7F",X"DD",X"00",X"E0",X"5F",X"DD",X"00",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"EE",X"00",X"EE",X"00",X"0E",X"00",
		X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"0E",X"00",
		X"00",X"DD",X"0E",X"00",X"00",X"DD",X"E0",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",
		X"E0",X"2D",X"00",X"00",X"7E",X"2D",X"00",X"E0",X"77",X"25",X"00",X"E0",X"77",X"55",X"00",X"E0",
		X"77",X"5F",X"00",X"E0",X"77",X"FF",X"00",X"E0",X"77",X"75",X"00",X"E0",X"77",X"77",X"00",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"EE",X"00",X"EE",X"00",X"EE",X"00",
		X"E0",X"00",X"E0",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",
		X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",
		X"08",X"00",X"00",X"00",X"08",X"00",X"D0",X"E0",X"08",X"00",X"D0",X"E0",X"EE",X"00",X"D0",X"E0",
		X"77",X"00",X"0E",X"E0",X"77",X"55",X"E0",X"E0",X"77",X"FF",X"20",X"E0",X"77",X"55",X"20",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"B0",
		X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"40",
		X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",
		X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",
		X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"44",
		X"00",X"00",X"00",X"44",X"00",X"00",X"55",X"44",X"00",X"0B",X"55",X"44",X"00",X"BB",X"FF",X"44",
		X"00",X"B0",X"55",X"44",X"00",X"00",X"55",X"44",X"00",X"00",X"50",X"44",X"00",X"00",X"00",X"44",
		X"00",X"00",X"4B",X"AB",X"00",X"00",X"4B",X"BB",X"00",X"00",X"4B",X"B0",X"00",X"00",X"4B",X"00",
		X"00",X"00",X"40",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"40",X"00",
		X"00",X"00",X"4B",X"00",X"00",X"00",X"4B",X"B0",X"00",X"00",X"4B",X"BB",X"00",X"00",X"4B",X"AB",
		X"55",X"3F",X"77",X"77",X"35",X"3F",X"77",X"77",X"33",X"3F",X"77",X"77",X"33",X"3F",X"77",X"77",
		X"43",X"3F",X"77",X"00",X"44",X"3F",X"77",X"00",X"44",X"00",X"77",X"00",X"44",X"00",X"77",X"00",
		X"44",X"00",X"70",X"00",X"44",X"00",X"70",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",
		X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"04",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"04",X"00",X"00",X"00",
		X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",
		X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",
		X"B0",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",
		X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",
		X"F5",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",
		X"04",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",
		X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",
		X"44",X"00",X"70",X"00",X"44",X"00",X"77",X"00",X"44",X"3F",X"77",X"00",X"43",X"3F",X"77",X"77",
		X"33",X"3F",X"77",X"77",X"33",X"3F",X"77",X"77",X"35",X"3F",X"77",X"77",X"55",X"3F",X"77",X"77",
		X"44",X"4F",X"77",X"22",X"44",X"3F",X"77",X"22",X"44",X"3F",X"77",X"22",X"44",X"3F",X"77",X"22",
		X"44",X"3F",X"77",X"22",X"44",X"3F",X"77",X"00",X"44",X"3F",X"77",X"00",X"44",X"40",X"77",X"00",
		X"40",X"40",X"70",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"44",X"40",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"40",X"00",
		X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"24",X"00",X"77",X"77",X"24",X"00",X"77",X"77",X"24",X"00",X"77",X"77",X"24",X"00",X"77",X"77",
		X"24",X"00",X"77",X"77",X"24",X"00",X"F7",X"77",X"24",X"03",X"F7",X"77",X"24",X"03",X"F7",X"77",
		X"24",X"33",X"F7",X"77",X"24",X"33",X"F7",X"07",X"24",X"33",X"F7",X"07",X"24",X"33",X"F7",X"00",
		X"04",X"33",X"F7",X"00",X"04",X"33",X"30",X"00",X"44",X"33",X"30",X"00",X"44",X"53",X"00",X"00",
		X"44",X"55",X"00",X"00",X"43",X"53",X"00",X"00",X"43",X"33",X"00",X"00",X"43",X"33",X"00",X"00",
		X"43",X"33",X"00",X"00",X"BB",X"33",X"44",X"44",X"BB",X"34",X"44",X"44",X"6B",X"34",X"44",X"44",
		X"BB",X"44",X"44",X"44",X"6A",X"44",X"44",X"00",X"AA",X"44",X"40",X"00",X"AA",X"44",X"00",X"00",
		X"AA",X"04",X"00",X"00",X"4A",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"DD",X"00",X"00",X"77",X"0D",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",
		X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"E0",X"EE",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"EE",X"00",X"00",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",
		X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"EE",X"00",X"00",X"EE",X"EE",X"00",
		X"00",X"E0",X"EE",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",
		X"EE",X"00",X"00",X"00",X"E0",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"EE",
		X"E0",X"00",X"00",X"EE",X"0E",X"00",X"0E",X"EE",X"00",X"00",X"0E",X"EE",X"00",X"00",X"E0",X"EE",
		X"00",X"00",X"00",X"E0",X"00",X"D0",X"00",X"E0",X"00",X"DD",X"00",X"E0",X"00",X"DD",X"00",X"00",
		X"00",X"DD",X"00",X"00",X"77",X"DD",X"00",X"00",X"77",X"DD",X"00",X"00",X"75",X"DD",X"EE",X"00",
		X"33",X"44",X"00",X"00",X"33",X"44",X"44",X"BB",X"34",X"44",X"44",X"00",X"34",X"44",X"44",X"00",
		X"44",X"44",X"44",X"00",X"44",X"44",X"00",X"B0",X"44",X"44",X"00",X"BB",X"44",X"00",X"00",X"00",
		X"34",X"00",X"00",X"00",X"33",X"50",X"00",X"00",X"33",X"50",X"00",X"00",X"A3",X"00",X"E0",X"00",
		X"AB",X"00",X"0E",X"00",X"BB",X"00",X"00",X"00",X"BB",X"40",X"00",X"00",X"BB",X"44",X"00",X"00",
		X"66",X"44",X"00",X"00",X"66",X"44",X"EE",X"00",X"BB",X"44",X"5E",X"00",X"BB",X"44",X"55",X"00",
		X"BB",X"44",X"FF",X"00",X"BB",X"44",X"55",X"00",X"BB",X"00",X"5F",X"00",X"00",X"00",X"F5",X"00",
		X"00",X"00",X"F5",X"00",X"00",X"00",X"55",X"B0",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",
		X"BB",X"DD",X"00",X"00",X"BB",X"DD",X"00",X"00",X"B5",X"00",X"00",X"00",X"55",X"00",X"00",X"00",
		X"55",X"00",X"00",X"00",X"0F",X"77",X"00",X"00",X"05",X"77",X"00",X"00",X"00",X"77",X"00",X"00",
		X"00",X"EE",X"77",X"00",X"00",X"EE",X"77",X"00",X"0E",X"00",X"77",X"00",X"0E",X"00",X"77",X"00",
		X"EE",X"77",X"77",X"00",X"E0",X"77",X"77",X"00",X"E0",X"77",X"E7",X"00",X"E0",X"77",X"EE",X"00",
		X"E7",X"77",X"EE",X"00",X"77",X"77",X"EE",X"00",X"77",X"77",X"0E",X"00",X"77",X"7E",X"00",X"00",
		X"77",X"7E",X"00",X"00",X"77",X"E0",X"00",X"00",X"77",X"E0",X"00",X"00",X"33",X"00",X"00",X"00",
		X"33",X"00",X"EE",X"00",X"33",X"00",X"00",X"0B",X"33",X"00",X"00",X"B0",X"33",X"EE",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"44",X"40",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"40",X"00",
		X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"04",X"FF",X"00",X"00",X"44",X"FF",X"00",X"00",
		X"44",X"44",X"00",X"00",X"FF",X"44",X"50",X"00",X"44",X"44",X"50",X"00",X"44",X"44",X"55",X"00",
		X"44",X"44",X"55",X"00",X"44",X"44",X"55",X"00",X"44",X"44",X"50",X"00",X"44",X"44",X"40",X"00",
		X"44",X"44",X"00",X"00",X"54",X"45",X"00",X"00",X"05",X"55",X"00",X"00",X"00",X"55",X"00",X"E0",
		X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"06",X"66",X"00",X"00",X"06",X"66",X"00",X"00",
		X"66",X"66",X"00",X"00",X"66",X"66",X"60",X"00",X"66",X"66",X"60",X"00",X"6F",X"66",X"66",X"00",
		X"66",X"66",X"66",X"00",X"66",X"66",X"DD",X"00",X"66",X"66",X"D0",X"00",X"66",X"66",X"60",X"00",
		X"86",X"66",X"00",X"00",X"06",X"6D",X"00",X"00",X"08",X"DD",X"00",X"00",X"00",X"DD",X"00",X"E0",
		X"00",X"DD",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"CC",X"CC",X"00",X"00",X"AA",X"AA",X"00",X"0C",X"AA",X"AA",X"00",
		X"CC",X"CC",X"AA",X"00",X"CA",X"FF",X"CC",X"00",X"AA",X"FF",X"CC",X"00",X"AA",X"CC",X"AA",X"00",
		X"AA",X"CC",X"AA",X"00",X"AA",X"CC",X"AA",X"00",X"AA",X"CC",X"AA",X"00",X"AA",X"CC",X"CC",X"00",
		X"AA",X"FF",X"CC",X"00",X"AA",X"FF",X"AA",X"00",X"AA",X"CC",X"AA",X"00",X"AA",X"CC",X"AA",X"00",
		X"AA",X"CC",X"AA",X"00",X"AA",X"CC",X"CC",X"00",X"CA",X"CC",X"CC",X"00",X"CC",X"AA",X"AA",X"00",
		X"0C",X"AA",X"AA",X"00",X"00",X"AA",X"AA",X"00",X"00",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"CC",X"CC",X"00",X"00",X"66",X"66",X"00",X"0C",X"66",X"66",X"00",
		X"CC",X"CC",X"66",X"00",X"C6",X"FF",X"CC",X"00",X"66",X"FF",X"CC",X"00",X"66",X"CC",X"66",X"00",
		X"66",X"CC",X"66",X"00",X"66",X"CC",X"66",X"00",X"66",X"CC",X"66",X"00",X"66",X"CC",X"CC",X"00",
		X"66",X"FF",X"CC",X"00",X"66",X"FF",X"66",X"00",X"66",X"CC",X"66",X"00",X"66",X"CC",X"66",X"00",
		X"66",X"CC",X"66",X"00",X"66",X"CC",X"CC",X"00",X"C6",X"CC",X"CC",X"00",X"CC",X"66",X"66",X"00",
		X"0C",X"66",X"66",X"00",X"00",X"66",X"66",X"00",X"00",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"CC",X"CC",X"00",X"00",X"BB",X"BB",X"00",X"0C",X"BB",X"BB",X"00",
		X"CC",X"CC",X"BB",X"00",X"CB",X"FF",X"CC",X"00",X"BB",X"FF",X"CC",X"00",X"BB",X"CC",X"BB",X"00",
		X"BB",X"CC",X"BB",X"00",X"BB",X"CC",X"BB",X"00",X"BB",X"CC",X"BB",X"00",X"BB",X"CC",X"CC",X"00",
		X"BB",X"FF",X"CC",X"00",X"BB",X"FF",X"BB",X"00",X"BB",X"CC",X"BB",X"00",X"BB",X"CC",X"BB",X"00",
		X"BB",X"CC",X"BB",X"00",X"BB",X"CC",X"CC",X"00",X"CB",X"CC",X"CC",X"00",X"CC",X"BB",X"BB",X"00",
		X"0C",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"00",X"00",
		X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"0A",X"FF",X"00",X"00",X"AA",X"FF",X"00",X"00",
		X"AA",X"FA",X"00",X"00",X"AF",X"AA",X"A0",X"00",X"FF",X"AA",X"A0",X"00",X"AA",X"AA",X"9A",X"00",
		X"AA",X"AA",X"AA",X"00",X"AA",X"AA",X"9A",X"00",X"AA",X"AA",X"90",X"00",X"AA",X"AA",X"A0",X"00",
		X"AA",X"A9",X"00",X"00",X"AA",X"99",X"00",X"00",X"0A",X"99",X"00",X"00",X"00",X"99",X"00",X"E0",
		X"00",X"99",X"00",X"00",X"00",X"A9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"0A",X"05",X"00",
		X"00",X"70",X"50",X"00",X"00",X"4A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"06",X"55",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"40",X"A0",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"04",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"66",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"A6",X"00",X"00",X"00",X"F6",X"00",X"00",X"0F",X"F6",X"00",X"00",
		X"00",X"FA",X"00",X"00",X"00",X"0A",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",
		X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"04",X"00",X"F5",X"04",X"40",X"00",X"00",X"04",X"00",X"00",X"00",X"A4",X"00",X"00",
		X"00",X"A4",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"6A",X"00",X"00",X"00",X"F6",X"00",X"00",
		X"04",X"46",X"00",X"00",X"00",X"66",X"44",X"00",X"00",X"04",X"00",X"00",X"00",X"05",X"00",X"00",
		X"00",X"05",X"00",X"00",X"05",X"00",X"00",X"00",X"55",X"50",X"00",X"00",X"0A",X"50",X"00",X"00",
		X"0A",X"50",X"A0",X"00",X"0A",X"40",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"44",X"40",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"04",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"04",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"40",X"00",
		X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"04",X"00",X"44",X"00",
		X"04",X"00",X"44",X"00",X"04",X"40",X"44",X"00",X"04",X"40",X"44",X"00",X"04",X"40",X"44",X"00",
		X"04",X"44",X"44",X"00",X"04",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"40",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"99",X"00",X"00",X"9A",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"09",X"9A",X"99",X"00",X"B9",X"99",X"99",X"00",
		X"09",X"9A",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"9A",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"90",X"00",
		X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"04",X"00",X"44",X"00",
		X"04",X"00",X"44",X"00",X"04",X"00",X"44",X"00",X"04",X"44",X"44",X"00",X"04",X"44",X"44",X"00",
		X"04",X"44",X"44",X"00",X"04",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"40",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"66",X"00",
		X"00",X"66",X"AA",X"00",X"00",X"6A",X"AA",X"00",X"00",X"6A",X"6A",X"00",X"00",X"6A",X"6A",X"00",
		X"00",X"6A",X"6A",X"00",X"00",X"6A",X"6A",X"00",X"00",X"AA",X"AA",X"00",X"00",X"AA",X"AA",X"00",
		X"00",X"66",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"66",X"06",X"00",X"00",X"AA",X"6A",X"00",X"00",X"AA",X"6A",X"00",
		X"00",X"66",X"6A",X"00",X"00",X"06",X"6A",X"00",X"00",X"06",X"6A",X"00",X"00",X"00",X"6A",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"66",X"00",
		X"00",X"66",X"AA",X"00",X"00",X"6A",X"AA",X"00",X"00",X"6A",X"6A",X"00",X"00",X"6A",X"6A",X"00",
		X"00",X"6A",X"6A",X"00",X"00",X"6A",X"6A",X"00",X"00",X"AA",X"AA",X"00",X"00",X"AA",X"AA",X"00",
		X"00",X"66",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"00",X"00",X"AA",X"AA",X"00",
		X"00",X"AA",X"AA",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"0A",X"00",
		X"00",X"00",X"0A",X"00",X"00",X"AA",X"AA",X"00",X"00",X"AA",X"AA",X"00",X"00",X"66",X"66",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"6A",X"00",X"00",X"66",X"6A",X"00",X"00",X"AA",X"AA",X"00",
		X"00",X"AA",X"AA",X"00",X"00",X"66",X"6A",X"00",X"00",X"A6",X"6A",X"00",X"00",X"A6",X"66",X"00",
		X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"66",X"00",X"00",X"66",X"AA",X"00",
		X"00",X"6A",X"AA",X"00",X"00",X"6A",X"6A",X"00",X"00",X"6A",X"6A",X"00",X"00",X"6A",X"6A",X"00",
		X"00",X"6A",X"6A",X"00",X"00",X"AA",X"AA",X"00",X"00",X"AA",X"AA",X"00",X"00",X"66",X"66",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"6A",X"00",X"00",X"66",X"6A",X"00",X"00",X"AA",X"AA",X"00",
		X"00",X"AA",X"AA",X"00",X"00",X"66",X"6A",X"00",X"00",X"A6",X"6A",X"00",X"00",X"A6",X"66",X"00",
		X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"00",
		X"00",X"AA",X"6A",X"00",X"00",X"AA",X"6A",X"00",X"00",X"66",X"6A",X"00",X"00",X"06",X"6A",X"00",
		X"00",X"00",X"6A",X"00",X"00",X"00",X"6A",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"60",X"00",X"00",X"A6",X"60",X"00",
		X"00",X"AA",X"60",X"00",X"00",X"6A",X"60",X"00",X"00",X"66",X"00",X"00",X"00",X"06",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"6A",X"60",X"00",X"00",X"AA",X"60",X"00",X"00",X"A6",X"60",X"00",
		X"00",X"66",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"00",
		X"00",X"AA",X"AA",X"00",X"00",X"AA",X"AA",X"00",X"00",X"66",X"6A",X"00",X"00",X"06",X"6A",X"00",
		X"00",X"06",X"6A",X"00",X"00",X"06",X"6A",X"00",X"00",X"06",X"AA",X"00",X"00",X"00",X"AA",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"60",X"00",X"00",X"A6",X"60",X"00",
		X"00",X"AA",X"60",X"00",X"00",X"6A",X"60",X"00",X"00",X"66",X"00",X"00",X"00",X"06",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"6A",X"60",X"00",X"00",X"AA",X"60",X"00",X"00",X"A6",X"60",X"00",
		X"00",X"66",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"06",X"66",X"66",X"00",X"06",X"AA",X"AA",X"00",X"06",X"AA",X"AA",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",
		X"00",X"AA",X"00",X"00",X"00",X"6A",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"06",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"60",X"00",X"00",X"A6",X"60",X"00",
		X"00",X"AA",X"60",X"00",X"00",X"6A",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"06",X"00",X"00",
		X"00",X"06",X"00",X"00",X"00",X"6A",X"60",X"00",X"00",X"AA",X"60",X"00",X"00",X"A6",X"60",X"00",
		X"00",X"66",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"66",X"00",
		X"00",X"66",X"AA",X"00",X"00",X"6A",X"AA",X"00",X"00",X"6A",X"6A",X"00",X"00",X"6A",X"6A",X"00",
		X"00",X"6A",X"6A",X"00",X"00",X"6A",X"6A",X"00",X"00",X"AA",X"AA",X"00",X"00",X"AA",X"AA",X"00",
		X"00",X"66",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"60",X"00",X"00",X"A6",X"60",X"00",
		X"00",X"AA",X"60",X"00",X"00",X"6A",X"60",X"00",X"00",X"66",X"00",X"00",X"00",X"06",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"6A",X"60",X"00",X"00",X"AA",X"60",X"00",X"00",X"A6",X"60",X"00",
		X"00",X"66",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"CC",X"CC",X"00",X"00",X"55",X"55",X"00",X"0C",X"55",X"55",X"00",
		X"CC",X"CC",X"55",X"00",X"C5",X"FF",X"CC",X"00",X"55",X"FF",X"CC",X"00",X"55",X"CC",X"55",X"00",
		X"55",X"CC",X"55",X"00",X"55",X"CC",X"55",X"00",X"55",X"CC",X"55",X"00",X"55",X"CC",X"CC",X"00",
		X"55",X"FF",X"CC",X"00",X"55",X"FF",X"55",X"00",X"55",X"CC",X"55",X"00",X"55",X"CC",X"55",X"00",
		X"55",X"CC",X"55",X"00",X"55",X"CC",X"CC",X"00",X"C5",X"CC",X"CC",X"00",X"CC",X"55",X"55",X"00",
		X"0C",X"55",X"55",X"00",X"00",X"55",X"55",X"00",X"00",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
