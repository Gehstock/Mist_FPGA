library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity travusa_chr_bit3 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of travusa_chr_bit3 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"00",X"00",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",
		X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"00",X"00",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"00",X"00",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"02",X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"00",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"3F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"40",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"BF",X"3F",X"7F",X"7F",X"7F",X"01",X"81",X"FF",X"81",X"01",X"7F",X"7F",X"7F",X"01",X"81",
		X"FF",X"01",X"01",X"E3",X"C7",X"E3",X"01",X"01",X"FF",X"01",X"01",X"DD",X"DD",X"DD",X"C1",X"E3",
		X"FF",X"FF",X"F3",X"3E",X"00",X"00",X"00",X"00",X"FF",X"FF",X"F9",X"67",X"00",X"00",X"00",X"00",
		X"3F",X"9F",X"9B",X"8E",X"00",X"00",X"00",X"00",X"FD",X"FE",X"CE",X"72",X"00",X"00",X"01",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"1C",X"1C",X"0C",X"08",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"A0",X"B0",X"F0",X"F8",X"78",X"E8",X"E8",X"B0",
		X"F0",X"E0",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0F",X"0F",X"0F",
		X"07",X"03",X"0B",X"0F",X"0F",X"05",X"05",X"05",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"C4",X"C7",X"BF",X"1F",X"3F",X"0F",X"0F",X"00",X"01",X"03",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"C0",X"BC",X"1E",X"3F",X"0F",X"0F",X"00",X"01",X"03",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"7F",X"1F",X"3F",X"0F",X"0F",X"27",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"7C",X"1E",X"3F",X"0F",X"0F",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"C0",X"80",X"C0",X"C0",X"C0",X"00",X"80",X"27",X"1F",X"1B",X"0E",X"00",X"00",X"00",X"00",
		X"CE",X"D7",X"DF",X"DE",X"DF",X"CF",X"EF",X"E7",X"F7",X"F5",X"F3",X"FB",X"FB",X"FB",X"FB",X"FB",
		X"FB",X"FB",X"FB",X"F3",X"F7",X"F7",X"E6",X"EE",X"CC",X"D4",X"DC",X"D8",X"D8",X"D8",X"98",X"A8",
		X"B8",X"B8",X"B8",X"98",X"DC",X"DC",X"DE",X"CE",X"EC",X"EE",X"EE",X"E6",X"EE",X"EE",X"EE",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"C0",X"C0",X"80",X"C0",X"C0",X"C0",X"C0",X"00",X"80",
		X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"04",X"07",X"07",X"07",X"07",X"07",X"07",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"01",X"01",X"01",X"02",X"03",X"03",X"03",X"04",X"07",X"0F",X"0F",X"1F",X"1B",X"0D",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3E",X"2F",X"1F",X"1F",X"1F",X"0B",X"0D",X"0F",X"0F",X"07",
		X"F7",X"F7",X"F7",X"F7",X"C7",X"F7",X"F7",X"77",X"F3",X"FB",X"FB",X"EB",X"D9",X"FD",X"FD",X"7D",
		X"B5",X"F9",X"FB",X"FB",X"FB",X"FB",X"EB",X"F3",X"F7",X"F7",X"E7",X"EF",X"CF",X"DF",X"DF",X"9F",
		X"BF",X"BF",X"BF",X"BF",X"9F",X"5F",X"DF",X"DF",X"DF",X"DF",X"CF",X"AF",X"EF",X"EF",X"E7",X"F7",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"DF",X"1F",X"8F",X"07",X"07",X"03",X"03",X"81",X"81",X"81",X"01",X"11",X"11",X"31",X"21",
		X"C0",X"81",X"C3",X"C0",X"C0",X"C0",X"00",X"80",X"00",X"C0",X"C0",X"BC",X"1E",X"3F",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"7C",X"1E",X"3F",X"0F",X"0F",X"06",X"00",
		X"03",X"03",X"07",X"07",X"07",X"07",X"0F",X"1F",X"80",X"81",X"03",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"C0",X"BC",X"1E",X"3F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"37",X"7F",X"1F",X"3F",X"0F",X"0F",X"07",X"05",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"3F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"6F",X"38",X"10",X"10",X"10",X"30",X"61",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"E3",X"81",X"01",X"01",X"01",X"01",X"01",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"60",X"F0",
		X"1C",X"00",X"01",X"01",X"01",X"03",X"06",X"04",X"00",X"00",X"00",X"01",X"81",X"03",X"C7",X"7F",
		X"1F",X"3F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"03",X"0E",X"08",X"80",X"C0",
		X"7E",X"30",X"18",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"1E",X"03",X"00",X"00",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"60",X"FC",X"01",X"01",X"01",X"03",
		X"06",X"64",X"C0",X"00",X"60",X"C1",X"83",X"FE",X"00",X"00",X"00",X"00",X"00",X"C8",X"1F",X"F9",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"A0",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"C0",X"E0",X"30",X"1C",X"16",X"00",X"00",X"03",X"00",X"00",X"80",X"80",X"08",X"48",X"CC",
		X"06",X"03",X"01",X"07",X"1C",X"00",X"C1",X"FF",X"08",X"08",X"08",X"1E",X"17",X"11",X"30",X"21",
		X"7F",X"18",X"0C",X"06",X"02",X"03",X"01",X"00",X"00",X"00",X"01",X"01",X"01",X"03",X"02",X"06",
		X"0C",X"08",X"08",X"1E",X"17",X"11",X"30",X"21",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"07",X"01",X"08",X"04",X"00",X"00",X"00",
		X"00",X"00",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0C",X"C4",X"04",X"04",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"C8",X"08",
		X"FF",X"FF",X"FC",X"80",X"00",X"06",X"80",X"80",X"F0",X"80",X"84",X"C4",X"40",X"60",X"20",X"20",
		X"7F",X"FF",X"FF",X"FF",X"FE",X"FC",X"F8",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"03",X"1F",X"7F",X"FF",X"FF",X"FE",X"F8",X"F0",X"91",X"11",X"18",X"08",X"C8",
		X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"3F",X"FF",X"FF",X"FE",X"EA",X"8B",X"09",
		X"FF",X"FF",X"FF",X"E0",X"04",X"22",X"40",X"00",X"FF",X"E0",X"AC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"24",X"46",X"6F",X"76",X"FE",X"FB",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"E0",X"E0",X"F0",X"A8",X"7C",X"52",X"FA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FB",X"FF",X"FF",X"FF",X"FF",X"7F",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"BC",X"FC",X"F8",X"F8",X"F0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"E0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"60",X"FC",X"FF",X"FF",X"FF",X"FF",X"E1",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"03",X"C7",X"F7",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F8",X"F8",X"3C",X"FC",X"9C",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"01",X"03",X"03",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"9F",X"FF",X"E7",X"FC",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CD",X"FD",X"FF",X"FF",X"FD",X"FD",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"F8",X"DC",X"5C",X"7C",X"FC",X"F0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"7F",X"9F",X"7F",X"FF",X"FF",X"7F",X"E7",X"FF",
		X"FE",X"F8",X"FF",X"FF",X"FB",X"F7",X"FE",X"FD",X"00",X"00",X"00",X"00",X"C0",X"C0",X"F0",X"F0",
		X"01",X"0F",X"FF",X"FF",X"FF",X"FF",X"F8",X"00",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",
		X"9F",X"FF",X"FF",X"FF",X"7B",X"39",X"00",X"00",X"BF",X"DE",X"7F",X"BF",X"FF",X"F8",X"F0",X"70",
		X"70",X"F0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"11",X"79",X"7F",
		X"01",X"13",X"BD",X"FF",X"CF",X"97",X"3E",X"3E",X"D8",X"FC",X"E0",X"8D",X"06",X"57",X"FF",X"F9",
		X"00",X"00",X"00",X"00",X"80",X"80",X"D0",X"F8",X"7E",X"FE",X"7E",X"FF",X"FF",X"7F",X"7F",X"FF",
		X"7F",X"3F",X"7F",X"7F",X"BF",X"FF",X"FF",X"FF",X"FC",X"F8",X"F1",X"E5",X"F7",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"7A",X"3F",X"BE",X"FE",X"FD",X"FF",X"FE",
		X"EF",X"1F",X"13",X"07",X"07",X"0F",X"0F",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FC",X"FE",X"FF",X"FF",X"FF",X"FE",X"FC",
		X"0F",X"07",X"02",X"01",X"03",X"01",X"00",X"00",X"FF",X"FF",X"FF",X"FB",X"FB",X"B9",X"3D",X"18",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EE",X"80",X"F8",X"F0",X"E0",X"E0",X"80",X"00",X"00",X"00",
		X"FF",X"FF",X"F8",X"C0",X"00",X"00",X"00",X"00",X"00",X"10",X"01",X"3F",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"18",X"00",X"01",X"FF",
		X"FF",X"FF",X"FE",X"F8",X"C0",X"00",X"00",X"00",X"00",X"90",X"91",X"87",X"FF",X"FF",X"BF",X"BE",
		X"00",X"00",X"00",X"00",X"10",X"18",X"09",X"8F",X"3F",X"7F",X"FF",X"FF",X"FE",X"F0",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"11",X"01",X"3F",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F0",X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",X"FC",X"FC",X"FC",X"FC",X"FE",X"FE",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"F8",X"F0",X"F0",X"F0",X"F4",X"F0",X"E0",X"E0",X"E0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"04",X"04",X"04",X"FC",X"FC",X"FC",X"FC",X"FE",X"FE",X"FE",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"04",X"4C",X"28",X"08",X"FC",X"FE",X"FF",
		X"00",X"00",X"00",X"40",X"82",X"04",X"01",X"FF",X"40",X"60",X"20",X"20",X"20",X"78",X"FE",X"FF",
		X"40",X"40",X"01",X"03",X"07",X"7F",X"FF",X"FF",X"7F",X"7F",X"7F",X"7F",X"3F",X"3F",X"3F",X"3F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"01",X"01",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"80",X"81",X"87",X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F0",X"C0",X"C0",X"C0",X"E0",X"E0",X"E0",X"E0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F0",X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FC",X"FC",X"FC",X"FC",X"FE",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C0",X"C0",X"C0",X"C0",X"E0",X"E0",X"E0",X"E0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C0",X"00",X"00",
		X"C0",X"80",X"88",X"90",X"83",X"9F",X"FF",X"FF",X"FF",X"FF",X"FE",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"0C",X"04",X"64",X"05",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"01",X"83",
		X"87",X"0F",X"FF",X"FF",X"FF",X"FF",X"FC",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"88",X"C8",X"43",X"5F",X"FF",X"FF",
		X"FF",X"FF",X"FE",X"F8",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"0C",X"C4",X"04",X"05",X"FF",X"BF",X"BF",X"BF",X"BE",
		X"F0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"0C",X"00",X"83",
		X"87",X"0F",X"FF",X"FF",X"FC",X"F0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"10",X"90",X"83",X"9F",X"FF",X"FF",X"FF",X"FC",X"E0",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"12",X"12",X"18",X"0B",X"8F",X"3F",X"FF",X"FF",X"FF",X"F8",X"E0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"03",X"05",X"00",X"00",X"02",X"04",X"03",X"FF",
		X"FF",X"FF",X"FF",X"7F",X"07",X"7F",X"FF",X"FF",X"FE",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FC",X"F0",X"F0",X"E0",X"E0",X"C0",X"FF",X"FF",X"FF",X"00",X"AA",X"00",X"AA",X"00",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"47",X"10",X"FE",X"FF",X"F0",X"FB",X"E0",X"FB",X"C0",X"FF",
		X"00",X"10",X"00",X"10",X"00",X"18",X"B9",X"B9",X"00",X"6D",X"00",X"6D",X"00",X"6D",X"00",X"FF",
		X"FF",X"C7",X"83",X"83",X"83",X"83",X"C7",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"07",X"03",X"07",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"9F",X"FF",X"FF",X"FE",X"FC",X"F8",X"F0",X"00",X"00",
		X"78",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"7F",X"2E",X"40",X"2E",X"40",X"3E",X"9F",
		X"FF",X"FF",X"7F",X"3F",X"1F",X"7F",X"FF",X"FF",X"03",X"07",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"03",X"05",X"00",X"00",X"02",X"04",X"00",X"00",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"FF",X"02",X"04",X"00",X"00",X"02",X"04",X"03",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"05",X"00",X"00",X"02",X"04",X"03",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"07",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"87",X"FF",
		X"07",X"FF",X"E7",X"E7",X"E7",X"E7",X"E7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"DF",X"8F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"03",X"05",X"00",X"00",X"02",X"04",X"03",X"FF",
		X"03",X"07",X"03",X"01",X"03",X"07",X"03",X"FF",X"FE",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"FE",X"FC",X"F0",X"F0",X"E0",X"E0",X"C0",X"FF",X"03",X"07",X"03",X"01",X"03",X"07",X"03",X"01",
		X"EF",X"FF",X"E8",X"FF",X"FF",X"FF",X"FF",X"FF",X"03",X"07",X"03",X"01",X"03",X"07",X"03",X"FF",
		X"FE",X"FC",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"FC",X"F0",X"F0",X"E0",X"E0",X"C0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"00",X"FF",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"FF",
		X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"FF",X"FE",X"FE",X"00",X"AA",X"00",X"AA",X"00",X"00",
		X"FA",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"EF",X"F8",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"03",X"05",X"00",X"00",X"02",X"04",X"03",X"FF",
		X"FE",X"FC",X"00",X"00",X"00",X"00",X"00",X"FF",X"03",X"07",X"03",X"01",X"03",X"07",X"03",X"FF",
		X"03",X"07",X"03",X"01",X"03",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"03",X"05",X"00",X"00",X"00",X"04",X"03",X"FF",X"03",X"07",X"03",X"01",X"03",X"07",X"03",X"FF",
		X"FE",X"FC",X"F0",X"F0",X"E0",X"E0",X"C0",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"FE",X"FC",X"F0",X"F0",X"E0",X"E0",X"C0",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"7F",X"1F",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FE",X"FC",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"03",X"01",X"00",X"12",X"03",X"03",X"FF",X"FF",X"FF",X"FF",X"70",X"18",X"8A",X"FF",
		X"FF",X"FF",X"E0",X"1E",X"03",X"31",X"1C",X"07",X"FF",X"FF",X"7E",X"1F",X"8F",X"CF",X"CF",X"EE",
		X"FC",X"02",X"7F",X"FF",X"FF",X"FF",X"FF",X"3F",X"DF",X"47",X"6F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"03",X"43",X"D7",X"DF",X"7F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"9F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EE",X"FF",X"FF",X"7F",X"BF",X"9F",X"EF",X"F7",
		X"BF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",
		X"01",X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"19",X"14",X"05",X"15",X"15",X"15",X"11",
		X"1F",X"9C",X"9B",X"11",X"14",X"04",X"48",X"48",X"FF",X"1F",X"63",X"81",X"00",X"0C",X"12",X"1A",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"10",X"D0",X"D0",X"10",X"D0",X"D5",X"15",X"D5",
		X"48",X"44",X"44",X"44",X"08",X"18",X"40",X"40",X"00",X"06",X"09",X"06",X"00",X"0F",X"08",X"00",
		X"3F",X"0F",X"0F",X"07",X"07",X"03",X"03",X"03",X"0F",X"09",X"06",X"00",X"0F",X"0D",X"08",X"00",
		X"1E",X"08",X"1E",X"00",X"81",X"62",X"1C",X"C1",X"00",X"00",X"03",X"07",X"07",X"0F",X"1E",X"1E",
		X"00",X"E0",X"F8",X"FE",X"FF",X"0F",X"07",X"07",X"1A",X"16",X"1E",X"DE",X"DC",X"1C",X"DC",X"D2",
		X"05",X"06",X"07",X"07",X"03",X"03",X"03",X"00",X"1C",X"DC",X"DC",X"1E",X"DE",X"D6",X"1A",X"1E",
		X"03",X"03",X"03",X"07",X"07",X"06",X"05",X"07",X"FF",X"1F",X"0F",X"0F",X"0F",X"0E",X"0C",X"0C",
		X"FF",X"FF",X"FF",X"FF",X"0F",X"47",X"93",X"AB",X"1E",X"1F",X"17",X"17",X"1B",X"1C",X"0F",X"09",
		X"07",X"0F",X"FF",X"FE",X"F8",X"E4",X"1C",X"FC",X"0C",X"0C",X"0C",X"08",X"08",X"0C",X"0C",X"0C",
		X"4B",X"03",X"D3",X"07",X"F7",X"07",X"EF",X"4F",X"DF",X"13",X"DF",X"17",X"1E",X"1F",X"0C",X"0F",
		X"94",X"F4",X"24",X"E4",X"44",X"C2",X"81",X"84",X"0D",X"0C",X"0E",X"0F",X"0F",X"17",X"E7",X"0F",
		X"2F",X"8F",X"5F",X"1F",X"FF",X"FF",X"FF",X"FF",X"07",X"07",X"07",X"07",X"FF",X"FF",X"40",X"18",
		X"01",X"02",X"04",X"08",X"13",X"04",X"0B",X"10",X"FF",X"07",X"00",X"F3",X"01",X"01",X"84",X"78",
		X"03",X"09",X"DC",X"9A",X"DA",X"EA",X"7C",X"3D",X"06",X"00",X"03",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"31",X"D7",X"11",X"00",X"E0",X"0B",X"01",X"00",X"27",X"52",X"27",X"00",X"00",
		X"FF",X"FF",X"7F",X"7F",X"1F",X"7B",X"4F",X"77",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"60",
		X"07",X"07",X"63",X"91",X"00",X"E0",X"50",X"E0",X"00",X"60",X"60",X"00",X"60",X"60",X"00",X"60",
		X"00",X"A0",X"50",X"00",X"F0",X"00",X"F0",X"60",X"FF",X"FF",X"9F",X"1F",X"9F",X"6F",X"9F",X"FF",
		X"F0",X"00",X"60",X"90",X"60",X"01",X"02",X"00",X"FF",X"FF",X"BF",X"3F",X"7F",X"9F",X"7F",X"0F",
		X"00",X"00",X"00",X"01",X"00",X"03",X"00",X"06",X"E2",X"01",X"04",X"C4",X"22",X"23",X"65",X"65",
		X"0F",X"FF",X"7F",X"9F",X"7F",X"3F",X"BF",X"FF",X"30",X"08",X"08",X"04",X"04",X"04",X"08",X"00",
		X"E6",X"EF",X"7E",X"7E",X"3E",X"3F",X"1F",X"1F",X"9F",X"0E",X"0C",X"08",X"98",X"FC",X"FF",X"FF",
		X"FF",X"FF",X"7F",X"7F",X"77",X"E3",X"C3",X"C3",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F3",X"E3",X"C7",X"C1",X"81",X"82",X"81",X"80",X"E7",X"FF",X"FF",X"7D",X"58",X"50",X"50",X"41",
		X"00",X"10",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"60",X"60",X"00",X"07",
		X"81",X"C7",X"C2",X"E0",X"F0",X"F1",X"F7",X"FF",X"9F",X"3F",X"7F",X"F7",X"E3",X"C3",X"C3",X"E7",
		X"01",X"01",X"03",X"03",X"03",X"07",X"07",X"07",X"F3",X"F8",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F0",X"F0",X"18",X"C8",X"E0",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"80",X"E0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"C7",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"0F",X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FC",X"3F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"C0",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"80",X"80",X"80",X"80",X"C0",X"C0",X"C0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"C0",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"0F",X"0F",
		X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F8",X"DB",X"C3",X"C3",X"C3",X"C3",X"C3",X"C3",X"C3",
		X"0F",X"0F",X"0F",X"0F",X"07",X"07",X"07",X"07",X"F8",X"F8",X"F8",X"F8",X"F8",X"FC",X"FC",X"FC",
		X"C3",X"F3",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"07",X"07",X"03",X"03",X"03",X"03",X"03",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"FC",X"FC",X"FE",X"B6",X"86",X"86",X"86",
		X"01",X"01",X"01",X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"F0",X"FC",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"78",X"78",X"78",X"38",X"38",X"78",X"78",X"78",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"7F",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"86",X"87",X"87",X"87",X"87",X"E7",X"FF",X"FE",X"FE",X"FE",X"FE",X"FC",X"FC",X"FC",X"FC",X"F8",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"3F",X"3F",X"8E",X"E0",X"FF",
		X"00",X"CF",X"E3",X"38",X"FF",X"FF",X"00",X"FF",X"00",X"FF",X"FF",X"00",X"CF",X"E3",X"F8",X"FF",
		X"00",X"F3",X"F8",X"FE",X"FF",X"FF",X"FF",X"FF",X"00",X"0F",X"03",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"FC",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"C7",X"F1",X"FC",X"FF",X"FF",X"FF",X"FF",
		X"00",X"F3",X"F8",X"FE",X"FF",X"FF",X"FF",X"FF",X"00",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"36",X"30",
		X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"3C",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"F0",X"7C",X"FF",X"3E",X"00",X"FF",X"00",X"00",X"3F",X"1E",X"1F",X"1C",X"1C",
		X"FF",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1C",X"1C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"04",X"04",X"04",X"04",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"78",X"78",X"78",X"F8",X"F8",X"78",X"78",X"F8",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"7F",X"1F",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"0F",X"1F",X"7F",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"1F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"0F",X"1F",X"7F",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"1F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"03",X"0F",X"1F",X"7F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"07",X"1F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"0F",X"1F",X"7F",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"0F",X"1F",X"7F",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"0F",X"1F",X"7F",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"0F",X"1F",X"7F",X"FF",X"FF",
		X"00",X"01",X"03",X"0F",X"1F",X"7F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"07",X"1F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"03",X"0F",X"1F",X"7F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"0F",X"1F",X"7F",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"0F",X"1F",X"7F",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"1F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"3F",X"00",X"01",X"03",X"0F",X"1F",X"7F",X"FF",X"FF",
		X"07",X"1F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"1F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"01",X"03",X"0F",X"1F",X"7F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"03",X"0F",X"1F",X"7F",X"FF",X"FF",X"00",X"01",X"03",X"0F",X"1F",X"7F",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"01",X"01",X"03",X"0F",X"1F",X"7F",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"01",X"03",X"0F",X"1F",X"7F",X"FF",X"FF",
		X"07",X"1F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"03",X"0F",X"1F",X"7F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"07",X"1F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"01",X"03",X"0F",X"1F",X"7F",X"FF",X"FF",
		X"00",X"01",X"03",X"0F",X"1F",X"7F",X"FF",X"FF",X"01",X"01",X"03",X"0F",X"1F",X"7F",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"3F",X"00",X"01",X"03",X"0F",X"1F",X"7F",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"1F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"01",X"03",X"0F",X"1F",X"7F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"07",X"1F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"3F",
		X"00",X"01",X"03",X"0F",X"1F",X"7F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"1F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"1F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"0F",X"1F",X"7F",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"3F",X"00",X"01",X"03",X"0F",X"1F",X"7F",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"3F",
		X"00",X"01",X"03",X"0F",X"1F",X"7F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"3F",
		X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"03",X"0F",X"1F",X"7F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"3F",
		X"00",X"01",X"03",X"0F",X"1F",X"7F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"3F",
		X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"3F",X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"3F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"3F",
		X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FD",X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"3F",X"0E",X"0C",X"00",X"0C",X"02",X"0E",X"02",
		X"FF",X"BF",X"BF",X"3F",X"BF",X"3F",X"BE",X"BE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"3F",X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"3F",
		X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"0F",X"1F",X"7F",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"4E",X"52",X"5E",X"7F",X"FF",X"F1",X"C0",X"2A",
		X"3F",X"BF",X"BF",X"FF",X"FF",X"60",X"00",X"AA",X"40",X"E0",X"E0",X"F0",X"A8",X"7C",X"52",X"FA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"70",X"3B",X"9F",X"CF",X"CF",X"EE",X"FF",X"FF",X"FF",X"FF",X"1F",X"CF",X"E7",X"33",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BE",X"7E",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"5F",X"47",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"63",X"81",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"81",X"62",X"1C",X"C1",X"00",X"E0",X"F8",X"FE",X"FF",X"0F",X"67",X"97",
		X"05",X"E6",X"57",X"E7",X"03",X"A3",X"53",X"00",X"F3",X"03",X"F3",X"67",X"F7",X"06",X"65",X"97",
		X"67",X"0F",X"FF",X"FE",X"F8",X"E4",X"1C",X"FC",X"FF",X"FF",X"77",X"47",X"03",X"43",X"47",X"77",
		X"9F",X"0E",X"0C",X"08",X"98",X"FC",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"77",X"E3",X"C3",X"C3",
		X"E7",X"FF",X"FF",X"7D",X"58",X"50",X"50",X"41",X"9F",X"3F",X"7F",X"F7",X"E3",X"C3",X"C3",X"E7",
		X"F0",X"F0",X"18",X"C8",X"E0",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"09",X"0D",X"00",X"0E",
		X"00",X"00",X"18",X"18",X"3C",X"3C",X"3C",X"3C",X"05",X"0E",X"40",X"4B",X"2D",X"20",X"18",X"00",
		X"3C",X"3C",X"7C",X"7C",X"3C",X"3C",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"0D",X"0F",X"0C",X"1C",X"B9",X"BF",X"FF",X"F7",X"A0",X"80",
		X"38",X"F0",X"F0",X"C0",X"C7",X"FF",X"A7",X"03",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"C0",
		X"1F",X"1F",X"3F",X"3E",X"3E",X"3F",X"7F",X"7F",X"80",X"00",X"00",X"02",X"83",X"87",X"05",X"0D",
		X"07",X"2F",X"BA",X"F0",X"E0",X"E1",X"C3",X"C3",X"E0",X"F0",X"38",X"18",X"C0",X"E0",X"C0",X"F4",
		X"7E",X"7E",X"7F",X"7F",X"3F",X"3F",X"2F",X"0F",X"0C",X"0C",X"1E",X"9E",X"8F",X"DF",X"DF",X"DD",
		X"E7",X"C6",X"CC",X"EC",X"FE",X"DE",X"9B",X"19",X"0E",X"1F",X"07",X"0C",X"00",X"08",X"5C",X"F0",
		X"0F",X"0F",X"0F",X"0B",X"03",X"01",X"01",X"00",X"FD",X"F9",X"F9",X"FC",X"EC",X"E4",X"F4",X"E8",
		X"58",X"CC",X"EF",X"FD",X"7E",X"3B",X"39",X"08",X"D8",X"00",X"30",X"98",X"00",X"00",X"80",X"C0",
		X"00",X"00",X"00",X"00",X"01",X"02",X"02",X"04",X"07",X"18",X"60",X"80",X"00",X"00",X"00",X"00",
		X"C0",X"30",X"08",X"06",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"60",X"10",X"08",
		X"04",X"04",X"04",X"08",X"08",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"04",X"02",X"02",X"02",X"01",X"01",X"01",
		X"08",X"08",X"08",X"08",X"08",X"08",X"04",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"02",
		X"04",X"02",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"87",X"78",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"60",X"1C",X"03",X"02",X"02",X"02",X"04",X"04",X"08",X"10",X"E0",
		X"00",X"00",X"00",X"00",X"10",X"38",X"38",X"11",X"00",X"00",X"40",X"60",X"60",X"20",X"0F",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"10",X"80",X"E0",X"03",X"07",X"07",X"0F",X"0F",X"0F",X"1F",X"3F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"F8",X"FC",X"FC",X"FC",X"FC",X"F9",X"F8",
		X"7E",X"7E",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F8",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"7F",X"1F",X"0F",X"03",X"01",X"20",X"00",X"18",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"01",X"00",X"F8",X"FC",X"FE",X"FE",X"FE",X"FE",X"FC",X"70",
		X"00",X"00",X"01",X"00",X"30",X"30",X"10",X"03",X"00",X"00",X"00",X"60",X"60",X"42",X"00",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"07",X"4F",X"1F",X"3F",X"7F",X"7F",X"7F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"40",X"70",X"F8",X"7C",X"7E",X"7F",X"7F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"E3",X"F3",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"F8",X"7F",X"3F",X"3F",X"1F",X"5F",X"07",X"11",X"00",
		X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7E",X"FC",X"FC",X"FC",X"FC",X"FD",X"F9",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"C0",X"20",X"18",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"07",X"0E",X"1C",X"1C",X"38",X"00",X"E0",X"80",X"00",X"3F",X"7F",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"F0",X"F8",X"FC",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"39",X"71",X"73",X"73",X"73",X"E3",X"E7",X"E7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"E7",X"E7",X"E7",X"E7",X"E7",X"E7",X"E7",X"E7",X"FF",X"FF",X"F9",X"F8",X"F9",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"9F",X"0F",X"9F",X"FF",X"FF",X"FF",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"00",X"60",X"FC",X"FF",X"FF",X"FF",X"FF",X"E1",X"01",X"01",X"03",X"C7",X"F7",X"FF",X"FF",X"FF",
		X"F0",X"F0",X"F8",X"F8",X"3C",X"FC",X"9C",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"70",
		X"00",X"00",X"00",X"01",X"03",X"13",X"7B",X"7F",X"01",X"13",X"BD",X"FF",X"CF",X"97",X"3E",X"3E",
		X"D8",X"FC",X"E0",X"8D",X"06",X"57",X"FF",X"F9",X"00",X"00",X"00",X"00",X"80",X"80",X"D0",X"F8",
		X"01",X"01",X"01",X"00",X"00",X"00",X"FF",X"FF",X"9F",X"FF",X"FF",X"FF",X"7B",X"39",X"FF",X"FF",
		X"BF",X"DE",X"7F",X"BF",X"FF",X"F8",X"FF",X"FF",X"70",X"F0",X"E0",X"C0",X"80",X"00",X"FF",X"FF",
		X"0F",X"07",X"02",X"01",X"03",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",X"FB",X"B9",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"F0",X"E0",X"E0",X"80",X"00",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
