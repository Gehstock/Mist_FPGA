-- generated with romgen by MikeJ
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ROM_SND_1 is
  port (
    CLK         : in    std_logic;
    ADDR        : in    std_logic_vector(10 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_SND_1 is


  type ROM_ARRAY is array(0 to 2047) of std_logic_vector(7 downto 0);
  constant ROM : ROM_ARRAY := (
    x"FE",x"0F",x"20",x"05",x"21",x"26",x"80",x"36", -- 0x0000
    x"00",x"47",x"CD",x"86",x"04",x"18",x"EA",x"CD", -- 0x0008
    x"10",x"05",x"D6",x"05",x"20",x"05",x"21",x"26", -- 0x0010
    x"80",x"36",x"00",x"47",x"CD",x"86",x"04",x"3A", -- 0x0018
    x"26",x"80",x"FE",x"00",x"20",x"D3",x"3A",x"27", -- 0x0020
    x"80",x"FE",x"44",x"20",x"CC",x"3E",x"FF",x"C9", -- 0x0028
    x"CD",x"7D",x"08",x"B7",x"20",x"02",x"18",x"C1", -- 0x0030
    x"21",x"26",x"80",x"36",x"02",x"18",x"BA",x"CD", -- 0x0038
    x"44",x"08",x"18",x"B5",x"CD",x"7D",x"08",x"B7", -- 0x0040
    x"C8",x"ED",x"5B",x"24",x"80",x"1A",x"32",x"23", -- 0x0048
    x"80",x"13",x"1A",x"6F",x"13",x"1A",x"67",x"13", -- 0x0050
    x"ED",x"53",x"24",x"80",x"CD",x"12",x"04",x"21", -- 0x0058
    x"27",x"80",x"34",x"21",x"26",x"80",x"36",x"01", -- 0x0060
    x"C9",x"CD",x"7D",x"08",x"B7",x"C8",x"3E",x"01", -- 0x0068
    x"32",x"23",x"80",x"21",x"27",x"80",x"34",x"21", -- 0x0070
    x"26",x"80",x"36",x"02",x"C9",x"21",x"22",x"80", -- 0x0078
    x"35",x"20",x"0C",x"3E",x"0B",x"77",x"21",x"23", -- 0x0080
    x"80",x"35",x"20",x"03",x"3E",x"FF",x"C9",x"AF", -- 0x0088
    x"C9",x"01",x"15",x"01",x"01",x"15",x"01",x"0B", -- 0x0090
    x"15",x"01",x"01",x"15",x"01",x"01",x"15",x"01", -- 0x0098
    x"03",x"15",x"01",x"03",x"4A",x"01",x"03",x"A0", -- 0x00A0
    x"01",x"03",x"4A",x"01",x"03",x"15",x"01",x"03", -- 0x00A8
    x"4A",x"01",x"03",x"15",x"01",x"03",x"D0",x"00", -- 0x00B0
    x"03",x"15",x"01",x"03",x"4A",x"01",x"03",x"A0", -- 0x00B8
    x"01",x"03",x"4A",x"01",x"03",x"15",x"01",x"03", -- 0x00C0
    x"4A",x"01",x"03",x"15",x"01",x"03",x"D0",x"00", -- 0x00C8
    x"0B",x"15",x"01",x"01",x"15",x"01",x"01",x"15", -- 0x00D0
    x"01",x"0B",x"15",x"01",x"01",x"15",x"01",x"01", -- 0x00D8
    x"15",x"01",x"0B",x"15",x"01",x"01",x"15",x"01", -- 0x00E0
    x"01",x"15",x"01",x"0B",x"15",x"01",x"01",x"15", -- 0x00E8
    x"01",x"01",x"15",x"01",x"20",x"15",x"01",x"3E", -- 0x00F0
    x"20",x"32",x"29",x"80",x"3E",x"08",x"32",x"2A", -- 0x00F8
    x"80",x"3E",x"FF",x"32",x"2B",x"80",x"AF",x"32", -- 0x0100
    x"2C",x"80",x"3E",x"0B",x"06",x"00",x"CD",x"0A", -- 0x0108
    x"05",x"3E",x"0C",x"06",x"20",x"CD",x"0A",x"05", -- 0x0110
    x"CD",x"EB",x"04",x"06",x"10",x"CD",x"86",x"04", -- 0x0118
    x"C9",x"3E",x"06",x"06",x"12",x"CD",x"0A",x"05", -- 0x0120
    x"3A",x"2C",x"80",x"FE",x"00",x"28",x"0C",x"FE", -- 0x0128
    x"01",x"28",x"16",x"21",x"2B",x"80",x"35",x"28", -- 0x0130
    x"2C",x"AF",x"C9",x"3E",x"0D",x"06",x"09",x"CD", -- 0x0138
    x"0A",x"05",x"3E",x"01",x"32",x"2C",x"80",x"18", -- 0x0140
    x"F0",x"21",x"29",x"80",x"35",x"20",x"EA",x"3E", -- 0x0148
    x"20",x"77",x"21",x"2A",x"80",x"35",x"20",x"07", -- 0x0150
    x"3E",x"02",x"32",x"2C",x"80",x"18",x"DA",x"AF", -- 0x0158
    x"32",x"2C",x"80",x"18",x"D4",x"3E",x"FF",x"C9", -- 0x0160
    x"3E",x"10",x"32",x"2E",x"80",x"21",x"F0",x"00", -- 0x0168
    x"CD",x"12",x"04",x"CD",x"58",x"04",x"06",x"0F", -- 0x0170
    x"CD",x"86",x"04",x"C9",x"21",x"2E",x"80",x"35", -- 0x0178
    x"20",x"0D",x"3E",x"10",x"77",x"CD",x"10",x"05", -- 0x0180
    x"3D",x"28",x"20",x"47",x"CD",x"86",x"04",x"CD", -- 0x0188
    x"35",x"04",x"B7",x"11",x"08",x"00",x"ED",x"52", -- 0x0190
    x"11",x"10",x"00",x"7C",x"BA",x"20",x"07",x"7D", -- 0x0198
    x"BB",x"20",x"03",x"21",x"F0",x"00",x"CD",x"12", -- 0x01A0
    x"04",x"AF",x"C9",x"3E",x"FF",x"C9",x"3E",x"08", -- 0x01A8
    x"32",x"30",x"80",x"3E",x"05",x"32",x"31",x"80", -- 0x01B0
    x"3E",x"0C",x"32",x"32",x"80",x"AF",x"32",x"33", -- 0x01B8
    x"80",x"21",x"50",x"00",x"CD",x"12",x"04",x"CD", -- 0x01C0
    x"58",x"04",x"06",x"00",x"CD",x"86",x"04",x"C9", -- 0x01C8
    x"3A",x"33",x"80",x"FE",x"00",x"28",x"18",x"FE", -- 0x01D0
    x"01",x"28",x"26",x"FE",x"02",x"28",x"27",x"FE", -- 0x01D8
    x"03",x"28",x"33",x"21",x"32",x"80",x"35",x"28", -- 0x01E0
    x"32",x"AF",x"32",x"33",x"80",x"AF",x"C9",x"CD", -- 0x01E8
    x"10",x"05",x"3C",x"FE",x"0F",x"20",x"04",x"21", -- 0x01F0
    x"33",x"80",x"34",x"47",x"CD",x"86",x"04",x"18", -- 0x01F8
    x"EC",x"CD",x"1E",x"0A",x"18",x"E7",x"CD",x"10", -- 0x0200
    x"05",x"3D",x"20",x"04",x"21",x"33",x"80",x"34", -- 0x0208
    x"47",x"CD",x"86",x"04",x"18",x"D7",x"CD",x"2B", -- 0x0210
    x"0A",x"18",x"D2",x"3E",x"FF",x"C9",x"21",x"30", -- 0x0218
    x"80",x"35",x"C0",x"3E",x"08",x"77",x"21",x"33", -- 0x0220
    x"80",x"34",x"C9",x"21",x"31",x"80",x"35",x"C0", -- 0x0228
    x"3E",x"05",x"77",x"21",x"33",x"80",x"34",x"C9", -- 0x0230
    x"3E",x"08",x"32",x"35",x"80",x"3E",x"01",x"32", -- 0x0238
    x"36",x"80",x"21",x"03",x"00",x"22",x"37",x"80", -- 0x0240
    x"AF",x"32",x"39",x"80",x"32",x"3A",x"80",x"21", -- 0x0248
    x"15",x"01",x"CD",x"12",x"04",x"CD",x"58",x"04", -- 0x0250
    x"06",x"0F",x"CD",x"86",x"04",x"C9",x"3A",x"39", -- 0x0258
    x"80",x"FE",x"01",x"28",x"14",x"FE",x"02",x"28", -- 0x0260
    x"24",x"3A",x"3A",x"80",x"FE",x"1C",x"28",x"3E", -- 0x0268
    x"E6",x"01",x"20",x"49",x"CD",x"E7",x"0A",x"AF", -- 0x0270
    x"C9",x"CD",x"10",x"05",x"C6",x"05",x"FE",x"0F", -- 0x0278
    x"20",x"05",x"21",x"39",x"80",x"36",x"00",x"47", -- 0x0280
    x"CD",x"86",x"04",x"18",x"EA",x"CD",x"10",x"05", -- 0x0288
    x"D6",x"01",x"20",x"05",x"21",x"39",x"80",x"36", -- 0x0290
    x"00",x"47",x"CD",x"86",x"04",x"3A",x"39",x"80", -- 0x0298
    x"FE",x"00",x"20",x"D3",x"3A",x"3A",x"80",x"FE", -- 0x02A0
    x"1C",x"20",x"CC",x"3E",x"FF",x"C9",x"CD",x"FB", -- 0x02A8
    x"0A",x"B7",x"20",x"02",x"18",x"C1",x"21",x"39", -- 0x02B0
    x"80",x"36",x"02",x"18",x"BA",x"CD",x"C2",x"0A", -- 0x02B8
    x"18",x"B5",x"CD",x"FB",x"0A",x"B7",x"C8",x"ED", -- 0x02C0
    x"5B",x"37",x"80",x"1A",x"32",x"36",x"80",x"13", -- 0x02C8
    x"1A",x"6F",x"13",x"1A",x"67",x"13",x"ED",x"53", -- 0x02D0
    x"37",x"80",x"CD",x"12",x"04",x"21",x"3A",x"80", -- 0x02D8
    x"34",x"21",x"39",x"80",x"36",x"01",x"C9",x"CD", -- 0x02E0
    x"FB",x"0A",x"B7",x"C8",x"3E",x"01",x"32",x"36", -- 0x02E8
    x"80",x"21",x"3A",x"80",x"34",x"21",x"39",x"80", -- 0x02F0
    x"36",x"02",x"C9",x"21",x"35",x"80",x"35",x"20", -- 0x02F8
    x"0C",x"3E",x"08",x"77",x"21",x"36",x"80",x"35", -- 0x0300
    x"20",x"03",x"3E",x"FF",x"C9",x"AF",x"C9",x"3E", -- 0x0308
    x"40",x"32",x"3C",x"80",x"3E",x"20",x"32",x"3D", -- 0x0310
    x"80",x"AF",x"32",x"3E",x"80",x"21",x"00",x"08", -- 0x0318
    x"CD",x"12",x"04",x"CD",x"58",x"04",x"06",x"0F", -- 0x0320
    x"CD",x"86",x"04",x"C9",x"3A",x"3E",x"80",x"FE", -- 0x0328
    x"00",x"28",x"20",x"FE",x"01",x"28",x"29",x"CD", -- 0x0330
    x"35",x"04",x"B7",x"11",x"20",x"00",x"ED",x"52", -- 0x0338
    x"11",x"00",x"02",x"7C",x"BA",x"20",x"07",x"7D", -- 0x0340
    x"BB",x"20",x"03",x"21",x"00",x"08",x"CD",x"12", -- 0x0348
    x"04",x"AF",x"C9",x"21",x"3C",x"80",x"35",x"20", -- 0x0350
    x"DE",x"3E",x"01",x"32",x"3E",x"80",x"18",x"D7", -- 0x0358
    x"21",x"3D",x"80",x"35",x"20",x"D1",x"3E",x"20", -- 0x0360
    x"77",x"CD",x"10",x"05",x"3D",x"28",x"06",x"47", -- 0x0368
    x"CD",x"86",x"04",x"18",x"C2",x"3E",x"FF",x"C9", -- 0x0370
    x"3E",x"05",x"32",x"40",x"80",x"21",x"50",x"00", -- 0x0378
    x"CD",x"12",x"04",x"CD",x"58",x"04",x"06",x"0F", -- 0x0380
    x"CD",x"86",x"04",x"C9",x"21",x"40",x"80",x"35", -- 0x0388
    x"20",x"0C",x"36",x"05",x"CD",x"10",x"05",x"3D", -- 0x0390
    x"28",x"06",x"47",x"CD",x"86",x"04",x"AF",x"C9", -- 0x0398
    x"3E",x"FF",x"C9",x"3E",x"04",x"32",x"42",x"80", -- 0x03A0
    x"3E",x"03",x"32",x"43",x"80",x"AF",x"32",x"44", -- 0x03A8
    x"80",x"CD",x"58",x"04",x"06",x"00",x"CD",x"86", -- 0x03B0
    x"04",x"C9",x"3A",x"44",x"80",x"FE",x"00",x"28", -- 0x03B8
    x"24",x"FE",x"01",x"28",x"31",x"CD",x"35",x"04", -- 0x03C0
    x"01",x"20",x"00",x"B7",x"09",x"CD",x"12",x"04", -- 0x03C8
    x"21",x"43",x"80",x"35",x"20",x"0D",x"36",x"03", -- 0x03D0
    x"CD",x"10",x"05",x"D6",x"03",x"28",x"23",x"47", -- 0x03D8
    x"CD",x"86",x"04",x"AF",x"C9",x"21",x"10",x"00", -- 0x03E0
    x"CD",x"12",x"04",x"06",x"0F",x"CD",x"86",x"04", -- 0x03E8
    x"21",x"44",x"80",x"34",x"18",x"ED",x"21",x"42", -- 0x03F0
    x"80",x"35",x"20",x"E7",x"21",x"44",x"80",x"34", -- 0x03F8
    x"18",x"E1",x"3E",x"FF",x"C9",x"3E",x"02",x"32", -- 0x0400
    x"46",x"80",x"3E",x"20",x"32",x"47",x"80",x"AF", -- 0x0408
    x"32",x"48",x"80",x"21",x"10",x"00",x"CD",x"12", -- 0x0410
    x"04",x"CD",x"58",x"04",x"06",x"00",x"CD",x"86", -- 0x0418
    x"04",x"C9",x"21",x"46",x"80",x"35",x"20",x"09", -- 0x0420
    x"36",x"02",x"CD",x"35",x"04",x"23",x"CD",x"12", -- 0x0428
    x"04",x"3A",x"48",x"80",x"FE",x"00",x"28",x"11", -- 0x0430
    x"FE",x"01",x"28",x"1F",x"21",x"47",x"80",x"35", -- 0x0438
    x"28",x"29",x"21",x"48",x"80",x"36",x"00",x"AF", -- 0x0440
    x"C9",x"CD",x"10",x"05",x"3C",x"FE",x"0F",x"20", -- 0x0448
    x"04",x"21",x"48",x"80",x"34",x"47",x"CD",x"86", -- 0x0450
    x"04",x"18",x"EC",x"CD",x"10",x"05",x"3D",x"20", -- 0x0458
    x"04",x"21",x"48",x"80",x"34",x"47",x"CD",x"86", -- 0x0460
    x"04",x"18",x"DC",x"3E",x"FF",x"C9",x"3E",x"03", -- 0x0468
    x"32",x"4A",x"80",x"21",x"00",x"04",x"22",x"4C", -- 0x0470
    x"80",x"AF",x"32",x"4B",x"80",x"21",x"00",x"02", -- 0x0478
    x"CD",x"12",x"04",x"CD",x"58",x"04",x"06",x"0A", -- 0x0480
    x"CD",x"86",x"04",x"C9",x"21",x"4A",x"80",x"35", -- 0x0488
    x"20",x"2E",x"36",x"03",x"CD",x"35",x"04",x"11", -- 0x0490
    x"20",x"00",x"19",x"ED",x"5B",x"4C",x"80",x"7C", -- 0x0498
    x"BA",x"20",x"18",x"7D",x"BB",x"20",x"14",x"3A", -- 0x04A0
    x"4B",x"80",x"B7",x"20",x"15",x"21",x"00",x"08", -- 0x04A8
    x"22",x"4C",x"80",x"3E",x"FF",x"32",x"4B",x"80", -- 0x04B0
    x"21",x"00",x"02",x"CD",x"12",x"04",x"AF",x"C9", -- 0x04B8
    x"AF",x"C9",x"21",x"00",x"04",x"22",x"4C",x"80", -- 0x04C0
    x"AF",x"32",x"4B",x"80",x"18",x"EA",x"3E",x"10", -- 0x04C8
    x"32",x"4F",x"80",x"AF",x"32",x"50",x"80",x"32", -- 0x04D0
    x"51",x"80",x"CD",x"58",x"04",x"06",x"00",x"CD", -- 0x04D8
    x"86",x"04",x"C9",x"3A",x"51",x"80",x"FE",x"00", -- 0x04E0
    x"CA",x"51",x"0D",x"FE",x"01",x"CA",x"5E",x"0D", -- 0x04E8
    x"FE",x"02",x"CA",x"69",x"0D",x"FE",x"03",x"CA", -- 0x04F0
    x"6F",x"0D",x"FE",x"04",x"CA",x"7A",x"0D",x"FE", -- 0x04F8
    x"05",x"CA",x"80",x"0D",x"FE",x"06",x"CA",x"8D", -- 0x0500
    x"0D",x"FE",x"07",x"CA",x"98",x"0D",x"FE",x"08", -- 0x0508
    x"CA",x"9E",x"0D",x"FE",x"09",x"CA",x"A9",x"0D", -- 0x0510
    x"FE",x"0A",x"CA",x"AF",x"0D",x"FE",x"0B",x"CA", -- 0x0518
    x"BC",x"0D",x"FE",x"0C",x"CA",x"C7",x"0D",x"FE", -- 0x0520
    x"0D",x"CA",x"CD",x"0D",x"FE",x"0E",x"CA",x"D8", -- 0x0528
    x"0D",x"FE",x"0F",x"CA",x"DE",x"0D",x"FE",x"10", -- 0x0530
    x"CA",x"EB",x"0D",x"FE",x"11",x"CA",x"F6",x"0D", -- 0x0538
    x"FE",x"12",x"CA",x"FC",x"0D",x"FE",x"13",x"CA", -- 0x0540
    x"07",x"0E",x"21",x"51",x"80",x"36",x"00",x"AF", -- 0x0548
    x"C9",x"21",x"E7",x"0B",x"CD",x"12",x"04",x"21", -- 0x0550
    x"51",x"80",x"34",x"C3",x"4F",x"0D",x"CD",x"0D", -- 0x0558
    x"0E",x"21",x"50",x"80",x"36",x"05",x"C3",x"4F", -- 0x0560
    x"0D",x"CD",x"21",x"0E",x"C3",x"4F",x"0D",x"CD", -- 0x0568
    x"17",x"0E",x"21",x"50",x"80",x"36",x"01",x"C3", -- 0x0570
    x"4F",x"0D",x"CD",x"21",x"0E",x"C3",x"4F",x"0D", -- 0x0578
    x"21",x"00",x"0A",x"CD",x"12",x"04",x"21",x"51", -- 0x0580
    x"80",x"34",x"C3",x"4F",x"0D",x"CD",x"0D",x"0E", -- 0x0588
    x"21",x"50",x"80",x"36",x"05",x"C3",x"4F",x"0D", -- 0x0590
    x"CD",x"21",x"0E",x"C3",x"4F",x"0D",x"CD",x"17", -- 0x0598
    x"0E",x"21",x"50",x"80",x"36",x"01",x"C3",x"4F", -- 0x05A0
    x"0D",x"CD",x"21",x"0E",x"C3",x"4F",x"0D",x"21", -- 0x05A8
    x"99",x"0A",x"CD",x"12",x"04",x"21",x"51",x"80", -- 0x05B0
    x"34",x"C3",x"4F",x"0D",x"CD",x"0D",x"0E",x"21", -- 0x05B8
    x"50",x"80",x"36",x"05",x"C3",x"4F",x"0D",x"CD", -- 0x05C0
    x"21",x"0E",x"C3",x"4F",x"0D",x"CD",x"17",x"0E", -- 0x05C8
    x"21",x"50",x"80",x"36",x"01",x"C3",x"4F",x"0D", -- 0x05D0
    x"CD",x"21",x"0E",x"C3",x"4F",x"0D",x"21",x"3B", -- 0x05D8
    x"0B",x"CD",x"12",x"04",x"21",x"51",x"80",x"34", -- 0x05E0
    x"C3",x"4F",x"0D",x"CD",x"0D",x"0E",x"21",x"50", -- 0x05E8
    x"80",x"36",x"05",x"C3",x"4F",x"0D",x"CD",x"21", -- 0x05F0
    x"0E",x"C3",x"4F",x"0D",x"CD",x"17",x"0E",x"21", -- 0x05F8
    x"50",x"80",x"36",x"01",x"C3",x"4F",x"0D",x"CD", -- 0x0600
    x"21",x"0E",x"C3",x"4F",x"0D",x"06",x"0A",x"CD", -- 0x0608
    x"86",x"04",x"21",x"51",x"80",x"34",x"C9",x"06", -- 0x0610
    x"00",x"CD",x"86",x"04",x"21",x"51",x"80",x"34", -- 0x0618
    x"C9",x"21",x"4F",x"80",x"35",x"C0",x"36",x"10", -- 0x0620
    x"21",x"50",x"80",x"35",x"C0",x"21",x"51",x"80", -- 0x0628
    x"34",x"C9",x"21",x"40",x"01",x"22",x"53",x"80", -- 0x0630
    x"11",x"01",x"00",x"ED",x"53",x"55",x"80",x"3E", -- 0x0638
    x"03",x"32",x"57",x"80",x"3E",x"20",x"32",x"58", -- 0x0640
    x"80",x"3E",x"40",x"32",x"59",x"80",x"32",x"5A", -- 0x0648
    x"80",x"AF",x"32",x"5B",x"80",x"CD",x"58",x"04", -- 0x0650
    x"06",x"00",x"CD",x"86",x"04",x"C9",x"3A",x"5B", -- 0x0658
    x"80",x"FE",x"00",x"28",x"29",x"FE",x"01",x"28", -- 0x0660
    x"31",x"FE",x"02",x"28",x"40",x"FE",x"03",x"28", -- 0x0668
    x"4F",x"FE",x"04",x"28",x"70",x"21",x"59",x"80", -- 0x0670
    x"35",x"20",x"11",x"3A",x"5A",x"80",x"32",x"59", -- 0x0678
    x"80",x"11",x"01",x"00",x"ED",x"53",x"55",x"80", -- 0x0680
    x"AF",x"32",x"5B",x"80",x"AF",x"C9",x"2A",x"53", -- 0x0688
    x"80",x"CD",x"12",x"04",x"21",x"5B",x"80",x"34", -- 0x0690
    x"18",x"F2",x"CD",x"10",x"05",x"C6",x"02",x"FE", -- 0x0698
    x"08",x"20",x"04",x"21",x"5B",x"80",x"34",x"47", -- 0x06A0
    x"CD",x"86",x"04",x"18",x"DF",x"CD",x"35",x"04", -- 0x06A8
    x"B7",x"ED",x"5B",x"55",x"80",x"ED",x"52",x"CD", -- 0x06B0
    x"12",x"04",x"21",x"5B",x"80",x"34",x"18",x"CC", -- 0x06B8
    x"21",x"57",x"80",x"35",x"20",x"0B",x"36",x"03", -- 0x06C0
    x"ED",x"5B",x"55",x"80",x"13",x"ED",x"53",x"55", -- 0x06C8
    x"80",x"21",x"58",x"80",x"35",x"20",x"08",x"36", -- 0x06D0
    x"20",x"21",x"5B",x"80",x"34",x"18",x"AD",x"21", -- 0x06D8
    x"5B",x"80",x"35",x"18",x"A7",x"CD",x"10",x"05", -- 0x06E0
    x"3D",x"20",x"04",x"21",x"5B",x"80",x"34",x"47", -- 0x06E8
    x"CD",x"86",x"04",x"18",x"97",x"21",x"20",x"01", -- 0x06F0
    x"22",x"53",x"80",x"11",x"01",x"00",x"ED",x"53", -- 0x06F8
    x"55",x"80",x"3E",x"03",x"32",x"57",x"80",x"3E", -- 0x0700
    x"20",x"32",x"58",x"80",x"3E",x"30",x"32",x"59", -- 0x0708
    x"80",x"32",x"5A",x"80",x"AF",x"32",x"5B",x"80", -- 0x0710
    x"CD",x"58",x"04",x"06",x"00",x"CD",x"86",x"04", -- 0x0718
    x"C9",x"C3",x"5E",x"0E",x"21",x"00",x"01",x"22", -- 0x0720
    x"53",x"80",x"11",x"01",x"00",x"ED",x"53",x"55", -- 0x0728
    x"80",x"3E",x"03",x"32",x"57",x"80",x"3E",x"20", -- 0x0730
    x"32",x"58",x"80",x"3E",x"20",x"32",x"59",x"80", -- 0x0738
    x"32",x"5A",x"80",x"AF",x"32",x"5B",x"80",x"CD", -- 0x0740
    x"58",x"04",x"06",x"00",x"CD",x"86",x"04",x"C9", -- 0x0748
    x"C3",x"5E",x"0E",x"3E",x"10",x"32",x"5D",x"80", -- 0x0750
    x"3E",x"03",x"32",x"5E",x"80",x"AF",x"32",x"5F", -- 0x0758
    x"80",x"21",x"E3",x"0F",x"22",x"60",x"80",x"21", -- 0x0760
    x"15",x"01",x"CD",x"12",x"04",x"CD",x"58",x"04", -- 0x0768
    x"06",x"0F",x"CD",x"86",x"04",x"C9",x"3A",x"5F", -- 0x0770
    x"80",x"FE",x"0A",x"20",x"08",x"CD",x"AA",x"0F", -- 0x0778
    x"B7",x"20",x"10",x"AF",x"C9",x"E6",x"01",x"28", -- 0x0780
    x"05",x"CD",x"BE",x"0F",x"18",x"F5",x"CD",x"96", -- 0x0788
    x"0F",x"18",x"F0",x"3E",x"FF",x"C9",x"CD",x"AA", -- 0x0790
    x"0F",x"B7",x"C8",x"3E",x"01",x"32",x"5E",x"80", -- 0x0798
    x"21",x"5F",x"80",x"34",x"06",x"00",x"CD",x"86", -- 0x07A0
    x"04",x"C9",x"21",x"5D",x"80",x"35",x"20",x"0C", -- 0x07A8
    x"3E",x"10",x"77",x"21",x"5E",x"80",x"35",x"20", -- 0x07B0
    x"03",x"3E",x"FF",x"C9",x"AF",x"C9",x"CD",x"AA", -- 0x07B8
    x"0F",x"B7",x"C8",x"ED",x"5B",x"60",x"80",x"1A", -- 0x07C0
    x"32",x"5E",x"80",x"13",x"1A",x"6F",x"13",x"1A", -- 0x07C8
    x"67",x"13",x"ED",x"53",x"60",x"80",x"CD",x"12", -- 0x07D0
    x"04",x"21",x"5F",x"80",x"34",x"06",x"0F",x"CD", -- 0x07D8
    x"86",x"04",x"C9",x"01",x"15",x"01",x"08",x"D0", -- 0x07E0
    x"00",x"03",x"15",x"01",x"01",x"D0",x"00",x"08", -- 0x07E8
    x"A5",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF"  -- 0x07F8
  );

begin

  p_rom : process
  begin
    wait until rising_edge(CLK);
     DATA <= ROM(to_integer(unsigned(ADDR)));
  end process;
end RTL;
