library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity popeye_sp_bits_2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of popeye_sp_bits_2 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"18",X"00",X"18",X"00",X"8E",X"00",X"9C",X"00",X"F0",X"00",X"60",X"00",X"00",X"00",X"00",
		X"CC",X"00",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"81",X"00",X"83",X"00",X"07",X"00",X"0F",X"00",X"07",X"00",X"03",
		X"00",X"00",X"00",X"C0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"0F",X"1D",X"18",X"1C",
		X"0E",X"0E",X"06",X"06",X"0C",X"8C",X"8C",X"8C",X"98",X"98",X"D8",X"F8",X"F0",X"70",X"30",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"3F",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C1",X"C1",X"C3",X"C3",X"C3",X"C3",
		X"46",X"46",X"24",X"38",X"F8",X"F0",X"FC",X"DE",X"8F",X"0F",X"CF",X"EF",X"FF",X"7F",X"3F",X"9F",
		X"DF",X"F7",X"EF",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"FC",X"F8",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",X"E0",X"E0",X"C0",X"C0",X"C0",X"E0",X"E0",X"E0",
		X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"80",X"C0",X"C0",X"40",X"00",X"00",X"80",X"80",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"EE",X"F8",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"07",X"03",X"07",X"07",
		X"07",X"07",X"07",X"03",X"00",X"37",X"57",X"7F",X"1F",X"0C",X"00",X"73",X"7D",X"3F",X"1F",X"01",
		X"04",X"44",X"63",X"63",X"E7",X"E6",X"C0",X"C3",X"FF",X"FE",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0E",X"07",X"03",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"38",X"3C",X"1C",X"0E",X"07",X"03",
		X"00",X"00",X"20",X"78",X"7F",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"04",X"08",X"09",X"1A",X"E6",X"20",X"00",
		X"00",X"00",X"01",X"6E",X"3C",X"00",X"00",X"11",X"E3",X"C7",X"0E",X"04",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"40",X"20",X"00",X"07",X"3C",X"FE",X"FE",X"C8",X"00",X"04",X"18",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"84",
		X"86",X"C3",X"E0",X"00",X"00",X"00",X"22",X"17",X"9F",X"07",X"03",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"03",X"23",X"61",X"70",X"30",X"18",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"1C",X"FE",X"FE",X"FE",X"FE",X"FC",X"FC",X"FC",X"FC",X"F8",X"F6",X"EF",X"DF",
		X"DF",X"DF",X"FF",X"FF",X"FE",X"FC",X"F8",X"F8",X"F0",X"F0",X"E0",X"E0",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"80",X"E0",X"A0",X"E0",X"C0",X"C0",X"C0",X"C0",X"80",X"00",X"40",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"03",X"0F",X"3F",X"FC",X"F0",X"F0",X"E0",X"60",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"80",X"3C",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"E3",X"E1",X"E1",X"E1",X"F8",X"78",X"F8",X"FC",X"FC",X"FE",X"3F",X"0F",X"0F",X"03",X"00",
		X"00",X"01",X"06",X"8F",X"4F",X"0F",X"0F",X"01",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",
		X"DF",X"DF",X"FF",X"FF",X"FE",X"FC",X"F8",X"F8",X"F0",X"F0",X"E0",X"E0",X"C0",X"C0",X"80",X"00",
		X"00",X"80",X"60",X"E0",X"E0",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"F1",X"E1",X"E1",X"E1",X"F1",X"70",X"78",X"BC",X"BE",X"DF",X"FF",X"FF",X"8F",X"81",
		X"00",X"01",X"03",X"03",X"07",X"86",X"00",X"00",X"80",X"01",X"1E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"E0",X"E0",X"E0",
		X"F0",X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F0",X"F0",
		X"F0",X"E0",X"E0",X"E0",X"C0",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"F0",X"FE",X"FF",X"FF",X"FF",X"3F",X"1F",X"CF",X"8F",X"0F",X"0F",X"1F",X"FF",X"FF",X"FF",
		X"1F",X"0F",X"87",X"C7",X"C7",X"C7",X"87",X"8F",X"8F",X"1F",X"1F",X"3F",X"7F",X"FF",X"7F",X"7F",
		X"3F",X"1F",X"1F",X"1F",X"1F",X"1F",X"3F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"E0",
		X"03",X"06",X"04",X"01",X"07",X"0F",X"1F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FE",X"FC",X"FC",X"FC",X"FC",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"FE",X"FF",X"7F",X"3F",X"0F",X"03",X"01",X"00",X"00",
		X"00",X"00",X"00",X"10",X"00",X"04",X"00",X"00",X"02",X"00",X"00",X"02",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"50",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"08",X"08",X"00",X"00",X"10",X"20",X"40",X"40",X"80",X"80",X"80",X"80",X"00",X"00",
		X"00",X"00",X"0F",X"0F",X"03",X"03",X"03",X"0F",X"0F",X"03",X"03",X"03",X"0F",X"0F",X"00",X"00",
		X"F8",X"FC",X"FE",X"FE",X"FE",X"FE",X"FC",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"04",X"04",X"04",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"C0",X"E0",X"F0",X"F8",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"3E",X"1C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"FC",X"00",X"00",X"00",X"00",X"00",X"60",X"60",X"60",X"60",X"60",X"60",X"20",X"00",X"00",
		X"F8",X"FC",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"00",
		X"78",X"7C",X"60",X"60",X"60",X"E0",X"E0",X"00",X"00",X"00",X"60",X"60",X"60",X"20",X"00",X"00",
		X"78",X"7C",X"7E",X"7E",X"7E",X"FE",X"FE",X"FE",X"FE",X"FE",X"7E",X"7E",X"3E",X"FE",X"FE",X"00",
		X"00",X"00",X"30",X"30",X"30",X"30",X"30",X"F0",X"F0",X"30",X"30",X"30",X"F0",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"F0",X"F0",X"C0",X"C0",X"F8",X"FC",X"FC",X"FE",X"FE",X"FE",X"FE",X"FC",X"3C",X"18",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"1F",X"0F",X"0F",X"07",X"07",X"87",X"F7",X"FE",X"7C",X"00",
		X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"E0",X"F8",X"FC",X"FE",X"FE",X"FF",X"FF",X"7F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3E",X"3E",X"3E",X"7C",X"FC",X"FC",X"F8",X"F0",X"EC",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",
		X"7E",X"7E",X"7E",X"7E",X"7C",X"7C",X"7C",X"78",X"70",X"60",X"F0",X"F0",X"E0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"83",X"DF",X"BF",X"FF",X"FF",X"FF",X"FF",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",
		X"3C",X"3C",X"0C",X"0E",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"30",X"30",X"32",X"32",X"32",X"32",X"32",X"32",X"30",X"30",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",
		X"00",X"03",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"33",X"33",X"33",X"33",X"03",X"03",
		X"33",X"33",X"33",X"33",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3C",X"3C",X"3F",X"3F",X"0C",X"CC",X"CF",X"CF",X"CC",X"CC",X"FF",X"FF",X"FF",X"FE",X"F0",X"00",
		X"FF",X"E7",X"3D",X"0F",X"0F",X"C7",X"FB",X"FF",X"FF",X"FF",X"DF",X"8F",X"07",X"03",X"01",X"00",
		X"00",X"00",X"00",X"00",X"21",X"73",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"67",X"67",X"FF",X"FF",X"67",X"67",X"67",X"67",X"67",X"67",X"FF",X"FF",X"FF",X"1F",X"0F",X"00",
		X"FF",X"E7",X"3D",X"0F",X"0F",X"C7",X"FB",X"FF",X"FF",X"FF",X"83",X"01",X"02",X"02",X"02",X"04",
		X"01",X"83",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"00",X"E0",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1E",X"00",X"3F",X"00",X"1E",
		X"00",X"D0",X"D0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F6",X"DF",X"DF",X"FC",X"FE",X"FE",X"FC",X"D8",
		X"00",X"80",X"C0",X"E0",X"F0",X"60",X"44",X"0C",X"7C",X"98",X"40",X"B0",X"FC",X"0E",X"07",X"03",
		X"00",X"68",X"64",X"32",X"20",X"00",X"18",X"18",X"40",X"E0",X"C0",X"F0",X"A0",X"C0",X"80",X"00",
		X"00",X"80",X"C0",X"E0",X"F0",X"60",X"C4",X"8C",X"1C",X"38",X"30",X"A0",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"06",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"42",X"4A",X"29",X"25",X"04",X"04",X"22",X"E2",X"82",X"10",X"00",X"10",X"98",X"90",X"C8",
		X"C8",X"90",X"90",X"00",X"10",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"20",X"A0",X"A0",X"A0",X"20",X"40",X"40",X"40",X"80",X"80",X"90",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"06",X"0C",X"38",X"EC",X"86",X"03",X"07",X"05",X"84",X"81",X"C4",X"C0",X"81",X"B0",X"0C",
		X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"04",
		X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"06",X"0C",X"38",X"EC",X"86",X"03",X"03",X"05",X"84",X"82",X"C0",X"C0",X"80",X"82",X"41",
		X"20",X"11",X"40",X"08",X"80",X"04",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"80",X"80",X"F3",X"DF",X"BE",X"F0",X"B0",X"60",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"90",X"90",X"10",X"20",X"20",X"20",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"48",X"50",X"90",X"20",X"20",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0D",X"17",X"07",X"26",X"2C",X"38",X"10",X"80",X"88",X"8C",X"9E",X"9E",X"9F",X"9F",X"9F",
		X"9F",X"9F",X"BF",X"BE",X"BC",X"B0",X"F0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"F8",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"7C",X"EE",X"C6",X"0C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"1F",X"3F",X"7F",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"0F",X"3F",X"F9",X"E3",X"C3",X"C3",X"C3",
		X"46",X"46",X"24",X"38",X"F8",X"F0",X"BC",X"9E",X"0F",X"CF",X"EF",X"FF",X"FF",X"7F",X"3F",X"9F",
		X"04",X"07",X"07",X"07",X"03",X"00",X"00",X"00",X"79",X"00",X"04",X"08",X"10",X"30",X"60",X"60",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"3C",X"18",X"18",X"3C",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D8",X"5C",X"4C",X"24",X"20",X"C0",X"F0",X"E0",
		X"C4",X"DE",X"7E",X"3E",X"26",X"70",X"F8",X"BC",X"3C",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"F0",X"FC",X"FE",X"FE",X"3F",X"1F",X"1F",X"3F",X"FE",X"FE",X"FC",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"7E",X"F8",X"C0",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"F8",X"FC",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"F8",
		X"F0",X"1C",X"06",X"7E",X"F8",X"C0",X"00",X"02",X"06",X"08",X"70",X"80",X"02",X"02",X"04",X"08",
		X"70",X"80",X"02",X"02",X"06",X"1C",X"F8",X"E8",X"A8",X"28",X"20",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F4",X"8C",X"F8",X"F0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"3F",X"7E",X"FD",X"FF",X"FF",X"FF",X"FF",
		X"F0",X"F0",X"E0",X"E0",X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",X"FC",X"FC",X"FC",X"FC",X"FC",X"FE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FD",X"F2",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FD",
		X"00",X"00",X"30",X"80",X"E0",X"F0",X"F0",X"F8",X"F8",X"78",X"BC",X"BC",X"BC",X"BC",X"DC",X"C0",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F7",X"FB",X"FD",X"FD",X"FD",X"FD",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FD",
		X"FD",X"FD",X"FB",X"F7",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"F8",X"F3",
		X"00",X"00",X"00",X"00",X"00",X"00",X"39",X"3B",X"B7",X"B7",X"76",X"77",X"7F",X"7F",X"FF",X"FF",
		X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"1F",X"07",X"01",X"01",X"01",X"01",
		X"FC",X"FE",X"FC",X"FB",X"CF",X"9F",X"BF",X"3B",X"87",X"00",X"18",X"34",X"0A",X"85",X"C3",X"89",
		X"FC",X"BC",X"5C",X"15",X"32",X"F7",X"E7",X"06",X"05",X"1F",X"FF",X"FF",X"7F",X"3C",X"00",X"00",
		X"F0",X"F0",X"F8",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"78",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"3F",X"7F",X"FF",X"FF",X"FE",X"FF",X"FF",X"F0",X"CF",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"04",X"00",X"00",X"E0",X"F0",X"F8",X"FC",X"7E",X"7F",X"7F",X"7F",X"BF",X"BE",X"BC",X"80",
		X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"F0",
		X"98",X"CC",X"EC",X"F6",X"FA",X"FD",X"7E",X"BE",X"DF",X"DF",X"DF",X"FF",X"FF",X"FB",X"FD",X"FD",
		X"FE",X"FE",X"FE",X"FE",X"FC",X"F8",X"C0",X"80",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"E0",
		X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",X"F0",X"F0",X"E0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"C0",X"F0",X"1C",X"E7",X"F9",X"FE",X"FF",X"FF",
		X"1F",X"CF",X"E7",X"EF",X"FD",X"FE",X"FF",X"7F",X"FF",X"DF",X"EF",X"F7",X"FB",X"FD",X"FE",X"FE",
		X"FF",X"FF",X"BF",X"BF",X"5F",X"5F",X"DF",X"BF",X"7E",X"7C",X"F2",X"F3",X"EB",X"D7",X"F7",X"CF",
		X"BF",X"FF",X"FF",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"00",X"00",X"00",
		X"00",X"04",X"04",X"04",X"04",X"84",X"70",X"00",X"FF",X"FF",X"00",X"7F",X"FF",X"FF",X"FF",X"9F",
		X"7C",X"FF",X"FF",X"FF",X"FF",X"FF",X"E0",X"DE",X"FF",X"FF",X"FF",X"7F",X"3F",X"FF",X"02",X"FE",
		X"FD",X"FD",X"FD",X"FD",X"FC",X"BC",X"7C",X"7D",X"3F",X"AF",X"9E",X"9E",X"9D",X"1B",X"0F",X"0F",
		X"07",X"01",X"00",X"00",X"30",X"39",X"3F",X"1F",X"FF",X"FF",X"3F",X"FF",X"FF",X"EE",X"9C",X"0C",
		X"98",X"B8",X"B0",X"F0",X"FE",X"FE",X"FC",X"F8",X"F0",X"F8",X"F8",X"F9",X"FB",X"FB",X"F9",X"F9",
		X"F8",X"F3",X"F7",X"FB",X"FB",X"FB",X"FB",X"F7",X"EE",X"DE",X"BC",X"FC",X"FC",X"FF",X"FF",X"FE",
		X"FF",X"FF",X"7F",X"B6",X"01",X"39",X"4C",X"46",X"63",X"11",X"08",X"04",X"63",X"F3",X"70",X"A0",
		X"7D",X"5A",X"36",X"EC",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"01",X"01",X"00",X"00",
		X"FF",X"3F",X"CF",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C7",
		X"E7",X"FF",X"FF",X"FF",X"FF",X"DB",X"E0",X"E0",X"CE",X"0A",X"1A",X"16",X"34",X"EC",X"99",X"73",
		X"4B",X"1F",X"18",X"01",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"1F",X"3F",X"7E",X"7D",X"FB",X"F7",X"EF",X"EF",X"FF",X"FF",X"FE",X"FE",
		X"EF",X"E5",X"CF",X"6F",X"0E",X"0F",X"06",X"05",X"07",X"07",X"07",X"07",X"03",X"01",X"03",X"03",
		X"0B",X"0D",X"1D",X"3E",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"F8",X"F0",
		X"E0",X"E0",X"F0",X"F0",X"78",X"38",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",
		X"00",X"06",X"04",X"02",X"0F",X"BF",X"BF",X"BF",X"7F",X"7F",X"BF",X"DF",X"FF",X"FF",X"C0",X"7F",
		X"00",X"00",X"3E",X"E0",X"00",X"00",X"06",X"7F",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FB",X"EF",X"DE",X"38",X"3B",X"3B",X"3B",X"3B",X"19",X"1E",X"1E",X"1C",X"0D",X"0D",X"0D",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0D",X"03",X"83",X"45",X"4E",X"4D",X"CF",X"8E",X"8F",X"2D",X"7A",X"65",X"00",X"00",X"00",X"00",
		X"80",X"80",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"C0",X"60",X"20",X"20",X"00",X"00",
		X"80",X"40",X"20",X"20",X"00",X"00",X"80",X"60",X"20",X"00",X"00",X"80",X"60",X"60",X"C0",X"00",
		X"FF",X"FF",X"FF",X"80",X"3F",X"FF",X"FF",X"FF",X"FF",X"F0",X"80",X"00",X"00",X"00",X"1F",X"E0",
		X"00",X"00",X"00",X"00",X"1F",X"E0",X"00",X"00",X"00",X"00",X"3F",X"FF",X"E0",X"00",X"80",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",X"F0",X"F0",X"F0",X"80",X"C0",X"E0",X"F0",X"F8",X"F8",
		X"C0",X"40",X"80",X"C0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"E0",X"C0",X"C0",X"C0",X"C0",
		X"80",X"80",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F1",X"CF",X"BF",X"FF",X"FF",X"FF",X"FF",X"E0",
		X"F7",X"EF",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"FF",
		X"FF",X"FF",X"FF",X"7F",X"DF",X"EF",X"F6",X"F8",X"FE",X"FF",X"FF",X"FF",X"FD",X"FE",X"FC",X"F0",
		X"F8",X"F0",X"F8",X"48",X"09",X"03",X"0E",X"0D",X"01",X"03",X"03",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"08",X"0C",X"00",X"00",X"00",X"01",X"01",X"03",X"03",X"03",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"01",X"03",X"06",X"07",X"07",X"07",X"03",X"03",X"01",X"60",X"66",X"67",
		X"67",X"77",X"BE",X"FF",X"FF",X"1F",X"0F",X"07",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7C",X"FE",X"FE",
		X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"FE",X"FE",X"FE",X"FE",X"FC",X"FC",X"FC",X"F8",X"F8",X"F0",
		X"F0",X"E0",X"E0",X"E0",X"C0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FB",X"FD",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F3",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"CF",X"D7",X"DB",X"9D",X"1E",X"9E",X"FF",X"FF",X"FF",X"FF",X"DF",X"BF",X"1B",X"07",
		X"06",X"06",X"0E",X"3E",X"FC",X"FA",X"FB",X"FB",X"FB",X"FD",X"FD",X"FE",X"FE",X"FF",X"FE",X"FE",
		X"FC",X"FC",X"F8",X"F8",X"F0",X"F0",X"F8",X"B8",X"7C",X"7C",X"7C",X"BC",X"C8",X"B0",X"70",X"E0",
		X"00",X"80",X"C0",X"80",X"C0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"C0",X"F0",X"F0",X"76",
		X"B0",X"D0",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",
		X"F8",X"F8",X"F8",X"F0",X"F0",X"F0",X"E0",X"E0",X"C0",X"80",X"80",X"80",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"F8",X"FF",X"FF",X"FF",X"18",X"E7",X"DE",X"3D",X"FB",X"FF",
		X"7F",X"BF",X"DF",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FE",X"FE",X"7F",X"77",X"7B",X"7D",
		X"7E",X"7E",X"7D",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"E0",X"E1",X"80",X"38",X"F8",X"F0",X"C0",X"80",X"C0",X"E0",X"F0",X"F0",X"F8",X"FC",X"FE",
		X"E9",X"E7",X"FF",X"DF",X"BF",X"BF",X"7F",X"7F",X"7F",X"BF",X"B7",X"8F",X"DF",X"FF",X"FF",X"FF",
		X"FF",X"7F",X"AD",X"83",X"00",X"7F",X"7A",X"0E",X"C2",X"E1",X"C4",X"7E",X"5E",X"AE",X"8A",X"99",
		X"FB",X"73",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"F0",X"F8",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"7C",X"F8",
		X"F8",X"F8",X"F8",X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",X"D8",X"D0",X"D0",X"E0",X"C0",X"80",X"00",
		X"60",X"38",X"1C",X"8C",X"CE",X"E6",X"F0",X"F8",X"30",X"DC",X"EE",X"F7",X"FF",X"FF",X"FF",X"80",
		X"FC",X"FE",X"FE",X"1F",X"EE",X"F4",X"F8",X"0C",X"F6",X"F7",X"FB",X"FB",X"F9",X"FA",X"FA",X"F6",
		X"F4",X"FD",X"FD",X"FD",X"FB",X"FB",X"FF",X"FF",X"FF",X"FF",X"CF",X"77",X"EB",X"1D",X"8D",X"8B",
		X"C7",X"45",X"42",X"C4",X"04",X"D8",X"9C",X"CC",X"E0",X"F0",X"E0",X"E0",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"1C",X"3C",X"3C",X"7D",X"7B",X"F7",X"FF",X"FF",
		X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"7F",X"7B",X"7D",X"3E",X"3F",X"1F",X"1F",X"1F",X"03",X"03",X"03",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"C0",X"C0",
		X"00",X"04",X"06",X"00",X"01",X"03",X"87",X"C7",X"E7",X"CF",X"FF",X"FF",X"FF",X"FF",X"80",X"9F",
		X"00",X"40",X"60",X"07",X"07",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"80",X"9F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"F0",X"F0",X"F8",X"F8",X"FC",X"FC",X"FE",X"FF",
		X"FF",X"FF",X"FF",X"FE",X"FE",X"FC",X"F8",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"60",X"01",X"03",X"0F",X"1F",X"07",X"00",X"00",X"C1",X"FF",X"FF",X"FF",X"80",X"9F",
		X"FB",X"FD",X"FE",X"FF",X"FF",X"EF",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C7",X"C2",X"86",X"26",X"74",X"F6",X"D6",X"E6",X"E0",X"B0",X"30",X"70",X"A0",X"00",X"00",X"00",
		X"0E",X"FE",X"FE",X"FE",X"FE",X"FE",X"3F",X"DF",X"FF",X"7F",X"3F",X"CE",X"E0",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",
		X"00",X"00",X"00",X"FC",X"F8",X"F0",X"F3",X"E7",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"80",X"9F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"80",X"C0",X"C0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"E0",X"E0",
		X"E0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"80",X"9F",
		X"FB",X"FD",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"EF",X"EF",X"D7",X"DB",X"DD",X"DE",X"1F",X"9F",X"FF",X"FF",X"FF",X"FF",X"DF",X"BF",X"1B",X"07",
		X"E3",X"C0",X"82",X"26",X"74",X"F6",X"D6",X"E6",X"60",X"30",X"70",X"F0",X"A0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"81",X"C1",X"01",X"01",X"01",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"1F",X"1D",X"1B",X"1B",X"1B",X"3B",X"3C",X"1F",X"1F",X"0C",X"0D",X"0D",X"05",X"06",
		X"7A",X"CE",X"B4",X"F2",X"E8",X"DA",X"77",X"6F",X"3D",X"1D",X"02",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"20",X"20",X"10",X"18",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"E0",X"F0",X"F0",
		X"F0",X"F8",X"FA",X"FA",X"FA",X"F6",X"77",X"77",X"76",X"7E",X"7E",X"7C",X"3C",X"38",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"04",X"F0",X"FE",X"FF",X"FF",X"1F",X"EF",X"77",X"FB",
		X"FB",X"FD",X"FD",X"FE",X"FE",X"FE",X"FF",X"FD",X"FC",X"78",X"38",X"30",X"20",X"40",X"D0",X"D8",
		X"D8",X"3C",X"FE",X"CF",X"3F",X"7F",X"FF",X"FF",X"FE",X"FE",X"FC",X"F8",X"E0",X"C0",X"C0",X"80",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"07",X"00",X"03",X"03",X"03",X"01",X"00",X"00",X"00",X"00",
		X"01",X"03",X"07",X"0F",X"31",X"F1",X"F9",X"FC",X"00",X"00",X"F9",X"F1",X"F3",X"F3",X"C6",X"C7",
		X"C7",X"C0",X"E0",X"E0",X"E0",X"E0",X"DC",X"1F",X"0F",X"07",X"3F",X"7F",X"67",X"0F",X"1D",X"19",
		X"18",X"B8",X"F6",X"FE",X"FC",X"F8",X"FE",X"FF",X"FF",X"38",X"98",X"58",X"70",X"70",X"70",X"E0",
		X"E0",X"E0",X"F8",X"7C",X"78",X"7B",X"37",X"0F",X"00",X"00",X"00",X"3C",X"66",X"67",X"6F",X"77",
		X"C3",X"DB",X"FB",X"DB",X"9B",X"79",X"EF",X"BE",X"BF",X"9F",X"FA",X"60",X"A0",X"10",X"00",X"00",
		X"E0",X"F0",X"30",X"30",X"F0",X"E0",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"F8",X"F8",X"FC",X"FC",X"C0",X"EA",X"BE",X"BF",
		X"3F",X"3F",X"5F",X"5F",X"7F",X"FF",X"FF",X"FE",X"FE",X"FE",X"5C",X"00",X"00",X"80",X"C4",X"FE",
		X"7F",X"3F",X"9C",X"9C",X"DC",X"EC",X"7C",X"7C",X"DE",X"DF",X"BF",X"F6",X"EE",X"DE",X"DE",X"8C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"0F",X"BF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"E7",X"F9",X"FE",X"FC",X"F1",X"03",X"1F",X"3F",X"3F",X"7F",X"7A",X"38",X"90",X"C0",
		X"E0",X"F0",X"C0",X"60",X"30",X"08",X"20",X"20",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"80",
		X"C0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"40",X"60",X"00",X"10",X"10",X"18",X"18",
		X"E0",X"F0",X"F8",X"F0",X"78",X"0C",X"00",X"18",X"10",X"40",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C7",X"63",X"73",X"33",X"33",X"33",X"33",X"33",X"33",X"63",X"C3",X"81",X"00",X"00",X"00",X"00",
		X"F8",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"F8",
		X"00",X"00",X"00",X"00",X"F0",X"19",X"1D",X"0C",X"0C",X"0C",X"FC",X"0C",X"0C",X"18",X"B0",X"E1",
		X"BE",X"E7",X"83",X"83",X"87",X"9E",X"BC",X"E0",X"80",X"86",X"CE",X"FC",X"00",X"00",X"00",X"00",
		X"1E",X"8C",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"8C",X"0E",X"08",X"00",X"00",X"0C",X"0C",
		X"1E",X"8C",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CE",X"8F",X"07",X"00",X"00",X"00",X"00",
		X"0E",X"1F",X"17",X"10",X"30",X"30",X"38",X"78",X"58",X"5C",X"CC",X"8C",X"8C",X"8E",X"06",X"8F",
		X"C0",X"E0",X"60",X"20",X"00",X"00",X"00",X"00",X"C0",X"E0",X"E0",X"60",X"60",X"E0",X"C0",X"80",
		X"C3",X"E6",X"6C",X"28",X"00",X"00",X"CF",X"EC",X"6C",X"66",X"63",X"C1",X"00",X"00",X"00",X"00",
		X"7B",X"31",X"31",X"31",X"31",X"31",X"31",X"71",X"71",X"F1",X"B9",X"21",X"00",X"00",X"00",X"00",
		X"38",X"7C",X"4C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"7F",X"0E",X"0C",X"08",X"08",
		X"87",X"CC",X"D8",X"D0",X"C0",X"80",X"1F",X"18",X"18",X"8C",X"86",X"03",X"00",X"00",X"00",X"00",
		X"7C",X"38",X"38",X"38",X"38",X"38",X"38",X"38",X"F8",X"38",X"38",X"38",X"38",X"38",X"38",X"FC",
		X"FE",X"87",X"83",X"E6",X"FC",X"3E",X"06",X"1C",X"78",X"CC",X"86",X"86",X"86",X"86",X"CC",X"78",
		X"DE",X"8C",X"8C",X"8C",X"8C",X"8C",X"8C",X"8C",X"8C",X"8C",X"CE",X"08",X"00",X"00",X"0C",X"0C",
		X"F8",X"70",X"70",X"70",X"70",X"70",X"F0",X"F0",X"F0",X"70",X"70",X"70",X"70",X"70",X"70",X"F8",
		X"06",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C3",X"E3",X"E3",X"F3",X"F3",X"F3",X"F3",X"F3",X"F3",X"E3",X"EF",X"CF",X"03",X"03",X"00",X"00",
		X"FC",X"FC",X"FC",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",
		X"00",X"00",X"00",X"00",X"F8",X"DC",X"8E",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8E",X"DC",X"F8",
		X"E0",X"F8",X"3C",X"1E",X"1E",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1E",X"1E",X"3C",X"F8",X"E0",
		X"0F",X"1D",X"38",X"78",X"78",X"00",X"00",X"78",X"78",X"38",X"1D",X"0F",X"00",X"00",X"00",X"00",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"EF",X"FF",X"F7",X"E7",X"00",X"00",X"00",X"00",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",
		X"01",X"83",X"87",X"CF",X"CF",X"C0",X"C0",X"CF",X"CF",X"87",X"83",X"01",X"00",X"00",X"00",X"00",
		X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"7B",X"7B",X"7B",X"03",X"00",X"78",X"78",X"78",
		X"1F",X"3B",X"71",X"F1",X"F1",X"01",X"FF",X"FF",X"F1",X"71",X"3B",X"1F",X"00",X"00",X"00",X"00",
		X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"BE",X"FF",X"DF",X"8E",X"00",X"00",X"00",X"00",
		X"E0",X"E0",X"E0",X"FF",X"FF",X"F0",X"F0",X"78",X"78",X"3D",X"3D",X"3F",X"1F",X"1F",X"0F",X"0F",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"07",X"07",X"01",X"01",X"07",X"07",
		X"F8",X"DC",X"8E",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8E",X"DC",X"F8",X"00",X"00",X"00",X"00",
		X"1F",X"3B",X"71",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"71",X"3B",X"1F",X"00",X"00",X"00",X"00",
		X"BC",X"FE",X"DE",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"DE",X"FE",X"BC",X"80",X"80",X"80",X"80",
		X"78",X"78",X"78",X"79",X"79",X"78",X"79",X"79",X"F9",X"F8",X"78",X"78",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"8F",X"CF",X"CF",X"CF",X"CF",X"CF",X"CF",X"8F",X"3F",X"3F",X"0F",X"0F",X"00",X"00",
		X"79",X"79",X"79",X"79",X"79",X"79",X"79",X"79",X"F9",X"F9",X"79",X"78",X"00",X"01",X"01",X"01",
		X"81",X"C1",X"C1",X"E1",X"E1",X"B1",X"B1",X"99",X"99",X"8D",X"8D",X"87",X"87",X"83",X"83",X"81",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"C0",X"F0",X"FC",X"C6",X"D9",X"FE",X"FF",X"CF",X"C3",X"C1",X"C0",X"C0",X"C0",X"C0",X"C1",
		X"C0",X"C0",X"C0",X"F0",X"F0",X"C0",X"C0",X"E0",X"70",X"30",X"30",X"30",X"30",X"60",X"40",X"00",
		X"00",X"40",X"60",X"30",X"30",X"30",X"30",X"30",X"30",X"60",X"40",X"00",X"00",X"40",X"60",X"30",
		X"00",X"00",X"01",X"02",X"05",X"05",X"8B",X"CB",X"D6",X"FE",X"FC",X"7F",X"7F",X"3C",X"30",X"00",
		X"E0",X"B0",X"10",X"B0",X"F0",X"78",X"7C",X"CC",X"8C",X"8C",X"9C",X"FC",X"F8",X"F8",X"F0",X"E0",
		X"EF",X"E7",X"A6",X"8C",X"EE",X"24",X"A6",X"F3",X"FF",X"2E",X"63",X"30",X"84",X"86",X"82",X"00",
		X"00",X"00",X"00",X"00",X"20",X"60",X"C0",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"02",X"00",X"00",X"00",X"01",X"03",X"03",X"0F",X"03",X"0D",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"0F",X"0F",X"07",X"0F",X"03",X"0D",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"8F",X"CF",X"C7",X"8F",X"83",X"0D",
		X"7E",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"3C",X"00",X"00",X"00",
		X"F8",X"1C",X"0C",X"30",X"70",X"38",X"3C",X"1C",X"0C",X"18",X"30",X"30",X"34",X"BC",X"1C",X"08",
		X"00",X"10",X"08",X"00",X"00",X"00",X"00",X"00",X"40",X"20",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"80",X"80",X"80",X"80",X"80",X"C0",X"C0",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"84",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"3E",X"7E",X"7C",X"7E",X"73",X"D9",X"DC",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"0F",
		X"0E",X"1C",X"19",X"13",X"17",X"37",X"2F",X"2F",X"EF",X"DF",X"DF",X"BF",X"AF",X"0F",X"07",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"01",X"00",
		X"00",X"03",X"07",X"0C",X"08",X"0A",X"08",X"08",X"09",X"0F",X"07",X"03",X"02",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"03",X"0D",X"1F",X"11",X"3F",X"7F",X"7F",X"1F",X"1F",X"2F",X"07",X"03",X"03",X"01",X"00",
		X"FE",X"86",X"00",X"00",X"C0",X"C0",X"E0",X"E1",X"43",X"06",X"0C",X"0C",X"8D",X"2F",X"07",X"02",
		X"00",X"00",X"18",X"BC",X"FC",X"7E",X"FE",X"FE",X"8E",X"8E",X"CE",X"FC",X"7C",X"38",X"F0",X"00",
		X"E0",X"F0",X"A0",X"00",X"00",X"54",X"FC",X"F8",X"34",X"18",X"50",X"D0",X"18",X"F8",X"F0",X"C0",
		X"00",X"00",X"F8",X"FC",X"A8",X"54",X"FC",X"F8",X"34",X"58",X"50",X"10",X"18",X"F8",X"F0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"C0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"00",X"0B",X"1F",X"1F",X"3C",X"70",X"00",
		X"07",X"0F",X"1F",X"1F",X"0F",X"0F",X"0F",X"07",X"07",X"07",X"07",X"03",X"03",X"03",X"03",X"03",
		X"00",X"00",X"00",X"10",X"78",X"5C",X"6C",X"74",X"6C",X"34",X"19",X"00",X"01",X"01",X"00",X"00",
		X"00",X"07",X"0F",X"0F",X"1F",X"3F",X"3F",X"0F",X"0F",X"17",X"03",X"07",X"0F",X"06",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"83",X"0F",X"1F",X"78",X"F0",
		X"60",X"C1",X"87",X"0F",X"1F",X"3F",X"1F",X"0F",X"0F",X"07",X"07",X"03",X"03",X"03",X"03",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"03",X"00",X"00",X"00",X"80",X"C0",X"00",X"00",X"00",X"04",X"02",X"01",X"0B",X"1E",
		X"7C",X"F8",X"C1",X"03",X"0F",X"3F",X"7F",X"7F",X"3F",X"1F",X"0F",X"07",X"07",X"03",X"03",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"C0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"1B",
		X"FE",X"FF",X"FF",X"FF",X"FF",X"7F",X"2F",X"0F",X"1F",X"07",X"03",X"07",X"0F",X"06",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"03",X"0F",X"1F",X"9E",X"0E",X"0C",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",
		X"00",X"07",X"0F",X"0F",X"1F",X"3F",X"3F",X"0F",X"17",X"07",X"03",X"07",X"0F",X"06",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"08",X"00",X"00",X"00",X"00",X"00",X"40",X"20",X"20",X"00",
		X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"FF",
		X"06",X"98",X"00",X"00",X"00",X"04",X"00",X"00",X"10",X"00",X"00",X"C0",X"C0",X"60",X"C0",X"80",
		X"00",X"00",X"04",X"04",X"04",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"8C",X"06",X"02",X"02",X"06",X"8C",X"F8",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"04",X"04",X"04",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"8C",X"06",X"02",X"02",X"06",X"8C",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F1",X"E7",X"C3",X"01",X"41",X"81",X"85",X"8D",X"8D",X"C5",X"C1",X"E3",X"FF",X"FC",X"FC",X"FC",
		X"FC",X"F8",X"F9",X"F9",X"F1",X"F3",X"F3",X"E3",X"E7",X"C7",X"C7",X"CF",X"8F",X"8F",X"1F",X"1F",
		X"8F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",
		X"F8",X"FA",X"FB",X"F3",X"F7",X"F7",X"E7",X"EF",X"EF",X"CF",X"CF",X"9F",X"9F",X"1F",X"3F",X"3F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"1F",X"00",X"0C",X"0F",X"1F",X"1F",X"3F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"00",X"C0",X"FF",
		X"C3",X"C1",X"E0",X"E0",X"F0",X"FC",X"FF",X"FE",X"F1",X"87",X"1F",X"7F",X"FF",X"FF",X"FF",X"FF",
		X"30",X"0F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",
		X"00",X"00",X"C0",X"C0",X"F0",X"F8",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"3F",X"0F",X"03",X"00",
		X"F8",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"80",X"DC",X"C0",X"E0",X"E0",X"E0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"E0",X"E0",X"E0",X"F0",X"F0",X"F8",X"F8",X"F8",X"D8",X"DC",
		X"54",X"8C",X"FC",X"FC",X"78",X"FC",X"FC",X"AC",X"54",X"50",X"30",X"00",X"00",X"00",X"00",X"00",
		X"6F",X"7F",X"7F",X"7E",X"7D",X"7B",X"7B",X"37",X"07",X"0F",X"07",X"07",X"0F",X"1F",X"1F",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"30",X"E0",X"EF",X"DF",X"DF",X"BF",X"BF",X"F0",X"EF",X"DF",X"9F",X"3F",X"7F",X"67",
		X"C1",X"83",X"0F",X"3F",X"5F",X"5F",X"4F",X"6F",X"67",X"73",X"79",X"BC",X"38",X"70",X"FC",X"FE",
		X"FF",X"8F",X"8F",X"07",X"05",X"ED",X"7B",X"DF",X"DF",X"3F",X"5F",X"17",X"0E",X"0D",X"0C",X"18",
		X"00",X"00",X"00",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"F0",X"80",X"80",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"00",X"00",X"00",X"00",X"00",X"40",
		X"20",X"A0",X"80",X"00",X"00",X"06",X"84",X"80",X"80",X"80",X"80",X"A0",X"A0",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"03",X"03",X"07",X"07",X"0F",X"0F",X"0F",X"0F",X"07",X"07",X"07",X"07",
		X"00",X"00",X"00",X"00",X"00",X"06",X"1E",X"07",X"3F",X"0F",X"03",X"07",X"0E",X"00",X"00",X"00",
		X"00",X"00",X"F0",X"78",X"78",X"1D",X"3F",X"FF",X"FE",X"FE",X"FE",X"FE",X"FD",X"F9",X"F8",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"06",X"4D",X"7F",X"3F",X"1E",X"1C",X"00",X"01",X"01",X"01",X"05",X"0C",X"1E",X"1E",X"1F",
		X"3F",X"3F",X"3F",X"3F",X"7F",X"7F",X"7F",X"3F",X"3F",X"1E",X"1E",X"1E",X"1E",X"1E",X"1C",X"1C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F8",X"FC",X"FE",X"FE",X"FF",X"FF",
		X"FF",X"FE",X"FE",X"FE",X"FE",X"FD",X"F1",X"01",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"F0",X"FC",X"7F",X"7D",X"2F",X"AF",X"EC",X"FE",X"FE",X"5C",X"DE",X"BE",X"F9",X"E6",X"7C",
		X"00",X"08",X"9C",X"7E",X"5E",X"5E",X"BE",X"BF",X"7D",X"7D",X"75",X"78",X"7D",X"3F",X"3F",X"3F",
		X"7E",X"DE",X"FE",X"FE",X"3E",X"7C",X"5C",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"E0",X"F0",X"F8",X"FC",X"FF",X"FF",X"FF",X"FF",X"7F",
		X"7F",X"00",X"3F",X"4F",X"3F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",X"E7",
		X"07",X"0F",X"1F",X"4F",X"67",X"73",X"79",X"3C",X"B3",X"AF",X"8F",X"BE",X"73",X"ED",X"DE",X"DE",
		X"DF",X"E6",X"58",X"0A",X"0D",X"07",X"03",X"C1",X"F9",X"DF",X"DF",X"82",X"6A",X"EA",X"FE",X"7C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"FF",X"1F",X"E3",X"FD",X"FE",X"FF",X"FD",X"FE",
		X"FE",X"FE",X"FC",X"F8",X"F0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"04",X"80",X"C0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"00",X"10",X"08",X"00",X"00",X"00",X"0D",X"3F",X"BC",X"9F",X"5C",X"FF",X"FD",X"F6",X"E0",X"C0",
		X"C3",X"81",X"11",X"D4",X"AF",X"6F",X"4F",X"C0",X"6F",X"6F",X"6F",X"E0",X"FE",X"FA",X"FD",X"F5",
		X"ED",X"1B",X"B7",X"5F",X"8F",X"3F",X"5B",X"27",X"1C",X"02",X"03",X"03",X"03",X"06",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"BC",X"7F",X"07",X"7F",X"BF",X"FF",X"FE",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"70",X"E8",X"D8",X"F0",X"EC",X"FC",X"F8",X"C0",
		X"E0",X"60",X"00",X"36",X"2A",X"7E",X"5F",X"5F",X"3F",X"1F",X"1F",X"3F",X"3F",X"71",X"6A",X"FB",
		X"FB",X"FA",X"7E",X"FE",X"FC",X"FC",X"F8",X"70",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"81",X"07",X"0F",X"9F",X"BE",X"71",X"6F",
		X"5F",X"BF",X"BF",X"7F",X"6F",X"DF",X"DF",X"DF",X"0F",X"0F",X"1F",X"16",X"19",X"1F",X"0F",X"06",
		X"09",X"0E",X"0F",X"0F",X"07",X"03",X"07",X"3F",X"7E",X"FC",X"CF",X"B7",X"FB",X"78",X"3F",X"08",
		X"0B",X"15",X"15",X"0E",X"3F",X"71",X"0E",X"0F",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"80",X"80",X"8C",X"9C",X"15",X"3B",X"BB",X"35",X"1E",X"3F",X"3F",X"3F",X"3F",X"3F",X"3E",
		X"3E",X"3E",X"3E",X"7C",X"7C",X"B8",X"E8",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"07",X"0B",
		X"0B",X"1B",X"1C",X"9B",X"D7",X"1B",X"0F",X"03",X"07",X"07",X"07",X"0F",X"0F",X"0F",X"1F",X"1F",
		X"1F",X"1F",X"EF",X"CF",X"AE",X"B6",X"BA",X"FC",X"3D",X"19",X"02",X"00",X"7E",X"FE",X"FE",X"F7",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"40",X"40",X"40",X"80",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"19",X"1F",X"37",X"2F",
		X"2F",X"7E",X"79",X"77",X"77",X"03",X"07",X"07",X"04",X"06",X"0E",X"0F",X"0F",X"1F",X"1F",X"1F",
		X"39",X"77",X"EF",X"EF",X"E7",X"58",X"DE",X"F8",X"5D",X"89",X"02",X"00",X"7E",X"FE",X"FE",X"F7",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",
		X"80",X"80",X"80",X"00",X"00",X"00",X"80",X"80",X"80",X"C0",X"C0",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"E0",X"D0",X"40",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"06",X"0E",X"1E",X"1F",X"3F",X"3F",X"3F",X"3F",X"3F",X"1F",
		X"0F",X"0E",X"01",X"C7",X"EF",X"E3",X"F3",X"CF",X"9A",X"AF",X"EF",X"F7",X"7F",X"7F",X"3F",X"1F",
		X"1B",X"5D",X"6D",X"3B",X"02",X"3A",X"3E",X"3C",X"1D",X"09",X"02",X"00",X"7E",X"FE",X"FE",X"F7",
		X"EB",X"FB",X"FB",X"F7",X"BF",X"1E",X"0D",X"03",X"03",X"03",X"83",X"07",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"08",X"14",X"2E",X"77",X"75",X"4B",X"FE",X"FC",X"FC",
		X"FC",X"FC",X"F8",X"F8",X"F0",X"E0",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"C6",X"E0",X"E0",X"C0",X"C0",X"C0",X"80",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"01",X"03",X"07",X"04",X"03",X"07",X"07",X"03",X"00",
		X"01",X"03",X"07",X"03",X"03",X"03",X"07",X"07",X"0F",X"0F",X"2F",X"FF",X"FE",X"FE",X"DE",X"46",
		X"C1",X"E7",X"A2",X"A9",X"AC",X"2E",X"27",X"97",X"03",X"01",X"03",X"1F",X"3F",X"7E",X"7C",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"04",X"C0",X"E8",X"E0",X"E0",X"E0",
		X"60",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"80",
		X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"1C",X"3E",X"3F",X"1F",X"1F",X"0F",X"0E",X"06",X"03",
		X"02",X"01",X"03",X"3F",X"7F",X"7F",X"FF",X"BF",X"7C",X"69",X"0A",X"0F",X"1F",X"1F",X"3F",X"72",
		X"00",X"46",X"67",X"63",X"69",X"6C",X"2E",X"27",X"17",X"03",X"01",X"03",X"1F",X"3F",X"7F",X"7F",
		X"80",X"80",X"80",X"80",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"40",X"00",X"00",X"00",X"40",X"00",X"40",X"00",
		X"00",X"00",X"00",X"00",X"80",X"00",X"30",X"3C",X"7E",X"7E",X"3E",X"3E",X"6C",X"44",X"6C",X"6C",
		X"6C",X"78",X"F8",X"F0",X"70",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"8F",X"0F",X"1F",X"1F",X"1F",X"1F",X"0F",X"0F",X"06",
		X"01",X"03",X"07",X"03",X"03",X"03",X"07",X"07",X"0F",X"0F",X"0F",X"1F",X"1F",X"3F",X"3F",X"82",
		X"81",X"67",X"E3",X"E9",X"EC",X"2E",X"27",X"17",X"03",X"01",X"03",X"1F",X"3F",X"7E",X"7C",X"FC",
		X"FD",X"C3",X"BB",X"76",X"7E",X"7A",X"33",X"01",X"00",X"00",X"01",X"00",X"18",X"1C",X"08",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"08",X"08",X"00",X"90",X"C0",X"C0",X"C0",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"E0",X"F0",X"F0",X"F0",X"F0",X"88",X"98",X"D8",X"E8",X"68",X"78",X"F8",
		X"70",X"A8",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"03",X"0F",X"1F",X"3F",X"3F",X"3E",X"3E",X"1D",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"7C",X"7F",X"7F",X"3F",X"3F",X"1F",X"1F",X"0F",
		X"06",X"01",X"03",X"07",X"03",X"03",X"03",X"07",X"07",X"0F",X"8F",X"CF",X"FF",X"FF",X"FF",X"32",
		X"01",X"47",X"67",X"63",X"69",X"6C",X"2E",X"27",X"17",X"03",X"01",X"03",X"1F",X"3F",X"7F",X"7F",
		X"07",X"07",X"00",X"07",X"0F",X"07",X"07",X"07",X"0F",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"BE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"80",X"80",X"80",X"80",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"0F",X"0F",X"9F",
		X"1F",X"0E",X"01",X"03",X"07",X"03",X"03",X"03",X"07",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",X"BE",
		X"91",X"03",X"47",X"67",X"63",X"69",X"6C",X"2E",X"27",X"17",X"03",X"01",X"03",X"1F",X"3F",X"7F",
		X"BE",X"FD",X"C3",X"BB",X"76",X"7F",X"7A",X"33",X"01",X"00",X"00",X"01",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
