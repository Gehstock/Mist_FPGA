library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity rom is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of rom is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"31",X"A0",X"20",X"97",X"00",X"C3",X"B6",X"00",X"C5",X"D5",X"E5",X"F5",X"C3",X"37",X"02",X"00",
		X"C3",X"08",X"00",X"C2",X"28",X"00",X"C9",X"00",X"C5",X"06",X"A0",X"0E",X"A0",X"0D",X"C2",X"1D",
		X"00",X"05",X"D3",X"06",X"C3",X"45",X"01",X"00",X"1A",X"77",X"13",X"23",X"05",X"C3",X"13",X"00",
		X"32",X"A1",X"20",X"32",X"A2",X"20",X"D3",X"01",X"00",X"06",X"0D",X"21",X"A3",X"20",X"11",X"FF",
		X"00",X"EF",X"C3",X"50",X"01",X"CD",X"CB",X"09",X"FB",X"CD",X"43",X"09",X"00",X"00",X"C3",X"D0",
		X"06",X"11",X"18",X"01",X"06",X"08",X"EF",X"21",X"40",X"21",X"06",X"08",X"EF",X"21",X"80",X"21",
		X"06",X"08",X"EF",X"21",X"C0",X"21",X"06",X"08",X"EF",X"06",X"05",X"21",X"F6",X"20",X"EF",X"21",
		X"00",X"00",X"22",X"ED",X"20",X"3E",X"05",X"32",X"00",X"22",X"21",X"01",X"20",X"36",X"00",X"23",
		X"7D",X"FE",X"24",X"DA",X"7D",X"00",X"21",X"20",X"26",X"36",X"00",X"23",X"7C",X"FE",X"3F",X"C2",
		X"89",X"00",X"21",X"27",X"00",X"22",X"03",X"20",X"D3",X"06",X"CD",X"AE",X"1E",X"3A",X"F5",X"20",
		X"A7",X"C2",X"42",X"03",X"3A",X"EF",X"20",X"FE",X"02",X"C2",X"98",X"00",X"C3",X"39",X"00",X"32",
		X"E8",X"20",X"C3",X"B9",X"06",X"00",X"32",X"F5",X"20",X"C3",X"30",X"00",X"3A",X"F5",X"20",X"A7",
		X"C3",X"84",X"03",X"C5",X"D5",X"E5",X"3A",X"E2",X"20",X"A7",X"C2",X"D3",X"00",X"2A",X"A5",X"20",
		X"C3",X"D6",X"00",X"2A",X"A9",X"20",X"78",X"01",X"20",X"00",X"FE",X"11",X"D2",X"EA",X"00",X"01",
		X"50",X"00",X"FE",X"0E",X"D2",X"EA",X"00",X"01",X"00",X"01",X"CD",X"2A",X"13",X"A7",X"C2",X"4A",
		X"01",X"22",X"A5",X"20",X"CD",X"40",X"0B",X"E1",X"D1",X"C1",X"3E",X"28",X"C3",X"31",X"13",X"2D",
		X"25",X"00",X"00",X"23",X"25",X"00",X"00",X"36",X"25",X"00",X"00",X"00",X"5D",X"29",X"00",X"18",
		X"41",X"27",X"00",X"1A",X"01",X"35",X"00",X"1A",X"82",X"3E",X"00",X"13",X"87",X"2F",X"00",X"13",
		X"FC",X"28",X"00",X"12",X"92",X"36",X"00",X"12",X"FC",X"3E",X"00",X"12",X"95",X"2F",X"00",X"12",
		X"F9",X"28",X"00",X"11",X"92",X"2F",X"00",X"11",X"00",X"08",X"48",X"88",X"C8",X"00",X"00",X"01",
		X"FE",X"00",X"00",X"FF",X"FF",X"C2",X"1B",X"00",X"C1",X"C9",X"22",X"A9",X"20",X"C3",X"7E",X"03",
		X"21",X"ED",X"20",X"11",X"3D",X"01",X"06",X"08",X"EF",X"C3",X"45",X"00",X"21",X"75",X"00",X"C3",
		X"03",X"09",X"00",X"00",X"00",X"00",X"3A",X"F1",X"20",X"FE",X"01",X"C2",X"FF",X"01",X"3A",X"E0",
		X"20",X"A7",X"CA",X"0C",X"06",X"3D",X"32",X"E0",X"20",X"3E",X"01",X"32",X"F5",X"20",X"E1",X"C9",
		X"00",X"3A",X"E2",X"20",X"A7",X"C2",X"B2",X"01",X"3A",X"E0",X"20",X"A7",X"C2",X"95",X"01",X"CD",
		X"DE",X"05",X"C3",X"A1",X"01",X"3D",X"32",X"E0",X"20",X"C3",X"A1",X"01",X"3E",X"03",X"C3",X"8F",
		X"04",X"3E",X"01",X"32",X"E2",X"20",X"CD",X"C7",X"03",X"11",X"98",X"0B",X"21",X"0C",X"31",X"C3",
		X"D5",X"01",X"97",X"32",X"E2",X"20",X"3A",X"E1",X"20",X"A7",X"C2",X"F8",X"01",X"00",X"00",X"00",
		X"00",X"CD",X"EC",X"05",X"3A",X"E0",X"20",X"A7",X"C2",X"CF",X"01",X"C3",X"AD",X"02",X"00",X"CD",
		X"C7",X"03",X"21",X"0C",X"31",X"0E",X"08",X"CD",X"F1",X"09",X"CD",X"73",X"04",X"11",X"ED",X"22",
		X"0E",X"50",X"CD",X"22",X"02",X"21",X"00",X"21",X"11",X"00",X"23",X"0E",X"FF",X"CD",X"CF",X"05",
		X"3E",X"01",X"32",X"F5",X"20",X"C3",X"29",X"03",X"3D",X"32",X"E1",X"20",X"C3",X"CF",X"01",X"97",
		X"D3",X"05",X"00",X"C3",X"81",X"01",X"7C",X"FE",X"27",X"C2",X"2A",X"19",X"7D",X"A7",X"C2",X"2A",
		X"19",X"C3",X"C6",X"1B",X"3E",X"01",X"32",X"D6",X"20",X"13",X"23",X"44",X"4D",X"E1",X"C9",X"00",
		X"00",X"00",X"7E",X"47",X"1A",X"77",X"78",X"12",X"13",X"23",X"0D",X"C2",X"22",X"02",X"C9",X"F3",
		X"76",X"CA",X"3D",X"03",X"C3",X"93",X"02",X"3A",X"F5",X"20",X"A7",X"CA",X"E4",X"17",X"C3",X"EA",
		X"17",X"C2",X"54",X"1F",X"CD",X"92",X"1F",X"C9",X"C2",X"ED",X"1E",X"CD",X"92",X"1F",X"C3",X"1E",
		X"1F",X"CD",X"D2",X"15",X"C3",X"D2",X"1D",X"3A",X"E6",X"20",X"3C",X"32",X"E6",X"20",X"C3",X"51",
		X"02",X"3A",X"E5",X"20",X"3C",X"32",X"E5",X"20",X"C3",X"51",X"02",X"3A",X"E4",X"20",X"3C",X"32",
		X"E4",X"20",X"C3",X"51",X"02",X"3A",X"E3",X"20",X"3C",X"32",X"E3",X"20",X"C3",X"51",X"02",X"21",
		X"00",X"21",X"97",X"32",X"E3",X"20",X"C9",X"97",X"32",X"E4",X"20",X"21",X"C0",X"21",X"C9",X"00",
		X"00",X"00",X"00",X"11",X"B0",X"20",X"2A",X"D3",X"20",X"E5",X"D5",X"CD",X"B4",X"15",X"D1",X"E1",
		X"3A",X"D6",X"20",X"A7",X"C2",X"D9",X"03",X"CD",X"96",X"15",X"C3",X"DE",X"15",X"3A",X"E1",X"20",
		X"A7",X"CA",X"EE",X"04",X"C3",X"A1",X"01",X"3A",X"E0",X"20",X"A7",X"CA",X"EE",X"04",X"C3",X"CF",
		X"01",X"3A",X"F6",X"20",X"FE",X"0A",X"DA",X"D6",X"06",X"11",X"00",X"14",X"CD",X"06",X"15",X"11",
		X"B0",X"20",X"21",X"F0",X"32",X"22",X"D3",X"20",X"CD",X"B4",X"15",X"3A",X"D6",X"20",X"FE",X"01",
		X"CA",X"1C",X"03",X"C3",X"78",X"03",X"00",X"CD",X"96",X"15",X"97",X"32",X"D1",X"20",X"32",X"DA",
		X"20",X"32",X"D7",X"20",X"32",X"D9",X"20",X"32",X"E8",X"20",X"3E",X"02",X"00",X"32",X"F5",X"20",
		X"3E",X"05",X"32",X"00",X"20",X"3E",X"10",X"32",X"D2",X"20",X"3E",X"02",X"32",X"DD",X"20",X"32",
		X"CF",X"20",X"3E",X"10",X"32",X"D5",X"20",X"3E",X"01",X"32",X"D8",X"20",X"97",X"32",X"D6",X"20",
		X"32",X"D0",X"20",X"00",X"00",X"00",X"C3",X"66",X"13",X"97",X"32",X"F6",X"20",X"C3",X"EE",X"08",
		X"FE",X"12",X"C2",X"94",X"03",X"78",X"A7",X"C2",X"1C",X"03",X"C3",X"9E",X"03",X"D5",X"C5",X"C3",
		X"C1",X"02",X"06",X"00",X"DB",X"01",X"E6",X"08",X"CA",X"4E",X"03",X"3E",X"21",X"47",X"3A",X"E8",
		X"20",X"A7",X"CA",X"5E",X"03",X"3D",X"32",X"E8",X"20",X"3E",X"22",X"C3",X"60",X"03",X"3E",X"20",
		X"B0",X"D3",X"03",X"C3",X"89",X"05",X"32",X"DA",X"20",X"00",X"3E",X"02",X"32",X"E8",X"20",X"21",
		X"EA",X"20",X"34",X"C3",X"41",X"16",X"00",X"00",X"01",X"60",X"00",X"C3",X"8E",X"03",X"CD",X"48",
		X"0B",X"C3",X"F7",X"00",X"CA",X"33",X"13",X"3E",X"20",X"D3",X"03",X"C3",X"C3",X"00",X"21",X"8D",
		X"31",X"5D",X"54",X"46",X"23",X"7E",X"B0",X"47",X"7D",X"E6",X"1F",X"C3",X"30",X"03",X"EB",X"09",
		X"7C",X"FE",X"34",X"C2",X"91",X"03",X"21",X"F0",X"32",X"11",X"B0",X"20",X"C3",X"E7",X"02",X"21",
		X"00",X"00",X"22",X"EB",X"20",X"22",X"DB",X"20",X"11",X"0C",X"01",X"21",X"C0",X"22",X"06",X"0C",
		X"EF",X"97",X"32",X"CE",X"22",X"C9",X"00",X"D3",X"06",X"21",X"20",X"26",X"36",X"00",X"23",X"7C",
		X"FE",X"3F",X"C2",X"CC",X"03",X"11",X"90",X"0B",X"C9",X"3E",X"24",X"D3",X"03",X"3A",X"AF",X"20",
		X"FE",X"A0",X"CA",X"96",X"13",X"3C",X"32",X"AF",X"20",X"C3",X"AE",X"13",X"97",X"32",X"AF",X"20",
		X"3E",X"00",X"D3",X"03",X"C3",X"D3",X"04",X"57",X"7B",X"E6",X"E0",X"5F",X"19",X"C3",X"B3",X"17",
		X"CD",X"48",X"0B",X"C3",X"F7",X"00",X"FE",X"A0",X"D2",X"9F",X"1F",X"3C",X"32",X"F6",X"20",X"C9",
		X"3A",X"EA",X"20",X"FE",X"20",X"DA",X"24",X"04",X"3E",X"20",X"32",X"EA",X"20",X"3E",X"10",X"D3",
		X"05",X"C3",X"9F",X"1F",X"3A",X"F6",X"20",X"C3",X"0B",X"04",X"97",X"32",X"EA",X"20",X"D3",X"05",
		X"C3",X"C8",X"18",X"3A",X"E2",X"20",X"2A",X"A5",X"20",X"A7",X"CA",X"40",X"04",X"2A",X"A9",X"20",
		X"3A",X"EF",X"20",X"01",X"00",X"02",X"FE",X"01",X"D2",X"4E",X"04",X"01",X"00",X"03",X"CD",X"EB",
		X"0B",X"3A",X"E2",X"20",X"A7",X"C2",X"61",X"04",X"22",X"A5",X"20",X"CD",X"40",X"0B",X"C3",X"67",
		X"04",X"22",X"A9",X"20",X"CD",X"48",X"0B",X"11",X"0C",X"01",X"06",X"0C",X"21",X"C0",X"20",X"EF",
		X"C3",X"C8",X"18",X"06",X"06",X"DF",X"05",X"C2",X"75",X"04",X"21",X"C0",X"20",X"11",X"C0",X"22",
		X"0E",X"10",X"CD",X"22",X"02",X"21",X"ED",X"20",X"C9",X"D3",X"02",X"DB",X"03",X"3E",X"12",X"6F",
		X"E6",X"30",X"0F",X"0F",X"B5",X"E6",X"0F",X"C9",X"E5",X"D5",X"11",X"80",X"00",X"19",X"7E",X"D1",
		X"E1",X"A7",X"C2",X"2A",X"19",X"C3",X"C6",X"1B",X"3E",X"20",X"D3",X"03",X"97",X"D3",X"05",X"C3",
		X"4E",X"00",X"23",X"7E",X"BA",X"00",X"00",X"00",X"C3",X"38",X"0B",X"97",X"32",X"EA",X"20",X"C3",
		X"AF",X"00",X"32",X"ED",X"20",X"32",X"EE",X"20",X"32",X"EA",X"20",X"D3",X"05",X"3E",X"05",X"32",
		X"00",X"22",X"C9",X"3E",X"01",X"32",X"DF",X"20",X"CD",X"88",X"17",X"26",X"20",X"3A",X"00",X"22",
		X"6F",X"CD",X"8D",X"18",X"97",X"32",X"DF",X"20",X"CD",X"88",X"17",X"C3",X"62",X"01",X"2A",X"A1",
		X"20",X"44",X"4D",X"2A",X"A5",X"20",X"EB",X"2A",X"A9",X"20",X"7A",X"BC",X"DA",X"08",X"05",X"C2",
		X"07",X"05",X"7B",X"BD",X"DA",X"08",X"05",X"EB",X"7C",X"B8",X"DA",X"18",X"05",X"C2",X"15",X"05",
		X"7D",X"B9",X"DA",X"18",X"05",X"22",X"A1",X"20",X"CD",X"4C",X"06",X"21",X"20",X"26",X"36",X"00",
		X"23",X"7C",X"FE",X"3F",X"C3",X"3F",X"06",X"0E",X"04",X"21",X"0E",X"2F",X"11",X"70",X"0B",X"CD",
		X"F1",X"09",X"3A",X"AD",X"20",X"FE",X"02",X"D2",X"4A",X"05",X"A7",X"CA",X"38",X"06",X"11",X"2D",
		X"09",X"C3",X"28",X"06",X"CD",X"F1",X"09",X"C3",X"30",X"06",X"11",X"74",X"0B",X"21",X"05",X"31",
		X"C3",X"23",X"06",X"31",X"9F",X"20",X"21",X"42",X"00",X"22",X"9F",X"20",X"00",X"C9",X"C3",X"7A",
		X"06",X"FE",X"04",X"D2",X"6E",X"06",X"DB",X"03",X"E6",X"80",X"C2",X"6E",X"06",X"11",X"B0",X"20",
		X"2A",X"D3",X"20",X"CD",X"B4",X"15",X"3A",X"CE",X"20",X"FE",X"01",X"CA",X"BC",X"05",X"FE",X"02",
		X"CA",X"C2",X"05",X"21",X"9A",X"29",X"C3",X"5F",X"06",X"3A",X"E3",X"20",X"47",X"3A",X"E4",X"20",
		X"B0",X"47",X"3A",X"E5",X"20",X"B0",X"47",X"3A",X"E6",X"20",X"B0",X"A7",X"CA",X"A8",X"04",X"C3",
		X"98",X"00",X"97",X"32",X"E5",X"20",X"21",X"40",X"21",X"C9",X"97",X"32",X"E6",X"20",X"21",X"80",
		X"21",X"C9",X"21",X"00",X"00",X"22",X"A5",X"20",X"22",X"A9",X"20",X"C9",X"21",X"42",X"3A",X"C3",
		X"86",X"05",X"21",X"83",X"2B",X"C3",X"86",X"05",X"97",X"32",X"CE",X"20",X"C3",X"71",X"06",X"CD",
		X"22",X"02",X"21",X"CE",X"20",X"11",X"CE",X"22",X"0E",X"01",X"CD",X"22",X"02",X"C9",X"21",X"0C",
		X"31",X"11",X"90",X"0B",X"0E",X"08",X"CD",X"F1",X"09",X"C3",X"F7",X"05",X"21",X"0C",X"31",X"11",
		X"98",X"0B",X"0E",X"08",X"CD",X"F1",X"09",X"21",X"0C",X"2F",X"11",X"03",X"06",X"0E",X"09",X"C3",
		X"18",X"06",X"C9",X"06",X"00",X"0C",X"04",X"26",X"0E",X"15",X"04",X"11",X"CD",X"DE",X"05",X"C3",
		X"EE",X"04",X"21",X"00",X"21",X"C3",X"51",X"00",X"CD",X"F1",X"09",X"06",X"06",X"DF",X"05",X"C2",
		X"1D",X"06",X"C9",X"0E",X"15",X"C3",X"44",X"05",X"21",X"08",X"31",X"0E",X"0F",X"C3",X"44",X"05",
		X"3E",X"01",X"32",X"F5",X"20",X"C3",X"3F",X"08",X"97",X"32",X"F5",X"20",X"C3",X"53",X"05",X"C2",
		X"1E",X"05",X"3A",X"AD",X"20",X"A7",X"CA",X"38",X"06",X"C3",X"27",X"05",X"97",X"D3",X"05",X"D3",
		X"03",X"00",X"00",X"00",X"00",X"CD",X"20",X"0B",X"CD",X"40",X"0B",X"CD",X"48",X"0B",X"C9",X"22",
		X"D3",X"20",X"3A",X"CE",X"20",X"3C",X"32",X"CE",X"20",X"3E",X"01",X"32",X"CD",X"20",X"E1",X"C9",
		X"00",X"32",X"CE",X"22",X"32",X"CD",X"20",X"C3",X"12",X"06",X"3A",X"CD",X"20",X"A7",X"C2",X"87",
		X"06",X"3A",X"CE",X"20",X"C3",X"61",X"05",X"DB",X"03",X"E6",X"80",X"CA",X"6E",X"06",X"97",X"32",
		X"CD",X"20",X"C3",X"6E",X"06",X"EB",X"7E",X"E6",X"FC",X"77",X"C3",X"A5",X"18",X"BC",X"D2",X"B1",
		X"06",X"2F",X"3C",X"84",X"FE",X"02",X"C9",X"BD",X"D2",X"B5",X"06",X"2F",X"3C",X"85",X"FE",X"E0",
		X"C9",X"94",X"C3",X"A4",X"06",X"95",X"C3",X"AE",X"06",X"11",X"0C",X"01",X"21",X"C0",X"20",X"06",
		X"0C",X"EF",X"C3",X"C8",X"05",X"3D",X"32",X"EE",X"20",X"E6",X"01",X"A7",X"C0",X"C3",X"5C",X"19",
		X"CD",X"CB",X"09",X"C3",X"BB",X"04",X"3E",X"23",X"CD",X"8F",X"04",X"67",X"CD",X"8D",X"04",X"84",
		X"67",X"C3",X"B8",X"0A",X"0A",X"CD",X"CB",X"09",X"C3",X"3F",X"08",X"00",X"00",X"82",X"82",X"FF",
		X"00",X"00",X"81",X"81",X"FF",X"00",X"00",X"42",X"5A",X"FF",X"00",X"00",X"3C",X"24",X"FF",X"FF",
		X"60",X"07",X"70",X"07",X"80",X"07",X"90",X"07",X"A0",X"07",X"B0",X"07",X"C0",X"07",X"D0",X"07",
		X"40",X"80",X"04",X"04",X"FF",X"80",X"40",X"03",X"05",X"FF",X"00",X"80",X"00",X"02",X"FF",X"FF",
		X"20",X"40",X"02",X"02",X"FF",X"C0",X"A0",X"01",X"02",X"FF",X"00",X"40",X"00",X"01",X"FF",X"FF",
		X"10",X"20",X"01",X"01",X"FF",X"E0",X"50",X"00",X"01",X"FF",X"00",X"A0",X"00",X"00",X"FF",X"FF",
		X"88",X"90",X"00",X"00",X"FF",X"70",X"A8",X"00",X"00",X"FF",X"00",X"50",X"00",X"00",X"FF",X"FF",
		X"44",X"48",X"00",X"00",X"FF",X"38",X"54",X"00",X"00",X"FF",X"00",X"28",X"00",X"00",X"FF",X"FF",
		X"22",X"14",X"00",X"00",X"FF",X"36",X"1C",X"00",X"00",X"FF",X"1C",X"00",X"00",X"00",X"FF",X"FF",
		X"44",X"28",X"00",X"00",X"FF",X"6C",X"38",X"00",X"00",X"FF",X"38",X"00",X"00",X"00",X"FF",X"FF",
		X"88",X"50",X"00",X"00",X"FF",X"D8",X"70",X"00",X"00",X"FF",X"70",X"00",X"00",X"00",X"FF",X"FF",
		X"10",X"A0",X"01",X"00",X"FF",X"B0",X"E0",X"01",X"00",X"FF",X"E0",X"00",X"00",X"00",X"FF",X"FF",
		X"20",X"40",X"02",X"01",X"FF",X"60",X"C0",X"03",X"01",X"FF",X"C0",X"00",X"01",X"00",X"FF",X"FF",
		X"40",X"80",X"04",X"02",X"FF",X"C0",X"80",X"06",X"03",X"FF",X"80",X"00",X"03",X"00",X"FF",X"FF",
		X"80",X"00",X"08",X"05",X"FF",X"80",X"00",X"0D",X"07",X"FF",X"00",X"00",X"07",X"00",X"FF",X"FF",
		X"00",X"00",X"11",X"0A",X"FF",X"00",X"00",X"1B",X"0E",X"FF",X"00",X"00",X"0E",X"00",X"FF",X"FF",
		X"40",X"40",X"10",X"10",X"FF",X"20",X"20",X"10",X"10",X"FF",X"40",X"40",X"08",X"0B",X"FF",X"80",
		X"80",X"07",X"04",X"FF",X"FF",X"11",X"B9",X"1C",X"CD",X"AA",X"1D",X"C3",X"17",X"13",X"00",X"00",
		X"FE",X"3F",X"C2",X"F8",X"17",X"0E",X"04",X"21",X"0E",X"2F",X"11",X"70",X"0B",X"CD",X"B0",X"0A",
		X"0E",X"0F",X"21",X"08",X"31",X"C3",X"0D",X"09",X"06",X"01",X"DF",X"05",X"C2",X"1A",X"08",X"CD",
		X"28",X"0A",X"C2",X"18",X"08",X"26",X"00",X"3A",X"AD",X"20",X"6F",X"0E",X"01",X"CD",X"EB",X"0B",
		X"7D",X"32",X"AD",X"20",X"CD",X"26",X"0B",X"3A",X"AD",X"20",X"FE",X"99",X"D2",X"53",X"08",X"DB",
		X"01",X"0F",X"DA",X"53",X"08",X"0E",X"15",X"11",X"74",X"0B",X"21",X"05",X"31",X"CD",X"F1",X"09",
		X"C3",X"18",X"08",X"3A",X"AD",X"20",X"FE",X"02",X"DA",X"62",X"08",X"DB",X"01",X"E6",X"02",X"C2",
		X"6E",X"08",X"DB",X"01",X"E6",X"04",X"CA",X"08",X"09",X"3E",X"01",X"C3",X"7B",X"08",X"CD",X"16",
		X"09",X"DB",X"00",X"E6",X"03",X"3C",X"32",X"E1",X"20",X"3E",X"02",X"32",X"F1",X"20",X"CD",X"16",
		X"09",X"CD",X"26",X"0B",X"DB",X"00",X"E6",X"03",X"3C",X"32",X"E0",X"20",X"21",X"40",X"26",X"36",
		X"00",X"23",X"7C",X"FE",X"3F",X"C2",X"8F",X"08",X"0E",X"08",X"21",X"0C",X"31",X"11",X"90",X"0B",
		X"CD",X"F1",X"09",X"C3",X"BC",X"08",X"4D",X"44",X"E5",X"7D",X"C6",X"DD",X"6F",X"24",X"7E",X"B8",
		X"00",X"00",X"00",X"23",X"7E",X"B9",X"00",X"00",X"00",X"C3",X"B2",X"04",X"CD",X"AF",X"03",X"21",
		X"00",X"23",X"06",X"08",X"EF",X"21",X"40",X"23",X"06",X"08",X"EF",X"21",X"80",X"23",X"06",X"08",
		X"EF",X"21",X"C0",X"23",X"06",X"08",X"EF",X"06",X"09",X"DF",X"05",X"C2",X"D9",X"08",X"21",X"F6",
		X"22",X"06",X"05",X"EF",X"06",X"08",X"21",X"ED",X"22",X"EF",X"97",X"CD",X"00",X"1C",X"31",X"9F",
		X"20",X"2A",X"A5",X"20",X"EB",X"2A",X"A9",X"20",X"7D",X"B4",X"B3",X"B2",X"A7",X"C2",X"5C",X"01",
		X"21",X"4E",X"00",X"22",X"9F",X"20",X"FB",X"C9",X"D3",X"06",X"C3",X"37",X"08",X"11",X"2D",X"09",
		X"CD",X"F1",X"09",X"C3",X"18",X"08",X"3A",X"AD",X"20",X"3D",X"47",X"E6",X"0F",X"FE",X"0F",X"C2",
		X"28",X"09",X"78",X"E6",X"F0",X"F6",X"09",X"47",X"78",X"32",X"AD",X"20",X"C9",X"1B",X"26",X"0F",
		X"0B",X"00",X"18",X"04",X"11",X"26",X"01",X"14",X"13",X"13",X"0E",X"0D",X"E5",X"CD",X"A7",X"0B",
		X"E1",X"23",X"C9",X"0E",X"04",X"21",X"0E",X"29",X"11",X"6C",X"0B",X"CD",X"BB",X"09",X"0E",X"08",
		X"21",X"0D",X"2C",X"11",X"F6",X"0B",X"CD",X"BB",X"09",X"21",X"07",X"31",X"CD",X"F7",X"0C",X"DF",
		X"21",X"11",X"31",X"1E",X"20",X"00",X"CD",X"D2",X"0B",X"DF",X"00",X"00",X"21",X"13",X"31",X"0E",
		X"07",X"11",X"A0",X"0B",X"CD",X"BB",X"09",X"21",X"07",X"34",X"CD",X"F5",X"10",X"DF",X"21",X"11",
		X"34",X"1E",X"50",X"00",X"CD",X"D2",X"0B",X"DF",X"00",X"00",X"21",X"13",X"34",X"0E",X"07",X"11",
		X"A0",X"0B",X"CD",X"BB",X"09",X"21",X"07",X"37",X"CD",X"F5",X"07",X"DF",X"21",X"0F",X"37",X"11",
		X"00",X"01",X"CD",X"CE",X"0B",X"DF",X"00",X"00",X"21",X"13",X"37",X"0E",X"07",X"11",X"A0",X"0B",
		X"CD",X"BB",X"09",X"06",X"03",X"DF",X"05",X"C2",X"B5",X"09",X"C9",X"1A",X"D5",X"E5",X"CD",X"A7",
		X"0B",X"E1",X"D1",X"DF",X"13",X"23",X"0D",X"C2",X"BB",X"09",X"C9",X"CD",X"F3",X"1C",X"0E",X"1C",
		X"21",X"01",X"24",X"11",X"50",X"0B",X"CD",X"F1",X"09",X"CD",X"40",X"0B",X"CD",X"20",X"0B",X"CD",
		X"48",X"0B",X"0E",X"07",X"21",X"16",X"3F",X"11",X"89",X"0B",X"CD",X"F1",X"09",X"CD",X"26",X"0B",
		X"C9",X"1A",X"D5",X"E5",X"CD",X"A7",X"0B",X"E1",X"D1",X"23",X"13",X"0D",X"C2",X"F1",X"09",X"C9",
		X"1E",X"21",X"21",X"21",X"3F",X"21",X"21",X"21",X"1F",X"21",X"21",X"1F",X"21",X"21",X"21",X"1F",
		X"1E",X"21",X"01",X"01",X"01",X"01",X"21",X"1E",X"1F",X"21",X"21",X"21",X"21",X"21",X"21",X"1F",
		X"3F",X"01",X"01",X"1F",X"01",X"01",X"01",X"3F",X"DB",X"01",X"E6",X"81",X"FE",X"81",X"C9",X"01",
		X"1E",X"21",X"01",X"01",X"39",X"21",X"21",X"1E",X"21",X"21",X"21",X"3F",X"21",X"21",X"21",X"21",
		X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"CD",X"9C",X"01",X"57",X"84",X"3D",X"3D",X"67",
		X"3D",X"3D",X"5F",X"87",X"87",X"C3",X"FC",X"1D",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"3F",
		X"21",X"33",X"2D",X"21",X"21",X"21",X"21",X"21",X"21",X"23",X"25",X"29",X"31",X"21",X"21",X"21",
		X"1E",X"21",X"21",X"21",X"21",X"21",X"21",X"1E",X"1F",X"21",X"21",X"1F",X"01",X"01",X"01",X"01",
		X"00",X"00",X"04",X"04",X"04",X"1F",X"1F",X"1F",X"1F",X"21",X"21",X"1F",X"09",X"11",X"21",X"21",
		X"1E",X"21",X"01",X"1E",X"20",X"20",X"21",X"1E",X"1F",X"04",X"04",X"04",X"04",X"04",X"04",X"04",
		X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"1E",X"21",X"21",X"21",X"21",X"21",X"21",X"0A",X"04",
		X"CD",X"F1",X"09",X"CD",X"CE",X"09",X"C9",X"14",X"CD",X"EB",X"19",X"84",X"67",X"C3",X"48",X"0A",
		X"11",X"11",X"11",X"11",X"0A",X"04",X"04",X"04",X"32",X"E2",X"20",X"3E",X"20",X"D3",X"03",X"C9",
		X"1E",X"21",X"23",X"25",X"29",X"31",X"21",X"1E",X"08",X"08",X"0C",X"08",X"08",X"08",X"08",X"08",
		X"1E",X"21",X"21",X"20",X"1C",X"02",X"01",X"3F",X"1E",X"21",X"20",X"1C",X"10",X"20",X"21",X"1E",
		X"10",X"18",X"14",X"12",X"11",X"3F",X"10",X"10",X"3F",X"01",X"01",X"1F",X"20",X"20",X"21",X"1F",
		X"1E",X"21",X"01",X"1D",X"23",X"21",X"21",X"1E",X"3F",X"21",X"20",X"10",X"08",X"04",X"02",X"01",
		X"1E",X"21",X"21",X"1E",X"21",X"21",X"21",X"1E",X"1E",X"21",X"21",X"31",X"2E",X"20",X"21",X"1E",
		X"21",X"A1",X"20",X"C3",X"C6",X"0B",X"3A",X"AD",X"20",X"5F",X"21",X"1D",X"3F",X"C3",X"D2",X"0B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"23",X"7E",X"BB",X"00",X"00",X"00",X"E1",X"E9",
		X"21",X"A5",X"20",X"C3",X"C6",X"0B",X"00",X"00",X"21",X"A9",X"20",X"C3",X"C6",X"0B",X"00",X"00",
		X"26",X"12",X"02",X"0E",X"11",X"04",X"26",X"1B",X"26",X"26",X"26",X"11",X"04",X"02",X"0E",X"11",
		X"03",X"26",X"26",X"26",X"12",X"02",X"0E",X"11",X"04",X"26",X"1C",X"26",X"0F",X"0B",X"00",X"18",
		X"0F",X"14",X"12",X"07",X"1B",X"26",X"0E",X"11",X"26",X"1C",X"26",X"0F",X"0B",X"00",X"18",X"04",
		X"11",X"12",X"26",X"01",X"14",X"13",X"13",X"0E",X"0D",X"02",X"11",X"04",X"03",X"08",X"13",X"26",
		X"0F",X"0B",X"00",X"18",X"04",X"11",X"26",X"1B",X"0F",X"0B",X"00",X"18",X"04",X"11",X"26",X"1C",
		X"26",X"0F",X"0E",X"08",X"0D",X"13",X"12",X"11",X"00",X"0A",X"E5",X"26",X"00",X"6F",X"29",X"29",
		X"29",X"19",X"EB",X"E1",X"06",X"08",X"D3",X"06",X"C5",X"1A",X"77",X"13",X"01",X"20",X"00",X"09",
		X"C1",X"05",X"C2",X"B8",X"0B",X"C9",X"5E",X"23",X"56",X"23",X"7E",X"23",X"66",X"6F",X"7A",X"CD",
		X"D3",X"0B",X"7B",X"D5",X"F5",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"CD",X"E6",X"0B",X"F1",X"E6",
		X"0F",X"CD",X"E6",X"0B",X"D1",X"C9",X"C6",X"1A",X"C3",X"3C",X"09",X"AF",X"7D",X"81",X"27",X"6F",
		X"7C",X"88",X"00",X"27",X"67",X"C9",X"00",X"12",X"13",X"11",X"0E",X"0F",X"00",X"0B",X"F3",X"76",
		X"7A",X"1E",X"8A",X"1E",X"9A",X"1E",X"10",X"07",X"20",X"07",X"30",X"07",X"40",X"07",X"50",X"07",
		X"00",X"00",X"41",X"41",X"FF",X"80",X"80",X"40",X"40",X"FF",X"00",X"00",X"21",X"2D",X"FF",X"00",
		X"00",X"1E",X"12",X"FF",X"FF",X"80",X"80",X"20",X"20",X"FF",X"40",X"40",X"20",X"20",X"FF",X"80",
		X"80",X"10",X"16",X"FF",X"00",X"00",X"0F",X"09",X"FF",X"FF",X"20",X"20",X"08",X"08",X"FF",X"10",
		X"10",X"08",X"08",X"FF",X"20",X"A0",X"04",X"05",X"FF",X"C0",X"40",X"03",X"02",X"FF",X"FF",X"10",
		X"10",X"04",X"04",X"FF",X"08",X"08",X"04",X"04",X"FF",X"10",X"D0",X"02",X"02",X"FF",X"E0",X"20",
		X"01",X"01",X"FF",X"FF",X"08",X"08",X"02",X"02",X"FF",X"04",X"04",X"02",X"02",X"FF",X"08",X"68",
		X"01",X"01",X"FF",X"F0",X"90",X"00",X"00",X"FF",X"FF",X"04",X"04",X"01",X"01",X"FF",X"02",X"02",
		X"01",X"01",X"FF",X"84",X"B4",X"00",X"00",X"FF",X"78",X"48",X"00",X"00",X"FF",X"FF",X"44",X"22",
		X"00",X"00",X"FF",X"92",X"41",X"00",X"00",X"FF",X"AA",X"5A",X"00",X"00",X"FF",X"44",X"34",X"00",
		X"00",X"FF",X"FF",X"88",X"44",X"00",X"00",X"FF",X"24",X"82",X"01",X"00",X"FF",X"54",X"B4",X"01",
		X"00",X"FF",X"88",X"48",X"00",X"00",X"FF",X"FF",X"10",X"88",X"01",X"00",X"FF",X"48",X"04",X"02",
		X"01",X"FF",X"A8",X"68",X"02",X"01",X"FF",X"10",X"90",X"01",X"00",X"FF",X"FF",X"20",X"10",X"02",
		X"01",X"FF",X"90",X"08",X"04",X"02",X"FF",X"50",X"D0",X"05",X"02",X"FF",X"20",X"20",X"02",X"01",
		X"FF",X"FF",X"40",X"20",X"04",X"02",X"FF",X"20",X"10",X"09",X"04",X"FF",X"A0",X"A0",X"0A",X"05",
		X"FF",X"40",X"40",X"04",X"02",X"FF",X"FF",X"11",X"41",X"1E",X"CD",X"AA",X"1D",X"C3",X"FA",X"0D",
		X"B9",X"1C",X"C9",X"1C",X"D9",X"1C",X"11",X"1D",X"21",X"1D",X"31",X"1D",X"41",X"1D",X"31",X"1E",
		X"80",X"40",X"08",X"04",X"FF",X"40",X"20",X"12",X"08",X"FF",X"40",X"40",X"15",X"0B",X"FF",X"80",
		X"80",X"08",X"04",X"FF",X"FF",X"00",X"80",X"11",X"08",X"FF",X"80",X"40",X"24",X"10",X"FF",X"80",
		X"80",X"2A",X"16",X"FF",X"00",X"00",X"11",X"09",X"FF",X"FF",X"00",X"00",X"22",X"11",X"FF",X"00",
		X"80",X"49",X"20",X"FF",X"00",X"00",X"55",X"2D",X"FF",X"00",X"00",X"22",X"12",X"FF",X"FF",X"84",
		X"04",X"40",X"40",X"00",X"00",X"FF",X"7C",X"04",X"40",X"40",X"00",X"00",X"FF",X"20",X"04",X"40",
		X"40",X"00",X"00",X"FF",X"10",X"08",X"43",X"20",X"00",X"00",X"FF",X"08",X"10",X"45",X"10",X"00",
		X"00",X"FF",X"10",X"20",X"25",X"08",X"00",X"00",X"FF",X"20",X"C0",X"19",X"07",X"00",X"00",X"FF",
		X"C0",X"00",X"01",X"00",X"00",X"00",X"FF",X"FF",X"08",X"08",X"81",X"80",X"00",X"00",X"FF",X"F8",
		X"08",X"80",X"80",X"00",X"00",X"FF",X"40",X"08",X"80",X"80",X"00",X"00",X"FF",X"20",X"10",X"86",
		X"40",X"00",X"00",X"FF",X"10",X"20",X"8A",X"20",X"00",X"00",X"FF",X"20",X"40",X"92",X"10",X"00",
		X"00",X"FF",X"40",X"80",X"62",X"0F",X"00",X"00",X"FF",X"80",X"00",X"03",X"00",X"00",X"00",X"FF",
		X"FF",X"10",X"10",X"02",X"00",X"01",X"01",X"FF",X"F0",X"10",X"01",X"00",X"01",X"01",X"FF",X"80",
		X"10",X"00",X"00",X"01",X"01",X"FF",X"40",X"20",X"0C",X"80",X"01",X"00",X"FF",X"20",X"40",X"14",
		X"40",X"01",X"00",X"FF",X"40",X"80",X"24",X"20",X"01",X"00",X"FF",X"80",X"00",X"C4",X"1F",X"00",
		X"00",X"FF",X"00",X"00",X"07",X"00",X"00",X"00",X"FF",X"FF",X"21",X"0A",X"31",X"C3",X"F4",X"0E",
		X"8E",X"0C",X"A3",X"0C",X"B8",X"0C",X"CD",X"0C",X"E2",X"0C",X"10",X"0D",X"25",X"0D",X"3A",X"0D",
		X"20",X"20",X"04",X"00",X"02",X"02",X"FF",X"E0",X"20",X"03",X"00",X"02",X"02",X"FF",X"00",X"20",
		X"01",X"00",X"02",X"02",X"FF",X"80",X"40",X"18",X"00",X"02",X"01",X"FF",X"40",X"80",X"28",X"80",
		X"02",X"00",X"FF",X"80",X"00",X"48",X"41",X"02",X"00",X"FF",X"00",X"00",X"89",X"3E",X"01",X"00",
		X"FF",X"00",X"00",X"0E",X"00",X"00",X"00",X"FF",X"FF",X"40",X"40",X"08",X"00",X"04",X"04",X"FF",
		X"C0",X"40",X"07",X"00",X"04",X"04",X"FF",X"00",X"40",X"02",X"00",X"04",X"04",X"FF",X"00",X"80",
		X"31",X"00",X"04",X"02",X"FF",X"80",X"00",X"50",X"01",X"04",X"01",X"FF",X"00",X"00",X"91",X"82",
		X"04",X"00",X"FF",X"00",X"00",X"12",X"7C",X"03",X"00",X"FF",X"00",X"00",X"1C",X"00",X"00",X"00",
		X"FF",X"FF",X"80",X"80",X"10",X"00",X"08",X"08",X"FF",X"80",X"80",X"0F",X"00",X"08",X"08",X"FF",
		X"00",X"80",X"04",X"00",X"08",X"08",X"FF",X"00",X"00",X"62",X"01",X"08",X"04",X"FF",X"00",X"00",
		X"A1",X"02",X"08",X"02",X"FF",X"00",X"00",X"22",X"04",X"09",X"01",X"FF",X"00",X"00",X"24",X"F8",
		X"06",X"00",X"FF",X"00",X"00",X"38",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"21",X"01",X"10",
		X"10",X"FF",X"00",X"00",X"1F",X"01",X"10",X"10",X"FF",X"00",X"00",X"08",X"01",X"10",X"10",X"FF",
		X"00",X"00",X"C4",X"02",X"10",X"08",X"FF",X"00",X"00",X"42",X"04",X"11",X"04",X"FF",X"00",X"00",
		X"44",X"08",X"12",X"02",X"FF",X"00",X"00",X"48",X"F0",X"0C",X"01",X"FF",X"00",X"00",X"70",X"00",
		X"00",X"00",X"FF",X"FF",X"11",X"A6",X"10",X"CD",X"AA",X"1D",X"21",X"0D",X"31",X"C3",X"F5",X"0F",
		X"EB",X"06",X"10",X"0C",X"25",X"0C",X"E0",X"07",X"3A",X"0C",X"4F",X"0C",X"64",X"0C",X"79",X"0C",
		X"00",X"00",X"01",X"02",X"10",X"10",X"FF",X"80",X"00",X"00",X"02",X"10",X"10",X"FF",X"00",X"00",
		X"01",X"02",X"08",X"10",X"FF",X"00",X"00",X"02",X"01",X"04",X"10",X"FF",X"00",X"00",X"04",X"62",
		X"02",X"08",X"FF",X"00",X"00",X"F8",X"94",X"01",X"04",X"FF",X"00",X"00",X"00",X"08",X"00",X"03",
		X"FF",X"FF",X"80",X"00",X"00",X"01",X"08",X"08",X"FF",X"40",X"00",X"00",X"01",X"08",X"08",X"FF",
		X"80",X"00",X"00",X"01",X"04",X"08",X"FF",X"00",X"80",X"01",X"00",X"02",X"08",X"FF",X"00",X"00",
		X"02",X"31",X"01",X"04",X"FF",X"00",X"00",X"FC",X"4A",X"00",X"02",X"FF",X"00",X"00",X"00",X"84",
		X"00",X"01",X"FF",X"FF",X"40",X"80",X"00",X"00",X"04",X"04",X"FF",X"20",X"80",X"00",X"00",X"04",
		X"04",X"FF",X"40",X"80",X"00",X"00",X"02",X"04",X"FF",X"80",X"40",X"00",X"00",X"01",X"04",X"FF",
		X"00",X"80",X"81",X"18",X"00",X"02",X"FF",X"00",X"00",X"7E",X"25",X"00",X"01",X"FF",X"00",X"00",
		X"00",X"C2",X"00",X"00",X"FF",X"FF",X"20",X"40",X"00",X"00",X"02",X"02",X"FF",X"10",X"40",X"00",
		X"00",X"02",X"02",X"FF",X"20",X"40",X"00",X"00",X"01",X"02",X"FF",X"40",X"20",X"80",X"00",X"00",
		X"02",X"FF",X"80",X"40",X"40",X"0C",X"00",X"01",X"FF",X"00",X"80",X"3F",X"92",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"61",X"00",X"00",X"FF",X"FF",X"00",X"00",X"01",X"0E",X"08",X"07",X"FF",X"80",
		X"00",X"BF",X"90",X"1F",X"00",X"FF",X"00",X"00",X"01",X"F0",X"08",X"00",X"FF",X"00",X"00",X"FE",
		X"00",X"07",X"00",X"FF",X"FF",X"11",X"10",X"11",X"CD",X"AA",X"1D",X"C9",X"00",X"00",X"00",X"00",
		X"11",X"1C",X"26",X"1C",X"3B",X"1C",X"50",X"1C",X"65",X"1C",X"7A",X"1C",X"8F",X"1C",X"A4",X"1C",
		X"10",X"20",X"00",X"00",X"01",X"01",X"FF",X"08",X"20",X"00",X"00",X"01",X"01",X"FF",X"10",X"20",
		X"80",X"00",X"00",X"01",X"FF",X"20",X"10",X"40",X"00",X"00",X"01",X"FF",X"40",X"20",X"20",X"86",
		X"00",X"00",X"FF",X"80",X"40",X"1F",X"49",X"00",X"00",X"FF",X"00",X"80",X"00",X"30",X"00",X"00",
		X"FF",X"FF",X"08",X"10",X"80",X"80",X"00",X"00",X"FF",X"04",X"10",X"80",X"80",X"00",X"00",X"FF",
		X"08",X"10",X"40",X"80",X"00",X"00",X"FF",X"10",X"08",X"20",X"80",X"00",X"00",X"FF",X"20",X"10",
		X"10",X"43",X"00",X"00",X"FF",X"C0",X"A0",X"0F",X"24",X"00",X"00",X"FF",X"00",X"40",X"00",X"18",
		X"00",X"00",X"FF",X"FF",X"04",X"08",X"40",X"40",X"00",X"00",X"FF",X"02",X"08",X"40",X"40",X"00",
		X"00",X"FF",X"04",X"08",X"20",X"40",X"00",X"00",X"FF",X"08",X"04",X"10",X"40",X"00",X"00",X"FF",
		X"10",X"88",X"08",X"21",X"00",X"00",X"FF",X"E0",X"50",X"07",X"12",X"00",X"00",X"FF",X"00",X"20",
		X"00",X"0C",X"00",X"00",X"FF",X"FF",X"02",X"04",X"20",X"20",X"00",X"00",X"FF",X"01",X"04",X"20",
		X"20",X"00",X"00",X"FF",X"02",X"04",X"10",X"20",X"00",X"00",X"FF",X"04",X"02",X"08",X"20",X"00",
		X"00",X"FF",X"08",X"C4",X"04",X"10",X"00",X"00",X"FF",X"F0",X"28",X"03",X"09",X"00",X"00",X"FF",
		X"00",X"10",X"00",X"06",X"00",X"00",X"FF",X"FF",X"80",X"00",X"00",X"87",X"04",X"03",X"FF",X"C0",
		X"00",X"DF",X"48",X"0F",X"00",X"FF",X"80",X"00",X"00",X"78",X"04",X"00",X"FF",X"00",X"00",X"DF",
		X"00",X"03",X"00",X"FF",X"FF",X"11",X"11",X"1C",X"CD",X"AA",X"1D",X"C3",X"F6",X"11",X"00",X"00",
		X"10",X"11",X"42",X"11",X"74",X"11",X"A6",X"12",X"A6",X"11",X"10",X"12",X"42",X"12",X"74",X"12",
		X"04",X"08",X"04",X"08",X"00",X"00",X"FF",X"02",X"04",X"08",X"10",X"00",X"00",X"FF",X"42",X"04",
		X"10",X"10",X"00",X"00",X"FF",X"A2",X"44",X"10",X"10",X"00",X"00",X"FF",X"14",X"A8",X"11",X"08",
		X"00",X"00",X"FF",X"08",X"10",X"0A",X"05",X"00",X"00",X"FF",X"00",X"00",X"04",X"02",X"00",X"00",
		X"FF",X"FF",X"08",X"10",X"08",X"10",X"00",X"00",X"FF",X"04",X"08",X"10",X"20",X"00",X"00",X"FF",
		X"84",X"08",X"20",X"20",X"00",X"00",X"FF",X"44",X"88",X"21",X"20",X"00",X"00",X"FF",X"28",X"50",
		X"22",X"11",X"00",X"00",X"FF",X"10",X"20",X"14",X"0A",X"00",X"00",X"FF",X"00",X"00",X"08",X"04",
		X"00",X"00",X"FF",X"FF",X"10",X"20",X"10",X"20",X"00",X"00",X"FF",X"08",X"10",X"20",X"40",X"00",
		X"00",X"FF",X"08",X"10",X"41",X"40",X"00",X"00",X"FF",X"88",X"10",X"42",X"41",X"00",X"00",X"FF",
		X"50",X"A0",X"44",X"22",X"00",X"00",X"FF",X"20",X"40",X"28",X"14",X"00",X"00",X"FF",X"00",X"00",
		X"10",X"08",X"00",X"00",X"FF",X"FF",X"40",X"80",X"40",X"80",X"00",X"00",X"FF",X"20",X"40",X"80",
		X"00",X"00",X"01",X"FF",X"20",X"40",X"04",X"00",X"01",X"01",X"FF",X"20",X"40",X"0A",X"04",X"01",
		X"01",X"FF",X"40",X"80",X"11",X"8A",X"01",X"00",X"FF",X"80",X"00",X"A0",X"51",X"00",X"00",X"FF",
		X"00",X"00",X"40",X"20",X"00",X"00",X"FF",X"FF",X"00",X"00",X"02",X"1C",X"10",X"0E",X"FF",X"00",
		X"00",X"7F",X"20",X"3F",X"01",X"FF",X"00",X"00",X"02",X"E0",X"10",X"01",X"FF",X"00",X"00",X"FC",
		X"00",X"0F",X"00",X"FF",X"FF",X"00",X"21",X"0A",X"34",X"11",X"79",X"0C",X"C3",X"F5",X"12",X"00",
		X"10",X"0F",X"42",X"0F",X"74",X"0F",X"A6",X"0F",X"10",X"10",X"42",X"10",X"74",X"10",X"A6",X"10",
		X"80",X"00",X"80",X"01",X"00",X"01",X"FF",X"40",X"80",X"00",X"00",X"01",X"02",X"FF",X"40",X"80",
		X"08",X"00",X"02",X"02",X"FF",X"40",X"80",X"14",X"08",X"02",X"02",X"FF",X"80",X"00",X"22",X"15",
		X"02",X"01",X"FF",X"00",X"00",X"41",X"A2",X"01",X"00",X"FF",X"00",X"00",X"80",X"40",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"01",X"02",X"01",X"02",X"FF",X"80",X"00",X"00",X"01",X"02",X"04",X"FF",
		X"80",X"00",X"10",X"01",X"04",X"04",X"FF",X"80",X"00",X"28",X"11",X"04",X"04",X"FF",X"00",X"00",
		X"45",X"2A",X"04",X"02",X"FF",X"00",X"00",X"82",X"44",X"02",X"01",X"FF",X"00",X"00",X"00",X"80",
		X"01",X"00",X"FF",X"FF",X"00",X"00",X"02",X"04",X"02",X"04",X"FF",X"00",X"00",X"01",X"02",X"04",
		X"08",X"FF",X"00",X"00",X"21",X"02",X"08",X"08",X"FF",X"00",X"00",X"51",X"22",X"08",X"08",X"FF",
		X"00",X"00",X"8A",X"54",X"08",X"04",X"FF",X"00",X"00",X"04",X"88",X"05",X"02",X"FF",X"00",X"00",
		X"00",X"00",X"02",X"01",X"FF",X"FF",X"20",X"40",X"20",X"40",X"00",X"00",X"FF",X"10",X"20",X"40",
		X"80",X"00",X"00",X"FF",X"10",X"20",X"82",X"80",X"00",X"00",X"FF",X"10",X"20",X"85",X"82",X"00",
		X"00",X"FF",X"A0",X"40",X"88",X"45",X"00",X"00",X"FF",X"40",X"80",X"50",X"28",X"00",X"00",X"FF",
		X"00",X"00",X"20",X"10",X"00",X"00",X"FF",X"FF",X"40",X"80",X"00",X"C3",X"02",X"01",X"FF",X"E0",
		X"00",X"EF",X"24",X"07",X"00",X"FF",X"40",X"00",X"00",X"3C",X"02",X"00",X"FF",X"80",X"00",X"EF",
		X"00",X"01",X"00",X"FF",X"FF",X"CD",X"AA",X"1D",X"21",X"0D",X"34",X"C3",X"10",X"13",X"00",X"00",
		X"41",X"1E",X"4F",X"0D",X"88",X"0D",X"C1",X"0D",X"10",X"0E",X"49",X"0E",X"82",X"0E",X"BB",X"0E",
		X"11",X"8E",X"0C",X"CD",X"AA",X"1D",X"C9",X"21",X"0A",X"37",X"11",X"50",X"07",X"CD",X"AA",X"1D",
		X"21",X"0D",X"37",X"11",X"60",X"07",X"CD",X"AA",X"1D",X"C9",X"CD",X"EB",X"0B",X"3A",X"E2",X"20",
		X"C9",X"D3",X"03",X"05",X"05",X"05",X"78",X"C9",X"23",X"97",X"77",X"C3",X"67",X"19",X"CD",X"BC",
		X"00",X"FE",X"0C",X"DA",X"60",X"13",X"3A",X"FA",X"20",X"CD",X"72",X"19",X"78",X"77",X"3D",X"FE",
		X"0B",X"C2",X"56",X"13",X"3E",X"07",X"12",X"13",X"23",X"7B",X"32",X"FA",X"20",X"C3",X"41",X"1F",
		X"23",X"97",X"77",X"C3",X"3E",X"1F",X"21",X"01",X"3F",X"11",X"86",X"13",X"3A",X"E2",X"20",X"A7",
		X"CA",X"79",X"13",X"3A",X"E1",X"20",X"C3",X"DC",X"13",X"3A",X"E0",X"20",X"C3",X"DC",X"13",X"CD",
		X"F1",X"09",X"C1",X"D1",X"E1",X"C9",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"26",X"26",X"26",
		X"26",X"26",X"26",X"26",X"26",X"26",X"11",X"C7",X"13",X"2A",X"D3",X"20",X"2B",X"CD",X"58",X"1D",
		X"21",X"00",X"3F",X"0E",X"09",X"11",X"8D",X"13",X"CD",X"F1",X"09",X"C3",X"EC",X"03",X"E6",X"01",
		X"2A",X"D3",X"20",X"2B",X"11",X"C7",X"13",X"A7",X"CA",X"C1",X"13",X"CD",X"58",X"1D",X"C3",X"7D",
		X"16",X"CD",X"AA",X"1D",X"C3",X"7D",X"16",X"80",X"80",X"01",X"01",X"FF",X"50",X"50",X"0A",X"0A",
		X"FF",X"28",X"28",X"14",X"14",X"FF",X"04",X"04",X"20",X"20",X"FF",X"FF",X"A7",X"CA",X"82",X"13",
		X"3D",X"A7",X"CA",X"82",X"13",X"4F",X"C3",X"7F",X"13",X"3E",X"02",X"C3",X"71",X"1F",X"CA",X"E2",
		X"18",X"FE",X"02",X"C2",X"57",X"18",X"3A",X"F5",X"20",X"A7",X"CA",X"E2",X"18",X"C3",X"33",X"04",
		X"07",X"C0",X"01",X"00",X"07",X"C0",X"01",X"00",X"07",X"C0",X"01",X"00",X"00",X"00",X"00",X"00",
		X"07",X"00",X"04",X"00",X"0F",X"C0",X"00",X"80",X"03",X"80",X"00",X"00",X"00",X"80",X"00",X"40",
		X"07",X"C0",X"0F",X"80",X"03",X"E0",X"07",X"40",X"01",X"C0",X"02",X"20",X"00",X"80",X"00",X"10",
		X"07",X"00",X"0E",X"40",X"07",X"00",X"02",X"10",X"03",X"80",X"00",X"00",X"02",X"00",X"00",X"00",
		X"07",X"E0",X"07",X"00",X"07",X"00",X"07",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"00",X"07",X"00",X"0E",X"00",X"04",X"00",X"1C",X"80",X"00",X"00",X"04",X"20",X"00",X"00",
		X"1F",X"00",X"0F",X"80",X"0E",X"80",X"07",X"C0",X"04",X"40",X"03",X"80",X"00",X"20",X"01",X"00",
		X"08",X"00",X"0E",X"00",X"01",X"00",X"1F",X"80",X"00",X"00",X"07",X"00",X"00",X"80",X"01",X"00",
		X"01",X"00",X"07",X"C0",X"01",X"00",X"07",X"C0",X"01",X"00",X"07",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"40",X"01",X"C0",X"02",X"00",X"07",X"E0",X"00",X"00",X"03",X"80",X"04",X"00",X"02",X"00",
		X"01",X"F0",X"03",X"E0",X"02",X"E0",X"07",X"C0",X"04",X"40",X"03",X"80",X"08",X"00",X"01",X"00",
		X"01",X"C0",X"01",X"C0",X"04",X"E0",X"03",X"80",X"10",X"80",X"00",X"80",X"00",X"00",X"00",X"00",
		X"07",X"E0",X"00",X"E0",X"00",X"E0",X"00",X"E0",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"C0",X"01",X"C0",X"03",X"80",X"04",X"E0",X"00",X"80",X"10",X"80",X"00",X"00",X"00",X"00",
		X"03",X"E0",X"01",X"F0",X"07",X"C0",X"02",X"E0",X"03",X"80",X"04",X"40",X"01",X"00",X"08",X"00",
		X"01",X"C0",X"00",X"40",X"07",X"E0",X"02",X"00",X"03",X"80",X"00",X"00",X"02",X"00",X"04",X"00",
		X"3A",X"D0",X"20",X"5F",X"16",X"14",X"21",X"B0",X"20",X"1A",X"77",X"7D",X"FE",X"BF",X"C8",X"13",
		X"23",X"C3",X"09",X"15",X"C5",X"06",X"00",X"11",X"B1",X"20",X"B7",X"1A",X"17",X"12",X"4F",X"1B",
		X"1A",X"17",X"12",X"79",X"B0",X"47",X"7B",X"FE",X"BE",X"CA",X"32",X"15",X"13",X"13",X"13",X"C3",
		X"1A",X"15",X"78",X"C1",X"A7",X"C0",X"23",X"C3",X"CC",X"17",X"00",X"00",X"1A",X"B6",X"77",X"13",
		X"2B",X"1A",X"B6",X"77",X"13",X"23",X"1A",X"E5",X"60",X"69",X"B6",X"77",X"13",X"2B",X"1A",X"B6",
		X"77",X"23",X"13",X"44",X"4D",X"E1",X"C9",X"1A",X"2F",X"A6",X"77",X"E6",X"07",X"CA",X"65",X"15",
		X"3E",X"01",X"32",X"D6",X"20",X"13",X"2B",X"1A",X"2F",X"A6",X"77",X"E6",X"E0",X"CA",X"75",X"15",
		X"3E",X"01",X"32",X"D6",X"20",X"13",X"23",X"1A",X"2F",X"E5",X"60",X"69",X"A6",X"77",X"E6",X"07",
		X"CA",X"88",X"15",X"3E",X"01",X"32",X"D6",X"20",X"13",X"2B",X"1A",X"2F",X"A6",X"77",X"E6",X"E0",
		X"CA",X"19",X"02",X"C3",X"14",X"02",X"7D",X"D6",X"20",X"4F",X"7C",X"DE",X"00",X"47",X"CD",X"3C",
		X"15",X"CD",X"82",X"1D",X"CD",X"3C",X"15",X"CD",X"82",X"1D",X"CD",X"3C",X"15",X"CD",X"82",X"1D",
		X"CD",X"3C",X"15",X"C9",X"7D",X"D6",X"20",X"4F",X"7C",X"DE",X"00",X"47",X"CD",X"57",X"15",X"CD",
		X"82",X"1D",X"CD",X"57",X"15",X"CD",X"82",X"1D",X"CD",X"57",X"15",X"CD",X"82",X"1D",X"CD",X"57",
		X"15",X"C9",X"3A",X"F5",X"20",X"A7",X"C8",X"FE",X"01",X"E5",X"C3",X"31",X"02",X"00",X"3A",X"D2",
		X"20",X"3D",X"32",X"D2",X"20",X"A7",X"C2",X"AA",X"16",X"3A",X"D7",X"20",X"A7",X"C2",X"AA",X"16",
		X"3E",X"10",X"32",X"D2",X"20",X"DB",X"01",X"07",X"07",X"D2",X"96",X"16",X"3A",X"D0",X"20",X"D6",
		X"10",X"32",X"D0",X"20",X"3A",X"D1",X"20",X"3D",X"3D",X"E6",X"1F",X"32",X"D1",X"20",X"3E",X"01",
		X"32",X"D8",X"20",X"11",X"B0",X"20",X"2A",X"D3",X"20",X"E5",X"D5",X"CD",X"B4",X"15",X"CD",X"00",
		X"15",X"D1",X"E1",X"3A",X"D6",X"20",X"A7",X"00",X"00",X"00",X"CD",X"96",X"15",X"3A",X"DA",X"20",
		X"A7",X"C2",X"87",X"16",X"DB",X"01",X"E6",X"10",X"A7",X"C2",X"7D",X"16",X"3E",X"03",X"C3",X"66",
		X"03",X"97",X"32",X"05",X"20",X"3A",X"D1",X"20",X"5F",X"16",X"17",X"1A",X"32",X"02",X"20",X"13",
		X"1A",X"32",X"01",X"20",X"2A",X"D3",X"20",X"7C",X"32",X"03",X"20",X"7D",X"32",X"04",X"20",X"CD",
		X"88",X"17",X"26",X"20",X"3A",X"DF",X"20",X"F5",X"97",X"32",X"DF",X"20",X"3A",X"00",X"22",X"6F",
		X"CD",X"8D",X"18",X"F1",X"32",X"DF",X"20",X"CD",X"88",X"17",X"C3",X"5E",X"05",X"3A",X"CF",X"20",
		X"A7",X"C2",X"87",X"1B",X"C3",X"12",X"1B",X"DB",X"01",X"E6",X"10",X"A7",X"CA",X"7D",X"16",X"21",
		X"DA",X"20",X"35",X"C3",X"7D",X"16",X"07",X"D2",X"AA",X"16",X"3A",X"D0",X"20",X"C6",X"10",X"32",
		X"D0",X"20",X"3A",X"D1",X"20",X"3C",X"3C",X"C3",X"09",X"16",X"3A",X"DD",X"20",X"47",X"3A",X"D5",
		X"20",X"90",X"D2",X"96",X"1B",X"3E",X"50",X"32",X"D5",X"20",X"DB",X"01",X"E6",X"08",X"A7",X"CA",
		X"6F",X"17",X"3A",X"D8",X"20",X"A7",X"C2",X"6F",X"17",X"3A",X"DD",X"20",X"FE",X"50",X"D2",X"D5",
		X"16",X"3C",X"32",X"DD",X"20",X"11",X"B0",X"20",X"2A",X"D3",X"20",X"E5",X"CD",X"B4",X"15",X"00",
		X"C3",X"33",X"18",X"00",X"00",X"00",X"E1",X"3A",X"D9",X"20",X"5F",X"16",X"17",X"1A",X"4F",X"B7",
		X"17",X"13",X"1A",X"CE",X"00",X"B7",X"17",X"17",X"17",X"17",X"17",X"5F",X"9F",X"C3",X"F7",X"03",
		X"00",X"FF",X"FF",X"FD",X"FF",X"FE",X"FE",X"FE",X"FE",X"FF",X"FE",X"00",X"FF",X"00",X"FF",X"01",
		X"00",X"01",X"01",X"02",X"01",X"01",X"02",X"01",X"02",X"00",X"02",X"FF",X"01",X"FF",X"01",X"FE",
		X"57",X"7B",X"E6",X"E0",X"26",X"3E",X"79",X"FE",X"03",X"DA",X"49",X"17",X"2F",X"3C",X"4F",X"A7",
		X"CA",X"63",X"17",X"CD",X"9C",X"1B",X"3A",X"D7",X"20",X"3C",X"E6",X"07",X"32",X"D7",X"20",X"3E",
		X"01",X"32",X"D2",X"20",X"0D",X"79",X"C3",X"2F",X"17",X"A7",X"CA",X"63",X"17",X"CD",X"14",X"15",
		X"3A",X"D7",X"20",X"3C",X"E6",X"07",X"32",X"D7",X"20",X"3E",X"01",X"32",X"D2",X"20",X"0D",X"79",
		X"C3",X"49",X"17",X"22",X"D3",X"20",X"11",X"B0",X"20",X"CD",X"96",X"15",X"C3",X"7D",X"1B",X"3A",
		X"DD",X"20",X"FE",X"03",X"DA",X"7B",X"17",X"3D",X"C3",X"D2",X"16",X"3A",X"D7",X"20",X"A7",X"C2",
		X"D5",X"16",X"3A",X"D1",X"20",X"C3",X"73",X"1B",X"3A",X"00",X"22",X"47",X"3A",X"00",X"20",X"32",
		X"00",X"22",X"78",X"32",X"00",X"20",X"2A",X"EB",X"20",X"EB",X"2A",X"DB",X"20",X"22",X"EB",X"20",
		X"EB",X"22",X"DB",X"20",X"3A",X"EE",X"20",X"47",X"3A",X"AE",X"20",X"32",X"EE",X"20",X"78",X"32",
		X"AE",X"20",X"C9",X"79",X"A7",X"C2",X"B9",X"17",X"19",X"7C",X"FE",X"27",X"DA",X"24",X"17",X"FE",
		X"3E",X"DA",X"26",X"17",X"CA",X"26",X"17",X"26",X"27",X"C3",X"26",X"17",X"E5",X"21",X"B1",X"20",
		X"11",X"B0",X"20",X"1A",X"47",X"7E",X"12",X"70",X"13",X"13",X"23",X"23",X"7D",X"FE",X"C1",X"C2",
		X"D3",X"17",X"E1",X"C9",X"CD",X"28",X"0A",X"C2",X"F0",X"17",X"F1",X"E1",X"D1",X"C1",X"FB",X"C9",
		X"3E",X"01",X"32",X"F5",X"20",X"21",X"40",X"26",X"36",X"00",X"23",X"7C",X"C3",X"00",X"08",X"00",
		X"88",X"1A",X"6B",X"1A",X"4E",X"1A",X"31",X"1A",X"D8",X"12",X"D8",X"10",X"D8",X"0F",X"D8",X"11",
		X"81",X"E6",X"0F",X"4F",X"D1",X"1B",X"12",X"A7",X"C2",X"42",X"1B",X"3A",X"F4",X"20",X"85",X"00",
		X"6F",X"3A",X"F3",X"20",X"8C",X"67",X"3A",X"F4",X"20",X"3D",X"C3",X"ED",X"1B",X"D1",X"24",X"24",
		X"C3",X"D2",X"1F",X"CD",X"88",X"17",X"26",X"20",X"3A",X"DF",X"20",X"F5",X"97",X"32",X"DF",X"20",
		X"3A",X"00",X"22",X"6F",X"C3",X"05",X"1B",X"00",X"00",X"1B",X"7C",X"12",X"1B",X"7D",X"12",X"3A",
		X"DF",X"20",X"FE",X"01",X"C3",X"EE",X"13",X"CD",X"A5",X"1D",X"3A",X"EE",X"20",X"A7",X"C2",X"C5",
		X"06",X"3E",X"0C",X"32",X"EE",X"20",X"97",X"32",X"05",X"22",X"3A",X"ED",X"20",X"5F",X"16",X"19",
		X"1A",X"32",X"02",X"22",X"13",X"1A",X"32",X"01",X"22",X"FE",X"02",X"D2",X"1B",X"19",X"C3",X"54",
		X"19",X"FE",X"01",X"CA",X"68",X"1B",X"C3",X"49",X"18",X"00",X"6F",X"26",X"22",X"7E",X"2B",X"FE",
		X"0C",X"CA",X"7A",X"1F",X"5E",X"2B",X"7E",X"A7",X"CA",X"F9",X"1F",X"57",X"97",X"77",X"2B",X"4E",
		X"2B",X"46",X"C3",X"95",X"06",X"3A",X"DF",X"20",X"00",X"A7",X"C2",X"F8",X"18",X"09",X"7C",X"FE",
		X"27",X"DA",X"C3",X"18",X"FE",X"3E",X"DA",X"BB",X"18",X"26",X"27",X"7E",X"A7",X"C2",X"06",X"02",
		X"C3",X"98",X"04",X"26",X"3E",X"C3",X"BB",X"18",X"3E",X"01",X"32",X"DF",X"20",X"3A",X"EF",X"20",
		X"3C",X"32",X"EF",X"20",X"97",X"32",X"F3",X"20",X"3E",X"01",X"32",X"F4",X"20",X"3E",X"02",X"32",
		X"F0",X"20",X"3A",X"00",X"22",X"FE",X"05",X"CA",X"ED",X"18",X"CD",X"8A",X"18",X"97",X"32",X"F6",
		X"20",X"32",X"DF",X"20",X"C3",X"C2",X"04",X"C9",X"EB",X"2B",X"7D",X"C3",X"E0",X"1B",X"00",X"00",
		X"FF",X"FF",X"00",X"FF",X"00",X"01",X"01",X"01",X"01",X"00",X"01",X"FF",X"00",X"FF",X"FF",X"FE",
		X"7D",X"C6",X"20",X"6F",X"7C",X"CE",X"00",X"67",X"C3",X"49",X"18",X"79",X"32",X"04",X"22",X"78",
		X"32",X"03",X"22",X"C3",X"5C",X"19",X"2B",X"C3",X"94",X"18",X"22",X"EB",X"20",X"C3",X"C6",X"1B",
		X"97",X"32",X"DF",X"20",X"3A",X"EC",X"20",X"CD",X"9D",X"06",X"D2",X"10",X"1A",X"3A",X"EB",X"20",
		X"CD",X"A7",X"06",X"D2",X"10",X"1A",X"E6",X"1F",X"FE",X"03",X"DA",X"F0",X"19",X"00",X"C3",X"10",
		X"1A",X"C3",X"E6",X"1D",X"7D",X"32",X"04",X"22",X"7C",X"32",X"03",X"22",X"3A",X"00",X"22",X"CD",
		X"8A",X"18",X"C9",X"CA",X"D0",X"19",X"23",X"23",X"23",X"23",X"3A",X"F9",X"20",X"BD",X"C3",X"41",
		X"02",X"00",X"5F",X"16",X"21",X"7E",X"12",X"13",X"23",X"7E",X"12",X"13",X"23",X"7E",X"12",X"13",
		X"23",X"C9",X"CD",X"BC",X"00",X"FE",X"0D",X"DA",X"9D",X"19",X"3A",X"F9",X"20",X"CD",X"72",X"19",
		X"78",X"77",X"3D",X"12",X"13",X"23",X"7B",X"32",X"F9",X"20",X"C3",X"D9",X"1E",X"23",X"97",X"77",
		X"C3",X"D6",X"1E",X"CD",X"BC",X"00",X"FE",X"07",X"DA",X"CA",X"19",X"3A",X"F8",X"20",X"CD",X"72",
		X"19",X"78",X"FE",X"0B",X"C2",X"BE",X"19",X"36",X"07",X"3E",X"0C",X"C3",X"C0",X"19",X"77",X"3C",
		X"12",X"13",X"23",X"7B",X"32",X"F8",X"20",X"C3",X"17",X"1F",X"23",X"97",X"77",X"C3",X"14",X"1F",
		X"CD",X"BC",X"00",X"FE",X"0C",X"DA",X"38",X"13",X"3A",X"F7",X"20",X"CD",X"72",X"19",X"78",X"77",
		X"3C",X"12",X"13",X"23",X"7B",X"32",X"F7",X"20",X"C3",X"6A",X"19",X"3E",X"30",X"C3",X"8F",X"04",
		X"97",X"57",X"32",X"EB",X"20",X"32",X"EC",X"20",X"32",X"DB",X"20",X"32",X"DC",X"20",X"C9",X"00",
		X"A5",X"1A",X"B5",X"1A",X"C5",X"1A",X"D5",X"1A",X"E5",X"1A",X"F5",X"1A",X"00",X"1D",X"00",X"1F",
		X"3A",X"DC",X"20",X"CD",X"9D",X"06",X"D2",X"29",X"1A",X"3A",X"DB",X"20",X"CD",X"A7",X"06",X"D2",
		X"29",X"1A",X"E6",X"1F",X"FE",X"03",X"DA",X"F0",X"19",X"3A",X"FB",X"20",X"C3",X"E6",X"1D",X"00",
		X"00",X"20",X"C0",X"00",X"E1",X"01",X"00",X"FF",X"F0",X"00",X"FD",X"12",X"03",X"00",X"FF",X"20",
		X"00",X"00",X"1E",X"01",X"00",X"FF",X"C0",X"00",X"FD",X"00",X"00",X"00",X"FF",X"FF",X"10",X"E0",
		X"80",X"70",X"00",X"00",X"FF",X"F8",X"00",X"FE",X"09",X"01",X"00",X"FF",X"10",X"00",X"80",X"0F",
		X"00",X"00",X"FF",X"E0",X"00",X"7F",X"00",X"00",X"00",X"FF",X"FF",X"08",X"70",X"40",X"38",X"00",
		X"00",X"FF",X"FC",X"80",X"FE",X"04",X"00",X"00",X"FF",X"08",X"80",X"40",X"07",X"00",X"00",X"FF",
		X"F0",X"00",X"3F",X"00",X"00",X"00",X"FF",X"FF",X"04",X"38",X"20",X"1C",X"00",X"00",X"FF",X"FE",
		X"40",X"7F",X"02",X"00",X"00",X"FF",X"04",X"C0",X"20",X"03",X"00",X"00",X"FE",X"F8",X"00",X"1F",
		X"00",X"00",X"00",X"FF",X"FF",X"EF",X"42",X"00",X"00",X"FF",X"42",X"3C",X"00",X"00",X"FF",X"3C",
		X"00",X"00",X"00",X"FF",X"FF",X"FE",X"84",X"01",X"00",X"FF",X"84",X"78",X"00",X"00",X"FF",X"78",
		X"00",X"00",X"00",X"FF",X"FF",X"FC",X"08",X"03",X"01",X"FF",X"08",X"F0",X"01",X"00",X"FF",X"F0",
		X"00",X"00",X"00",X"FF",X"FF",X"F8",X"10",X"07",X"02",X"FF",X"10",X"E0",X"02",X"01",X"FF",X"E0",
		X"00",X"01",X"00",X"FF",X"FF",X"F0",X"20",X"0F",X"04",X"FF",X"20",X"C0",X"04",X"03",X"FF",X"C0",
		X"00",X"03",X"00",X"FF",X"FF",X"E0",X"40",X"1F",X"08",X"FF",X"40",X"80",X"08",X"07",X"FF",X"80",
		X"00",X"07",X"00",X"FF",X"FF",X"CD",X"8D",X"18",X"F1",X"32",X"DF",X"20",X"CD",X"88",X"17",X"C3",
		X"E6",X"16",X"3A",X"D1",X"20",X"A7",X"CA",X"C0",X"1B",X"FE",X"80",X"CA",X"C0",X"1B",X"C3",X"8E",
		X"1B",X"E5",X"24",X"7E",X"23",X"B6",X"23",X"B6",X"E1",X"A7",X"CA",X"10",X"19",X"FE",X"01",X"CA",
		X"10",X"19",X"7D",X"D6",X"20",X"6F",X"7C",X"DE",X"00",X"67",X"C3",X"49",X"18",X"EB",X"2B",X"C3",
		X"DD",X"1B",X"7D",X"E6",X"1F",X"FE",X"19",X"D2",X"49",X"18",X"FE",X"15",X"D2",X"5C",X"1B",X"FE",
		X"10",X"D2",X"49",X"18",X"FE",X"09",X"DA",X"21",X"1B",X"C3",X"49",X"18",X"E5",X"25",X"7E",X"23",
		X"B6",X"23",X"B6",X"E1",X"A7",X"C2",X"81",X"18",X"7D",X"D6",X"20",X"6F",X"7C",X"DE",X"00",X"67",
		X"C3",X"49",X"18",X"32",X"D9",X"20",X"97",X"32",X"D8",X"20",X"C3",X"2D",X"16",X"3A",X"D7",X"20",
		X"A7",X"CA",X"2D",X"16",X"C3",X"7D",X"16",X"3D",X"32",X"CF",X"20",X"C3",X"5E",X"05",X"3E",X"0F",
		X"32",X"CF",X"20",X"C3",X"5F",X"16",X"32",X"D5",X"20",X"C3",X"7D",X"1B",X"C5",X"06",X"00",X"11",
		X"B0",X"20",X"B7",X"1A",X"1F",X"12",X"4F",X"13",X"1A",X"1F",X"12",X"79",X"B0",X"47",X"7B",X"FE",
		X"BF",X"CA",X"B8",X"1B",X"13",X"C3",X"A2",X"1B",X"78",X"C1",X"A7",X"C0",X"2B",X"C3",X"CC",X"17",
		X"3E",X"08",X"C3",X"90",X"1B",X"00",X"3E",X"03",X"77",X"EB",X"23",X"23",X"23",X"23",X"7E",X"3C",
		X"23",X"70",X"23",X"71",X"23",X"72",X"23",X"73",X"23",X"77",X"7D",X"D6",X"0A",X"6F",X"00",X"00",
		X"A7",X"C2",X"26",X"19",X"3A",X"00",X"22",X"C6",X"05",X"32",X"00",X"22",X"C9",X"81",X"E6",X"0F",
		X"4F",X"12",X"3A",X"ED",X"20",X"3C",X"3C",X"E6",X"0F",X"32",X"ED",X"20",X"C3",X"21",X"1B",X"00",
		X"CD",X"C8",X"0A",X"CD",X"B2",X"05",X"CD",X"CB",X"09",X"C9",X"D3",X"02",X"D3",X"00",X"C3",X"A6",
		X"08",X"8F",X"81",X"00",X"00",X"FF",X"B4",X"81",X"00",X"00",X"FF",X"D2",X"42",X"00",X"00",X"FF",
		X"1C",X"3C",X"00",X"00",X"FF",X"FF",X"1E",X"02",X"01",X"01",X"FF",X"68",X"02",X"01",X"01",X"FF",
		X"A4",X"84",X"00",X"00",X"FF",X"38",X"78",X"00",X"00",X"FF",X"FF",X"3C",X"04",X"02",X"02",X"FF",
		X"D0",X"04",X"02",X"02",X"FF",X"48",X"08",X"03",X"01",X"FF",X"70",X"F0",X"00",X"00",X"FF",X"FF",
		X"78",X"08",X"04",X"04",X"FF",X"A0",X"08",X"05",X"04",X"FF",X"90",X"10",X"06",X"02",X"FF",X"E0",
		X"E0",X"00",X"01",X"FF",X"FF",X"F0",X"10",X"08",X"08",X"FF",X"40",X"10",X"0B",X"08",X"FF",X"20",
		X"20",X"0D",X"04",X"FF",X"C0",X"C0",X"01",X"03",X"FF",X"FF",X"E0",X"20",X"11",X"10",X"FF",X"80",
		X"20",X"16",X"10",X"FF",X"40",X"40",X"1A",X"08",X"FF",X"80",X"80",X"03",X"07",X"FF",X"FF",X"C0",
		X"40",X"23",X"20",X"FF",X"00",X"40",X"2D",X"20",X"FF",X"80",X"80",X"34",X"10",X"FF",X"00",X"00",
		X"07",X"0F",X"FF",X"FF",X"80",X"80",X"47",X"40",X"FF",X"00",X"80",X"5A",X"40",X"FF",X"00",X"00",
		X"69",X"21",X"FF",X"00",X"00",X"0E",X"1E",X"FF",X"FF",X"26",X"24",X"00",X"00",X"FF",X"2A",X"1C",
		X"00",X"00",X"FF",X"14",X"00",X"00",X"00",X"FF",X"FF",X"4C",X"48",X"00",X"00",X"FF",X"54",X"38",
		X"00",X"00",X"FF",X"28",X"00",X"00",X"00",X"FF",X"FF",X"98",X"90",X"00",X"00",X"FF",X"A8",X"70",
		X"00",X"00",X"FF",X"50",X"00",X"00",X"00",X"FF",X"FF",X"02",X"B6",X"D1",X"C3",X"66",X"1F",X"00",
		X"00",X"00",X"00",X"21",X"00",X"24",X"36",X"00",X"23",X"7C",X"FE",X"40",X"C2",X"F6",X"1C",X"C9",
		X"C0",X"80",X"3F",X"10",X"FF",X"80",X"00",X"10",X"0F",X"FF",X"00",X"00",X"0F",X"00",X"FF",X"FF",
		X"00",X"30",X"20",X"01",X"01",X"FF",X"50",X"E0",X"01",X"00",X"FF",X"A0",X"00",X"00",X"00",X"FF",
		X"FF",X"60",X"40",X"02",X"02",X"FF",X"A0",X"C0",X"02",X"01",X"FF",X"40",X"00",X"01",X"00",X"FF",
		X"FF",X"C0",X"80",X"04",X"04",X"FF",X"40",X"80",X"05",X"03",X"FF",X"80",X"00",X"02",X"00",X"FF",
		X"FF",X"80",X"00",X"09",X"09",X"FF",X"80",X"00",X"0A",X"07",X"FF",X"00",X"00",X"05",X"00",X"FF",
		X"FF",X"00",X"00",X"0A",X"5F",X"03",X"0A",X"57",X"7D",X"D6",X"20",X"4F",X"7C",X"DE",X"00",X"47",
		X"E5",X"C5",X"1A",X"2F",X"A6",X"77",X"13",X"D5",X"1A",X"2F",X"5F",X"0A",X"A3",X"C3",X"E9",X"1C",
		X"1A",X"FE",X"FF",X"C2",X"63",X"1D",X"C1",X"E1",X"CD",X"81",X"1D",X"FE",X"FF",X"C2",X"60",X"1D",
		X"C9",X"13",X"7D",X"C6",X"20",X"6F",X"7C",X"CE",X"00",X"67",X"79",X"D6",X"20",X"4F",X"78",X"DE",
		X"00",X"47",X"FE",X"27",X"DA",X"F0",X"1F",X"7C",X"FE",X"3F",X"DA",X"9F",X"1D",X"26",X"27",X"1A",
		X"C9",X"06",X"3E",X"1A",X"C9",X"0A",X"5F",X"03",X"0A",X"57",X"7D",X"D6",X"20",X"4F",X"7C",X"DE",
		X"00",X"47",X"E5",X"C5",X"1A",X"B6",X"77",X"13",X"D5",X"C3",X"2A",X"1E",X"02",X"D1",X"03",X"13",
		X"23",X"1A",X"FE",X"FF",X"C2",X"B5",X"1D",X"C1",X"E1",X"CD",X"81",X"1D",X"FE",X"FF",X"C2",X"B2",
		X"1D",X"C9",X"5E",X"23",X"56",X"23",X"4E",X"23",X"46",X"EB",X"C5",X"D5",X"E5",X"CD",X"53",X"1D",
		X"E1",X"D1",X"C1",X"C3",X"30",X"19",X"81",X"E6",X"0F",X"1B",X"12",X"4F",X"C2",X"02",X"1E",X"3A",
		X"FD",X"20",X"85",X"6F",X"3A",X"FC",X"20",X"8C",X"67",X"C3",X"02",X"1E",X"C6",X"3A",X"6F",X"C3",
		X"0A",X"1C",X"3A",X"FF",X"20",X"85",X"6F",X"3A",X"FE",X"20",X"8C",X"67",X"FE",X"27",X"DA",X"25",
		X"1E",X"FE",X"3E",X"DA",X"1B",X"1E",X"CA",X"1B",X"1E",X"26",X"27",X"1B",X"7C",X"12",X"1B",X"7D",
		X"12",X"CD",X"A5",X"1D",X"C9",X"26",X"3E",X"C3",X"1B",X"1E",X"1A",X"5F",X"0A",X"B3",X"C3",X"BC",
		X"1D",X"00",X"00",X"13",X"12",X"FF",X"00",X"00",X"15",X"0E",X"FF",X"00",X"00",X"0A",X"00",X"FF",
		X"FF",X"42",X"02",X"20",X"20",X"00",X"00",X"FF",X"3E",X"02",X"20",X"20",X"00",X"00",X"FF",X"10",
		X"02",X"20",X"20",X"00",X"00",X"FF",X"88",X"04",X"21",X"10",X"00",X"00",X"FF",X"84",X"08",X"22",
		X"08",X"00",X"00",X"FF",X"88",X"10",X"12",X"04",X"00",X"00",X"FF",X"90",X"E0",X"0C",X"03",X"00",
		X"00",X"FF",X"E0",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"22",X"24",X"FF",X"00",
		X"00",X"1C",X"2A",X"FF",X"00",X"00",X"00",X"14",X"FF",X"FF",X"00",X"00",X"11",X"12",X"FF",X"00",
		X"00",X"0E",X"15",X"FF",X"00",X"00",X"00",X"0A",X"FF",X"FF",X"80",X"00",X"08",X"09",X"FF",X"00",
		X"80",X"07",X"0A",X"FF",X"00",X"00",X"00",X"05",X"FF",X"FF",X"97",X"EB",X"E9",X"00",X"3E",X"02",
		X"32",X"FB",X"20",X"21",X"00",X"01",X"22",X"FC",X"20",X"21",X"FF",X"E0",X"22",X"FE",X"20",X"CD",
		X"7F",X"02",X"00",X"23",X"7E",X"A7",X"CA",X"D6",X"1E",X"00",X"2B",X"E5",X"CD",X"75",X"02",X"E1",
		X"7A",X"A7",X"CA",X"82",X"19",X"23",X"23",X"23",X"23",X"3A",X"F7",X"20",X"BD",X"C2",X"C2",X"1E",
		X"00",X"CD",X"92",X"1F",X"21",X"00",X"20",X"22",X"FE",X"20",X"CD",X"87",X"02",X"23",X"7E",X"A7",
		X"CA",X"14",X"1F",X"2B",X"E5",X"CD",X"6B",X"02",X"E1",X"7A",X"A7",X"C3",X"10",X"1F",X"00",X"00",
		X"80",X"00",X"7F",X"21",X"FF",X"00",X"00",X"21",X"1E",X"FF",X"00",X"00",X"1E",X"00",X"FF",X"FF",
		X"CA",X"A3",X"19",X"23",X"23",X"23",X"23",X"3A",X"FA",X"20",X"BD",X"C3",X"48",X"02",X"3E",X"02",
		X"32",X"FB",X"20",X"21",X"FF",X"FF",X"22",X"FC",X"20",X"CD",X"A2",X"05",X"23",X"7E",X"A7",X"CA",
		X"3E",X"1F",X"2B",X"E5",X"CD",X"61",X"02",X"E1",X"7A",X"A7",X"CA",X"3E",X"13",X"23",X"23",X"23",
		X"23",X"3A",X"F8",X"20",X"BD",X"C2",X"2C",X"1F",X"CD",X"92",X"1F",X"21",X"FF",X"E0",X"22",X"FE",
		X"20",X"CD",X"AA",X"05",X"23",X"7E",X"A7",X"CA",X"67",X"19",X"2B",X"E5",X"CD",X"57",X"02",X"E1",
		X"7A",X"A7",X"C3",X"63",X"19",X"00",X"A7",X"CA",X"74",X"1F",X"FE",X"03",X"CA",X"E9",X"13",X"3E",
		X"01",X"32",X"DF",X"20",X"03",X"13",X"23",X"C3",X"70",X"1D",X"5E",X"2B",X"56",X"97",X"BA",X"CA",
		X"8B",X"1F",X"12",X"77",X"C3",X"8B",X"1F",X"1E",X"AA",X"03",X"1C",X"2B",X"2B",X"2B",X"7D",X"C3",
		X"EA",X"1F",X"3A",X"F5",X"20",X"A7",X"C2",X"10",X"04",X"3A",X"F6",X"20",X"C3",X"06",X"04",X"3A",
		X"EF",X"20",X"FE",X"01",X"CA",X"B2",X"1F",X"FE",X"02",X"CA",X"B8",X"1F",X"21",X"C8",X"20",X"C3",
		X"BB",X"1F",X"21",X"C0",X"20",X"C3",X"BB",X"1F",X"21",X"C4",X"20",X"5E",X"23",X"56",X"23",X"4E",
		X"23",X"46",X"EB",X"C5",X"D5",X"E5",X"CD",X"53",X"1D",X"E1",X"D1",X"C1",X"7D",X"E6",X"1F",X"CA",
		X"2A",X"04",X"D5",X"54",X"5D",X"3A",X"F4",X"20",X"8B",X"5F",X"3A",X"F3",X"20",X"8A",X"57",X"1A",
		X"A7",X"C2",X"2D",X"18",X"3A",X"F0",X"20",X"C3",X"10",X"18",X"32",X"00",X"22",X"C3",X"DE",X"1B",
		X"79",X"FE",X"20",X"DA",X"A1",X"1D",X"C3",X"97",X"1D",X"2B",X"2B",X"2B",X"7D",X"C3",X"DE",X"1B");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
