library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity b1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of b1 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"20",X"A1",X"6F",X"20",X"B8",X"7B",X"2C",X"0F",X"0C",X"30",X"49",X"A9",X"01",X"8D",X"00",X"0C",
		X"8D",X"01",X"0C",X"20",X"A2",X"79",X"20",X"F8",X"7C",X"90",X"25",X"A0",X"01",X"20",X"75",X"77",
		X"F0",X"1E",X"A5",X"B5",X"30",X"04",X"C6",X"B5",X"D0",X"E1",X"A0",X"01",X"B9",X"0D",X"0C",X"10",
		X"0F",X"B9",X"05",X"0C",X"10",X"0A",X"88",X"10",X"F3",X"A0",X"00",X"2C",X"07",X"0C",X"30",X"07",
		X"98",X"29",X"01",X"A8",X"A9",X"01",X"2C",X"A9",X"00",X"99",X"08",X"0C",X"20",X"A1",X"7E",X"20",
		X"82",X"70",X"F0",X"AC",X"20",X"96",X"6F",X"20",X"B2",X"6F",X"20",X"26",X"70",X"20",X"85",X"70",
		X"2C",X"0F",X"0C",X"10",X"F5",X"60",X"20",X"96",X"6F",X"20",X"00",X"68",X"20",X"B2",X"6F",X"E6",
		X"C7",X"A5",X"CA",X"85",X"A4",X"58",X"A5",X"CB",X"F0",X"08",X"20",X"45",X"6C",X"20",X"13",X"6E",
		X"F0",X"09",X"20",X"45",X"6C",X"20",X"64",X"6E",X"20",X"23",X"6F",X"20",X"27",X"71",X"20",X"54",
		X"73",X"20",X"C9",X"6F",X"20",X"78",X"6C",X"A5",X"B8",X"D0",X"06",X"20",X"2A",X"71",X"A2",X"01",
		X"2C",X"A2",X"00",X"8E",X"0A",X"0C",X"A2",X"01",X"8E",X"0F",X"0C",X"A2",X"FF",X"86",X"5E",X"A5",
		X"8B",X"C5",X"2C",X"F0",X"FA",X"85",X"2C",X"C6",X"59",X"C6",X"5A",X"A2",X"00",X"A5",X"59",X"D0",
		X"03",X"8E",X"0D",X"0C",X"A5",X"5A",X"D0",X"03",X"8E",X"0C",X"0C",X"A5",X"5C",X"F0",X"0F",X"C6",
		X"5C",X"A5",X"5C",X"A2",X"01",X"29",X"08",X"D0",X"02",X"A2",X"00",X"8E",X"09",X"0C",X"A9",X"00",
		X"85",X"14",X"A2",X"0A",X"B5",X"3C",X"F0",X"37",X"E6",X"14",X"20",X"C4",X"73",X"B5",X"47",X"86",
		X"24",X"10",X"70",X"29",X"7F",X"D0",X"36",X"8A",X"0A",X"AA",X"A0",X"00",X"20",X"57",X"74",X"9D",
		X"60",X"02",X"20",X"55",X"74",X"9D",X"60",X"02",X"A0",X"20",X"20",X"56",X"74",X"9D",X"60",X"02",
		X"20",X"55",X"74",X"9D",X"60",X"02",X"A9",X"14",X"20",X"16",X"74",X"A6",X"24",X"F6",X"47",X"CA",
		X"CA",X"10",X"C1",X"4C",X"FC",X"6A",X"A9",X"18",X"AC",X"A9",X"1C",X"D0",X"EB",X"C9",X"09",X"F0",
		X"F5",X"C9",X"12",X"F0",X"F4",X"C9",X"1B",X"D0",X"E4",X"8A",X"0A",X"AA",X"A0",X"00",X"BD",X"60",
		X"02",X"91",X"28",X"E8",X"C8",X"BD",X"60",X"02",X"91",X"28",X"A0",X"20",X"E8",X"BD",X"60",X"02",
		X"91",X"28",X"E8",X"C8",X"BD",X"60",X"02",X"91",X"28",X"A6",X"24",X"A0",X"00",X"94",X"3C",X"94",
		X"47",X"F0",X"BC",X"D0",X"5E",X"38",X"B5",X"3B",X"E9",X"21",X"B0",X"02",X"D6",X"3C",X"95",X"3B",
		X"20",X"C6",X"73",X"20",X"64",X"74",X"A0",X"03",X"20",X"2C",X"74",X"9D",X"00",X"02",X"E8",X"88",
		X"10",X"F6",X"20",X"6E",X"74",X"C6",X"23",X"D0",X"ED",X"38",X"A5",X"28",X"E9",X"5F",X"B0",X"02",
		X"C6",X"29",X"85",X"28",X"A9",X"18",X"4C",X"18",X"69",X"A2",X"20",X"2C",X"A2",X"30",X"A0",X"04",
		X"84",X"23",X"A0",X"03",X"8A",X"91",X"28",X"AA",X"E8",X"88",X"10",X"F8",X"20",X"6E",X"74",X"C6",
		X"23",X"D0",X"EF",X"4C",X"1B",X"69",X"A0",X"00",X"20",X"FE",X"6C",X"A0",X"20",X"20",X"FE",X"6C",
		X"4C",X"59",X"69",X"C9",X"09",X"F0",X"D2",X"C9",X"12",X"F0",X"D1",X"C9",X"1B",X"F0",X"CA",X"C9",
		X"24",X"F0",X"07",X"C9",X"60",X"F0",X"DF",X"4C",X"1D",X"69",X"20",X"64",X"74",X"A0",X"03",X"BD",
		X"00",X"02",X"91",X"28",X"E8",X"88",X"10",X"F7",X"20",X"6E",X"74",X"C6",X"23",X"D0",X"EE",X"A6",
		X"24",X"B5",X"48",X"10",X"0E",X"29",X"40",X"F0",X"07",X"A9",X"EC",X"85",X"2E",X"20",X"05",X"74",
		X"4C",X"5B",X"69",X"18",X"B5",X"3B",X"69",X"21",X"90",X"02",X"F6",X"3C",X"95",X"3B",X"20",X"C6",
		X"73",X"B5",X"48",X"AA",X"24",X"B5",X"10",X"03",X"09",X"70",X"2C",X"09",X"60",X"A0",X"00",X"91",
		X"28",X"A0",X"20",X"18",X"69",X"01",X"91",X"28",X"E0",X"0A",X"D0",X"09",X"A9",X"80",X"20",X"34",
		X"76",X"A9",X"80",X"D0",X"03",X"BD",X"25",X"6C",X"20",X"34",X"76",X"C6",X"A5",X"E6",X"A7",X"20",
		X"76",X"6D",X"86",X"8E",X"4C",X"1B",X"69",X"20",X"0D",X"6D",X"A9",X"00",X"8D",X"0F",X"0C",X"A5",
		X"B8",X"D0",X"0E",X"A0",X"D9",X"A2",X"61",X"20",X"9A",X"73",X"A0",X"E0",X"A2",X"61",X"20",X"9A",
		X"73",X"20",X"94",X"70",X"A5",X"B8",X"F0",X"76",X"24",X"13",X"70",X"21",X"C6",X"A4",X"F0",X"1D",
		X"A5",X"A7",X"85",X"A6",X"C9",X"14",X"90",X"07",X"20",X"22",X"71",X"A9",X"00",X"85",X"90",X"A9",
		X"00",X"85",X"A5",X"A5",X"B4",X"F0",X"5F",X"20",X"57",X"6C",X"4C",X"A1",X"68",X"24",X"B5",X"10",
		X"14",X"A0",X"69",X"A2",X"61",X"20",X"9A",X"73",X"A0",X"E7",X"A2",X"61",X"20",X"9A",X"73",X"A0",
		X"EE",X"A2",X"61",X"D0",X"1D",X"A0",X"4A",X"A2",X"61",X"20",X"9A",X"73",X"A4",X"B5",X"F0",X"07",
		X"A0",X"3C",X"A2",X"61",X"20",X"9A",X"73",X"A0",X"D9",X"A2",X"61",X"20",X"9A",X"73",X"A0",X"E0",
		X"A2",X"61",X"20",X"9A",X"73",X"A9",X"80",X"A4",X"B5",X"F0",X"01",X"4A",X"05",X"B4",X"C9",X"C0",
		X"D0",X"12",X"A5",X"B5",X"D0",X"05",X"20",X"C9",X"6F",X"30",X"03",X"20",X"CC",X"6F",X"20",X"9A",
		X"70",X"4C",X"6C",X"68",X"85",X"B4",X"A2",X"00",X"A5",X"B5",X"D0",X"08",X"A2",X"7F",X"24",X"CD",
		X"10",X"02",X"A2",X"FF",X"86",X"B5",X"20",X"6E",X"6C",X"4C",X"A1",X"68",X"A5",X"53",X"05",X"54",
		X"F0",X"56",X"F8",X"18",X"A2",X"FD",X"B5",X"56",X"75",X"A3",X"95",X"A3",X"E8",X"D0",X"F7",X"D8",
		X"A9",X"00",X"85",X"53",X"85",X"54",X"A5",X"9F",X"30",X"09",X"A5",X"A1",X"C5",X"CC",X"90",X"03",
		X"20",X"94",X"6D",X"A2",X"03",X"CA",X"30",X"1B",X"B5",X"A0",X"D5",X"C3",X"90",X"15",X"F0",X"F5",
		X"B5",X"A0",X"95",X"C3",X"CA",X"10",X"F9",X"24",X"B5",X"10",X"05",X"20",X"FA",X"71",X"D0",X"03",
		X"20",X"E2",X"71",X"A2",X"02",X"A5",X"B5",X"F0",X"07",X"10",X"0A",X"20",X"EC",X"71",X"D0",X"08",
		X"20",X"DC",X"71",X"D0",X"03",X"20",X"D4",X"71",X"A5",X"14",X"D0",X"22",X"A5",X"13",X"F0",X"03",
		X"4C",X"47",X"6A",X"A5",X"A7",X"C9",X"14",X"90",X"15",X"20",X"0D",X"6D",X"A9",X"00",X"8D",X"0F",
		X"0C",X"20",X"22",X"71",X"A9",X"00",X"85",X"90",X"20",X"57",X"6C",X"4C",X"A1",X"68",X"A5",X"8D",
		X"C9",X"3C",X"90",X"0E",X"A9",X"00",X"85",X"8D",X"E6",X"8E",X"E6",X"8F",X"E6",X"91",X"D0",X"02",
		X"E6",X"92",X"A5",X"92",X"D0",X"17",X"A0",X"01",X"A5",X"91",X"C9",X"14",X"F0",X"0A",X"C9",X"28",
		X"F0",X"05",X"C9",X"3C",X"D0",X"07",X"C8",X"C8",X"84",X"26",X"20",X"53",X"71",X"A5",X"A6",X"C9",
		X"14",X"B0",X"0E",X"A5",X"A5",X"C5",X"99",X"B0",X"08",X"A5",X"8E",X"C5",X"9A",X"90",X"02",X"66",
		X"57",X"A5",X"13",X"D0",X"42",X"A0",X"04",X"A5",X"8B",X"29",X"20",X"F0",X"02",X"A0",X"00",X"84",
		X"2E",X"20",X"05",X"74",X"2C",X"0F",X"0C",X"30",X"03",X"4C",X"43",X"7D",X"A5",X"B8",X"F0",X"2B",
		X"A5",X"8B",X"29",X"10",X"F0",X"18",X"A5",X"B5",X"D0",X"06",X"A0",X"91",X"A2",X"60",X"D0",X"11",
		X"30",X"06",X"A0",X"97",X"A2",X"60",X"D0",X"09",X"A0",X"9D",X"A2",X"60",X"D0",X"03",X"20",X"2E",
		X"6C",X"20",X"9A",X"73",X"4C",X"AF",X"68",X"A5",X"B8",X"D0",X"F3",X"A0",X"D9",X"A2",X"61",X"20",
		X"9A",X"73",X"A0",X"E0",X"A2",X"61",X"20",X"9A",X"73",X"A5",X"C0",X"F0",X"E1",X"A9",X"00",X"8D",
		X"0F",X"0C",X"4C",X"6C",X"68",X"03",X"00",X"06",X"00",X"15",X"00",X"30",X"00",X"80",X"A5",X"B5",
		X"D0",X"06",X"A0",X"A3",X"A2",X"60",X"D0",X"0C",X"30",X"06",X"A0",X"A9",X"A2",X"60",X"D0",X"04",
		X"A0",X"AF",X"A2",X"60",X"60",X"20",X"06",X"70",X"20",X"EC",X"6D",X"4C",X"96",X"71",X"20",X"06",
		X"70",X"20",X"FF",X"6D",X"4C",X"B6",X"71",X"20",X"9A",X"70",X"A5",X"B5",X"F0",X"08",X"20",X"CC",
		X"6F",X"20",X"94",X"72",X"F0",X"62",X"20",X"C9",X"6F",X"20",X"8E",X"72",X"F0",X"0D",X"20",X"9A",
		X"70",X"A5",X"B5",X"D0",X"4D",X"20",X"94",X"72",X"20",X"CC",X"6F",X"20",X"B5",X"6F",X"A5",X"B5",
		X"D0",X"06",X"20",X"DC",X"6F",X"4C",X"8B",X"6C",X"20",X"DF",X"6F",X"A5",X"B8",X"F0",X"0D",X"20",
		X"45",X"6C",X"20",X"8B",X"6E",X"24",X"90",X"30",X"0A",X"20",X"85",X"6E",X"20",X"0E",X"73",X"A9",
		X"80",X"85",X"90",X"20",X"97",X"70",X"20",X"45",X"6C",X"20",X"EA",X"70",X"20",X"B1",X"6D",X"20",
		X"49",X"6D",X"20",X"E8",X"6E",X"20",X"E9",X"6F",X"A5",X"B5",X"D0",X"03",X"4C",X"B8",X"72",X"4C",
		X"BE",X"72",X"20",X"C9",X"6F",X"20",X"8E",X"72",X"24",X"B5",X"10",X"AF",X"20",X"B5",X"6F",X"20",
		X"DF",X"6F",X"20",X"4E",X"6C",X"20",X"C3",X"6E",X"24",X"90",X"30",X"0A",X"20",X"A4",X"6E",X"20",
		X"58",X"73",X"A9",X"80",X"85",X"90",X"20",X"97",X"70",X"20",X"4E",X"6C",X"20",X"EA",X"70",X"20",
		X"A2",X"6D",X"20",X"40",X"6D",X"20",X"E3",X"6E",X"20",X"EF",X"6F",X"4C",X"BE",X"72",X"B1",X"28",
		X"C9",X"11",X"90",X"04",X"C9",X"60",X"90",X"04",X"A9",X"00",X"91",X"28",X"60",X"A9",X"06",X"85",
		X"8A",X"24",X"13",X"70",X"07",X"A9",X"00",X"85",X"2E",X"20",X"05",X"74",X"20",X"2E",X"6C",X"20",
		X"9A",X"73",X"A5",X"8A",X"D0",X"FC",X"60",X"A2",X"09",X"A0",X"9E",X"86",X"29",X"84",X"28",X"A5",
		X"A7",X"60",X"A2",X"0B",X"A0",X"80",X"86",X"29",X"84",X"28",X"A9",X"14",X"38",X"E5",X"A7",X"60",
		X"20",X"32",X"6D",X"A2",X"FE",X"A0",X"FF",X"D0",X"07",X"20",X"27",X"6D",X"A2",X"CF",X"A0",X"CE",
		X"85",X"26",X"84",X"24",X"86",X"25",X"A2",X"0A",X"A0",X"00",X"C6",X"26",X"30",X"03",X"A5",X"25",
		X"2C",X"A5",X"24",X"91",X"28",X"C8",X"C0",X"02",X"90",X"F0",X"20",X"7A",X"74",X"CA",X"D0",X"E8",
		X"60",X"20",X"32",X"6D",X"10",X"0A",X"24",X"B5",X"30",X"F7",X"20",X"27",X"6D",X"38",X"E9",X"01",
		X"4A",X"A0",X"00",X"90",X"01",X"C8",X"AA",X"F0",X"06",X"20",X"7A",X"74",X"CA",X"D0",X"FA",X"A9",
		X"CF",X"91",X"28",X"60",X"A9",X"80",X"85",X"9F",X"A9",X"49",X"85",X"5C",X"E6",X"A4",X"24",X"B5",
		X"10",X"0F",X"A9",X"86",X"38",X"E5",X"A4",X"85",X"23",X"A0",X"60",X"A2",X"09",X"A9",X"48",X"D0",
		X"0B",X"A6",X"A4",X"CA",X"86",X"23",X"A0",X"7E",X"A2",X"0B",X"A9",X"4C",X"84",X"28",X"86",X"29",
		X"A2",X"05",X"86",X"24",X"85",X"25",X"A6",X"23",X"CA",X"30",X"10",X"A5",X"25",X"20",X"16",X"74",
		X"20",X"7A",X"74",X"20",X"7A",X"74",X"C6",X"24",X"D0",X"EE",X"60",X"A9",X"00",X"A8",X"91",X"28",
		X"C8",X"91",X"28",X"A0",X"20",X"91",X"28",X"C8",X"91",X"28",X"D0",X"E4",X"A2",X"60",X"A0",X"B5",
		X"20",X"9A",X"73",X"A5",X"C9",X"D0",X"01",X"60",X"A2",X"60",X"A0",X"97",X"4C",X"9A",X"73",X"A2",
		X"60",X"A0",X"CE",X"D0",X"F7",X"80",X"61",X"8A",X"61",X"A0",X"61",X"B1",X"61",X"B6",X"61",X"CA",
		X"61",X"CF",X"61",X"A5",X"C0",X"D0",X"E0",X"A2",X"0C",X"86",X"5D",X"BC",X"05",X"6E",X"BD",X"06",
		X"6E",X"AA",X"20",X"9A",X"73",X"A6",X"5D",X"CA",X"CA",X"10",X"EE",X"20",X"03",X"6F",X"A0",X"00",
		X"84",X"2F",X"B9",X"25",X"6C",X"85",X"AB",X"A0",X"B5",X"A9",X"09",X"A2",X"0B",X"20",X"14",X"6F",
		X"A9",X"A0",X"8D",X"95",X"09",X"20",X"94",X"70",X"8D",X"D5",X"09",X"8D",X"B5",X"09",X"8D",X"95",
		X"09",X"20",X"A3",X"70",X"A4",X"2F",X"C8",X"C8",X"C0",X"0A",X"D0",X"D4",X"A9",X"AA",X"8D",X"B5",
		X"09",X"A9",X"00",X"60",X"A2",X"60",X"A0",X"FC",X"20",X"9A",X"73",X"A6",X"CC",X"30",X"10",X"A2",
		X"61",X"A0",X"10",X"20",X"9A",X"73",X"A0",X"72",X"A9",X"09",X"A2",X"2C",X"20",X"14",X"6F",X"A0",
		X"2B",X"A2",X"61",X"D0",X"1C",X"A0",X"42",X"A2",X"61",X"D0",X"1D",X"A2",X"61",X"A0",X"4A",X"20",
		X"9A",X"73",X"A5",X"B5",X"F0",X"07",X"A2",X"61",X"A0",X"3C",X"20",X"9A",X"73",X"A2",X"61",X"A0",
		X"57",X"4C",X"9A",X"73",X"A2",X"61",X"A0",X"61",X"20",X"D0",X"6E",X"A5",X"B5",X"30",X"06",X"A0",
		X"8E",X"A9",X"09",X"D0",X"5F",X"A0",X"51",X"A9",X"0A",X"84",X"2A",X"85",X"2B",X"A9",X"20",X"A0",
		X"00",X"F0",X"59",X"A2",X"61",X"A0",X"69",X"20",X"9A",X"73",X"A0",X"76",X"A2",X"61",X"D0",X"D1",
		X"20",X"9A",X"73",X"A5",X"B8",X"D0",X"03",X"A6",X"E3",X"2C",X"A6",X"A3",X"86",X"AA",X"A2",X"0A",
		X"4C",X"A4",X"7B",X"20",X"E8",X"73",X"D0",X"03",X"20",X"D5",X"73",X"20",X"D3",X"6E",X"A5",X"B5",
		X"10",X"06",X"A0",X"00",X"A9",X"0A",X"D0",X"C1",X"A0",X"DF",X"D0",X"B5",X"A2",X"60",X"A0",X"E7",
		X"4C",X"9A",X"73",X"A5",X"CB",X"F0",X"F5",X"A2",X"60",X"A0",X"F3",X"20",X"9A",X"73",X"A2",X"20",
		X"A0",X"7F",X"A9",X"0A",X"84",X"2A",X"85",X"2B",X"A9",X"E0",X"A0",X"20",X"85",X"25",X"A9",X"00",
		X"4C",X"16",X"72",X"20",X"03",X"6F",X"A9",X"FF",X"85",X"B8",X"A5",X"CB",X"D0",X"0D",X"20",X"73",
		X"77",X"D0",X"08",X"A2",X"03",X"20",X"A4",X"7B",X"20",X"E8",X"6E",X"A5",X"27",X"49",X"01",X"85",
		X"27",X"A6",X"C0",X"E0",X"01",X"F0",X"03",X"8D",X"01",X"0C",X"8D",X"00",X"0C",X"A0",X"10",X"20",
		X"B4",X"70",X"A6",X"C0",X"0E",X"0D",X"0C",X"6A",X"0E",X"0E",X"0C",X"6A",X"85",X"5F",X"24",X"5F",
		X"50",X"0A",X"10",X"05",X"88",X"D0",X"E8",X"F0",X"BA",X"E0",X"02",X"AD",X"E0",X"01",X"A5",X"CB",
		X"F0",X"02",X"90",X"F0",X"A0",X"00",X"70",X"02",X"A0",X"40",X"84",X"B4",X"84",X"C9",X"A5",X"CB",
		X"F0",X"08",X"50",X"03",X"20",X"AE",X"7B",X"20",X"AE",X"7B",X"A2",X"FF",X"86",X"B8",X"E8",X"8E",
		X"01",X"0C",X"8E",X"00",X"0C",X"60",X"A2",X"18",X"A9",X"00",X"9D",X"00",X"0C",X"CA",X"10",X"FA",
		X"60",X"A2",X"F0",X"A9",X"00",X"CA",X"95",X"10",X"8D",X"18",X"0C",X"D0",X"F8",X"F0",X"12",X"A2",
		X"00",X"2C",X"A2",X"C0",X"2C",X"A2",X"9F",X"A9",X"00",X"CA",X"95",X"00",X"8D",X"18",X"0C",X"D0",
		X"F8",X"8E",X"09",X"0C",X"E8",X"8E",X"0A",X"0C",X"60",X"A9",X"87",X"2C",X"A9",X"9F",X"85",X"23",
		X"A2",X"00",X"A9",X"90",X"A4",X"B8",X"F0",X"2D",X"A0",X"17",X"D0",X"1B",X"A9",X"D0",X"2C",X"A9",
		X"E8",X"A2",X"00",X"A0",X"47",X"84",X"23",X"D0",X"EB",X"A2",X"66",X"A9",X"23",X"D0",X"04",X"A2",
		X"66",X"A9",X"32",X"A0",X"0E",X"84",X"23",X"86",X"1F",X"85",X"1E",X"A6",X"23",X"B1",X"1E",X"95");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
