library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity sound is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of sound is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"B7",X"60",X"00",X"96",X"40",X"B7",X"30",X"00",X"81",X"11",X"26",X"F7",X"4F",X"8E",X"E0",X"00",
		X"B7",X"30",X"00",X"AB",X"80",X"8C",X"00",X"00",X"26",X"F6",X"81",X"00",X"27",X"02",X"86",X"01",
		X"B7",X"03",X"80",X"86",X"22",X"97",X"40",X"8E",X"00",X"00",X"CC",X"00",X"00",X"10",X"BE",X"30",
		X"00",X"ED",X"81",X"8C",X"03",X"00",X"25",X"F5",X"8E",X"E3",X"EF",X"CE",X"00",X"A0",X"EC",X"81",
		X"ED",X"C1",X"8C",X"E4",X"0F",X"25",X"F7",X"10",X"CE",X"04",X"00",X"1C",X"EF",X"B7",X"40",X"00",
		X"B7",X"20",X"07",X"20",X"FE",X"B7",X"60",X"00",X"B7",X"30",X"00",X"8E",X"00",X"80",X"CE",X"00",
		X"03",X"EC",X"81",X"ED",X"C1",X"EC",X"81",X"ED",X"C4",X"33",X"46",X"11",X"83",X"00",X"43",X"26",
		X"F0",X"8E",X"00",X"80",X"6F",X"80",X"8C",X"00",X"A0",X"26",X"F9",X"96",X"40",X"27",X"09",X"86",
		X"00",X"97",X"C0",X"BD",X"E2",X"33",X"20",X"02",X"0F",X"60",X"96",X"41",X"27",X"06",X"0F",X"41",
		X"0F",X"61",X"20",X"04",X"96",X"61",X"27",X"07",X"86",X"01",X"97",X"C0",X"BD",X"E2",X"33",X"96",
		X"42",X"27",X"09",X"86",X"02",X"97",X"C0",X"BD",X"E2",X"33",X"20",X"02",X"0F",X"62",X"96",X"43",
		X"27",X"09",X"86",X"03",X"97",X"C0",X"BD",X"E2",X"33",X"20",X"02",X"0F",X"63",X"96",X"44",X"27",
		X"09",X"86",X"04",X"97",X"C0",X"BD",X"E2",X"33",X"20",X"02",X"0F",X"64",X"96",X"45",X"27",X"09",
		X"86",X"05",X"97",X"C0",X"BD",X"E2",X"33",X"20",X"02",X"0F",X"65",X"96",X"46",X"27",X"09",X"86",
		X"06",X"97",X"C0",X"BD",X"E2",X"33",X"20",X"02",X"0F",X"66",X"96",X"47",X"27",X"06",X"0F",X"47",
		X"0F",X"67",X"20",X"04",X"96",X"67",X"27",X"07",X"86",X"07",X"97",X"C0",X"BD",X"E2",X"33",X"96",
		X"48",X"27",X"09",X"86",X"08",X"97",X"C0",X"BD",X"E2",X"33",X"20",X"02",X"0F",X"68",X"96",X"49",
		X"27",X"09",X"86",X"09",X"97",X"C0",X"BD",X"E2",X"33",X"20",X"02",X"0F",X"69",X"96",X"4A",X"27",
		X"06",X"0F",X"4A",X"0F",X"6A",X"20",X"04",X"96",X"6A",X"27",X"07",X"86",X"0A",X"97",X"C0",X"BD",
		X"E2",X"33",X"96",X"4B",X"27",X"06",X"0F",X"4B",X"0F",X"6B",X"20",X"04",X"96",X"6B",X"27",X"07",
		X"86",X"0B",X"97",X"C0",X"BD",X"E2",X"33",X"96",X"4C",X"27",X"06",X"0F",X"4C",X"0F",X"6C",X"20",
		X"04",X"96",X"6C",X"27",X"07",X"86",X"0C",X"97",X"C0",X"BD",X"E2",X"33",X"96",X"4D",X"27",X"06",
		X"0F",X"4D",X"0F",X"6D",X"20",X"04",X"96",X"6D",X"27",X"07",X"86",X"0D",X"97",X"C0",X"BD",X"E2",
		X"33",X"96",X"4E",X"27",X"06",X"0F",X"4E",X"0F",X"6E",X"20",X"04",X"96",X"6E",X"27",X"07",X"86",
		X"0E",X"97",X"C0",X"BD",X"E2",X"33",X"96",X"4F",X"27",X"09",X"86",X"0F",X"97",X"C0",X"BD",X"E2",
		X"33",X"20",X"02",X"0F",X"6F",X"96",X"50",X"27",X"09",X"86",X"10",X"97",X"C0",X"BD",X"E2",X"33",
		X"20",X"02",X"0F",X"70",X"96",X"51",X"27",X"09",X"86",X"11",X"97",X"C0",X"BD",X"E2",X"33",X"20",
		X"02",X"0F",X"71",X"96",X"52",X"27",X"09",X"86",X"12",X"97",X"C0",X"BD",X"E2",X"33",X"20",X"02",
		X"0F",X"72",X"96",X"53",X"27",X"09",X"86",X"13",X"97",X"C0",X"BD",X"E2",X"33",X"20",X"02",X"0F",
		X"73",X"96",X"54",X"27",X"09",X"86",X"14",X"97",X"C0",X"BD",X"E2",X"33",X"20",X"02",X"0F",X"74",
		X"96",X"55",X"27",X"09",X"86",X"15",X"97",X"C0",X"BD",X"E2",X"33",X"20",X"02",X"0F",X"75",X"96",
		X"56",X"27",X"09",X"86",X"16",X"97",X"C0",X"BD",X"E2",X"33",X"20",X"02",X"0F",X"76",X"96",X"57",
		X"27",X"09",X"86",X"17",X"97",X"C0",X"BD",X"E2",X"33",X"20",X"02",X"0F",X"77",X"96",X"58",X"27",
		X"09",X"86",X"18",X"97",X"C0",X"BD",X"E2",X"33",X"20",X"02",X"0F",X"78",X"96",X"59",X"27",X"09",
		X"86",X"19",X"97",X"C0",X"BD",X"E2",X"33",X"20",X"02",X"0F",X"79",X"86",X"01",X"97",X"C2",X"B7",
		X"40",X"00",X"3B",X"8E",X"E3",X"D5",X"D6",X"C0",X"A6",X"85",X"97",X"C1",X"8E",X"E4",X"09",X"58",
		X"AE",X"85",X"CE",X"00",X"60",X"54",X"A6",X"C5",X"26",X"35",X"6C",X"C5",X"CE",X"E4",X"3D",X"58",
		X"EE",X"C5",X"34",X"10",X"EC",X"C1",X"81",X"11",X"27",X"21",X"ED",X"84",X"10",X"AE",X"84",X"A6",
		X"C0",X"48",X"A7",X"02",X"EC",X"A1",X"ED",X"03",X"10",X"AF",X"84",X"BD",X"E3",X"09",X"30",X"0C",
		X"CC",X"00",X"00",X"ED",X"81",X"ED",X"81",X"A7",X"80",X"20",X"D9",X"A7",X"1F",X"35",X"10",X"A6",
		X"05",X"81",X"F0",X"27",X"55",X"CE",X"E5",X"D2",X"A6",X"04",X"48",X"EE",X"C6",X"E6",X"0A",X"A6",
		X"C5",X"81",X"10",X"25",X"45",X"33",X"C5",X"84",X"0F",X"10",X"8E",X"E2",X"9F",X"6E",X"B6",X"E2",
		X"CC",X"E2",X"D0",X"E2",X"C8",X"E2",X"A7",X"A6",X"0B",X"81",X"FF",X"27",X"14",X"E6",X"41",X"5C",
		X"D7",X"C3",X"91",X"C3",X"26",X"06",X"C6",X"FF",X"E7",X"0B",X"20",X"1E",X"4A",X"A7",X"0B",X"20",
		X"1B",X"A6",X"5F",X"4A",X"A7",X"0B",X"20",X"14",X"6F",X"0A",X"20",X"B9",X"A6",X"5F",X"20",X"0C",
		X"A6",X"5F",X"A1",X"09",X"23",X"06",X"A6",X"09",X"20",X"02",X"6C",X"0A",X"A7",X"05",X"CE",X"00",
		X"80",X"D6",X"C1",X"58",X"58",X"33",X"C5",X"EC",X"05",X"A7",X"C4",X"E7",X"43",X"EC",X"07",X"A7",
		X"42",X"E7",X"41",X"6A",X"09",X"26",X"02",X"8D",X"10",X"A6",X"88",X"10",X"81",X"11",X"26",X"01",
		X"39",X"0C",X"C1",X"30",X"88",X"11",X"7E",X"E2",X"7F",X"34",X"40",X"A6",X"94",X"81",X"F0",X"24",
		X"58",X"84",X"F0",X"81",X"C0",X"27",X"32",X"6F",X"05",X"CE",X"E6",X"D2",X"E6",X"02",X"EE",X"C5",
		X"44",X"44",X"44",X"97",X"C3",X"44",X"9B",X"C3",X"33",X"C6",X"EC",X"C4",X"ED",X"06",X"A6",X"42",
		X"A7",X"08",X"A6",X"94",X"84",X"0F",X"27",X"09",X"64",X"06",X"66",X"07",X"66",X"08",X"4A",X"26",
		X"F7",X"A6",X"03",X"AA",X"06",X"A7",X"06",X"20",X"04",X"86",X"F0",X"A7",X"05",X"EE",X"84",X"10",
		X"8E",X"00",X"A0",X"D6",X"C0",X"A6",X"A5",X"E6",X"41",X"3D",X"E7",X"09",X"33",X"42",X"EF",X"84",
		X"6F",X"0A",X"86",X"FF",X"A7",X"0B",X"35",X"40",X"39",X"EE",X"84",X"E6",X"41",X"10",X"8E",X"E3",
		X"76",X"84",X"0F",X"48",X"6E",X"B6",X"E3",X"BF",X"E3",X"8A",X"E3",X"8E",X"E3",X"98",X"E3",X"92",
		X"E3",X"AE",X"E3",X"A4",X"E3",X"86",X"EE",X"41",X"20",X"30",X"E7",X"03",X"20",X"06",X"E7",X"04",
		X"20",X"02",X"E7",X"0D",X"33",X"42",X"20",X"22",X"A6",X"0D",X"26",X"1C",X"6C",X"0C",X"E1",X"0C",
		X"27",X"16",X"20",X"10",X"6C",X"0F",X"E1",X"0F",X"26",X"0E",X"6F",X"0F",X"20",X"06",X"6C",X"0E",
		X"E1",X"0E",X"26",X"04",X"EE",X"42",X"20",X"02",X"33",X"44",X"EF",X"84",X"7E",X"E3",X"0B",X"8E",
		X"00",X"40",X"D6",X"C0",X"3A",X"C1",X"16",X"27",X"04",X"6F",X"84",X"20",X"02",X"6A",X"84",X"6F",
		X"88",X"20",X"35",X"50",X"39",X"00",X"00",X"01",X"00",X"00",X"01",X"00",X"00",X"04",X"04",X"04",
		X"05",X"05",X"05",X"04",X"02",X"02",X"02",X"01",X"02",X"00",X"00",X"00",X"00",X"03",X"04",X"02",
		X"01",X"01",X"03",X"01",X"02",X"07",X"01",X"05",X"02",X"03",X"02",X"01",X"01",X"01",X"01",X"04",
		X"05",X"05",X"01",X"03",X"06",X"02",X"01",X"04",X"01",X"01",X"00",X"02",X"21",X"01",X"00",X"01",
		X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"02",X"21",X"01",X"00",X"02",X"A9",X"02",X"A9",X"01",
		X"EE",X"01",X"DD",X"01",X"CC",X"01",X"AA",X"03",X"0F",X"02",X"ED",X"01",X"88",X"01",X"00",X"01",
		X"88",X"01",X"00",X"02",X"65",X"02",X"65",X"01",X"00",X"01",X"00",X"03",X"0F",X"E4",X"71",X"E4",
		X"8A",X"E4",X"97",X"E4",X"AA",X"E4",X"C0",X"E4",X"D6",X"E5",X"55",X"E5",X"B8",X"E4",X"F6",X"E5",
		X"03",X"E5",X"68",X"E5",X"3E",X"E5",X"2F",X"E5",X"33",X"E5",X"37",X"E5",X"48",X"E5",X"10",X"E5",
		X"17",X"E5",X"1E",X"E5",X"28",X"E5",X"75",X"E5",X"8E",X"E5",X"9B",X"E4",X"E9",X"E5",X"A8",X"E5",
		X"C5",X"E7",X"77",X"00",X"E7",X"D2",X"00",X"E8",X"5D",X"00",X"E8",X"C2",X"00",X"E8",X"FF",X"00",
		X"E9",X"3C",X"00",X"E9",X"42",X"00",X"E8",X"5D",X"01",X"11",X"E9",X"48",X"00",X"E9",X"6D",X"01",
		X"E9",X"90",X"02",X"E9",X"B5",X"02",X"11",X"E9",X"D8",X"00",X"E9",X"FD",X"00",X"EA",X"22",X"00",
		X"EA",X"47",X"00",X"EA",X"6A",X"00",X"EA",X"83",X"00",X"11",X"EA",X"9C",X"00",X"ED",X"98",X"01",
		X"EB",X"17",X"00",X"EB",X"A0",X"01",X"EB",X"A0",X"02",X"EC",X"A7",X"00",X"EB",X"17",X"02",X"11",
		X"ED",X"9E",X"00",X"ED",X"F7",X"00",X"EE",X"59",X"00",X"EE",X"F9",X"00",X"EF",X"B0",X"00",X"ED",
		X"9E",X"02",X"EE",X"59",X"02",X"11",X"F0",X"68",X"00",X"F0",X"7D",X"00",X"F0",X"92",X"00",X"F0",
		X"A9",X"00",X"F0",X"C0",X"00",X"F0",X"DF",X"00",X"11",X"E7",X"47",X"00",X"E7",X"4C",X"00",X"E7",
		X"47",X"01",X"E7",X"4C",X"01",X"11",X"E7",X"61",X"00",X"E7",X"6C",X"00",X"E7",X"61",X"01",X"E7",
		X"6C",X"01",X"11",X"F2",X"3C",X"00",X"F2",X"E1",X"01",X"F3",X"84",X"00",X"F3",X"8B",X"01",X"11",
		X"F3",X"92",X"00",X"F3",X"D3",X"01",X"11",X"F4",X"0E",X"00",X"F4",X"1B",X"01",X"11",X"F4",X"28",
		X"00",X"F4",X"37",X"00",X"F4",X"28",X"01",X"11",X"F4",X"46",X"00",X"F4",X"5F",X"01",X"11",X"F4",
		X"78",X"00",X"11",X"F7",X"75",X"00",X"11",X"F5",X"29",X"00",X"F5",X"E6",X"02",X"11",X"F8",X"4C",
		X"00",X"F8",X"4C",X"01",X"F8",X"4C",X"02",X"11",X"F8",X"69",X"00",X"F8",X"A2",X"00",X"F8",X"69",
		X"01",X"F8",X"A2",X"01",X"11",X"E7",X"51",X"00",X"E7",X"5C",X"00",X"E7",X"51",X"01",X"E7",X"5C",
		X"01",X"E7",X"51",X"02",X"E7",X"5C",X"02",X"11",X"F5",X"EE",X"00",X"F5",X"FB",X"00",X"F5",X"EE",
		X"01",X"F5",X"FB",X"01",X"11",X"F9",X"79",X"00",X"F9",X"9E",X"00",X"F9",X"A5",X"00",X"F9",X"FF",
		X"00",X"FA",X"0E",X"00",X"F9",X"79",X"01",X"F9",X"A5",X"01",X"F9",X"A5",X"02",X"11",X"F8",X"DB",
		X"00",X"F8",X"EA",X"00",X"F8",X"DB",X"01",X"F8",X"EA",X"01",X"11",X"F8",X"FB",X"00",X"F9",X"3A",
		X"00",X"F8",X"FB",X"02",X"F9",X"3A",X"02",X"11",X"F6",X"FC",X"00",X"F7",X"05",X"00",X"F7",X"0E",
		X"00",X"F7",X"33",X"00",X"F7",X"58",X"00",X"11",X"F6",X"08",X"00",X"F6",X"4F",X"01",X"F6",X"96",
		X"00",X"F6",X"C9",X"01",X"11",X"FA",X"1D",X"00",X"FA",X"1D",X"00",X"FA",X"1D",X"00",X"FA",X"1D",
		X"00",X"11",X"E6",X"10",X"E6",X"12",X"E6",X"14",X"E6",X"16",X"E6",X"18",X"E6",X"1A",X"E6",X"1C",
		X"E6",X"1E",X"E6",X"23",X"E6",X"28",X"E6",X"2D",X"E6",X"32",X"E6",X"37",X"E6",X"3C",X"E6",X"46",
		X"E6",X"4F",X"E6",X"54",X"E6",X"5C",X"E6",X"63",X"E6",X"6C",X"E6",X"6E",X"E6",X"70",X"E6",X"72",
		X"E6",X"85",X"E6",X"87",X"E6",X"94",X"E6",X"A2",X"E6",X"AB",X"E6",X"BA",X"E6",X"C6",X"E6",X"CA",
		X"0F",X"10",X"0C",X"10",X"0A",X"10",X"07",X"10",X"05",X"10",X"03",X"10",X"02",X"10",X"0A",X"0A",
		X"03",X"03",X"14",X"0F",X"0F",X"16",X"05",X"10",X"0C",X"0C",X"16",X"03",X"10",X"0C",X"0C",X"16",
		X"05",X"10",X"07",X"07",X"16",X"00",X"10",X"07",X"07",X"16",X"04",X"10",X"06",X"08",X"0A",X"0C",
		X"0F",X"0F",X"0F",X"16",X"05",X"10",X"04",X"06",X"08",X"0A",X"0A",X"0A",X"16",X"03",X"10",X"04",
		X"08",X"0A",X"0A",X"12",X"0F",X"0C",X"0A",X"08",X"05",X"03",X"00",X"10",X"0A",X"08",X"06",X"04",
		X"02",X"00",X"10",X"08",X"07",X"06",X"05",X"04",X"03",X"02",X"00",X"10",X"0F",X"12",X"0A",X"12",
		X"07",X"12",X"0F",X"0F",X"0F",X"06",X"06",X"06",X"0A",X"0A",X"0A",X"04",X"04",X"04",X"07",X"07",
		X"07",X"02",X"02",X"02",X"10",X"05",X"12",X"0A",X"0C",X"0F",X"0F",X"0F",X"0C",X"0A",X"07",X"05",
		X"03",X"01",X"00",X"10",X"08",X"09",X"0A",X"0B",X"0B",X"0B",X"0A",X"08",X"06",X"04",X"02",X"01",
		X"00",X"10",X"05",X"06",X"07",X"07",X"07",X"07",X"16",X"00",X"10",X"03",X"04",X"05",X"05",X"05",
		X"05",X"05",X"04",X"04",X"03",X"03",X"02",X"01",X"00",X"10",X"0F",X"0F",X"0F",X"0E",X"0C",X"0A",
		X"08",X"06",X"04",X"02",X"00",X"10",X"0A",X"16",X"00",X"10",X"0A",X"0C",X"0A",X"08",X"06",X"16",
		X"00",X"10",X"E6",X"D8",X"E6",X"FD",X"E7",X"22",X"02",X"54",X"A8",X"02",X"78",X"28",X"02",X"9D",
		X"B4",X"02",X"C5",X"78",X"02",X"EF",X"CB",X"03",X"1C",X"82",X"03",X"4B",X"C8",X"03",X"7D",X"F6",
		X"03",X"B3",X"35",X"03",X"EB",X"87",X"04",X"27",X"17",X"04",X"66",X"69",X"00",X"02",X"58",X"C0",
		X"02",X"7C",X"6C",X"02",X"A2",X"4F",X"02",X"CA",X"6B",X"02",X"F4",X"EA",X"03",X"21",X"F8",X"03",
		X"51",X"96",X"03",X"84",X"1A",X"03",X"B9",X"B1",X"03",X"F2",X"5B",X"04",X"2E",X"6E",X"04",X"6E",
		X"17",X"00",X"02",X"5C",X"D9",X"02",X"80",X"DC",X"02",X"A6",X"EB",X"02",X"CF",X"5E",X"02",X"FA",
		X"08",X"03",X"27",X"6E",X"03",X"57",X"63",X"03",X"8A",X"3F",X"03",X"C0",X"2E",X"03",X"F9",X"2E",
		X"04",X"35",X"C5",X"04",X"75",X"C5",X"00",X"10",X"07",X"32",X"04",X"F0",X"40",X"07",X"B3",X"04",
		X"F0",X"10",X"00",X"22",X"05",X"A3",X"05",X"F3",X"04",X"E7",X"53",X"F0",X"40",X"07",X"F7",X"E7",
		X"53",X"40",X"11",X"B3",X"01",X"02",X"01",X"B3",X"01",X"02",X"01",X"F0",X"40",X"11",X"83",X"01",
		X"93",X"01",X"83",X"01",X"93",X"01",X"F0",X"10",X"08",X"73",X"09",X"F2",X"10",X"53",X"03",X"F2",
		X"08",X"53",X"0C",X"C0",X"06",X"23",X"03",X"33",X"03",X"73",X"03",X"53",X"03",X"43",X"03",X"53",
		X"03",X"02",X"09",X"F2",X"10",X"A3",X"03",X"F2",X"08",X"A3",X"0C",X"C0",X"06",X"A3",X"03",X"02",
		X"03",X"32",X"03",X"22",X"03",X"02",X"03",X"A3",X"03",X"F1",X"40",X"F2",X"10",X"72",X"03",X"52",
		X"03",X"52",X"03",X"72",X"03",X"72",X"03",X"52",X"03",X"52",X"03",X"72",X"03",X"73",X"03",X"53",
		X"03",X"53",X"03",X"73",X"03",X"F2",X"00",X"74",X"04",X"54",X"04",X"74",X"04",X"F2",X"0D",X"94",
		X"30",X"F0",X"70",X"0B",X"A5",X"03",X"95",X"03",X"75",X"03",X"55",X"03",X"A5",X"03",X"95",X"03",
		X"75",X"03",X"55",X"03",X"A5",X"03",X"95",X"03",X"75",X"03",X"55",X"03",X"A5",X"03",X"95",X"03",
		X"75",X"03",X"55",X"03",X"64",X"03",X"54",X"03",X"34",X"03",X"14",X"03",X"64",X"03",X"54",X"03",
		X"34",X"03",X"14",X"03",X"64",X"03",X"54",X"03",X"34",X"03",X"14",X"03",X"64",X"03",X"54",X"03",
		X"34",X"03",X"24",X"03",X"A4",X"03",X"94",X"03",X"74",X"03",X"54",X"03",X"A4",X"03",X"94",X"03",
		X"74",X"03",X"54",X"03",X"A5",X"03",X"95",X"03",X"75",X"03",X"55",X"03",X"A5",X"03",X"95",X"03",
		X"75",X"03",X"55",X"03",X"F2",X"10",X"F1",X"40",X"91",X"03",X"61",X"03",X"21",X"03",X"92",X"03",
		X"21",X"03",X"92",X"03",X"62",X"03",X"22",X"03",X"F2",X"11",X"22",X"03",X"93",X"03",X"63",X"03",
		X"23",X"03",X"F2",X"12",X"23",X"03",X"94",X"03",X"64",X"03",X"24",X"03",X"F0",X"30",X"11",X"A4",
		X"06",X"54",X"02",X"54",X"02",X"54",X"02",X"A4",X"06",X"54",X"02",X"54",X"02",X"54",X"02",X"A4",
		X"06",X"54",X"02",X"54",X"02",X"54",X"02",X"A4",X"06",X"54",X"02",X"54",X"02",X"54",X"02",X"13",
		X"06",X"64",X"02",X"64",X"02",X"64",X"02",X"13",X"06",X"64",X"02",X"64",X"02",X"64",X"02",X"13",
		X"06",X"64",X"02",X"64",X"02",X"64",X"02",X"64",X"06",X"34",X"02",X"34",X"02",X"34",X"02",X"A4",
		X"06",X"54",X"02",X"54",X"02",X"54",X"02",X"A4",X"06",X"54",X"02",X"54",X"02",X"54",X"02",X"A4",
		X"06",X"54",X"02",X"54",X"02",X"54",X"02",X"A4",X"06",X"54",X"02",X"54",X"02",X"54",X"02",X"24",
		X"30",X"F0",X"30",X"0A",X"23",X"09",X"23",X"03",X"23",X"0C",X"C0",X"06",X"23",X"06",X"23",X"0C",
		X"63",X"09",X"63",X"03",X"63",X"0C",X"C0",X"06",X"63",X"06",X"A3",X"06",X"63",X"06",X"22",X"03",
		X"22",X"03",X"22",X"03",X"22",X"03",X"22",X"03",X"22",X"03",X"22",X"03",X"22",X"03",X"23",X"03",
		X"23",X"03",X"23",X"03",X"23",X"03",X"24",X"04",X"24",X"04",X"24",X"04",X"64",X"30",X"F0",X"10",
		X"0A",X"94",X"09",X"94",X"03",X"94",X"0C",X"C0",X"06",X"94",X"06",X"A4",X"0C",X"13",X"09",X"13",
		X"03",X"13",X"0C",X"C0",X"06",X"13",X"06",X"63",X"06",X"34",X"06",X"93",X"03",X"A3",X"03",X"A3",
		X"03",X"A3",X"03",X"93",X"03",X"A3",X"03",X"A3",X"03",X"A3",X"03",X"94",X"03",X"A4",X"03",X"A4",
		X"03",X"A4",X"03",X"A5",X"04",X"A5",X"04",X"A5",X"04",X"14",X"30",X"F0",X"20",X"08",X"F7",X"E7",
		X"79",X"F0",X"40",X"08",X"F7",X"E7",X"79",X"F0",X"20",X"00",X"42",X"01",X"32",X"01",X"42",X"01",
		X"C0",X"01",X"32",X"02",X"22",X"02",X"12",X"02",X"02",X"02",X"B3",X"02",X"F2",X"02",X"A3",X"01",
		X"83",X"01",X"63",X"01",X"F2",X"03",X"43",X"01",X"23",X"01",X"B4",X"01",X"F0",X"50",X"03",X"C0",
		X"02",X"43",X"01",X"33",X"01",X"43",X"01",X"F2",X"04",X"C0",X"01",X"33",X"02",X"23",X"02",X"13",
		X"02",X"03",X"01",X"B4",X"01",X"F2",X"05",X"A4",X"01",X"84",X"01",X"64",X"01",X"24",X"01",X"F0",
		X"10",X"00",X"02",X"01",X"B3",X"01",X"02",X"01",X"C0",X"01",X"B3",X"02",X"A3",X"02",X"93",X"02",
		X"83",X"01",X"73",X"01",X"F2",X"02",X"63",X"01",X"43",X"01",X"23",X"01",X"F2",X"03",X"03",X"01",
		X"A4",X"01",X"74",X"01",X"F0",X"40",X"03",X"C0",X"02",X"03",X"01",X"B4",X"01",X"03",X"01",X"F2",
		X"04",X"C0",X"01",X"B4",X"02",X"A4",X"02",X"94",X"02",X"84",X"01",X"74",X"01",X"F2",X"05",X"64",
		X"01",X"44",X"01",X"24",X"01",X"B5",X"01",X"F0",X"00",X"08",X"A5",X"06",X"04",X"06",X"A5",X"06",
		X"75",X"06",X"A5",X"06",X"34",X"06",X"54",X"06",X"74",X"06",X"A4",X"06",X"33",X"06",X"53",X"06",
		X"73",X"06",X"F2",X"11",X"B3",X"0C",X"93",X"06",X"F2",X"13",X"B3",X"36",X"F0",X"00",X"09",X"75",
		X"06",X"85",X"06",X"75",X"06",X"C0",X"06",X"75",X"06",X"A5",X"06",X"34",X"06",X"54",X"06",X"74",
		X"06",X"A4",X"06",X"33",X"06",X"53",X"06",X"F2",X"11",X"73",X"0C",X"63",X"06",X"F2",X"13",X"73",
		X"36",X"F0",X"40",X"1D",X"C0",X"02",X"A5",X"06",X"04",X"06",X"A5",X"06",X"C0",X"0A",X"75",X"06",
		X"A5",X"06",X"34",X"06",X"54",X"06",X"74",X"06",X"A4",X"06",X"33",X"06",X"F2",X"11",X"23",X"0C",
		X"23",X"06",X"F2",X"13",X"23",X"36",X"F0",X"40",X"0B",X"C0",X"02",X"75",X"06",X"85",X"06",X"75",
		X"06",X"C0",X"10",X"75",X"06",X"A5",X"06",X"34",X"06",X"54",X"06",X"74",X"06",X"A4",X"06",X"F2",
		X"11",X"B4",X"0C",X"94",X"06",X"F2",X"13",X"B4",X"36",X"F0",X"40",X"0B",X"C0",X"2A",X"75",X"06",
		X"A5",X"06",X"34",X"06",X"54",X"06",X"74",X"06",X"F2",X"11",X"74",X"0C",X"64",X"06",X"F2",X"13",
		X"74",X"36",X"F0",X"40",X"05",X"C0",X"30",X"75",X"06",X"A5",X"06",X"34",X"06",X"54",X"06",X"F1",
		X"20",X"F2",X"11",X"24",X"0C",X"24",X"06",X"F2",X"13",X"24",X"36",X"F0",X"20",X"08",X"73",X"04",
		X"A4",X"02",X"F2",X"13",X"73",X"0A",X"F2",X"08",X"73",X"02",X"53",X"02",X"13",X"02",X"53",X"02",
		X"73",X"04",X"A4",X"02",X"F2",X"13",X"73",X"0C",X"F2",X"08",X"93",X"02",X"A3",X"02",X"02",X"02",
		X"22",X"04",X"53",X"02",X"F2",X"13",X"22",X"0A",X"F2",X"08",X"22",X"02",X"02",X"02",X"83",X"02",
		X"02",X"02",X"22",X"04",X"53",X"02",X"F2",X"13",X"22",X"12",X"F2",X"08",X"52",X"04",X"02",X"02",
		X"52",X"0C",X"32",X"02",X"22",X"02",X"02",X"02",X"A3",X"04",X"73",X"02",X"F2",X"13",X"A3",X"12",
		X"F2",X"08",X"A3",X"04",X"63",X"02",X"F2",X"13",X"A3",X"12",X"F2",X"12",X"F1",X"40",X"C0",X"02",
		X"93",X"02",X"93",X"02",X"C0",X"02",X"73",X"02",X"73",X"02",X"53",X"02",X"73",X"02",X"93",X"02",
		X"53",X"02",X"73",X"02",X"83",X"02",X"F0",X"10",X"0E",X"33",X"04",X"74",X"02",X"F2",X"14",X"33",
		X"0A",X"F2",X"0E",X"33",X"02",X"84",X"02",X"84",X"01",X"84",X"01",X"84",X"01",X"84",X"01",X"33",
		X"04",X"74",X"02",X"F2",X"14",X"33",X"0C",X"F2",X"0E",X"63",X"02",X"63",X"01",X"63",X"01",X"63",
		X"01",X"63",X"01",X"53",X"04",X"23",X"02",X"F2",X"14",X"53",X"0A",X"F2",X"0E",X"53",X"02",X"33",
		X"02",X"33",X"01",X"33",X"01",X"33",X"01",X"33",X"01",X"53",X"04",X"23",X"02",X"F2",X"14",X"53",
		X"12",X"F2",X"0E",X"83",X"04",X"83",X"02",X"83",X"0C",X"73",X"02",X"53",X"02",X"33",X"02",X"73",
		X"04",X"23",X"02",X"F2",X"14",X"73",X"12",X"F2",X"13",X"63",X"04",X"13",X"02",X"F2",X"14",X"63",
		X"12",X"F1",X"40",X"F2",X"12",X"C0",X"02",X"53",X"02",X"53",X"02",X"C0",X"02",X"43",X"02",X"43",
		X"02",X"F2",X"03",X"03",X"02",X"43",X"02",X"53",X"02",X"03",X"02",X"33",X"02",X"53",X"02",X"F0",
		X"40",X"10",X"34",X"02",X"34",X"01",X"34",X"01",X"A5",X"01",X"A5",X"01",X"34",X"02",X"A5",X"02",
		X"34",X"02",X"A5",X"02",X"34",X"02",X"A5",X"02",X"14",X"02",X"14",X"01",X"14",X"01",X"14",X"01",
		X"14",X"01",X"34",X"02",X"34",X"01",X"34",X"01",X"A5",X"01",X"A5",X"01",X"34",X"02",X"A5",X"02",
		X"34",X"02",X"A5",X"02",X"34",X"02",X"A5",X"02",X"24",X"02",X"24",X"01",X"24",X"01",X"04",X"01",
		X"04",X"01",X"A5",X"02",X"A5",X"01",X"A5",X"01",X"54",X"01",X"54",X"01",X"A5",X"02",X"54",X"02",
		X"A5",X"02",X"54",X"02",X"A5",X"02",X"54",X"02",X"85",X"02",X"85",X"01",X"85",X"01",X"85",X"01",
		X"85",X"01",X"A5",X"02",X"A5",X"01",X"A5",X"01",X"54",X"01",X"54",X"01",X"A5",X"02",X"54",X"02",
		X"A5",X"02",X"54",X"02",X"A5",X"02",X"54",X"02",X"A5",X"02",X"A5",X"01",X"A5",X"01",X"24",X"01",
		X"24",X"01",X"54",X"02",X"54",X"01",X"54",X"01",X"04",X"01",X"04",X"01",X"F2",X"00",X"54",X"02",
		X"84",X"02",X"A4",X"02",X"03",X"02",X"84",X"02",X"04",X"02",X"54",X"06",X"F2",X"10",X"74",X"02",
		X"74",X"01",X"74",X"01",X"24",X"01",X"24",X"01",X"74",X"02",X"24",X"02",X"74",X"02",X"24",X"02",
		X"74",X"02",X"24",X"02",X"74",X"02",X"24",X"01",X"24",X"01",X"74",X"01",X"74",X"01",X"64",X"02",
		X"64",X"01",X"64",X"01",X"14",X"01",X"14",X"01",X"64",X"02",X"14",X"02",X"64",X"02",X"14",X"02",
		X"64",X"02",X"14",X"02",X"64",X"02",X"14",X"01",X"14",X"01",X"64",X"01",X"64",X"01",X"54",X"02",
		X"54",X"01",X"54",X"01",X"04",X"01",X"04",X"01",X"44",X"02",X"44",X"01",X"44",X"01",X"04",X"01",
		X"04",X"01",X"54",X"02",X"54",X"01",X"54",X"01",X"04",X"01",X"04",X"01",X"A5",X"02",X"A5",X"01",
		X"A5",X"01",X"24",X"01",X"24",X"01",X"F0",X"40",X"11",X"74",X"02",X"74",X"01",X"74",X"01",X"34",
		X"01",X"34",X"01",X"74",X"02",X"34",X"02",X"74",X"02",X"34",X"02",X"74",X"02",X"34",X"02",X"54",
		X"02",X"54",X"01",X"54",X"01",X"54",X"01",X"54",X"01",X"74",X"02",X"74",X"01",X"74",X"01",X"34",
		X"01",X"34",X"01",X"74",X"02",X"34",X"02",X"74",X"02",X"34",X"02",X"74",X"02",X"34",X"02",X"94",
		X"02",X"94",X"01",X"94",X"01",X"24",X"01",X"24",X"01",X"24",X"02",X"24",X"01",X"24",X"01",X"A4",
		X"01",X"A4",X"01",X"24",X"02",X"A4",X"02",X"24",X"02",X"A4",X"02",X"24",X"02",X"A4",X"02",X"04",
		X"02",X"04",X"01",X"04",X"01",X"04",X"01",X"04",X"01",X"24",X"02",X"24",X"01",X"24",X"01",X"A4",
		X"01",X"A4",X"01",X"24",X"02",X"A4",X"02",X"24",X"02",X"A4",X"02",X"24",X"02",X"A4",X"02",X"24",
		X"02",X"24",X"01",X"24",X"01",X"54",X"01",X"54",X"01",X"84",X"02",X"84",X"01",X"84",X"01",X"54",
		X"01",X"54",X"01",X"03",X"04",X"C0",X"02",X"03",X"04",X"03",X"02",X"84",X"06",X"A4",X"02",X"A4",
		X"01",X"A4",X"01",X"74",X"01",X"74",X"01",X"A4",X"02",X"74",X"02",X"A4",X"02",X"74",X"02",X"A4",
		X"02",X"74",X"02",X"A4",X"02",X"74",X"01",X"74",X"01",X"A4",X"01",X"A4",X"01",X"A4",X"02",X"A4",
		X"01",X"A4",X"01",X"64",X"01",X"64",X"01",X"A4",X"02",X"64",X"02",X"A4",X"02",X"64",X"02",X"A4",
		X"02",X"64",X"02",X"A4",X"02",X"64",X"01",X"64",X"01",X"A4",X"01",X"A4",X"01",X"F2",X"12",X"C0",
		X"02",X"03",X"02",X"03",X"02",X"C0",X"02",X"03",X"02",X"03",X"02",X"53",X"02",X"73",X"02",X"93",
		X"02",X"53",X"02",X"73",X"02",X"83",X"02",X"F0",X"30",X"08",X"F7",X"EA",X"9E",X"F0",X"20",X"0D",
		X"73",X"0F",X"A3",X"0F",X"33",X"14",X"A4",X"0F",X"03",X"0F",X"73",X"50",X"83",X"0F",X"02",X"0F",
		X"53",X"14",X"03",X"0F",X"53",X"0F",X"83",X"28",X"63",X"14",X"53",X"14",X"F3",X"02",X"ED",X"A0",
		X"F2",X"10",X"A3",X"05",X"A3",X"05",X"F2",X"00",X"93",X"02",X"83",X"02",X"F2",X"02",X"73",X"02",
		X"F2",X"03",X"63",X"02",X"F2",X"04",X"53",X"02",X"C0",X"1E",X"F2",X"0D",X"12",X"0F",X"B3",X"0F",
		X"A3",X"28",X"13",X"14",X"33",X"14",X"A3",X"28",X"B3",X"14",X"12",X"14",X"32",X"28",X"C0",X"0A",
		X"22",X"0A",X"C0",X"05",X"A3",X"0F",X"F0",X"20",X"0E",X"33",X"0F",X"73",X"0F",X"74",X"14",X"74",
		X"14",X"74",X"0A",X"A4",X"50",X"03",X"0F",X"53",X"0F",X"84",X"14",X"54",X"14",X"84",X"0A",X"F5",
		X"02",X"EE",X"1C",X"B4",X"28",X"84",X"14",X"23",X"14",X"F7",X"ED",X"F9",X"B4",X"28",X"84",X"14",
		X"B4",X"14",X"F2",X"10",X"13",X"05",X"13",X"05",X"F2",X"00",X"03",X"02",X"B4",X"02",X"F2",X"02",
		X"A4",X"02",X"F2",X"03",X"94",X"02",X"F2",X"04",X"84",X"02",X"C0",X"1E",X"F2",X"0E",X"A3",X"0F",
		X"83",X"0F",X"63",X"28",X"A4",X"14",X"A4",X"14",X"63",X"28",X"63",X"14",X"63",X"14",X"53",X"28",
		X"C0",X"0A",X"53",X"0A",X"C0",X"05",X"23",X"0F",X"F0",X"00",X"09",X"35",X"0F",X"35",X"05",X"35",
		X"0F",X"35",X"05",X"A5",X"0F",X"A5",X"05",X"A5",X"0F",X"A5",X"05",X"75",X"0F",X"75",X"05",X"45",
		X"0F",X"45",X"05",X"05",X"0F",X"05",X"05",X"75",X"0F",X"75",X"05",X"55",X"0F",X"55",X"05",X"55",
		X"0F",X"55",X"05",X"04",X"0F",X"04",X"05",X"04",X"0F",X"04",X"05",X"F5",X"02",X"EE",X"A2",X"B5",
		X"0F",X"B5",X"05",X"85",X"0F",X"85",X"05",X"55",X"0F",X"55",X"05",X"25",X"0F",X"25",X"05",X"F7",
		X"EE",X"5B",X"B5",X"05",X"25",X"0A",X"25",X"0A",X"25",X"0A",X"25",X"05",X"B5",X"05",X"25",X"0A",
		X"25",X"0A",X"25",X"0A",X"25",X"05",X"65",X"0F",X"65",X"05",X"14",X"0F",X"14",X"05",X"55",X"0F",
		X"55",X"05",X"14",X"0F",X"14",X"05",X"35",X"0F",X"35",X"05",X"A5",X"0F",X"A5",X"05",X"15",X"0F",
		X"15",X"05",X"A5",X"0F",X"A5",X"05",X"B6",X"0F",X"B6",X"05",X"A5",X"0F",X"A5",X"05",X"A6",X"0F",
		X"A6",X"05",X"65",X"0F",X"65",X"05",X"85",X"05",X"35",X"0A",X"35",X"0A",X"35",X"0A",X"35",X"05",
		X"C0",X"0A",X"A5",X"0A",X"C0",X"05",X"A5",X"0F",X"F0",X"40",X"08",X"33",X"0A",X"F2",X"10",X"33",
		X"05",X"33",X"05",X"33",X"05",X"33",X"05",X"33",X"05",X"33",X"05",X"F2",X"08",X"33",X"0A",X"F2",
		X"10",X"33",X"05",X"33",X"05",X"33",X"05",X"33",X"05",X"33",X"05",X"33",X"05",X"F2",X"08",X"43",
		X"14",X"43",X"0F",X"F2",X"10",X"03",X"05",X"C0",X"0A",X"F2",X"08",X"73",X"0A",X"C0",X"05",X"43",
		X"0F",X"53",X"0A",X"F2",X"10",X"53",X"05",X"53",X"05",X"53",X"05",X"53",X"05",X"53",X"05",X"53",
		X"05",X"F2",X"08",X"53",X"0A",X"F2",X"10",X"53",X"05",X"53",X"05",X"53",X"05",X"53",X"05",X"53",
		X"05",X"53",X"05",X"F5",X"02",X"EF",X"6E",X"F2",X"08",X"23",X"14",X"23",X"0F",X"F2",X"10",X"23",
		X"05",X"C0",X"0A",X"F2",X"08",X"B4",X"0A",X"C0",X"05",X"B4",X"0F",X"F7",X"EE",X"FB",X"F2",X"08",
		X"53",X"14",X"53",X"0F",X"F2",X"10",X"53",X"05",X"C0",X"0A",X"F2",X"08",X"23",X"0A",X"C0",X"05",
		X"23",X"0F",X"F2",X"09",X"63",X"14",X"63",X"0F",X"63",X"05",X"C0",X"0A",X"A3",X"0F",X"83",X"0F",
		X"63",X"14",X"63",X"0F",X"63",X"05",X"C0",X"0A",X"13",X"0A",X"C0",X"05",X"33",X"0F",X"33",X"14",
		X"33",X"0F",X"33",X"05",X"C0",X"0A",X"B4",X"0A",X"C0",X"05",X"13",X"0F",X"53",X"53",X"28",X"F0",
		X"40",X"08",X"74",X"0A",X"F2",X"10",X"74",X"05",X"74",X"05",X"74",X"05",X"74",X"05",X"74",X"05",
		X"74",X"05",X"F2",X"08",X"74",X"0A",X"F2",X"10",X"74",X"05",X"74",X"05",X"74",X"05",X"74",X"05",
		X"74",X"05",X"74",X"05",X"F2",X"08",X"74",X"14",X"74",X"0F",X"F2",X"10",X"74",X"05",X"C0",X"0A",
		X"F2",X"08",X"03",X"0A",X"C0",X"05",X"74",X"0F",X"84",X"0A",X"F2",X"10",X"84",X"05",X"84",X"05",
		X"84",X"05",X"84",X"05",X"84",X"05",X"84",X"05",X"F2",X"08",X"84",X"0A",X"F2",X"10",X"84",X"05",
		X"84",X"05",X"84",X"05",X"84",X"05",X"84",X"05",X"84",X"05",X"F5",X"02",X"F0",X"25",X"F2",X"08",
		X"54",X"14",X"54",X"0F",X"F2",X"10",X"54",X"05",X"C0",X"0A",X"F2",X"08",X"84",X"0A",X"C0",X"05",
		X"A4",X"0F",X"F7",X"EF",X"B2",X"F2",X"08",X"84",X"14",X"84",X"0F",X"F2",X"10",X"84",X"05",X"C0",
		X"0A",X"F2",X"08",X"84",X"0A",X"C0",X"05",X"84",X"0F",X"F2",X"09",X"A4",X"14",X"A4",X"0F",X"A4",
		X"05",X"C0",X"0A",X"13",X"0F",X"B4",X"0F",X"A4",X"14",X"A4",X"0F",X"A4",X"05",X"C0",X"0A",X"64",
		X"0A",X"C0",X"05",X"64",X"0F",X"B4",X"14",X"B4",X"0F",X"B4",X"05",X"C0",X"0A",X"64",X"0A",X"C0",
		X"05",X"64",X"0F",X"B4",X"28",X"A4",X"28",X"F0",X"10",X"00",X"A5",X"03",X"34",X"03",X"54",X"03",
		X"74",X"03",X"A4",X"04",X"33",X"06",X"53",X"08",X"F2",X"0F",X"A3",X"18",X"F0",X"10",X"01",X"75",
		X"03",X"A5",X"03",X"24",X"03",X"34",X"03",X"74",X"04",X"A4",X"06",X"33",X"08",X"F2",X"0F",X"53",
		X"18",X"F0",X"10",X"02",X"C0",X"03",X"A5",X"03",X"34",X"03",X"54",X"03",X"74",X"03",X"A4",X"04",
		X"33",X"06",X"53",X"08",X"F2",X"0F",X"33",X"18",X"F0",X"40",X"03",X"C0",X"03",X"75",X"03",X"A5",
		X"03",X"24",X"03",X"34",X"03",X"74",X"04",X"A4",X"06",X"33",X"08",X"F2",X"0F",X"A4",X"18",X"F0",
		X"50",X"04",X"C0",X"0C",X"A5",X"03",X"34",X"03",X"54",X"03",X"74",X"03",X"A4",X"03",X"33",X"03",
		X"53",X"03",X"73",X"03",X"A3",X"03",X"32",X"03",X"52",X"03",X"72",X"03",X"A2",X"0C",X"F0",X"50",
		X"05",X"C0",X"0C",X"75",X"03",X"A5",X"03",X"24",X"03",X"34",X"03",X"74",X"03",X"A4",X"03",X"23",
		X"03",X"33",X"03",X"73",X"03",X"A3",X"03",X"22",X"03",X"32",X"03",X"72",X"0C",X"F0",X"20",X"08",
		X"74",X"02",X"84",X"01",X"A4",X"01",X"03",X"01",X"A4",X"02",X"74",X"01",X"84",X"01",X"A4",X"01",
		X"03",X"01",X"A4",X"01",X"84",X"01",X"74",X"01",X"54",X"01",X"34",X"02",X"54",X"01",X"74",X"01",
		X"84",X"01",X"74",X"02",X"34",X"01",X"54",X"01",X"74",X"01",X"84",X"01",X"74",X"01",X"54",X"01",
		X"34",X"01",X"F6",X"02",X"F1",X"65",X"24",X"01",X"04",X"02",X"54",X"02",X"24",X"01",X"A5",X"01",
		X"04",X"02",X"54",X"02",X"24",X"01",X"A5",X"01",X"F2",X"1C",X"C0",X"01",X"04",X"01",X"54",X"01",
		X"24",X"01",X"A5",X"01",X"04",X"01",X"54",X"01",X"24",X"01",X"A5",X"01",X"F3",X"02",X"F1",X"56",
		X"F2",X"08",X"F7",X"F1",X"00",X"74",X"01",X"84",X"02",X"33",X"01",X"B4",X"01",X"53",X"01",X"83",
		X"01",X"73",X"03",X"53",X"01",X"33",X"01",X"23",X"01",X"F2",X"10",X"33",X"01",X"33",X"01",X"33",
		X"01",X"33",X"01",X"C0",X"02",X"33",X"01",X"C0",X"01",X"33",X"02",X"33",X"01",X"33",X"01",X"33",
		X"02",X"C0",X"02",X"F0",X"50",X"15",X"A5",X"03",X"A5",X"03",X"A5",X"03",X"A5",X"03",X"85",X"03",
		X"75",X"03",X"75",X"03",X"75",X"03",X"75",X"03",X"55",X"03",X"F6",X"02",X"F1",X"BD",X"35",X"03",
		X"55",X"03",X"F3",X"03",X"F1",X"AE",X"75",X"03",X"85",X"03",X"F7",X"F1",X"96",X"F0",X"50",X"15",
		X"75",X"03",X"75",X"03",X"75",X"03",X"75",X"03",X"55",X"03",X"35",X"03",X"35",X"03",X"35",X"03",
		X"35",X"03",X"25",X"03",X"F6",X"02",X"F1",X"E7",X"05",X"03",X"25",X"03",X"F3",X"03",X"F1",X"D8",
		X"35",X"03",X"55",X"03",X"F7",X"F1",X"C0",X"F0",X"50",X"15",X"35",X"03",X"35",X"03",X"35",X"03",
		X"35",X"03",X"15",X"03",X"25",X"03",X"15",X"03",X"05",X"03",X"05",X"03",X"A6",X"03",X"F6",X"02",
		X"F2",X"11",X"86",X"03",X"A6",X"03",X"F3",X"03",X"F2",X"02",X"05",X"03",X"25",X"03",X"F7",X"F1",
		X"EA",X"F0",X"50",X"15",X"35",X"03",X"25",X"03",X"15",X"03",X"05",X"03",X"B6",X"03",X"A6",X"03",
		X"A6",X"03",X"A6",X"03",X"86",X"03",X"76",X"03",X"F6",X"02",X"F2",X"3B",X"56",X"03",X"76",X"03",
		X"F3",X"03",X"F2",X"2C",X"86",X"03",X"A6",X"03",X"F7",X"F2",X"14",X"F0",X"20",X"05",X"F1",X"20",
		X"13",X"01",X"23",X"01",X"33",X"01",X"43",X"01",X"53",X"01",X"63",X"01",X"73",X"01",X"83",X"01",
		X"93",X"01",X"C0",X"01",X"93",X"01",X"83",X"01",X"73",X"01",X"63",X"01",X"53",X"01",X"43",X"01",
		X"33",X"01",X"C0",X"02",X"73",X"01",X"63",X"01",X"53",X"01",X"43",X"01",X"33",X"01",X"23",X"01",
		X"13",X"01",X"C0",X"02",X"F1",X"40",X"84",X"01",X"94",X"01",X"A4",X"01",X"B4",X"01",X"03",X"01",
		X"13",X"01",X"23",X"01",X"33",X"01",X"43",X"01",X"C0",X"01",X"43",X"01",X"33",X"01",X"23",X"01",
		X"13",X"01",X"03",X"01",X"B4",X"01",X"A4",X"01",X"C0",X"02",X"23",X"01",X"13",X"01",X"03",X"01",
		X"B4",X"01",X"A4",X"01",X"94",X"01",X"84",X"01",X"C0",X"02",X"F1",X"70",X"03",X"01",X"13",X"01",
		X"23",X"01",X"33",X"01",X"43",X"01",X"53",X"01",X"63",X"01",X"73",X"01",X"83",X"01",X"C0",X"01",
		X"83",X"01",X"73",X"01",X"63",X"01",X"53",X"01",X"43",X"01",X"33",X"01",X"23",X"01",X"C0",X"02",
		X"63",X"01",X"53",X"01",X"43",X"01",X"33",X"01",X"23",X"01",X"13",X"01",X"03",X"01",X"C0",X"02",
		X"F0",X"20",X"06",X"14",X"01",X"24",X"01",X"34",X"01",X"44",X"01",X"54",X"01",X"64",X"01",X"74",
		X"01",X"84",X"01",X"94",X"01",X"C0",X"01",X"34",X"01",X"44",X"01",X"54",X"01",X"64",X"01",X"74",
		X"01",X"84",X"01",X"94",X"01",X"C0",X"02",X"34",X"01",X"44",X"01",X"54",X"01",X"64",X"01",X"74",
		X"01",X"84",X"01",X"94",X"01",X"C0",X"02",X"F1",X"40",X"85",X"01",X"95",X"01",X"A5",X"01",X"B5",
		X"01",X"04",X"01",X"14",X"01",X"24",X"01",X"34",X"01",X"44",X"01",X"C0",X"01",X"A5",X"01",X"B5",
		X"01",X"04",X"01",X"14",X"01",X"24",X"01",X"34",X"01",X"44",X"01",X"C0",X"02",X"A5",X"01",X"B5",
		X"01",X"04",X"01",X"14",X"01",X"24",X"01",X"34",X"01",X"44",X"01",X"C0",X"02",X"F1",X"70",X"04",
		X"01",X"14",X"01",X"24",X"01",X"34",X"01",X"44",X"01",X"54",X"01",X"64",X"01",X"74",X"01",X"84",
		X"01",X"C0",X"01",X"24",X"01",X"34",X"01",X"44",X"01",X"54",X"01",X"64",X"01",X"74",X"01",X"84",
		X"01",X"C0",X"02",X"24",X"01",X"34",X"01",X"44",X"01",X"54",X"01",X"64",X"01",X"74",X"01",X"84",
		X"01",X"C0",X"02",X"F0",X"20",X"06",X"C0",X"03",X"F7",X"F2",X"3E",X"20",X"05",X"C0",X"03",X"F7",
		X"F2",X"E3",X"40",X"00",X"72",X"01",X"62",X"01",X"52",X"01",X"42",X"01",X"32",X"01",X"22",X"01",
		X"62",X"01",X"52",X"01",X"42",X"01",X"32",X"01",X"22",X"01",X"12",X"01",X"52",X"01",X"42",X"01",
		X"32",X"01",X"22",X"01",X"12",X"01",X"02",X"01",X"42",X"01",X"32",X"01",X"22",X"01",X"12",X"01",
		X"02",X"01",X"B3",X"01",X"32",X"01",X"22",X"01",X"12",X"01",X"02",X"01",X"B3",X"01",X"A3",X"01",
		X"C0",X"01",X"F0",X"40",X"02",X"C0",X"03",X"73",X"01",X"63",X"01",X"53",X"01",X"43",X"01",X"33",
		X"01",X"23",X"01",X"63",X"01",X"53",X"01",X"43",X"01",X"33",X"01",X"23",X"01",X"13",X"01",X"53",
		X"01",X"43",X"01",X"33",X"01",X"23",X"01",X"13",X"01",X"03",X"01",X"43",X"01",X"33",X"01",X"23",
		X"01",X"13",X"01",X"03",X"01",X"B4",X"01",X"33",X"01",X"23",X"01",X"13",X"01",X"F0",X"20",X"00",
		X"73",X"01",X"02",X"01",X"42",X"01",X"F3",X"08",X"F4",X"10",X"F0",X"20",X"00",X"43",X"01",X"73",
		X"01",X"02",X"01",X"F3",X"08",X"F4",X"1D",X"F0",X"50",X"00",X"42",X"01",X"52",X"01",X"12",X"01",
		X"52",X"01",X"F3",X"06",X"F4",X"2A",X"F0",X"50",X"00",X"02",X"01",X"12",X"01",X"83",X"01",X"12",
		X"01",X"F3",X"06",X"F4",X"39",X"F0",X"20",X"0D",X"04",X"12",X"F2",X"10",X"73",X"06",X"73",X"06",
		X"43",X"06",X"F1",X"50",X"F2",X"0D",X"B3",X"02",X"F2",X"13",X"02",X"16",X"C0",X"0C",X"F0",X"40",
		X"0D",X"04",X"12",X"F2",X"10",X"43",X"06",X"43",X"06",X"03",X"06",X"F1",X"70",X"F2",X"0D",X"B2",
		X"02",X"F2",X"13",X"01",X"16",X"C0",X"0C",X"F0",X"40",X"02",X"C0",X"04",X"32",X"01",X"52",X"01",
		X"32",X"01",X"52",X"01",X"32",X"01",X"C0",X"02",X"F2",X"01",X"01",X"01",X"B2",X"01",X"A2",X"01",
		X"92",X"01",X"F2",X"00",X"82",X"01",X"72",X"01",X"62",X"01",X"52",X"01",X"82",X"01",X"72",X"01",
		X"62",X"01",X"52",X"01",X"42",X"01",X"32",X"01",X"22",X"01",X"12",X"01",X"42",X"01",X"32",X"01",
		X"22",X"01",X"12",X"01",X"02",X"01",X"B3",X"01",X"A3",X"01",X"93",X"01",X"F2",X"01",X"12",X"01",
		X"02",X"01",X"B3",X"01",X"A3",X"01",X"93",X"01",X"83",X"01",X"73",X"01",X"63",X"01",X"A3",X"01",
		X"93",X"01",X"83",X"01",X"73",X"01",X"63",X"01",X"53",X"01",X"43",X"01",X"33",X"01",X"F2",X"02",
		X"63",X"01",X"53",X"01",X"43",X"01",X"33",X"01",X"23",X"01",X"13",X"01",X"03",X"01",X"B4",X"01",
		X"F2",X"03",X"03",X"01",X"B4",X"01",X"A4",X"01",X"94",X"01",X"84",X"01",X"74",X"01",X"64",X"01",
		X"54",X"01",X"F2",X"04",X"74",X"01",X"64",X"01",X"54",X"01",X"44",X"01",X"34",X"01",X"24",X"01",
		X"14",X"01",X"04",X"01",X"F2",X"05",X"14",X"01",X"04",X"01",X"B5",X"01",X"A5",X"01",X"95",X"01",
		X"85",X"01",X"75",X"01",X"65",X"01",X"C0",X"04",X"F0",X"10",X"00",X"42",X"01",X"02",X"01",X"22",
		X"01",X"B3",X"01",X"C0",X"01",X"02",X"01",X"73",X"01",X"93",X"01",X"43",X"01",X"C0",X"01",X"63",
		X"01",X"33",X"01",X"43",X"01",X"03",X"01",X"C0",X"01",X"23",X"01",X"A4",X"01",X"03",X"01",X"94",
		X"01",X"C0",X"01",X"A4",X"01",X"74",X"01",X"94",X"01",X"54",X"01",X"C0",X"01",X"74",X"01",X"54",
		X"01",X"44",X"01",X"24",X"01",X"04",X"01",X"A5",X"01",X"95",X"01",X"75",X"01",X"C0",X"01",X"65",
		X"01",X"B5",X"01",X"95",X"01",X"24",X"01",X"C0",X"01",X"04",X"01",X"54",X"01",X"34",X"01",X"84",
		X"01",X"C0",X"01",X"F2",X"01",X"64",X"01",X"B4",X"01",X"94",X"01",X"23",X"01",X"C0",X"01",X"04",
		X"01",X"54",X"01",X"34",X"01",X"84",X"01",X"C0",X"01",X"F2",X"02",X"64",X"01",X"B4",X"01",X"94",
		X"01",X"23",X"01",X"C0",X"01",X"04",X"01",X"54",X"01",X"34",X"01",X"84",X"01",X"C0",X"01",X"F2",
		X"03",X"64",X"01",X"B4",X"01",X"94",X"01",X"23",X"01",X"C0",X"01",X"04",X"01",X"54",X"01",X"34",
		X"01",X"84",X"01",X"C0",X"01",X"F2",X"04",X"64",X"01",X"B4",X"01",X"94",X"01",X"23",X"01",X"C0",
		X"01",X"04",X"01",X"54",X"01",X"34",X"01",X"84",X"01",X"C0",X"01",X"64",X"01",X"B4",X"01",X"94",
		X"01",X"23",X"01",X"C0",X"01",X"F0",X"10",X"00",X"C0",X"03",X"F7",X"F5",X"2B",X"F0",X"10",X"08",
		X"32",X"04",X"B3",X"02",X"12",X"04",X"62",X"02",X"C0",X"01",X"F0",X"40",X"08",X"B3",X"04",X"63",
		X"02",X"A3",X"04",X"12",X"02",X"C0",X"01",X"F0",X"20",X"00",X"44",X"01",X"34",X"01",X"24",X"01",
		X"34",X"01",X"44",X"01",X"54",X"01",X"64",X"01",X"C0",X"01",X"33",X"01",X"23",X"01",X"13",X"01",
		X"03",X"01",X"B4",X"01",X"A4",X"01",X"94",X"01",X"F2",X"02",X"84",X"01",X"74",X"01",X"F2",X"03",
		X"64",X"01",X"54",X"01",X"F2",X"04",X"44",X"01",X"34",X"01",X"24",X"01",X"04",X"01",X"A5",X"01",
		X"85",X"01",X"65",X"01",X"45",X"01",X"25",X"01",X"05",X"01",X"A6",X"01",X"86",X"01",X"F0",X"70",
		X"00",X"73",X"01",X"63",X"01",X"53",X"01",X"63",X"01",X"73",X"01",X"83",X"01",X"93",X"01",X"C0",
		X"01",X"62",X"01",X"52",X"01",X"42",X"01",X"32",X"01",X"22",X"01",X"12",X"01",X"03",X"01",X"F2",
		X"02",X"A3",X"01",X"93",X"01",X"F2",X"03",X"73",X"01",X"53",X"01",X"F2",X"04",X"13",X"01",X"B4",
		X"01",X"94",X"01",X"74",X"01",X"44",X"01",X"34",X"01",X"B5",X"01",X"85",X"01",X"65",X"01",X"45",
		X"01",X"25",X"01",X"C0",X"01",X"F0",X"10",X"00",X"C0",X"0A",X"24",X"01",X"14",X"01",X"04",X"01",
		X"14",X"01",X"24",X"01",X"34",X"01",X"44",X"01",X"C0",X"01",X"F2",X"02",X"B3",X"01",X"A3",X"01",
		X"93",X"01",X"83",X"01",X"73",X"01",X"F2",X"04",X"63",X"01",X"53",X"01",X"43",X"01",X"33",X"01",
		X"23",X"01",X"13",X"01",X"03",X"01",X"B4",X"01",X"F0",X"50",X"00",X"C0",X"0A",X"74",X"01",X"64",
		X"01",X"54",X"01",X"64",X"01",X"74",X"01",X"84",X"01",X"94",X"01",X"C0",X"01",X"F2",X"02",X"63",
		X"01",X"53",X"01",X"43",X"01",X"33",X"01",X"23",X"01",X"F2",X"04",X"13",X"01",X"03",X"01",X"B4",
		X"01",X"A4",X"01",X"94",X"01",X"84",X"01",X"74",X"01",X"64",X"01",X"F0",X"50",X"10",X"35",X"06",
		X"45",X"06",X"F7",X"F6",X"FE",X"50",X"10",X"A6",X"03",X"25",X"03",X"F7",X"F7",X"07",X"40",X"14",
		X"C0",X"30",X"A5",X"24",X"F2",X"10",X"A5",X"04",X"A5",X"04",X"A5",X"04",X"F2",X"14",X"95",X"24",
		X"F2",X"01",X"55",X"0C",X"F2",X"14",X"85",X"30",X"F2",X"10",X"75",X"04",X"F2",X"01",X"35",X"02",
		X"75",X"2A",X"F0",X"40",X"14",X"C0",X"30",X"65",X"24",X"F2",X"10",X"65",X"04",X"65",X"04",X"65",
		X"04",X"F2",X"14",X"55",X"24",X"F2",X"01",X"05",X"0C",X"F2",X"14",X"55",X"30",X"F2",X"10",X"35",
		X"04",X"F2",X"01",X"A6",X"02",X"35",X"2A",X"F0",X"40",X"03",X"C0",X"32",X"A5",X"24",X"A5",X"04",
		X"A5",X"04",X"A5",X"04",X"95",X"24",X"55",X"0C",X"85",X"2E",X"F2",X"11",X"75",X"04",X"F2",X"03",
		X"35",X"02",X"75",X"2A",X"F0",X"40",X"02",X"32",X"01",X"22",X"01",X"12",X"01",X"02",X"01",X"B3",
		X"01",X"A3",X"01",X"93",X"01",X"83",X"01",X"12",X"01",X"02",X"01",X"B3",X"01",X"A3",X"01",X"93",
		X"01",X"83",X"01",X"73",X"01",X"63",X"01",X"B3",X"01",X"A3",X"01",X"93",X"01",X"83",X"01",X"73",
		X"01",X"63",X"01",X"53",X"01",X"43",X"01",X"93",X"01",X"83",X"01",X"73",X"01",X"63",X"01",X"53",
		X"01",X"43",X"01",X"33",X"01",X"23",X"01",X"73",X"01",X"63",X"01",X"53",X"01",X"43",X"01",X"33",
		X"01",X"23",X"01",X"13",X"01",X"03",X"01",X"53",X"01",X"43",X"01",X"33",X"01",X"23",X"01",X"13",
		X"01",X"03",X"01",X"B4",X"01",X"A4",X"01",X"33",X"01",X"23",X"01",X"13",X"01",X"03",X"01",X"B4",
		X"01",X"A4",X"01",X"94",X"01",X"84",X"01",X"13",X"01",X"03",X"01",X"B4",X"01",X"A4",X"01",X"94",
		X"01",X"84",X"01",X"74",X"01",X"64",X"01",X"B4",X"01",X"A4",X"01",X"94",X"01",X"84",X"01",X"74",
		X"01",X"64",X"01",X"54",X"01",X"44",X"01",X"94",X"01",X"84",X"01",X"74",X"01",X"64",X"01",X"54",
		X"01",X"44",X"01",X"34",X"01",X"24",X"01",X"74",X"01",X"64",X"01",X"54",X"01",X"44",X"01",X"34",
		X"01",X"24",X"01",X"14",X"01",X"04",X"01",X"F2",X"03",X"54",X"01",X"44",X"01",X"34",X"01",X"24",
		X"01",X"14",X"01",X"04",X"01",X"B5",X"01",X"A5",X"01",X"F2",X"04",X"34",X"01",X"24",X"01",X"14",
		X"01",X"04",X"01",X"B5",X"01",X"A5",X"01",X"95",X"01",X"85",X"01",X"F0",X"10",X"00",X"A3",X"01",
		X"B3",X"01",X"A3",X"01",X"B3",X"01",X"C0",X"02",X"63",X"01",X"73",X"01",X"83",X"01",X"C0",X"01",
		X"02",X"01",X"22",X"01",X"52",X"01",X"92",X"01",X"F0",X"20",X"03",X"72",X"07",X"42",X"07",X"52",
		X"07",X"22",X"07",X"F2",X"02",X"72",X"06",X"42",X"06",X"52",X"06",X"22",X"06",X"F2",X"01",X"72",
		X"05",X"42",X"05",X"52",X"05",X"22",X"05",X"F2",X"00",X"72",X"04",X"42",X"04",X"52",X"04",X"22",
		X"04",X"72",X"04",X"42",X"04",X"52",X"04",X"22",X"04",X"72",X"04",X"42",X"04",X"52",X"04",X"22",
		X"04",X"F0",X"30",X"03",X"04",X"07",X"75",X"07",X"B5",X"07",X"75",X"07",X"F2",X"02",X"03",X"06",
		X"74",X"06",X"B4",X"06",X"74",X"06",X"F2",X"01",X"03",X"05",X"74",X"05",X"B4",X"05",X"74",X"05",
		X"F2",X"00",X"02",X"04",X"73",X"04",X"B3",X"04",X"73",X"04",X"02",X"04",X"73",X"04",X"B3",X"04",
		X"73",X"04",X"02",X"04",X"73",X"04",X"B3",X"04",X"73",X"04",X"F0",X"50",X"08",X"93",X"02",X"53",
		X"01",X"73",X"02",X"F2",X"07",X"02",X"06",X"C0",X"01",X"F0",X"00",X"08",X"53",X"01",X"03",X"01",
		X"94",X"01",X"03",X"02",X"F2",X"03",X"03",X"06",X"C0",X"01",X"F0",X"00",X"08",X"35",X"01",X"45",
		X"01",X"55",X"01",X"45",X"01",X"35",X"02",X"35",X"01",X"45",X"01",X"55",X"01",X"65",X"01",X"73",
		X"01",X"63",X"01",X"53",X"01",X"43",X"01",X"33",X"02",X"33",X"01",X"43",X"01",X"53",X"01",X"63",
		X"01",X"73",X"01",X"83",X"01",X"93",X"01",X"A3",X"01",X"93",X"01",X"83",X"01",X"73",X"01",X"63",
		X"01",X"53",X"01",X"43",X"01",X"33",X"02",X"C0",X"05",X"F0",X"00",X"08",X"05",X"01",X"15",X"01",
		X"25",X"01",X"15",X"01",X"05",X"02",X"03",X"01",X"13",X"01",X"23",X"01",X"33",X"01",X"43",X"01",
		X"33",X"01",X"23",X"01",X"13",X"01",X"03",X"02",X"03",X"01",X"13",X"01",X"23",X"01",X"33",X"01",
		X"43",X"01",X"53",X"01",X"63",X"01",X"73",X"01",X"63",X"01",X"53",X"01",X"43",X"01",X"33",X"01",
		X"23",X"01",X"13",X"01",X"03",X"02",X"C0",X"05",X"F0",X"10",X"00",X"12",X"12",X"B3",X"03",X"12",
		X"03",X"32",X"06",X"B3",X"06",X"12",X"03",X"83",X"03",X"C0",X"03",X"53",X"03",X"12",X"0C",X"B3",
		X"04",X"12",X"04",X"B3",X"04",X"A3",X"24",X"A3",X"24",X"A3",X"0C",X"C0",X"18",X"F0",X"10",X"03",
		X"C0",X"02",X"F7",X"F9",X"7B",X"10",X"18",X"85",X"06",X"F2",X"1E",X"85",X"02",X"85",X"02",X"85",
		X"02",X"F2",X"18",X"85",X"06",X"F2",X"1E",X"85",X"02",X"85",X"02",X"85",X"02",X"85",X"02",X"85",
		X"02",X"85",X"02",X"85",X"02",X"85",X"02",X"85",X"02",X"F6",X"02",X"F9",X"D0",X"F7",X"F9",X"A7",
		X"F2",X"18",X"A5",X"06",X"F2",X"1E",X"A5",X"02",X"A5",X"02",X"A5",X"02",X"F2",X"18",X"A5",X"06",
		X"F2",X"1E",X"A5",X"02",X"A5",X"02",X"A5",X"02",X"A5",X"02",X"A5",X"02",X"A5",X"02",X"A5",X"02",
		X"A5",X"02",X"A5",X"02",X"F3",X"02",X"F9",X"D0",X"F2",X"04",X"A5",X"0C",X"C0",X"18",X"F0",X"10",
		X"03",X"63",X"24",X"63",X"24",X"53",X"24",X"53",X"24",X"53",X"0C",X"C0",X"18",X"F0",X"10",X"03",
		X"33",X"24",X"33",X"24",X"23",X"24",X"23",X"24",X"23",X"0C",X"C0",X"18",X"F0",X"40",X"02",X"55",
		X"02",X"75",X"02",X"95",X"02",X"C0",X"03",X"04",X"02",X"24",X"02",X"44",X"02",X"C0",X"03",X"74",
		X"02",X"94",X"02",X"B4",X"02",X"C0",X"03",X"F1",X"70",X"F2",X"10",X"83",X"08",X"F0",X"31",X"39",
		X"38",X"34",X"20",X"4E",X"41",X"4D",X"43",X"4F",X"20",X"41",X"4C",X"4C",X"20",X"52",X"49",X"47",
		X"48",X"54",X"53",X"20",X"52",X"45",X"53",X"45",X"52",X"56",X"45",X"44",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"46",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E0",X"55",X"FF",X"FF",X"FF",X"FF",X"E0",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
