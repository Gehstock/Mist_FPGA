library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity a1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of a1 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"C0",X"40",X"C0",X"40",X"01",X"01",X"FC",X"01",X"01",X"FE",X"C0",X"30",X"A0",X"12",X"50",X"02",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"50",X"C0",X"50",X"01",X"01",X"FC",X"01",X"01",X"FE",X"C0",X"30",X"A0",X"12",X"50",X"02",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"08",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"08",X"00",X"00",X"C0",X"9C",X"01",X"00",X"00",X"08",X"08",X"00",X"00",X"C0",X"80",
		X"01",X"00",X"00",X"08",X"08",X"8E",X"E3",X"00",X"41",X"80",X"E3",X"38",X"08",X"08",X"51",X"14",
		X"01",X"3E",X"40",X"14",X"45",X"08",X"08",X"51",X"14",X"41",X"22",X"41",X"14",X"45",X"08",X"08",
		X"51",X"14",X"41",X"2A",X"41",X"14",X"45",X"08",X"08",X"51",X"14",X"41",X"22",X"41",X"14",X"45",
		X"08",X"08",X"51",X"14",X"01",X"3E",X"40",X"14",X"45",X"08",X"08",X"8E",X"E3",X"00",X"41",X"80",
		X"E3",X"38",X"08",X"08",X"00",X"00",X"C0",X"80",X"01",X"00",X"00",X"08",X"08",X"00",X"00",X"C0",
		X"9C",X"01",X"00",X"00",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",
		X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"08",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"08",X"00",X"00",X"C0",X"9C",X"01",X"00",X"00",X"08",X"08",X"00",X"00",X"C0",X"80",
		X"01",X"00",X"00",X"08",X"08",X"9F",X"E3",X"00",X"41",X"C0",X"E7",X"38",X"08",X"08",X"41",X"14",
		X"01",X"3E",X"40",X"10",X"45",X"08",X"08",X"4F",X"14",X"41",X"22",X"C1",X"13",X"45",X"08",X"08",
		X"50",X"14",X"41",X"2A",X"01",X"14",X"45",X"08",X"08",X"50",X"14",X"41",X"22",X"01",X"14",X"45",
		X"08",X"08",X"51",X"14",X"01",X"3E",X"40",X"14",X"45",X"08",X"08",X"8E",X"E3",X"00",X"41",X"80",
		X"E3",X"38",X"08",X"08",X"00",X"00",X"C0",X"80",X"01",X"00",X"00",X"08",X"08",X"00",X"00",X"C0",
		X"9C",X"01",X"00",X"00",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",
		X"FC",X"90",X"31",X"46",X"02",X"51",X"4A",X"C9",X"31",X"52",X"4A",X"49",X"49",X"52",X"4A",X"49",
		X"09",X"52",X"4A",X"49",X"09",X"92",X"33",X"09",X"09",X"12",X"4A",X"49",X"49",X"12",X"4A",X"C9",
		X"31",X"12",X"4A",X"49",X"02",X"11",X"4A",X"49",X"FC",X"10",X"32",X"46",X"35",X"25",X"05",X"55",
		X"55",X"05",X"55",X"75",X"02",X"55",X"57",X"02",X"35",X"55",X"02",X"00",X"00",X"00",X"DD",X"B9",
		X"03",X"45",X"88",X"02",X"4D",X"89",X"02",X"45",X"89",X"02",X"C5",X"B9",X"0B",X"37",X"37",X"1D",
		X"51",X"51",X"09",X"31",X"53",X"09",X"51",X"51",X"09",X"57",X"37",X"09",X"F0",X"FF",X"01",X"10",
		X"00",X"01",X"10",X"00",X"01",X"10",X"00",X"01",X"10",X"00",X"01",X"10",X"00",X"01",X"10",X"00",
		X"01",X"10",X"00",X"01",X"10",X"00",X"01",X"10",X"00",X"01",X"F0",X"FF",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C3",X"8F",X"5A",X"C3",X"99",X"5A",X"C3",X"CA",X"5A",X"C3",X"46",X"5B",X"C3",X"90",X"5B",X"3A",
		X"8C",X"21",X"FE",X"02",X"D8",X"CD",X"83",X"5A",X"C9",X"7E",X"B7",X"C8",X"23",X"A6",X"C0",X"7D",
		X"D6",X"08",X"6F",X"7E",X"FE",X"70",X"D0",X"7D",X"D6",X"07",X"6F",X"3A",X"6A",X"20",X"96",X"DA",
		X"C0",X"5A",X"07",X"07",X"07",X"E6",X"07",X"C6",X"04",X"47",X"7D",X"C6",X"04",X"6F",X"70",X"C9",
		X"07",X"07",X"07",X"F6",X"F8",X"D6",X"04",X"C3",X"B9",X"5A",X"DB",X"02",X"E6",X"30",X"FE",X"30",
		X"C8",X"21",X"CB",X"5B",X"11",X"E0",X"20",X"06",X"09",X"FF",X"DB",X"02",X"E6",X"03",X"4F",X"07",
		X"07",X"07",X"81",X"4F",X"06",X"00",X"21",X"D8",X"57",X"09",X"CD",X"0E",X"5B",X"CD",X"03",X"5B",
		X"CD",X"03",X"5B",X"EB",X"36",X"FF",X"21",X"E0",X"20",X"22",X"80",X"21",X"21",X"A2",X"29",X"22",
		X"82",X"21",X"C9",X"EB",X"36",X"2C",X"23",X"36",X"20",X"23",X"EB",X"23",X"23",X"23",X"23",X"23",
		X"CD",X"2F",X"5B",X"2B",X"CD",X"1C",X"5B",X"2B",X"CD",X"1C",X"5B",X"C9",X"7E",X"07",X"07",X"07",
		X"07",X"E6",X"0F",X"C6",X"30",X"12",X"13",X"7E",X"E6",X"0F",X"C6",X"30",X"12",X"13",X"C9",X"7E",
		X"07",X"07",X"07",X"07",X"E6",X"0F",X"CA",X"3D",X"5B",X"C6",X"30",X"12",X"13",X"7E",X"E6",X"0F",
		X"C8",X"C6",X"30",X"12",X"13",X"C9",X"2A",X"80",X"21",X"7D",X"B4",X"C0",X"CD",X"7A",X"5B",X"DA",
		X"70",X"5B",X"3E",X"20",X"21",X"E0",X"20",X"BE",X"C8",X"06",X"1F",X"77",X"23",X"05",X"C2",X"5B",
		X"5B",X"36",X"FF",X"21",X"E0",X"20",X"22",X"80",X"21",X"21",X"A2",X"29",X"22",X"82",X"21",X"C9",
		X"3A",X"E0",X"20",X"FE",X"20",X"C0",X"CD",X"86",X"5A",X"C9",X"3E",X"34",X"21",X"03",X"22",X"BE",
		X"D0",X"21",X"23",X"22",X"BE",X"D0",X"21",X"43",X"22",X"BE",X"D0",X"21",X"63",X"22",X"BE",X"C9",
		X"3A",X"04",X"20",X"B7",X"CA",X"B2",X"5B",X"3A",X"12",X"20",X"0F",X"0F",X"0F",X"E6",X"0E",X"21",
		X"BB",X"5B",X"85",X"D2",X"A7",X"5B",X"24",X"6F",X"7E",X"32",X"82",X"22",X"23",X"7E",X"32",X"A2",
		X"22",X"C9",X"3A",X"8C",X"21",X"FE",X"01",X"D8",X"C3",X"97",X"5B",X"30",X"D8",X"D8",X"D8",X"40",
		X"D0",X"D0",X"20",X"D0",X"D0",X"E0",X"C0",X"30",X"20",X"E0",X"20",X"42",X"4F",X"4E",X"55",X"53",
		X"20",X"41",X"54",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F3",X"C3",X"2E",X"5C",X"C6",X"A4",X"5A",X"09",X"67",X"4A",X"B7",X"FA",X"A3",X"66",X"72",X"03",
		X"C1",X"DA",X"54",X"10",X"C3",X"B3",X"5E",X"C3",X"B4",X"5E",X"C3",X"B6",X"5E",X"C3",X"2D",X"5C",
		X"C3",X"2C",X"5C",X"C3",X"58",X"5E",X"C3",X"B7",X"5E",X"C3",X"BA",X"5E",X"C9",X"C9",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"06",X"00",X"21",
		X"00",X"20",X"70",X"7E",X"A8",X"4F",X"7D",X"E6",X"01",X"79",X"CA",X"52",X"5C",X"B3",X"5F",X"C3",
		X"54",X"5C",X"B2",X"57",X"78",X"2F",X"77",X"AE",X"4F",X"7D",X"E6",X"01",X"79",X"CA",X"65",X"5C",
		X"B3",X"5F",X"C3",X"67",X"5C",X"B2",X"57",X"23",X"7C",X"FE",X"40",X"C2",X"42",X"5C",X"D3",X"02",
		X"21",X"00",X"20",X"06",X"00",X"70",X"04",X"C2",X"7B",X"5C",X"04",X"23",X"7C",X"FE",X"40",X"C2",
		X"75",X"5C",X"D3",X"02",X"21",X"00",X"20",X"06",X"00",X"7E",X"A8",X"4F",X"7D",X"E6",X"01",X"79",
		X"CA",X"98",X"5C",X"B3",X"5F",X"C3",X"9A",X"5C",X"B2",X"57",X"04",X"C2",X"9F",X"5C",X"04",X"23",
		X"7C",X"FE",X"40",X"C2",X"89",X"5C",X"D3",X"02",X"21",X"00",X"20",X"AF",X"77",X"23",X"7C",X"FE",
		X"40",X"C2",X"AB",X"5C",X"3E",X"08",X"32",X"43",X"20",X"D3",X"00",X"7B",X"B2",X"C2",X"2B",X"5E",
		X"21",X"DE",X"5C",X"22",X"80",X"21",X"21",X"10",X"2D",X"22",X"82",X"21",X"CD",X"1F",X"5E",X"C3",
		X"ED",X"5C",X"D3",X"02",X"DB",X"00",X"E6",X"80",X"C2",X"D2",X"5C",X"C3",X"ED",X"5C",X"52",X"41",
		X"4D",X"20",X"54",X"45",X"53",X"54",X"53",X"20",X"47",X"4F",X"4F",X"44",X"FF",X"21",X"4F",X"5E",
		X"22",X"80",X"21",X"21",X"81",X"2B",X"22",X"82",X"21",X"CD",X"1F",X"5E",X"21",X"00",X"00",X"22",
		X"70",X"23",X"AF",X"32",X"72",X"23",X"CD",X"30",X"5D",X"CD",X"30",X"5D",X"CD",X"30",X"5D",X"CD",
		X"30",X"5D",X"21",X"00",X"40",X"22",X"70",X"23",X"CD",X"30",X"5D",X"CD",X"30",X"5D",X"CD",X"30",
		X"5D",X"CD",X"78",X"5D",X"D3",X"02",X"DB",X"00",X"E6",X"40",X"C2",X"24",X"5D",X"C3",X"C9",X"01",
		X"CD",X"37",X"5D",X"CD",X"6A",X"5D",X"C9",X"2A",X"70",X"23",X"44",X"4D",X"21",X"00",X"00",X"11",
		X"00",X"00",X"0A",X"5F",X"19",X"03",X"79",X"B7",X"C2",X"42",X"5D",X"78",X"E6",X"07",X"C2",X"42",
		X"5D",X"EB",X"60",X"69",X"22",X"70",X"23",X"21",X"72",X"23",X"7E",X"34",X"34",X"21",X"04",X"5C",
		X"85",X"D2",X"65",X"5D",X"24",X"6F",X"4E",X"23",X"46",X"C9",X"79",X"BB",X"C2",X"D9",X"5D",X"78",
		X"BA",X"C2",X"D9",X"5D",X"CD",X"BE",X"5D",X"C9",X"CD",X"37",X"5D",X"60",X"69",X"78",X"06",X"00",
		X"09",X"4F",X"09",X"44",X"4D",X"CD",X"6A",X"5D",X"C9",X"3A",X"72",X"23",X"11",X"80",X"01",X"21",
		X"03",X"2D",X"19",X"D6",X"02",X"C2",X"92",X"5D",X"E5",X"3A",X"72",X"23",X"D6",X"02",X"0F",X"47",
		X"3E",X"48",X"90",X"EB",X"CD",X"A9",X"5D",X"E1",X"C9",X"D5",X"D6",X"20",X"26",X"00",X"6F",X"29",
		X"29",X"29",X"01",X"02",X"0A",X"09",X"EB",X"06",X"08",X"CD",X"0A",X"0E",X"D1",X"C9",X"CD",X"89",
		X"5D",X"23",X"23",X"22",X"82",X"21",X"21",X"D0",X"5D",X"22",X"80",X"21",X"CD",X"1F",X"5E",X"C9",
		X"47",X"4F",X"4F",X"44",X"FF",X"42",X"41",X"44",X"FF",X"D5",X"CD",X"89",X"5D",X"23",X"23",X"22",
		X"82",X"21",X"21",X"D5",X"5D",X"22",X"80",X"21",X"CD",X"1F",X"5E",X"2A",X"82",X"21",X"23",X"22",
		X"82",X"21",X"EB",X"C1",X"78",X"0F",X"0F",X"0F",X"0F",X"CD",X"0D",X"5E",X"78",X"CD",X"0D",X"5E",
		X"79",X"0F",X"0F",X"0F",X"0F",X"CD",X"0D",X"5E",X"79",X"CD",X"0D",X"5E",X"C9",X"C5",X"E6",X"0F",
		X"C6",X"30",X"FE",X"3A",X"DA",X"19",X"5E",X"C6",X"07",X"CD",X"A9",X"5D",X"13",X"C1",X"C9",X"CD",
		X"77",X"0D",X"2A",X"80",X"21",X"7C",X"B5",X"C2",X"1F",X"5E",X"C9",X"EB",X"F9",X"11",X"00",X"24",
		X"06",X"40",X"21",X"00",X"00",X"39",X"0E",X"10",X"AF",X"29",X"DA",X"3E",X"5E",X"2F",X"12",X"13",
		X"3E",X"18",X"12",X"13",X"0D",X"C2",X"38",X"5E",X"05",X"C2",X"32",X"5E",X"C3",X"D2",X"5C",X"52",
		X"4F",X"4D",X"20",X"54",X"45",X"53",X"54",X"FF",X"AF",X"32",X"D0",X"21",X"32",X"A0",X"21",X"3E",
		X"0A",X"D3",X"00",X"21",X"00",X"20",X"01",X"E0",X"20",X"AF",X"77",X"23",X"0D",X"C2",X"6A",X"5E",
		X"05",X"C2",X"6A",X"5E",X"21",X"00",X"24",X"0E",X"1A",X"CD",X"92",X"5E",X"16",X"07",X"CD",X"A4",
		X"5E",X"15",X"C2",X"7E",X"5E",X"0D",X"C2",X"79",X"5E",X"CD",X"92",X"5E",X"00",X"00",X"00",X"C3",
		X"8C",X"5E",X"23",X"23",X"06",X"1B",X"3E",X"FF",X"77",X"23",X"05",X"C2",X"98",X"5E",X"36",X"01",
		X"23",X"23",X"23",X"C9",X"23",X"23",X"06",X"1C",X"3E",X"01",X"77",X"23",X"05",X"C2",X"AA",X"5E",
		X"23",X"23",X"C9",X"C9",X"C9",X"C9",X"C9",X"3E",X"00",X"C9",X"06",X"10",X"0E",X"09",X"C9",X"43",
		X"4F",X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"20",X"31",X"39",X"38",X"30",X"2C",X"20",X"44",
		X"41",X"56",X"45",X"20",X"4E",X"45",X"45",X"44",X"4C",X"45",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
