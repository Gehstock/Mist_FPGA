library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity satans_hollow_sp_bits_3 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of satans_hollow_sp_bits_3 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"76",X"00",
		X"00",X"00",X"76",X"00",X"00",X"00",X"76",X"00",X"00",X"00",X"76",X"00",X"00",X"DE",X"77",X"0D",
		X"00",X"DD",X"DD",X"77",X"00",X"77",X"66",X"07",X"00",X"7D",X"77",X"00",X"00",X"7D",X"76",X"00",
		X"00",X"7D",X"07",X"00",X"00",X"DE",X"00",X"00",X"00",X"DD",X"00",X"00",X"ED",X"66",X"E0",X"00",
		X"D7",X"66",X"D0",X"00",X"00",X"77",X"00",X"00",X"00",X"7D",X"00",X"00",X"00",X"7D",X"07",X"00",
		X"00",X"7D",X"76",X"00",X"00",X"DE",X"76",X"00",X"00",X"77",X"76",X"0D",X"00",X"77",X"76",X"77",
		X"00",X"7D",X"76",X"07",X"00",X"00",X"76",X"00",X"00",X"00",X"76",X"00",X"00",X"00",X"76",X"00",
		X"00",X"00",X"76",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"76",X"00",
		X"00",X"00",X"76",X"00",X"00",X"00",X"76",X"00",X"00",X"00",X"76",X"00",X"00",X"DE",X"77",X"0D",
		X"00",X"DD",X"DD",X"77",X"00",X"77",X"66",X"07",X"00",X"7D",X"77",X"00",X"00",X"7D",X"76",X"00",
		X"00",X"7D",X"07",X"00",X"00",X"DE",X"00",X"00",X"00",X"DD",X"00",X"00",X"DD",X"66",X"E0",X"00",
		X"77",X"66",X"D0",X"00",X"00",X"77",X"00",X"00",X"00",X"7D",X"00",X"00",X"00",X"7D",X"07",X"00",
		X"00",X"7D",X"76",X"00",X"00",X"DE",X"76",X"00",X"00",X"77",X"76",X"0D",X"00",X"77",X"76",X"77",
		X"00",X"7D",X"76",X"07",X"00",X"00",X"76",X"00",X"00",X"00",X"76",X"00",X"00",X"00",X"76",X"00",
		X"00",X"00",X"76",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"76",X"00",
		X"00",X"00",X"76",X"00",X"00",X"00",X"76",X"00",X"00",X"00",X"76",X"00",X"00",X"DE",X"77",X"0D",
		X"00",X"DD",X"DD",X"77",X"00",X"77",X"66",X"07",X"00",X"7D",X"77",X"00",X"00",X"7D",X"76",X"00",
		X"00",X"7D",X"07",X"00",X"00",X"DE",X"00",X"00",X"00",X"DD",X"00",X"00",X"ED",X"66",X"E0",X"00",
		X"D7",X"66",X"D0",X"00",X"00",X"77",X"00",X"00",X"00",X"7D",X"00",X"00",X"00",X"7D",X"07",X"00",
		X"00",X"7D",X"76",X"00",X"00",X"DE",X"76",X"00",X"00",X"77",X"76",X"0D",X"00",X"77",X"76",X"77",
		X"00",X"7D",X"76",X"07",X"00",X"00",X"76",X"00",X"00",X"00",X"76",X"00",X"00",X"00",X"76",X"00",
		X"00",X"00",X"76",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"76",X"00",
		X"00",X"00",X"76",X"00",X"00",X"00",X"76",X"00",X"00",X"00",X"76",X"00",X"00",X"DE",X"77",X"0D",
		X"DD",X"DD",X"DD",X"77",X"77",X"77",X"66",X"07",X"00",X"7D",X"77",X"00",X"00",X"7D",X"76",X"00",
		X"00",X"7D",X"07",X"00",X"00",X"DE",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"66",X"E0",X"00",
		X"00",X"66",X"D0",X"00",X"00",X"77",X"00",X"00",X"00",X"7D",X"00",X"00",X"00",X"7D",X"07",X"00",
		X"00",X"7D",X"76",X"00",X"00",X"DE",X"76",X"00",X"00",X"77",X"76",X"0D",X"00",X"77",X"76",X"77",
		X"00",X"7D",X"76",X"07",X"00",X"00",X"76",X"00",X"00",X"00",X"76",X"00",X"00",X"00",X"76",X"00",
		X"00",X"00",X"76",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"76",X"00",
		X"00",X"00",X"76",X"00",X"00",X"00",X"76",X"00",X"00",X"00",X"76",X"00",X"00",X"DE",X"77",X"0D",
		X"00",X"DD",X"DD",X"77",X"00",X"77",X"66",X"07",X"00",X"7D",X"77",X"00",X"00",X"7D",X"76",X"00",
		X"00",X"7D",X"07",X"00",X"00",X"DE",X"00",X"00",X"00",X"DD",X"00",X"00",X"ED",X"66",X"E0",X"00",
		X"D7",X"66",X"D0",X"00",X"00",X"77",X"00",X"00",X"00",X"7D",X"00",X"00",X"00",X"7D",X"07",X"00",
		X"00",X"7D",X"76",X"00",X"00",X"DE",X"76",X"00",X"00",X"77",X"76",X"0D",X"00",X"77",X"76",X"77",
		X"00",X"7D",X"76",X"07",X"00",X"00",X"76",X"00",X"00",X"00",X"76",X"00",X"00",X"00",X"76",X"00",
		X"00",X"00",X"76",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"76",X"00",
		X"00",X"00",X"76",X"00",X"00",X"00",X"76",X"00",X"00",X"00",X"76",X"00",X"00",X"DE",X"77",X"0D",
		X"ED",X"7D",X"DD",X"77",X"D7",X"77",X"66",X"07",X"00",X"7D",X"77",X"00",X"00",X"7D",X"76",X"00",
		X"00",X"7D",X"07",X"00",X"00",X"DE",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"66",X"E0",X"00",
		X"00",X"66",X"D0",X"00",X"00",X"77",X"00",X"00",X"00",X"7D",X"00",X"00",X"00",X"7D",X"07",X"00",
		X"00",X"7D",X"76",X"00",X"00",X"DE",X"76",X"00",X"ED",X"77",X"76",X"0D",X"D7",X"77",X"76",X"77",
		X"00",X"7D",X"76",X"07",X"00",X"00",X"76",X"00",X"00",X"00",X"76",X"00",X"00",X"00",X"76",X"00",
		X"00",X"00",X"76",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"10",X"00",X"00",X"44",X"10",X"00",X"00",X"23",X"31",X"00",X"00",X"31",X"10",X"01",
		X"00",X"31",X"11",X"14",X"11",X"32",X"14",X"14",X"3F",X"32",X"13",X"24",X"31",X"12",X"32",X"14",
		X"43",X"12",X"42",X"14",X"14",X"93",X"24",X"01",X"14",X"C9",X"22",X"00",X"14",X"93",X"22",X"00",
		X"43",X"13",X"24",X"00",X"31",X"32",X"42",X"10",X"3F",X"22",X"22",X"31",X"11",X"32",X"24",X"11",
		X"00",X"32",X"44",X"33",X"00",X"23",X"11",X"11",X"00",X"23",X"00",X"31",X"00",X"31",X"00",X"10",
		X"10",X"10",X"00",X"00",X"11",X"10",X"00",X"00",X"33",X"00",X"00",X"00",X"22",X"00",X"00",X"00",
		X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"C0",X"00",X"00",X"0C",X"99",X"00",X"00",X"CC",X"09",X"00",X"00",X"99",X"09",
		X"00",X"00",X"99",X"09",X"00",X"9F",X"99",X"09",X"00",X"C9",X"99",X"09",X"00",X"CC",X"90",X"09",
		X"00",X"C0",X"90",X"09",X"00",X"00",X"90",X"09",X"00",X"00",X"09",X"09",X"00",X"0F",X"C9",X"0C",
		X"00",X"0F",X"9F",X"CC",X"00",X"0F",X"FF",X"0C",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"09",
		X"00",X"CC",X"0F",X"99",X"00",X"C0",X"9F",X"0C",X"00",X"00",X"9F",X"0C",X"00",X"00",X"9F",X"0C",
		X"00",X"00",X"9F",X"00",X"00",X"00",X"FF",X"9F",X"00",X"0F",X"CC",X"F0",X"00",X"F9",X"99",X"00",
		X"00",X"99",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"CC",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"90",X"9F",X"00",X"00",X"9F",X"00",X"00",X"0F",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"09",X"00",
		X"00",X"99",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"09",X"09",X"09",X"99",X"99",
		X"99",X"99",X"99",X"99",X"96",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"00",
		X"96",X"99",X"99",X"00",X"99",X"99",X"99",X"99",X"09",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"09",X"99",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"FC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"0C",X"CC",X"00",X"00",X"0C",X"CC",X"00",
		X"00",X"0C",X"CC",X"00",X"00",X"0C",X"CC",X"00",X"00",X"0C",X"CC",X"00",X"00",X"0C",X"CC",X"00",
		X"00",X"0C",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"50",X"90",X"00",X"99",X"05",X"66",X"00",
		X"09",X"55",X"CC",X"00",X"05",X"59",X"CC",X"00",X"00",X"55",X"CC",X"00",X"00",X"F5",X"CC",X"00",
		X"5F",X"F0",X"CC",X"00",X"95",X"06",X"CC",X"00",X"00",X"66",X"C6",X"00",X"00",X"6C",X"66",X"00",
		X"00",X"CC",X"6C",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"66",X"00",X"00",X"C6",X"66",X"00",
		X"00",X"CC",X"6C",X"00",X"00",X"CC",X"66",X"00",X"00",X"6C",X"C6",X"00",X"00",X"66",X"66",X"00",
		X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",
		X"0B",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"C0",X"00",X"BB",X"BB",X"00",X"00",
		X"0B",X"BB",X"00",X"00",X"CC",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DD",X"9C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DD",X"90",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"92",X"00",
		X"44",X"00",X"99",X"00",X"94",X"00",X"92",X"99",X"14",X"99",X"22",X"00",X"94",X"29",X"99",X"00",
		X"44",X"22",X"99",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"99",X"00",X"00",X"92",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"29",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",
		X"99",X"99",X"00",X"00",X"BB",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"1B",X"B9",X"B0",X"00",
		X"00",X"BB",X"1B",X"00",X"09",X"BB",X"B1",X"00",X"99",X"B9",X"BB",X"00",X"1B",X"1B",X"1B",X"00",
		X"1A",X"11",X"B1",X"00",X"AA",X"11",X"BB",X"00",X"BA",X"C1",X"B1",X"90",X"BB",X"C1",X"BB",X"9B",
		X"BB",X"11",X"BB",X"1B",X"BB",X"11",X"1B",X"19",X"BB",X"99",X"11",X"19",X"BB",X"BB",X"11",X"19",
		X"BB",X"BB",X"1B",X"19",X"BB",X"1B",X"BB",X"1B",X"BB",X"C1",X"BB",X"9B",X"B9",X"C1",X"BB",X"90",
		X"BA",X"11",X"BB",X"00",X"AA",X"11",X"BB",X"00",X"1A",X"1B",X"1B",X"00",X"1B",X"BB",X"BB",X"00",
		X"9B",X"BB",X"BB",X"00",X"9B",X"BB",X"B0",X"00",X"09",X"B9",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"9A",X"9B",X"00",X"00",X"11",X"90",X"00",X"00",X"99",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"BA",
		X"00",X"00",X"00",X"BA",X"00",X"00",X"00",X"9A",X"00",X"00",X"00",X"9A",X"00",X"00",X"00",X"9A",
		X"00",X"00",X"00",X"BA",X"00",X"00",X"00",X"BA",X"FF",X"00",X"0B",X"0B",X"7F",X"00",X"9B",X"00",
		X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"91",X"00",X"90",X"00",X"91",X"00",
		X"99",X"00",X"91",X"00",X"79",X"77",X"99",X"00",X"FF",X"FF",X"99",X"00",X"90",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"F7",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"BB",X"99",X"00",X"09",X"BB",X"11",X"00",X"00",X"BB",X"11",X"00",X"00",X"BB",X"C1",
		X"00",X"00",X"BB",X"C1",X"00",X"00",X"AB",X"C1",X"00",X"00",X"AB",X"11",X"00",X"00",X"BB",X"11",
		X"00",X"00",X"19",X"11",X"00",X"00",X"99",X"1B",X"00",X"00",X"99",X"BB",X"00",X"00",X"B9",X"BB",
		X"00",X"00",X"9B",X"B9",X"00",X"00",X"BB",X"99",X"00",X"00",X"B9",X"99",X"00",X"00",X"B9",X"00",
		X"00",X"09",X"90",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"19",X"00",X"00",X"1B",X"19",X"00",X"00",X"BB",X"19",X"00",X"00",X"BB",X"19",X"00",X"00",
		X"BB",X"90",X"00",X"00",X"BB",X"00",X"00",X"00",X"9B",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",
		X"B1",X"00",X"00",X"00",X"1B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"99",X"88",X"88",X"88",X"99",X"88",X"88",X"F9",X"99",
		X"88",X"88",X"98",X"77",X"88",X"88",X"98",X"77",X"88",X"88",X"FF",X"97",X"88",X"88",X"F9",X"99",
		X"88",X"88",X"98",X"99",X"88",X"88",X"89",X"CC",X"88",X"88",X"88",X"CC",X"88",X"88",X"99",X"AA",
		X"88",X"88",X"99",X"CC",X"88",X"8F",X"79",X"CC",X"88",X"88",X"99",X"7C",X"88",X"88",X"F9",X"9C",
		X"88",X"88",X"88",X"AC",X"88",X"88",X"88",X"A9",X"88",X"88",X"88",X"9C",X"88",X"88",X"89",X"CC",
		X"88",X"88",X"99",X"CA",X"88",X"88",X"F9",X"9C",X"88",X"88",X"88",X"99",X"88",X"88",X"88",X"9A",
		X"88",X"88",X"F9",X"99",X"88",X"88",X"99",X"99",X"88",X"88",X"99",X"99",X"88",X"88",X"99",X"99",
		X"88",X"88",X"88",X"F9",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"00",X"B9",X"BB",X"99",X"00",X"BB",X"BB",X"11",X"00",X"9B",X"BB",X"11",X"00",X"BB",X"BB",X"C1",
		X"00",X"B9",X"BB",X"C1",X"00",X"BB",X"BB",X"C1",X"00",X"9B",X"BB",X"1B",X"00",X"BB",X"B9",X"1B",
		X"00",X"BB",X"B9",X"1B",X"00",X"BB",X"91",X"BB",X"00",X"9A",X"91",X"BB",X"00",X"AA",X"11",X"BB",
		X"00",X"AA",X"1C",X"B9",X"00",X"0B",X"C1",X"99",X"00",X"00",X"BB",X"99",X"00",X"00",X"B9",X"99",
		X"00",X"09",X"BB",X"91",X"00",X"99",X"00",X"99",X"00",X"BB",X"00",X"91",X"00",X"11",X"B0",X"99",
		X"00",X"99",X"B0",X"00",X"00",X"00",X"9B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"11",X"1B",X"00",X"91",X"C1",X"1B",X"00",X"19",X"11",X"BB",X"00",X"99",X"11",X"BB",X"00",
		X"91",X"11",X"B0",X"00",X"B1",X"C1",X"B0",X"00",X"BB",X"11",X"00",X"00",X"BB",X"11",X"00",X"00",
		X"B1",X"91",X"00",X"00",X"BB",X"1B",X"00",X"00",X"BB",X"10",X"00",X"00",X"BB",X"00",X"00",X"00",
		X"BB",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"1B",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"DD",X"D0",X"00",
		X"00",X"DD",X"EE",X"00",X"00",X"FD",X"EE",X"00",X"00",X"DD",X"EE",X"00",X"00",X"DD",X"EE",X"00",
		X"00",X"DD",X"EE",X"00",X"00",X"DD",X"EE",X"00",X"00",X"DD",X"EE",X"00",X"00",X"DD",X"DE",X"00",
		X"00",X"EE",X"EE",X"00",X"00",X"EE",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",
		X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",
		X"00",X"00",X"23",X"00",X"00",X"44",X"23",X"00",X"00",X"49",X"22",X"00",X"00",X"40",X"02",X"30",
		X"00",X"49",X"32",X"33",X"00",X"44",X"33",X"22",X"00",X"00",X"22",X"00",X"00",X"33",X"33",X"00",
		X"00",X"22",X"33",X"00",X"00",X"02",X"23",X"34",X"00",X"00",X"22",X"00",X"00",X"00",X"32",X"00",
		X"00",X"00",X"22",X"00",X"00",X"00",X"23",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",
		X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",
		X"00",X"02",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"23",X"00",X"00",X"00",X"33",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"99",X"CC",X"00",
		X"00",X"99",X"CC",X"00",X"00",X"CC",X"55",X"00",X"00",X"CC",X"55",X"00",X"00",X"00",X"50",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"5C",X"CC",X"00",X"00",X"5C",X"CC",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"C5",X"00",X"00",X"00",X"99",X"C0",X"00",X"00",X"99",X"C5",X"00",
		X"00",X"C9",X"05",X"00",X"00",X"5C",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"CC",X"CC",X"00",X"99",X"CC",X"CC",X"00",X"99",
		X"99",X"CC",X"00",X"00",X"99",X"CC",X"00",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"CC",X"55",X"55",X"00",X"CC",X"55",X"55",X"00",X"00",X"55",X"99",X"00",X"00",X"55",X"99",X"00",
		X"99",X"59",X"55",X"00",X"99",X"99",X"55",X"00",X"99",X"99",X"99",X"55",X"99",X"99",X"99",X"55",
		X"00",X"CC",X"CC",X"99",X"00",X"C9",X"CC",X"99",X"00",X"99",X"55",X"00",X"00",X"99",X"55",X"00",
		X"00",X"55",X"99",X"00",X"00",X"55",X"99",X"00",X"CC",X"55",X"00",X"00",X"CC",X"55",X"00",X"00",
		X"CC",X"55",X"00",X"00",X"CC",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"55",X"00",X"00",X"CC",X"55",X"00",X"00",X"CC",
		X"55",X"CC",X"00",X"55",X"55",X"CC",X"00",X"55",X"CC",X"55",X"CC",X"CC",X"CC",X"55",X"CC",X"CC",
		X"00",X"99",X"55",X"CC",X"00",X"99",X"55",X"CC",X"CC",X"99",X"55",X"CC",X"CC",X"99",X"55",X"CC",
		X"55",X"99",X"99",X"00",X"55",X"99",X"99",X"00",X"99",X"99",X"99",X"CC",X"99",X"F9",X"FF",X"CC",
		X"55",X"FF",X"F9",X"55",X"55",X"FF",X"99",X"55",X"55",X"99",X"99",X"CC",X"55",X"99",X"99",X"CC",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"55",X"99",X"99",X"CC",X"55",X"59",X"99",X"CC",
		X"00",X"55",X"99",X"55",X"00",X"55",X"99",X"55",X"CC",X"CC",X"55",X"CC",X"CC",X"CC",X"55",X"CC",
		X"CC",X"00",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"55",X"00",X"CC",X"00",X"55",X"00",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"90",X"FF",X"99",X"00",X"90",X"99",X"99",
		X"09",X"99",X"90",X"99",X"9F",X"00",X"99",X"90",X"9F",X"00",X"99",X"99",X"CC",X"00",X"99",X"99",
		X"CC",X"99",X"FF",X"00",X"99",X"9F",X"CC",X"CC",X"CC",X"99",X"CC",X"9C",X"CC",X"99",X"CC",X"99",
		X"CC",X"CC",X"CF",X"99",X"9F",X"FC",X"FF",X"00",X"FF",X"FF",X"99",X"00",X"99",X"CF",X"CC",X"90",
		X"99",X"99",X"99",X"99",X"99",X"CC",X"99",X"00",X"99",X"FF",X"99",X"00",X"99",X"99",X"00",X"00",
		X"00",X"99",X"00",X"90",X"00",X"99",X"00",X"99",X"00",X"90",X"00",X"99",X"00",X"99",X"00",X"09",
		X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"09",X"00",X"90",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"90",
		X"99",X"99",X"00",X"00",X"99",X"FF",X"99",X"00",X"99",X"CC",X"99",X"00",X"99",X"99",X"99",X"99",
		X"99",X"CF",X"CC",X"90",X"9F",X"F9",X"99",X"00",X"9F",X"FC",X"FF",X"00",X"9C",X"CC",X"CF",X"99",
		X"99",X"99",X"9C",X"99",X"CC",X"99",X"CC",X"9C",X"99",X"9F",X"CC",X"CC",X"CC",X"99",X"FF",X"00",
		X"99",X"90",X"99",X"99",X"9F",X"00",X"99",X"00",X"9F",X"00",X"99",X"00",X"09",X"99",X"90",X"90",
		X"00",X"90",X"99",X"90",X"00",X"90",X"FF",X"99",X"00",X"00",X"99",X"99",X"00",X"99",X"00",X"99",
		X"00",X"99",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"09",X"09",X"00",X"C9",X"09",X"99",X"90",X"09",X"99",X"00",X"90",X"90",X"09",X"09",X"99",
		X"99",X"90",X"CC",X"99",X"99",X"99",X"99",X"99",X"C9",X"09",X"99",X"90",X"C9",X"09",X"99",X"90",
		X"CC",X"09",X"09",X"F0",X"9C",X"99",X"09",X"FF",X"9C",X"99",X"00",X"0F",X"9C",X"CC",X"00",X"0F",
		X"0F",X"00",X"00",X"0F",X"09",X"00",X"00",X"99",X"09",X"00",X"00",X"99",X"99",X"00",X"00",X"99",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"90",X"99",X"00",X"00",X"F9",X"99",
		X"00",X"00",X"FF",X"99",X"00",X"00",X"CC",X"99",X"00",X"00",X"0C",X"F9",X"00",X"00",X"0C",X"F9",
		X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",
		X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"32",X"00",X"00",X"00",X"32",X"00",
		X"44",X"00",X"33",X"00",X"94",X"00",X"32",X"33",X"14",X"33",X"22",X"00",X"94",X"23",X"33",X"00",
		X"44",X"22",X"33",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"33",X"00",X"00",X"32",X"00",
		X"00",X"00",X"33",X"00",X"00",X"00",X"32",X"00",X"00",X"00",X"32",X"00",X"00",X"00",X"23",X"00",
		X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",
		X"00",X"00",X"30",X"00",X"00",X"40",X"33",X"00",X"00",X"93",X"33",X"00",X"00",X"13",X"33",X"00",
		X"00",X"93",X"23",X"00",X"00",X"40",X"23",X"00",X"00",X"00",X"23",X"00",X"00",X"00",X"23",X"00",
		X"00",X"20",X"33",X"00",X"00",X"22",X"23",X"00",X"00",X"33",X"22",X"00",X"00",X"03",X"22",X"00",
		X"00",X"00",X"22",X"00",X"00",X"00",X"32",X"00",X"00",X"00",X"33",X"00",X"00",X"22",X"33",X"30",
		X"00",X"23",X"33",X"30",X"00",X"33",X"23",X"30",X"22",X"32",X"33",X"04",X"00",X"22",X"33",X"00",
		X"00",X"33",X"33",X"00",X"00",X"33",X"33",X"00",X"00",X"33",X"33",X"00",X"00",X"00",X"33",X"00",
		X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"34",X"02",X"00",
		X"00",X"44",X"02",X"00",X"00",X"24",X"02",X"00",X"00",X"04",X"02",X"00",X"00",X"00",X"22",X"00",
		X"00",X"00",X"23",X"00",X"00",X"00",X"23",X"00",X"00",X"00",X"23",X"00",X"00",X"20",X"23",X"00",
		X"00",X"33",X"33",X"00",X"00",X"03",X"33",X"00",X"00",X"00",X"32",X"00",X"22",X"00",X"22",X"00",
		X"03",X"00",X"22",X"00",X"00",X"22",X"32",X"00",X"00",X"32",X"33",X"00",X"00",X"33",X"33",X"00",
		X"00",X"33",X"33",X"00",X"00",X"33",X"33",X"00",X"00",X"33",X"23",X"00",X"00",X"33",X"33",X"00",
		X"00",X"03",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"30",X"00",
		X"00",X"00",X"30",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"13",X"00",X"00",X"00",X"12",X"90",
		X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"30",X"00",
		X"00",X"20",X"30",X"00",X"00",X"32",X"30",X"00",X"00",X"33",X"30",X"00",X"00",X"33",X"30",X"00",
		X"00",X"33",X"33",X"00",X"00",X"33",X"33",X"00",X"00",X"03",X"33",X"00",X"00",X"03",X"33",X"00",
		X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",
		X"00",X"66",X"33",X"00",X"00",X"66",X"33",X"00",X"00",X"66",X"33",X"00",X"00",X"66",X"03",X"00",
		X"00",X"66",X"03",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"06",X"00",X"00",
		X"00",X"00",X"40",X"00",X"00",X"00",X"93",X"00",X"00",X"00",X"13",X"00",X"00",X"00",X"93",X"00",
		X"00",X"00",X"40",X"00",X"00",X"03",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"03",X"00",X"00",
		X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"32",X"00",X"00",
		X"00",X"32",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",
		X"00",X"23",X"00",X"00",X"00",X"23",X"00",X"00",X"00",X"23",X"00",X"00",X"00",X"02",X"00",X"00",
		X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"20",X"04",X"00",X"00",X"20",X"04",X"00",X"00",X"20",X"44",X"00",
		X"00",X"20",X"04",X"00",X"00",X"20",X"04",X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",
		X"00",X"20",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"32",X"02",X"00",X"00",X"32",X"23",X"00",
		X"00",X"32",X"33",X"00",X"00",X"32",X"33",X"00",X"00",X"32",X"30",X"00",X"00",X"32",X"30",X"00",
		X"00",X"32",X"00",X"00",X"00",X"32",X"00",X"00",X"00",X"32",X"06",X"00",X"00",X"33",X"66",X"00",
		X"00",X"33",X"66",X"00",X"00",X"33",X"66",X"00",X"00",X"33",X"66",X"00",X"00",X"33",X"60",X"00",
		X"00",X"33",X"66",X"00",X"00",X"33",X"60",X"00",X"00",X"33",X"66",X"00",X"00",X"33",X"66",X"00",
		X"00",X"33",X"60",X"00",X"00",X"33",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"03",X"99",X"00",X"00",X"30",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",
		X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"23",X"00",X"00",
		X"00",X"33",X"02",X"00",X"00",X"33",X"22",X"00",X"00",X"33",X"33",X"00",X"00",X"32",X"33",X"00",
		X"03",X"32",X"33",X"00",X"03",X"22",X"33",X"00",X"03",X"32",X"30",X"00",X"03",X"33",X"00",X"00",
		X"03",X"33",X"00",X"00",X"40",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",
		X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"32",X"00",X"00",X"00",X"32",X"00",X"00",
		X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"03",X"90",
		X"00",X"20",X"32",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",
		X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"22",X"00",X"00",X"03",X"23",X"00",X"00",
		X"03",X"33",X"00",X"00",X"33",X"33",X"00",X"00",X"33",X"33",X"00",X"00",X"33",X"32",X"00",X"00",
		X"33",X"22",X"22",X"00",X"33",X"22",X"33",X"00",X"00",X"22",X"33",X"20",X"00",X"22",X"22",X"00",
		X"00",X"23",X"33",X"00",X"00",X"23",X"33",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",
		X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0D",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0D",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",
		X"00",X"00",X"0C",X"F9",X"00",X"00",X"0C",X"F9",X"00",X"00",X"CC",X"F9",X"00",X"00",X"FF",X"C9",
		X"00",X"00",X"F9",X"C9",X"00",X"00",X"90",X"C9",X"00",X"00",X"00",X"C9",X"00",X"00",X"00",X"99",
		X"99",X"00",X"00",X"99",X"09",X"00",X"00",X"99",X"09",X"00",X"00",X"99",X"0F",X"00",X"00",X"0F",
		X"9C",X"CC",X"00",X"0F",X"9C",X"99",X"00",X"0F",X"9C",X"99",X"09",X"FF",X"C9",X"09",X"09",X"F0",
		X"C9",X"09",X"99",X"90",X"99",X"09",X"99",X"90",X"99",X"99",X"99",X"99",X"99",X"90",X"CC",X"09",
		X"90",X"09",X"09",X"99",X"09",X"99",X"99",X"90",X"C9",X"00",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"F0",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",
		X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",
		X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",
		X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"0F",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",
		X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"88",X"00",X"00",X"08",X"88",X"00",X"00",
		X"88",X"88",X"00",X"00",X"88",X"88",X"80",X"00",X"88",X"88",X"88",X"00",X"88",X"88",X"88",X"00",
		X"88",X"88",X"88",X"00",X"88",X"88",X"88",X"00",X"88",X"88",X"88",X"00",X"88",X"88",X"88",X"00",
		X"88",X"88",X"88",X"00",X"88",X"88",X"88",X"80",X"88",X"CC",X"88",X"88",X"88",X"99",X"88",X"88",
		X"88",X"CC",X"88",X"88",X"88",X"85",X"98",X"88",X"88",X"88",X"88",X"80",X"88",X"8C",X"88",X"00",
		X"88",X"98",X"88",X"00",X"88",X"89",X"88",X"00",X"88",X"58",X"88",X"00",X"88",X"C8",X"88",X"00",
		X"88",X"89",X"88",X"00",X"88",X"88",X"88",X"00",X"88",X"88",X"80",X"00",X"88",X"88",X"00",X"00",
		X"08",X"88",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"09",X"00",
		X"00",X"99",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"09",X"09",X"09",X"99",X"99",
		X"99",X"99",X"99",X"99",X"96",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"00",
		X"96",X"99",X"99",X"00",X"99",X"99",X"99",X"99",X"09",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"09",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"D0",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0C",X"00",X"00",X"00",X"9C",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"09",X"99",X"00",X"00",X"9F",X"00",X"00",X"00",X"C9",X"00",X"00",
		X"00",X"C9",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"0C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0C",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"9F",X"00",X"00",X"00",X"C9",X"99",X"00",
		X"00",X"C9",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"0C",X"90",X"00",
		X"00",X"00",X"C0",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"FF",X"50",X"00",X"00",X"5F",X"55",X"00",X"00",X"55",X"F5",X"00",X"00",
		X"05",X"FF",X"00",X"00",X"05",X"FF",X"00",X"00",X"00",X"5F",X"00",X"00",X"00",X"55",X"00",X"00",
		X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"90",X"00",X"00",X"40",X"99",X"00",X"00",X"93",X"99",X"00",X"00",X"13",X"99",X"00",
		X"00",X"93",X"29",X"00",X"00",X"40",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",
		X"00",X"20",X"99",X"00",X"00",X"22",X"29",X"00",X"00",X"99",X"22",X"00",X"00",X"09",X"22",X"00",
		X"00",X"00",X"22",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"99",X"00",X"00",X"22",X"99",X"90",
		X"00",X"29",X"99",X"90",X"00",X"99",X"29",X"90",X"22",X"92",X"99",X"04",X"00",X"22",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EF",X"00",X"00",X"00",X"EF",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"0E",X"FF",X"00",X"00",X"0E",X"FF",X"00",X"00",X"E0",X"EF",
		X"00",X"00",X"E0",X"EF",X"00",X"00",X"0E",X"EF",X"00",X"00",X"0E",X"EF",X"00",X"00",X"0F",X"EF",
		X"00",X"00",X"FF",X"EF",X"00",X"00",X"FF",X"EF",X"99",X"99",X"99",X"EF",X"00",X"00",X"F0",X"EF",
		X"00",X"00",X"FF",X"EF",X"00",X"00",X"FF",X"EF",X"00",X"00",X"EF",X"EF",X"00",X"00",X"E0",X"EF",
		X"00",X"00",X"00",X"EF",X"00",X"00",X"00",X"EF",X"00",X"00",X"E0",X"EF",X"00",X"00",X"E0",X"FF",
		X"00",X"00",X"EE",X"FF",X"00",X"00",X"0E",X"FF",X"00",X"00",X"00",X"EF",X"00",X"00",X"00",X"EF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"94",X"02",X"00",
		X"00",X"44",X"02",X"00",X"00",X"94",X"02",X"00",X"00",X"04",X"02",X"00",X"00",X"00",X"22",X"00",
		X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"20",X"29",X"00",
		X"00",X"99",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"92",X"00",X"22",X"00",X"22",X"00",
		X"09",X"00",X"22",X"00",X"00",X"22",X"92",X"00",X"00",X"92",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"99",X"00",
		X"00",X"09",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"12",X"90",
		X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",
		X"00",X"20",X"90",X"00",X"00",X"92",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"66",X"99",X"00",X"00",X"66",X"99",X"00",X"00",X"66",X"99",X"00",X"00",X"66",X"09",X"00",
		X"00",X"66",X"09",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"06",X"00",X"00",
		X"00",X"00",X"40",X"00",X"00",X"00",X"93",X"00",X"00",X"00",X"13",X"00",X"00",X"00",X"93",X"00",
		X"00",X"00",X"40",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"92",X"00",X"00",
		X"00",X"92",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"02",X"00",X"00",
		X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"20",X"04",X"00",X"00",X"20",X"04",X"00",X"00",X"20",X"44",X"00",
		X"00",X"20",X"04",X"00",X"00",X"20",X"04",X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",
		X"00",X"20",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"92",X"02",X"00",X"00",X"92",X"29",X"00",
		X"00",X"92",X"99",X"00",X"00",X"92",X"99",X"00",X"00",X"92",X"90",X"00",X"00",X"92",X"90",X"00",
		X"00",X"92",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"92",X"06",X"00",X"00",X"99",X"66",X"00",
		X"00",X"99",X"66",X"00",X"00",X"99",X"66",X"00",X"00",X"99",X"66",X"00",X"00",X"99",X"60",X"00",
		X"00",X"99",X"66",X"00",X"00",X"99",X"60",X"00",X"00",X"99",X"66",X"00",X"00",X"99",X"66",X"00",
		X"00",X"99",X"60",X"00",X"00",X"99",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"09",X"99",X"00",X"00",X"90",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",
		X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"29",X"00",X"00",
		X"00",X"99",X"02",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"99",X"00",X"00",X"92",X"99",X"00",
		X"09",X"92",X"99",X"00",X"09",X"22",X"99",X"00",X"09",X"92",X"90",X"00",X"09",X"99",X"00",X"00",
		X"09",X"99",X"00",X"00",X"40",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"92",X"00",X"00",
		X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"09",X"90",
		X"00",X"20",X"92",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",
		X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"22",X"00",X"00",X"09",X"29",X"00",X"00",
		X"09",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"92",X"00",X"00",
		X"99",X"22",X"22",X"00",X"99",X"22",X"99",X"00",X"00",X"22",X"99",X"20",X"00",X"22",X"29",X"00",
		X"00",X"29",X"99",X"00",X"00",X"29",X"99",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
