library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity cs50xx_prog is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of cs50xx_prog is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"68",X"40",X"50",X"1B",X"51",X"48",X"F0",X"55",X"5B",X"80",X"0D",X"04",X"5A",X"98",X"0F",X"0B",
		X"3F",X"04",X"D4",X"0D",X"21",X"01",X"08",X"0D",X"23",X"01",X"08",X"25",X"DE",X"DB",X"25",X"DE",
		X"14",X"0C",X"B0",X"D3",X"9F",X"21",X"01",X"23",X"01",X"55",X"51",X"1B",X"50",X"3E",X"04",X"3C",
		X"59",X"54",X"12",X"0A",X"55",X"80",X"13",X"55",X"0A",X"54",X"51",X"1B",X"50",X"3E",X"04",X"3C",
		X"58",X"80",X"90",X"1B",X"0A",X"C4",X"1B",X"71",X"B8",X"C3",X"3E",X"04",X"57",X"59",X"90",X"0B",
		X"08",X"3D",X"02",X"18",X"14",X"57",X"58",X"84",X"2E",X"DB",X"CC",X"72",X"04",X"57",X"90",X"59",
		X"0B",X"B0",X"E4",X"CC",X"08",X"3D",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"68",X"53",X"00",X"00",X"68",X"C0",X"00",X"00",X"69",X"02",X"00",X"00",X"69",X"0C",X"00",X"00",
		X"69",X"16",X"00",X"00",X"69",X"20",X"00",X"00",X"0D",X"69",X"30",X"00",X"0D",X"69",X"39",X"00",
		X"0D",X"69",X"3E",X"00",X"0D",X"69",X"4F",X"00",X"0D",X"69",X"60",X"00",X"0D",X"69",X"71",X"00",
		X"0D",X"69",X"82",X"00",X"0D",X"69",X"93",X"00",X"0D",X"69",X"A4",X"00",X"0D",X"69",X"B5",X"00",
		X"08",X"57",X"5A",X"80",X"90",X"0A",X"C5",X"5D",X"0A",X"C8",X"5E",X"0A",X"CB",X"5F",X"0A",X"CE",
		X"95",X"52",X"81",X"56",X"5B",X"81",X"64",X"E2",X"95",X"52",X"89",X"56",X"5B",X"81",X"64",X"E2",
		X"96",X"52",X"81",X"56",X"5B",X"89",X"64",X"E2",X"96",X"52",X"89",X"56",X"5B",X"89",X"64",X"E2",
		X"97",X"52",X"81",X"56",X"58",X"89",X"64",X"E2",X"97",X"52",X"89",X"56",X"58",X"89",X"64",X"E2",
		X"68",X"4C",X"93",X"52",X"56",X"81",X"56",X"65",X"30",X"57",X"68",X"4C",X"93",X"52",X"56",X"89",
		X"56",X"65",X"30",X"57",X"68",X"4C",X"90",X"52",X"56",X"89",X"56",X"65",X"30",X"57",X"68",X"4C",
		X"94",X"52",X"56",X"81",X"56",X"65",X"30",X"57",X"89",X"56",X"81",X"5C",X"64",X"E2",X"68",X"4C",
		X"08",X"57",X"5B",X"80",X"1D",X"88",X"1D",X"6C",X"3F",X"08",X"57",X"53",X"68",X"4C",X"08",X"57",
		X"5B",X"80",X"52",X"0D",X"77",X"04",X"52",X"5A",X"53",X"B0",X"69",X"C6",X"53",X"3D",X"08",X"08",
		X"57",X"5B",X"80",X"52",X"0D",X"76",X"04",X"52",X"5A",X"53",X"B0",X"69",X"C6",X"53",X"3D",X"08",
		X"08",X"57",X"5B",X"80",X"52",X"0D",X"75",X"04",X"52",X"5A",X"53",X"B0",X"69",X"C6",X"53",X"3D",
		X"08",X"08",X"57",X"5B",X"80",X"52",X"0D",X"77",X"04",X"52",X"5A",X"53",X"B0",X"69",X"C9",X"53",
		X"3D",X"09",X"08",X"57",X"5B",X"80",X"52",X"0D",X"76",X"04",X"52",X"5A",X"53",X"B0",X"69",X"C9",
		X"53",X"3D",X"09",X"08",X"57",X"5B",X"80",X"52",X"0D",X"75",X"04",X"52",X"5A",X"53",X"B0",X"69",
		X"C9",X"53",X"3D",X"09",X"08",X"57",X"5B",X"80",X"52",X"0D",X"77",X"04",X"52",X"5A",X"53",X"B0",
		X"69",X"CC",X"53",X"3D",X"0A",X"08",X"57",X"5B",X"80",X"52",X"0D",X"76",X"04",X"52",X"5A",X"53",
		X"B0",X"69",X"CC",X"53",X"3D",X"0A",X"53",X"3D",X"0D",X"53",X"3D",X"0E",X"53",X"3D",X"0F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"95",X"6A",X"EC",X"00",X"91",X"6A",X"EB",X"00",X"91",X"6A",X"D2",X"00",X"92",X"6A",X"EB",X"00",
		X"92",X"6A",X"D2",X"00",X"93",X"6A",X"EB",X"00",X"94",X"6A",X"EB",X"00",X"95",X"6A",X"EB",X"00",
		X"96",X"6A",X"EB",X"00",X"97",X"6A",X"EB",X"00",X"98",X"6A",X"EB",X"00",X"99",X"6A",X"EB",X"00",
		X"91",X"18",X"6A",X"EB",X"92",X"18",X"6A",X"EB",X"93",X"18",X"6A",X"EB",X"95",X"18",X"6A",X"EB",
		X"91",X"6A",X"EB",X"00",X"92",X"6A",X"EB",X"00",X"93",X"6A",X"EB",X"00",X"94",X"6A",X"EB",X"00",
		X"95",X"6A",X"EB",X"00",X"96",X"6A",X"EB",X"00",X"98",X"6A",X"EB",X"00",X"91",X"18",X"6A",X"EB",
		X"91",X"18",X"6A",X"C6",X"91",X"18",X"6A",X"CC",X"91",X"18",X"6A",X"D8",X"91",X"18",X"6A",X"E4",
		X"92",X"18",X"6A",X"EB",X"94",X"18",X"6A",X"EB",X"96",X"18",X"6A",X"EB",X"91",X"18",X"6A",X"EA",
		X"91",X"6A",X"D2",X"00",X"93",X"6A",X"EB",X"00",X"94",X"6A",X"D2",X"00",X"96",X"6A",X"EB",X"00",
		X"97",X"6A",X"D2",X"00",X"99",X"6A",X"EB",X"00",X"91",X"18",X"6A",X"C6",X"91",X"18",X"6A",X"D2",
		X"91",X"18",X"6A",X"E4",X"92",X"18",X"6A",X"C0",X"92",X"18",X"6A",X"CC",X"92",X"18",X"6A",X"DE",
		X"93",X"18",X"6A",X"EB",X"96",X"18",X"6A",X"EB",X"99",X"18",X"6A",X"EB",X"91",X"18",X"18",X"D2",
		X"0B",X"71",X"10",X"0B",X"18",X"ED",X"0B",X"72",X"10",X"0B",X"18",X"ED",X"0B",X"74",X"10",X"0B",
		X"18",X"ED",X"0B",X"75",X"10",X"0B",X"18",X"ED",X"0B",X"76",X"10",X"0B",X"18",X"ED",X"0B",X"77",
		X"10",X"0B",X"18",X"ED",X"0B",X"78",X"10",X"0B",X"18",X"ED",X"18",X"18",X"23",X"0E",X"F2",X"10",
		X"1A",X"F6",X"10",X"6B",X"0B",X"1A",X"0D",X"71",X"10",X"6B",X"0B",X"1A",X"14",X"23",X"0C",X"B0",
		X"6A",X"F6",X"08",X"99",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"95",X"1D",X"6C",X"3F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"95",X"6C",X"24",X"00",X"91",X"6C",X"23",X"00",X"91",X"6C",X"0C",X"00",X"92",X"6C",X"23",X"00",
		X"92",X"6C",X"0C",X"00",X"93",X"6C",X"23",X"00",X"94",X"6C",X"23",X"00",X"95",X"6C",X"23",X"00",
		X"96",X"6C",X"23",X"00",X"97",X"6C",X"23",X"00",X"98",X"6C",X"23",X"00",X"99",X"6C",X"23",X"00",
		X"91",X"18",X"6C",X"23",X"92",X"18",X"6C",X"23",X"93",X"18",X"6C",X"23",X"95",X"18",X"6C",X"23",
		X"91",X"6C",X"23",X"00",X"92",X"6C",X"23",X"00",X"93",X"6C",X"23",X"00",X"94",X"6C",X"23",X"00",
		X"95",X"6C",X"23",X"00",X"96",X"6C",X"23",X"00",X"98",X"6C",X"23",X"00",X"91",X"18",X"6C",X"23",
		X"91",X"18",X"6C",X"04",X"91",X"18",X"6C",X"08",X"91",X"18",X"6C",X"10",X"91",X"18",X"6C",X"18",
		X"92",X"18",X"6C",X"23",X"94",X"18",X"6C",X"23",X"96",X"18",X"6C",X"23",X"91",X"18",X"6C",X"22",
		X"91",X"6C",X"0C",X"00",X"93",X"6C",X"23",X"00",X"94",X"6C",X"0C",X"00",X"96",X"6C",X"23",X"00",
		X"97",X"6C",X"0C",X"00",X"99",X"6C",X"23",X"00",X"91",X"18",X"6C",X"04",X"91",X"18",X"6C",X"0C",
		X"91",X"18",X"6C",X"18",X"92",X"18",X"6C",X"00",X"92",X"18",X"6C",X"08",X"92",X"18",X"6C",X"14",
		X"93",X"18",X"6C",X"23",X"96",X"18",X"6C",X"23",X"99",X"18",X"6C",X"23",X"91",X"18",X"18",X"CC",
		X"0B",X"7F",X"DD",X"DB",X"0B",X"7E",X"DD",X"DB",X"0B",X"7C",X"DD",X"DB",X"0B",X"7B",X"DD",X"DB",
		X"0B",X"7A",X"DD",X"DB",X"0B",X"79",X"DD",X"DB",X"0B",X"78",X"DD",X"23",X"DE",X"21",X"11",X"0B",
		X"18",X"E5",X"18",X"18",X"23",X"1E",X"11",X"FC",X"1A",X"23",X"91",X"1E",X"11",X"FC",X"1A",X"14",
		X"23",X"0C",X"B0",X"E9",X"08",X"90",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"1D",X"6C",X"3F",X"94",
		X"52",X"5B",X"80",X"0D",X"04",X"56",X"04",X"08",X"5A",X"64",X"CD",X"5A",X"80",X"52",X"90",X"1D",
		X"88",X"1D",X"52",X"B0",X"6C",X"6A",X"56",X"33",X"94",X"52",X"08",X"94",X"52",X"56",X"81",X"56",
		X"64",X"E2",X"5C",X"94",X"52",X"89",X"56",X"81",X"64",X"E2",X"95",X"52",X"5B",X"80",X"0D",X"04",
		X"56",X"04",X"5D",X"0D",X"B0",X"6C",X"8B",X"08",X"5A",X"64",X"CD",X"B0",X"6C",X"8B",X"5A",X"56",
		X"32",X"95",X"52",X"14",X"77",X"04",X"56",X"5B",X"87",X"65",X"85",X"96",X"52",X"5B",X"80",X"0D",
		X"04",X"56",X"04",X"5E",X"0D",X"B0",X"EA",X"08",X"5A",X"64",X"CD",X"B0",X"EA",X"5A",X"56",X"31",
		X"96",X"52",X"14",X"77",X"04",X"56",X"5B",X"8F",X"65",X"85",X"97",X"52",X"5B",X"80",X"0D",X"04",
		X"56",X"04",X"5F",X"0D",X"B0",X"68",X"4C",X"08",X"5A",X"64",X"CD",X"B0",X"68",X"4C",X"5A",X"56",
		X"30",X"97",X"52",X"14",X"77",X"04",X"56",X"58",X"8F",X"65",X"85",X"68",X"4C",X"0D",X"1B",X"52",
		X"1B",X"2E",X"DC",X"1B",X"52",X"1B",X"08",X"14",X"0C",X"B0",X"CD",X"2C",X"90",X"28",X"E0",X"2C",
		X"91",X"2C",X"0D",X"1B",X"52",X"56",X"1B",X"0A",X"1B",X"52",X"56",X"1B",X"08",X"0D",X"1B",X"52",
		X"56",X"1B",X"0A",X"1B",X"52",X"56",X"1B",X"08",X"0D",X"1B",X"52",X"56",X"1B",X"0A",X"1B",X"52",
		X"56",X"1B",X"08",X"0D",X"1B",X"52",X"56",X"1B",X"0A",X"1B",X"52",X"56",X"1B",X"08",X"0D",X"1B",
		X"52",X"56",X"1B",X"0A",X"1B",X"52",X"56",X"1B",X"08",X"0D",X"1B",X"52",X"56",X"1B",X"0A",X"1B",
		X"52",X"56",X"1B",X"08",X"0D",X"1B",X"52",X"56",X"1B",X"0A",X"1B",X"52",X"56",X"1B",X"08",X"2C",
		X"0D",X"1B",X"52",X"56",X"1B",X"0A",X"1B",X"52",X"56",X"1B",X"90",X"0A",X"0D",X"1B",X"52",X"56",
		X"1B",X"0A",X"1B",X"52",X"56",X"1B",X"90",X"0A",X"0D",X"1B",X"52",X"56",X"1B",X"0A",X"1B",X"52",
		X"56",X"1B",X"90",X"0A",X"0D",X"1B",X"52",X"56",X"1B",X"0A",X"1B",X"52",X"56",X"1B",X"90",X"0A",
		X"0D",X"1B",X"52",X"56",X"1B",X"0A",X"1B",X"52",X"56",X"1B",X"90",X"0A",X"0D",X"1B",X"52",X"56",
		X"1B",X"0A",X"1B",X"52",X"56",X"1B",X"90",X"0A",X"0D",X"1B",X"52",X"56",X"1B",X"0A",X"1B",X"52",
		X"56",X"1B",X"90",X"0A",X"2C",X"0D",X"1B",X"52",X"56",X"1B",X"0E",X"CF",X"10",X"21",X"D0",X"10",
		X"1A",X"1B",X"52",X"56",X"1B",X"18",X"0D",X"1B",X"52",X"56",X"1B",X"0E",X"E0",X"10",X"21",X"E1",
		X"10",X"1A",X"1B",X"52",X"56",X"1B",X"18",X"0D",X"1B",X"52",X"56",X"1B",X"0E",X"F1",X"10",X"21",
		X"F2",X"10",X"1A",X"1B",X"52",X"56",X"1B",X"18",X"0D",X"1B",X"52",X"56",X"1B",X"0E",X"6D",X"C3",
		X"10",X"21",X"C4",X"10",X"1A",X"1B",X"52",X"56",X"1B",X"18",X"0D",X"1B",X"52",X"56",X"1B",X"0E",
		X"D4",X"10",X"21",X"D5",X"10",X"1A",X"1B",X"52",X"56",X"1B",X"18",X"0D",X"1B",X"52",X"56",X"1B",
		X"0E",X"E5",X"10",X"21",X"E6",X"10",X"1A",X"1B",X"52",X"56",X"1B",X"18",X"0D",X"1B",X"52",X"56",
		X"1B",X"0E",X"F6",X"10",X"21",X"F7",X"10",X"1A",X"90",X"0E",X"1D",X"1B",X"52",X"56",X"1B",X"18",
		X"2C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
