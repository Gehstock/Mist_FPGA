library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity time_pilot_sound_prog2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of time_pilot_sound_prog2 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"21",X"00",X"30",X"06",X"00",X"C3",X"7C",X"01",X"32",X"00",X"50",X"3A",X"00",X"40",X"C9",X"FF",
		X"32",X"00",X"70",X"3A",X"00",X"60",X"C9",X"FF",X"78",X"CF",X"79",X"32",X"00",X"40",X"C9",X"FF",
		X"78",X"D7",X"79",X"32",X"00",X"60",X"C9",X"FF",X"87",X"85",X"6F",X"7C",X"CE",X"00",X"67",X"7E",
		X"23",X"66",X"6F",X"E9",X"FF",X"FF",X"FF",X"FF",X"D9",X"08",X"CD",X"40",X"00",X"08",X"D9",X"C9",
		X"3E",X"0E",X"CF",X"B7",X"28",X"26",X"32",X"0B",X"30",X"CD",X"2D",X"01",X"3A",X"0B",X"30",X"CB",
		X"77",X"20",X"3F",X"3A",X"06",X"30",X"B7",X"3A",X"0B",X"30",X"C2",X"E6",X"00",X"21",X"06",X"30",
		X"36",X"00",X"B7",X"F2",X"FE",X"00",X"CB",X"BF",X"CD",X"89",X"00",X"C9",X"21",X"00",X"30",X"06",
		X"04",X"AF",X"77",X"23",X"10",X"FC",X"C9",X"21",X"00",X"30",X"06",X"02",X"0E",X"03",X"BE",X"28",
		X"05",X"23",X"23",X"10",X"F9",X"41",X"79",X"90",X"C9",X"CD",X"77",X"00",X"C8",X"AF",X"77",X"23",
		X"77",X"C9",X"3A",X"06",X"30",X"B7",X"20",X"27",X"3A",X"09",X"30",X"2A",X"07",X"30",X"BD",X"D8",
		X"BC",X"D8",X"3E",X"FF",X"32",X"06",X"30",X"06",X"00",X"21",X"00",X"30",X"3A",X"0B",X"30",X"77",
		X"23",X"70",X"23",X"70",X"23",X"70",X"3E",X"01",X"32",X"04",X"30",X"CD",X"BE",X"02",X"C9",X"3A",
		X"0B",X"30",X"CB",X"B7",X"CD",X"77",X"00",X"28",X"04",X"23",X"36",X"00",X"C9",X"3A",X"09",X"30",
		X"47",X"3A",X"07",X"30",X"B8",X"D0",X"21",X"00",X"30",X"3A",X"0B",X"30",X"77",X"23",X"36",X"00",
		X"3E",X"FF",X"32",X"06",X"30",X"C9",X"3A",X"09",X"30",X"47",X"3A",X"07",X"30",X"B8",X"D0",X"AF",
		X"32",X"06",X"30",X"3A",X"0B",X"30",X"21",X"00",X"30",X"77",X"23",X"36",X"00",X"C9",X"32",X"0B",
		X"30",X"CD",X"77",X"00",X"28",X"04",X"23",X"36",X"00",X"C9",X"AF",X"CD",X"77",X"00",X"28",X"08",
		X"3A",X"0B",X"30",X"77",X"23",X"36",X"00",X"C9",X"CD",X"2D",X"01",X"21",X"00",X"30",X"B7",X"C8",
		X"3D",X"87",X"4F",X"06",X"00",X"09",X"3A",X"0B",X"30",X"77",X"23",X"70",X"C9",X"3A",X"00",X"30",
		X"CD",X"4F",X"01",X"32",X"07",X"30",X"3A",X"02",X"30",X"CD",X"4F",X"01",X"32",X"08",X"30",X"3A",
		X"0B",X"30",X"CD",X"4F",X"01",X"32",X"09",X"30",X"CD",X"61",X"01",X"32",X"0A",X"30",X"C9",X"21",
		X"AD",X"05",X"CB",X"77",X"28",X"05",X"CB",X"B7",X"21",X"AD",X"05",X"06",X"00",X"4F",X"09",X"7E",
		X"C9",X"2A",X"07",X"30",X"7C",X"BD",X"38",X"09",X"3A",X"09",X"30",X"BD",X"38",X"0C",X"3E",X"01",
		X"C9",X"3A",X"09",X"30",X"BC",X"38",X"03",X"3E",X"02",X"C9",X"AF",X"C9",X"70",X"23",X"7C",X"FE",
		X"34",X"20",X"F9",X"F9",X"ED",X"56",X"21",X"00",X"80",X"22",X"0C",X"30",X"77",X"01",X"3F",X"07",
		X"DF",X"E7",X"32",X"0E",X"30",X"32",X"0F",X"30",X"CD",X"A2",X"02",X"CD",X"A6",X"02",X"CD",X"AA",
		X"02",X"CD",X"B0",X"02",X"CD",X"B4",X"02",X"CD",X"B8",X"02",X"3A",X"06",X"30",X"B7",X"28",X"06",
		X"FB",X"00",X"00",X"F3",X"18",X"0F",X"FB",X"3E",X"0F",X"CF",X"E6",X"40",X"20",X"F9",X"3E",X"0F",
		X"CF",X"E6",X"40",X"28",X"F9",X"F3",X"3A",X"06",X"30",X"B7",X"20",X"2E",X"3E",X"00",X"32",X"04",
		X"30",X"3A",X"01",X"30",X"B7",X"3A",X"00",X"30",X"28",X"05",X"CD",X"85",X"02",X"18",X"03",X"CD",
		X"68",X"02",X"3E",X"01",X"32",X"04",X"30",X"3A",X"03",X"30",X"B7",X"3A",X"02",X"30",X"28",X"05",
		X"CD",X"85",X"02",X"18",X"B5",X"CD",X"68",X"02",X"18",X"B0",X"3E",X"00",X"32",X"04",X"30",X"3A",
		X"01",X"30",X"B7",X"3A",X"00",X"30",X"28",X"05",X"CD",X"3C",X"02",X"18",X"9D",X"CD",X"12",X"02",
		X"18",X"98",X"CB",X"B7",X"32",X"00",X"30",X"CD",X"BE",X"02",X"3A",X"00",X"30",X"21",X"F9",X"04",
		X"EF",X"B7",X"20",X"6B",X"21",X"01",X"30",X"36",X"01",X"11",X"53",X"05",X"3A",X"00",X"30",X"6F",
		X"26",X"00",X"29",X"19",X"5E",X"23",X"56",X"ED",X"53",X"10",X"30",X"C9",X"B7",X"C8",X"2A",X"10",
		X"30",X"CD",X"33",X"00",X"B7",X"C8",X"21",X"00",X"30",X"3D",X"28",X"06",X"36",X"00",X"AF",X"32",
		X"06",X"30",X"23",X"36",X"00",X"C9",X"B7",X"C8",X"E6",X"03",X"C5",X"47",X"3A",X"04",X"30",X"4F",
		X"87",X"81",X"80",X"32",X"05",X"30",X"C1",X"C9",X"F5",X"CD",X"BE",X"02",X"F1",X"E6",X"3F",X"21",
		X"F9",X"04",X"EF",X"B7",X"C2",X"8F",X"02",X"21",X"01",X"30",X"3A",X"04",X"30",X"87",X"5F",X"16",
		X"00",X"19",X"36",X"01",X"C9",X"B7",X"C8",X"E6",X"3F",X"21",X"53",X"05",X"EF",X"B7",X"C8",X"57",
		X"21",X"00",X"30",X"3A",X"04",X"30",X"4F",X"06",X"00",X"09",X"09",X"15",X"28",X"01",X"70",X"23",
		X"70",X"C9",X"06",X"08",X"18",X"06",X"06",X"09",X"18",X"02",X"06",X"0A",X"0E",X"00",X"DF",X"C9",
		X"06",X"08",X"18",X"06",X"06",X"09",X"18",X"02",X"06",X"0A",X"0E",X"00",X"E7",X"C9",X"01",X"00",
		X"08",X"3A",X"04",X"30",X"B7",X"20",X"0C",X"DF",X"04",X"DF",X"04",X"DF",X"0E",X"3F",X"CD",X"2D",
		X"03",X"AF",X"C9",X"E7",X"04",X"E7",X"04",X"E7",X"0E",X"3F",X"CD",X"39",X"03",X"AF",X"C9",X"CD",
		X"56",X"02",X"3A",X"05",X"30",X"3D",X"21",X"EB",X"02",X"EF",X"C9",X"F7",X"02",X"00",X"03",X"09",
		X"03",X"12",X"03",X"1B",X"03",X"24",X"03",X"CD",X"A2",X"02",X"0E",X"09",X"CD",X"2D",X"03",X"C9",
		X"CD",X"A6",X"02",X"0E",X"12",X"CD",X"2D",X"03",X"C9",X"CD",X"AA",X"02",X"0E",X"24",X"CD",X"2D",
		X"03",X"C9",X"CD",X"B0",X"02",X"0E",X"09",X"CD",X"39",X"03",X"C9",X"CD",X"B4",X"02",X"0E",X"12",
		X"CD",X"39",X"03",X"C9",X"CD",X"B8",X"02",X"0E",X"24",X"CD",X"39",X"03",X"C9",X"3A",X"0E",X"30",
		X"B1",X"32",X"0E",X"30",X"06",X"07",X"4F",X"DF",X"C9",X"3A",X"0F",X"30",X"B1",X"32",X"0F",X"30",
		X"06",X"07",X"4F",X"E7",X"C9",X"06",X"06",X"3A",X"04",X"30",X"B7",X"20",X"02",X"DF",X"C9",X"E7",
		X"C9",X"06",X"06",X"3A",X"04",X"30",X"B7",X"20",X"04",X"78",X"CF",X"4F",X"C9",X"78",X"D7",X"4F",
		X"C9",X"3A",X"0E",X"30",X"A0",X"B1",X"32",X"0E",X"30",X"4F",X"06",X"07",X"DF",X"C9",X"3A",X"0F",
		X"30",X"A0",X"B1",X"32",X"0F",X"30",X"4F",X"06",X"07",X"E7",X"C9",X"21",X"91",X"03",X"3D",X"87",
		X"5F",X"16",X"00",X"19",X"5E",X"23",X"56",X"4B",X"42",X"3A",X"04",X"30",X"B7",X"28",X"D2",X"18",
		X"DD",X"08",X"FE",X"10",X"FD",X"20",X"FB",X"21",X"AD",X"03",X"3D",X"87",X"5F",X"16",X"00",X"19",
		X"5E",X"23",X"56",X"4B",X"42",X"3A",X"04",X"30",X"B7",X"28",X"B6",X"18",X"C1",X"01",X"F7",X"02",
		X"EF",X"04",X"DF",X"21",X"C9",X"03",X"3D",X"87",X"5F",X"16",X"00",X"19",X"5E",X"23",X"56",X"4B",
		X"42",X"3A",X"04",X"30",X"B7",X"28",X"9A",X"18",X"A5",X"00",X"F6",X"00",X"ED",X"00",X"DB",X"21",
		X"E7",X"03",X"3D",X"87",X"5F",X"16",X"00",X"19",X"5E",X"23",X"56",X"4B",X"42",X"3A",X"04",X"30",
		X"B7",X"CA",X"61",X"03",X"C3",X"6E",X"03",X"09",X"FF",X"12",X"FF",X"24",X"FF",X"C6",X"07",X"47",
		X"3A",X"04",X"30",X"B7",X"20",X"02",X"DF",X"C9",X"E7",X"C9",X"C6",X"07",X"47",X"3A",X"04",X"30",
		X"B7",X"78",X"20",X"02",X"CF",X"C9",X"D7",X"C9",X"3D",X"87",X"47",X"4D",X"3A",X"04",X"30",X"B7",
		X"20",X"05",X"DF",X"4C",X"04",X"DF",X"C9",X"E7",X"4C",X"04",X"E7",X"C9",X"3D",X"87",X"67",X"3A",
		X"04",X"30",X"B7",X"7C",X"20",X"07",X"CF",X"6F",X"7C",X"3C",X"CF",X"67",X"C9",X"D7",X"6F",X"7C",
		X"3C",X"D7",X"67",X"C9",X"CD",X"56",X"02",X"7D",X"FE",X"04",X"D0",X"F5",X"21",X"83",X"04",X"3A",
		X"05",X"30",X"3D",X"87",X"5F",X"16",X"00",X"19",X"5E",X"23",X"56",X"2A",X"0C",X"30",X"7B",X"A5",
		X"6F",X"7A",X"A4",X"67",X"22",X"0C",X"30",X"F1",X"B7",X"20",X"02",X"77",X"C9",X"21",X"83",X"04",
		X"87",X"87",X"4F",X"87",X"81",X"4F",X"06",X"00",X"09",X"3A",X"05",X"30",X"3D",X"87",X"5F",X"16",
		X"00",X"19",X"5E",X"23",X"56",X"2A",X"0C",X"30",X"7B",X"B5",X"6F",X"7A",X"B4",X"67",X"22",X"0C",
		X"30",X"77",X"C9",X"3F",X"FF",X"FF",X"FC",X"FF",X"F3",X"FC",X"FF",X"F3",X"FF",X"CF",X"FF",X"80",
		X"00",X"00",X"02",X"00",X"08",X"02",X"00",X"08",X"00",X"20",X"00",X"40",X"00",X"00",X"01",X"00",
		X"04",X"01",X"00",X"04",X"00",X"10",X"00",X"C0",X"00",X"00",X"03",X"00",X"0C",X"03",X"00",X"0C",
		X"00",X"30",X"00",X"0E",X"10",X"C6",X"07",X"47",X"3A",X"04",X"30",X"B7",X"20",X"02",X"DF",X"C9",
		X"E7",X"C9",X"06",X"0B",X"4D",X"3A",X"04",X"30",X"B7",X"20",X"05",X"DF",X"04",X"4C",X"DF",X"C9",
		X"E7",X"04",X"4C",X"E7",X"C9",X"3A",X"04",X"30",X"B7",X"3E",X"0B",X"47",X"20",X"07",X"CF",X"6F",
		X"78",X"3C",X"CF",X"67",X"C9",X"D7",X"6F",X"78",X"3C",X"D7",X"67",X"C9",X"4F",X"06",X"0D",X"3A",
		X"04",X"30",X"B7",X"20",X"02",X"DF",X"C9",X"E7",X"C9",X"BE",X"02",X"B0",X"0F",X"7D",X"0F",X"8E",
		X"0F",X"5A",X"10",X"F4",X"0F",X"DA",X"05",X"08",X"17",X"DA",X"05",X"82",X"1B",X"99",X"16",X"D2",
		X"0F",X"2F",X"16",X"76",X"17",X"DA",X"05",X"27",X"1B",X"B6",X"1D",X"DA",X"05",X"9D",X"1C",X"DA",
		X"05",X"DA",X"05",X"2A",X"1C",X"DA",X"05",X"DA",X"05",X"DA",X"05",X"DA",X"05",X"DA",X"05",X"05",
		X"10",X"16",X"10",X"9F",X"0F",X"DA",X"05",X"DA",X"05",X"DA",X"05",X"27",X"10",X"38",X"10",X"49",
		X"10",X"DA",X"05",X"C1",X"0F",X"DA",X"05",X"DA",X"05",X"DA",X"05",X"DA",X"05",X"DA",X"05",X"DA",
		X"05",X"48",X"1D",X"00",X"00",X"BD",X"0F",X"8A",X"0F",X"9B",X"0F",X"67",X"10",X"01",X"10",X"DD",
		X"05",X"3B",X"17",X"DD",X"05",X"BE",X"1B",X"CB",X"16",X"DF",X"0F",X"62",X"16",X"8E",X"17",X"DD",
		X"05",X"44",X"1B",X"F0",X"1D",X"DD",X"05",X"D5",X"1C",X"DD",X"05",X"DD",X"05",X"55",X"1C",X"DD",
		X"05",X"DD",X"05",X"DD",X"05",X"DD",X"05",X"DD",X"05",X"12",X"10",X"23",X"10",X"AC",X"0F",X"DD",
		X"05",X"DD",X"05",X"DD",X"05",X"34",X"10",X"45",X"10",X"56",X"10",X"DD",X"05",X"CE",X"0F",X"DD",
		X"05",X"DD",X"05",X"DD",X"05",X"DD",X"05",X"DD",X"05",X"DD",X"05",X"6F",X"1D",X"00",X"98",X"A0",
		X"A8",X"D8",X"60",X"00",X"EC",X"00",X"B0",X"78",X"F0",X"C0",X"E8",X"00",X"B2",X"00",X"00",X"E0",
		X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"70",X"68",X"B8",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"C8",X"3E",X"00",X"C9",X"3E",X"FF",X"C9",
		X"DD",X"7E",X"00",X"FE",X"FF",X"C8",X"DD",X"36",X"09",X"01",X"CD",X"4C",X"06",X"AF",X"C9",X"DD",
		X"7E",X"00",X"FE",X"FF",X"28",X"09",X"DD",X"36",X"09",X"02",X"CD",X"4C",X"06",X"AF",X"C9",X"0E",
		X"00",X"3E",X"02",X"CD",X"ED",X"03",X"3E",X"FF",X"C9",X"DD",X"7E",X"00",X"FE",X"FF",X"28",X"09",
		X"DD",X"36",X"09",X"03",X"CD",X"4C",X"06",X"AF",X"C9",X"0E",X"00",X"3E",X"03",X"CD",X"ED",X"03",
		X"3E",X"FF",X"C9",X"DD",X"7E",X"0A",X"FE",X"FF",X"C8",X"DD",X"36",X"09",X"04",X"CD",X"72",X"07",
		X"AF",X"C9",X"DD",X"7E",X"0A",X"FE",X"FF",X"C8",X"DD",X"36",X"09",X"05",X"CD",X"72",X"07",X"AF",
		X"C9",X"DD",X"7E",X"00",X"FE",X"FF",X"C8",X"CD",X"3E",X"08",X"AF",X"C9",X"DD",X"35",X"01",X"C0",
		X"3A",X"48",X"30",X"DD",X"77",X"01",X"DD",X"CB",X"00",X"46",X"C2",X"6F",X"06",X"DD",X"7E",X"07",
		X"D6",X"01",X"FA",X"6F",X"06",X"DD",X"77",X"07",X"4F",X"DD",X"7E",X"09",X"CD",X"ED",X"03",X"DD",
		X"35",X"00",X"C0",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"7E",X"47",X"E6",X"1F",X"CA",X"37",X"07",
		X"FE",X"1F",X"C2",X"45",X"07",X"23",X"DD",X"75",X"02",X"DD",X"74",X"03",X"78",X"E6",X"E0",X"0F",
		X"0F",X"0F",X"0F",X"4F",X"06",X"00",X"21",X"9F",X"06",X"09",X"5E",X"23",X"56",X"EB",X"E9",X"AF",
		X"06",X"E5",X"06",X"07",X"07",X"FB",X"06",X"2A",X"07",X"2A",X"07",X"2A",X"07",X"2A",X"07",X"DD",
		X"6E",X"02",X"DD",X"66",X"03",X"4E",X"CB",X"21",X"06",X"00",X"21",X"34",X"09",X"09",X"5E",X"23",
		X"56",X"ED",X"53",X"44",X"30",X"DD",X"73",X"04",X"DD",X"72",X"05",X"DD",X"6E",X"02",X"DD",X"66",
		X"03",X"4E",X"CB",X"21",X"06",X"00",X"21",X"60",X"09",X"09",X"5E",X"23",X"56",X"DD",X"73",X"0B",
		X"DD",X"72",X"0C",X"18",X"35",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"4E",X"06",X"00",X"21",X"7C",
		X"0A",X"09",X"7E",X"32",X"48",X"30",X"DD",X"77",X"01",X"18",X"1F",X"DD",X"6E",X"02",X"DD",X"66",
		X"03",X"7E",X"DD",X"77",X"08",X"18",X"13",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"7E",X"DD",X"77",
		X"06",X"DD",X"77",X"07",X"DD",X"77",X"0D",X"DD",X"77",X"0E",X"DD",X"6E",X"02",X"DD",X"66",X"03",
		X"23",X"DD",X"75",X"02",X"DD",X"74",X"03",X"C3",X"73",X"06",X"DD",X"7E",X"09",X"0E",X"00",X"CD",
		X"ED",X"03",X"DD",X"36",X"00",X"FF",X"C9",X"CD",X"02",X"09",X"DD",X"7E",X"09",X"0E",X"00",X"CD",
		X"ED",X"03",X"C3",X"26",X"09",X"C5",X"CD",X"02",X"09",X"C1",X"78",X"E6",X"1F",X"3D",X"07",X"4F",
		X"06",X"00",X"DD",X"6E",X"04",X"DD",X"66",X"05",X"09",X"5E",X"23",X"56",X"EB",X"DD",X"7E",X"09",
		X"CD",X"08",X"04",X"DD",X"4E",X"06",X"DD",X"71",X"07",X"DD",X"7E",X"09",X"CD",X"ED",X"03",X"C3",
		X"26",X"09",X"DD",X"35",X"0F",X"C0",X"3A",X"48",X"30",X"DD",X"77",X"0F",X"DD",X"CB",X"0A",X"46",
		X"C2",X"A5",X"07",X"DD",X"7E",X"0E",X"D6",X"01",X"FA",X"A5",X"07",X"DD",X"77",X"0E",X"DD",X"7E",
		X"09",X"FE",X"04",X"28",X"08",X"DD",X"4E",X"0E",X"3E",X"02",X"CD",X"ED",X"03",X"DD",X"4E",X"0E",
		X"3E",X"03",X"CD",X"ED",X"03",X"DD",X"35",X"0A",X"C0",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"2B",
		X"7E",X"47",X"E6",X"1F",X"28",X"1E",X"FE",X"1F",X"20",X"33",X"DD",X"7E",X"09",X"FE",X"04",X"28",
		X"07",X"3E",X"02",X"0E",X"00",X"CD",X"ED",X"03",X"3E",X"03",X"0E",X"00",X"CD",X"ED",X"03",X"DD",
		X"36",X"0A",X"FF",X"C9",X"CD",X"14",X"09",X"DD",X"7E",X"09",X"FE",X"04",X"28",X"07",X"3E",X"02",
		X"0E",X"00",X"CD",X"ED",X"03",X"3E",X"03",X"0E",X"00",X"CD",X"ED",X"03",X"C9",X"C5",X"CD",X"14",
		X"09",X"C1",X"78",X"E6",X"1F",X"3D",X"07",X"4F",X"06",X"00",X"DD",X"7E",X"09",X"FE",X"04",X"28",
		X"12",X"DD",X"6E",X"04",X"DD",X"66",X"05",X"09",X"5E",X"23",X"56",X"EB",X"C5",X"3E",X"02",X"CD",
		X"08",X"04",X"C1",X"DD",X"6E",X"0B",X"DD",X"66",X"0C",X"09",X"5E",X"23",X"56",X"EB",X"3E",X"03",
		X"CD",X"08",X"04",X"DD",X"4E",X"0D",X"DD",X"71",X"0E",X"DD",X"7E",X"09",X"FE",X"04",X"28",X"05",
		X"3E",X"02",X"CD",X"ED",X"03",X"3E",X"03",X"DD",X"4E",X"0D",X"CD",X"ED",X"03",X"C9",X"DD",X"35",
		X"01",X"C0",X"3A",X"48",X"30",X"DD",X"77",X"01",X"DD",X"CB",X"00",X"46",X"C2",X"5A",X"08",X"DD",
		X"7E",X"07",X"D6",X"01",X"FA",X"5A",X"08",X"DD",X"77",X"07",X"DD",X"35",X"00",X"C0",X"DD",X"6E",
		X"02",X"DD",X"66",X"03",X"7E",X"47",X"E6",X"1F",X"CA",X"F0",X"08",X"FE",X"1F",X"C2",X"F6",X"08",
		X"23",X"DD",X"75",X"02",X"DD",X"74",X"03",X"78",X"E6",X"E0",X"0F",X"0F",X"0F",X"0F",X"4F",X"06",
		X"00",X"21",X"8A",X"08",X"09",X"5E",X"23",X"56",X"EB",X"E9",X"9A",X"08",X"B8",X"08",X"CE",X"08",
		X"EB",X"08",X"EB",X"08",X"EB",X"08",X"EB",X"08",X"EB",X"08",X"DD",X"6E",X"02",X"DD",X"66",X"03",
		X"4E",X"CB",X"21",X"06",X"00",X"21",X"34",X"09",X"09",X"5E",X"23",X"56",X"ED",X"53",X"44",X"30",
		X"DD",X"73",X"04",X"DD",X"72",X"05",X"18",X"23",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"4E",X"06",
		X"00",X"21",X"7C",X"0A",X"09",X"7E",X"32",X"48",X"30",X"DD",X"77",X"01",X"18",X"0D",X"DD",X"6E",
		X"02",X"DD",X"66",X"03",X"7E",X"DD",X"77",X"06",X"DD",X"77",X"07",X"DD",X"6E",X"02",X"DD",X"66",
		X"03",X"23",X"DD",X"75",X"02",X"DD",X"74",X"03",X"C3",X"5E",X"08",X"DD",X"36",X"00",X"FF",X"C9",
		X"CD",X"02",X"09",X"C3",X"26",X"09",X"CD",X"02",X"09",X"DD",X"4E",X"06",X"DD",X"71",X"07",X"C3",
		X"26",X"09",X"78",X"E6",X"E0",X"07",X"07",X"07",X"47",X"3E",X"01",X"18",X"01",X"07",X"10",X"FD",
		X"DD",X"77",X"00",X"C9",X"78",X"E6",X"E0",X"07",X"07",X"07",X"47",X"3E",X"01",X"18",X"01",X"07",
		X"10",X"FD",X"DD",X"77",X"0A",X"C9",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"23",X"DD",X"75",X"02",
		X"DD",X"74",X"03",X"C9",X"8C",X"09",X"90",X"09",X"94",X"09",X"98",X"09",X"9C",X"09",X"A0",X"09",
		X"A4",X"09",X"A8",X"09",X"AC",X"09",X"B0",X"09",X"B4",X"09",X"B8",X"09",X"BC",X"09",X"C0",X"09",
		X"C4",X"09",X"C8",X"09",X"CC",X"09",X"D0",X"09",X"D4",X"09",X"D8",X"09",X"DC",X"09",X"E0",X"09",
		X"04",X"0A",X"08",X"0A",X"0C",X"0A",X"10",X"0A",X"14",X"0A",X"18",X"0A",X"1C",X"0A",X"20",X"0A",
		X"24",X"0A",X"28",X"0A",X"2C",X"0A",X"30",X"0A",X"34",X"0A",X"38",X"0A",X"3C",X"0A",X"40",X"0A",
		X"44",X"0A",X"48",X"0A",X"4C",X"0A",X"50",X"0A",X"54",X"0A",X"58",X"0A",X"6B",X"08",X"F2",X"07",
		X"80",X"07",X"14",X"07",X"AE",X"06",X"4E",X"06",X"F3",X"05",X"9E",X"05",X"4E",X"05",X"01",X"05",
		X"B9",X"04",X"76",X"04",X"36",X"04",X"F9",X"03",X"C0",X"03",X"8A",X"03",X"57",X"03",X"27",X"03",
		X"FA",X"02",X"CF",X"02",X"A7",X"02",X"81",X"02",X"5D",X"02",X"3B",X"02",X"1B",X"02",X"FD",X"01",
		X"E0",X"01",X"C5",X"01",X"AC",X"01",X"94",X"01",X"7D",X"01",X"68",X"01",X"53",X"01",X"40",X"01",
		X"2E",X"01",X"1D",X"01",X"0D",X"01",X"FE",X"00",X"F0",X"00",X"E3",X"00",X"D6",X"00",X"CA",X"00",
		X"BE",X"00",X"B4",X"00",X"AA",X"00",X"A0",X"00",X"97",X"00",X"8F",X"00",X"87",X"00",X"7F",X"00",
		X"78",X"00",X"71",X"00",X"6B",X"00",X"65",X"00",X"5F",X"00",X"5A",X"00",X"55",X"00",X"50",X"00",
		X"4C",X"00",X"47",X"00",X"6A",X"08",X"F1",X"07",X"7F",X"07",X"15",X"07",X"AD",X"06",X"4D",X"06",
		X"F2",X"05",X"9D",X"05",X"4D",X"05",X"00",X"05",X"B8",X"04",X"75",X"04",X"35",X"04",X"F8",X"03",
		X"BF",X"03",X"89",X"03",X"56",X"03",X"26",X"03",X"F9",X"02",X"CE",X"02",X"A6",X"02",X"80",X"02",
		X"5C",X"02",X"3A",X"02",X"1A",X"02",X"FC",X"01",X"DF",X"01",X"C4",X"01",X"AB",X"01",X"93",X"01",
		X"7C",X"01",X"67",X"01",X"52",X"01",X"3F",X"01",X"2D",X"01",X"1C",X"01",X"0C",X"01",X"FD",X"00",
		X"EF",X"00",X"E2",X"00",X"D5",X"00",X"C9",X"00",X"BD",X"00",X"B3",X"00",X"A9",X"00",X"9F",X"00",
		X"96",X"00",X"8E",X"00",X"86",X"00",X"7E",X"00",X"77",X"00",X"70",X"00",X"6A",X"00",X"64",X"00",
		X"5E",X"00",X"59",X"00",X"54",X"00",X"4F",X"00",X"4B",X"00",X"46",X"00",X"46",X"3F",X"38",X"31",
		X"2B",X"26",X"21",X"1C",X"18",X"15",X"12",X"0F",X"0D",X"0C",X"0B",X"0A",X"3A",X"04",X"30",X"FE",
		X"00",X"C2",X"F5",X"0D",X"3E",X"01",X"2E",X"00",X"CD",X"34",X"04",X"3E",X"02",X"2E",X"00",X"CD",
		X"34",X"04",X"3E",X"03",X"2E",X"00",X"CD",X"34",X"04",X"3E",X"01",X"CD",X"7B",X"03",X"3E",X"02",
		X"CD",X"7B",X"03",X"3E",X"03",X"CD",X"7B",X"03",X"21",X"EA",X"0A",X"11",X"14",X"30",X"01",X"30",
		X"00",X"ED",X"B0",X"3A",X"12",X"30",X"07",X"4F",X"07",X"81",X"4F",X"06",X"00",X"21",X"F3",X"0E",
		X"09",X"11",X"16",X"30",X"CD",X"E0",X"0A",X"11",X"26",X"30",X"CD",X"E0",X"0A",X"11",X"36",X"30",
		X"7E",X"12",X"CD",X"E7",X"0A",X"7E",X"12",X"23",X"13",X"C9",X"01",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3A",X"04",X"30",X"FE",X"00",X"C2",
		X"7B",X"0E",X"DD",X"21",X"14",X"30",X"CD",X"E0",X"05",X"DD",X"7E",X"08",X"FE",X"01",X"28",X"28",
		X"FE",X"02",X"28",X"3B",X"DD",X"21",X"24",X"30",X"CD",X"EF",X"05",X"DD",X"21",X"34",X"30",X"CD",
		X"09",X"06",X"3C",X"28",X"02",X"AF",X"C9",X"DD",X"21",X"14",X"30",X"3E",X"FF",X"DD",X"BE",X"00",
		X"20",X"04",X"DD",X"BE",X"10",X"C8",X"AF",X"C9",X"DD",X"21",X"14",X"30",X"CD",X"32",X"06",X"DD",
		X"21",X"34",X"30",X"CD",X"41",X"06",X"DD",X"21",X"24",X"30",X"CD",X"41",X"06",X"18",X"15",X"DD",
		X"21",X"14",X"30",X"CD",X"23",X"06",X"DD",X"21",X"24",X"30",X"CD",X"EF",X"05",X"DD",X"21",X"34",
		X"30",X"CD",X"41",X"06",X"DD",X"21",X"14",X"30",X"3E",X"FF",X"DD",X"BE",X"00",X"20",X"09",X"DD",
		X"BE",X"0A",X"20",X"04",X"DD",X"BE",X"10",X"C8",X"AF",X"C9",X"DD",X"7E",X"00",X"FE",X"FF",X"C8",
		X"DD",X"36",X"09",X"01",X"CD",X"06",X"0C",X"AF",X"C9",X"DD",X"7E",X"00",X"FE",X"FF",X"28",X"09",
		X"DD",X"36",X"09",X"02",X"CD",X"06",X"0C",X"AF",X"C9",X"0E",X"00",X"3E",X"02",X"CD",X"ED",X"03",
		X"3E",X"FF",X"C9",X"DD",X"7E",X"00",X"FE",X"FF",X"28",X"09",X"DD",X"36",X"09",X"03",X"CD",X"06",
		X"0C",X"AF",X"C9",X"0E",X"00",X"3E",X"03",X"CD",X"ED",X"03",X"3E",X"FF",X"C9",X"DD",X"7E",X"0A",
		X"FE",X"FF",X"C8",X"DD",X"36",X"09",X"04",X"CD",X"E4",X"0C",X"AF",X"C9",X"DD",X"7E",X"0A",X"FE",
		X"FF",X"C8",X"DD",X"36",X"09",X"05",X"CD",X"E4",X"0C",X"AF",X"C9",X"DD",X"7E",X"00",X"FE",X"FF",
		X"C8",X"CD",X"48",X"0D",X"AF",X"C9",X"DD",X"35",X"01",X"C0",X"3A",X"7E",X"30",X"DD",X"77",X"01",
		X"DD",X"CB",X"00",X"46",X"C2",X"29",X"0C",X"DD",X"7E",X"07",X"D6",X"01",X"FA",X"6F",X"06",X"DD",
		X"77",X"07",X"4F",X"DD",X"7E",X"09",X"CD",X"ED",X"03",X"DD",X"35",X"00",X"C0",X"DD",X"6E",X"02",
		X"DD",X"66",X"03",X"7E",X"47",X"E6",X"1F",X"CA",X"37",X"07",X"FE",X"1F",X"C2",X"45",X"07",X"23",
		X"DD",X"75",X"02",X"DD",X"74",X"03",X"78",X"E6",X"E0",X"0F",X"0F",X"0F",X"0F",X"4F",X"06",X"00",
		X"21",X"59",X"0C",X"09",X"5E",X"23",X"56",X"EB",X"E9",X"69",X"0C",X"9F",X"0C",X"C1",X"0C",X"B5",
		X"0C",X"2A",X"07",X"2A",X"07",X"2A",X"07",X"2A",X"07",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"4E",
		X"CB",X"21",X"06",X"00",X"21",X"34",X"09",X"09",X"5E",X"23",X"56",X"ED",X"53",X"7A",X"30",X"DD",
		X"73",X"04",X"DD",X"72",X"05",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"4E",X"CB",X"21",X"06",X"00",
		X"21",X"60",X"09",X"09",X"5E",X"23",X"56",X"DD",X"73",X"0B",X"DD",X"72",X"0C",X"18",X"35",X"DD",
		X"6E",X"02",X"DD",X"66",X"03",X"4E",X"06",X"00",X"21",X"7C",X"0A",X"09",X"7E",X"32",X"7E",X"30",
		X"DD",X"77",X"01",X"18",X"1F",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"7E",X"DD",X"77",X"08",X"18",
		X"13",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"7E",X"DD",X"77",X"06",X"DD",X"77",X"07",X"DD",X"77",
		X"0D",X"DD",X"77",X"0E",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"23",X"DD",X"75",X"02",X"DD",X"74",
		X"03",X"C3",X"2D",X"0C",X"DD",X"35",X"0F",X"C0",X"3A",X"7E",X"30",X"DD",X"77",X"0F",X"DD",X"CB",
		X"0A",X"46",X"C2",X"17",X"0D",X"DD",X"7E",X"0E",X"D6",X"01",X"FA",X"17",X"0D",X"DD",X"77",X"0E",
		X"DD",X"7E",X"09",X"FE",X"04",X"28",X"08",X"DD",X"4E",X"0E",X"3E",X"02",X"CD",X"ED",X"03",X"DD",
		X"4E",X"0E",X"3E",X"03",X"CD",X"ED",X"03",X"DD",X"35",X"0A",X"C0",X"DD",X"6E",X"02",X"DD",X"66",
		X"03",X"2B",X"7E",X"47",X"E6",X"1F",X"CA",X"D4",X"07",X"FE",X"1F",X"C2",X"ED",X"07",X"DD",X"7E",
		X"09",X"FE",X"04",X"28",X"07",X"3E",X"02",X"0E",X"00",X"CD",X"ED",X"03",X"3E",X"03",X"0E",X"00",
		X"CD",X"ED",X"03",X"DD",X"36",X"0A",X"FF",X"C9",X"DD",X"35",X"01",X"C0",X"3A",X"7E",X"30",X"DD",
		X"77",X"01",X"DD",X"CB",X"00",X"46",X"C2",X"64",X"0D",X"DD",X"7E",X"07",X"D6",X"01",X"FA",X"64",
		X"0D",X"DD",X"77",X"07",X"DD",X"35",X"00",X"C0",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"7E",X"47",
		X"E6",X"1F",X"CA",X"F0",X"08",X"FE",X"1F",X"C2",X"F6",X"08",X"23",X"DD",X"75",X"02",X"DD",X"74",
		X"03",X"78",X"E6",X"E0",X"0F",X"0F",X"0F",X"0F",X"4F",X"06",X"00",X"21",X"94",X"0D",X"09",X"5E",
		X"23",X"56",X"EB",X"E9",X"A4",X"0D",X"C2",X"0D",X"D8",X"0D",X"EB",X"08",X"EB",X"08",X"EB",X"08",
		X"EB",X"08",X"EB",X"08",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"4E",X"CB",X"21",X"06",X"00",X"21",
		X"34",X"09",X"09",X"5E",X"23",X"56",X"ED",X"53",X"7A",X"30",X"DD",X"73",X"04",X"DD",X"72",X"05",
		X"18",X"23",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"4E",X"06",X"00",X"21",X"7C",X"0A",X"09",X"7E",
		X"32",X"7E",X"30",X"DD",X"77",X"01",X"18",X"0D",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"7E",X"DD",
		X"77",X"06",X"DD",X"77",X"07",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"23",X"DD",X"75",X"02",X"DD",
		X"74",X"03",X"C3",X"68",X"0D",X"3E",X"01",X"2E",X"00",X"CD",X"34",X"04",X"3E",X"02",X"2E",X"00",
		X"CD",X"34",X"04",X"3E",X"03",X"2E",X"00",X"CD",X"34",X"04",X"3E",X"01",X"CD",X"7B",X"03",X"3E",
		X"02",X"CD",X"7B",X"03",X"3E",X"03",X"CD",X"7B",X"03",X"21",X"4B",X"0E",X"11",X"4A",X"30",X"01",
		X"30",X"00",X"ED",X"B0",X"3A",X"80",X"30",X"07",X"4F",X"07",X"81",X"4F",X"06",X"00",X"21",X"F3",
		X"0E",X"09",X"11",X"4C",X"30",X"CD",X"41",X"0E",X"11",X"5C",X"30",X"CD",X"41",X"0E",X"11",X"6C",
		X"30",X"7E",X"12",X"CD",X"48",X"0E",X"7E",X"12",X"23",X"13",X"C9",X"01",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DD",X"21",X"4A",X"30",X"CD",
		X"9A",X"0B",X"DD",X"7E",X"08",X"FE",X"01",X"28",X"28",X"FE",X"02",X"28",X"3B",X"DD",X"21",X"5A",
		X"30",X"CD",X"A9",X"0B",X"DD",X"21",X"6A",X"30",X"CD",X"C3",X"0B",X"3C",X"28",X"02",X"AF",X"C9",
		X"DD",X"21",X"4A",X"30",X"3E",X"FF",X"DD",X"BE",X"00",X"20",X"04",X"DD",X"BE",X"10",X"C8",X"AF",
		X"C9",X"DD",X"21",X"4A",X"30",X"CD",X"EC",X"0B",X"DD",X"21",X"6A",X"30",X"CD",X"FB",X"0B",X"DD",
		X"21",X"5A",X"30",X"CD",X"FB",X"0B",X"18",X"15",X"DD",X"21",X"4A",X"30",X"CD",X"DD",X"0B",X"DD",
		X"21",X"5A",X"30",X"CD",X"A9",X"0B",X"DD",X"21",X"6A",X"30",X"CD",X"FB",X"0B",X"DD",X"21",X"4A",
		X"30",X"3E",X"FF",X"DD",X"BE",X"00",X"20",X"09",X"DD",X"BE",X"0A",X"20",X"04",X"DD",X"BE",X"10",
		X"C8",X"AF",X"C9",X"6B",X"10",X"81",X"10",X"95",X"10",X"9D",X"10",X"CD",X"10",X"FB",X"10",X"BD",
		X"13",X"0F",X"14",X"5F",X"14",X"23",X"11",X"34",X"11",X"43",X"11",X"6B",X"10",X"81",X"10",X"95",
		X"10",X"52",X"11",X"EC",X"11",X"24",X"12",X"5C",X"12",X"AE",X"12",X"FE",X"12",X"6B",X"10",X"81",
		X"10",X"95",X"10",X"BF",X"14",X"D1",X"14",X"0A",X"15",X"6B",X"10",X"81",X"10",X"95",X"10",X"FC",
		X"10",X"11",X"11",X"22",X"11",X"6B",X"10",X"81",X"10",X"95",X"10",X"60",X"14",X"90",X"14",X"BE",
		X"14",X"FF",X"12",X"15",X"13",X"29",X"13",X"31",X"13",X"40",X"13",X"49",X"13",X"4A",X"13",X"59",
		X"13",X"62",X"13",X"6B",X"10",X"81",X"10",X"95",X"10",X"6B",X"10",X"81",X"10",X"95",X"10",X"63",
		X"13",X"7F",X"13",X"80",X"13",X"81",X"13",X"9D",X"13",X"9E",X"13",X"9F",X"13",X"BB",X"13",X"BC",
		X"13",X"6B",X"10",X"81",X"10",X"95",X"10",X"6B",X"10",X"81",X"10",X"95",X"10",X"3E",X"00",X"32",
		X"12",X"30",X"32",X"80",X"30",X"CD",X"8C",X"0A",X"AF",X"C9",X"CD",X"1A",X"0B",X"C9",X"3E",X"01",
		X"32",X"12",X"30",X"32",X"80",X"30",X"CD",X"8C",X"0A",X"AF",X"C9",X"CD",X"1A",X"0B",X"C9",X"3E",
		X"08",X"32",X"12",X"30",X"32",X"80",X"30",X"CD",X"8C",X"0A",X"AF",X"C9",X"CD",X"1A",X"0B",X"C9",
		X"3E",X"03",X"32",X"12",X"30",X"32",X"80",X"30",X"CD",X"8C",X"0A",X"AF",X"C9",X"CD",X"1A",X"0B",
		X"C9",X"3E",X"0C",X"32",X"12",X"30",X"32",X"80",X"30",X"CD",X"8C",X"0A",X"AF",X"C9",X"CD",X"1A",
		X"0B",X"C9",X"3E",X"05",X"32",X"12",X"30",X"32",X"80",X"30",X"CD",X"8C",X"0A",X"AF",X"C9",X"CD",
		X"1A",X"0B",X"C9",X"3E",X"06",X"32",X"12",X"30",X"32",X"80",X"30",X"CD",X"8C",X"0A",X"AF",X"C9",
		X"CD",X"1A",X"0B",X"C9",X"3E",X"0A",X"32",X"12",X"30",X"32",X"80",X"30",X"CD",X"8C",X"0A",X"AF",
		X"C9",X"CD",X"1A",X"0B",X"C9",X"3E",X"0E",X"32",X"12",X"30",X"32",X"80",X"30",X"CD",X"8C",X"0A",
		X"AF",X"C9",X"CD",X"1A",X"0B",X"C9",X"3E",X"0F",X"32",X"12",X"30",X"32",X"80",X"30",X"CD",X"8C",
		X"0A",X"AF",X"C9",X"CD",X"1A",X"0B",X"C9",X"3E",X"12",X"32",X"12",X"30",X"32",X"80",X"30",X"CD",
		X"8C",X"0A",X"AF",X"C9",X"CD",X"1A",X"0B",X"C9",X"3E",X"13",X"32",X"12",X"30",X"32",X"80",X"30",
		X"CD",X"8C",X"0A",X"AF",X"C9",X"CD",X"1A",X"0B",X"C9",X"3E",X"14",X"32",X"12",X"30",X"32",X"80",
		X"30",X"CD",X"8C",X"0A",X"AF",X"C9",X"CD",X"1A",X"0B",X"C9",X"3E",X"02",X"32",X"12",X"30",X"32",
		X"80",X"30",X"CD",X"8C",X"0A",X"AF",X"C9",X"CD",X"1A",X"0B",X"C9",X"1F",X"0F",X"3F",X"0F",X"5F",
		X"09",X"7F",X"00",X"22",X"23",X"24",X"25",X"23",X"24",X"25",X"26",X"24",X"25",X"26",X"27",X"A8",
		X"FF",X"1F",X"0F",X"3F",X"0F",X"5F",X"09",X"26",X"27",X"28",X"29",X"27",X"28",X"29",X"2A",X"28",
		X"29",X"2A",X"2B",X"AC",X"FF",X"1F",X"08",X"3F",X"0F",X"5F",X"08",X"A2",X"FF",X"1F",X"0D",X"3F",
		X"0A",X"5F",X"09",X"7F",X"00",X"2E",X"2E",X"20",X"30",X"30",X"20",X"32",X"32",X"20",X"30",X"30",
		X"20",X"32",X"32",X"20",X"33",X"33",X"20",X"32",X"32",X"20",X"33",X"33",X"20",X"35",X"35",X"20",
		X"33",X"33",X"20",X"35",X"35",X"20",X"37",X"37",X"20",X"3F",X"05",X"B5",X"FF",X"1F",X"0D",X"3F",
		X"0A",X"5F",X"09",X"32",X"32",X"20",X"33",X"33",X"20",X"35",X"35",X"20",X"33",X"33",X"20",X"35",
		X"35",X"20",X"37",X"37",X"20",X"35",X"35",X"20",X"37",X"37",X"20",X"39",X"39",X"20",X"37",X"37",
		X"20",X"39",X"39",X"20",X"3A",X"3A",X"20",X"3F",X"05",X"B2",X"FF",X"FF",X"1F",X"0E",X"3F",X"0F",
		X"5F",X"09",X"7F",X"02",X"6B",X"60",X"80",X"70",X"60",X"80",X"74",X"60",X"80",X"3F",X"05",X"B7",
		X"FF",X"1F",X"0E",X"3F",X"0F",X"5F",X"09",X"64",X"60",X"80",X"6B",X"60",X"80",X"70",X"60",X"80",
		X"B4",X"FF",X"FF",X"1F",X"0E",X"3F",X"0C",X"5F",X"09",X"7F",X"00",X"4E",X"52",X"55",X"5A",X"52",
		X"55",X"5A",X"5E",X"FF",X"1F",X"0E",X"3F",X"0C",X"5F",X"09",X"49",X"4E",X"52",X"55",X"4E",X"52",
		X"55",X"5A",X"FF",X"1F",X"08",X"3F",X"0C",X"5F",X"08",X"46",X"49",X"4E",X"52",X"49",X"4E",X"52",
		X"55",X"FF",X"1F",X"0E",X"3F",X"0B",X"5F",X"09",X"7F",X"02",X"70",X"7F",X"00",X"70",X"7F",X"02",
		X"72",X"7F",X"00",X"70",X"7F",X"02",X"73",X"7F",X"00",X"70",X"7F",X"02",X"75",X"7F",X"00",X"70",
		X"7F",X"02",X"73",X"7F",X"00",X"70",X"7F",X"02",X"72",X"7F",X"00",X"70",X"7F",X"02",X"70",X"7F",
		X"00",X"70",X"7F",X"02",X"6E",X"7F",X"00",X"70",X"7F",X"02",X"70",X"7F",X"00",X"70",X"7F",X"02",
		X"72",X"7F",X"00",X"70",X"7F",X"02",X"73",X"7F",X"00",X"70",X"7F",X"02",X"75",X"7F",X"00",X"70",
		X"7F",X"02",X"73",X"7F",X"00",X"70",X"7F",X"02",X"72",X"7F",X"00",X"70",X"7F",X"02",X"70",X"7F",
		X"00",X"70",X"7F",X"02",X"6E",X"7F",X"00",X"70",X"7F",X"02",X"70",X"7F",X"00",X"70",X"7F",X"02",
		X"72",X"7F",X"00",X"70",X"7F",X"02",X"6E",X"7F",X"00",X"70",X"7F",X"02",X"70",X"7F",X"00",X"70",
		X"7F",X"02",X"72",X"7F",X"00",X"70",X"7F",X"02",X"6E",X"7F",X"00",X"70",X"7F",X"02",X"70",X"7F",
		X"00",X"70",X"7F",X"02",X"72",X"7F",X"00",X"70",X"7F",X"02",X"B0",X"FF",X"1F",X"08",X"3F",X"0B",
		X"5F",X"08",X"70",X"70",X"72",X"70",X"73",X"70",X"75",X"70",X"73",X"70",X"72",X"70",X"70",X"70",
		X"6E",X"70",X"70",X"70",X"72",X"70",X"73",X"70",X"75",X"70",X"73",X"70",X"72",X"70",X"70",X"70",
		X"6E",X"70",X"70",X"70",X"72",X"70",X"6E",X"70",X"70",X"70",X"72",X"70",X"6E",X"70",X"70",X"70",
		X"72",X"70",X"B0",X"FF",X"1F",X"02",X"3F",X"0B",X"5F",X"08",X"70",X"70",X"72",X"70",X"73",X"70",
		X"75",X"70",X"73",X"70",X"72",X"70",X"70",X"70",X"6E",X"70",X"70",X"70",X"72",X"70",X"73",X"70",
		X"75",X"70",X"73",X"70",X"72",X"70",X"70",X"70",X"6E",X"70",X"70",X"70",X"72",X"70",X"6E",X"70",
		X"70",X"70",X"72",X"70",X"6E",X"70",X"70",X"70",X"72",X"70",X"B0",X"FF",X"1F",X"0E",X"3F",X"0A",
		X"5F",X"09",X"7F",X"02",X"77",X"75",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"37",
		X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"37",
		X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"B7",X"60",
		X"75",X"73",X"72",X"70",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"30",X"30",X"30",X"30",
		X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"B0",X"FF",X"1F",X"02",
		X"3F",X"0A",X"5F",X"08",X"77",X"75",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"37",
		X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"37",
		X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"B7",X"60",
		X"75",X"73",X"72",X"70",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"30",X"30",X"30",X"30",
		X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"B0",X"FF",X"FF",X"1F",
		X"0E",X"3F",X"07",X"5F",X"09",X"7F",X"00",X"22",X"23",X"24",X"25",X"26",X"27",X"28",X"29",X"2A");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
