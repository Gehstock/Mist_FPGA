library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity sol_sound_cpu is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of sol_sound_cpu is
	type rom is array(0 to  12287) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"F3",X"00",X"00",X"00",X"31",X"F6",X"83",X"ED",X"56",X"18",X"55",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F5",X"E5",X"C5",X"3A",X"00",X"E0",X"CD",X"D9",
		X"01",X"3A",X"76",X"83",X"3D",X"28",X"08",X"32",X"76",X"83",X"C1",X"E1",X"F1",X"FB",X"C9",X"3C",
		X"32",X"75",X"83",X"3E",X"04",X"32",X"76",X"83",X"C1",X"E1",X"F1",X"FB",X"C9",X"FF",X"FF",X"FF",
		X"21",X"00",X"B0",X"36",X"0F",X"21",X"02",X"B0",X"36",X"F0",X"3A",X"00",X"F0",X"CB",X"47",X"20",
		X"4F",X"CB",X"4F",X"20",X"2E",X"AF",X"32",X"78",X"83",X"CD",X"31",X"04",X"CD",X"EA",X"04",X"3A",
		X"78",X"83",X"FE",X"00",X"28",X"1D",X"CB",X"67",X"20",X"05",X"01",X"00",X"10",X"18",X"03",X"01",
		X"00",X"80",X"11",X"01",X"00",X"60",X"69",X"32",X"00",X"D0",X"37",X"3F",X"ED",X"52",X"20",X"FC",
		X"2F",X"18",X"F2",X"3E",X"FF",X"32",X"00",X"D0",X"3A",X"00",X"F0",X"CB",X"57",X"20",X"08",X"CD",
		X"5F",X"03",X"18",X"EF",X"3A",X"00",X"F0",X"CB",X"5F",X"20",X"F9",X"CD",X"86",X"03",X"18",X"F4",
		X"06",X"00",X"CD",X"41",X"05",X"06",X"FF",X"CD",X"41",X"05",X"06",X"55",X"CD",X"41",X"05",X"06",
		X"AA",X"CD",X"41",X"05",X"AF",X"32",X"78",X"83",X"CD",X"31",X"04",X"CD",X"EA",X"04",X"3A",X"78",
		X"83",X"32",X"00",X"C0",X"CD",X"E7",X"00",X"31",X"F6",X"83",X"F3",X"ED",X"56",X"CD",X"0C",X"01",
		X"CD",X"81",X"0F",X"FB",X"AF",X"32",X"75",X"83",X"CD",X"F6",X"01",X"CD",X"7B",X"01",X"CD",X"F0",
		X"0A",X"CD",X"81",X"0F",X"3A",X"75",X"83",X"B7",X"28",X"FA",X"18",X"E8",X"21",X"32",X"11",X"06",
		X"20",X"11",X"20",X"80",X"DD",X"21",X"00",X"80",X"7E",X"DD",X"77",X"00",X"2F",X"12",X"13",X"23",
		X"DD",X"23",X"10",X"F4",X"06",X"06",X"11",X"09",X"00",X"DD",X"21",X"BC",X"82",X"DD",X"36",X"00",
		X"FF",X"DD",X"36",X"01",X"FF",X"DD",X"36",X"02",X"00",X"DD",X"36",X"03",X"00",X"DD",X"36",X"04",
		X"00",X"DD",X"36",X"05",X"00",X"DD",X"36",X"06",X"00",X"DD",X"19",X"10",X"E0",X"06",X"03",X"21",
		X"6B",X"83",X"36",X"00",X"23",X"10",X"FB",X"3E",X"01",X"32",X"0C",X"83",X"32",X"20",X"83",X"3D",
		X"32",X"1F",X"83",X"3A",X"00",X"90",X"E6",X"80",X"32",X"6E",X"83",X"3E",X"55",X"32",X"71",X"83",
		X"3E",X"04",X"32",X"76",X"83",X"3E",X"40",X"32",X"77",X"83",X"C9",X"3A",X"6E",X"83",X"47",X"3A",
		X"00",X"90",X"A8",X"CB",X"7F",X"20",X"31",X"CB",X"40",X"28",X"1E",X"CB",X"80",X"78",X"32",X"6E",
		X"83",X"CD",X"5E",X"05",X"3A",X"70",X"83",X"CB",X"47",X"28",X"0E",X"CD",X"0F",X"06",X"CD",X"1C",
		X"07",X"CD",X"7F",X"07",X"CD",X"9C",X"08",X"18",X"23",X"CD",X"1C",X"07",X"3A",X"6F",X"83",X"CB",
		X"47",X"28",X"19",X"CD",X"9C",X"08",X"18",X"14",X"78",X"2F",X"CB",X"C7",X"32",X"6E",X"83",X"CD",
		X"1C",X"07",X"3A",X"6F",X"83",X"CB",X"47",X"28",X"03",X"CD",X"9C",X"08",X"3E",X"01",X"32",X"20",
		X"83",X"32",X"0C",X"83",X"3D",X"32",X"1F",X"83",X"C9",X"3A",X"00",X"F0",X"47",X"E6",X"10",X"20",
		X"08",X"21",X"F8",X"83",X"BE",X"77",X"20",X"05",X"C9",X"32",X"F8",X"83",X"C9",X"78",X"E6",X"0F",
		X"F6",X"80",X"32",X"F9",X"83",X"C9",X"3A",X"F9",X"83",X"B7",X"FA",X"FE",X"01",X"C9",X"E6",X"0F",
		X"32",X"F9",X"83",X"47",X"3A",X"FE",X"83",X"B7",X"F2",X"5C",X"02",X"CB",X"77",X"CA",X"38",X"02",
		X"21",X"FA",X"83",X"16",X"00",X"E6",X"03",X"5F",X"19",X"7E",X"E6",X"F0",X"B0",X"77",X"3A",X"FE",
		X"83",X"E6",X"7F",X"32",X"FE",X"83",X"E6",X"03",X"FE",X"03",X"28",X"07",X"3A",X"FE",X"83",X"3C",
		X"32",X"FE",X"83",X"3E",X"50",X"C3",X"49",X"03",X"21",X"FA",X"83",X"16",X"00",X"3A",X"FE",X"83",
		X"E6",X"03",X"5F",X"19",X"78",X"07",X"07",X"07",X"07",X"47",X"7E",X"E6",X"0F",X"B0",X"77",X"3A",
		X"FE",X"83",X"CB",X"F7",X"32",X"FE",X"83",X"3E",X"50",X"C3",X"49",X"03",X"78",X"FE",X"0F",X"C2",
		X"71",X"02",X"3A",X"FE",X"83",X"E6",X"03",X"F6",X"80",X"32",X"FE",X"83",X"3E",X"F0",X"C3",X"49",
		X"03",X"FE",X"0E",X"C2",X"B2",X"02",X"3A",X"FB",X"83",X"32",X"01",X"90",X"3A",X"FC",X"83",X"32",
		X"02",X"90",X"3A",X"FD",X"83",X"32",X"03",X"90",X"3A",X"00",X"90",X"EE",X"80",X"E6",X"80",X"47",
		X"3A",X"FA",X"83",X"E6",X"7F",X"5F",X"3A",X"F7",X"83",X"BB",X"3E",X"00",X"28",X"0F",X"7B",X"32",
		X"F7",X"83",X"4F",X"0F",X"E6",X"38",X"57",X"79",X"E6",X"07",X"B2",X"F6",X"40",X"B0",X"32",X"00",
		X"90",X"C9",X"FE",X"0D",X"C2",X"D1",X"02",X"3E",X"83",X"32",X"FE",X"83",X"3A",X"FB",X"83",X"F6",
		X"80",X"32",X"FB",X"83",X"3A",X"FC",X"83",X"F6",X"80",X"32",X"FC",X"83",X"3E",X"F0",X"C3",X"49",
		X"03",X"FE",X"0C",X"C2",X"F0",X"02",X"3E",X"83",X"32",X"FE",X"83",X"3A",X"FB",X"83",X"F6",X"80",
		X"32",X"FB",X"83",X"3A",X"FC",X"83",X"E6",X"7F",X"32",X"FC",X"83",X"3E",X"F0",X"C3",X"49",X"03",
		X"FE",X"0A",X"C2",X"1D",X"03",X"AF",X"32",X"02",X"90",X"32",X"FA",X"83",X"32",X"FB",X"83",X"32",
		X"FC",X"83",X"32",X"FD",X"83",X"32",X"03",X"90",X"3E",X"02",X"32",X"01",X"90",X"3A",X"00",X"90",
		X"E6",X"80",X"EE",X"80",X"32",X"00",X"90",X"3E",X"01",X"32",X"FE",X"83",X"C9",X"FE",X"0B",X"C2",
		X"39",X"03",X"3E",X"01",X"32",X"FE",X"83",X"AF",X"32",X"FA",X"83",X"32",X"FB",X"83",X"32",X"FC",
		X"83",X"32",X"FD",X"83",X"3E",X"F0",X"C3",X"49",X"03",X"FE",X"00",X"C2",X"48",X"03",X"3E",X"80",
		X"32",X"FE",X"83",X"3E",X"F0",X"C3",X"49",X"03",X"C9",X"32",X"03",X"90",X"3E",X"AC",X"32",X"01",
		X"90",X"3E",X"80",X"32",X"02",X"90",X"3A",X"00",X"90",X"EE",X"80",X"32",X"00",X"90",X"C9",X"06",
		X"00",X"CD",X"C0",X"03",X"0E",X"00",X"3E",X"AD",X"CD",X"00",X"04",X"0E",X"01",X"3E",X"07",X"CD",
		X"00",X"04",X"06",X"01",X"CD",X"C0",X"03",X"0E",X"00",X"3E",X"AD",X"CD",X"00",X"04",X"0E",X"01",
		X"3E",X"77",X"CD",X"00",X"04",X"C9",X"F3",X"CD",X"5F",X"03",X"16",X"10",X"AF",X"1E",X"FF",X"06",
		X"00",X"0E",X"00",X"CD",X"00",X"04",X"2F",X"0E",X"01",X"CD",X"00",X"04",X"06",X"01",X"32",X"72",
		X"83",X"E6",X"7F",X"CD",X"00",X"04",X"3A",X"72",X"83",X"2F",X"0E",X"00",X"CD",X"00",X"04",X"3C",
		X"E6",X"0F",X"47",X"07",X"07",X"07",X"07",X"B0",X"1D",X"20",X"FD",X"15",X"20",X"CF",X"FB",X"C9",
		X"CD",X"17",X"04",X"36",X"00",X"DD",X"36",X"00",X"F4",X"36",X"01",X"DD",X"36",X"00",X"01",X"36",
		X"02",X"DD",X"36",X"00",X"FA",X"36",X"03",X"DD",X"36",X"00",X"00",X"36",X"04",X"DD",X"36",X"00",
		X"7D",X"36",X"05",X"DD",X"36",X"00",X"00",X"36",X"08",X"DD",X"36",X"00",X"0B",X"36",X"09",X"DD",
		X"36",X"00",X"0B",X"36",X"0A",X"DD",X"36",X"00",X"0B",X"36",X"07",X"DD",X"36",X"00",X"F8",X"C9",
		X"CD",X"17",X"04",X"32",X"73",X"83",X"AF",X"A9",X"28",X"09",X"36",X"0F",X"3A",X"73",X"83",X"DD",
		X"77",X"00",X"C9",X"36",X"0E",X"18",X"F5",X"32",X"73",X"83",X"AF",X"A8",X"3A",X"73",X"83",X"20",
		X"08",X"21",X"00",X"A0",X"DD",X"21",X"02",X"A0",X"C9",X"21",X"00",X"B0",X"DD",X"21",X"02",X"B0",
		X"C9",X"DD",X"21",X"DA",X"04",X"AF",X"F5",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"7C",X"B5",X"20",
		X"0A",X"F1",X"47",X"3A",X"78",X"83",X"B0",X"32",X"78",X"83",X"C9",X"DD",X"5E",X"04",X"DD",X"56",
		X"05",X"DD",X"4E",X"02",X"DD",X"46",X"03",X"ED",X"B0",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"DD",
		X"5E",X"02",X"DD",X"56",X"03",X"7A",X"B3",X"28",X"11",X"06",X"02",X"3E",X"00",X"77",X"BE",X"C2",
		X"D5",X"04",X"F6",X"FF",X"10",X"F7",X"23",X"1B",X"18",X"EB",X"DD",X"66",X"01",X"DD",X"6E",X"00",
		X"DD",X"5E",X"02",X"DD",X"56",X"03",X"7A",X"B3",X"28",X"06",X"36",X"00",X"23",X"1B",X"18",X"F6",
		X"DD",X"6E",X"00",X"DD",X"66",X"01",X"DD",X"5E",X"02",X"DD",X"56",X"03",X"7A",X"B3",X"28",X"15",
		X"7E",X"FE",X"00",X"C2",X"D5",X"04",X"3E",X"01",X"77",X"BE",X"C2",X"D5",X"04",X"CB",X"27",X"30",
		X"F7",X"23",X"1B",X"18",X"E7",X"AF",X"DD",X"66",X"05",X"DD",X"6E",X"04",X"DD",X"56",X"01",X"DD",
		X"5E",X"00",X"DD",X"4E",X"02",X"DD",X"46",X"03",X"ED",X"B0",X"47",X"F1",X"B0",X"11",X"07",X"00",
		X"DD",X"19",X"C3",X"36",X"04",X"DD",X"7E",X"06",X"18",X"DC",X"00",X"80",X"00",X"02",X"00",X"80",
		X"10",X"00",X"82",X"00",X"02",X"00",X"80",X"0A",X"00",X"00",X"DD",X"21",X"26",X"05",X"16",X"00",
		X"DD",X"6E",X"02",X"DD",X"66",X"03",X"DD",X"4E",X"00",X"DD",X"46",X"01",X"78",X"B1",X"28",X"1A",
		X"AF",X"86",X"23",X"0D",X"20",X"FB",X"05",X"20",X"F8",X"DD",X"BE",X"04",X"28",X"05",X"7A",X"DD",
		X"B6",X"05",X"57",X"01",X"06",X"00",X"DD",X"09",X"18",X"D6",X"7A",X"B7",X"C8",X"47",X"3A",X"78",
		X"83",X"B0",X"32",X"78",X"83",X"C9",X"00",X"10",X"00",X"00",X"00",X"01",X"00",X"10",X"00",X"10",
		X"F0",X"02",X"00",X"10",X"00",X"20",X"60",X"04",X"00",X"10",X"00",X"30",X"00",X"08",X"00",X"00",
		X"5A",X"3A",X"00",X"90",X"B8",X"20",X"FA",X"3A",X"01",X"90",X"B8",X"20",X"F4",X"3A",X"02",X"90",
		X"B8",X"20",X"EE",X"3A",X"03",X"90",X"B8",X"20",X"E8",X"78",X"32",X"00",X"C0",X"C9",X"3E",X"01",
		X"32",X"70",X"83",X"DD",X"21",X"00",X"90",X"DD",X"46",X"00",X"CB",X"70",X"28",X"23",X"FD",X"21",
		X"00",X"80",X"FD",X"7E",X"0F",X"E6",X"8F",X"4F",X"78",X"17",X"E6",X"70",X"B1",X"FD",X"77",X"0F",
		X"FD",X"7E",X"1F",X"E6",X"8F",X"4F",X"78",X"17",X"17",X"17",X"17",X"E6",X"70",X"B1",X"FD",X"77",
		X"1F",X"DD",X"7E",X"01",X"4F",X"FE",X"00",X"28",X"22",X"CB",X"7F",X"28",X"6A",X"DD",X"7E",X"02",
		X"CB",X"7F",X"20",X"63",X"79",X"E6",X"7F",X"4F",X"06",X"06",X"FD",X"21",X"BC",X"82",X"11",X"09",
		X"00",X"FD",X"7E",X"06",X"B9",X"28",X"23",X"FD",X"19",X"10",X"F6",X"FD",X"21",X"6B",X"83",X"DD",
		X"46",X"02",X"78",X"E6",X"7F",X"28",X"21",X"FD",X"77",X"01",X"DD",X"7E",X"01",X"CB",X"7F",X"C0",
		X"DD",X"7E",X"03",X"FE",X"00",X"C8",X"FD",X"77",X"02",X"C9",X"DD",X"7E",X"03",X"E5",X"FD",X"6E",
		X"07",X"FD",X"66",X"08",X"77",X"E1",X"18",X"D3",X"DD",X"4E",X"01",X"79",X"FE",X"00",X"20",X"09",
		X"DD",X"7E",X"03",X"FE",X"00",X"20",X"D3",X"18",X"09",X"CB",X"79",X"28",X"CD",X"CB",X"78",X"20",
		X"C9",X"AF",X"32",X"70",X"83",X"18",X"C3",X"79",X"E6",X"7F",X"32",X"6B",X"83",X"18",X"AC",X"06",
		X"03",X"21",X"6B",X"83",X"C5",X"7E",X"4F",X"FE",X"00",X"CA",X"DF",X"06",X"3A",X"77",X"83",X"91",
		X"DA",X"DF",X"06",X"79",X"FE",X"33",X"20",X"04",X"F3",X"C3",X"00",X"00",X"79",X"FE",X"01",X"20",
		X"0C",X"DD",X"21",X"00",X"80",X"DD",X"7E",X"1F",X"F6",X"80",X"DD",X"77",X"1F",X"79",X"FE",X"02",
		X"20",X"0F",X"DD",X"21",X"00",X"80",X"DD",X"7E",X"1F",X"E6",X"7F",X"DD",X"77",X"1F",X"CD",X"E6",
		X"06",X"79",X"FE",X"03",X"20",X"02",X"0E",X"04",X"79",X"FE",X"50",X"20",X"07",X"3E",X"40",X"32",
		X"77",X"83",X"18",X"0A",X"79",X"FE",X"50",X"20",X"05",X"3E",X"40",X"32",X"77",X"83",X"79",X"D9",
		X"6F",X"26",X"00",X"54",X"5D",X"29",X"29",X"19",X"19",X"19",X"11",X"11",X"12",X"19",X"EB",X"1A",
		X"FE",X"00",X"20",X"1F",X"01",X"0C",X"83",X"60",X"69",X"3E",X"06",X"08",X"13",X"1A",X"FE",X"00",
		X"28",X"4A",X"7E",X"CD",X"BC",X"0F",X"1A",X"77",X"60",X"69",X"34",X"08",X"3D",X"FE",X"00",X"20",
		X"EA",X"18",X"39",X"3E",X"06",X"21",X"20",X"83",X"08",X"13",X"1A",X"FE",X"00",X"28",X"2D",X"7E",
		X"CD",X"BC",X"0F",X"1A",X"77",X"26",X"00",X"6F",X"29",X"01",X"DE",X"15",X"09",X"01",X"20",X"83",
		X"0A",X"CB",X"27",X"E5",X"21",X"33",X"83",X"CD",X"BC",X"0F",X"EB",X"E3",X"7E",X"12",X"23",X"13",
		X"7E",X"12",X"0A",X"3C",X"02",X"D1",X"60",X"69",X"08",X"3D",X"20",X"CC",X"D9",X"AF",X"77",X"23",
		X"C1",X"05",X"C2",X"14",X"06",X"C9",X"D9",X"DD",X"21",X"BC",X"82",X"01",X"09",X"00",X"11",X"0C",
		X"83",X"3E",X"01",X"12",X"62",X"6B",X"3E",X"06",X"08",X"DD",X"7E",X"03",X"FE",X"00",X"28",X"0B",
		X"1A",X"CD",X"BC",X"0F",X"DD",X"7E",X"03",X"77",X"62",X"6B",X"34",X"DD",X"09",X"08",X"3D",X"20",
		X"E7",X"3E",X"00",X"32",X"1F",X"83",X"3C",X"32",X"20",X"83",X"D9",X"C9",X"AF",X"32",X"6F",X"83",
		X"21",X"0C",X"83",X"7E",X"D6",X"01",X"28",X"2A",X"11",X"09",X"00",X"4F",X"DD",X"21",X"BC",X"82",
		X"06",X"06",X"23",X"7E",X"DD",X"BE",X"04",X"20",X"13",X"AF",X"DD",X"77",X"06",X"DD",X"77",X"04",
		X"DD",X"77",X"05",X"3C",X"32",X"6F",X"83",X"0D",X"20",X"E2",X"18",X"06",X"DD",X"19",X"10",X"E4",
		X"18",X"F5",X"21",X"1F",X"83",X"7E",X"4F",X"FE",X"00",X"C8",X"3E",X"01",X"32",X"6F",X"83",X"06",
		X"06",X"21",X"5B",X"11",X"DD",X"21",X"BC",X"82",X"11",X"09",X"00",X"79",X"A6",X"28",X"0A",X"AF",
		X"DD",X"77",X"06",X"DD",X"77",X"04",X"DD",X"77",X"05",X"DD",X"19",X"23",X"10",X"ED",X"C9",X"3A",
		X"20",X"83",X"D6",X"01",X"C8",X"08",X"CD",X"B1",X"07",X"CD",X"CD",X"07",X"79",X"CB",X"27",X"21",
		X"33",X"83",X"CD",X"BC",X"0F",X"7A",X"FE",X"00",X"20",X"11",X"CB",X"7E",X"20",X"0A",X"E5",X"CD",
		X"0E",X"08",X"E1",X"7A",X"FE",X"00",X"20",X"03",X"CD",X"47",X"08",X"23",X"36",X"00",X"08",X"18",
		X"D1",X"06",X"00",X"0E",X"01",X"16",X"01",X"3A",X"20",X"83",X"5F",X"21",X"33",X"83",X"23",X"7A",
		X"BB",X"C8",X"23",X"23",X"78",X"BE",X"30",X"02",X"46",X"4A",X"14",X"18",X"F2",X"79",X"CB",X"27",
		X"21",X"33",X"83",X"CD",X"BC",X"0F",X"C5",X"06",X"06",X"4E",X"11",X"09",X"00",X"21",X"5B",X"11",
		X"DD",X"21",X"BC",X"82",X"7E",X"A1",X"28",X"1D",X"DD",X"7E",X"04",X"FE",X"00",X"20",X"16",X"21",
		X"20",X"83",X"C1",X"79",X"CD",X"BC",X"0F",X"7E",X"DD",X"77",X"04",X"DD",X"70",X"05",X"AF",X"DD",
		X"77",X"03",X"16",X"01",X"C9",X"DD",X"19",X"23",X"10",X"DA",X"16",X"00",X"C1",X"C9",X"26",X"06",
		X"11",X"09",X"00",X"DD",X"21",X"BC",X"82",X"DD",X"7E",X"04",X"FE",X"00",X"20",X"15",X"79",X"21",
		X"20",X"83",X"CD",X"BC",X"0F",X"7E",X"DD",X"77",X"04",X"DD",X"70",X"05",X"AF",X"DD",X"77",X"03",
		X"16",X"01",X"C9",X"DD",X"19",X"25",X"20",X"DF",X"16",X"00",X"21",X"33",X"83",X"79",X"CB",X"27",
		X"CD",X"BC",X"0F",X"F6",X"3F",X"77",X"C9",X"16",X"FF",X"1E",X"00",X"E5",X"C5",X"4E",X"06",X"00",
		X"DD",X"21",X"BC",X"82",X"21",X"5B",X"11",X"7E",X"A1",X"28",X"08",X"DD",X"7E",X"05",X"BA",X"30",
		X"02",X"57",X"58",X"D5",X"11",X"09",X"00",X"DD",X"19",X"D1",X"23",X"04",X"78",X"FE",X"06",X"20",
		X"E6",X"C1",X"7A",X"B8",X"28",X"02",X"30",X"22",X"21",X"20",X"83",X"79",X"CD",X"BC",X"0F",X"4E",
		X"6B",X"26",X"00",X"54",X"5D",X"29",X"29",X"29",X"19",X"EB",X"DD",X"21",X"BC",X"82",X"DD",X"19",
		X"DD",X"71",X"04",X"DD",X"70",X"05",X"AF",X"DD",X"77",X"03",X"E1",X"C9",X"DD",X"21",X"BC",X"82",
		X"06",X"00",X"DD",X"7E",X"04",X"DD",X"BE",X"03",X"28",X"49",X"DD",X"77",X"03",X"DD",X"36",X"02",
		X"01",X"26",X"00",X"DD",X"6E",X"04",X"29",X"54",X"5D",X"19",X"19",X"11",X"BC",X"13",X"19",X"5E",
		X"23",X"56",X"DD",X"E5",X"E5",X"EB",X"11",X"CB",X"08",X"D5",X"E9",X"E1",X"DD",X"E1",X"23",X"7E",
		X"DD",X"77",X"00",X"23",X"7E",X"DD",X"77",X"01",X"DD",X"7E",X"04",X"FE",X"00",X"28",X"14",X"23",
		X"23",X"7E",X"FE",X"FF",X"28",X"0D",X"DD",X"E5",X"57",X"2B",X"5E",X"EB",X"11",X"F1",X"08",X"D5",
		X"E9",X"DD",X"E1",X"11",X"09",X"00",X"DD",X"19",X"04",X"78",X"FE",X"06",X"20",X"A4",X"C9",X"50",
		X"1E",X"36",X"CD",X"C1",X"0F",X"11",X"EE",X"0F",X"19",X"E5",X"FD",X"E1",X"DD",X"E3",X"DD",X"CB",
		X"00",X"46",X"20",X"10",X"FD",X"7E",X"09",X"2F",X"4F",X"FD",X"5E",X"06",X"FD",X"56",X"07",X"1A",
		X"B1",X"12",X"18",X"0B",X"FD",X"5E",X"06",X"FD",X"56",X"07",X"1A",X"FD",X"A6",X"09",X"12",X"DD",
		X"CB",X"00",X"66",X"20",X"0A",X"FD",X"7E",X"08",X"2F",X"4F",X"1A",X"B1",X"12",X"18",X"05",X"1A",
		X"FD",X"A6",X"08",X"12",X"DD",X"4E",X"01",X"FD",X"7E",X"14",X"FE",X"0F",X"20",X"0A",X"79",X"CB",
		X"27",X"CB",X"27",X"CB",X"27",X"CB",X"27",X"4F",X"FD",X"5E",X"12",X"FD",X"56",X"13",X"1A",X"FD",
		X"A6",X"14",X"B1",X"12",X"DD",X"7E",X"02",X"4F",X"FE",X"FF",X"28",X"2F",X"26",X"00",X"68",X"5D",
		X"54",X"29",X"29",X"29",X"19",X"11",X"BC",X"82",X"19",X"11",X"01",X"90",X"3E",X"06",X"CD",X"BC",
		X"0F",X"1A",X"E6",X"7F",X"77",X"23",X"FD",X"E5",X"D1",X"EB",X"79",X"CD",X"BC",X"0F",X"7E",X"12",
		X"23",X"13",X"66",X"6F",X"EB",X"72",X"21",X"03",X"90",X"7E",X"12",X"DD",X"E5",X"E1",X"1E",X"03",
		X"16",X"00",X"19",X"D9",X"FD",X"E5",X"D1",X"D9",X"7E",X"FE",X"FF",X"28",X"12",X"D9",X"62",X"6B",
		X"CD",X"BC",X"0F",X"4E",X"23",X"46",X"D9",X"23",X"7E",X"D9",X"02",X"D9",X"23",X"18",X"E9",X"23",
		X"D1",X"E5",X"C9",X"DD",X"E1",X"48",X"DD",X"5E",X"00",X"CD",X"D0",X"0F",X"DD",X"5E",X"01",X"FD",
		X"E5",X"16",X"00",X"FD",X"19",X"FD",X"7E",X"00",X"77",X"23",X"FD",X"7E",X"01",X"77",X"FD",X"E1",
		X"DD",X"5E",X"02",X"FD",X"E5",X"FD",X"19",X"FD",X"7E",X"00",X"23",X"77",X"23",X"FD",X"7E",X"01",
		X"77",X"1E",X"03",X"DD",X"19",X"FD",X"E1",X"DD",X"E5",X"C9",X"DD",X"E1",X"FD",X"E5",X"E1",X"16",
		X"00",X"DD",X"5E",X"01",X"19",X"E5",X"48",X"DD",X"5E",X"00",X"CD",X"D0",X"0F",X"16",X"00",X"1E",
		X"02",X"19",X"D1",X"1A",X"77",X"13",X"23",X"1A",X"77",X"16",X"00",X"1E",X"02",X"DD",X"19",X"DD",
		X"E5",X"C9",X"DD",X"E1",X"DD",X"5E",X"00",X"48",X"CD",X"D0",X"0F",X"EB",X"21",X"0D",X"00",X"19",
		X"FD",X"7E",X"00",X"77",X"FD",X"7E",X"01",X"23",X"77",X"21",X"0F",X"00",X"19",X"FD",X"7E",X"0A",
		X"77",X"FD",X"7E",X"0B",X"23",X"77",X"DD",X"23",X"DD",X"E5",X"C9",X"DD",X"E1",X"26",X"00",X"68",
		X"29",X"54",X"5D",X"29",X"29",X"19",X"E5",X"DD",X"6E",X"00",X"26",X"00",X"54",X"5D",X"29",X"29",
		X"19",X"D1",X"19",X"11",X"44",X"82",X"19",X"DD",X"5E",X"01",X"16",X"00",X"FD",X"E5",X"FD",X"19",
		X"FD",X"7E",X"00",X"77",X"23",X"FD",X"7E",X"01",X"77",X"1E",X"02",X"19",X"FD",X"E1",X"FD",X"E5",
		X"DD",X"5E",X"02",X"FD",X"19",X"FD",X"7E",X"01",X"77",X"2B",X"FD",X"7E",X"00",X"77",X"23",X"23",
		X"72",X"1E",X"03",X"DD",X"19",X"FD",X"E1",X"DD",X"E5",X"C9",X"DD",X"E1",X"21",X"04",X"83",X"16",
		X"00",X"DD",X"7E",X"00",X"B7",X"28",X"03",X"1E",X"04",X"19",X"DD",X"5E",X"01",X"FD",X"E5",X"FD",
		X"19",X"FD",X"7E",X"00",X"77",X"23",X"FD",X"7E",X"01",X"77",X"23",X"DD",X"7E",X"02",X"77",X"23",
		X"DD",X"7E",X"03",X"77",X"1E",X"04",X"DD",X"19",X"FD",X"E1",X"DD",X"E5",X"C9",X"DD",X"E1",X"FD",
		X"E5",X"E1",X"DD",X"5E",X"00",X"16",X"00",X"19",X"E5",X"68",X"26",X"00",X"54",X"5D",X"29",X"19",
		X"11",X"F2",X"82",X"19",X"D1",X"1A",X"77",X"13",X"23",X"1A",X"77",X"DD",X"23",X"DD",X"E5",X"C9",
		X"06",X"06",X"11",X"09",X"00",X"DD",X"21",X"BC",X"82",X"DD",X"7E",X"01",X"FE",X"FF",X"28",X"13",
		X"DD",X"4E",X"02",X"21",X"0C",X"0B",X"E5",X"DD",X"6E",X"00",X"67",X"E9",X"11",X"09",X"00",X"DD",
		X"36",X"02",X"00",X"DD",X"19",X"10",X"E2",X"C9",X"FD",X"E1",X"C5",X"3E",X"06",X"90",X"4F",X"FD",
		X"5E",X"02",X"CD",X"D0",X"0F",X"C1",X"C5",X"E5",X"DD",X"E3",X"79",X"FE",X"00",X"28",X"33",X"DD",
		X"6E",X"00",X"DD",X"66",X"01",X"DD",X"5E",X"02",X"DD",X"56",X"03",X"7E",X"12",X"FD",X"CB",X"03",
		X"4E",X"28",X"04",X"23",X"13",X"7E",X"12",X"FD",X"7E",X"06",X"DD",X"77",X"04",X"FD",X"7E",X"05",
		X"DD",X"77",X"05",X"AF",X"DD",X"77",X"06",X"FD",X"7E",X"04",X"DD",X"77",X"07",X"DD",X"E1",X"C3",
		X"20",X"0C",X"DD",X"35",X"04",X"28",X"05",X"DD",X"E1",X"C3",X"20",X"0C",X"FD",X"46",X"03",X"CB",
		X"48",X"26",X"00",X"DD",X"6E",X"06",X"54",X"5D",X"20",X"04",X"0E",X"03",X"18",X"03",X"0E",X"04",
		X"29",X"19",X"19",X"16",X"00",X"1E",X"05",X"19",X"EB",X"FD",X"E5",X"FD",X"19",X"DD",X"6E",X"00",
		X"DD",X"66",X"01",X"DD",X"5E",X"02",X"DD",X"56",X"03",X"CB",X"48",X"20",X"07",X"FD",X"7E",X"02",
		X"86",X"12",X"18",X"10",X"C5",X"4E",X"23",X"46",X"FD",X"6E",X"02",X"FD",X"66",X"03",X"09",X"C1",
		X"EB",X"73",X"23",X"72",X"DD",X"35",X"05",X"20",X"5D",X"DD",X"34",X"06",X"16",X"00",X"59",X"FD",
		X"19",X"FD",X"7E",X"00",X"FE",X"00",X"20",X"3C",X"DD",X"7E",X"07",X"FE",X"00",X"28",X"1D",X"FE",
		X"FF",X"28",X"03",X"DD",X"35",X"07",X"AF",X"DD",X"77",X"06",X"FD",X"E1",X"FD",X"7E",X"05",X"DD",
		X"77",X"05",X"FD",X"7E",X"06",X"DD",X"77",X"04",X"DD",X"E1",X"18",X"34",X"FD",X"E1",X"DD",X"E1",
		X"C1",X"3E",X"06",X"90",X"21",X"5B",X"11",X"16",X"00",X"5F",X"19",X"3A",X"1F",X"83",X"B6",X"32",
		X"1F",X"83",X"18",X"1D",X"FD",X"7E",X"01",X"DD",X"77",X"04",X"FD",X"7E",X"00",X"DD",X"77",X"05",
		X"FD",X"E1",X"DD",X"E1",X"18",X"0A",X"FD",X"7E",X"01",X"DD",X"77",X"04",X"FD",X"E1",X"DD",X"E1",
		X"C1",X"FD",X"6E",X"00",X"FD",X"66",X"01",X"E5",X"C9",X"FD",X"E1",X"C5",X"3E",X"06",X"90",X"4F",
		X"FD",X"5E",X"02",X"CD",X"D0",X"0F",X"C1",X"E5",X"DD",X"E3",X"79",X"FE",X"00",X"28",X"2A",X"FD",
		X"7E",X"06",X"DD",X"5E",X"02",X"DD",X"56",X"03",X"12",X"FD",X"CB",X"03",X"4E",X"28",X"05",X"13",
		X"FD",X"7E",X"07",X"12",X"FD",X"7E",X"05",X"DD",X"77",X"04",X"AF",X"DD",X"77",X"06",X"FD",X"7E",
		X"04",X"DD",X"77",X"07",X"DD",X"E1",X"C3",X"FD",X"0C",X"DD",X"35",X"04",X"28",X"05",X"DD",X"E1",
		X"C3",X"FD",X"0C",X"DD",X"34",X"06",X"C5",X"FD",X"46",X"03",X"CB",X"48",X"26",X"00",X"DD",X"6E",
		X"06",X"54",X"5D",X"29",X"28",X"01",X"19",X"FD",X"E5",X"16",X"00",X"1E",X"05",X"19",X"EB",X"FD",
		X"19",X"FD",X"7E",X"00",X"FE",X"00",X"28",X"1D",X"DD",X"77",X"04",X"FD",X"7E",X"01",X"DD",X"5E",
		X"02",X"DD",X"56",X"03",X"12",X"CB",X"48",X"28",X"05",X"FD",X"7E",X"02",X"13",X"12",X"FD",X"E1",
		X"C1",X"DD",X"E1",X"18",X"48",X"DD",X"7E",X"07",X"FE",X"00",X"28",X"2B",X"FE",X"FF",X"28",X"03",
		X"DD",X"35",X"07",X"AF",X"DD",X"77",X"06",X"FD",X"E1",X"FD",X"7E",X"05",X"DD",X"77",X"04",X"FD",
		X"7E",X"06",X"DD",X"5E",X"02",X"DD",X"56",X"03",X"12",X"CB",X"48",X"28",X"05",X"FD",X"7E",X"07",
		X"13",X"12",X"C1",X"DD",X"E1",X"18",X"16",X"FD",X"E1",X"C1",X"DD",X"E1",X"3E",X"06",X"90",X"21",
		X"5B",X"11",X"16",X"00",X"5F",X"19",X"3A",X"1F",X"83",X"B6",X"32",X"1F",X"83",X"FD",X"6E",X"00",
		X"FD",X"66",X"01",X"E5",X"C9",X"FD",X"E1",X"C5",X"3E",X"06",X"90",X"4F",X"FD",X"5E",X"02",X"CD",
		X"D0",X"0F",X"C1",X"E5",X"DD",X"E3",X"79",X"FE",X"00",X"28",X"0C",X"FD",X"7E",X"03",X"DD",X"77",
		X"00",X"CD",X"27",X"0E",X"C3",X"DA",X"0D",X"DD",X"35",X"0C",X"C2",X"DA",X"0D",X"DD",X"5E",X"09",
		X"DD",X"56",X"0A",X"21",X"02",X"00",X"19",X"7E",X"DD",X"6E",X"0F",X"DD",X"66",X"10",X"86",X"77",
		X"DD",X"35",X"0B",X"C2",X"D2",X"0D",X"21",X"03",X"00",X"19",X"DD",X"75",X"09",X"DD",X"74",X"0A",
		X"7E",X"FE",X"00",X"20",X"70",X"DD",X"5E",X"05",X"DD",X"56",X"06",X"21",X"03",X"00",X"19",X"DD",
		X"75",X"05",X"DD",X"74",X"06",X"7E",X"FE",X"00",X"20",X"54",X"DD",X"6E",X"01",X"DD",X"66",X"02",
		X"23",X"23",X"DD",X"75",X"01",X"DD",X"74",X"02",X"23",X"7E",X"FE",X"00",X"20",X"26",X"DD",X"7E",
		X"00",X"FE",X"00",X"20",X"13",X"3E",X"06",X"90",X"21",X"5B",X"11",X"16",X"00",X"5F",X"19",X"3A",
		X"1F",X"83",X"B6",X"32",X"1F",X"83",X"18",X"42",X"FE",X"FF",X"28",X"03",X"DD",X"35",X"00",X"CD",
		X"27",X"0E",X"18",X"36",X"DD",X"6E",X"01",X"DD",X"66",X"02",X"5E",X"23",X"56",X"DD",X"73",X"03",
		X"DD",X"72",X"04",X"DD",X"73",X"05",X"DD",X"72",X"06",X"CD",X"E4",X"0D",X"18",X"1C",X"54",X"5D",
		X"CD",X"E4",X"0D",X"18",X"15",X"DD",X"77",X"0B",X"11",X"01",X"00",X"19",X"7E",X"DD",X"77",X"0C",
		X"18",X"08",X"21",X"01",X"00",X"19",X"7E",X"DD",X"77",X"0C",X"DD",X"E1",X"FD",X"6E",X"00",X"FD",
		X"66",X"01",X"E5",X"C9",X"13",X"DD",X"6E",X"0D",X"DD",X"66",X"0E",X"1A",X"77",X"13",X"23",X"1A",
		X"77",X"1B",X"1B",X"26",X"00",X"1A",X"6F",X"11",X"00",X"12",X"19",X"5E",X"23",X"56",X"DD",X"73",
		X"07",X"DD",X"72",X"08",X"21",X"00",X"00",X"19",X"7E",X"DD",X"6E",X"0F",X"DD",X"66",X"10",X"77",
		X"21",X"01",X"00",X"19",X"DD",X"75",X"09",X"DD",X"74",X"0A",X"7E",X"DD",X"77",X"0B",X"11",X"01",
		X"00",X"19",X"7E",X"DD",X"77",X"0C",X"C9",X"FD",X"E5",X"E1",X"11",X"04",X"00",X"19",X"DD",X"75",
		X"01",X"DD",X"74",X"02",X"FD",X"7E",X"04",X"DD",X"77",X"03",X"DD",X"77",X"05",X"6F",X"FD",X"7E",
		X"05",X"DD",X"77",X"04",X"DD",X"77",X"06",X"67",X"23",X"DD",X"5E",X"0D",X"DD",X"56",X"0E",X"7E",
		X"12",X"23",X"13",X"7E",X"12",X"2B",X"2B",X"16",X"00",X"5E",X"21",X"00",X"12",X"19",X"5E",X"DD",
		X"73",X"07",X"23",X"56",X"DD",X"72",X"08",X"21",X"00",X"00",X"19",X"7E",X"DD",X"6E",X"0F",X"DD",
		X"66",X"10",X"77",X"21",X"01",X"00",X"19",X"DD",X"75",X"09",X"DD",X"74",X"0A",X"7E",X"DD",X"77",
		X"0B",X"11",X"01",X"00",X"19",X"7E",X"DD",X"77",X"0C",X"C9",X"3E",X"06",X"90",X"6F",X"26",X"00",
		X"54",X"5D",X"29",X"19",X"FD",X"21",X"F2",X"82",X"EB",X"FD",X"19",X"FD",X"6E",X"00",X"FD",X"66",
		X"01",X"FD",X"7E",X"02",X"96",X"D8",X"3E",X"01",X"77",X"C9",X"3E",X"06",X"90",X"6F",X"26",X"00",
		X"29",X"54",X"5D",X"29",X"29",X"19",X"11",X"44",X"82",X"19",X"FD",X"E1",X"E5",X"26",X"00",X"FD",
		X"6E",X"02",X"54",X"5D",X"29",X"29",X"19",X"DD",X"E3",X"EB",X"DD",X"19",X"DD",X"7E",X"04",X"FE",
		X"00",X"28",X"05",X"DD",X"35",X"04",X"18",X"35",X"3A",X"71",X"83",X"C5",X"4F",X"E6",X"33",X"EA",
		X"E3",X"0E",X"37",X"79",X"1F",X"32",X"71",X"83",X"47",X"FD",X"7E",X"03",X"DD",X"77",X"04",X"DD",
		X"6E",X"00",X"DD",X"66",X"01",X"5E",X"16",X"00",X"21",X"52",X"11",X"19",X"4E",X"79",X"A0",X"47",
		X"79",X"2F",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"4E",X"A1",X"B0",X"77",X"C1",X"DD",X"E1",X"FD",
		X"6E",X"00",X"FD",X"66",X"01",X"E5",X"C9",X"C5",X"3E",X"06",X"90",X"47",X"57",X"1E",X"36",X"CD",
		X"C1",X"0F",X"EB",X"FD",X"21",X"EE",X"0F",X"FD",X"19",X"16",X"00",X"58",X"21",X"3E",X"82",X"19",
		X"FD",X"7E",X"14",X"4F",X"FE",X"0F",X"7E",X"20",X"17",X"CB",X"27",X"CB",X"27",X"CB",X"27",X"CB",
		X"27",X"E6",X"F0",X"47",X"FD",X"6E",X"12",X"FD",X"66",X"13",X"7E",X"A1",X"B0",X"77",X"C1",X"C9",
		X"E6",X"0F",X"18",X"EF",X"FD",X"E1",X"21",X"04",X"83",X"FD",X"7E",X"00",X"B7",X"28",X"05",X"16",
		X"00",X"1E",X"04",X"19",X"5E",X"23",X"56",X"1A",X"17",X"17",X"17",X"17",X"E6",X"70",X"23",X"5E",
		X"23",X"56",X"67",X"1A",X"E6",X"8F",X"B4",X"12",X"1E",X"01",X"16",X"00",X"FD",X"19",X"FD",X"E5",
		X"C9",X"01",X"1F",X"00",X"21",X"00",X"80",X"11",X"20",X"80",X"09",X"EB",X"09",X"06",X"0F",X"DD",
		X"21",X"00",X"B0",X"1A",X"BE",X"28",X"07",X"77",X"DD",X"70",X"00",X"32",X"02",X"B0",X"1B",X"2B",
		X"05",X"F2",X"93",X"0F",X"06",X"0F",X"DD",X"21",X"00",X"A0",X"1A",X"BE",X"28",X"07",X"77",X"DD",
		X"70",X"00",X"32",X"02",X"A0",X"1B",X"2B",X"05",X"F2",X"AA",X"0F",X"C9",X"85",X"6F",X"D0",X"24",
		X"C9",X"C5",X"42",X"21",X"00",X"00",X"54",X"78",X"B7",X"28",X"03",X"19",X"10",X"FD",X"C1",X"C9",
		X"21",X"6D",X"11",X"16",X"00",X"19",X"56",X"21",X"61",X"11",X"79",X"CB",X"27",X"5F",X"7A",X"16",
		X"00",X"19",X"5E",X"23",X"56",X"6F",X"26",X"00",X"19",X"11",X"40",X"80",X"19",X"C9",X"00",X"80",
		X"01",X"80",X"06",X"80",X"07",X"80",X"F7",X"FE",X"08",X"80",X"0B",X"80",X"0C",X"80",X"0D",X"80",
		X"0E",X"80",X"F0",X"00",X"48",X"80",X"59",X"80",X"6A",X"80",X"7B",X"80",X"8C",X"80",X"44",X"80",
		X"55",X"80",X"66",X"80",X"77",X"80",X"88",X"80",X"3E",X"82",X"F4",X"82",X"49",X"80",X"5A",X"80",
		X"6B",X"80",X"7C",X"80",X"02",X"80",X"03",X"80",X"06",X"80",X"07",X"80",X"EF",X"FD",X"09",X"80",
		X"0B",X"80",X"0C",X"80",X"0D",X"80",X"0E",X"80",X"0F",X"00",X"9D",X"80",X"AE",X"80",X"BF",X"80",
		X"D0",X"80",X"E1",X"80",X"99",X"80",X"AA",X"80",X"BB",X"80",X"CC",X"80",X"DD",X"80",X"3F",X"82",
		X"F7",X"82",X"9E",X"80",X"AF",X"80",X"C0",X"80",X"D1",X"80",X"04",X"80",X"05",X"80",X"06",X"80",
		X"07",X"80",X"DF",X"FB",X"0A",X"80",X"0B",X"80",X"0C",X"80",X"0D",X"80",X"0F",X"80",X"F0",X"00",
		X"F2",X"80",X"03",X"81",X"14",X"81",X"25",X"81",X"36",X"81",X"EE",X"80",X"FF",X"80",X"10",X"81",
		X"21",X"81",X"32",X"81",X"40",X"82",X"FA",X"82",X"F3",X"80",X"04",X"81",X"15",X"81",X"26",X"81",
		X"10",X"80",X"11",X"80",X"16",X"80",X"17",X"80",X"F7",X"FE",X"18",X"80",X"1B",X"80",X"1C",X"80",
		X"1D",X"80",X"1E",X"80",X"F0",X"00",X"47",X"81",X"58",X"81",X"69",X"81",X"7A",X"81",X"8B",X"81",
		X"43",X"81",X"54",X"81",X"65",X"81",X"76",X"81",X"87",X"81",X"41",X"82",X"FD",X"82",X"48",X"81",
		X"59",X"81",X"6A",X"81",X"7B",X"81",X"12",X"80",X"13",X"80",X"16",X"80",X"17",X"80",X"EF",X"FD",
		X"19",X"80",X"1B",X"80",X"1C",X"80",X"1D",X"80",X"1E",X"80",X"0F",X"00",X"9C",X"81",X"AD",X"81",
		X"BE",X"81",X"CF",X"81",X"E0",X"81",X"98",X"81",X"A9",X"81",X"BA",X"81",X"CB",X"81",X"DC",X"81",
		X"42",X"82",X"00",X"83",X"9D",X"81",X"AE",X"81",X"BF",X"81",X"D0",X"81",X"14",X"80",X"15",X"80",
		X"16",X"80",X"17",X"80",X"DF",X"FB",X"1A",X"80",X"1B",X"80",X"1C",X"80",X"1D",X"80",X"1F",X"80",
		X"F0",X"00",X"F1",X"81",X"02",X"82",X"13",X"82",X"24",X"82",X"35",X"82",X"ED",X"81",X"FE",X"81",
		X"0F",X"82",X"20",X"82",X"31",X"82",X"43",X"82",X"03",X"83",X"F2",X"81",X"03",X"82",X"14",X"82",
		X"25",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"70",X"00",X"01",X"03",X"07",X"0F",X"1F",X"3F",X"7F",X"FF",X"01",X"02",X"04",X"08",X"10",
		X"20",X"00",X"00",X"55",X"00",X"AA",X"00",X"FF",X"00",X"54",X"01",X"A9",X"01",X"00",X"11",X"22",
		X"33",X"44",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"9E",X"16",X"A6",X"16",X"AE",X"16",X"B9",X"16",X"1D",X"2B",X"2B",X"2B",X"36",X"2B",X"44",
		X"2B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"18",X"00",
		X"00",X"00",X"00",X"00",X"01",X"06",X"00",X"00",X"00",X"00",X"00",X"01",X"49",X"00",X"00",X"00",
		X"00",X"00",X"01",X"27",X"00",X"00",X"00",X"00",X"00",X"00",X"49",X"00",X"00",X"00",X"00",X"00",
		X"01",X"15",X"00",X"00",X"00",X"00",X"00",X"01",X"09",X"0A",X"00",X"00",X"00",X"00",X"01",X"31",
		X"32",X"00",X"00",X"00",X"00",X"01",X"41",X"00",X"00",X"00",X"00",X"00",X"01",X"22",X"00",X"00",
		X"00",X"00",X"00",X"01",X"0C",X"0D",X"0E",X"00",X"00",X"00",X"00",X"0C",X"0D",X"0E",X"00",X"00",
		X"00",X"01",X"42",X"00",X"00",X"00",X"00",X"00",X"01",X"11",X"12",X"13",X"00",X"00",X"00",X"01",
		X"22",X"00",X"00",X"00",X"00",X"00",X"01",X"43",X"00",X"00",X"00",X"00",X"00",X"01",X"44",X"00",
		X"00",X"00",X"00",X"00",X"00",X"29",X"29",X"29",X"29",X"29",X"29",X"00",X"27",X"00",X"00",X"00",
		X"00",X"00",X"01",X"02",X"00",X"00",X"00",X"00",X"00",X"01",X"45",X"00",X"00",X"00",X"00",X"00",
		X"01",X"46",X"00",X"00",X"00",X"00",X"00",X"01",X"47",X"00",X"00",X"00",X"00",X"00",X"01",X"2B",
		X"00",X"00",X"00",X"00",X"00",X"01",X"1C",X"21",X"1D",X"1E",X"1F",X"20",X"01",X"2D",X"00",X"00",
		X"00",X"00",X"00",X"01",X"28",X"00",X"00",X"00",X"00",X"00",X"01",X"23",X"23",X"23",X"23",X"23",
		X"23",X"01",X"48",X"4A",X"00",X"00",X"00",X"00",X"01",X"4A",X"4B",X"00",X"00",X"00",X"00",X"01",
		X"2E",X"00",X"00",X"00",X"00",X"00",X"01",X"4A",X"4C",X"00",X"00",X"00",X"00",X"01",X"37",X"37",
		X"37",X"37",X"37",X"37",X"00",X"37",X"37",X"37",X"37",X"37",X"37",X"01",X"29",X"00",X"00",X"00",
		X"00",X"00",X"01",X"3C",X"00",X"00",X"00",X"00",X"00",X"01",X"04",X"00",X"00",X"00",X"00",X"00",
		X"00",X"1C",X"21",X"1D",X"1E",X"1F",X"20",X"01",X"26",X"00",X"00",X"00",X"00",X"00",X"01",X"3D",
		X"00",X"00",X"00",X"00",X"00",X"01",X"2C",X"00",X"00",X"00",X"00",X"00",X"01",X"24",X"24",X"24",
		X"24",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"40",X"40",X"00",X"00",X"00",
		X"00",X"01",X"2F",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"00",X"00",X"00",X"00",X"00",X"01",
		X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"4F",X"50",
		X"51",X"52",X"53",X"54",X"01",X"35",X"00",X"00",X"00",X"00",X"00",X"01",X"55",X"56",X"57",X"58",
		X"00",X"00",X"01",X"59",X"5A",X"00",X"00",X"00",X"00",X"01",X"10",X"00",X"00",X"00",X"00",X"00",
		X"01",X"14",X"00",X"00",X"00",X"00",X"00",X"01",X"16",X"17",X"16",X"17",X"16",X"17",X"01",X"19",
		X"00",X"00",X"00",X"00",X"00",X"01",X"05",X"00",X"00",X"00",X"00",X"00",X"94",X"16",X"FF",X"FF",
		X"FF",X"FF",X"C8",X"16",X"DC",X"16",X"D6",X"16",X"FE",X"16",X"16",X"17",X"0C",X"17",X"83",X"17",
		X"9B",X"17",X"91",X"17",X"D9",X"17",X"F1",X"17",X"E7",X"17",X"A1",X"24",X"BC",X"24",X"AF",X"24",
		X"5E",X"18",X"77",X"18",X"6A",X"18",X"98",X"18",X"98",X"18",X"98",X"18",X"98",X"18",X"98",X"18",
		X"98",X"18",X"98",X"18",X"B3",X"18",X"A6",X"18",X"98",X"18",X"D0",X"18",X"A6",X"18",X"E1",X"18",
		X"E1",X"18",X"E1",X"18",X"E1",X"18",X"FC",X"18",X"EF",X"18",X"1B",X"19",X"29",X"19",X"EF",X"18",
		X"48",X"19",X"56",X"19",X"EF",X"18",X"75",X"19",X"92",X"19",X"85",X"19",X"A8",X"19",X"C3",X"19",
		X"B6",X"19",X"E4",X"19",X"FF",X"19",X"F2",X"19",X"1B",X"1A",X"29",X"1A",X"F2",X"19",X"45",X"1A",
		X"53",X"1A",X"F2",X"19",X"6F",X"1A",X"84",X"1A",X"7D",X"1A",X"A6",X"1A",X"C7",X"1A",X"B4",X"1A",
		X"FE",X"1A",X"21",X"1B",X"0E",X"1B",X"71",X"1B",X"21",X"1B",X"0E",X"1B",X"81",X"1B",X"96",X"1B",
		X"8F",X"1B",X"AC",X"1B",X"C5",X"1B",X"B8",X"1B",X"E6",X"1B",X"E6",X"1B",X"E6",X"1B",X"E6",X"1B",
		X"E6",X"1B",X"E6",X"1B",X"E6",X"1B",X"FF",X"1B",X"F4",X"1B",X"98",X"1C",X"AC",X"1C",X"A6",X"1C",
		X"FD",X"1D",X"11",X"1E",X"0B",X"1E",X"F3",X"1E",X"0C",X"1F",X"01",X"1F",X"79",X"20",X"92",X"20",
		X"87",X"20",X"E6",X"1B",X"36",X"21",X"F4",X"1B",X"93",X"21",X"BC",X"21",X"A3",X"21",X"E4",X"21",
		X"FF",X"21",X"F2",X"21",X"27",X"22",X"42",X"22",X"35",X"22",X"5F",X"22",X"74",X"22",X"6D",X"22",
		X"93",X"22",X"AE",X"22",X"A1",X"22",X"CA",X"22",X"EF",X"22",X"DC",X"22",X"21",X"23",X"44",X"23",
		X"31",X"23",X"7E",X"23",X"A7",X"23",X"94",X"23",X"CF",X"23",X"E4",X"23",X"DD",X"23",X"F4",X"23",
		X"02",X"24",X"DD",X"23",X"14",X"24",X"27",X"24",X"20",X"24",X"3A",X"24",X"4F",X"24",X"48",X"24",
		X"3A",X"24",X"6F",X"24",X"48",X"24",X"81",X"24",X"6F",X"24",X"48",X"24",X"61",X"24",X"8F",X"24",
		X"48",X"24",X"DA",X"24",X"F5",X"24",X"E8",X"24",X"13",X"25",X"2E",X"25",X"21",X"25",X"4C",X"25",
		X"4C",X"25",X"21",X"25",X"4C",X"25",X"4C",X"25",X"21",X"25",X"4C",X"25",X"67",X"25",X"5A",X"25",
		X"86",X"25",X"86",X"25",X"86",X"25",X"86",X"25",X"9B",X"25",X"94",X"25",X"AD",X"25",X"AD",X"25",
		X"AD",X"25",X"AD",X"25",X"C6",X"25",X"B9",X"25",X"AD",X"25",X"E3",X"25",X"B9",X"25",X"3B",X"26",
		X"F4",X"25",X"4B",X"26",X"F4",X"25",X"18",X"26",X"04",X"26",X"3B",X"26",X"56",X"26",X"4B",X"26",
		X"3B",X"26",X"23",X"27",X"4B",X"26",X"3B",X"26",X"23",X"27",X"4B",X"26",X"23",X"27",X"36",X"27",
		X"2F",X"27",X"49",X"27",X"4F",X"27",X"4C",X"27",X"56",X"27",X"5C",X"27",X"59",X"27",X"63",X"27",
		X"7E",X"27",X"71",X"27",X"A2",X"27",X"B7",X"27",X"B0",X"27",X"C9",X"27",X"DE",X"27",X"D7",X"27",
		X"09",X"28",X"1C",X"28",X"15",X"28",X"4A",X"28",X"49",X"27",X"49",X"27",X"4D",X"28",X"77",X"28",
		X"5D",X"28",X"BC",X"28",X"DF",X"28",X"CC",X"28",X"15",X"29",X"36",X"29",X"23",X"29",X"64",X"29",
		X"77",X"28",X"5D",X"28",X"72",X"29",X"77",X"28",X"5D",X"28",X"80",X"29",X"80",X"29",X"80",X"29",
		X"80",X"29",X"80",X"29",X"80",X"29",X"80",X"29",X"95",X"29",X"8E",X"29",X"A8",X"29",X"B6",X"29",
		X"8E",X"29",X"CB",X"29",X"D9",X"29",X"8E",X"29",X"EE",X"29",X"FC",X"29",X"8E",X"29",X"11",X"2A",
		X"1F",X"2A",X"8E",X"29",X"34",X"2A",X"42",X"2A",X"8E",X"29",X"5A",X"2A",X"69",X"2A",X"64",X"2A",
		X"5A",X"2A",X"74",X"2A",X"64",X"2A",X"5A",X"2A",X"7F",X"2A",X"64",X"2A",X"5A",X"2A",X"8A",X"2A",
		X"64",X"2A",X"4A",X"2B",X"59",X"2B",X"54",X"2B",X"4A",X"2B",X"64",X"2B",X"54",X"2B",X"00",X"00",
		X"1F",X"FE",X"A0",X"FA",X"A0",X"FA",X"BF",X"FA",X"BF",X"F0",X"1F",X"80",X"00",X"00",X"00",X"00",
		X"1F",X"80",X"1F",X"80",X"00",X"00",X"1F",X"C8",X"1F",X"C8",X"1F",X"C8",X"00",X"00",X"BF",X"FA",
		X"1F",X"C8",X"1F",X"C8",X"1F",X"C8",X"BF",X"F9",X"1F",X"F9",X"BF",X"FF",X"BF",X"FF",X"1F",X"FE",
		X"BF",X"C8",X"00",X"00",X"00",X"00",X"BF",X"FE",X"BF",X"FE",X"BF",X"FE",X"BF",X"FE",X"BF",X"FE",
		X"BF",X"FE",X"1F",X"E1",X"BF",X"FE",X"1F",X"E1",X"00",X"00",X"88",X"FF",X"1F",X"80",X"A0",X"F9",
		X"81",X"FF",X"00",X"00",X"00",X"00",X"BF",X"FF",X"1F",X"F9",X"1F",X"F9",X"BF",X"FA",X"BF",X"F9",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BF",X"FB",X"00",X"00",X"BF",X"FA",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"81",X"FE",X"BF",X"FE",X"00",X"00",X"00",X"00",X"BF",X"FA",
		X"1F",X"80",X"1F",X"80",X"1F",X"80",X"1F",X"80",X"1F",X"80",X"1F",X"80",X"00",X"00",X"1F",X"F9",
		X"A0",X"0A",X"1F",X"F9",X"1F",X"F9",X"1F",X"F9",X"00",X"00",X"00",X"00",X"81",X"32",X"82",X"32",
		X"84",X"32",X"88",X"32",X"90",X"32",X"A0",X"32",X"9E",X"55",X"9E",X"55",X"9E",X"55",X"9E",X"55",
		X"BF",X"FE",X"BF",X"FE",X"CD",X"FF",X"08",X"00",X"00",X"FF",X"0A",X"00",X"FF",X"C9",X"07",X"05",
		X"01",X"01",X"01",X"02",X"F8",X"00",X"07",X"05",X"01",X"01",X"01",X"09",X"F8",X"00",X"04",X"08",
		X"01",X"01",X"01",X"20",X"00",X"02",X"01",X"FC",X"00",X"04",X"08",X"01",X"01",X"01",X"66",X"00",
		X"02",X"01",X"FC",X"00",X"00",X"00",X"00",X"00",X"CD",X"FF",X"08",X"01",X"08",X"FF",X"0A",X"0D",
		X"00",X"52",X"02",X"01",X"FF",X"C9",X"CD",X"FA",X"09",X"00",X"00",X"C9",X"CD",X"29",X"0C",X"FD",
		X"16",X"00",X"02",X"00",X"0A",X"70",X"00",X"0A",X"90",X"00",X"0A",X"60",X"00",X"0A",X"A0",X"00",
		X"0A",X"50",X"00",X"0A",X"B0",X"00",X"0A",X"40",X"00",X"0A",X"C0",X"00",X"00",X"C9",X"CD",X"FF",
		X"08",X"01",X"08",X"2C",X"0A",X"0F",X"00",X"52",X"02",X"01",X"FF",X"C9",X"CD",X"FA",X"09",X"00",
		X"00",X"CD",X"CD",X"0A",X"20",X"C9",X"CD",X"29",X"0C",X"7F",X"17",X"00",X"02",X"FF",X"7F",X"FB",
		X"04",X"7F",X"01",X"00",X"7F",X"B4",X"04",X"7F",X"01",X"00",X"7F",X"FB",X"04",X"7F",X"01",X"00",
		X"7F",X"38",X"02",X"7F",X"01",X"00",X"7F",X"FB",X"04",X"7F",X"01",X"00",X"7F",X"B4",X"04",X"7F",
		X"01",X"00",X"7F",X"FB",X"04",X"7F",X"01",X"00",X"7F",X"DE",X"01",X"7F",X"01",X"00",X"7F",X"FB",
		X"04",X"7F",X"01",X"00",X"7F",X"B4",X"04",X"7F",X"01",X"00",X"7F",X"FB",X"04",X"7F",X"01",X"00",
		X"7F",X"FA",X"01",X"7F",X"01",X"00",X"7F",X"FB",X"04",X"7F",X"01",X"00",X"7F",X"B4",X"04",X"7F",
		X"01",X"00",X"7F",X"FB",X"04",X"7F",X"01",X"00",X"7F",X"C3",X"01",X"7F",X"01",X"00",X"00",X"CD",
		X"8A",X"0E",X"C9",X"CD",X"FF",X"08",X"01",X"08",X"2C",X"0A",X"0F",X"00",X"52",X"02",X"01",X"FF",
		X"C9",X"CD",X"FA",X"09",X"00",X"00",X"CD",X"CD",X"0A",X"20",X"C9",X"CD",X"29",X"0C",X"D5",X"17",
		X"00",X"02",X"FF",X"7F",X"98",X"05",X"7F",X"01",X"00",X"7F",X"68",X"09",X"7F",X"01",X"00",X"7F",
		X"98",X"05",X"7F",X"01",X"00",X"7F",X"CC",X"02",X"7F",X"01",X"00",X"7F",X"98",X"05",X"7F",X"01",
		X"00",X"7F",X"61",X"08",X"7F",X"01",X"00",X"7F",X"98",X"05",X"7F",X"01",X"00",X"7F",X"F6",X"02",
		X"7F",X"01",X"00",X"00",X"00",X"CD",X"8A",X"0E",X"C9",X"CD",X"FF",X"08",X"01",X"08",X"2C",X"0A",
		X"0F",X"00",X"52",X"02",X"01",X"FF",X"C9",X"CD",X"FA",X"09",X"00",X"00",X"CD",X"CD",X"0A",X"20",
		X"C9",X"CD",X"29",X"0C",X"5A",X"18",X"00",X"02",X"FF",X"7F",X"7F",X"02",X"7F",X"01",X"00",X"7F",
		X"5A",X"02",X"7F",X"01",X"00",X"7F",X"7F",X"02",X"7F",X"01",X"00",X"7F",X"38",X"02",X"7F",X"01",
		X"00",X"7F",X"7F",X"02",X"7F",X"01",X"00",X"7F",X"5A",X"02",X"7F",X"01",X"00",X"7F",X"7F",X"02",
		X"7F",X"01",X"00",X"7F",X"DE",X"01",X"7F",X"01",X"00",X"7F",X"7F",X"02",X"7F",X"01",X"00",X"7F",
		X"5A",X"02",X"7F",X"01",X"00",X"7F",X"7F",X"02",X"7F",X"01",X"00",X"7F",X"FA",X"01",X"7F",X"01",
		X"00",X"7F",X"7F",X"02",X"7F",X"01",X"00",X"7F",X"5A",X"02",X"7F",X"01",X"00",X"7F",X"7F",X"02",
		X"7F",X"01",X"00",X"7F",X"C3",X"01",X"7F",X"01",X"00",X"00",X"CD",X"8A",X"0E",X"C9",X"CD",X"FF",
		X"08",X"01",X"08",X"00",X"0A",X"0F",X"02",X"00",X"FF",X"C9",X"CD",X"C3",X"09",X"00",X"00",X"00",
		X"CD",X"C3",X"09",X"01",X"0A",X"0A",X"C9",X"CD",X"18",X"0B",X"88",X"18",X"00",X"02",X"FF",X"05",
		X"01",X"F7",X"FF",X"05",X"01",X"09",X"00",X"00",X"CD",X"18",X"0B",X"97",X"18",X"01",X"01",X"00",
		X"0F",X"01",X"00",X"0F",X"03",X"FF",X"00",X"C9",X"CD",X"FF",X"08",X"01",X"01",X"FF",X"0A",X"0C",
		X"00",X"00",X"02",X"00",X"FF",X"C9",X"CD",X"C3",X"09",X"00",X"00",X"00",X"CD",X"C3",X"09",X"01",
		X"0A",X"0A",X"C9",X"CD",X"18",X"0B",X"C0",X"18",X"00",X"02",X"00",X"50",X"01",X"10",X"00",X"00",
		X"CD",X"18",X"0B",X"CF",X"18",X"01",X"01",X"00",X"01",X"50",X"00",X"0A",X"01",X"FF",X"00",X"C9",
		X"CD",X"18",X"0B",X"C0",X"18",X"00",X"02",X"00",X"01",X"03",X"00",X"00",X"50",X"01",X"10",X"00",
		X"00",X"CD",X"FF",X"08",X"01",X"05",X"FF",X"0A",X"0B",X"00",X"28",X"02",X"00",X"FF",X"C9",X"CD",
		X"C3",X"09",X"00",X"0A",X"0A",X"CD",X"C3",X"09",X"01",X"0A",X"0A",X"C9",X"CD",X"18",X"0B",X"0B",
		X"19",X"00",X"01",X"FF",X"01",X"02",X"01",X"01",X"02",X"FF",X"00",X"CD",X"18",X"0B",X"1A",X"19",
		X"01",X"01",X"FF",X"08",X"02",X"FF",X"01",X"01",X"08",X"00",X"C9",X"CD",X"FF",X"08",X"01",X"03",
		X"FF",X"0A",X"0B",X"00",X"3C",X"02",X"00",X"FF",X"C9",X"CD",X"18",X"0B",X"38",X"19",X"00",X"01",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"FF",X"00",X"CD",X"18",X"0B",X"47",X"19",X"01",X"01",X"FF",
		X"08",X"02",X"FF",X"01",X"01",X"08",X"00",X"C9",X"CD",X"FF",X"08",X"01",X"03",X"FF",X"0A",X"0B",
		X"00",X"50",X"02",X"00",X"FF",X"C9",X"CD",X"18",X"0B",X"65",X"19",X"00",X"01",X"FF",X"01",X"03",
		X"01",X"01",X"03",X"FF",X"00",X"CD",X"18",X"0B",X"74",X"19",X"01",X"01",X"FF",X"08",X"02",X"FF",
		X"01",X"01",X"08",X"00",X"C9",X"CD",X"FF",X"08",X"11",X"00",X"FF",X"04",X"1F",X"0A",X"0C",X"00",
		X"1C",X"02",X"01",X"FF",X"C9",X"CD",X"C3",X"09",X"00",X"2A",X"2A",X"CD",X"C3",X"09",X"01",X"0A",
		X"0A",X"C9",X"CD",X"18",X"0B",X"9E",X"19",X"00",X"01",X"00",X"0F",X"03",X"01",X"00",X"CD",X"18",
		X"0B",X"A7",X"19",X"01",X"01",X"00",X"00",X"C9",X"CD",X"FF",X"08",X"01",X"00",X"FF",X"00",X"EC",
		X"02",X"00",X"0A",X"0F",X"FF",X"C9",X"CD",X"C3",X"09",X"00",X"00",X"00",X"CD",X"C3",X"09",X"01",
		X"0A",X"0A",X"C9",X"CD",X"18",X"0B",X"D4",X"19",X"00",X"02",X"0F",X"01",X"02",X"9C",X"FF",X"01",
		X"02",X"74",X"00",X"00",X"CD",X"18",X"0B",X"E3",X"19",X"01",X"01",X"00",X"28",X"01",X"00",X"05",
		X"04",X"FD",X"00",X"C9",X"CD",X"FF",X"08",X"01",X"05",X"FF",X"0A",X"0B",X"00",X"28",X"02",X"00",
		X"FF",X"C9",X"CD",X"C3",X"09",X"00",X"0A",X"0A",X"CD",X"C3",X"09",X"01",X"0A",X"0A",X"C9",X"CD",
		X"18",X"0B",X"0E",X"1A",X"00",X"01",X"FF",X"01",X"02",X"01",X"01",X"02",X"FF",X"00",X"CD",X"18",
		X"0B",X"1A",X"1A",X"01",X"01",X"00",X"0B",X"05",X"FF",X"00",X"C9",X"CD",X"FF",X"08",X"01",X"05",
		X"FF",X"0A",X"0B",X"00",X"3C",X"02",X"00",X"FF",X"C9",X"CD",X"18",X"0B",X"38",X"1A",X"00",X"01",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"FF",X"00",X"CD",X"18",X"0B",X"44",X"1A",X"01",X"01",X"00",
		X"0B",X"05",X"FF",X"00",X"C9",X"CD",X"FF",X"08",X"01",X"03",X"FF",X"0A",X"0B",X"00",X"50",X"02",
		X"00",X"FF",X"C9",X"CD",X"18",X"0B",X"62",X"1A",X"00",X"01",X"FF",X"01",X"03",X"01",X"01",X"03",
		X"FF",X"00",X"CD",X"18",X"0B",X"6E",X"1A",X"01",X"01",X"00",X"0B",X"05",X"FF",X"00",X"C9",X"CD",
		X"FF",X"08",X"01",X"01",X"FF",X"0A",X"0F",X"02",X"00",X"00",X"4C",X"FF",X"C9",X"CD",X"C3",X"09",
		X"00",X"00",X"00",X"C9",X"CD",X"18",X"0B",X"A5",X"1A",X"00",X"02",X"03",X"03",X"02",X"F0",X"FF",
		X"03",X"02",X"10",X"00",X"01",X"01",X"A1",X"00",X"03",X"02",X"F0",X"FF",X"03",X"02",X"10",X"00",
		X"01",X"01",X"5F",X"FF",X"00",X"C9",X"CD",X"FF",X"08",X"10",X"0F",X"FF",X"2A",X"00",X"04",X"1F",
		X"0A",X"00",X"FF",X"C9",X"CD",X"C3",X"09",X"00",X"0A",X"0A",X"CD",X"C3",X"09",X"01",X"2A",X"2A",
		X"CD",X"C3",X"09",X"02",X"04",X"04",X"C9",X"CD",X"18",X"0B",X"D9",X"1A",X"00",X"01",X"00",X"0F",
		X"01",X"01",X"24",X"01",X"00",X"01",X"01",X"F1",X"00",X"CD",X"18",X"0B",X"E8",X"1A",X"01",X"01",
		X"00",X"0F",X"02",X"FF",X"01",X"0C",X"00",X"00",X"CD",X"18",X"0B",X"FA",X"1A",X"02",X"01",X"00",
		X"0F",X"02",X"FF",X"10",X"01",X"FF",X"01",X"01",X"1D",X"00",X"CD",X"17",X"0F",X"C9",X"CD",X"FF",
		X"08",X"01",X"01",X"FF",X"0A",X"0E",X"02",X"04",X"00",X"70",X"2A",X"01",X"FF",X"C9",X"CD",X"C3",
		X"09",X"00",X"0A",X"0A",X"CD",X"C3",X"09",X"01",X"02",X"02",X"CD",X"C3",X"09",X"02",X"2A",X"2A",
		X"C9",X"CD",X"18",X"0B",X"30",X"1B",X"00",X"01",X"FF",X"01",X"01",X"01",X"01",X"01",X"FF",X"00",
		X"CD",X"18",X"0B",X"3C",X"1B",X"00",X"01",X"0D",X"01",X"1E",X"FF",X"00",X"CD",X"18",X"0B",X"4D",
		X"1B",X"01",X"02",X"FF",X"32",X"01",X"FF",X"FF",X"32",X"01",X"01",X"00",X"00",X"CD",X"18",X"0B",
		X"5E",X"1B",X"01",X"02",X"FF",X"0A",X"01",X"FF",X"FF",X"0A",X"01",X"01",X"00",X"00",X"CD",X"18",
		X"0B",X"6D",X"1B",X"02",X"01",X"FF",X"0A",X"01",X"01",X"0A",X"01",X"FF",X"00",X"CD",X"17",X"0F",
		X"C9",X"CD",X"FF",X"08",X"01",X"01",X"FF",X"0A",X"0E",X"02",X"01",X"00",X"FA",X"2A",X"01",X"FF",
		X"C9",X"CD",X"FF",X"08",X"01",X"03",X"FF",X"0A",X"00",X"02",X"00",X"00",X"30",X"FF",X"C9",X"CD",
		X"C3",X"09",X"00",X"0A",X"0A",X"C9",X"CD",X"18",X"0B",X"AB",X"1B",X"00",X"01",X"08",X"0B",X"01",
		X"00",X"01",X"01",X"0F",X"0B",X"01",X"00",X"01",X"01",X"F1",X"00",X"C9",X"CD",X"FF",X"08",X"01",
		X"03",X"00",X"0A",X"0F",X"02",X"00",X"FF",X"C9",X"CD",X"C3",X"09",X"00",X"00",X"00",X"CD",X"C3",
		X"09",X"01",X"0A",X"0A",X"C9",X"CD",X"18",X"0B",X"D4",X"1B",X"01",X"01",X"00",X"01",X"0D",X"00",
		X"0F",X"0D",X"FF",X"00",X"CD",X"18",X"0B",X"E5",X"1B",X"00",X"02",X"FF",X"0A",X"01",X"03",X"00",
		X"0A",X"01",X"FD",X"FF",X"00",X"C9",X"CD",X"FF",X"08",X"01",X"00",X"FF",X"0A",X"00",X"00",X"52",
		X"02",X"01",X"FF",X"C9",X"CD",X"FA",X"09",X"00",X"00",X"CD",X"FA",X"09",X"01",X"0A",X"C9",X"CD",
		X"29",X"0C",X"5C",X"1C",X"00",X"02",X"00",X"28",X"00",X"00",X"28",X"00",X"00",X"28",X"00",X"00",
		X"28",X"00",X"00",X"14",X"52",X"01",X"1E",X"FD",X"00",X"0A",X"52",X"01",X"14",X"FD",X"00",X"3C",
		X"D5",X"00",X"3C",X"FD",X"00",X"1E",X"D5",X"00",X"0A",X"FD",X"00",X"14",X"D5",X"00",X"3C",X"A9",
		X"00",X"3C",X"D5",X"00",X"1E",X"A9",X"00",X"0A",X"D5",X"00",X"14",X"A9",X"00",X"3C",X"8E",X"00",
		X"3C",X"1C",X"01",X"1E",X"D5",X"00",X"0A",X"1C",X"01",X"14",X"D5",X"00",X"3C",X"A9",X"00",X"3C",
		X"A9",X"00",X"3C",X"A9",X"00",X"3C",X"A9",X"00",X"3C",X"A9",X"00",X"00",X"CD",X"29",X"0C",X"97",
		X"1C",X"01",X"01",X"FF",X"3C",X"00",X"3C",X"00",X"28",X"00",X"14",X"0A",X"3C",X"0A",X"3C",X"0A",
		X"3C",X"0A",X"3C",X"0A",X"3C",X"0A",X"3C",X"0A",X"3C",X"0A",X"3C",X"0A",X"3C",X"0A",X"3C",X"0A",
		X"3C",X"0A",X"3C",X"0A",X"14",X"0C",X"14",X"0B",X"14",X"0A",X"14",X"09",X"14",X"07",X"14",X"06",
		X"14",X"05",X"14",X"03",X"14",X"01",X"00",X"C9",X"CD",X"FF",X"08",X"01",X"00",X"FF",X"0A",X"0A",
		X"00",X"54",X"02",X"00",X"FF",X"C9",X"CD",X"FA",X"09",X"00",X"00",X"C9",X"CD",X"29",X"0C",X"FC",
		X"1D",X"00",X"02",X"00",X"08",X"54",X"00",X"08",X"6A",X"00",X"08",X"7F",X"00",X"08",X"A9",X"00",
		X"08",X"D5",X"00",X"14",X"FD",X"00",X"08",X"7F",X"00",X"08",X"A9",X"00",X"08",X"D5",X"00",X"08",
		X"FD",X"00",X"08",X"52",X"01",X"14",X"AA",X"01",X"08",X"A9",X"00",X"08",X"D5",X"00",X"08",X"FD",
		X"00",X"08",X"52",X"01",X"08",X"AA",X"01",X"14",X"FA",X"01",X"08",X"54",X"00",X"08",X"6A",X"00",
		X"08",X"7F",X"00",X"08",X"A9",X"00",X"08",X"D5",X"00",X"14",X"FD",X"00",X"08",X"7F",X"00",X"08",
		X"A9",X"00",X"08",X"D5",X"00",X"08",X"FD",X"00",X"08",X"52",X"01",X"14",X"AA",X"01",X"08",X"A9",
		X"00",X"08",X"D5",X"00",X"08",X"FD",X"00",X"08",X"52",X"01",X"08",X"AA",X"01",X"14",X"FA",X"01",
		X"08",X"54",X"00",X"08",X"6A",X"00",X"08",X"7F",X"00",X"08",X"A9",X"00",X"08",X"D5",X"00",X"14",
		X"FD",X"00",X"08",X"7F",X"00",X"08",X"A9",X"00",X"08",X"D5",X"00",X"08",X"FD",X"00",X"08",X"52",
		X"01",X"14",X"AA",X"01",X"08",X"A9",X"00",X"08",X"D5",X"00",X"08",X"FD",X"00",X"08",X"52",X"01",
		X"08",X"AA",X"01",X"14",X"FA",X"01",X"08",X"47",X"00",X"08",X"54",X"00",X"08",X"6A",X"00",X"08",
		X"8E",X"00",X"08",X"A9",X"00",X"14",X"D5",X"00",X"08",X"6A",X"00",X"08",X"8E",X"00",X"08",X"A9",
		X"00",X"08",X"D5",X"00",X"08",X"1C",X"01",X"14",X"52",X"01",X"07",X"8E",X"00",X"07",X"BE",X"00",
		X"07",X"E1",X"00",X"07",X"1C",X"01",X"06",X"7B",X"01",X"06",X"C3",X"01",X"14",X"38",X"02",X"08",
		X"47",X"00",X"08",X"54",X"00",X"08",X"6A",X"00",X"08",X"8E",X"00",X"08",X"A9",X"00",X"14",X"D5",
		X"00",X"08",X"6A",X"00",X"08",X"8E",X"00",X"08",X"A9",X"00",X"08",X"D5",X"00",X"08",X"1C",X"01",
		X"14",X"52",X"01",X"08",X"8E",X"00",X"08",X"A9",X"00",X"08",X"D5",X"00",X"08",X"1C",X"01",X"08",
		X"52",X"01",X"14",X"AA",X"01",X"08",X"47",X"00",X"08",X"54",X"00",X"08",X"6A",X"00",X"08",X"8E",
		X"00",X"08",X"A9",X"00",X"14",X"D5",X"00",X"08",X"6A",X"00",X"08",X"8E",X"00",X"08",X"A9",X"00",
		X"08",X"D5",X"00",X"08",X"1C",X"01",X"14",X"52",X"01",X"08",X"8E",X"00",X"08",X"A9",X"00",X"08",
		X"D5",X"00",X"08",X"1C",X"01",X"08",X"52",X"01",X"14",X"AA",X"01",X"00",X"C9",X"CD",X"FF",X"08",
		X"01",X"03",X"FF",X"0A",X"0B",X"00",X"A9",X"02",X"00",X"FF",X"C9",X"CD",X"FA",X"09",X"00",X"00",
		X"C9",X"CD",X"29",X"0C",X"F2",X"1E",X"00",X"01",X"00",X"0A",X"54",X"0A",X"50",X"0A",X"54",X"0A",
		X"50",X"0A",X"54",X"0A",X"50",X"0A",X"54",X"0A",X"50",X"0A",X"54",X"0A",X"50",X"0A",X"54",X"0A",
		X"50",X"0A",X"54",X"0A",X"50",X"0A",X"54",X"0A",X"50",X"0A",X"54",X"0A",X"50",X"0A",X"54",X"0A",
		X"50",X"0A",X"54",X"0A",X"50",X"0A",X"54",X"0A",X"50",X"0A",X"54",X"0A",X"50",X"0A",X"54",X"0A",
		X"50",X"0A",X"54",X"0A",X"50",X"0A",X"54",X"0A",X"50",X"0A",X"54",X"0A",X"50",X"0A",X"54",X"0A",
		X"50",X"0A",X"54",X"0A",X"50",X"0A",X"54",X"0A",X"50",X"0A",X"54",X"0A",X"50",X"0A",X"54",X"0A",
		X"50",X"0A",X"54",X"0A",X"50",X"0A",X"54",X"0A",X"50",X"0A",X"54",X"0A",X"50",X"0A",X"54",X"0A",
		X"50",X"0A",X"54",X"0A",X"50",X"0A",X"47",X"0A",X"3F",X"0A",X"47",X"0A",X"3F",X"0A",X"47",X"0A",
		X"3F",X"0A",X"47",X"0A",X"3F",X"0A",X"47",X"0A",X"3F",X"0A",X"47",X"0A",X"3F",X"0A",X"47",X"0A",
		X"3F",X"0A",X"47",X"0A",X"3F",X"0A",X"47",X"0A",X"3F",X"0A",X"47",X"0A",X"3F",X"0A",X"47",X"0A",
		X"3F",X"0A",X"47",X"0A",X"3F",X"0A",X"47",X"0A",X"3F",X"0A",X"47",X"0A",X"3F",X"0A",X"47",X"0A",
		X"3F",X"0A",X"47",X"0A",X"3F",X"0A",X"47",X"0A",X"3F",X"0A",X"47",X"0A",X"3F",X"0A",X"47",X"0A",
		X"3F",X"0A",X"47",X"0A",X"3F",X"0A",X"47",X"0A",X"3F",X"0A",X"47",X"0A",X"3F",X"0A",X"47",X"0A",
		X"3F",X"0A",X"47",X"0A",X"3F",X"0A",X"47",X"0A",X"3F",X"0A",X"47",X"0A",X"3F",X"0A",X"47",X"0A",
		X"3F",X"00",X"C9",X"CD",X"FF",X"08",X"01",X"02",X"FF",X"0A",X"09",X"00",X"FA",X"02",X"01",X"FF",
		X"C9",X"CD",X"FA",X"09",X"00",X"00",X"CD",X"FA",X"09",X"01",X"0A",X"C9",X"CD",X"29",X"0C",X"23",
		X"20",X"00",X"02",X"00",X"28",X"FA",X"01",X"05",X"FD",X"00",X"05",X"E1",X"00",X"05",X"D5",X"00",
		X"05",X"BE",X"00",X"28",X"A9",X"00",X"05",X"7F",X"00",X"05",X"71",X"00",X"05",X"6A",X"00",X"05",
		X"5F",X"00",X"28",X"54",X"00",X"05",X"52",X"01",X"05",X"7B",X"01",X"05",X"AA",X"01",X"05",X"C3",
		X"01",X"28",X"FA",X"01",X"05",X"FD",X"00",X"05",X"E1",X"00",X"05",X"D5",X"00",X"05",X"BE",X"00",
		X"28",X"A9",X"00",X"05",X"7F",X"00",X"05",X"71",X"00",X"05",X"6A",X"00",X"05",X"5F",X"00",X"28",
		X"54",X"00",X"05",X"52",X"01",X"05",X"7B",X"01",X"05",X"AA",X"01",X"05",X"C3",X"01",X"28",X"FA",
		X"01",X"05",X"FD",X"00",X"05",X"E1",X"00",X"05",X"D5",X"00",X"05",X"BE",X"00",X"28",X"A9",X"00",
		X"05",X"7F",X"00",X"05",X"71",X"00",X"05",X"6A",X"00",X"05",X"5F",X"00",X"28",X"54",X"00",X"05",
		X"AA",X"01",X"05",X"C3",X"01",X"05",X"DE",X"01",X"05",X"FA",X"01",X"28",X"38",X"02",X"05",X"D5",
		X"00",X"05",X"E1",X"00",X"05",X"EF",X"00",X"05",X"FD",X"00",X"28",X"1C",X"01",X"05",X"6A",X"00",
		X"05",X"71",X"00",X"05",X"77",X"00",X"05",X"7F",X"00",X"28",X"8E",X"00",X"05",X"1C",X"01",X"05",
		X"3F",X"01",X"05",X"52",X"01",X"05",X"7B",X"01",X"28",X"AA",X"01",X"05",X"D5",X"00",X"05",X"BE",
		X"00",X"05",X"A9",X"00",X"05",X"9F",X"00",X"28",X"8E",X"00",X"05",X"6A",X"00",X"05",X"5F",X"00",
		X"05",X"54",X"00",X"05",X"50",X"00",X"28",X"47",X"00",X"05",X"1C",X"01",X"05",X"3F",X"01",X"05",
		X"52",X"01",X"05",X"7B",X"01",X"28",X"AA",X"01",X"05",X"D5",X"00",X"05",X"BE",X"00",X"05",X"A9",
		X"00",X"05",X"9F",X"00",X"28",X"8E",X"00",X"05",X"6A",X"00",X"05",X"5F",X"00",X"05",X"54",X"00",
		X"05",X"50",X"00",X"28",X"47",X"00",X"05",X"1C",X"01",X"05",X"3F",X"01",X"05",X"52",X"01",X"05",
		X"7B",X"01",X"00",X"CD",X"29",X"0C",X"78",X"20",X"01",X"01",X"FF",X"14",X"0A",X"14",X"00",X"28",
		X"0A",X"14",X"00",X"28",X"0A",X"14",X"00",X"28",X"0A",X"14",X"00",X"28",X"0A",X"14",X"00",X"28",
		X"0A",X"14",X"00",X"28",X"0A",X"14",X"00",X"28",X"0A",X"14",X"00",X"28",X"0A",X"14",X"00",X"14",
		X"0A",X"28",X"0A",X"28",X"0A",X"14",X"00",X"28",X"0A",X"14",X"00",X"14",X"0A",X"14",X"0A",X"14",
		X"00",X"28",X"0A",X"14",X"00",X"28",X"0A",X"14",X"00",X"28",X"0A",X"14",X"00",X"28",X"0A",X"14",
		X"00",X"28",X"0A",X"14",X"00",X"14",X"0A",X"00",X"C9",X"CD",X"FF",X"08",X"01",X"06",X"FF",X"0A",
		X"00",X"00",X"F4",X"02",X"03",X"FF",X"C9",X"CD",X"FA",X"09",X"00",X"00",X"CD",X"FA",X"09",X"01",
		X"0A",X"C9",X"CD",X"29",X"0C",X"18",X"21",X"00",X"02",X"00",X"3C",X"F4",X"03",X"1E",X"F4",X"03",
		X"0A",X"FA",X"01",X"14",X"A4",X"02",X"1E",X"A4",X"02",X"0A",X"52",X"01",X"14",X"FA",X"01",X"3C",
		X"F4",X"03",X"1E",X"F4",X"03",X"0A",X"FA",X"01",X"14",X"A4",X"02",X"1E",X"A4",X"02",X"0A",X"52",
		X"01",X"14",X"FA",X"01",X"3C",X"F4",X"03",X"1E",X"F4",X"03",X"0A",X"FA",X"01",X"14",X"A4",X"02",
		X"1E",X"A4",X"02",X"0A",X"52",X"01",X"14",X"FA",X"01",X"3C",X"70",X"04",X"1E",X"70",X"04",X"0A",
		X"AA",X"01",X"14",X"38",X"02",X"1E",X"38",X"02",X"0A",X"1C",X"01",X"14",X"7B",X"01",X"3C",X"53",
		X"03",X"1E",X"53",X"03",X"0A",X"AA",X"01",X"14",X"38",X"02",X"1E",X"38",X"02",X"0A",X"1C",X"01",
		X"14",X"AA",X"01",X"3C",X"53",X"03",X"1E",X"53",X"03",X"0A",X"AA",X"01",X"14",X"38",X"02",X"1E",
		X"38",X"02",X"0A",X"1C",X"01",X"14",X"AA",X"01",X"CD",X"29",X"0C",X"35",X"21",X"01",X"01",X"FF",
		X"3C",X"00",X"28",X"0A",X"0A",X"0A",X"05",X"0A",X"05",X"00",X"28",X"0A",X"05",X"0B",X"05",X"09",
		X"05",X"07",X"05",X"04",X"00",X"C9",X"CD",X"29",X"0C",X"5C",X"1C",X"00",X"02",X"00",X"28",X"00",
		X"00",X"28",X"00",X"00",X"28",X"00",X"00",X"28",X"00",X"00",X"14",X"51",X"01",X"1E",X"FC",X"00",
		X"0A",X"51",X"01",X"14",X"FC",X"00",X"3C",X"D4",X"00",X"3C",X"FC",X"00",X"1E",X"D4",X"00",X"0A",
		X"FC",X"00",X"14",X"D4",X"00",X"3C",X"A8",X"00",X"3C",X"D4",X"00",X"1E",X"A8",X"00",X"0A",X"D4",
		X"00",X"14",X"A8",X"00",X"3C",X"8D",X"00",X"3C",X"1B",X"01",X"1E",X"D4",X"00",X"0A",X"1B",X"01",
		X"14",X"D4",X"00",X"3C",X"A8",X"00",X"3C",X"A8",X"00",X"3C",X"A8",X"00",X"3C",X"A8",X"00",X"3C",
		X"A8",X"00",X"00",X"CD",X"FF",X"08",X"01",X"05",X"FF",X"02",X"0C",X"18",X"01",X"16",X"08",X"0A",
		X"0C",X"FF",X"C9",X"CD",X"4B",X"0A",X"00",X"16",X"00",X"CD",X"4B",X"0A",X"01",X"18",X"02",X"CD",
		X"C3",X"09",X"01",X"0A",X"0A",X"CD",X"C3",X"09",X"00",X"00",X"02",X"C9",X"CD",X"AA",X"0E",X"C3",
		X"21",X"00",X"18",X"CD",X"18",X"0B",X"D4",X"21",X"00",X"02",X"02",X"04",X"01",X"02",X"00",X"04",
		X"01",X"FE",X"FF",X"00",X"CD",X"18",X"0B",X"E3",X"21",X"01",X"01",X"00",X"01",X"01",X"00",X"06",
		X"04",X"FF",X"00",X"C9",X"CD",X"FF",X"08",X"10",X"0B",X"FF",X"2A",X"0A",X"0A",X"0E",X"04",X"1F",
		X"FF",X"C9",X"CD",X"C3",X"09",X"00",X"0A",X"0A",X"CD",X"C3",X"09",X"01",X"2A",X"2A",X"C9",X"CD",
		X"18",X"0B",X"11",X"22",X"00",X"01",X"00",X"04",X"07",X"FF",X"01",X"01",X"05",X"0F",X"19",X"FF",
		X"00",X"CD",X"18",X"0B",X"23",X"22",X"01",X"01",X"00",X"03",X"09",X"00",X"01",X"01",X"FD",X"0F",
		X"19",X"00",X"00",X"CD",X"17",X"0F",X"C9",X"CD",X"FF",X"08",X"01",X"08",X"FF",X"0A",X"01",X"02",
		X"02",X"00",X"38",X"FF",X"C9",X"CD",X"C3",X"09",X"00",X"0A",X"0A",X"CD",X"C3",X"09",X"01",X"00",
		X"00",X"C9",X"CD",X"18",X"0B",X"51",X"22",X"00",X"01",X"05",X"01",X"01",X"0E",X"0E",X"01",X"FF",
		X"00",X"CD",X"18",X"0B",X"5E",X"22",X"01",X"02",X"FF",X"01",X"01",X"F6",X"FF",X"00",X"C9",X"CD",
		X"FF",X"08",X"01",X"08",X"FF",X"0A",X"0D",X"02",X"04",X"00",X"70",X"FF",X"C9",X"CD",X"C3",X"09",
		X"00",X"00",X"00",X"C9",X"CD",X"18",X"0B",X"85",X"22",X"00",X"02",X"FF",X"0A",X"02",X"01",X"00",
		X"0A",X"02",X"FF",X"FF",X"00",X"CD",X"18",X"0B",X"92",X"22",X"00",X"02",X"FF",X"19",X"01",X"FF",
		X"FF",X"00",X"C9",X"CD",X"FF",X"08",X"01",X"00",X"FF",X"00",X"FF",X"02",X"00",X"0A",X"0F",X"FF",
		X"C9",X"CD",X"C3",X"09",X"00",X"00",X"00",X"CD",X"C3",X"09",X"01",X"0A",X"0A",X"C9",X"CD",X"18",
		X"0B",X"BD",X"22",X"00",X"01",X"64",X"04",X"01",X"DD",X"04",X"01",X"18",X"00",X"CD",X"18",X"0B",
		X"C9",X"22",X"01",X"01",X"0D",X"01",X"3C",X"FF",X"00",X"C9",X"CD",X"FF",X"08",X"11",X"00",X"FF",
		X"00",X"00",X"02",X"00",X"0A",X"01",X"04",X"1F",X"2A",X"00",X"FF",X"C9",X"CD",X"C3",X"09",X"00",
		X"2A",X"2A",X"CD",X"C3",X"09",X"01",X"0A",X"0A",X"CD",X"C3",X"09",X"02",X"00",X"00",X"C9",X"CD",
		X"18",X"0B",X"FB",X"22",X"00",X"01",X"00",X"0F",X"07",X"01",X"00",X"CD",X"18",X"0B",X"10",X"23",
		X"01",X"01",X"00",X"01",X"01",X"0E",X"02",X"02",X"00",X"01",X"50",X"00",X"0D",X"01",X"FF",X"00",
		X"CD",X"18",X"0B",X"1D",X"23",X"02",X"02",X"00",X"43",X"01",X"28",X"00",X"00",X"CD",X"17",X"0F",
		X"C9",X"CD",X"FF",X"08",X"11",X"05",X"00",X"2A",X"00",X"04",X"1F",X"02",X"00",X"0A",X"0F",X"FF",
		X"C9",X"CD",X"C3",X"09",X"00",X"00",X"00",X"CD",X"C3",X"09",X"01",X"0A",X"0A",X"CD",X"C3",X"09",
		X"02",X"2A",X"2A",X"C9",X"CD",X"18",X"0B",X"65",X"23",X"01",X"01",X"00",X"06",X"01",X"FF",X"06",
		X"01",X"01",X"06",X"01",X"FF",X"06",X"01",X"01",X"06",X"01",X"FF",X"06",X"01",X"01",X"06",X"01",
		X"FF",X"06",X"01",X"01",X"00",X"CD",X"18",X"0B",X"71",X"23",X"01",X"01",X"00",X"06",X"08",X"FF",
		X"00",X"CD",X"18",X"0B",X"7D",X"23",X"02",X"01",X"00",X"0C",X"04",X"01",X"00",X"C9",X"CD",X"FF",
		X"08",X"01",X"03",X"FF",X"2E",X"05",X"32",X"05",X"16",X"ED",X"1A",X"ED",X"0A",X"0D",X"02",X"05",
		X"00",X"ED",X"FF",X"C9",X"CD",X"C3",X"09",X"00",X"16",X"00",X"CD",X"C3",X"09",X"01",X"1A",X"00",
		X"CD",X"C3",X"09",X"02",X"1A",X"1A",X"C9",X"CD",X"18",X"0B",X"B4",X"23",X"00",X"02",X"C8",X"01",
		X"19",X"00",X"00",X"00",X"CD",X"18",X"0B",X"C1",X"23",X"01",X"02",X"C8",X"01",X"32",X"00",X"00",
		X"00",X"CD",X"18",X"0B",X"CE",X"23",X"02",X"02",X"FF",X"01",X"01",X"FF",X"FF",X"00",X"C9",X"CD",
		X"FF",X"08",X"01",X"00",X"FF",X"0A",X"0F",X"02",X"00",X"00",X"26",X"FF",X"C9",X"CD",X"C3",X"09",
		X"00",X"00",X"00",X"C9",X"CD",X"18",X"0B",X"F3",X"23",X"00",X"01",X"09",X"01",X"01",X"0F",X"01",
		X"01",X"F1",X"00",X"C9",X"CD",X"FF",X"08",X"01",X"08",X"FF",X"0A",X"0F",X"02",X"03",X"00",X"26",
		X"FF",X"C9",X"CD",X"18",X"0B",X"13",X"24",X"00",X"02",X"04",X"07",X"01",X"0A",X"00",X"01",X"01",
		X"C9",X"FF",X"00",X"C9",X"CD",X"FF",X"08",X"01",X"00",X"00",X"0A",X"00",X"02",X"00",X"FF",X"C9",
		X"CD",X"C3",X"09",X"00",X"0A",X"0A",X"C9",X"CD",X"18",X"0B",X"39",X"24",X"00",X"01",X"00",X"01",
		X"01",X"0E",X"0A",X"01",X"00",X"0E",X"01",X"FF",X"00",X"C9",X"CD",X"FF",X"08",X"01",X"01",X"FF",
		X"0A",X"0F",X"02",X"01",X"00",X"1C",X"FF",X"C9",X"CD",X"C3",X"09",X"00",X"00",X"00",X"C9",X"CD",
		X"18",X"0B",X"60",X"24",X"00",X"02",X"19",X"06",X"01",X"F8",X"FF",X"06",X"01",X"08",X"00",X"00",
		X"C9",X"CD",X"FF",X"08",X"01",X"01",X"FF",X"0A",X"0F",X"02",X"00",X"00",X"ED",X"FF",X"C9",X"CD",
		X"18",X"0B",X"80",X"24",X"00",X"02",X"04",X"06",X"01",X"F8",X"FF",X"06",X"01",X"08",X"00",X"00",
		X"C9",X"CD",X"FF",X"08",X"01",X"01",X"FF",X"0A",X"0F",X"02",X"00",X"00",X"4C",X"FF",X"C9",X"CD",
		X"18",X"0B",X"A0",X"24",X"00",X"02",X"0C",X"06",X"02",X"F8",X"FF",X"06",X"02",X"08",X"00",X"00",
		X"C9",X"CD",X"FF",X"08",X"01",X"02",X"FF",X"0A",X"0F",X"00",X"F6",X"02",X"02",X"FF",X"C9",X"CD",
		X"C3",X"09",X"00",X"0A",X"0A",X"CD",X"C3",X"09",X"01",X"00",X"00",X"C9",X"CD",X"18",X"0B",X"C8",
		X"24",X"00",X"01",X"0F",X"01",X"13",X"FF",X"00",X"CD",X"18",X"0B",X"D9",X"24",X"01",X"02",X"FF",
		X"05",X"02",X"F6",X"FF",X"05",X"02",X"0A",X"00",X"00",X"C9",X"CD",X"FF",X"08",X"01",X"08",X"FF",
		X"0A",X"0F",X"00",X"FF",X"02",X"00",X"FF",X"C9",X"CD",X"C3",X"09",X"00",X"00",X"00",X"CD",X"C3",
		X"09",X"01",X"0A",X"0A",X"C9",X"CD",X"18",X"0B",X"12",X"25",X"00",X"02",X"04",X"0A",X"01",X"FF",
		X"FF",X"0A",X"01",X"01",X"00",X"00",X"CD",X"18",X"0B",X"12",X"25",X"01",X"01",X"00",X"0F",X"07",
		X"FF",X"00",X"C9",X"CD",X"FF",X"08",X"01",X"08",X"FF",X"0A",X"0F",X"00",X"FF",X"02",X"00",X"FF",
		X"C9",X"CD",X"C3",X"09",X"00",X"00",X"00",X"CD",X"C3",X"09",X"01",X"0A",X"0A",X"C9",X"CD",X"18",
		X"0B",X"4B",X"25",X"00",X"02",X"04",X"0A",X"01",X"01",X"00",X"0A",X"01",X"FF",X"FF",X"00",X"CD",
		X"18",X"0B",X"4B",X"25",X"01",X"01",X"00",X"0F",X"07",X"FF",X"00",X"C9",X"CD",X"FF",X"08",X"10",
		X"05",X"FF",X"2A",X"05",X"04",X"00",X"0A",X"0B",X"FF",X"C9",X"CD",X"C3",X"09",X"00",X"0A",X"0A",
		X"CD",X"C3",X"09",X"01",X"2A",X"2A",X"C9",X"CD",X"18",X"0B",X"76",X"25",X"00",X"01",X"00",X"04",
		X"03",X"01",X"08",X"01",X"FF",X"00",X"CD",X"18",X"0B",X"82",X"25",X"01",X"01",X"00",X"05",X"04",
		X"FF",X"00",X"CD",X"17",X"0F",X"C9",X"CD",X"FF",X"08",X"01",X"08",X"FF",X"0A",X"0F",X"00",X"80",
		X"02",X"00",X"FF",X"C9",X"CD",X"C3",X"09",X"00",X"00",X"00",X"C9",X"CD",X"18",X"0B",X"AC",X"25",
		X"00",X"02",X"FF",X"28",X"02",X"FE",X"FF",X"28",X"02",X"02",X"00",X"00",X"C9",X"CD",X"FF",X"08",
		X"01",X"01",X"02",X"0A",X"0A",X"00",X"00",X"FF",X"C9",X"CD",X"C3",X"09",X"00",X"00",X"00",X"CD",
		X"C3",X"09",X"01",X"0A",X"0A",X"C9",X"CD",X"18",X"0B",X"D3",X"25",X"00",X"02",X"00",X"70",X"01",
		X"10",X"00",X"00",X"CD",X"18",X"0B",X"E2",X"25",X"01",X"01",X"00",X"01",X"70",X"00",X"0A",X"01",
		X"FF",X"00",X"C9",X"CD",X"18",X"0B",X"D3",X"25",X"00",X"02",X"00",X"01",X"03",X"00",X"00",X"70",
		X"01",X"10",X"00",X"00",X"CD",X"FF",X"08",X"01",X"08",X"FF",X"16",X"00",X"0A",X"0F",X"00",X"C0",
		X"02",X"00",X"FF",X"C9",X"CD",X"C3",X"09",X"00",X"0A",X"0A",X"CD",X"C3",X"09",X"01",X"16",X"16",
		X"CD",X"9A",X"0A",X"00",X"16",X"0F",X"80",X"C9",X"CD",X"18",X"0B",X"27",X"26",X"00",X"01",X"0C",
		X"01",X"32",X"F1",X"01",X"32",X"0F",X"00",X"CD",X"18",X"0B",X"36",X"26",X"01",X"01",X"FF",X"01",
		X"64",X"0F",X"01",X"64",X"F1",X"00",X"CD",X"54",X"0F",X"00",X"C9",X"CD",X"FF",X"08",X"01",X"00",
		X"FF",X"0A",X"0C",X"00",X"FB",X"02",X"04",X"2C",X"10",X"FF",X"C9",X"CD",X"FA",X"09",X"00",X"00",
		X"00",X"CD",X"CD",X"0A",X"20",X"C9",X"CD",X"29",X"0C",X"1F",X"27",X"00",X"02",X"00",X"1C",X"FB",
		X"04",X"1C",X"53",X"03",X"1C",X"F4",X"03",X"1C",X"CC",X"02",X"1C",X"53",X"03",X"1C",X"7F",X"02",
		X"1C",X"CC",X"02",X"1C",X"FA",X"01",X"1C",X"7F",X"02",X"1C",X"AA",X"01",X"1C",X"FA",X"01",X"1C",
		X"66",X"01",X"1C",X"AA",X"01",X"1C",X"3F",X"01",X"1C",X"66",X"01",X"1C",X"FD",X"00",X"1C",X"3F",
		X"01",X"1C",X"D5",X"00",X"1C",X"FD",X"00",X"1C",X"B3",X"00",X"1C",X"D5",X"00",X"1C",X"9F",X"00",
		X"1C",X"B3",X"00",X"1C",X"7F",X"00",X"1C",X"9F",X"00",X"1C",X"6A",X"00",X"1C",X"7F",X"00",X"1C",
		X"59",X"00",X"1C",X"6A",X"00",X"1C",X"50",X"00",X"1C",X"59",X"00",X"1C",X"3F",X"00",X"1C",X"50",
		X"00",X"1C",X"3B",X"00",X"1C",X"3F",X"00",X"1C",X"47",X"00",X"1C",X"50",X"00",X"1C",X"59",X"00",
		X"1C",X"5F",X"00",X"1C",X"6A",X"00",X"1C",X"77",X"00",X"1C",X"3B",X"00",X"1C",X"3F",X"00",X"1C",
		X"47",X"00",X"1C",X"50",X"00",X"1C",X"59",X"00",X"1C",X"5F",X"00",X"1C",X"6A",X"00",X"1C",X"77",
		X"00",X"1C",X"EF",X"00",X"1C",X"D5",X"00",X"1C",X"BE",X"00",X"1C",X"B3",X"00",X"1C",X"9F",X"00",
		X"1C",X"8E",X"00",X"1C",X"7F",X"00",X"1C",X"77",X"00",X"1C",X"6A",X"00",X"1C",X"5F",X"00",X"1C",
		X"59",X"00",X"1C",X"50",X"00",X"1C",X"47",X"00",X"1C",X"3F",X"00",X"1C",X"3B",X"00",X"00",X"CD",
		X"8A",X"0E",X"C9",X"CD",X"FF",X"08",X"10",X"00",X"FF",X"0A",X"09",X"04",X"1F",X"FF",X"C9",X"CD",
		X"C3",X"09",X"00",X"0A",X"0A",X"C9",X"CD",X"18",X"0B",X"48",X"27",X"00",X"01",X"00",X"02",X"01",
		X"03",X"05",X"01",X"00",X"0F",X"03",X"FF",X"00",X"C9",X"CD",X"FF",X"08",X"CD",X"C3",X"09",X"CD",
		X"18",X"0B",X"CD",X"18",X"0B",X"C9",X"CD",X"FF",X"08",X"CD",X"C3",X"09",X"CD",X"18",X"0B",X"CD",
		X"18",X"0B",X"C9",X"CD",X"FF",X"08",X"01",X"08",X"FF",X"0A",X"00",X"00",X"FF",X"02",X"00",X"FF",
		X"C9",X"CD",X"C3",X"09",X"00",X"0A",X"0A",X"CD",X"C3",X"09",X"01",X"00",X"00",X"C9",X"CD",X"18",
		X"0B",X"90",X"27",X"00",X"01",X"00",X"0E",X"03",X"01",X"01",X"02",X"01",X"01",X"01",X"F1",X"00",
		X"CD",X"18",X"0B",X"A1",X"27",X"01",X"02",X"09",X"03",X"01",X"FA",X"FF",X"02",X"01",X"05",X"00",
		X"00",X"C9",X"CD",X"FF",X"08",X"01",X"08",X"FF",X"0A",X"0F",X"00",X"80",X"02",X"01",X"FF",X"C9",
		X"CD",X"C3",X"09",X"00",X"00",X"00",X"C9",X"CD",X"18",X"0B",X"C8",X"27",X"00",X"02",X"0A",X"1E",
		X"01",X"FF",X"FF",X"01",X"01",X"0F",X"00",X"00",X"C9",X"CD",X"FF",X"08",X"01",X"08",X"FF",X"0A",
		X"0F",X"02",X"04",X"00",X"80",X"FF",X"C9",X"CD",X"C3",X"09",X"00",X"0A",X"0A",X"C9",X"CD",X"18",
		X"0B",X"08",X"28",X"00",X"01",X"00",X"0F",X"02",X"FF",X"01",X"01",X"0E",X"0E",X"02",X"FF",X"01",
		X"01",X"0D",X"0D",X"01",X"FF",X"01",X"01",X"0C",X"0C",X"01",X"FF",X"01",X"01",X"0B",X"0B",X"01",
		X"FF",X"01",X"01",X"0A",X"0A",X"01",X"FF",X"00",X"C9",X"CD",X"FF",X"08",X"10",X"08",X"FF",X"0A",
		X"00",X"04",X"1F",X"FF",X"C9",X"CD",X"C3",X"09",X"00",X"0A",X"0A",X"C9",X"CD",X"18",X"0B",X"49",
		X"28",X"00",X"01",X"00",X"01",X"01",X"0F",X"0F",X"02",X"FF",X"01",X"01",X"0E",X"0E",X"02",X"FF",
		X"01",X"01",X"0D",X"0D",X"01",X"FF",X"01",X"01",X"0C",X"0C",X"01",X"FF",X"01",X"01",X"0B",X"0B",
		X"01",X"FF",X"01",X"01",X"0A",X"0A",X"01",X"FF",X"00",X"C9",X"CD",X"FF",X"08",X"CD",X"FF",X"08",
		X"01",X"00",X"00",X"16",X"00",X"2A",X"00",X"0A",X"0D",X"02",X"00",X"FF",X"C9",X"CD",X"C3",X"09",
		X"00",X"0A",X"0A",X"CD",X"C3",X"09",X"01",X"00",X"00",X"CD",X"C3",X"09",X"02",X"2A",X"2A",X"CD",
		X"9A",X"0A",X"00",X"16",X"0F",X"80",X"C9",X"CD",X"18",X"0B",X"86",X"28",X"00",X"01",X"00",X"02",
		X"0A",X"FF",X"01",X"01",X"00",X"00",X"CD",X"18",X"0B",X"93",X"28",X"01",X"02",X"00",X"15",X"01",
		X"07",X"00",X"00",X"CD",X"18",X"0B",X"A2",X"28",X"02",X"01",X"03",X"05",X"01",X"01",X"02",X"01",
		X"00",X"00",X"CD",X"18",X"0B",X"B4",X"28",X"03",X"01",X"00",X"03",X"01",X"00",X"01",X"0F",X"01",
		X"03",X"01",X"00",X"00",X"CD",X"17",X"0F",X"CD",X"54",X"0F",X"00",X"C9",X"CD",X"FF",X"08",X"11",
		X"08",X"FF",X"04",X"1F",X"0A",X"01",X"02",X"70",X"00",X"04",X"FF",X"C9",X"CD",X"C3",X"09",X"00",
		X"0A",X"0A",X"CD",X"C3",X"09",X"01",X"00",X"00",X"CD",X"C3",X"09",X"02",X"2A",X"2A",X"C9",X"CD",
		X"18",X"0B",X"F1",X"28",X"00",X"01",X"FF",X"0E",X"18",X"01",X"0E",X"0C",X"00",X"0E",X"0C",X"FF",
		X"00",X"CD",X"18",X"0B",X"02",X"29",X"01",X"02",X"FF",X"A8",X"02",X"FF",X"FF",X"A8",X"02",X"01",
		X"00",X"00",X"CD",X"18",X"0B",X"11",X"29",X"02",X"01",X"FF",X"08",X"2A",X"01",X"08",X"2A",X"FF",
		X"00",X"CD",X"17",X"0F",X"C9",X"CD",X"FF",X"08",X"10",X"00",X"FF",X"04",X"0A",X"2A",X"00",X"0A",
		X"0A",X"FF",X"C9",X"CD",X"C3",X"09",X"00",X"0A",X"0A",X"CD",X"C3",X"09",X"01",X"2A",X"2A",X"CD",
		X"C3",X"09",X"02",X"04",X"04",X"C9",X"CD",X"18",X"0B",X"45",X"29",X"00",X"01",X"00",X"02",X"0A",
		X"FF",X"01",X"01",X"00",X"00",X"CD",X"18",X"0B",X"54",X"29",X"01",X"01",X"03",X"05",X"01",X"01",
		X"02",X"01",X"00",X"00",X"CD",X"18",X"0B",X"60",X"29",X"02",X"01",X"00",X"14",X"01",X"01",X"00",
		X"CD",X"17",X"0F",X"C9",X"CD",X"FF",X"08",X"01",X"00",X"00",X"2A",X"00",X"0A",X"0D",X"02",X"01",
		X"FF",X"C9",X"CD",X"FF",X"08",X"01",X"00",X"00",X"2A",X"00",X"0A",X"0D",X"02",X"02",X"FF",X"C9",
		X"CD",X"FF",X"08",X"01",X"02",X"FF",X"0A",X"01",X"00",X"DE",X"02",X"01",X"FF",X"C9",X"CD",X"C3",
		X"09",X"00",X"0A",X"0A",X"C9",X"CD",X"18",X"0B",X"A7",X"29",X"00",X"01",X"00",X"04",X"01",X"03",
		X"01",X"34",X"00",X"04",X"01",X"FD",X"00",X"C9",X"CD",X"FF",X"08",X"01",X"02",X"FF",X"0A",X"01",
		X"00",X"AA",X"02",X"01",X"FF",X"C9",X"CD",X"18",X"0B",X"A7",X"29",X"00",X"01",X"00",X"01",X"3C",
		X"00",X"04",X"01",X"03",X"01",X"34",X"00",X"04",X"01",X"FD",X"00",X"CD",X"FF",X"08",X"01",X"02",
		X"FF",X"0A",X"01",X"00",X"7B",X"02",X"01",X"FF",X"C9",X"CD",X"18",X"0B",X"A7",X"29",X"00",X"01",
		X"00",X"01",X"78",X"00",X"04",X"01",X"03",X"01",X"34",X"00",X"04",X"01",X"FD",X"00",X"CD",X"FF",
		X"08",X"01",X"02",X"FF",X"0A",X"01",X"00",X"52",X"02",X"01",X"FF",X"C9",X"CD",X"18",X"0B",X"A7",
		X"29",X"00",X"01",X"00",X"01",X"B4",X"00",X"04",X"01",X"03",X"01",X"34",X"00",X"04",X"01",X"FD",
		X"00",X"CD",X"FF",X"08",X"01",X"02",X"FF",X"0A",X"01",X"00",X"2D",X"02",X"01",X"FF",X"C9",X"CD",
		X"18",X"0B",X"A7",X"29",X"00",X"01",X"00",X"01",X"F0",X"00",X"04",X"01",X"03",X"01",X"34",X"00",
		X"04",X"01",X"FD",X"00",X"CD",X"FF",X"08",X"01",X"02",X"FF",X"0A",X"01",X"00",X"0C",X"02",X"01",
		X"FF",X"C9",X"CD",X"18",X"0B",X"A7",X"29",X"00",X"01",X"00",X"01",X"C8",X"00",X"01",X"64",X"00",
		X"04",X"01",X"03",X"01",X"34",X"00",X"04",X"01",X"FD",X"00",X"CD",X"FF",X"08",X"01",X"01",X"FF",
		X"0A",X"00",X"FF",X"C9",X"CD",X"22",X"0A",X"00",X"C9",X"CD",X"05",X"0D",X"A7",X"29",X"00",X"00",
		X"95",X"2A",X"00",X"00",X"CD",X"05",X"0D",X"A7",X"29",X"00",X"00",X"B7",X"2A",X"00",X"00",X"CD",
		X"05",X"0D",X"A7",X"29",X"00",X"00",X"D9",X"2A",X"00",X"00",X"CD",X"05",X"0D",X"A7",X"29",X"00",
		X"00",X"FB",X"2A",X"00",X"00",X"0D",X"EF",X"00",X"0F",X"00",X"00",X"0D",X"EF",X"00",X"0D",X"EF",
		X"00",X"0B",X"BE",X"00",X"0B",X"EF",X"00",X"0B",X"BE",X"00",X"0B",X"9F",X"00",X"0B",X"BE",X"00",
		X"0B",X"9F",X"00",X"09",X"77",X"00",X"00",X"0D",X"3F",X"01",X"0F",X"00",X"00",X"0D",X"3F",X"01",
		X"0D",X"3F",X"01",X"0B",X"EF",X"00",X"0B",X"3F",X"01",X"0B",X"EF",X"00",X"0B",X"3F",X"01",X"0B",
		X"EF",X"00",X"0B",X"EF",X"00",X"09",X"BE",X"00",X"00",X"0D",X"F6",X"02",X"0F",X"00",X"00",X"0D",
		X"F6",X"02",X"0D",X"F6",X"02",X"0B",X"7F",X"02",X"0B",X"F6",X"02",X"0B",X"7F",X"02",X"0B",X"7F",
		X"02",X"0B",X"7F",X"02",X"0B",X"DE",X"01",X"09",X"DE",X"01",X"00",X"0D",X"BC",X"03",X"0F",X"00",
		X"00",X"0D",X"BC",X"03",X"0D",X"BC",X"03",X"0B",X"F6",X"02",X"0B",X"BC",X"03",X"0B",X"F6",X"02",
		X"0B",X"7F",X"02",X"0B",X"F6",X"02",X"0B",X"7F",X"02",X"09",X"7F",X"02",X"00",X"05",X"02",X"01",
		X"03",X"02",X"04",X"FF",X"01",X"25",X"FE",X"01",X"01",X"FE",X"00",X"05",X"02",X"01",X"03",X"02",
		X"06",X"FF",X"02",X"01",X"FF",X"00",X"05",X"02",X"01",X"03",X"01",X"04",X"FF",X"01",X"05",X"FE",
		X"01",X"01",X"FE",X"00",X"00",X"01",X"0C",X"00",X"00",X"00",X"CD",X"FF",X"08",X"01",X"01",X"FF",
		X"0A",X"00",X"FF",X"C9",X"CD",X"22",X"0A",X"00",X"C9",X"CD",X"05",X"0D",X"A7",X"29",X"00",X"05",
		X"6F",X"2B",X"00",X"00",X"CD",X"05",X"0D",X"A7",X"29",X"00",X"00",X"88",X"2B",X"00",X"00",X"0D",
		X"2F",X"0B",X"0D",X"2F",X"0B",X"0D",X"F7",X"09",X"0D",X"2F",X"0B",X"0D",X"68",X"09",X"0D",X"2F",
		X"0B",X"0D",X"E1",X"08",X"0D",X"2F",X"0B",X"00",X"09",X"68",X"09",X"00",X"68",X"09",X"0D",X"68",
		X"09",X"0D",X"2F",X"0B",X"09",X"2F",X"0B",X"09",X"68",X"09",X"09",X"61",X"08",X"09",X"E9",X"07",
		X"09",X"E9",X"07",X"09",X"E9",X"07",X"09",X"E9",X"07",X"09",X"61",X"08",X"09",X"68",X"09",X"09",
		X"2F",X"0B",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
