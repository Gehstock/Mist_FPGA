library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity bg_graphx_3 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of bg_graphx_3 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"F0",X"C0",X"00",X"70",X"7C",X"7E",X"7E",X"7C",X"70",X"00",X"C0",X"F0",X"C0",X"00",
		X"E3",X"CF",X"03",X"6F",X"03",X"00",X"00",X"3B",X"3B",X"00",X"00",X"03",X"6F",X"03",X"CF",X"E3",
		X"FF",X"FC",X"FE",X"FC",X"F8",X"F8",X"F0",X"00",X"08",X"E8",X"C4",X"C4",X"C2",X"C2",X"81",X"01",
		X"80",X"81",X"43",X"41",X"23",X"23",X"17",X"10",X"00",X"0F",X"1F",X"1F",X"1F",X"7F",X"FF",X"FF",
		X"01",X"C1",X"C2",X"82",X"C4",X"C4",X"E8",X"08",X"00",X"F0",X"F8",X"F8",X"F8",X"FC",X"FC",X"FF",
		X"FF",X"FF",X"7F",X"1F",X"1F",X"1F",X"0F",X"00",X"10",X"17",X"23",X"23",X"41",X"43",X"80",X"80",
		X"FF",X"FE",X"FE",X"FC",X"F8",X"F0",X"F0",X"F8",X"F8",X"F0",X"C0",X"C0",X"80",X"80",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"01",X"01",X"01",X"01",X"01",X"03",X"03",X"03",X"03",X"03",X"07",X"1F",X"0F",X"3F",X"7F",X"7F",
		X"01",X"01",X"02",X"02",X"04",X"04",X"08",X"08",X"10",X"10",X"20",X"20",X"40",X"40",X"80",X"80",
		X"00",X"00",X"80",X"80",X"80",X"00",X"00",X"C0",X"E0",X"E0",X"F0",X"F0",X"F8",X"FC",X"FE",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"7F",X"7F",X"3F",X"3F",X"1F",X"3F",X"1F",X"0F",X"0F",X"07",X"07",X"07",X"01",X"01",X"01",
		X"80",X"80",X"40",X"40",X"20",X"20",X"10",X"10",X"08",X"08",X"04",X"04",X"02",X"02",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"40",X"40",X"20",X"10",X"10",X"08",X"04",X"02",X"04",X"04",X"02",X"02",X"02",X"01",
		X"80",X"80",X"40",X"20",X"18",X"04",X"08",X"08",X"04",X"04",X"02",X"04",X"02",X"02",X"01",X"01",
		X"80",X"80",X"40",X"40",X"20",X"20",X"10",X"10",X"08",X"08",X"04",X"04",X"02",X"02",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"02",X"01",X"02",X"04",X"04",X"02",X"04",X"08",X"08",X"10",X"20",X"40",X"40",X"80",X"80",
		X"01",X"01",X"02",X"02",X"04",X"04",X"06",X"08",X"10",X"20",X"10",X"20",X"20",X"40",X"80",X"80",
		X"01",X"01",X"02",X"02",X"04",X"04",X"08",X"08",X"10",X"10",X"20",X"20",X"40",X"40",X"80",X"80",
		X"FF",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FC",X"FC",X"F8",X"F8",X"F0",X"C0",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"81",X"81",X"43",X"43",X"27",X"27",X"1F",X"1F",X"1F",X"1F",X"3F",X"3F",X"7F",X"7F",X"FF",X"FF",
		X"01",X"01",X"02",X"02",X"04",X"04",X"08",X"08",X"10",X"10",X"20",X"20",X"40",X"40",X"80",X"80",
		X"00",X"C0",X"F0",X"F8",X"F8",X"FC",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"7F",X"7F",X"3F",X"3F",X"1F",X"1F",X"1F",X"1F",X"27",X"27",X"43",X"43",X"81",X"81",
		X"80",X"80",X"40",X"40",X"20",X"20",X"10",X"10",X"08",X"08",X"04",X"04",X"02",X"02",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"04",X"06",X"0C",X"03",X"02",X"03",X"02",X"0E",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"09",X"05",X"07",X"0D",X"02",X"03",X"02",X"0E",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0C",X"03",X"02",X"03",X"02",X"0E",X"04",X"0E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"02",X"06",X"04",X"03",X"0F",X"05",X"0F",X"0B",X"0A",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0C",X"03",X"07",X"05",X"02",X"03",X"02",X"03",X"02",X"0E",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"0E",X"04",X"03",X"02",X"06",X"0C",X"03",X"0A",X"00",X"00",X"00",
		X"00",X"00",X"08",X"09",X"05",X"0F",X"05",X"02",X"03",X"07",X"0D",X"02",X"03",X"0A",X"00",X"00",
		X"00",X"00",X"0C",X"03",X"02",X"03",X"02",X"03",X"02",X"0E",X"04",X"03",X"02",X"0E",X"00",X"00",
		X"00",X"00",X"00",X"0C",X"03",X"02",X"03",X"02",X"03",X"0F",X"05",X"02",X"0E",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"0E",X"0C",X"06",X"04",X"03",X"02",X"0E",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"09",X"0D",X"07",X"05",X"02",X"0E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"03",X"02",X"0E",X"04",X"03",X"0F",X"0B",X"0A",X"00",X"00",X"00",
		X"00",X"00",X"08",X"09",X"0D",X"02",X"03",X"0F",X"05",X"02",X"03",X"02",X"0E",X"00",X"00",X"00",
		X"00",X"00",X"0C",X"03",X"02",X"03",X"02",X"03",X"02",X"03",X"02",X"0E",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0C",X"03",X"02",X"06",X"04",X"0E",X"04",X"03",X"0F",X"0B",X"0A",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"03",X"07",X"05",X"0F",X"05",X"02",X"03",X"02",X"0E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"02",X"03",X"02",X"03",X"02",X"03",X"02",X"0E",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"02",X"06",X"0C",X"03",X"02",X"03",X"02",X"0E",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0C",X"03",X"07",X"0D",X"02",X"03",X"02",X"03",X"0A",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"02",X"03",X"02",X"06",X"0C",X"03",X"02",X"0E",X"00",X"00",X"00",X"00",
		X"00",X"00",X"08",X"02",X"06",X"0C",X"03",X"07",X"0D",X"02",X"03",X"0F",X"0B",X"0A",X"00",X"00",
		X"00",X"00",X"0C",X"03",X"07",X"0D",X"02",X"06",X"04",X"03",X"02",X"03",X"02",X"03",X"0A",X"00",
		X"00",X"00",X"00",X"04",X"03",X"02",X"03",X"07",X"05",X"02",X"0E",X"04",X"03",X"02",X"0E",X"00",
		X"00",X"08",X"09",X"05",X"02",X"03",X"02",X"03",X"02",X"03",X"0F",X"05",X"02",X"03",X"0A",X"00",
		X"00",X"0C",X"03",X"02",X"06",X"0C",X"06",X"04",X"03",X"02",X"0E",X"04",X"03",X"02",X"0E",X"00",
		X"00",X"00",X"0C",X"03",X"07",X"0D",X"07",X"05",X"02",X"03",X"0F",X"05",X"02",X"03",X"0A",X"00",
		X"08",X"09",X"0D",X"02",X"03",X"02",X"03",X"02",X"03",X"02",X"03",X"02",X"03",X"02",X"06",X"00",
		X"02",X"03",X"02",X"06",X"0C",X"03",X"02",X"06",X"04",X"03",X"02",X"0E",X"04",X"03",X"07",X"0B",
		X"03",X"02",X"03",X"07",X"0D",X"02",X"03",X"07",X"05",X"02",X"03",X"0F",X"05",X"02",X"06",X"04",
		X"02",X"03",X"02",X"06",X"04",X"03",X"02",X"06",X"04",X"03",X"02",X"06",X"04",X"03",X"07",X"05",
		X"03",X"02",X"03",X"07",X"05",X"02",X"03",X"07",X"05",X"02",X"03",X"07",X"05",X"02",X"03",X"02",
		X"02",X"03",X"02",X"03",X"02",X"03",X"02",X"03",X"02",X"03",X"02",X"03",X"02",X"03",X"02",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"0A",X"00",X"0C",X"03",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"03",X"09",X"0D",X"02",X"0E",X"00",X"08",X"0A",X"00",X"00",X"00",
		X"00",X"00",X"08",X"09",X"0D",X"02",X"03",X"02",X"0E",X"00",X"00",X"0C",X"03",X"0A",X"00",X"00",
		X"00",X"08",X"02",X"03",X"02",X"0E",X"0C",X"0E",X"00",X"08",X"09",X"0D",X"02",X"03",X"0A",X"00",
		X"00",X"0C",X"03",X"02",X"03",X"0F",X"0B",X"0A",X"08",X"02",X"06",X"04",X"03",X"02",X"0E",X"00",
		X"00",X"08",X"02",X"06",X"0C",X"03",X"02",X"06",X"0C",X"03",X"07",X"05",X"02",X"03",X"0A",X"00",
		X"00",X"0C",X"03",X"07",X"0D",X"02",X"03",X"07",X"0D",X"02",X"0E",X"0C",X"03",X"02",X"0E",X"00",
		X"00",X"00",X"0C",X"0E",X"0C",X"03",X"02",X"0E",X"0C",X"0E",X"00",X"00",X"0C",X"03",X"0A",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"0E",X"00",X"08",X"0A",X"08",X"09",X"0D",X"02",X"0E",X"00",
		X"00",X"00",X"00",X"08",X"0A",X"08",X"0A",X"08",X"02",X"0E",X"04",X"03",X"02",X"0E",X"00",X"00",
		X"00",X"00",X"00",X"0C",X"06",X"04",X"03",X"02",X"03",X"0F",X"05",X"02",X"0E",X"00",X"00",X"00",
		X"00",X"08",X"09",X"0D",X"07",X"05",X"02",X"0E",X"0C",X"0E",X"0C",X"0E",X"00",X"00",X"00",X"00",
		X"00",X"0C",X"03",X"02",X"06",X"0C",X"06",X"00",X"00",X"00",X"08",X"0A",X"08",X"0A",X"00",X"00",
		X"00",X"00",X"0C",X"03",X"07",X"0D",X"07",X"0B",X"09",X"0B",X"02",X"03",X"02",X"03",X"0A",X"00",
		X"00",X"00",X"08",X"02",X"03",X"02",X"03",X"02",X"0E",X"0C",X"03",X"02",X"03",X"02",X"0E",X"00",
		X"00",X"00",X"0C",X"03",X"02",X"03",X"02",X"0E",X"00",X"00",X"0C",X"06",X"0C",X"03",X"0A",X"00",
		X"00",X"00",X"00",X"0C",X"0E",X"0C",X"0E",X"00",X"08",X"09",X"0D",X"07",X"0D",X"02",X"0E",X"00",
		X"00",X"00",X"00",X"08",X"0A",X"08",X"0A",X"08",X"02",X"03",X"02",X"03",X"02",X"0E",X"00",X"00",
		X"00",X"00",X"08",X"02",X"06",X"0C",X"03",X"02",X"03",X"02",X"0E",X"0C",X"0E",X"00",X"00",X"00",
		X"00",X"00",X"0C",X"03",X"07",X"0D",X"02",X"03",X"02",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"08",X"02",X"06",X"0C",X"06",X"0C",X"0E",X"00",X"08",X"0A",X"00",X"00",X"00",X"00",
		X"00",X"08",X"02",X"03",X"07",X"0D",X"07",X"0B",X"0A",X"08",X"02",X"0E",X"00",X"00",X"00",X"00",
		X"00",X"0C",X"03",X"02",X"0E",X"04",X"0E",X"04",X"03",X"02",X"03",X"0F",X"0B",X"0A",X"00",X"00",
		X"00",X"00",X"0C",X"03",X"0F",X"05",X"0F",X"05",X"02",X"0E",X"0C",X"03",X"02",X"03",X"0A",X"00",
		X"00",X"00",X"00",X"0C",X"0E",X"0C",X"0E",X"0C",X"0E",X"00",X"00",X"0C",X"03",X"02",X"0E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"0A",X"08",X"09",X"0D",X"02",X"0E",X"00",X"00",
		X"00",X"00",X"08",X"09",X"0B",X"0A",X"08",X"02",X"03",X"02",X"03",X"02",X"0E",X"00",X"00",X"00",
		X"00",X"08",X"02",X"06",X"0C",X"03",X"02",X"03",X"02",X"06",X"04",X"0E",X"00",X"00",X"00",X"00",
		X"00",X"0C",X"03",X"07",X"0D",X"02",X"03",X"02",X"03",X"07",X"05",X"0F",X"0B",X"0A",X"00",X"00",
		X"00",X"08",X"02",X"03",X"02",X"0E",X"0C",X"06",X"0C",X"0E",X"0C",X"03",X"02",X"0E",X"00",X"00",
		X"00",X"0C",X"03",X"02",X"03",X"0F",X"0D",X"07",X"0B",X"0A",X"00",X"0C",X"0E",X"00",X"00",X"00",
		X"00",X"00",X"0C",X"03",X"02",X"0E",X"04",X"03",X"02",X"03",X"0A",X"08",X"0A",X"00",X"00",X"00",
		X"08",X"09",X"0D",X"02",X"03",X"0F",X"05",X"02",X"0E",X"04",X"03",X"02",X"03",X"0A",X"08",X"0A",
		X"02",X"03",X"02",X"03",X"02",X"06",X"04",X"03",X"0F",X"05",X"02",X"06",X"04",X"03",X"02",X"03",
		X"03",X"02",X"03",X"02",X"03",X"07",X"05",X"02",X"03",X"02",X"03",X"07",X"05",X"02",X"03",X"02",
		X"04",X"03",X"02",X"03",X"02",X"06",X"04",X"03",X"02",X"03",X"02",X"03",X"02",X"03",X"02",X"03");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
