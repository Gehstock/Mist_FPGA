library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity travusa_sound is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of travusa_sound is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"76",X"BB",X"5A",X"0F",X"55",X"00",X"54",X"5B",X"14",X"30",X"04",X"14",X"33",X"04",X"14",X"36",
		X"04",X"14",X"39",X"04",X"14",X"3D",X"04",X"14",X"40",X"04",X"14",X"44",X"04",X"14",X"48",X"04",
		X"14",X"4D",X"04",X"14",X"50",X"04",X"14",X"56",X"04",X"14",X"5B",X"04",X"14",X"60",X"04",X"14",
		X"66",X"04",X"14",X"6C",X"04",X"14",X"73",X"04",X"14",X"7A",X"04",X"14",X"81",X"04",X"14",X"88",
		X"04",X"14",X"90",X"04",X"14",X"99",X"04",X"14",X"A1",X"04",X"14",X"AB",X"04",X"14",X"B6",X"04",
		X"5A",X"00",X"77",X"04",X"FF",X"04",X"14",X"0E",X"04",X"14",X"0F",X"04",X"14",X"10",X"04",X"14",
		X"11",X"04",X"14",X"12",X"04",X"14",X"13",X"04",X"14",X"14",X"04",X"14",X"15",X"04",X"14",X"16",
		X"04",X"14",X"17",X"04",X"14",X"18",X"04",X"14",X"19",X"04",X"14",X"1A",X"04",X"14",X"1B",X"04",
		X"14",X"1C",X"04",X"14",X"1E",X"04",X"14",X"20",X"04",X"14",X"22",X"04",X"14",X"24",X"04",X"14",
		X"26",X"04",X"14",X"28",X"04",X"14",X"2A",X"04",X"5A",X"00",X"77",X"04",X"FF",X"76",X"BB",X"5A",
		X"0F",X"55",X"00",X"54",X"48",X"14",X"45",X"04",X"14",X"4F",X"04",X"14",X"4D",X"04",X"14",X"4E",
		X"04",X"14",X"45",X"04",X"14",X"43",X"04",X"14",X"4B",X"04",X"14",X"48",X"04",X"14",X"49",X"04",
		X"14",X"4A",X"04",X"14",X"43",X"04",X"14",X"4F",X"04",X"14",X"4C",X"04",X"14",X"45",X"04",X"14",
		X"40",X"04",X"14",X"49",X"04",X"14",X"48",X"04",X"14",X"4F",X"04",X"14",X"4D",X"04",X"14",X"4F",
		X"04",X"14",X"4B",X"04",X"14",X"48",X"04",X"14",X"47",X"04",X"14",X"4A",X"04",X"14",X"44",X"04",
		X"14",X"4D",X"04",X"14",X"45",X"04",X"14",X"41",X"04",X"14",X"4A",X"04",X"14",X"4C",X"04",X"14",
		X"48",X"04",X"14",X"45",X"04",X"14",X"4D",X"04",X"14",X"4A",X"04",X"14",X"45",X"04",X"14",X"46",
		X"04",X"14",X"47",X"04",X"14",X"4F",X"04",X"14",X"48",X"04",X"14",X"40",X"04",X"14",X"4C",X"04",
		X"14",X"4D",X"04",X"14",X"49",X"04",X"14",X"43",X"04",X"14",X"42",X"04",X"14",X"49",X"04",X"14",
		X"4A",X"04",X"14",X"4E",X"04",X"14",X"4A",X"04",X"14",X"4B",X"04",X"14",X"48",X"04",X"5A",X"00",
		X"77",X"04",X"FF",X"76",X"BD",X"59",X"10",X"5B",X"00",X"5C",X"01",X"5D",X"0D",X"53",X"00",X"FE",
		X"E1",X"5F",X"FE",X"E1",X"5F",X"FE",X"E1",X"58",X"59",X"00",X"5C",X"00",X"77",X"02",X"FF",X"12",
		X"64",X"04",X"12",X"63",X"04",X"12",X"62",X"04",X"12",X"61",X"04",X"12",X"60",X"12",X"12",X"48",
		X"04",X"12",X"47",X"04",X"12",X"46",X"04",X"12",X"45",X"04",X"12",X"44",X"12",X"FD",X"20",X"44",
		X"00",X"12",X"FD",X"6C",X"14",X"6D",X"14",X"6E",X"0A",X"42",X"DD",X"43",X"01",X"4A",X"10",X"46",
		X"00",X"4B",X"18",X"4C",X"06",X"66",X"9C",X"FE",X"E1",X"9D",X"47",X"BF",X"FF",X"40",X"6C",X"41",
		X"00",X"42",X"D9",X"43",X"00",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"30",X"68",X"0F",X"69",X"0F",
		X"0D",X"09",X"18",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"18",X"40",X"90",X"42",X"21",X"43",X"01",
		X"68",X"0F",X"69",X"0F",X"0D",X"09",X"30",X"40",X"7A",X"42",X"F3",X"43",X"00",X"68",X"0F",X"69",
		X"0F",X"0D",X"09",X"18",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"18",X"68",X"0F",X"69",X"0F",X"0D",
		X"09",X"30",X"40",X"90",X"42",X"21",X"43",X"01",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"18",X"68",
		X"0F",X"69",X"0F",X"0D",X"09",X"18",X"40",X"7A",X"42",X"F3",X"43",X"00",X"68",X"0F",X"69",X"0F",
		X"0D",X"09",X"30",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"18",X"68",X"0F",X"69",X"0F",X"0D",X"09",
		X"18",X"40",X"90",X"42",X"21",X"43",X"01",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"30",X"40",X"A1",
		X"42",X"43",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"18",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"18",
		X"40",X"AB",X"42",X"56",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"30",X"40",X"D9",X"42",X"B2",X"68",
		X"0F",X"69",X"0F",X"0D",X"09",X"18",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"18",X"68",X"0F",X"69",
		X"0F",X"0D",X"09",X"30",X"40",X"7A",X"42",X"F3",X"43",X"00",X"68",X"0F",X"69",X"0F",X"0D",X"09",
		X"18",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"18",X"40",X"6C",X"42",X"D9",X"68",X"0F",X"69",X"0F",
		X"0D",X"09",X"18",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"18",X"68",X"00",X"69",X"00",X"0D",X"09",
		X"18",X"68",X"00",X"69",X"00",X"0D",X"09",X"18",X"FD",X"66",X"F8",X"48",X"10",X"49",X"00",X"4B",
		X"00",X"4C",X"0A",X"20",X"48",X"00",X"24",X"20",X"60",X"00",X"24",X"20",X"7A",X"00",X"18",X"20",
		X"4D",X"00",X"24",X"20",X"66",X"00",X"24",X"20",X"81",X"00",X"18",X"20",X"50",X"00",X"24",X"20",
		X"6C",X"00",X"24",X"20",X"88",X"00",X"18",X"20",X"56",X"00",X"24",X"20",X"73",X"00",X"24",X"20",
		X"90",X"00",X"18",X"20",X"60",X"00",X"48",X"20",X"6C",X"00",X"18",X"20",X"73",X"00",X"48",X"20",
		X"90",X"00",X"18",X"20",X"90",X"00",X"60",X"20",X"21",X"01",X"30",X"48",X"00",X"49",X"00",X"4A",
		X"00",X"20",X"00",X"00",X"30",X"67",X"07",X"FF",X"76",X"BD",X"59",X"10",X"5B",X"00",X"5C",X"01",
		X"5D",X"0D",X"53",X"00",X"12",X"2D",X"20",X"12",X"3D",X"20",X"12",X"2D",X"20",X"12",X"3D",X"20",
		X"12",X"2D",X"20",X"12",X"3D",X"20",X"59",X"00",X"5C",X"00",X"77",X"02",X"FF",X"22",X"04",X"12",
		X"00",X"04",X"53",X"01",X"12",X"C2",X"04",X"12",X"00",X"04",X"12",X"D0",X"04",X"12",X"00",X"04",
		X"12",X"E6",X"04",X"12",X"00",X"04",X"12",X"FF",X"04",X"12",X"00",X"04",X"53",X"02",X"12",X"22",
		X"04",X"12",X"00",X"04",X"12",X"65",X"04",X"12",X"00",X"04",X"12",X"3E",X"04",X"12",X"00",X"04",
		X"12",X"84",X"04",X"12",X"00",X"04",X"12",X"AB",X"04",X"12",X"00",X"04",X"12",X"D0",X"04",X"12",
		X"00",X"04",X"12",X"FB",X"04",X"12",X"00",X"04",X"59",X"00",X"5C",X"00",X"77",X"02",X"FF",X"76",
		X"BD",X"52",X"36",X"53",X"00",X"19",X"0F",X"18",X"59",X"00",X"77",X"06",X"FF",X"24",X"19",X"00",
		X"24",X"19",X"0F",X"24",X"19",X"00",X"24",X"19",X"0F",X"24",X"19",X"00",X"24",X"59",X"00",X"77",
		X"06",X"FF",X"76",X"BB",X"5A",X"10",X"5B",X"00",X"5C",X"0A",X"55",X"00",X"54",X"33",X"1D",X"09",
		X"12",X"54",X"39",X"1D",X"09",X"12",X"54",X"40",X"1D",X"09",X"12",X"54",X"4D",X"1D",X"09",X"12",
		X"5A",X"00",X"77",X"04",X"FF",X"54",X"81",X"1D",X"09",X"18",X"54",X"88",X"1D",X"09",X"0C",X"54",
		X"81",X"1D",X"09",X"18",X"54",X"88",X"1D",X"09",X"0C",X"54",X"81",X"1D",X"09",X"18",X"54",X"88",
		X"1D",X"09",X"0C",X"54",X"81",X"1D",X"09",X"18",X"5A",X"00",X"77",X"04",X"FF",X"76",X"AF",X"59",
		X"0F",X"53",X"00",X"52",X"56",X"16",X"2A",X"03",X"16",X"2D",X"03",X"16",X"30",X"03",X"16",X"33",
		X"03",X"16",X"36",X"03",X"16",X"39",X"03",X"16",X"3D",X"03",X"16",X"40",X"03",X"16",X"44",X"03",
		X"16",X"48",X"03",X"16",X"4D",X"03",X"16",X"50",X"03",X"16",X"56",X"03",X"16",X"5B",X"03",X"16",
		X"60",X"03",X"16",X"66",X"03",X"16",X"6C",X"03",X"16",X"73",X"03",X"16",X"7A",X"03",X"16",X"81",
		X"03",X"16",X"88",X"03",X"16",X"90",X"03",X"59",X"00",X"77",X"B8",X"FF",X"03",X"16",X"AB",X"03",
		X"16",X"B6",X"03",X"16",X"C1",X"03",X"16",X"CB",X"03",X"16",X"D9",X"03",X"16",X"E5",X"03",X"16",
		X"F3",X"03",X"16",X"FB",X"03",X"59",X"00",X"77",X"B8",X"FF",X"5D",X"00",X"77",X"B8",X"FF",X"77",
		X"B8",X"FF",X"46",X"10",X"66",X"C7",X"48",X"10",X"49",X"10",X"4A",X"10",X"4B",X"10",X"4C",X"09",
		X"40",X"32",X"41",X"01",X"0D",X"09",X"C0",X"67",X"38",X"FF",X"76",X"BD",X"59",X"10",X"5B",X"00",
		X"5C",X"01",X"5D",X"0D",X"53",X"00",X"12",X"2A",X"12",X"12",X"20",X"12",X"12",X"26",X"12",X"12",
		X"1C",X"12",X"59",X"00",X"5C",X"00",X"77",X"02",X"FF",X"0F",X"09",X"19",X"00",X"03",X"19",X"0F",
		X"09",X"19",X"00",X"03",X"19",X"0F",X"09",X"19",X"00",X"03",X"19",X"0F",X"09",X"19",X"00",X"03",
		X"19",X"0F",X"09",X"19",X"00",X"03",X"59",X"00",X"77",X"06",X"FF",X"6C",X"14",X"6D",X"14",X"6E",
		X"0A",X"4A",X"10",X"46",X"00",X"4B",X"00",X"4C",X"04",X"66",X"9C",X"FE",X"E4",X"B7",X"FE",X"E4",
		X"B7",X"FE",X"E5",X"4D",X"FE",X"E4",X"AB",X"40",X"90",X"41",X"00",X"42",X"7F",X"43",X"04",X"68",
		X"0F",X"69",X"0F",X"0D",X"09",X"30",X"69",X"00",X"0D",X"09",X"18",X"0D",X"09",X"18",X"40",X"C1",
		X"42",X"7F",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"30",X"40",X"81",X"68",X"0F",X"69",X"00",X"0D",
		X"09",X"18",X"0D",X"09",X"18",X"42",X"7F",X"69",X"0F",X"0D",X"09",X"30",X"40",X"A1",X"68",X"0F",
		X"69",X"00",X"0D",X"09",X"18",X"0D",X"09",X"18",X"40",X"90",X"42",X"7F",X"68",X"0F",X"69",X"0F",
		X"0D",X"09",X"30",X"69",X"00",X"0D",X"09",X"18",X"0D",X"09",X"18",X"40",X"C1",X"42",X"7F",X"68",
		X"0F",X"69",X"0F",X"0D",X"09",X"30",X"40",X"D9",X"68",X"0F",X"69",X"00",X"0D",X"09",X"18",X"0D",
		X"09",X"18",X"42",X"7F",X"69",X"0F",X"0D",X"09",X"30",X"40",X"F3",X"68",X"0F",X"69",X"00",X"0D",
		X"09",X"18",X"0D",X"09",X"18",X"40",X"D9",X"42",X"7F",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"30",
		X"40",X"C1",X"68",X"0F",X"69",X"00",X"0D",X"09",X"18",X"0D",X"09",X"18",X"FD",X"40",X"F3",X"42",
		X"7F",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"30",X"69",X"00",X"0D",X"09",X"18",X"0D",X"09",X"18",
		X"40",X"21",X"41",X"01",X"42",X"7F",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"30",X"40",X"D9",X"41",
		X"00",X"68",X"0F",X"69",X"00",X"0D",X"09",X"18",X"0D",X"04",X"18",X"42",X"7F",X"69",X"0F",X"0D",
		X"09",X"30",X"40",X"C1",X"68",X"0F",X"69",X"00",X"0D",X"09",X"18",X"0D",X"09",X"18",X"42",X"7F",
		X"69",X"0F",X"0D",X"09",X"30",X"40",X"21",X"41",X"01",X"68",X"0F",X"69",X"00",X"0D",X"09",X"18",
		X"0D",X"09",X"18",X"40",X"21",X"42",X"7F",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"30",X"69",X"00",
		X"0D",X"09",X"18",X"0D",X"09",X"18",X"40",X"F3",X"41",X"00",X"42",X"7F",X"68",X"0F",X"69",X"0F",
		X"0D",X"09",X"30",X"40",X"D9",X"68",X"0F",X"69",X"00",X"0D",X"09",X"18",X"0D",X"09",X"18",X"42",
		X"7F",X"69",X"0F",X"0D",X"09",X"30",X"40",X"C1",X"68",X"0F",X"69",X"00",X"0D",X"09",X"18",X"0D",
		X"09",X"18",X"40",X"A1",X"42",X"7F",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"30",X"40",X"90",X"68",
		X"0F",X"69",X"00",X"0D",X"09",X"18",X"0D",X"09",X"18",X"FD",X"10",X"20",X"B6",X"00",X"18",X"68",
		X"00",X"49",X"00",X"4A",X"00",X"20",X"00",X"00",X"0C",X"68",X"0F",X"49",X"10",X"4A",X"10",X"20",
		X"B6",X"00",X"18",X"68",X"00",X"49",X"00",X"4A",X"00",X"20",X"00",X"00",X"0C",X"68",X"0F",X"49",
		X"10",X"4A",X"10",X"20",X"B6",X"00",X"18",X"68",X"00",X"49",X"00",X"4A",X"00",X"20",X"00",X"00",
		X"0C",X"68",X"0F",X"49",X"10",X"4A",X"10",X"20",X"04",X"01",X"18",X"68",X"00",X"49",X"00",X"4A",
		X"00",X"20",X"00",X"00",X"0C",X"68",X"0F",X"49",X"10",X"4A",X"10",X"20",X"04",X"01",X"18",X"68",
		X"00",X"49",X"00",X"4A",X"00",X"20",X"00",X"00",X"0C",X"68",X"0F",X"49",X"10",X"4A",X"10",X"20",
		X"04",X"01",X"18",X"68",X"00",X"49",X"00",X"4A",X"00",X"20",X"00",X"00",X"0C",X"68",X"0F",X"49",
		X"10",X"4A",X"10",X"20",X"04",X"01",X"24",X"68",X"00",X"49",X"00",X"4A",X"00",X"20",X"00",X"00",
		X"0C",X"68",X"0F",X"49",X"10",X"4A",X"10",X"20",X"04",X"01",X"24",X"68",X"00",X"49",X"00",X"4A",
		X"00",X"20",X"00",X"00",X"0C",X"68",X"0F",X"49",X"10",X"4A",X"10",X"20",X"04",X"01",X"24",X"68",
		X"00",X"49",X"00",X"4A",X"00",X"20",X"00",X"00",X"0C",X"68",X"0F",X"49",X"10",X"4A",X"10",X"20",
		X"F3",X"00",X"24",X"68",X"00",X"49",X"00",X"4A",X"00",X"20",X"00",X"00",X"0C",X"68",X"0F",X"49",
		X"10",X"4A",X"10",X"20",X"F3",X"00",X"24",X"68",X"00",X"49",X"00",X"4A",X"00",X"20",X"00",X"00",
		X"0C",X"68",X"0F",X"49",X"10",X"4A",X"10",X"20",X"D9",X"00",X"24",X"68",X"00",X"49",X"00",X"4A",
		X"00",X"20",X"00",X"00",X"0C",X"68",X"0F",X"49",X"10",X"4A",X"10",X"20",X"C1",X"00",X"30",X"68",
		X"00",X"49",X"00",X"4A",X"00",X"20",X"00",X"00",X"60",X"67",X"07",X"FF",X"66",X"B9",X"6C",X"14",
		X"6D",X"14",X"6E",X"0A",X"FE",X"E7",X"0A",X"FE",X"E7",X"04",X"42",X"5B",X"43",X"00",X"45",X"01",
		X"69",X"0E",X"6A",X"0E",X"04",X"6C",X"30",X"69",X"00",X"6A",X"00",X"04",X"00",X"30",X"42",X"5B",
		X"45",X"00",X"69",X"0E",X"6A",X"0E",X"04",X"B6",X"30",X"69",X"00",X"6A",X"00",X"04",X"00",X"30",
		X"42",X"88",X"45",X"01",X"69",X"0E",X"6A",X"0E",X"04",X"10",X"30",X"69",X"0E",X"6A",X"00",X"04",
		X"00",X"18",X"42",X"7A",X"69",X"0E",X"6A",X"00",X"04",X"00",X"18",X"42",X"6C",X"45",X"00",X"69",
		X"0E",X"6A",X"0E",X"04",X"D9",X"30",X"69",X"00",X"6A",X"00",X"04",X"00",X"30",X"42",X"5B",X"45",
		X"01",X"69",X"0E",X"6A",X"0E",X"04",X"6C",X"30",X"69",X"00",X"6A",X"00",X"04",X"00",X"30",X"42",
		X"5B",X"45",X"00",X"69",X"0E",X"6A",X"0E",X"04",X"B6",X"30",X"69",X"00",X"6A",X"00",X"04",X"00",
		X"30",X"42",X"88",X"45",X"01",X"69",X"0E",X"6A",X"0E",X"04",X"10",X"30",X"69",X"0E",X"6A",X"00",
		X"04",X"00",X"18",X"42",X"7A",X"69",X"0E",X"6A",X"00",X"04",X"00",X"18",X"42",X"6C",X"45",X"00",
		X"69",X"0E",X"6A",X"0E",X"04",X"D9",X"24",X"42",X"60",X"69",X"0E",X"6A",X"00",X"04",X"00",X"24",
		X"42",X"5B",X"69",X"0E",X"6A",X"00",X"04",X"00",X"18",X"42",X"60",X"45",X"01",X"69",X"0E",X"6A",
		X"0E",X"04",X"7F",X"30",X"69",X"00",X"6A",X"00",X"04",X"00",X"30",X"42",X"60",X"45",X"00",X"69",
		X"0E",X"6A",X"0E",X"04",X"C1",X"30",X"69",X"00",X"6A",X"00",X"04",X"00",X"30",X"42",X"90",X"45",
		X"01",X"69",X"0E",X"6A",X"0E",X"04",X"21",X"30",X"69",X"0E",X"6A",X"00",X"04",X"00",X"18",X"42",
		X"88",X"69",X"0E",X"6A",X"00",X"04",X"00",X"18",X"42",X"7A",X"45",X"00",X"69",X"0E",X"6A",X"0E",
		X"04",X"F3",X"30",X"69",X"00",X"6A",X"00",X"04",X"00",X"30",X"42",X"60",X"45",X"01",X"69",X"0E",
		X"6A",X"0E",X"04",X"7F",X"30",X"69",X"00",X"6A",X"00",X"04",X"00",X"30",X"42",X"60",X"45",X"00",
		X"69",X"0E",X"6A",X"0E",X"04",X"C1",X"30",X"69",X"00",X"6A",X"00",X"04",X"00",X"30",X"42",X"90",
		X"45",X"01",X"69",X"0E",X"6A",X"0E",X"04",X"21",X"30",X"69",X"0E",X"6A",X"00",X"04",X"00",X"18",
		X"42",X"88",X"69",X"0E",X"6A",X"00",X"04",X"00",X"18",X"42",X"7A",X"45",X"00",X"69",X"0E",X"6A",
		X"0E",X"04",X"F3",X"24",X"42",X"6C",X"69",X"0E",X"6A",X"00",X"04",X"00",X"24",X"42",X"60",X"69",
		X"0E",X"6A",X"00",X"04",X"00",X"18",X"FD",X"66",X"B9",X"6D",X"14",X"6E",X"0A",X"FE",X"E8",X"7C",
		X"FE",X"E8",X"7C",X"FE",X"E9",X"89",X"FE",X"E9",X"89",X"FE",X"E8",X"6D",X"42",X"90",X"43",X"00",
		X"45",X"01",X"69",X"0E",X"6A",X"0E",X"04",X"B2",X"30",X"42",X"A1",X"69",X"0E",X"6A",X"0E",X"04",
		X"B2",X"30",X"42",X"AB",X"69",X"0E",X"6A",X"0E",X"04",X"B2",X"30",X"42",X"D9",X"69",X"0E",X"6A",
		X"0E",X"04",X"B2",X"30",X"69",X"00",X"6A",X"0E",X"04",X"B2",X"30",X"69",X"00",X"6A",X"0E",X"04",
		X"B2",X"30",X"42",X"7A",X"69",X"0E",X"6A",X"0E",X"04",X"E6",X"30",X"42",X"81",X"69",X"0E",X"6A",
		X"0E",X"04",X"E6",X"30",X"42",X"90",X"69",X"0E",X"6A",X"0E",X"04",X"E6",X"30",X"42",X"A1",X"69",
		X"0E",X"6A",X"0E",X"04",X"E6",X"30",X"69",X"00",X"6A",X"0E",X"04",X"E6",X"30",X"42",X"81",X"69",
		X"0E",X"6A",X"0E",X"04",X"E6",X"30",X"42",X"7A",X"69",X"0E",X"6A",X"0E",X"04",X"E6",X"30",X"42",
		X"6C",X"69",X"0E",X"6A",X"0E",X"04",X"E6",X"30",X"42",X"60",X"69",X"0E",X"6A",X"0E",X"04",X"E6",
		X"30",X"69",X"00",X"6A",X"0E",X"04",X"E6",X"30",X"42",X"6C",X"69",X"0E",X"6A",X"0E",X"04",X"B2",
		X"30",X"69",X"00",X"6A",X"0E",X"04",X"B2",X"30",X"42",X"81",X"69",X"0E",X"6A",X"0E",X"04",X"B2",
		X"30",X"69",X"00",X"6A",X"0E",X"04",X"B2",X"30",X"69",X"00",X"6A",X"0E",X"04",X"B2",X"30",X"69",
		X"00",X"6A",X"0E",X"04",X"B2",X"30",X"69",X"00",X"6A",X"0E",X"04",X"B2",X"30",X"42",X"6C",X"69",
		X"0E",X"6A",X"0E",X"04",X"B2",X"30",X"42",X"60",X"69",X"0E",X"6A",X"0E",X"04",X"E6",X"30",X"69",
		X"00",X"6A",X"0E",X"04",X"E6",X"30",X"42",X"7A",X"69",X"0E",X"6A",X"0E",X"04",X"E6",X"30",X"42",
		X"6C",X"69",X"0E",X"6A",X"0E",X"04",X"E6",X"30",X"69",X"00",X"6A",X"0E",X"04",X"E6",X"30",X"42",
		X"81",X"69",X"0E",X"6A",X"0E",X"04",X"E6",X"30",X"42",X"7A",X"69",X"0E",X"6A",X"0E",X"04",X"E6",
		X"30",X"69",X"00",X"6A",X"0E",X"04",X"E6",X"30",X"FD",X"42",X"6C",X"45",X"01",X"69",X"0E",X"6A",
		X"0E",X"04",X"43",X"18",X"69",X"00",X"6A",X"00",X"04",X"00",X"18",X"42",X"40",X"69",X"0E",X"6A",
		X"0E",X"04",X"43",X"18",X"69",X"00",X"6A",X"00",X"04",X"00",X"18",X"42",X"50",X"69",X"0E",X"6A",
		X"0E",X"04",X"43",X"18",X"69",X"00",X"6A",X"00",X"04",X"00",X"18",X"42",X"6C",X"69",X"0E",X"6A",
		X"0E",X"04",X"43",X"18",X"69",X"00",X"6A",X"00",X"04",X"00",X"18",X"42",X"40",X"69",X"0E",X"6A",
		X"0E",X"04",X"43",X"18",X"69",X"00",X"6A",X"00",X"04",X"00",X"18",X"42",X"50",X"69",X"0E",X"6A",
		X"0E",X"04",X"43",X"18",X"69",X"00",X"6A",X"00",X"04",X"00",X"18",X"42",X"D9",X"69",X"0E",X"6A",
		X"0E",X"04",X"43",X"18",X"69",X"00",X"6A",X"00",X"04",X"00",X"18",X"42",X"40",X"69",X"0E",X"6A",
		X"0E",X"04",X"43",X"18",X"69",X"00",X"6A",X"00",X"04",X"00",X"18",X"42",X"50",X"69",X"0E",X"6A",
		X"0E",X"04",X"6C",X"18",X"69",X"00",X"6A",X"00",X"04",X"00",X"18",X"42",X"6C",X"69",X"0E",X"6A",
		X"0E",X"04",X"6C",X"18",X"69",X"00",X"6A",X"00",X"04",X"00",X"18",X"42",X"40",X"69",X"0E",X"6A",
		X"0E",X"04",X"6C",X"18",X"69",X"00",X"6A",X"00",X"04",X"00",X"18",X"42",X"50",X"69",X"0E",X"6A",
		X"0E",X"04",X"6C",X"18",X"69",X"00",X"6A",X"00",X"04",X"00",X"18",X"42",X"6C",X"69",X"0E",X"6A",
		X"0E",X"04",X"6C",X"18",X"69",X"00",X"6A",X"00",X"04",X"00",X"18",X"42",X"40",X"69",X"0E",X"6A",
		X"0E",X"04",X"6C",X"18",X"69",X"00",X"6A",X"00",X"04",X"00",X"18",X"42",X"50",X"69",X"0E",X"6A",
		X"0E",X"04",X"6C",X"18",X"69",X"00",X"6A",X"00",X"04",X"00",X"18",X"42",X"6C",X"69",X"0E",X"6A",
		X"0E",X"04",X"6C",X"18",X"69",X"00",X"6A",X"00",X"04",X"00",X"18",X"42",X"48",X"69",X"0E",X"6A",
		X"0E",X"04",X"B2",X"18",X"69",X"00",X"6A",X"00",X"04",X"00",X"18",X"42",X"56",X"69",X"0E",X"6A",
		X"0E",X"04",X"B2",X"18",X"69",X"00",X"6A",X"00",X"04",X"00",X"18",X"42",X"6C",X"69",X"0E",X"6A",
		X"0E",X"04",X"B2",X"18",X"69",X"00",X"6A",X"00",X"04",X"00",X"18",X"42",X"48",X"69",X"0E",X"6A",
		X"0E",X"04",X"B2",X"18",X"69",X"00",X"6A",X"00",X"04",X"00",X"18",X"42",X"56",X"69",X"0E",X"6A",
		X"0E",X"04",X"B2",X"18",X"69",X"00",X"6A",X"00",X"04",X"00",X"18",X"42",X"6C",X"69",X"0E",X"6A",
		X"0E",X"04",X"B2",X"18",X"69",X"00",X"6A",X"00",X"04",X"00",X"18",X"42",X"48",X"69",X"0E",X"6A",
		X"0E",X"04",X"B2",X"18",X"69",X"00",X"6A",X"00",X"04",X"00",X"18",X"42",X"56",X"69",X"0E",X"6A",
		X"0E",X"04",X"B2",X"18",X"69",X"00",X"6A",X"00",X"04",X"00",X"18",X"42",X"6C",X"45",X"02",X"69",
		X"0E",X"6A",X"0E",X"04",X"3E",X"18",X"69",X"00",X"6A",X"00",X"04",X"00",X"18",X"42",X"48",X"69",
		X"0E",X"6A",X"0E",X"04",X"3E",X"18",X"69",X"00",X"6A",X"00",X"04",X"00",X"18",X"42",X"56",X"69",
		X"0E",X"6A",X"0E",X"04",X"3E",X"18",X"69",X"00",X"6A",X"00",X"04",X"00",X"18",X"42",X"6C",X"69",
		X"0E",X"6A",X"0E",X"04",X"3E",X"18",X"69",X"00",X"6A",X"00",X"04",X"00",X"18",X"42",X"48",X"69",
		X"0E",X"6A",X"0E",X"04",X"3E",X"18",X"69",X"00",X"6A",X"00",X"04",X"00",X"18",X"42",X"56",X"69",
		X"0E",X"6A",X"0E",X"04",X"3E",X"18",X"69",X"00",X"6A",X"00",X"04",X"00",X"18",X"42",X"D9",X"69",
		X"0E",X"6A",X"0E",X"04",X"3E",X"18",X"69",X"00",X"6A",X"00",X"04",X"00",X"18",X"42",X"90",X"69",
		X"0E",X"6A",X"0E",X"04",X"3E",X"18",X"69",X"00",X"6A",X"00",X"04",X"00",X"18",X"FD",X"6C",X"14",
		X"6D",X"14",X"6E",X"0A",X"4A",X"00",X"46",X"00",X"4B",X"00",X"4C",X"00",X"66",X"9C",X"FE",X"EB",
		X"A4",X"47",X"BF",X"FF",X"40",X"7A",X"41",X"00",X"42",X"E6",X"43",X"01",X"68",X"0F",X"69",X"0F",
		X"0D",X"09",X"24",X"42",X"43",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"0C",X"40",X"A1",X"68",X"0F",
		X"69",X"0F",X"0D",X"09",X"18",X"40",X"88",X"42",X"10",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"24",
		X"42",X"43",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"0C",X"40",X"7A",X"68",X"0F",X"69",X"0F",X"0D",
		X"09",X"18",X"42",X"E6",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"24",X"42",X"43",X"68",X"0F",X"69",
		X"0F",X"0D",X"09",X"0C",X"40",X"88",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"18",X"40",X"90",X"42",
		X"6C",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"18",X"40",X"A1",X"68",X"0F",X"69",X"0F",X"0D",X"09",
		X"0C",X"42",X"43",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"0C",X"40",X"88",X"68",X"0F",X"69",X"0F",
		X"0D",X"09",X"18",X"40",X"7A",X"42",X"E6",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"24",X"42",X"6C",
		X"68",X"0F",X"69",X"0F",X"0D",X"09",X"0C",X"40",X"B6",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"18",
		X"40",X"90",X"42",X"21",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"24",X"42",X"6C",X"68",X"0F",X"69",
		X"0F",X"0D",X"09",X"0C",X"40",X"7A",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"18",X"42",X"E6",X"68",
		X"0F",X"69",X"0F",X"0D",X"09",X"24",X"42",X"43",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"0C",X"40",
		X"88",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"18",X"40",X"90",X"42",X"6C",X"68",X"0F",X"69",X"0F",
		X"0D",X"09",X"18",X"40",X"A1",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"0C",X"42",X"43",X"68",X"0F",
		X"69",X"0F",X"0D",X"09",X"0C",X"40",X"88",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"18",X"40",X"7A",
		X"42",X"E6",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"24",X"42",X"6C",X"68",X"0F",X"69",X"0F",X"0D",
		X"09",X"0C",X"40",X"90",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"18",X"40",X"66",X"42",X"92",X"68",
		X"0F",X"69",X"0F",X"0D",X"09",X"18",X"68",X"00",X"69",X"0F",X"0D",X"09",X"0C",X"42",X"D9",X"43",
		X"00",X"68",X"00",X"69",X"0F",X"0D",X"09",X"0C",X"40",X"6C",X"68",X"0F",X"69",X"0F",X"0D",X"09",
		X"18",X"42",X"B2",X"43",X"01",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"18",X"68",X"00",X"69",X"0F",
		X"0D",X"09",X"0C",X"42",X"F3",X"43",X"00",X"68",X"00",X"69",X"0F",X"0D",X"09",X"0C",X"40",X"7A",
		X"68",X"0F",X"69",X"0F",X"0D",X"09",X"18",X"42",X"E6",X"43",X"01",X"68",X"0F",X"69",X"0F",X"0D",
		X"09",X"24",X"42",X"10",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"0C",X"40",X"88",X"68",X"0F",X"69",
		X"0F",X"0D",X"09",X"18",X"42",X"22",X"43",X"02",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"24",X"42",
		X"43",X"43",X"01",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"0C",X"40",X"A1",X"68",X"0F",X"69",X"0F",
		X"0D",X"09",X"18",X"40",X"90",X"42",X"21",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"24",X"42",X"B2",
		X"68",X"0F",X"69",X"0F",X"0D",X"09",X"0C",X"40",X"88",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"18",
		X"42",X"43",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"24",X"42",X"21",X"68",X"0F",X"69",X"0F",X"0D",
		X"09",X"0C",X"40",X"90",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"18",X"40",X"A1",X"42",X"43",X"68",
		X"0F",X"69",X"0F",X"0D",X"09",X"24",X"42",X"22",X"43",X"02",X"68",X"0F",X"69",X"0F",X"0D",X"09",
		X"0C",X"40",X"D9",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"18",X"40",X"F3",X"42",X"E6",X"43",X"01",
		X"68",X"0F",X"69",X"0F",X"0D",X"09",X"18",X"40",X"D9",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"18",
		X"40",X"C1",X"68",X"0F",X"69",X"00",X"0D",X"09",X"18",X"40",X"B6",X"42",X"6C",X"68",X"0F",X"69",
		X"0F",X"0D",X"09",X"18",X"40",X"A1",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"18",X"40",X"90",X"68",
		X"0F",X"69",X"00",X"0D",X"09",X"18",X"40",X"88",X"42",X"10",X"68",X"0F",X"69",X"0F",X"0D",X"09",
		X"18",X"40",X"7A",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"18",X"40",X"6C",X"68",X"0F",X"69",X"00",
		X"0D",X"09",X"18",X"40",X"60",X"42",X"C1",X"43",X"00",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"18",
		X"40",X"5B",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"18",X"40",X"50",X"68",X"0F",X"69",X"00",X"0D",
		X"09",X"18",X"40",X"5B",X"42",X"B6",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"30",X"40",X"50",X"42",
		X"A1",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"18",X"40",X"5B",X"42",X"B6",X"68",X"0F",X"69",X"0F",
		X"0D",X"09",X"24",X"68",X"00",X"69",X"00",X"0D",X"09",X"0C",X"40",X"5B",X"42",X"B6",X"68",X"0F",
		X"69",X"0F",X"0D",X"09",X"48",X"40",X"50",X"42",X"A1",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"18",
		X"40",X"5B",X"42",X"B6",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"24",X"68",X"00",X"69",X"00",X"0D",
		X"09",X"0C",X"40",X"44",X"42",X"88",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"48",X"40",X"48",X"42",
		X"90",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"18",X"40",X"50",X"42",X"A1",X"68",X"0F",X"69",X"0F",
		X"0D",X"09",X"30",X"40",X"5B",X"42",X"B6",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"60",X"FD",X"44",
		X"B2",X"69",X"00",X"6A",X"0E",X"02",X"00",X"30",X"44",X"43",X"69",X"0E",X"6A",X"0E",X"02",X"81",
		X"30",X"44",X"B2",X"69",X"00",X"6A",X"0E",X"02",X"00",X"30",X"44",X"B2",X"69",X"0E",X"6A",X"0E",
		X"02",X"90",X"30",X"44",X"B2",X"69",X"00",X"6A",X"0E",X"02",X"00",X"30",X"44",X"B2",X"69",X"00",
		X"6A",X"0E",X"02",X"00",X"30",X"44",X"E6",X"69",X"0E",X"6A",X"0E",X"02",X"7A",X"30",X"44",X"E6",
		X"69",X"00",X"6A",X"0E",X"02",X"00",X"30",X"44",X"B2",X"69",X"0E",X"6A",X"0E",X"02",X"81",X"30",
		X"44",X"B2",X"69",X"00",X"6A",X"0E",X"02",X"00",X"30",X"44",X"B2",X"69",X"0E",X"6A",X"0E",X"02",
		X"90",X"30",X"44",X"B2",X"69",X"00",X"6A",X"0E",X"02",X"00",X"30",X"44",X"B2",X"69",X"0E",X"6A",
		X"0E",X"02",X"90",X"30",X"44",X"7F",X"69",X"0E",X"6A",X"0E",X"02",X"A1",X"30",X"44",X"56",X"69",
		X"0E",X"6A",X"0E",X"02",X"AB",X"30",X"FD",X"76",X"BB",X"5A",X"0F",X"55",X"02",X"54",X"22",X"14",
		X"AB",X"03",X"14",X"65",X"03",X"55",X"01",X"14",X"FF",X"03",X"14",X"C2",X"03",X"14",X"92",X"03",
		X"14",X"56",X"03",X"14",X"32",X"03",X"14",X"04",X"03",X"55",X"00",X"14",X"E5",X"03",X"14",X"CB",
		X"03",X"5A",X"00",X"77",X"04",X"FF",X"14",X"D9",X"03",X"14",X"F3",X"03",X"14",X"E5",X"03",X"5A",
		X"00",X"77",X"04",X"FF",X"6A",X"03",X"14",X"8F",X"03",X"14",X"D0",X"03",X"14",X"E0",X"03",X"5A",
		X"00",X"77",X"04",X"FF",X"8F",X"32",X"38",X"DF",X"84",X"97",X"A4",X"7F",X"00",X"80",X"7F",X"00",
		X"8C",X"86",X"BE",X"9A",X"BA",X"97",X"BA",X"39",X"81",X"22",X"2A",X"03",X"7E",X"FF",X"67",X"80",
		X"20",X"97",X"DB",X"39",X"81",X"0E",X"26",X"08",X"7F",X"00",X"D9",X"39",X"86",X"03",X"97",X"DC",
		X"86",X"0C",X"97",X"DB",X"86",X"01",X"97",X"D9",X"39",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FA",X"80",X"FA",X"80",X"FA",X"80",X"FA",X"80",X"FC",X"6D",X"FA",X"80",X"FB",X"59",X"FA",X"80",
		X"6C",X"14",X"6D",X"14",X"6E",X"0A",X"42",X"6A",X"43",X"03",X"4A",X"10",X"46",X"00",X"4B",X"00",
		X"4C",X"04",X"66",X"9C",X"FE",X"F0",X"17",X"68",X"00",X"69",X"0F",X"0D",X"09",X"30",X"68",X"00",
		X"69",X"00",X"0D",X"09",X"18",X"0D",X"09",X"18",X"FE",X"F0",X"14",X"29",X"0F",X"30",X"42",X"B2",
		X"68",X"00",X"29",X"0F",X"30",X"42",X"B2",X"68",X"00",X"29",X"0F",X"30",X"40",X"43",X"41",X"01",
		X"42",X"84",X"43",X"02",X"68",X"0F",X"29",X"0F",X"30",X"40",X"10",X"42",X"84",X"68",X"0F",X"29",
		X"0F",X"30",X"42",X"22",X"68",X"0F",X"29",X"0F",X"30",X"42",X"22",X"68",X"00",X"29",X"0F",X"30",
		X"42",X"FF",X"43",X"01",X"68",X"00",X"29",X"0F",X"30",X"42",X"FF",X"68",X"00",X"29",X"0F",X"30",
		X"42",X"E6",X"68",X"00",X"29",X"0F",X"30",X"42",X"E6",X"68",X"00",X"29",X"0F",X"30",X"40",X"43",
		X"42",X"84",X"43",X"02",X"68",X"0F",X"29",X"0F",X"30",X"40",X"10",X"42",X"84",X"68",X"0F",X"29",
		X"0F",X"30",X"42",X"22",X"68",X"0F",X"29",X"0F",X"30",X"42",X"22",X"68",X"00",X"29",X"0F",X"30",
		X"40",X"43",X"42",X"FF",X"43",X"01",X"68",X"0F",X"29",X"0F",X"30",X"40",X"10",X"42",X"FF",X"68",
		X"0F",X"29",X"0F",X"30",X"42",X"E6",X"68",X"0F",X"29",X"0F",X"30",X"40",X"43",X"42",X"E6",X"68",
		X"0F",X"29",X"0F",X"30",X"42",X"22",X"43",X"02",X"68",X"00",X"29",X"0F",X"30",X"40",X"43",X"42",
		X"22",X"68",X"0F",X"29",X"0F",X"30",X"42",X"3E",X"68",X"00",X"29",X"0F",X"30",X"40",X"56",X"42",
		X"3E",X"68",X"0F",X"29",X"0F",X"30",X"42",X"65",X"68",X"00",X"29",X"0F",X"30",X"40",X"56",X"42",
		X"65",X"68",X"0F",X"29",X"0F",X"30",X"68",X"00",X"29",X"00",X"30",X"40",X"6C",X"42",X"D5",X"68",
		X"0F",X"29",X"0F",X"30",X"40",X"6C",X"42",X"D5",X"68",X"0F",X"29",X"0F",X"30",X"68",X"00",X"29",
		X"00",X"30",X"FD",X"76",X"BB",X"5A",X"10",X"5B",X"00",X"5C",X"10",X"55",X"00",X"54",X"7A",X"1D",
		X"09",X"30",X"5A",X"00",X"1D",X"09",X"C0",X"5A",X"10",X"1D",X"09",X"30",X"5A",X"00",X"1D",X"09",
		X"C0",X"5A",X"10",X"1D",X"09",X"30",X"5A",X"00",X"1D",X"09",X"C0",X"5A",X"10",X"54",X"3D",X"1D",
		X"09",X"C0",X"5A",X"00",X"77",X"04",X"FF",X"6C",X"14",X"6D",X"14",X"6E",X"0A",X"4A",X"00",X"46",
		X"00",X"4B",X"00",X"4C",X"00",X"66",X"9C",X"FE",X"F1",X"72",X"FE",X"F1",X"72",X"FE",X"F1",X"72",
		X"FE",X"F1",X"72",X"FE",X"F1",X"C7",X"FE",X"F1",X"C7",X"FE",X"F1",X"C7",X"FE",X"F2",X"20",X"FE",
		X"F1",X"57",X"40",X"88",X"41",X"00",X"42",X"FF",X"43",X"01",X"68",X"0F",X"69",X"0F",X"0D",X"09",
		X"0C",X"40",X"81",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"24",X"40",X"88",X"42",X"04",X"68",X"0F",
		X"69",X"0F",X"0D",X"09",X"18",X"40",X"81",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"18",X"40",X"60",
		X"42",X"FF",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"18",X"40",X"81",X"68",X"0F",X"69",X"0F",X"0D",
		X"09",X"18",X"40",X"88",X"42",X"04",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"18",X"40",X"81",X"68",
		X"0F",X"69",X"0F",X"0D",X"09",X"18",X"FD",X"40",X"A1",X"42",X"65",X"43",X"02",X"68",X"0F",X"69",
		X"0F",X"0D",X"09",X"0C",X"40",X"99",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"24",X"40",X"A1",X"42",
		X"32",X"43",X"01",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"18",X"40",X"99",X"68",X"0F",X"69",X"0F",
		X"0D",X"09",X"18",X"40",X"73",X"42",X"65",X"43",X"02",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"18",
		X"40",X"99",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"18",X"40",X"A1",X"42",X"32",X"43",X"01",X"68",
		X"0F",X"69",X"0F",X"0D",X"09",X"18",X"40",X"99",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"18",X"FD",
		X"40",X"A1",X"42",X"65",X"43",X"02",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"0C",X"40",X"99",X"68",
		X"0F",X"69",X"0F",X"0D",X"09",X"24",X"40",X"A1",X"42",X"32",X"43",X"01",X"68",X"0F",X"69",X"0F",
		X"0D",X"09",X"18",X"40",X"99",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"18",X"40",X"73",X"42",X"65",
		X"43",X"02",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"18",X"40",X"99",X"68",X"0F",X"69",X"0F",X"0D",
		X"09",X"18",X"40",X"90",X"42",X"32",X"43",X"01",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"18",X"40",
		X"88",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"18",X"40",X"88",X"42",X"FF",X"68",X"0F",X"69",X"0F",
		X"0D",X"09",X"0C",X"40",X"81",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"24",X"40",X"88",X"42",X"04",
		X"68",X"0F",X"69",X"0F",X"0D",X"09",X"0C",X"40",X"81",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"24",
		X"40",X"66",X"42",X"FF",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"0C",X"40",X"60",X"68",X"0F",X"69",
		X"0F",X"0D",X"09",X"24",X"40",X"88",X"42",X"04",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"0C",X"40",
		X"81",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"24",X"40",X"A1",X"42",X"65",X"43",X"02",X"68",X"0F",
		X"69",X"0F",X"0D",X"09",X"0C",X"40",X"99",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"24",X"40",X"A1",
		X"42",X"32",X"43",X"01",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"0C",X"40",X"99",X"68",X"0F",X"69",
		X"0F",X"0D",X"09",X"24",X"40",X"7A",X"42",X"65",X"43",X"02",X"68",X"0F",X"69",X"0F",X"0D",X"09",
		X"0C",X"40",X"73",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"24",X"40",X"A1",X"42",X"32",X"43",X"01",
		X"68",X"0F",X"69",X"0F",X"0D",X"09",X"0C",X"40",X"99",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"24",
		X"40",X"88",X"42",X"FF",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"0C",X"40",X"81",X"68",X"0F",X"69",
		X"0F",X"0D",X"09",X"24",X"40",X"B6",X"42",X"AB",X"43",X"02",X"68",X"0F",X"69",X"0F",X"0D",X"09",
		X"0C",X"40",X"AB",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"24",X"40",X"A1",X"42",X"65",X"68",X"0F",
		X"69",X"0F",X"0D",X"09",X"0C",X"42",X"99",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"24",X"40",X"D9",
		X"42",X"29",X"43",X"03",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"0C",X"40",X"CB",X"68",X"0F",X"69",
		X"0F",X"0D",X"09",X"24",X"40",X"B6",X"42",X"AB",X"43",X"02",X"68",X"0F",X"69",X"0F",X"0D",X"09",
		X"0C",X"40",X"AB",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"24",X"40",X"F3",X"42",X"8F",X"43",X"03",
		X"68",X"0F",X"69",X"0F",X"0D",X"09",X"0C",X"40",X"E5",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"24",
		X"40",X"D9",X"42",X"29",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"0C",X"40",X"CB",X"68",X"0F",X"69",
		X"0F",X"0D",X"09",X"24",X"40",X"10",X"41",X"01",X"42",X"01",X"43",X"04",X"68",X"0F",X"69",X"0F",
		X"0D",X"09",X"0C",X"40",X"04",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"24",X"FD",X"54",X"69",X"0E",
		X"6A",X"0E",X"04",X"58",X"30",X"42",X"4F",X"69",X"0E",X"6A",X"0E",X"04",X"7D",X"30",X"42",X"59",
		X"69",X"0E",X"6A",X"0E",X"04",X"38",X"30",X"42",X"5E",X"69",X"0E",X"6A",X"0E",X"04",X"16",X"30",
		X"42",X"6A",X"45",X"01",X"69",X"0E",X"6A",X"0E",X"04",X"FC",X"30",X"FD",X"76",X"BB",X"55",X"00",
		X"54",X"70",X"5A",X"10",X"5B",X"00",X"5C",X"08",X"1D",X"09",X"E0",X"5A",X"00",X"77",X"04",X"FF",
		X"76",X"BD",X"52",X"20",X"53",X"00",X"19",X"0F",X"60",X"59",X"00",X"77",X"06",X"FF",X"76",X"BD",
		X"52",X"7F",X"53",X"00",X"19",X"0F",X"30",X"19",X"00",X"90",X"19",X"0F",X"30",X"19",X"00",X"90",
		X"19",X"0F",X"30",X"19",X"00",X"90",X"52",X"2F",X"19",X"0F",X"70",X"59",X"00",X"77",X"06",X"FF",
		X"66",X"F8",X"48",X"10",X"49",X"00",X"4B",X"00",X"4C",X"0A",X"20",X"9F",X"00",X"20",X"20",X"5E",
		X"00",X"20",X"20",X"9F",X"00",X"20",X"20",X"A8",X"00",X"20",X"20",X"64",X"00",X"20",X"20",X"A8",
		X"00",X"20",X"20",X"B3",X"00",X"20",X"20",X"6A",X"00",X"20",X"20",X"B3",X"00",X"20",X"42",X"77",
		X"43",X"00",X"6D",X"10",X"69",X"0F",X"20",X"BD",X"00",X"40",X"67",X"02",X"20",X"9F",X"00",X"20",
		X"20",X"8E",X"00",X"20",X"0D",X"09",X"20",X"20",X"86",X"00",X"80",X"67",X"07",X"FF",X"66",X"FC",
		X"6C",X"14",X"6D",X"14",X"FE",X"F4",X"CB",X"02",X"1C",X"20",X"40",X"8E",X"68",X"0F",X"29",X"0F",
		X"20",X"40",X"7E",X"42",X"51",X"68",X"0F",X"29",X"0F",X"40",X"40",X"8E",X"68",X"0F",X"29",X"0F",
		X"20",X"FE",X"F4",X"CB",X"42",X"FC",X"29",X"0F",X"20",X"29",X"0F",X"20",X"42",X"DD",X"29",X"0F",
		X"40",X"42",X"C1",X"68",X"0F",X"29",X"0F",X"20",X"FE",X"F4",X"94",X"40",X"6A",X"41",X"00",X"42",
		X"A9",X"43",X"01",X"68",X"0F",X"29",X"0F",X"40",X"40",X"8E",X"68",X"0F",X"29",X"0F",X"20",X"40",
		X"7E",X"42",X"51",X"68",X"0F",X"29",X"0F",X"40",X"40",X"77",X"68",X"0F",X"29",X"0F",X"20",X"42",
		X"1C",X"29",X"0F",X"20",X"FD",X"FE",X"F4",X"94",X"66",X"F8",X"68",X"0F",X"49",X"10",X"4A",X"10",
		X"4B",X"00",X"4C",X"10",X"6C",X"14",X"FE",X"F5",X"0F",X"FE",X"F5",X"0F",X"67",X"07",X"FF",X"20",
		X"6A",X"00",X"30",X"20",X"7E",X"00",X"30",X"20",X"8E",X"00",X"30",X"20",X"6A",X"00",X"60",X"FD",
		X"76",X"BB",X"5A",X"0F",X"55",X"00",X"54",X"58",X"14",X"50",X"04",X"14",X"59",X"04",X"14",X"57",
		X"04",X"14",X"5F",X"04",X"14",X"56",X"04",X"14",X"55",X"04",X"14",X"59",X"04",X"14",X"56",X"04",
		X"14",X"5A",X"04",X"14",X"57",X"04",X"14",X"50",X"04",X"14",X"5C",X"04",X"14",X"59",X"04",X"14",
		X"57",X"04",X"14",X"53",X"04",X"14",X"5C",X"04",X"14",X"58",X"04",X"5A",X"00",X"77",X"04",X"FF",
		X"76",X"BB",X"55",X"00",X"54",X"38",X"5A",X"0F",X"14",X"36",X"04",X"14",X"38",X"04",X"14",X"36",
		X"04",X"14",X"3A",X"04",X"14",X"33",X"04",X"14",X"37",X"04",X"14",X"3F",X"04",X"14",X"36",X"04",
		X"14",X"38",X"04",X"14",X"3C",X"04",X"14",X"34",X"04",X"14",X"39",X"04",X"14",X"3F",X"04",X"14",
		X"35",X"04",X"14",X"3D",X"04",X"14",X"38",X"04",X"14",X"33",X"04",X"14",X"3F",X"04",X"5A",X"00",
		X"77",X"04",X"FF",X"76",X"AF",X"59",X"10",X"5C",X"01",X"5D",X"0D",X"16",X"1E",X"01",X"16",X"1D",
		X"01",X"16",X"1C",X"01",X"16",X"1B",X"01",X"16",X"1A",X"01",X"16",X"19",X"01",X"16",X"18",X"01",
		X"16",X"17",X"01",X"16",X"16",X"01",X"16",X"15",X"01",X"16",X"14",X"01",X"16",X"13",X"01",X"16",
		X"12",X"01",X"16",X"11",X"01",X"16",X"10",X"01",X"5B",X"A1",X"5C",X"07",X"5D",X"09",X"16",X"0F",
		X"01",X"16",X"FE",X"01",X"16",X"0D",X"01",X"16",X"0C",X"01",X"16",X"0B",X"01",X"16",X"0A",X"01",
		X"16",X"09",X"01",X"16",X"08",X"01",X"16",X"07",X"01",X"16",X"06",X"01",X"16",X"05",X"01",X"16",
		X"04",X"01",X"16",X"03",X"01",X"16",X"02",X"01",X"16",X"01",X"01",X"56",X"00",X"59",X"00",X"5B",
		X"00",X"5C",X"00",X"5D",X"00",X"77",X"B8",X"FF",X"76",X"BB",X"55",X"00",X"54",X"70",X"5A",X"10",
		X"5B",X"00",X"5C",X"10",X"1D",X"09",X"E0",X"5A",X"00",X"77",X"04",X"FF",X"6C",X"14",X"6D",X"14",
		X"6E",X"0A",X"42",X"DD",X"43",X"01",X"4A",X"10",X"46",X"00",X"4B",X"00",X"4C",X"04",X"66",X"9C",
		X"FE",X"F6",X"46",X"47",X"BF",X"FF",X"40",X"9F",X"41",X"00",X"42",X"D4",X"43",X"00",X"68",X"0F",
		X"69",X"0F",X"0D",X"09",X"15",X"0D",X"09",X"15",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"15",X"40",
		X"FD",X"42",X"65",X"43",X"01",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"15",X"0D",X"09",X"15",X"0D",
		X"09",X"15",X"40",X"EE",X"42",X"3E",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"15",X"0D",X"09",X"15",
		X"0D",X"09",X"15",X"40",X"E1",X"42",X"2C",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"15",X"0D",X"09",
		X"15",X"0D",X"09",X"15",X"40",X"D4",X"42",X"1C",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"15",X"0D",
		X"09",X"15",X"0D",X"09",X"15",X"40",X"BD",X"42",X"FD",X"43",X"00",X"68",X"0F",X"69",X"0F",X"0D",
		X"09",X"15",X"0D",X"09",X"15",X"0D",X"09",X"15",X"40",X"B3",X"42",X"EE",X"68",X"0F",X"69",X"0F",
		X"0D",X"09",X"15",X"0D",X"09",X"15",X"0D",X"09",X"15",X"40",X"A8",X"42",X"E1",X"68",X"0F",X"69",
		X"0F",X"0D",X"09",X"15",X"0D",X"09",X"15",X"0D",X"09",X"15",X"40",X"9F",X"42",X"D4",X"68",X"0F",
		X"69",X"0F",X"0D",X"09",X"15",X"0D",X"09",X"15",X"0D",X"09",X"15",X"40",X"7E",X"42",X"B3",X"68",
		X"0F",X"69",X"0F",X"0D",X"09",X"15",X"0D",X"09",X"15",X"0D",X"09",X"15",X"40",X"77",X"42",X"9F",
		X"68",X"0F",X"69",X"0F",X"0D",X"09",X"15",X"0D",X"09",X"15",X"0D",X"09",X"15",X"40",X"70",X"42",
		X"96",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"15",X"0D",X"09",X"15",X"0D",X"09",X"15",X"40",X"6A",
		X"42",X"8E",X"69",X"0F",X"68",X"0F",X"0D",X"09",X"15",X"0D",X"09",X"15",X"0D",X"09",X"15",X"40",
		X"5E",X"42",X"7E",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"15",X"0D",X"09",X"15",X"0D",X"09",X"15",
		X"40",X"59",X"42",X"77",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"15",X"0D",X"09",X"15",X"0D",X"09",
		X"15",X"40",X"54",X"42",X"70",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"15",X"0D",X"09",X"15",X"0D",
		X"09",X"15",X"40",X"4F",X"42",X"6A",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"15",X"0D",X"09",X"15",
		X"0D",X"09",X"15",X"FD",X"66",X"F8",X"68",X"0F",X"49",X"10",X"4A",X"10",X"4B",X"00",X"4C",X"10",
		X"20",X"9F",X"00",X"30",X"20",X"BD",X"00",X"18",X"20",X"EE",X"00",X"48",X"20",X"BD",X"00",X"48",
		X"20",X"9F",X"00",X"48",X"20",X"77",X"00",X"90",X"20",X"5E",X"00",X"30",X"20",X"6A",X"00",X"18",
		X"20",X"77",X"00",X"48",X"20",X"BD",X"00",X"48",X"20",X"A8",X"00",X"48",X"20",X"9F",X"00",X"90",
		X"20",X"9F",X"00",X"24",X"20",X"9F",X"00",X"24",X"20",X"5E",X"00",X"60",X"20",X"6A",X"00",X"18",
		X"20",X"77",X"00",X"48",X"20",X"7E",X"00",X"90",X"20",X"8E",X"00",X"24",X"20",X"7E",X"00",X"24",
		X"20",X"77",X"00",X"48",X"20",X"77",X"00",X"48",X"20",X"9F",X"00",X"48",X"20",X"EE",X"00",X"90",
		X"FE",X"F7",X"80",X"46",X"10",X"66",X"C7",X"48",X"10",X"49",X"10",X"4A",X"10",X"4B",X"00",X"4C",
		X"0A",X"0D",X"09",X"20",X"67",X"38",X"FF",X"80",X"88",X"08",X"80",X"80",X"80",X"80",X"00",X"81",
		X"80",X"80",X"90",X"80",X"04",X"41",X"FF",X"8C",X"D7",X"24",X"0A",X"E8",X"08",X"29",X"80",X"22",
		X"E0",X"81",X"51",X"CC",X"0B",X"42",X"00",X"58",X"A9",X"EA",X"02",X"51",X"29",X"A9",X"BC",X"91",
		X"27",X"38",X"9A",X"B9",X"0B",X"17",X"03",X"8A",X"C0",X"80",X"00",X"00",X"49",X"B0",X"00",X"60",
		X"D9",X"0A",X"40",X"00",X"58",X"AA",X"CA",X"15",X"21",X"29",X"AA",X"CE",X"01",X"17",X"08",X"98",
		X"A8",X"8A",X"15",X"21",X"9A",X"B8",X"00",X"92",X"10",X"7A",X"A0",X"00",X"40",X"E8",X"08",X"28",
		X"01",X"59",X"9C",X"BA",X"27",X"01",X"29",X"A9",X"CC",X"02",X"37",X"09",X"89",X"B8",X"98",X"26",
		X"38",X"AA",X"A8",X"08",X"83",X"14",X"3F",X"90",X"80",X"4A",X"98",X"00",X"00",X"02",X"79",X"9D",
		X"99",X"34",X"02",X"19",X"B9",X"FB",X"12",X"53",X"0A",X"99",X"D8",X"A1",X"27",X"18",X"9A",X"A0",
		X"09",X"13",X"05",X"0D",X"90",X"00",X"3C",X"80",X"18",X"80",X"02",X"79",X"BB",X"AA",X"72",X"82",
		X"2A",X"A9",X"FA",X"12",X"43",X"0A",X"9A",X"D9",X"91",X"47",X"09",X"8A",X"90",X"8A",X"32",X"14",
		X"9C",X"90",X"80",X"3B",X"00",X"5B",X"80",X"02",X"79",X"D8",X"98",X"50",X"83",X"09",X"AB",X"F8",
		X"14",X"12",X"89",X"9A",X"CB",X"02",X"57",X"88",X"99",X"98",X"89",X"32",X"31",X"AE",X"80",X"80",
		X"18",X"00",X"5C",X"80",X"02",X"3C",X"C0",X"A2",X"30",X"06",X"0A",X"9E",X"B0",X"25",X"03",X"8A",
		X"9A",X"DA",X"12",X"72",X"89",X"9B",X"90",X"A0",X"61",X"39",X"9C",X"88",X"00",X"00",X"04",X"0D",
		X"08",X"03",X"2E",X"90",X"A3",X"10",X"07",X"89",X"AC",X"B1",X"43",X"04",X"8A",X"9C",X"D8",X"12",
		X"71",X"98",X"9A",X"98",X"91",X"52",X"19",X"9C",X"88",X"09",X"30",X"16",X"AB",X"00",X"03",X"2F",
		X"88",X"82",X"00",X"87",X"89",X"BA",X"B1",X"71",X"02",X"99",X"9B",X"F0",X"12",X"50",X"89",X"9B",
		X"8A",X"82",X"72",X"09",X"AB",X"80",X"0A",X"50",X"13",X"CA",X"80",X"04",X"9B",X"00",X"00",X"01",
		X"07",X"1B",X"E9",X"A3",X"50",X"12",X"9A",X"AF",X"A0",X"25",X"30",X"A9",X"9C",X"8B",X"12",X"72",
		X"89",X"9B",X"80",X"A1",X"58",X"40",X"C9",X"80",X"04",X"B8",X"01",X"88",X"00",X"17",X"8B",X"B9",
		X"B7",X"10",X"21",X"9A",X"9F",X"A1",X"24",X"30",X"A9",X"AD",X"9A",X"22",X"72",X"8A",X"9B",X"08",
		X"B3",X"50",X"48",X"C9",X"08",X"02",X"A0",X"05",X"B8",X"00",X"07",X"8C",X"98",X"95",X"00",X"11",
		X"99",X"AF",X"91",X"41",X"20",X"A9",X"9D",X"A0",X"13",X"71",X"99",X"9B",X"08",X"A3",X"43",X"2A",
		X"DA",X"00",X"00",X"81",X"07",X"B8",X"80",X"00",X"00",X"00",X"01",X"F7",X"F7",X"01",X"80",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"F4",X"8D",X"F4",X"8D",X"EF",
		X"17",X"F1",X"13",X"E4",X"5A",X"E3",X"82",X"E2",X"E8",X"E3",X"5F",X"E0",X"00",X"E0",X"9D",X"EF",
		X"17",X"E3",X"CD",X"F0",X"00",X"E2",X"89",X"E1",X"83",X"E1",X"43",X"E4",X"9B",X"E4",X"42",X"EB",
		X"8E",X"E6",X"FC",X"F1",X"47",X"E8",X"67",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"8E",X"00",X"FF",X"BD",X"FC",X"7A",X"86",X"BF",X"C6",X"07",X"BD",X"FC",X"BA",X"86",X"13",
		X"C6",X"0F",X"BD",X"FC",X"BA",X"BD",X"FC",X"8F",X"7F",X"90",X"00",X"0F",X"BD",X"FB",X"C8",X"96",
		X"BC",X"2B",X"07",X"BD",X"FE",X"C3",X"86",X"FF",X"97",X"BC",X"0E",X"CE",X"00",X"00",X"DF",X"D1",
		X"96",X"80",X"26",X"0B",X"DE",X"84",X"D6",X"8C",X"BD",X"FD",X"BE",X"DF",X"84",X"97",X"80",X"7C",
		X"00",X"D2",X"96",X"81",X"26",X"0B",X"DE",X"86",X"D6",X"8D",X"BD",X"FD",X"BE",X"DF",X"86",X"97",
		X"81",X"7C",X"00",X"D2",X"96",X"82",X"26",X"0B",X"DE",X"88",X"D6",X"8E",X"BD",X"FD",X"BE",X"DF",
		X"88",X"97",X"82",X"7C",X"00",X"D2",X"96",X"83",X"26",X"0B",X"DE",X"8A",X"D6",X"8F",X"BD",X"FD",
		X"BE",X"DF",X"8A",X"97",X"83",X"96",X"A8",X"27",X"08",X"7F",X"00",X"A8",X"C6",X"08",X"BD",X"FD",
		X"1C",X"96",X"A9",X"27",X"08",X"7F",X"00",X"A9",X"C6",X"09",X"BD",X"FD",X"1C",X"96",X"AA",X"27",
		X"08",X"7F",X"00",X"AA",X"C6",X"0A",X"BD",X"FD",X"1C",X"96",X"AB",X"27",X"08",X"7F",X"00",X"AB",
		X"C6",X"18",X"BD",X"FD",X"35",X"96",X"AC",X"27",X"08",X"7F",X"00",X"AC",X"C6",X"19",X"BD",X"FD",
		X"35",X"96",X"AD",X"27",X"08",X"7F",X"00",X"AD",X"C6",X"1A",X"BD",X"FD",X"35",X"96",X"BE",X"16",
		X"9A",X"D8",X"0F",X"97",X"D8",X"54",X"24",X"09",X"D6",X"CB",X"C1",X"02",X"26",X"03",X"5C",X"D7",
		X"BC",X"C6",X"0F",X"BD",X"FC",X"C0",X"7E",X"FA",X"9B",X"96",X"C1",X"B7",X"08",X"01",X"96",X"C2",
		X"B7",X"08",X"02",X"7C",X"00",X"BD",X"96",X"BF",X"4C",X"97",X"BF",X"44",X"24",X"32",X"DE",X"C3",
		X"09",X"27",X"1E",X"DF",X"C3",X"DE",X"C7",X"A6",X"00",X"44",X"44",X"44",X"44",X"97",X"C1",X"DE",
		X"C5",X"09",X"27",X"15",X"DF",X"C5",X"DE",X"C9",X"A6",X"00",X"44",X"44",X"44",X"44",X"97",X"C2",
		X"3B",X"86",X"01",X"9A",X"BE",X"97",X"BE",X"20",X"E6",X"86",X"02",X"9A",X"BE",X"97",X"BE",X"3B",
		X"96",X"C7",X"81",X"A0",X"25",X"09",X"DE",X"C7",X"A6",X"00",X"97",X"C1",X"08",X"DF",X"C7",X"96",
		X"C9",X"81",X"A0",X"25",X"09",X"DE",X"C9",X"A6",X"00",X"97",X"C2",X"08",X"DF",X"C9",X"96",X"BF",
		X"84",X"0E",X"26",X"CC",X"7C",X"00",X"C0",X"3B",X"96",X"C0",X"27",X"41",X"7A",X"00",X"C0",X"BD",
		X"FC",X"19",X"96",X"80",X"27",X"06",X"4C",X"27",X"03",X"7A",X"00",X"80",X"96",X"81",X"27",X"06",
		X"4C",X"27",X"03",X"7A",X"00",X"81",X"96",X"82",X"27",X"06",X"4C",X"27",X"03",X"7A",X"00",X"82",
		X"96",X"83",X"27",X"06",X"4C",X"27",X"03",X"7A",X"00",X"83",X"CE",X"00",X"06",X"A6",X"AD",X"27",
		X"09",X"4A",X"26",X"04",X"6C",X"A7",X"A6",X"B3",X"A7",X"AD",X"09",X"26",X"F0",X"39",X"C6",X"17",
		X"96",X"BB",X"8A",X"B1",X"97",X"BB",X"7E",X"FC",X"C0",X"96",X"D9",X"98",X"DA",X"27",X"13",X"96",
		X"D9",X"97",X"DA",X"27",X"E9",X"C6",X"17",X"96",X"BB",X"8A",X"BE",X"84",X"BE",X"97",X"BB",X"BD",
		X"FC",X"C0",X"DE",X"DC",X"96",X"DB",X"91",X"DC",X"27",X"2F",X"2A",X"08",X"09",X"09",X"09",X"09",
		X"09",X"7E",X"FC",X"47",X"C6",X"0A",X"3A",X"DF",X"DC",X"96",X"D9",X"27",X"C0",X"D6",X"09",X"D4",
		X"7F",X"3A",X"DF",X"D5",X"96",X"D5",X"C6",X"11",X"BD",X"FC",X"C0",X"96",X"D6",X"C6",X"10",X"BD",
		X"FC",X"C0",X"86",X"0F",X"C6",X"18",X"7E",X"FC",X"C0",X"7F",X"00",X"D9",X"39",X"B7",X"90",X"00",
		X"C6",X"0E",X"BD",X"FD",X"02",X"84",X"3F",X"97",X"BC",X"3B",X"CE",X"FF",X"FF",X"DF",X"00",X"C6",
		X"4F",X"08",X"86",X"00",X"A7",X"80",X"08",X"5A",X"26",X"FA",X"86",X"13",X"97",X"D8",X"39",X"BD",
		X"FC",X"A5",X"86",X"BF",X"97",X"BB",X"C6",X"FF",X"D7",X"82",X"D7",X"B1",X"D7",X"B2",X"D7",X"B3",
		X"C6",X"17",X"7E",X"FC",X"C0",X"86",X"BF",X"97",X"BA",X"C6",X"FF",X"D7",X"80",X"D7",X"81",X"D7",
		X"AE",X"D7",X"AF",X"D7",X"B0",X"C6",X"07",X"7E",X"FC",X"C0",X"7C",X"00",X"BD",X"20",X"04",X"0F",
		X"7F",X"00",X"BD",X"37",X"36",X"C1",X"10",X"2A",X"19",X"86",X"0D",X"97",X"03",X"D7",X"02",X"C6",
		X"08",X"D7",X"03",X"5C",X"32",X"97",X"02",X"96",X"BD",X"27",X"FC",X"D7",X"03",X"5A",X"D7",X"03",
		X"33",X"39",X"86",X"15",X"97",X"03",X"C4",X"0F",X"D7",X"02",X"C6",X"10",X"20",X"E3",X"37",X"20",
		X"E4",X"37",X"86",X"15",X"97",X"03",X"C4",X"0F",X"D7",X"02",X"C6",X"14",X"20",X"0D",X"C1",X"10",
		X"2A",X"EF",X"37",X"86",X"0D",X"97",X"03",X"D7",X"02",X"C6",X"0C",X"4F",X"97",X"03",X"97",X"00",
		X"D7",X"03",X"96",X"02",X"5F",X"D7",X"03",X"5A",X"D7",X"00",X"33",X"39",X"0F",X"BD",X"FD",X"02",
		X"C6",X"09",X"7F",X"00",X"BD",X"84",X"1F",X"81",X"10",X"2A",X"08",X"4A",X"81",X"07",X"2B",X"03",
		X"BD",X"FC",X"EE",X"0E",X"39",X"0F",X"BD",X"FC",X"F1",X"C6",X"11",X"20",X"E5",X"17",X"84",X"0F",
		X"81",X"08",X"2A",X"08",X"A6",X"94",X"AB",X"98",X"A7",X"94",X"20",X"67",X"CB",X"38",X"DE",X"CD",
		X"A6",X"05",X"36",X"DE",X"D1",X"AB",X"94",X"A7",X"94",X"32",X"2B",X"0C",X"24",X"02",X"6C",X"98",
		X"BD",X"FC",X"BF",X"5C",X"A6",X"94",X"20",X"4B",X"25",X"F6",X"6A",X"98",X"20",X"F2",X"6F",X"8C",
		X"DE",X"CD",X"C1",X"A0",X"2B",X"02",X"08",X"08",X"08",X"08",X"08",X"C1",X"C0",X"2B",X"08",X"17",
		X"84",X"0F",X"81",X"08",X"2B",X"01",X"08",X"86",X"01",X"39",X"DF",X"CD",X"DE",X"D1",X"6A",X"90",
		X"27",X"DC",X"C1",X"A0",X"2A",X"10",X"C4",X"1F",X"A6",X"94",X"36",X"DE",X"CD",X"A6",X"03",X"BD",
		X"FC",X"BF",X"0E",X"32",X"08",X"39",X"C1",X"C0",X"2A",X"93",X"A6",X"90",X"44",X"A6",X"94",X"25",
		X"02",X"A6",X"98",X"C4",X"1F",X"BD",X"FC",X"BF",X"0E",X"DE",X"CD",X"A6",X"04",X"39",X"26",X"CA",
		X"DF",X"CD",X"E6",X"00",X"2A",X"03",X"7E",X"FE",X"75",X"C4",X"3F",X"C1",X"20",X"2A",X"11",X"A6",
		X"01",X"BD",X"FC",X"BF",X"0E",X"E6",X"00",X"08",X"08",X"58",X"2B",X"E4",X"A6",X"00",X"08",X"39",
		X"C4",X"1F",X"17",X"84",X"0F",X"26",X"31",X"A6",X"01",X"97",X"CE",X"A6",X"02",X"97",X"CD",X"BD",
		X"FE",X"B6",X"DC",X"CD",X"04",X"DD",X"CD",X"E6",X"00",X"C4",X"1F",X"5C",X"5C",X"BD",X"FE",X"B6",
		X"7C",X"00",X"CE",X"26",X"03",X"7C",X"00",X"CD",X"BD",X"FE",X"B6",X"CB",X"07",X"86",X"09",X"BD",
		X"FC",X"C0",X"0E",X"E6",X"00",X"08",X"20",X"BF",X"80",X"08",X"2B",X"29",X"DD",X"CF",X"84",X"03",
		X"C1",X"30",X"2B",X"02",X"8B",X"03",X"16",X"A6",X"01",X"CE",X"00",X"00",X"3A",X"D6",X"CF",X"C1",
		X"04",X"2A",X"0B",X"A6",X"B4",X"A7",X"AE",X"DE",X"CD",X"D6",X"D0",X"7E",X"FD",X"CF",X"A7",X"B4",
		X"DE",X"CD",X"7E",X"FD",X"D5",X"4C",X"27",X"17",X"5C",X"C1",X"10",X"2A",X"09",X"96",X"BA",X"A4",
		X"01",X"97",X"BA",X"7E",X"FD",X"D1",X"96",X"BB",X"A4",X"01",X"97",X"BB",X"7E",X"FD",X"D1",X"C1",
		X"10",X"2A",X"09",X"96",X"BA",X"AA",X"01",X"97",X"BA",X"7E",X"FD",X"D1",X"96",X"BB",X"AA",X"01",
		X"97",X"BB",X"7E",X"FD",X"D1",X"C1",X"F0",X"2A",X"17",X"A6",X"01",X"EE",X"02",X"3C",X"DE",X"D1",
		X"E7",X"8C",X"4C",X"A7",X"90",X"32",X"A7",X"94",X"32",X"A7",X"98",X"DE",X"CD",X"86",X"01",X"39",
		X"5C",X"27",X"12",X"DE",X"D1",X"5C",X"26",X"10",X"DC",X"CD",X"A7",X"9C",X"E7",X"A0",X"DE",X"CD",
		X"EE",X"01",X"86",X"01",X"39",X"86",X"FF",X"39",X"A6",X"9C",X"E6",X"A0",X"DD",X"CD",X"DE",X"CD",
		X"08",X"08",X"08",X"86",X"01",X"39",X"96",X"CE",X"BD",X"FC",X"BF",X"5C",X"96",X"CD",X"BD",X"FC",
		X"C0",X"5C",X"39",X"26",X"0E",X"BD",X"FC",X"7A",X"7F",X"00",X"D9",X"CE",X"0F",X"00",X"DF",X"DC",
		X"7E",X"FC",X"8F",X"81",X"0E",X"2B",X"03",X"7E",X"FF",X"0F",X"97",X"CB",X"96",X"D8",X"8A",X"01",
		X"16",X"C4",X"FE",X"D7",X"D8",X"C6",X"0F",X"BD",X"FC",X"C0",X"86",X"05",X"7F",X"00",X"BD",X"D6",
		X"BD",X"27",X"FC",X"4A",X"26",X"F6",X"D6",X"CB",X"58",X"58",X"CE",X"F9",X"77",X"3A",X"3C",X"EE",
		X"00",X"DF",X"C7",X"38",X"EE",X"02",X"DF",X"C3",X"96",X"BE",X"84",X"02",X"97",X"BE",X"39",X"16",
		X"58",X"CE",X"F9",X"9F",X"3A",X"EE",X"00",X"81",X"10",X"2B",X"21",X"27",X"6F",X"81",X"16",X"2A",
		X"1C",X"D6",X"82",X"5C",X"27",X"06",X"91",X"A6",X"27",X"02",X"2A",X"10",X"97",X"A6",X"DF",X"88",
		X"7F",X"00",X"82",X"7F",X"00",X"8E",X"C6",X"B8",X"DA",X"BB",X"D7",X"BB",X"39",X"81",X"15",X"27",
		X"26",X"81",X"1A",X"2A",X"11",X"DF",X"8A",X"97",X"A7",X"7F",X"00",X"83",X"7F",X"00",X"8F",X"86",
		X"BE",X"9A",X"BB",X"97",X"BB",X"39",X"81",X"20",X"2A",X"1E",X"3C",X"36",X"BD",X"FC",X"7A",X"7F",
		X"00",X"D9",X"BD",X"FC",X"8F",X"32",X"38",X"DF",X"84",X"97",X"A4",X"7F",X"00",X"80",X"7F",X"00",
		X"8C",X"86",X"BE",X"9A",X"BA",X"97",X"BA",X"39",X"81",X"24",X"2A",X"03",X"7E",X"FF",X"67",X"80",
		X"20",X"97",X"DB",X"39",X"81",X"0E",X"26",X"08",X"7F",X"00",X"D9",X"39",X"86",X"03",X"97",X"DC",
		X"86",X"0C",X"97",X"DB",X"86",X"01",X"97",X"D9",X"39",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FA",X"80",X"FA",X"80",X"FA",X"80",X"FA",X"80",X"FC",X"6D",X"FA",X"80",X"FB",X"59",X"FA",X"80");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
