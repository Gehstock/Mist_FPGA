library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity twotiger_bg_bits_2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of twotiger_bg_bits_2 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"55",X"5A",X"55",X"5A",X"55",X"5A",X"55",X"5A",X"7E",X"AA",X"56",X"AA",
		X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",
		X"AB",X"CA",X"AE",X"B2",X"75",X"71",X"55",X"71",X"75",X"51",X"75",X"75",X"55",X"55",X"55",X"55",
		X"55",X"6A",X"55",X"6A",X"55",X"6A",X"55",X"6A",X"55",X"6A",X"55",X"6A",X"55",X"6A",X"55",X"6A",
		X"AA",X"A6",X"AA",X"AE",X"A6",X"66",X"A9",X"AE",X"A9",X"A6",X"55",X"AE",X"56",X"A6",X"55",X"DE",
		X"56",X"AA",X"56",X"AA",X"56",X"AA",X"56",X"AA",X"56",X"AA",X"56",X"AA",X"56",X"AA",X"56",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",
		X"5A",X"AA",X"5A",X"BE",X"59",X"EA",X"57",X"AA",X"5F",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",
		X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"6A",X"55",X"6A",X"75",X"5A",X"7D",X"56",X"55",X"55",
		X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AB",X"EA",X"AF",X"AA",X"5E",X"AA",X"56",X"AA",
		X"55",X"55",X"55",X"55",X"55",X"5A",X"75",X"5A",X"75",X"DA",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"5A",X"55",X"5A",X"55",X"5A",X"55",X"5A",X"AA",X"AA",X"AA",X"BA",X"AB",X"AA",X"BA",X"AA",
		X"55",X"5A",X"55",X"5A",X"55",X"5A",X"55",X"5A",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"55",X"56",X"55",X"56",X"55",X"56",X"55",X"56",X"55",X"56",X"55",X"56",
		X"55",X"AA",X"55",X"AA",X"56",X"AA",X"55",X"55",X"55",X"55",X"55",X"55",X"5D",X"55",X"55",X"55",
		X"55",X"56",X"55",X"56",X"55",X"56",X"55",X"56",X"55",X"56",X"55",X"56",X"55",X"56",X"55",X"56",
		X"55",X"6A",X"55",X"6A",X"55",X"5A",X"55",X"5A",X"55",X"56",X"55",X"56",X"55",X"55",X"55",X"55",
		X"A5",X"55",X"B9",X"5D",X"A9",X"55",X"EA",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"6A",X"55",X"5A",X"55",X"6A",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A5",X"AA",X"A5",X"AA",X"A6",
		X"AA",X"A6",X"AA",X"9A",X"AA",X"9A",X"AA",X"9A",X"AA",X"9A",X"AA",X"9A",X"AA",X"9A",X"AA",X"9A",
		X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",
		X"AA",X"6A",X"AA",X"6A",X"AA",X"6A",X"AA",X"5A",X"AA",X"56",X"AA",X"56",X"AA",X"96",X"AA",X"96",
		X"AA",X"9A",X"AA",X"A6",X"AA",X"A6",X"AA",X"A6",X"AA",X"A6",X"AA",X"A9",X"AA",X"A9",X"AA",X"A9",
		X"AA",X"A9",X"AA",X"A9",X"AA",X"A9",X"AA",X"A6",X"AA",X"A6",X"AA",X"A6",X"AA",X"A6",X"AA",X"9A",
		X"AA",X"9A",X"AA",X"99",X"AA",X"6A",X"AA",X"6A",X"AA",X"6A",X"AA",X"6A",X"AA",X"5A",X"AA",X"5A",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"55",X"6A",X"A9",X"AA",X"A6",X"AA",X"9A",X"AA",X"9A",X"AA",
		X"AA",X"AA",X"AA",X"A9",X"AA",X"A9",X"AA",X"A6",X"AA",X"A6",X"AA",X"9A",X"AA",X"9A",X"AA",X"9A",
		X"AA",X"6A",X"AA",X"6A",X"AA",X"6A",X"AA",X"6A",X"A9",X"AA",X"A9",X"AA",X"A9",X"AA",X"A9",X"AA",
		X"A6",X"AA",X"96",X"AA",X"A6",X"AA",X"A6",X"AA",X"A6",X"AA",X"A6",X"AA",X"A6",X"AA",X"A6",X"AA",
		X"9A",X"AA",X"9A",X"AA",X"9A",X"AA",X"9A",X"AA",X"9A",X"AA",X"9A",X"AA",X"9A",X"AA",X"9A",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"55",X"5A",X"AA",X"6A",X"A9",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A6",X"AA",X"9A",X"AA",X"6A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"99",X"99",X"A9",X"56",X"A5",X"65",X"9A",X"55",X"A9",X"A6",X"A6",X"5A",X"A9",X"6A",X"A9",X"AA",
		X"56",X"AA",X"5A",X"AA",X"6A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"A9",X"AA",X"66",X"AA",X"A9",X"AA",X"65",X"AA",X"96",X"AA",X"56",X"AA",X"5A",X"AA",X"9A",
		X"AA",X"6A",X"A9",X"AA",X"A9",X"AA",X"A6",X"AA",X"9A",X"AA",X"9A",X"AA",X"6A",X"AA",X"6A",X"AA",
		X"AA",X"A9",X"AA",X"A9",X"5A",X"A6",X"AA",X"A6",X"5A",X"A6",X"66",X"9A",X"5A",X"9A",X"55",X"9A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"56",X"AA",X"5A",X"AA",X"6A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"A9",X"AA",X"66",X"AA",X"A9",X"AA",X"65",X"AA",X"96",X"AA",X"56",X"AA",X"5A",X"AA",X"9A",
		X"AA",X"6A",X"A9",X"AA",X"A9",X"AA",X"A6",X"AA",X"9A",X"AA",X"9A",X"AA",X"6A",X"AA",X"6A",X"AA",
		X"AA",X"A9",X"AA",X"A9",X"5A",X"A6",X"AA",X"A6",X"5A",X"A6",X"66",X"9A",X"5A",X"9A",X"55",X"9A",
		X"55",X"55",X"55",X"55",X"A6",X"A9",X"65",X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"55",X"55",X"55",X"55",X"AA",X"A6",X"99",X"6A",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"95",X"55",X"56",X"A5",X"6A",X"AA",X"A5",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"55",X"55",X"55",X"9A",X"AA",X"A9",X"59",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A5",X"55",X"55",X"AA",X"5A",X"55",X"A9",X"55",
		X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"FC",X"FF",X"03",X"00",X"03",X"00",X"03",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A5",X"55",X"A5",X"AA",X"A6",X"69",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A5",X"55",X"56",X"A9",X"6A",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"55",X"55",X"A5",X"65",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"55",X"55",X"69",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"A5",X"55",X"A5",X"55",X"A5",X"55",X"A5",X"55",X"AA",X"95",X"AA",X"95",
		X"AA",X"A5",X"AA",X"A5",X"AA",X"A5",X"AA",X"A5",X"AA",X"A5",X"AA",X"A5",X"AA",X"A5",X"AA",X"A5",
		X"AA",X"AA",X"AA",X"AA",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"A9",X"55",X"A9",X"55",X"A9",X"55",X"A9",X"55",X"A9",X"55",X"A9",X"5D",X"A9",X"55",X"A9",X"55",
		X"AA",X"6A",X"AA",X"AA",X"AA",X"AA",X"AA",X"EA",X"AA",X"6A",X"AA",X"E5",X"AA",X"D5",X"AA",X"95",
		X"AA",X"95",X"AA",X"95",X"AA",X"95",X"AA",X"95",X"AA",X"95",X"AA",X"95",X"AA",X"95",X"AA",X"95",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"95",X"A9",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"B5",X"AA",X"A5",X"AB",X"A5",X"AA",X"A5",X"BA",X"A5",X"AA",X"B5",
		X"AA",X"B5",X"AA",X"A5",X"AA",X"A5",X"AA",X"A5",X"AA",X"A5",X"AB",X"55",X"AA",X"55",X"AA",X"55",
		X"AA",X"55",X"AA",X"55",X"AA",X"55",X"A9",X"55",X"A9",X"55",X"A5",X"55",X"95",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A5",X"AA",X"95",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"55",X"A5",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"D5",X"A5",X"55",X"AD",X"55",X"AD",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"A5",X"55",X"A5",X"55",X"A5",X"55",X"AD",X"55",X"AE",X"AA",X"AA",X"BA",X"AA",X"AB",X"AA",X"AA",
		X"A5",X"55",X"A5",X"55",X"A5",X"55",X"A5",X"55",X"AA",X"A5",X"AA",X"A5",X"AA",X"A5",X"AA",X"A5",
		X"56",X"95",X"56",X"95",X"56",X"95",X"56",X"D5",X"56",X"95",X"57",X"95",X"D6",X"95",X"56",X"95",
		X"AA",X"AA",X"AA",X"AA",X"95",X"55",X"95",X"55",X"95",X"55",X"95",X"55",X"95",X"55",X"95",X"55",
		X"AA",X"55",X"AA",X"55",X"AA",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"57",X"55",X"55",X"55",
		X"95",X"55",X"95",X"55",X"95",X"55",X"95",X"55",X"95",X"55",X"95",X"55",X"95",X"55",X"95",X"55",
		X"A9",X"55",X"A9",X"55",X"A5",X"55",X"A5",X"55",X"95",X"55",X"95",X"55",X"55",X"55",X"55",X"55",
		X"55",X"5A",X"55",X"6A",X"55",X"6A",X"55",X"AA",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"95",X"56",X"95",X"56",X"95",X"56",X"55",X"56",X"55",X"6A",X"55",X"6E",X"55",X"7A",X"55",X"EA",
		X"55",X"55",X"FD",X"55",X"AB",X"F5",X"A9",X"55",X"A9",X"55",X"55",X"55",X"55",X"5D",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"6A",X"A5",X"FF",X"D5",X"9A",X"95",X"DA",X"A9",X"B6",X"AD",X"AE",X"BA",X"AB",X"E9",X"5E",X"B5",
		X"AA",X"A9",X"7F",X"F7",X"5A",X"96",X"9A",X"E5",X"AB",X"A9",X"AE",X"AA",X"7A",X"A9",X"FF",X"F5",
		X"AA",X"AB",X"FF",X"FD",X"56",X"A5",X"AB",X"A6",X"AB",X"EA",X"AE",X"B9",X"7A",X"AF",X"DF",X"F6",
		X"5A",X"A9",X"A7",X"FD",X"96",X"A6",X"EA",X"A7",X"7A",X"9E",X"AE",X"BA",X"AB",X"EA",X"5E",X"B5",
		X"6A",X"A9",X"FF",X"D5",X"9A",X"95",X"5A",X"A9",X"55",X"AE",X"6D",X"BA",X"AB",X"EA",X"5E",X"B5",
		X"59",X"66",X"56",X"5A",X"59",X"66",X"55",X"AA",X"56",X"66",X"56",X"AA",X"55",X"6A",X"5A",X"AA",
		X"AA",X"AA",X"9A",X"A5",X"AA",X"95",X"AA",X"99",X"9A",X"95",X"55",X"65",X"99",X"95",X"AA",X"55",
		X"55",X"56",X"55",X"55",X"57",X"55",X"5F",X"D5",X"5F",X"D5",X"57",X"55",X"55",X"56",X"9A",X"6A",
		X"55",X"FF",X"55",X"D7",X"55",X"D7",X"55",X"5F",X"55",X"5D",X"55",X"75",X"55",X"55",X"55",X"55",
		X"6A",X"9A",X"AA",X"AA",X"69",X"9A",X"AA",X"AA",X"6A",X"AA",X"5A",X"9A",X"5A",X"AA",X"55",X"9A",
		X"6A",X"AA",X"AA",X"AA",X"6A",X"AA",X"AA",X"A9",X"6A",X"AA",X"6A",X"AA",X"6A",X"AA",X"59",X"9A",
		X"55",X"55",X"55",X"55",X"95",X"66",X"9A",X"59",X"99",X"95",X"AA",X"A6",X"A9",X"99",X"AA",X"AA",
		X"55",X"55",X"57",X"75",X"55",X"55",X"55",X"55",X"FF",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"F7",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"AB",X"F7",X"B7",X"DA",X"FD",X"FF",X"AA",X"AA",
		X"FF",X"FF",X"FA",X"AA",X"FF",X"FF",X"AA",X"AE",X"AF",X"F7",X"B7",X"FA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"AA",X"AA",X"FF",X"FF",X"F7",X"FF",X"AB",X"7F",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FA",X"AA",X"FF",X"FF",X"FF",X"FF",X"AB",X"7F",X"B3",X"FA",X"AA",X"AA",X"AA",X"AA",
		X"7F",X"FF",X"AA",X"AA",X"FF",X"AB",X"F7",X"FF",X"A9",X"A7",X"AA",X"AA",X"FF",X"FA",X"AA",X"AA",
		X"FF",X"FF",X"DF",X"FF",X"7D",X"AB",X"FF",X"5F",X"FB",X"AF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"DF",X"F7",X"AB",X"E5",X"FA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"EA",X"D7",X"A5",X"7B",X"AA",X"AA",X"FF",X"FA",X"AA",X"AA",X"AB",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"77",X"FF",X"AF",X"FB",X"BF",X"5E",X"F5",X"FA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FE",X"BF",X"AA",X"FF",X"FF",X"AF",X"FB",X"AF",X"FE",X"AB",X"FA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"88",X"A8",X"00",X"80",X"00",X"80",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"0A",X"AA",X"02",X"2A",X"00",X"02",X"00",X"0A",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A2",X"A8",X"80",X"A0",X"00",X"A0",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"2A",X"AA",X"00",X"AA",X"02",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"0A",X"A8",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"2A",X"AA",X"08",X"AA",X"00",X"02",X"00",X"0A",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"22",X"A2",X"00",X"80",X"00",X"80",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"2A",X"AA",X"00",X"2A",X"00",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"8A",X"AA",X"02",X"80",X"00",X"80",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"2A",X"AA",X"00",X"2A",X"00",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A2",X"AA",X"A0",X"A8",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A2",X"AA",X"82",X"AA",X"00",X"AA",X"00",X"00",X"00",X"02",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"28",X"02",X"88",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A2",X"AA",X"22",X"AA",X"00",X"2A",X"00",X"00",X"00",X"02",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A2",X"AA",X"A0",X"82",X"A2",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"2A",X"AA",X"AA",X"AA",X"00",X"2A",X"00",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"AA",X"AA",X"00",X"00",X"A0",X"00",X"A0",X"00",
		X"3A",X"AC",X"0E",X"B0",X"83",X"C2",X"00",X"0A",X"0C",X"3A",X"30",X"0C",X"C0",X"03",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"02",X"00",X"0A",X"00",X"2A",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"AA",X"A0",X"00",X"00",X"A0",X"00",X"80",X"00",X"80",X"00",
		X"8A",X"AA",X"82",X"AA",X"82",X"AA",X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"2A",X"00",X"AA",X"02",X"AA",
		X"00",X"00",X"0C",X"0C",X"0F",X"33",X"0C",X"C3",X"C0",X"03",X"00",X"0C",X"00",X"30",X"AA",X"8A",
		X"30",X"00",X"FC",X"0C",X"FF",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FF",X"F0",X"AA",X"AA",
		X"59",X"66",X"56",X"5A",X"59",X"66",X"55",X"AA",X"56",X"66",X"56",X"AA",X"55",X"6A",X"5A",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"AA",X"A6",X"BA",X"AE",X"ED",X"F7",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"9A",X"69",X"B7",X"5E",X"F9",X"EB",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"96",X"AA",X"A9",X"AA",X"AA",X"6A",X"AA",X"96",X"AA",X"A9",X"AA",X"AA",X"AA",X"AA",
		X"55",X"55",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"6A",X"AA",X"9A",X"AA",
		X"A5",X"55",X"A9",X"55",X"A9",X"55",X"AA",X"55",X"AA",X"95",X"AA",X"A5",X"AA",X"A9",X"AA",X"A9",
		X"A6",X"AA",X"A9",X"AA",X"A9",X"AA",X"AA",X"6A",X"AA",X"9A",X"AA",X"A6",X"AA",X"A9",X"AA",X"A9",
		X"AA",X"A6",X"AA",X"A6",X"AA",X"A9",X"AA",X"A9",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"6A",X"AA",X"6A",X"AA",X"9A",X"AA",X"9A",X"AA",
		X"A6",X"AA",X"A6",X"AA",X"A9",X"AA",X"A9",X"AA",X"AA",X"6A",X"AA",X"6A",X"AA",X"9A",X"AA",X"9A",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"5A",X"AA",X"5A",X"AA",X"9A",X"AA",
		X"9A",X"AA",X"A6",X"AA",X"A6",X"AA",X"A6",X"AA",X"A6",X"AA",X"A6",X"AA",X"A6",X"AA",X"A6",X"AA",
		X"A9",X"AA",X"A9",X"AA",X"A9",X"AA",X"A9",X"AA",X"A9",X"AA",X"A9",X"AA",X"A9",X"AA",X"A9",X"AA",
		X"A9",X"AA",X"A9",X"AA",X"A9",X"AA",X"A5",X"AA",X"95",X"AA",X"95",X"AA",X"96",X"AA",X"96",X"AA",
		X"A6",X"AA",X"9A",X"AA",X"9A",X"AA",X"9A",X"AA",X"9A",X"AA",X"6A",X"AA",X"6A",X"AA",X"6A",X"AA",
		X"6A",X"AA",X"6A",X"AA",X"6A",X"AA",X"9A",X"AA",X"9A",X"AA",X"9A",X"AA",X"9A",X"AA",X"A6",X"AA",
		X"A6",X"AA",X"66",X"AA",X"A9",X"AA",X"A9",X"AA",X"A9",X"AA",X"A9",X"AA",X"A5",X"AA",X"A5",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"A9",X"FB",X"AF",X"DF",X"BF",X"BB",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"EA",X"AA",X"99",X"EB",X"FF",X"DF",X"7F",X"BF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FD",X"9B",X"BE",X"FE",
		X"FF",X"55",X"D7",X"55",X"D7",X"55",X"F5",X"55",X"75",X"55",X"5D",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"AA",X"AA",X"AA",X"AA",X"AA",X"59",X"AA",X"9A",X"AA",X"A6",X"AA",X"A9",X"AA",X"99",
		X"55",X"55",X"AA",X"AA",X"AA",X"AA",X"95",X"55",X"65",X"55",X"99",X"55",X"95",X"55",X"65",X"95",
		X"55",X"55",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"55",X"55",
		X"55",X"55",X"AA",X"96",X"AA",X"6A",X"A9",X"AA",X"96",X"AA",X"6A",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"55",X"55",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A9",X"AA",X"A6",
		X"55",X"5A",X"55",X"6A",X"55",X"6A",X"55",X"AA",X"56",X"AA",X"5A",X"AA",X"6A",X"AA",X"6A",X"AA",
		X"AA",X"9A",X"AA",X"6A",X"AA",X"6A",X"A9",X"AA",X"A6",X"AA",X"9A",X"AA",X"6A",X"AA",X"6A",X"AA",
		X"9A",X"AA",X"9A",X"AA",X"6A",X"AA",X"6A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A9",X"AA",X"A9",X"AA",X"A6",X"AA",X"A6",
		X"AA",X"9A",X"AA",X"9A",X"AA",X"6A",X"AA",X"6A",X"A9",X"AA",X"A9",X"AA",X"A6",X"AA",X"A6",X"AA",
		X"55",X"55",X"AA",X"AA",X"AA",X"AA",X"65",X"AA",X"A6",X"AA",X"9A",X"AA",X"6A",X"AA",X"66",X"AA",
		X"55",X"55",X"AA",X"AA",X"AA",X"AA",X"55",X"A6",X"55",X"99",X"99",X"66",X"66",X"56",X"66",X"9A",
		X"55",X"55",X"AA",X"AA",X"AA",X"AA",X"55",X"56",X"55",X"59",X"55",X"66",X"55",X"56",X"56",X"59",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"9A",X"AA",X"EF",X"6A",X"F7",X"FA",X"EE",X"FE",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AB",X"EB",X"66",X"F7",X"FF",X"FE",X"FD",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"E6",X"7F",X"BF",X"BE",
		X"5A",X"6A",X"69",X"AA",X"5A",X"66",X"A6",X"AA",X"99",X"AA",X"AA",X"AA",X"E6",X"7F",X"7F",X"7E",
		X"A9",X"A6",X"AA",X"69",X"AA",X"A5",X"AA",X"AA",X"AA",X"A6",X"AA",X"AA",X"B9",X"9B",X"FD",X"FD",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"77",X"5D",X"DB",X"E7",
		X"A9",X"65",X"A6",X"59",X"A9",X"96",X"9A",X"69",X"A6",X"A5",X"AA",X"65",X"A9",X"AA",X"AA",X"99",
		X"65",X"55",X"95",X"55",X"69",X"55",X"99",X"59",X"66",X"95",X"9A",X"65",X"69",X"9A",X"9A",X"95",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"D5",X"7D",X"75",X"5D",X"5D",X"55",X"57",X"55",X"55",X"55",X"5D",X"D5",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"5D",X"55",X"5D",X"D5",X"55",X"55",X"55",X"7F",X"55",X"D5",X"57",X"7D",X"5D",X"75",X"75",X"55",
		X"55",X"57",X"55",X"55",X"55",X"75",X"55",X"55",X"57",X"55",X"55",X"55",X"75",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"FC",X"0C",X"0C",X"0C",X"0C",X"30",X"0C",X"C0",X"0C",X"C0",X"0C",X"C0",X"0C",X"F0",X"0C",
		X"30",X"0C",X"30",X"0C",X"30",X"0C",X"30",X"0C",X"30",X"0C",X"30",X"0C",X"30",X"0C",X"30",X"0C",
		X"30",X"0C",X"30",X"0C",X"30",X"0C",X"30",X"0C",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"FF",X"FF",
		X"00",X"FF",X"03",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"03",X"0C",X"03",X"0C",X"03",
		X"0C",X"03",X"0C",X"03",X"0C",X"03",X"0C",X"03",X"0C",X"03",X"0C",X"03",X"0C",X"03",X"0C",X"03",
		X"0C",X"03",X"0C",X"03",X"0C",X"03",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"03",X"00",X"00",X"FF",
		X"FF",X"F0",X"00",X"0C",X"00",X"03",X"00",X"03",X"F0",X"03",X"0C",X"03",X"0C",X"03",X"0C",X"03",
		X"0C",X"03",X"0C",X"03",X"0C",X"03",X"0C",X"03",X"0C",X"03",X"0C",X"03",X"0C",X"03",X"0C",X"03",
		X"0C",X"03",X"0C",X"03",X"0C",X"03",X"F0",X"03",X"00",X"03",X"00",X"03",X"00",X"0C",X"FF",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"0D",X"00",X"35",X"00",X"D5",X"03",X"55",X"0D",X"55",
		X"35",X"55",X"D5",X"55",X"D5",X"5F",X"D5",X"55",X"3F",X"57",X"3F",X"DF",X"0F",X"FD",X"03",X"FD",
		X"00",X"FF",X"00",X"3F",X"00",X"3F",X"00",X"0F",X"00",X"03",X"00",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"0D",X"00",X"35",X"00",X"D5",X"03",X"55",X"0D",X"57",
		X"3F",X"57",X"D5",X"D7",X"F5",X"FF",X"55",X"D7",X"57",X"D7",X"5C",X"D7",X"70",X"F5",X"70",X"35",
		X"C0",X"FD",X"C0",X"D5",X"C0",X"37",X"C0",X"3D",X"C0",X"0D",X"70",X"0D",X"5F",X"3F",X"55",X"FF",
		X"55",X"7F",X"55",X"75",X"D5",X"5D",X"F5",X"5D",X"F5",X"5D",X"FD",X"5D",X"FD",X"75",X"3F",X"75",
		X"3F",X"75",X"0F",X"DF",X"0F",X"D5",X"03",X"F5",X"00",X"F7",X"00",X"F7",X"00",X"F7",X"00",X"37",
		X"00",X"35",X"00",X"35",X"00",X"35",X"00",X"35",X"00",X"35",X"00",X"35",X"00",X"D5",X"00",X"D5",
		X"00",X"D5",X"03",X"D5",X"0D",X"D7",X"35",X"7F",X"35",X"7F",X"D5",X"5F",X"D5",X"57",X"D5",X"55",
		X"35",X"55",X"35",X"55",X"0D",X"55",X"0D",X"55",X"35",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",
		X"D5",X"55",X"35",X"55",X"35",X"55",X"35",X"55",X"0D",X"55",X"0D",X"55",X"03",X"55",X"03",X"55",
		X"03",X"55",X"03",X"55",X"00",X"FF",X"03",X"FF",X"03",X"FF",X"03",X"FF",X"0F",X"FF",X"0F",X"FF",
		X"0F",X"FF",X"0F",X"FF",X"03",X"FF",X"03",X"FF",X"03",X"FF",X"03",X"FF",X"00",X"FF",X"00",X"FF",
		X"00",X"FF",X"03",X"FF",X"03",X"FF",X"03",X"FF",X"00",X"FF",X"03",X"FF",X"03",X"FF",X"00",X"FF",
		X"3F",X"C0",X"DD",X"70",X"75",X"C0",X"D7",X"C0",X"5E",X"B3",X"5E",X"AF",X"57",X"A7",X"57",X"B5",
		X"57",X"DF",X"7F",X"DD",X"D5",X"DD",X"7F",X"5F",X"D5",X"75",X"7F",X"7F",X"7F",X"57",X"55",X"57",
		X"55",X"55",X"55",X"FD",X"D7",X"57",X"DD",X"57",X"75",X"57",X"55",X"5F",X"55",X"F5",X"D7",X"5F",
		X"FD",X"7D",X"FD",X"55",X"7F",X"55",X"7F",X"FF",X"5F",X"FF",X"57",X"FF",X"55",X"FF",X"5F",X"FF",
		X"F5",X"7F",X"55",X"7F",X"55",X"7F",X"55",X"5F",X"FF",X"DF",X"00",X"D7",X"00",X"D5",X"FF",X"D5",
		X"CF",X"55",X"C3",X"57",X"C3",X"5D",X"FD",X"75",X"55",X"D5",X"5F",X"55",X"5D",X"55",X"5F",X"FF",
		X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FF",X"FC",
		X"55",X"5C",X"55",X"5C",X"55",X"5C",X"55",X"5C",X"FD",X"5C",X"75",X"57",X"75",X"57",X"75",X"57",
		X"75",X"57",X"75",X"55",X"75",X"55",X"75",X"55",X"D5",X"55",X"F5",X"55",X"CD",X"55",X"C3",X"55",
		X"C3",X"55",X"C0",X"D5",X"C0",X"D5",X"C0",X"FF",X"C3",X"FF",X"C3",X"FF",X"CF",X"FF",X"CF",X"FF",
		X"CF",X"FF",X"C3",X"FF",X"C3",X"FF",X"03",X"FF",X"03",X"FC",X"03",X"FC",X"03",X"FC",X"03",X"FC",
		X"03",X"FC",X"03",X"FF",X"C3",X"FF",X"CF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"AC",X"00",X"AC",X"00",X"EC",X"00",
		X"70",X"00",X"F0",X"00",X"5C",X"00",X"D7",X"00",X"77",X"00",X"DC",X"00",X"DC",X"00",X"5C",X"00",
		X"D7",X"00",X"D7",X"00",X"D7",X"00",X"7C",X"00",X"5F",X"00",X"57",X"00",X"D7",X"00",X"77",X"00",
		X"FC",X"00",X"C0",X"00",X"F0",X"00",X"FF",X"C0",X"FD",X"70",X"FF",X"5C",X"FF",X"57",X"FF",X"57",
		X"FF",X"D7",X"FF",X"DC",X"FF",X"DC",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",
		X"FF",X"D7",X"FF",X"D7",X"FF",X"DC",X"FF",X"DC",X"FD",X"5C",X"7D",X"5C",X"55",X"70",X"55",X"C0",
		X"FF",X"C0",X"FD",X"C0",X"F5",X"C0",X"F5",X"C0",X"F5",X"C0",X"FF",X"00",X"F7",X"00",X"F7",X"00",
		X"FD",X"F0",X"D5",X"5C",X"D5",X"57",X"D7",X"D7",X"DD",X"17",X"D7",X"37",X"37",X"DC",X"37",X"30",
		X"37",X"C0",X"CF",X"C0",X"CF",X"C0",X"7F",X"C0",X"7F",X"C0",X"5F",X"C0",X"5F",X"C0",X"5F",X"C0",
		X"5F",X"C0",X"5F",X"C0",X"7F",X"C0",X"CF",X"C0",X"CF",X"C0",X"CF",X"C0",X"CF",X"C0",X"CF",X"C0",
		X"0F",X"C0",X"0F",X"C0",X"0F",X"C0",X"0F",X"C0",X"0F",X"C0",X"0F",X"C0",X"0F",X"C0",X"0F",X"C0",
		X"0F",X"C0",X"0F",X"C0",X"CF",X"C0",X"FF",X"C0",X"FF",X"C0",X"FF",X"F0",X"FF",X"F0",X"FF",X"C0",
		X"00",X"03",X"00",X"03",X"00",X"0D",X"00",X"35",X"00",X"37",X"00",X"35",X"00",X"3D",X"00",X"D7",
		X"00",X"DD",X"03",X"57",X"03",X"75",X"00",X"F5",X"00",X"0F",X"00",X"03",X"03",X"FF",X"0D",X"7F",
		X"0D",X"FF",X"0D",X"FD",X"03",X"FD",X"0D",X"FD",X"35",X"FD",X"37",X"FD",X"37",X"FD",X"37",X"FD",
		X"37",X"FD",X"37",X"FD",X"37",X"FD",X"3B",X"FE",X"0F",X"FE",X"0F",X"FE",X"03",X"FE",X"03",X"FE",
		X"03",X"FD",X"03",X"FF",X"03",X"FC",X"03",X"FC",X"00",X"FC",X"00",X"F0",X"00",X"00",X"00",X"03",
		X"00",X"D0",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"0F",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"3C",X"00",X"EB",X"3F",X"EB",X"EA",X"FF",X"EA",X"FF",X"7F",X"FF",X"57",X"D7",X"55",X"55",X"D5",
		X"D5",X"75",X"FD",X"ED",X"F5",X"FF",X"D5",X"FD",X"55",X"55",X"F5",X"57",X"55",X"57",X"57",X"55",
		X"FD",X"55",X"55",X"5F",X"55",X"5C",X"7F",X"FF",X"FF",X"FD",X"FF",X"F5",X"FF",X"D5",X"FF",X"55",
		X"55",X"55",X"55",X"55",X"5F",X"FD",X"5C",X"0D",X"5C",X"0D",X"5F",X"FD",X"7F",X"D5",X"7F",X"D5",
		X"7F",X"D5",X"5F",X"55",X"55",X"55",X"95",X"55",X"95",X"55",X"A5",X"55",X"A9",X"55",X"AA",X"55",
		X"AA",X"5F",X"FF",X"FF",X"F0",X"FF",X"F0",X"FF",X"FF",X"F5",X"D5",X"55",X"DD",X"55",X"5D",X"55",
		X"5D",X"55",X"5D",X"55",X"FD",X"55",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",
		X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"0F",X"FF",X"03",X"FF",
		X"0F",X"FF",X"0F",X"FF",X"0F",X"FF",X"0F",X"FF",X"0F",X"FF",X"0F",X"FF",X"0F",X"FF",X"0F",X"FF",
		X"03",X"FF",X"03",X"FF",X"03",X"FF",X"03",X"FF",X"03",X"FF",X"03",X"FF",X"03",X"FF",X"03",X"FF",
		X"0F",X"FF",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"3F",X"C0",X"0F",
		X"00",X"00",X"00",X"00",X"3C",X"00",X"C3",X"F0",X"F0",X"C0",X"C3",X"00",X"C0",X"F0",X"70",X"0C",
		X"5C",X"0C",X"57",X"FC",X"5D",X"5F",X"FA",X"55",X"CE",X"95",X"03",X"A5",X"00",X"E9",X"C3",X"3A",
		X"CC",X"0F",X"0C",X"3A",X"3C",X"F9",X"D7",X"E5",X"5D",X"55",X"75",X"56",X"55",X"5A",X"55",X"6A",
		X"55",X"6A",X"55",X"AB",X"56",X"AC",X"5A",X"B0",X"6A",X"B0",X"6A",X"C0",X"6B",X"00",X"6C",X"00",
		X"70",X"00",X"70",X"00",X"70",X"00",X"70",X"00",X"70",X"00",X"7C",X"00",X"7F",X"00",X"FF",X"00",
		X"FF",X"00",X"F5",X"C0",X"D5",X"70",X"55",X"5C",X"55",X"5C",X"55",X"57",X"55",X"57",X"55",X"57",
		X"55",X"57",X"55",X"FC",X"7F",X"C0",X"FF",X"C0",X"FF",X"C0",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FC",X"00",X"FC",X"00",X"FC",X"00",X"FC",X"00",
		X"FC",X"00",X"FC",X"00",X"FC",X"00",X"FC",X"00",X"FC",X"00",X"FC",X"00",X"F0",X"00",X"C0",X"00",
		X"F0",X"00",X"F0",X"00",X"FC",X"00",X"FC",X"00",X"FC",X"00",X"FC",X"00",X"FC",X"00",X"FC",X"00",
		X"FC",X"00",X"FC",X"00",X"FC",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",
		X"F0",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"FC",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"70",X"00",X"5F",X"00",X"55",X"C0",X"55",X"70",
		X"55",X"AC",X"56",X"B0",X"5A",X"C0",X"6A",X"C0",X"AB",X"00",X"AC",X"00",X"B0",X"00",X"B0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"35",X"00",X"35",
		X"00",X"35",X"00",X"35",X"00",X"35",X"00",X"35",X"00",X"35",X"00",X"35",X"00",X"35",X"00",X"35",
		X"00",X"35",X"00",X"35",X"00",X"35",X"00",X"35",X"00",X"35",X"00",X"35",X"00",X"35",X"F0",X"35",
		X"EC",X"35",X"EC",X"3D",X"3B",X"37",X"0E",X"F5",X"0E",X"B5",X"03",X"DF",X"03",X"55",X"03",X"57",
		X"03",X"5C",X"03",X"5C",X"00",X"D7",X"00",X"35",X"00",X"0D",X"00",X"03",X"00",X"00",X"00",X"00",
		X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"0F",X"00",X"3F",X"00",X"FF",X"00",X"FF",
		X"AB",X"FF",X"AB",X"FF",X"BB",X"FF",X"AA",X"FF",X"AA",X"AF",X"FE",X"AF",X"AA",X"FE",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"3B",X"00",X"EA",X"03",X"6A",X"03",X"7F",X"03",X"D5",
		X"35",X"FF",X"D7",X"5D",X"5D",X"57",X"57",X"D5",X"5D",X"7D",X"57",X"7F",X"57",X"5F",X"57",X"55",
		X"57",X"5F",X"5D",X"75",X"77",X"D5",X"75",X"57",X"5D",X"5F",X"57",X"F7",X"55",X"75",X"55",X"75",
		X"5D",X"5F",X"5D",X"55",X"5D",X"55",X"73",X"55",X"73",X"5F",X"73",X"5D",X"70",X"DD",X"70",X"DD",
		X"70",X"DD",X"70",X"DD",X"70",X"FD",X"70",X"DF",X"70",X"D5",X"73",X"55",X"73",X"55",X"73",X"55",
		X"73",X"57",X"7D",X"55",X"7D",X"55",X"75",X"55",X"75",X"55",X"DD",X"55",X"57",X"55",X"D7",X"55",
		X"37",X"55",X"37",X"55",X"DD",X"55",X"75",X"55",X"F5",X"55",X"35",X"55",X"0D",X"55",X"0D",X"55",
		X"03",X"55",X"0F",X"FF",X"3F",X"FF",X"3F",X"FF",X"FF",X"FC",X"FF",X"FC",X"FF",X"F0",X"FF",X"F0",
		X"FF",X"C0",X"FF",X"C0",X"FF",X"00",X"FF",X"00",X"FC",X"00",X"FC",X"00",X"FC",X"00",X"F0",X"00",
		X"FA",X"AA",X"FF",X"FF",X"FF",X"AF",X"FF",X"FA",X"FF",X"FA",X"FF",X"FA",X"FF",X"EA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"F0",X"FE",X"AC",X"DE",X"AC",X"F7",X"EC",X"F5",X"70",
		X"5F",X"FF",X"57",X"55",X"FD",X"57",X"75",X"7F",X"75",X"F5",X"5F",X"F7",X"57",X"F7",X"55",X"57",
		X"DF",X"D7",X"DD",X"75",X"75",X"5F",X"FF",X"55",X"F0",X"D5",X"FF",X"7F",X"55",X"5D",X"55",X"5D",
		X"55",X"F5",X"FF",X"55",X"5D",X"55",X"F5",X"55",X"55",X"55",X"D5",X"D5",X"55",X"57",X"55",X"57",
		X"D5",X"D7",X"55",X"57",X"55",X"5F",X"FF",X"F7",X"55",X"57",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"55",X"75",X"55",X"75",X"55",X"75",X"55",X"75",X"55",X"75",X"55",X"75",X"57",X"75",X"57",
		X"75",X"57",X"75",X"57",X"75",X"55",X"75",X"55",X"75",X"55",X"75",X"55",X"75",X"55",X"75",X"55",
		X"75",X"57",X"CF",X"FF",X"0F",X"FF",X"0F",X"FF",X"03",X"FF",X"03",X"FF",X"00",X"FF",X"00",X"FF",
		X"00",X"3F",X"00",X"3F",X"00",X"0F",X"00",X"0F",X"00",X"03",X"00",X"03",X"00",X"00",X"00",X"00",
		X"AA",X"AB",X"AF",X"FA",X"AA",X"AA",X"BE",X"BF",X"AA",X"FF",X"AA",X"FF",X"AA",X"BF",X"AA",X"AA",
		X"00",X"00",X"F0",X"00",X"5C",X"00",X"57",X"00",X"D5",X"C0",X"55",X"C0",X"55",X"70",X"55",X"70",
		X"55",X"70",X"D5",X"70",X"75",X"70",X"75",X"70",X"D5",X"70",X"55",X"70",X"55",X"70",X"55",X"70",
		X"D5",X"70",X"D5",X"70",X"D5",X"70",X"D5",X"70",X"F5",X"70",X"35",X"70",X"35",X"70",X"35",X"70",
		X"35",X"70",X"35",X"70",X"35",X"70",X"35",X"70",X"35",X"70",X"35",X"70",X"F5",X"70",X"F5",X"70",
		X"F5",X"70",X"75",X"70",X"77",X"F0",X"75",X"70",X"75",X"70",X"DF",X"F0",X"55",X"70",X"55",X"70",
		X"5D",X"70",X"FD",X"70",X"D5",X"70",X"D7",X"C0",X"FC",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",
		X"00",X"00",X"C0",X"00",X"C0",X"00",X"F0",X"00",X"FC",X"00",X"FC",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"C0",X"FF",X"C0",X"FF",X"F0",X"FF",X"F0",X"FF",X"FC",X"3F",X"FF",
		X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"AA",X"FF",X"BE",X"FE",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"F0",X"0F",X"00",X"F0",X"00",
		X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"03",X"C3",X"03",X"FF",X"03",X"03",X"03",X"03",X"03",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"FF",
		X"00",X"0F",X"00",X"F3",X"0C",X"C3",X"FC",X"C3",X"0C",X"C3",X"0C",X"C3",X"0C",X"C3",X"0C",X"C0",
		X"0C",X"30",X"0C",X"30",X"3C",X"30",X"C0",X"30",X"00",X"30",X"00",X"30",X"00",X"30",X"00",X"30",
		X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",
		X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"FC",X"0F",X"0C",X"0C",X"0C",
		X"0C",X"03",X"0C",X"03",X"0C",X"03",X"0C",X"03",X"0C",X"03",X"0C",X"03",X"0C",X"03",X"0C",X"03",
		X"CC",X"03",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"F0",X"30",X"F0",X"30",X"30",X"30",
		X"30",X"30",X"30",X"30",X"00",X"30",X"00",X"30",X"00",X"CC",X"00",X"CC",X"00",X"CC",X"00",X"CC",
		X"03",X"0C",X"03",X"0C",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"FF",X"03",
		X"00",X"0C",X"00",X"FC",X"0F",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",
		X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"30",X"0C",X"30",X"0C",X"30",X"0C",X"30",X"0C",X"30",X"30",
		X"30",X"30",X"F0",X"30",X"F0",X"30",X"F0",X"30",X"C0",X"30",X"C0",X"30",X"C0",X"30",X"C0",X"30",
		X"00",X"30",X"00",X"30",X"00",X"30",X"00",X"30",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",
		X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"FF",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"3C",X"03",X"C0",X"0C",X"00",X"30",X"00",
		X"30",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"0F",
		X"C0",X"30",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"3F",X"C0",X"00",X"C0",X"00",X"C0",X"00",
		X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"30",X"00",X"0F",X"FF",
		X"00",X"00",X"03",X"F0",X"3C",X"0C",X"C0",X"0C",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",
		X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",
		X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",
		X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"0C",X"00",X"0C",X"00",X"30",X"FF",X"C0",
		X"FC",X"00",X"C3",X"F0",X"C0",X"0F",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",
		X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"FC",X"00",X"03",X"FC",X"00",X"0C",X"00",X"0C",
		X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",
		X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0F",
		X"00",X"00",X"00",X"00",X"C0",X"00",X"3F",X"00",X"00",X"FC",X"00",X"03",X"00",X"03",X"00",X"03",
		X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"03",X"C3",
		X"03",X"3F",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",
		X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",
		X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"00",X"30",X"FC",
		X"30",X"0C",X"30",X"0C",X"30",X"0C",X"30",X"0C",X"30",X"0C",X"30",X"0C",X"30",X"0C",X"30",X"0C",
		X"30",X"0C",X"30",X"0C",X"30",X"0C",X"30",X"0C",X"30",X"0C",X"30",X"0C",X"30",X"0C",X"3F",X"FC",
		X"00",X"00",X"0F",X"00",X"30",X"F0",X"C0",X"0F",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",
		X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"C0",X"C3",X"30",X"C3",X"0C",X"C3",X"0C",X"C3",X"0F",
		X"C3",X"00",X"C3",X"3C",X"C3",X"33",X"C3",X"30",X"C3",X"30",X"C3",X"30",X"C3",X"30",X"C3",X"30",
		X"C3",X"30",X"C3",X"3C",X"C3",X"0C",X"C3",X"0C",X"C3",X"0C",X"C3",X"0C",X"C0",X"F0",X"C0",X"00",
		X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"0F",X"30",X"33",X"0F",X"C3",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"33",X"FC",X"33",X"03",X"33",X"00",
		X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"0F",
		X"F3",X"0C",X"03",X"0C",X"C3",X"0C",X"33",X"0C",X"33",X"0F",X"33",X"00",X"33",X"00",X"33",X"00",
		X"33",X"00",X"33",X"0F",X"33",X"0C",X"33",X"0C",X"33",X"0C",X"33",X"0C",X"33",X"0C",X"33",X"0C",
		X"33",X"0F",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"F3",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"0F",X"00",
		X"03",X"3F",X"03",X"30",X"03",X"30",X"03",X"30",X"03",X"30",X"03",X"30",X"03",X"30",X"F3",X"30",
		X"0F",X"30",X"00",X"30",X"00",X"30",X"00",X"30",X"FF",X"30",X"03",X"30",X"03",X"30",X"03",X"30",
		X"03",X"30",X"03",X"30",X"FF",X"30",X"00",X"30",X"00",X"30",X"00",X"30",X"00",X"30",X"00",X"30",
		X"FF",X"30",X"03",X"30",X"03",X"30",X"03",X"30",X"03",X"30",X"03",X"30",X"03",X"30",X"FF",X"3F",
		X"00",X"00",X"F0",X"00",X"0C",X"00",X"03",X"00",X"00",X"C0",X"00",X"C3",X"00",X"3C",X"00",X"3C",
		X"00",X"3C",X"F0",X"3C",X"CC",X"3C",X"CC",X"3C",X"CC",X"3C",X"F0",X"3C",X"00",X"3C",X"00",X"3C",
		X"00",X"CC",X"03",X"0C",X"00",X"CC",X"F0",X"33",X"CC",X"30",X"CC",X"30",X"CC",X"3F",X"CC",X"3C",
		X"CC",X"3C",X"CC",X"3C",X"CC",X"3C",X"CC",X"3C",X"CC",X"3C",X"CC",X"33",X"CC",X"33",X"CC",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"00",X"03",X"F0",X"00",X"0C",X"00",X"03",
		X"00",X"03",X"00",X"03",X"00",X"03",X"0F",X"03",X"30",X"C3",X"30",X"FF",X"30",X"00",X"0C",X"00",
		X"03",X"FC",X"00",X"03",X"00",X"03",X"C0",X"03",X"3F",X"03",X"00",X"C3",X"F0",X"C3",X"30",X"C3",
		X"0F",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"0C",X"00",X"0C",X"FF",X"F0",
		X"A8",X"00",X"AA",X"80",X"AA",X"E0",X"AA",X"A8",X"AA",X"AE",X"AA",X"A8",X"A8",X"00",X"AA",X"80",
		X"AA",X"80",X"A8",X"00",X"AA",X"A8",X"AA",X"AE",X"AA",X"A8",X"AA",X"E0",X"AA",X"80",X"A8",X"00",
		X"02",X"AA",X"00",X"2A",X"2A",X"AA",X"BA",X"AA",X"2A",X"AA",X"0B",X"AA",X"02",X"AA",X"00",X"2A",
		X"00",X"2A",X"0A",X"AA",X"2B",X"AA",X"AA",X"AA",X"BA",X"AA",X"2A",X"AA",X"0A",X"AA",X"02",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"3C",X"0F",X"C0",
		X"30",X"00",X"30",X"0F",X"33",X"F5",X"3D",X"57",X"35",X"5C",X"CF",X"F0",X"C0",X"CF",X"3F",X"75",
		X"3F",X"DF",X"37",X"5F",X"37",X"55",X"0D",X"55",X"0F",X"D5",X"0D",X"55",X"37",X"FF",X"35",X"7F",
		X"DD",X"7F",X"D5",X"5F",X"DD",X"55",X"35",X"5F",X"0F",X"F0",X"00",X"00",X"0C",X"00",X"37",X"00",
		X"35",X"C0",X"D7",X"70",X"D5",X"70",X"D5",X"F3",X"D7",X"5D",X"D7",X"5D",X"3E",X"9D",X"0E",X"95",
		X"03",X"A9",X"00",X"EA",X"00",X"3A",X"00",X"0E",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"0F",X"00",X"0F",X"00",X"3F",X"00",X"3F",
		X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",
		X"AA",X"AA",X"AA",X"AF",X"AA",X"BF",X"AA",X"BF",X"AA",X"AF",X"AA",X"AB",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"33",X"F0",X"3C",X"30",
		X"00",X"30",X"C0",X"0C",X"70",X"0C",X"5C",X"0C",X"D7",X"03",X"37",X"0C",X"D7",X"0C",X"57",X"03",
		X"DC",X"00",X"D7",X"00",X"55",X"C0",X"55",X"C0",X"55",X"C3",X"55",X"7E",X"55",X"EB",X"D5",X"ED",
		X"D7",X"F5",X"57",X"55",X"5D",X"55",X"F5",X"55",X"35",X"55",X"35",X"55",X"0D",X"55",X"0D",X"55",
		X"35",X"55",X"35",X"55",X"D5",X"55",X"D5",X"5E",X"D5",X"7A",X"D5",X"FA",X"57",X"0E",X"57",X"03",
		X"5C",X"03",X"5C",X"03",X"70",X"03",X"C0",X"03",X"00",X"0E",X"00",X"0E",X"00",X"3F",X"00",X"FF",
		X"0F",X"FF",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CF",X"FF",X"C3",
		X"FF",X"C0",X"FF",X"C0",X"FF",X"C0",X"FF",X"C0",X"FF",X"F0",X"3F",X"F0",X"3F",X"F0",X"3F",X"F0",
		X"FF",X"FA",X"FF",X"FA",X"FF",X"FA",X"FF",X"FA",X"FF",X"FA",X"FF",X"FA",X"AF",X"EA",X"AA",X"AA",
		X"C0",X"00",X"C0",X"00",X"C0",X"3C",X"C3",X"D7",X"3D",X"55",X"D5",X"55",X"55",X"55",X"55",X"57",
		X"55",X"57",X"55",X"57",X"55",X"57",X"55",X"57",X"55",X"57",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"95",X"55",X"95",X"55",X"A5",X"55",X"A5",X"55",X"A5",X"55",X"A5",X"5F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"99",X"55",X"A5",X"55",X"A5",X"55",X"A5",X"55",X"E5",X"55",
		X"E9",X"55",X"FD",X"55",X"FF",X"55",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FF",X"F0",
		X"FF",X"C0",X"FF",X"00",X"FF",X"00",X"FF",X"C0",X"FF",X"C0",X"FF",X"F0",X"FF",X"FC",X"FF",X"FC",
		X"FF",X"FF",X"3F",X"FF",X"0F",X"FF",X"0F",X"FF",X"03",X"FF",X"00",X"FF",X"00",X"3F",X"00",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"7C",X"00",X"57",X"C0",X"55",X"70",
		X"A5",X"5C",X"A9",X"5B",X"EF",X"6B",X"35",X"AC",X"3E",X"AC",X"EA",X"B0",X"EA",X"B0",X"EA",X"C0",
		X"EB",X"00",X"EB",X"00",X"7C",X"00",X"70",X"00",X"70",X"00",X"70",X"00",X"F0",X"00",X"F0",X"00",
		X"70",X"00",X"DC",X"00",X"57",X"00",X"57",X"00",X"75",X"C0",X"75",X"C0",X"7D",X"70",X"7D",X"70",
		X"7D",X"70",X"FD",X"C0",X"FF",X"00",X"F0",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"C0",X"00",X"F0",X"00",X"FC",X"00",X"FC",X"00",
		X"FF",X"AA",X"FF",X"AA",X"FF",X"AA",X"FF",X"AA",X"FF",X"AA",X"FF",X"AA",X"FE",X"AA",X"AA",X"AA",
		X"6E",X"4A",X"FE",X"7A",X"01",X"C5",X"61",X"45",X"31",X"25",X"EA",X"49",X"2E",X"F9",X"75",X"FB",
		X"4D",X"C9",X"3B",X"39",X"27",X"7E",X"1C",X"3F",X"CC",X"7B",X"6E",X"49",X"FB",X"E5",X"49",X"A1",
		X"26",X"25",X"3B",X"B7",X"35",X"C9",X"1E",X"D9",X"47",X"69",X"2E",X"DE",X"0E",X"F8",X"FB",X"2B",
		X"C6",X"45",X"26",X"21",X"29",X"FB",X"4E",X"1E",X"44",X"B5",X"CE",X"42",X"6E",X"F9",X"09",X"19",
		X"22",X"71",X"45",X"36",X"D8",X"A9",X"2A",X"09",X"7A",X"E1",X"E9",X"29",X"EE",X"0E",X"D2",X"FB",
		X"02",X"39",X"49",X"C8",X"2F",X"75",X"28",X"CD",X"7E",X"F8",X"E6",X"F8",X"BD",X"6A",X"CD",X"F1",
		X"7A",X"E9",X"06",X"F8",X"B9",X"B5",X"08",X"9D",X"0C",X"74",X"69",X"09",X"21",X"4F",X"09",X"34",
		X"FE",X"3A",X"E7",X"11",X"E1",X"5A",X"48",X"FD",X"E2",X"38",X"66",X"21",X"E5",X"FA",X"FB",X"DD",
		X"C9",X"07",X"0B",X"85",X"66",X"D9",X"7A",X"F9",X"C5",X"4A",X"62",X"F8",X"0E",X"31",X"E5",X"0A",
		X"35",X"03",X"26",X"E9",X"47",X"C9",X"39",X"39",X"ED",X"C2",X"01",X"F0",X"EC",X"DA",X"6C",X"41",
		X"ED",X"03",X"2A",X"A7",X"65",X"99",X"39",X"F9",X"C8",X"C9",X"06",X"B9",X"66",X"BA",X"2F",X"F8",
		X"E1",X"07",X"47",X"BB",X"C6",X"89",X"6A",X"99",X"68",X"E1",X"E3",X"F3",X"A6",X"11",X"A5",X"79",
		X"F9",X"CD",X"16",X"C5",X"3C",X"18",X"69",X"3B",X"EA",X"D9",X"F8",X"0A",X"05",X"F1",X"E6",X"15",
		X"7E",X"00",X"78",X"39",X"09",X"3B",X"4D",X"C9",X"02",X"E9",X"39",X"BB",X"C6",X"F4",X"AE",X"C9",
		X"4B",X"2B",X"B9",X"3A",X"7E",X"F9",X"86",X"F1",X"FA",X"83",X"34",X"01",X"6A",X"79",X"EC",X"FD",
		X"6D",X"E7",X"67",X"FB",X"6E",X"29",X"F9",X"2D",X"75",X"37",X"33",X"4B",X"3F",X"D1",X"22",X"39");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
