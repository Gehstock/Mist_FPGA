library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity spr_rom is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of spr_rom is
	type rom is array(0 to  32767) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"22",X"22",X"22",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"02",X"22",X"22",X"53",X"8C",X"00",X"00",X"00",X"00",X"00",X"FF",X"22",X"2D",X"E2",X"C3",
		X"85",X"50",X"00",X"00",X"00",X"00",X"FF",X"22",X"2D",X"E2",X"55",X"53",X"33",X"00",X"00",X"00",
		X"00",X"FF",X"22",X"22",X"22",X"53",X"35",X"55",X"55",X"50",X"00",X"00",X"FF",X"22",X"22",X"22",
		X"25",X"55",X"25",X"BB",X"55",X"50",X"00",X"FF",X"22",X"22",X"23",X"35",X"55",X"55",X"7B",X"B5",
		X"C5",X"00",X"FF",X"02",X"22",X"33",X"35",X"55",X"25",X"17",X"B5",X"CC",X"50",X"FF",X"00",X"22",
		X"33",X"35",X"55",X"55",X"77",X"B5",X"C6",X"C5",X"FF",X"00",X"00",X"33",X"35",X"55",X"25",X"77",
		X"B5",X"C1",X"65",X"FF",X"00",X"00",X"33",X"25",X"55",X"55",X"17",X"55",X"C1",X"65",X"FF",X"00",
		X"00",X"33",X"22",X"35",X"55",X"55",X"55",X"C6",X"65",X"FF",X"00",X"00",X"32",X"55",X"53",X"55",
		X"55",X"5C",X"C1",X"C5",X"FF",X"00",X"22",X"22",X"53",X"85",X"35",X"55",X"55",X"CC",X"C5",X"FF",
		X"02",X"22",X"22",X"53",X"85",X"53",X"55",X"55",X"5C",X"50",X"FF",X"22",X"2D",X"E2",X"55",X"CC",
		X"53",X"55",X"77",X"55",X"50",X"FF",X"22",X"2D",X"E2",X"25",X"CC",X"C3",X"45",X"B7",X"B5",X"00",
		X"FF",X"22",X"22",X"22",X"22",X"5C",X"C2",X"34",X"5B",X"50",X"00",X"FF",X"22",X"22",X"22",X"22",
		X"25",X"C2",X"23",X"35",X"00",X"00",X"FF",X"22",X"22",X"22",X"22",X"25",X"35",X"55",X"33",X"27",
		X"00",X"FF",X"02",X"B9",X"99",X"B2",X"52",X"5C",X"CC",X"55",X"71",X"00",X"FF",X"00",X"BB",X"BB",
		X"B2",X"22",X"55",X"5C",X"C5",X"27",X"00",X"FF",X"00",X"00",X"00",X"02",X"22",X"22",X"25",X"C5",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"02",X"22",X"22",X"22",X"50",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"02",X"2B",X"99",X"B2",X"20",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"2B",X"BB",X"B2",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"25",X"83",X"50",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"02",X"25",X"83",X"CC",X"A0",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"22",X"25",X"CC",X"C5",X"30",X"00",X"00",X"00",X"00",X"00",X"FF",X"22",X"25",X"55",X"33",X"55",
		X"55",X"53",X"3C",X"C0",X"00",X"FF",X"22",X"25",X"53",X"55",X"55",X"B5",X"55",X"53",X"CC",X"00",
		X"FF",X"22",X"22",X"25",X"52",X"5B",X"BB",X"55",X"55",X"3C",X"00",X"FF",X"22",X"22",X"55",X"55",
		X"5B",X"77",X"55",X"C6",X"5C",X"00",X"FF",X"02",X"23",X"55",X"52",X"5B",X"17",X"55",X"C1",X"C5",
		X"00",X"FF",X"00",X"23",X"55",X"55",X"5B",X"71",X"55",X"C1",X"15",X"27",X"FF",X"00",X"03",X"55",
		X"52",X"5B",X"17",X"55",X"C6",X"15",X"71",X"FF",X"00",X"03",X"55",X"55",X"55",X"75",X"55",X"C6",
		X"C5",X"27",X"FF",X"00",X"03",X"55",X"55",X"55",X"55",X"55",X"5C",X"55",X"00",X"FF",X"00",X"02",
		X"25",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"FF",X"00",X"23",X"33",X"35",X"55",X"55",X"55",
		X"55",X"55",X"00",X"FF",X"02",X"25",X"55",X"53",X"33",X"55",X"77",X"B5",X"50",X"27",X"FF",X"22",
		X"25",X"83",X"CC",X"52",X"55",X"55",X"55",X"32",X"71",X"FF",X"22",X"25",X"83",X"CC",X"C2",X"22",
		X"33",X"33",X"30",X"27",X"FF",X"22",X"25",X"55",X"5C",X"C5",X"23",X"55",X"55",X"55",X"00",X"FF",
		X"22",X"22",X"55",X"55",X"55",X"25",X"5C",X"CC",X"CC",X"00",X"FF",X"22",X"22",X"22",X"22",X"25",
		X"25",X"5C",X"CC",X"CC",X"00",X"FF",X"02",X"B9",X"99",X"B2",X"00",X"22",X"22",X"22",X"2C",X"00",
		X"FF",X"00",X"BB",X"BB",X"B0",X"00",X"22",X"B9",X"9B",X"22",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"02",X"BB",X"BB",X"20",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"22",X"22",
		X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"02",X"22",X"22",X"53",X"80",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"22",X"2D",X"E2",X"C3",X"8C",X"00",X"00",X"00",X"00",X"00",X"FF",X"22",X"2D",
		X"E2",X"C5",X"55",X"50",X"00",X"00",X"00",X"00",X"FF",X"22",X"22",X"22",X"55",X"33",X"35",X"00",
		X"00",X"00",X"00",X"FF",X"22",X"22",X"22",X"33",X"35",X"55",X"55",X"00",X"00",X"00",X"FF",X"22",
		X"22",X"22",X"25",X"55",X"C5",X"55",X"5C",X"00",X"00",X"FF",X"02",X"22",X"32",X"55",X"5C",X"CC",
		X"25",X"55",X"C0",X"00",X"FF",X"00",X"23",X"32",X"55",X"CC",X"CC",X"55",X"BB",X"5C",X"00",X"FF",
		X"00",X"03",X"32",X"55",X"CC",X"CC",X"25",X"1B",X"BC",X"C0",X"FF",X"00",X"03",X"32",X"55",X"5C",
		X"CC",X"55",X"71",X"BC",X"C0",X"FF",X"00",X"03",X"32",X"33",X"55",X"C5",X"25",X"17",X"BC",X"C0",
		X"FF",X"00",X"03",X"32",X"55",X"35",X"55",X"55",X"71",X"5C",X"C0",X"FF",X"00",X"22",X"22",X"53",
		X"83",X"55",X"55",X"55",X"5C",X"C0",X"FF",X"02",X"22",X"22",X"53",X"85",X"35",X"55",X"55",X"CC",
		X"C0",X"FF",X"22",X"2D",X"E2",X"55",X"CC",X"35",X"55",X"55",X"5C",X"C0",X"FF",X"22",X"2D",X"E2",
		X"25",X"5C",X"35",X"55",X"17",X"BC",X"00",X"FF",X"22",X"22",X"22",X"22",X"5C",X"35",X"55",X"77",
		X"BC",X"00",X"FF",X"22",X"22",X"22",X"22",X"5C",X"35",X"55",X"BB",X"C0",X"00",X"FF",X"22",X"22",
		X"22",X"22",X"5C",X"23",X"55",X"5C",X"00",X"00",X"FF",X"02",X"B9",X"99",X"B2",X"C2",X"33",X"55",
		X"00",X"00",X"00",X"FF",X"00",X"BB",X"BB",X"BC",X"C2",X"53",X"70",X"00",X"00",X"00",X"FF",X"00",
		X"02",X"22",X"55",X"55",X"55",X"10",X"00",X"00",X"00",X"FF",X"00",X"02",X"22",X"22",X"25",X"55",
		X"70",X"00",X"00",X"00",X"FF",X"00",X"02",X"22",X"22",X"22",X"25",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"02",X"2B",X"99",X"B2",X"20",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"2B",X"BB",X"B2",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"22",X"22",X"25",X"71",X"70",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"02",X"22",X"22",X"25",X"71",X"7C",X"A0",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"22",X"21",X"22",X"25",X"C7",X"C5",X"30",X"00",X"00",X"00",X"00",X"00",X"FF",X"22",
		X"21",X"22",X"25",X"55",X"33",X"55",X"55",X"53",X"3C",X"C0",X"00",X"FF",X"22",X"22",X"22",X"25",
		X"53",X"55",X"55",X"B5",X"55",X"53",X"CC",X"00",X"FF",X"22",X"22",X"22",X"22",X"25",X"52",X"5B",
		X"BB",X"55",X"55",X"3C",X"00",X"FF",X"22",X"22",X"22",X"22",X"55",X"55",X"5B",X"77",X"55",X"C6",
		X"5C",X"00",X"FF",X"02",X"BB",X"BB",X"B3",X"55",X"52",X"5B",X"17",X"55",X"C1",X"C5",X"00",X"FF",
		X"00",X"BB",X"BB",X"B3",X"55",X"55",X"5B",X"71",X"55",X"C1",X"15",X"27",X"FF",X"00",X"00",X"00",
		X"03",X"55",X"52",X"5B",X"17",X"55",X"C6",X"15",X"71",X"FF",X"00",X"00",X"00",X"03",X"55",X"55",
		X"55",X"75",X"55",X"C6",X"C5",X"27",X"FF",X"00",X"00",X"00",X"03",X"55",X"55",X"55",X"55",X"55",
		X"5C",X"55",X"00",X"FF",X"00",X"00",X"00",X"02",X"25",X"55",X"55",X"55",X"55",X"55",X"55",X"00",
		X"FF",X"00",X"22",X"22",X"23",X"33",X"35",X"55",X"55",X"55",X"55",X"55",X"00",X"FF",X"02",X"22",
		X"22",X"25",X"57",X"53",X"33",X"55",X"77",X"B5",X"50",X"27",X"FF",X"22",X"21",X"22",X"25",X"71",
		X"7C",X"52",X"55",X"55",X"55",X"32",X"71",X"FF",X"22",X"21",X"22",X"25",X"71",X"7C",X"C2",X"22",
		X"33",X"33",X"30",X"27",X"FF",X"22",X"22",X"22",X"25",X"57",X"5C",X"C5",X"23",X"55",X"55",X"55",
		X"00",X"FF",X"22",X"22",X"22",X"22",X"55",X"55",X"55",X"25",X"5C",X"CC",X"CC",X"00",X"FF",X"22",
		X"22",X"22",X"22",X"20",X"22",X"33",X"25",X"5C",X"CC",X"CC",X"00",X"FF",X"02",X"B1",X"11",X"B2",
		X"00",X"22",X"22",X"22",X"55",X"55",X"CC",X"00",X"FF",X"00",X"BB",X"BB",X"B0",X"00",X"22",X"B1",
		X"1B",X"22",X"00",X"50",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"02",X"BB",X"BB",X"20",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"71",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"22",X"22",X"21",X"11",X"70",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"02",X"22",X"22",X"27",X"11",X"1C",X"A0",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"22",X"21",X"22",X"25",X"17",X"C5",X"30",X"00",X"00",X"00",X"00",X"00",X"FF",X"22",X"21",
		X"22",X"25",X"55",X"33",X"55",X"55",X"53",X"3C",X"C0",X"00",X"FF",X"22",X"22",X"22",X"25",X"53",
		X"55",X"55",X"B5",X"55",X"53",X"CC",X"00",X"FF",X"22",X"22",X"22",X"22",X"25",X"52",X"5B",X"BB",
		X"55",X"55",X"3C",X"00",X"FF",X"22",X"22",X"22",X"22",X"55",X"55",X"5B",X"77",X"55",X"C6",X"5C",
		X"00",X"FF",X"02",X"BB",X"BB",X"B3",X"55",X"52",X"5B",X"17",X"55",X"C1",X"C5",X"00",X"FF",X"00",
		X"BB",X"BB",X"B3",X"55",X"55",X"5B",X"71",X"55",X"C1",X"15",X"27",X"FF",X"00",X"00",X"00",X"03",
		X"55",X"52",X"5B",X"17",X"55",X"C6",X"15",X"71",X"FF",X"00",X"00",X"00",X"03",X"55",X"55",X"55",
		X"75",X"55",X"C6",X"C5",X"27",X"FF",X"00",X"00",X"00",X"03",X"55",X"55",X"55",X"55",X"55",X"5C",
		X"55",X"00",X"FF",X"00",X"00",X"00",X"02",X"25",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"FF",
		X"00",X"22",X"22",X"23",X"33",X"35",X"55",X"55",X"55",X"55",X"55",X"00",X"FF",X"02",X"22",X"22",
		X"25",X"71",X"53",X"33",X"55",X"77",X"B5",X"50",X"27",X"FF",X"22",X"21",X"22",X"21",X"11",X"7C",
		X"52",X"55",X"55",X"55",X"32",X"71",X"FF",X"22",X"21",X"22",X"27",X"11",X"1C",X"C2",X"22",X"33",
		X"33",X"30",X"27",X"FF",X"22",X"22",X"22",X"25",X"17",X"5C",X"C5",X"23",X"55",X"55",X"55",X"00",
		X"FF",X"22",X"22",X"22",X"22",X"55",X"55",X"55",X"25",X"5C",X"CC",X"CC",X"00",X"FF",X"22",X"22",
		X"22",X"22",X"20",X"22",X"33",X"25",X"5C",X"CC",X"CC",X"00",X"FF",X"02",X"B1",X"11",X"B2",X"00",
		X"22",X"22",X"22",X"55",X"55",X"CC",X"00",X"FF",X"00",X"BB",X"BB",X"B0",X"00",X"22",X"B1",X"1B",
		X"22",X"00",X"50",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"02",X"BB",X"BB",X"20",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"22",X"22",X"20",X"01",X"11",X"10",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"02",X"22",X"22",X"22",X"11",X"11",X"11",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"22",X"21",X"22",X"22",X"11",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"22",X"21",X"22",X"22",X"21",X"11",X"13",X"30",X"00",X"00",X"00",X"00",X"FF",X"22",X"22",X"22",
		X"22",X"25",X"11",X"55",X"55",X"55",X"00",X"00",X"00",X"FF",X"22",X"22",X"22",X"22",X"22",X"55",
		X"52",X"5B",X"B5",X"55",X"00",X"00",X"FF",X"22",X"22",X"22",X"22",X"33",X"55",X"55",X"57",X"BB",
		X"5C",X"50",X"00",X"FF",X"02",X"BB",X"BB",X"B3",X"33",X"55",X"52",X"51",X"7B",X"5C",X"C5",X"00",
		X"FF",X"00",X"BB",X"BB",X"B3",X"33",X"55",X"55",X"57",X"7B",X"5C",X"6C",X"50",X"FF",X"00",X"00",
		X"00",X"03",X"33",X"55",X"52",X"57",X"7B",X"5C",X"16",X"50",X"FF",X"00",X"00",X"00",X"03",X"32",
		X"55",X"55",X"51",X"75",X"5C",X"16",X"50",X"FF",X"00",X"00",X"00",X"03",X"32",X"11",X"55",X"55",
		X"55",X"5C",X"66",X"50",X"FF",X"00",X"00",X"00",X"00",X"31",X"11",X"15",X"55",X"55",X"CC",X"1C",
		X"50",X"FF",X"00",X"22",X"22",X"20",X"11",X"11",X"11",X"55",X"55",X"5C",X"CC",X"50",X"FF",X"02",
		X"22",X"22",X"22",X"11",X"11",X"11",X"35",X"55",X"55",X"C5",X"00",X"FF",X"22",X"21",X"22",X"22",
		X"21",X"11",X"15",X"35",X"57",X"75",X"55",X"00",X"FF",X"22",X"21",X"22",X"22",X"20",X"11",X"CC",
		X"34",X"5B",X"7B",X"50",X"00",X"FF",X"22",X"22",X"22",X"22",X"20",X"05",X"CC",X"23",X"45",X"B5",
		X"00",X"00",X"FF",X"22",X"22",X"22",X"22",X"20",X"03",X"5C",X"22",X"33",X"50",X"00",X"00",X"FF",
		X"22",X"22",X"22",X"22",X"20",X"03",X"53",X"55",X"53",X"32",X"70",X"00",X"FF",X"02",X"B1",X"11",
		X"B2",X"22",X"25",X"25",X"CC",X"C5",X"57",X"10",X"00",X"FF",X"00",X"BB",X"BB",X"B2",X"22",X"22",
		X"25",X"55",X"CC",X"52",X"70",X"00",X"FF",X"00",X"00",X"00",X"02",X"22",X"22",X"22",X"20",X"5C",
		X"50",X"00",X"00",X"FF",X"00",X"00",X"00",X"02",X"22",X"22",X"22",X"20",X"05",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"02",X"2B",X"11",X"B2",X"20",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"2B",X"BB",X"B2",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"22",X"22",X"20",X"00",X"71",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"02",
		X"22",X"22",X"22",X"01",X"11",X"70",X"00",X"00",X"00",X"00",X"00",X"FF",X"22",X"21",X"22",X"22",
		X"27",X"11",X"15",X"00",X"00",X"00",X"00",X"00",X"FF",X"22",X"21",X"22",X"22",X"25",X"17",X"33",
		X"30",X"00",X"00",X"00",X"00",X"FF",X"22",X"22",X"22",X"22",X"25",X"33",X"55",X"55",X"55",X"00",
		X"00",X"00",X"FF",X"22",X"22",X"22",X"22",X"22",X"55",X"52",X"5B",X"B5",X"55",X"00",X"00",X"FF",
		X"22",X"22",X"22",X"22",X"33",X"55",X"55",X"57",X"BB",X"5C",X"50",X"00",X"FF",X"02",X"BB",X"BB",
		X"B3",X"33",X"55",X"52",X"51",X"7B",X"5C",X"C5",X"00",X"FF",X"00",X"BB",X"BB",X"B3",X"33",X"55",
		X"55",X"57",X"7B",X"5C",X"6C",X"50",X"FF",X"00",X"00",X"00",X"03",X"33",X"55",X"52",X"57",X"7B",
		X"5C",X"16",X"50",X"FF",X"00",X"00",X"00",X"03",X"32",X"55",X"55",X"51",X"75",X"5C",X"16",X"50",
		X"FF",X"00",X"00",X"00",X"03",X"32",X"23",X"55",X"55",X"55",X"5C",X"66",X"50",X"FF",X"00",X"00",
		X"00",X"00",X"35",X"71",X"35",X"55",X"55",X"CC",X"1C",X"50",X"FF",X"00",X"22",X"22",X"20",X"31",
		X"11",X"73",X"55",X"55",X"5C",X"CC",X"50",X"FF",X"02",X"22",X"22",X"22",X"37",X"11",X"15",X"35",
		X"55",X"55",X"C5",X"00",X"FF",X"22",X"21",X"22",X"22",X"25",X"17",X"C5",X"35",X"57",X"75",X"55",
		X"00",X"FF",X"22",X"21",X"22",X"22",X"20",X"5C",X"CC",X"34",X"5B",X"7B",X"50",X"00",X"FF",X"22",
		X"22",X"22",X"22",X"20",X"05",X"CC",X"23",X"45",X"B5",X"00",X"00",X"FF",X"22",X"22",X"22",X"22",
		X"20",X"03",X"5C",X"22",X"33",X"50",X"00",X"00",X"FF",X"22",X"22",X"22",X"22",X"20",X"03",X"53",
		X"55",X"53",X"32",X"70",X"00",X"FF",X"02",X"B1",X"11",X"B2",X"22",X"25",X"25",X"CC",X"C5",X"57",
		X"10",X"00",X"FF",X"00",X"BB",X"BB",X"B2",X"22",X"22",X"25",X"55",X"CC",X"52",X"70",X"00",X"FF",
		X"00",X"00",X"00",X"02",X"22",X"22",X"22",X"20",X"5C",X"50",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"02",X"22",X"22",X"22",X"20",X"05",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"02",X"2B",X"11",
		X"B2",X"20",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"2B",X"BB",X"B2",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"22",
		X"22",X"20",X"00",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"02",X"22",X"22",X"22",X"03",
		X"53",X"10",X"00",X"00",X"00",X"00",X"00",X"FF",X"22",X"21",X"22",X"22",X"23",X"C1",X"71",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"22",X"21",X"22",X"22",X"23",X"C1",X"71",X"50",X"00",X"00",X"00",
		X"00",X"FF",X"22",X"22",X"22",X"22",X"23",X"55",X"13",X"35",X"00",X"00",X"00",X"00",X"FF",X"22",
		X"22",X"22",X"22",X"23",X"33",X"35",X"55",X"55",X"00",X"00",X"00",X"FF",X"22",X"22",X"22",X"22",
		X"22",X"25",X"55",X"C5",X"55",X"5C",X"00",X"00",X"FF",X"02",X"BB",X"BB",X"B2",X"32",X"55",X"5C",
		X"CC",X"25",X"55",X"C0",X"00",X"FF",X"00",X"BB",X"BB",X"B3",X"32",X"55",X"CC",X"CC",X"55",X"BB",
		X"5C",X"00",X"FF",X"00",X"00",X"22",X"23",X"32",X"55",X"CC",X"CC",X"25",X"1B",X"BC",X"C0",X"FF",
		X"00",X"00",X"22",X"23",X"32",X"55",X"5C",X"CC",X"55",X"71",X"BC",X"C0",X"FF",X"00",X"00",X"02",
		X"23",X"32",X"33",X"55",X"C5",X"25",X"17",X"BC",X"C0",X"FF",X"00",X"00",X"00",X"03",X"32",X"55",
		X"15",X"55",X"55",X"71",X"5C",X"C0",X"FF",X"00",X"22",X"22",X"23",X"32",X"51",X"71",X"55",X"55",
		X"55",X"5C",X"C0",X"FF",X"02",X"22",X"22",X"22",X"32",X"51",X"71",X"35",X"55",X"55",X"CC",X"C0",
		X"FF",X"22",X"21",X"22",X"22",X"22",X"55",X"1C",X"35",X"55",X"55",X"5C",X"C0",X"FF",X"22",X"21",
		X"22",X"22",X"22",X"35",X"5C",X"35",X"55",X"17",X"BC",X"00",X"FF",X"22",X"22",X"22",X"22",X"23",
		X"33",X"5C",X"35",X"55",X"77",X"BC",X"00",X"FF",X"22",X"22",X"22",X"22",X"20",X"33",X"5C",X"35",
		X"55",X"BB",X"C0",X"00",X"FF",X"22",X"22",X"22",X"22",X"20",X"33",X"5C",X"23",X"55",X"5C",X"00",
		X"00",X"FF",X"02",X"B1",X"11",X"B2",X"00",X"33",X"C2",X"33",X"55",X"00",X"00",X"00",X"FF",X"00",
		X"BB",X"BB",X"B2",X"22",X"3C",X"C2",X"53",X"70",X"00",X"00",X"00",X"FF",X"00",X"00",X"22",X"22",
		X"22",X"55",X"55",X"55",X"10",X"00",X"00",X"00",X"FF",X"00",X"00",X"22",X"22",X"22",X"22",X"05",
		X"55",X"70",X"00",X"00",X"00",X"FF",X"00",X"00",X"22",X"22",X"22",X"22",X"00",X"35",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"22",X"B1",X"1B",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"02",X"BB",X"BB",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"22",X"22",X"20",X"55",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"02",X"22",X"22",X"22",X"57",X"10",X"00",X"00",X"00",X"00",X"00",X"FF",X"22",X"21",
		X"22",X"22",X"C7",X"1C",X"00",X"00",X"00",X"00",X"00",X"FF",X"22",X"21",X"22",X"22",X"C5",X"55",
		X"50",X"00",X"00",X"00",X"00",X"FF",X"22",X"22",X"22",X"22",X"55",X"33",X"35",X"00",X"00",X"00",
		X"00",X"FF",X"22",X"22",X"22",X"22",X"33",X"35",X"55",X"55",X"00",X"00",X"00",X"FF",X"22",X"22",
		X"22",X"22",X"25",X"55",X"C5",X"55",X"5C",X"00",X"00",X"FF",X"02",X"BB",X"BB",X"32",X"55",X"5C",
		X"CC",X"25",X"55",X"C0",X"00",X"FF",X"00",X"BB",X"B3",X"32",X"55",X"CC",X"CC",X"55",X"BB",X"5C",
		X"00",X"FF",X"00",X"00",X"03",X"32",X"55",X"CC",X"CC",X"25",X"1B",X"BC",X"C0",X"FF",X"00",X"00",
		X"03",X"32",X"55",X"5C",X"CC",X"55",X"71",X"BC",X"C0",X"FF",X"00",X"00",X"03",X"32",X"33",X"55",
		X"C5",X"25",X"17",X"BC",X"C0",X"FF",X"00",X"00",X"03",X"32",X"55",X"35",X"55",X"55",X"71",X"5C",
		X"C0",X"FF",X"00",X"22",X"22",X"22",X"57",X"13",X"55",X"55",X"55",X"5C",X"C0",X"FF",X"02",X"22",
		X"22",X"22",X"57",X"15",X"35",X"55",X"55",X"CC",X"C0",X"FF",X"22",X"21",X"22",X"22",X"55",X"CC",
		X"35",X"55",X"55",X"5C",X"C0",X"FF",X"22",X"21",X"22",X"22",X"25",X"5C",X"35",X"55",X"17",X"BC",
		X"00",X"FF",X"22",X"22",X"22",X"22",X"23",X"5C",X"35",X"55",X"77",X"BC",X"00",X"FF",X"22",X"22",
		X"22",X"22",X"23",X"5C",X"35",X"55",X"BB",X"C0",X"00",X"FF",X"22",X"22",X"22",X"22",X"23",X"5C",
		X"23",X"55",X"5C",X"00",X"00",X"FF",X"02",X"B1",X"11",X"B2",X"33",X"C2",X"33",X"55",X"00",X"00",
		X"00",X"FF",X"00",X"BB",X"BB",X"B2",X"2C",X"C2",X"53",X"70",X"00",X"00",X"00",X"FF",X"00",X"02",
		X"22",X"22",X"55",X"55",X"55",X"10",X"00",X"00",X"00",X"FF",X"00",X"02",X"22",X"22",X"22",X"25",
		X"55",X"70",X"00",X"00",X"00",X"FF",X"00",X"02",X"22",X"22",X"22",X"20",X"35",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"02",X"2B",X"11",X"B2",X"20",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"2B",X"BB",X"B2",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"02",X"22",
		X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"22",X"22",X"22",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"22",X"22",X"14",X"22",X"22",X"20",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"22",X"22",X"14",X"22",X"22",X"22",X"00",X"00",X"00",X"00",X"00",X"FF",X"22",X"22",
		X"22",X"22",X"24",X"12",X"20",X"00",X"00",X"00",X"00",X"FF",X"26",X"A2",X"22",X"22",X"24",X"12",
		X"20",X"00",X"00",X"00",X"00",X"FF",X"26",X"AA",X"22",X"22",X"24",X"12",X"20",X"00",X"00",X"00",
		X"00",X"FF",X"26",X"AA",X"AA",X"92",X"22",X"22",X"20",X"00",X"00",X"00",X"00",X"FF",X"06",X"A7",
		X"AA",X"99",X"88",X"88",X"88",X"80",X"00",X"00",X"00",X"FF",X"06",X"A7",X"77",X"79",X"88",X"3C",
		X"C8",X"8A",X"00",X"00",X"00",X"FF",X"06",X"A7",X"77",X"7D",X"DD",X"3C",X"CD",X"7A",X"A0",X"00",
		X"00",X"FF",X"06",X"AA",X"77",X"7D",X"DD",X"3C",X"CD",X"77",X"22",X"20",X"00",X"FF",X"06",X"AA",
		X"AA",X"9D",X"DD",X"3C",X"CD",X"77",X"22",X"22",X"00",X"FF",X"06",X"6A",X"AA",X"99",X"88",X"3C",
		X"C8",X"87",X"77",X"02",X"20",X"FF",X"00",X"66",X"AA",X"99",X"88",X"3C",X"C8",X"8A",X"A7",X"00",
		X"20",X"FF",X"02",X"22",X"22",X"69",X"88",X"88",X"88",X"8A",X"22",X"20",X"00",X"FF",X"22",X"22",
		X"22",X"26",X"66",X"66",X"66",X"6A",X"22",X"22",X"00",X"FF",X"22",X"22",X"22",X"22",X"22",X"26",
		X"CC",X"66",X"AA",X"02",X"20",X"FF",X"22",X"22",X"14",X"22",X"22",X"22",X"6C",X"C6",X"6A",X"00",
		X"20",X"FF",X"22",X"22",X"14",X"22",X"22",X"22",X"26",X"66",X"66",X"00",X"00",X"FF",X"22",X"22",
		X"22",X"22",X"22",X"22",X"26",X"60",X"00",X"00",X"00",X"FF",X"22",X"22",X"22",X"22",X"24",X"12",
		X"20",X"00",X"00",X"00",X"00",X"FF",X"22",X"5E",X"52",X"22",X"24",X"12",X"20",X"00",X"00",X"00",
		X"00",X"FF",X"02",X"22",X"22",X"22",X"24",X"12",X"20",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"22",X"22",X"22",X"22",X"20",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"22",X"22",X"22",X"22",
		X"20",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"02",X"25",X"E5",X"22",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"22",X"22",X"20",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"02",X"22",X"22",X"00",X"02",X"22",X"22",X"00",X"00",X"00",X"FF",X"22",X"21",X"42",X"20",X"22",
		X"22",X"22",X"20",X"00",X"00",X"FF",X"22",X"21",X"42",X"22",X"22",X"22",X"41",X"22",X"00",X"00",
		X"FF",X"22",X"22",X"22",X"22",X"22",X"22",X"41",X"22",X"00",X"00",X"FF",X"8A",X"22",X"22",X"22",
		X"22",X"88",X"91",X"22",X"00",X"00",X"FF",X"8A",X"AA",X"22",X"22",X"88",X"8C",X"9A",X"A2",X"22",
		X"00",X"FF",X"87",X"AA",X"AA",X"98",X"88",X"3C",X"DA",X"22",X"22",X"20",X"FF",X"87",X"77",X"AA",
		X"98",X"DD",X"3C",X"D7",X"22",X"AA",X"22",X"FF",X"87",X"77",X"77",X"7D",X"DD",X"3C",X"D7",X"77",
		X"7A",X"02",X"FF",X"8A",X"77",X"77",X"7D",X"DD",X"3C",X"97",X"72",X"22",X"00",X"FF",X"8A",X"AA",
		X"77",X"7D",X"88",X"3C",X"9A",X"22",X"22",X"20",X"FF",X"8A",X"AA",X"AA",X"98",X"88",X"38",X"9A",
		X"22",X"A7",X"22",X"FF",X"66",X"AA",X"AA",X"98",X"88",X"88",X"89",X"AA",X"AA",X"02",X"FF",X"66",
		X"66",X"AA",X"98",X"88",X"66",X"66",X"69",X"AA",X"00",X"FF",X"06",X"66",X"66",X"66",X"66",X"66",
		X"6C",X"C6",X"66",X"00",X"FF",X"02",X"22",X"22",X"66",X"62",X"22",X"22",X"CC",X"60",X"00",X"FF",
		X"22",X"22",X"22",X"26",X"22",X"22",X"22",X"26",X"60",X"00",X"FF",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"00",X"00",X"FF",X"22",X"21",X"42",X"22",X"22",X"22",X"22",X"22",X"00",X"00",
		X"FF",X"22",X"21",X"42",X"22",X"22",X"22",X"41",X"22",X"00",X"00",X"FF",X"22",X"22",X"22",X"22",
		X"22",X"22",X"41",X"22",X"00",X"00",X"FF",X"22",X"22",X"22",X"22",X"22",X"22",X"41",X"22",X"00",
		X"00",X"FF",X"22",X"5E",X"52",X"22",X"22",X"22",X"22",X"22",X"00",X"00",X"FF",X"02",X"22",X"22",
		X"02",X"22",X"22",X"22",X"22",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"22",X"5E",X"52",X"20",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"02",X"22",X"22",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"02",X"22",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"22",X"22",X"22",
		X"22",X"00",X"00",X"00",X"00",X"00",X"FF",X"22",X"22",X"14",X"22",X"20",X"00",X"00",X"00",X"00",
		X"FF",X"22",X"22",X"14",X"22",X"22",X"00",X"00",X"00",X"00",X"FF",X"22",X"8A",X"22",X"24",X"12",
		X"00",X"00",X"00",X"00",X"FF",X"22",X"9A",X"A2",X"24",X"12",X"00",X"00",X"00",X"00",X"FF",X"22",
		X"97",X"A9",X"24",X"12",X"00",X"00",X"00",X"00",X"FF",X"22",X"97",X"79",X"98",X"22",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"97",X"77",X"98",X"88",X"88",X"8A",X"00",X"00",X"FF",X"00",X"9A",X"77",
		X"7D",X"88",X"8C",X"38",X"A0",X"00",X"FF",X"00",X"9A",X"A7",X"7D",X"DD",X"DC",X"38",X"A0",X"00",
		X"FF",X"00",X"9A",X"A9",X"7D",X"DD",X"DC",X"3D",X"AA",X"00",X"FF",X"00",X"66",X"A9",X"98",X"DD",
		X"DC",X"3D",X"72",X"20",X"FF",X"00",X"86",X"69",X"98",X"88",X"8C",X"3D",X"72",X"22",X"FF",X"00",
		X"06",X"66",X"66",X"88",X"8C",X"38",X"77",X"02",X"FF",X"02",X"22",X"22",X"66",X"66",X"68",X"88",
		X"A7",X"02",X"FF",X"22",X"22",X"22",X"22",X"66",X"66",X"66",X"A2",X"20",X"FF",X"22",X"22",X"22",
		X"22",X"26",X"6C",X"C6",X"82",X"22",X"FF",X"22",X"22",X"14",X"22",X"22",X"66",X"CC",X"6A",X"02",
		X"FF",X"22",X"22",X"14",X"22",X"22",X"66",X"66",X"6A",X"02",X"FF",X"22",X"22",X"22",X"24",X"12",
		X"66",X"00",X"00",X"02",X"FF",X"22",X"22",X"22",X"24",X"12",X"00",X"00",X"00",X"00",X"FF",X"22",
		X"5E",X"52",X"24",X"12",X"00",X"00",X"00",X"00",X"FF",X"02",X"22",X"22",X"22",X"22",X"00",X"00",
		X"00",X"00",X"FF",X"02",X"22",X"22",X"22",X"22",X"00",X"00",X"00",X"00",X"FF",X"00",X"22",X"5E",
		X"52",X"20",X"00",X"00",X"00",X"00",X"FF",X"00",X"02",X"22",X"22",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"22",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"02",X"22",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"22",X"22",X"32",X"22",
		X"20",X"00",X"00",X"00",X"00",X"00",X"FF",X"22",X"23",X"32",X"22",X"22",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"22",X"23",X"22",X"22",X"22",X"20",X"00",X"00",X"00",X"00",X"FF",X"22",X"22",X"26",
		X"A2",X"22",X"22",X"00",X"00",X"00",X"00",X"FF",X"22",X"22",X"26",X"A2",X"23",X"22",X"00",X"00",
		X"00",X"00",X"FF",X"22",X"22",X"66",X"A2",X"33",X"22",X"00",X"00",X"00",X"00",X"FF",X"02",X"22",
		X"66",X"A9",X"32",X"22",X"00",X"00",X"00",X"00",X"FF",X"00",X"22",X"66",X"A9",X"98",X"88",X"90",
		X"00",X"00",X"00",X"FF",X"00",X"22",X"66",X"A7",X"98",X"C3",X"9A",X"00",X"00",X"00",X"FF",X"00",
		X"22",X"66",X"A7",X"77",X"C3",X"7A",X"A0",X"00",X"00",X"FF",X"00",X"02",X"66",X"A7",X"77",X"C3",
		X"77",X"22",X"20",X"00",X"FF",X"00",X"00",X"66",X"99",X"77",X"C3",X"77",X"22",X"22",X"20",X"FF",
		X"00",X"22",X"66",X"69",X"98",X"C3",X"97",X"70",X"00",X"00",X"FF",X"02",X"22",X"26",X"66",X"68",
		X"C3",X"9A",X"70",X"00",X"00",X"FF",X"22",X"23",X"22",X"66",X"66",X"68",X"9A",X"22",X"20",X"00",
		X"FF",X"22",X"23",X"32",X"22",X"26",X"66",X"69",X"22",X"22",X"20",X"FF",X"22",X"22",X"32",X"22",
		X"22",X"66",X"66",X"90",X"00",X"00",X"FF",X"22",X"22",X"22",X"22",X"22",X"26",X"66",X"60",X"00",
		X"00",X"FF",X"22",X"22",X"22",X"22",X"32",X"26",X"60",X"00",X"00",X"00",X"FF",X"22",X"22",X"E2",
		X"22",X"33",X"22",X"00",X"00",X"00",X"00",X"FF",X"02",X"2E",X"22",X"22",X"23",X"22",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"22",X"22",X"22",X"22",X"22",X"00",X"00",X"00",X"00",X"FF",X"00",X"22",
		X"22",X"22",X"22",X"22",X"00",X"00",X"00",X"00",X"FF",X"00",X"22",X"22",X"22",X"2E",X"22",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"02",X"22",X"22",X"E2",X"20",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"22",X"22",X"22",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"02",X"22",X"20",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"02",X"22",X"22",X"22",X"20",X"00",X"91",X"10",
		X"00",X"00",X"00",X"FF",X"22",X"23",X"42",X"22",X"22",X"01",X"12",X"81",X"00",X"00",X"00",X"FF",
		X"22",X"23",X"42",X"22",X"21",X"19",X"12",X"81",X"00",X"00",X"00",X"FF",X"22",X"22",X"22",X"21",
		X"11",X"97",X"12",X"81",X"00",X"00",X"00",X"FF",X"22",X"22",X"21",X"11",X"97",X"78",X"81",X"10",
		X"00",X"00",X"00",X"FF",X"22",X"27",X"11",X"97",X"78",X"82",X"22",X"22",X"20",X"00",X"00",X"FF",
		X"02",X"29",X"97",X"78",X"22",X"22",X"21",X"12",X"22",X"BB",X"B0",X"FF",X"00",X"09",X"98",X"22",
		X"22",X"21",X"12",X"81",X"22",X"BB",X"B0",X"FF",X"00",X"00",X"AA",X"22",X"21",X"19",X"12",X"81",
		X"22",X"00",X"20",X"FF",X"00",X"00",X"AA",X"21",X"11",X"97",X"12",X"81",X"22",X"AA",X"20",X"FF",
		X"00",X"00",X"A1",X"19",X"77",X"78",X"81",X"12",X"22",X"00",X"00",X"FF",X"00",X"09",X"97",X"77",
		X"88",X"88",X"22",X"22",X"22",X"BB",X"B0",X"FF",X"00",X"09",X"78",X"88",X"52",X"22",X"22",X"22",
		X"22",X"BB",X"B0",X"FF",X"02",X"22",X"22",X"22",X"25",X"22",X"22",X"22",X"22",X"00",X"20",X"FF",
		X"22",X"23",X"42",X"22",X"22",X"52",X"22",X"22",X"22",X"AA",X"20",X"FF",X"22",X"23",X"42",X"22",
		X"22",X"52",X"2C",X"CC",X"22",X"00",X"00",X"FF",X"22",X"22",X"22",X"22",X"22",X"52",X"22",X"C2",
		X"20",X"00",X"00",X"FF",X"22",X"22",X"22",X"22",X"22",X"55",X"22",X"22",X"00",X"00",X"00",X"FF",
		X"22",X"29",X"11",X"92",X"22",X"55",X"52",X"20",X"00",X"00",X"00",X"FF",X"02",X"22",X"22",X"22",
		X"22",X"22",X"25",X"22",X"22",X"00",X"00",X"FF",X"00",X"00",X"00",X"22",X"22",X"22",X"22",X"50",
		X"22",X"00",X"00",X"FF",X"00",X"00",X"00",X"22",X"22",X"22",X"22",X"50",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"22",X"91",X"19",X"22",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"02",
		X"22",X"22",X"20",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"09",X"11",
		X"10",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"11",X"88",X"81",X"00",X"00",X"00",X"FF",
		X"02",X"22",X"22",X"21",X"11",X"22",X"81",X"00",X"00",X"00",X"FF",X"22",X"34",X"22",X"19",X"81",
		X"22",X"81",X"00",X"00",X"00",X"FF",X"22",X"34",X"21",X"97",X"78",X"11",X"12",X"2B",X"D0",X"00",
		X"FF",X"22",X"22",X"19",X"77",X"88",X"88",X"22",X"BB",X"DD",X"00",X"FF",X"22",X"29",X"97",X"78",
		X"29",X"11",X"15",X"B2",X"5D",X"00",X"FF",X"22",X"99",X"77",X"82",X"11",X"88",X"81",X"22",X"50",
		X"00",X"FF",X"02",X"97",X"78",X"21",X"11",X"22",X"81",X"22",X"52",X"00",X"FF",X"00",X"99",X"8A",
		X"11",X"81",X"22",X"81",X"2B",X"D2",X"20",X"FF",X"00",X"00",X"A1",X"19",X"77",X"11",X"12",X"BB",
		X"DD",X"20",X"FF",X"00",X"00",X"91",X"97",X"78",X"88",X"22",X"B2",X"5D",X"22",X"FF",X"00",X"09",
		X"19",X"77",X"88",X"22",X"55",X"22",X"52",X"22",X"FF",X"00",X"99",X"87",X"78",X"22",X"22",X"22",
		X"52",X"52",X"22",X"FF",X"00",X"99",X"78",X"55",X"52",X"22",X"22",X"25",X"52",X"22",X"FF",X"02",
		X"22",X"22",X"22",X"25",X"22",X"2C",X"22",X"52",X"22",X"FF",X"22",X"34",X"22",X"22",X"22",X"52",
		X"CC",X"C2",X"52",X"22",X"FF",X"22",X"34",X"22",X"22",X"22",X"52",X"22",X"22",X"52",X"22",X"FF",
		X"22",X"22",X"22",X"22",X"22",X"55",X"55",X"55",X"22",X"22",X"FF",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"52",X"22",X"FF",X"22",X"29",X"11",X"92",X"22",X"22",X"22",X"22",X"25",X"22",
		X"FF",X"02",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"25",X"20",X"FF",X"00",X"00",X"00",X"00",
		X"02",X"29",X"11",X"92",X"20",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"22",X"22",X"22",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"02",X"22",X"22",X"22",X"20",X"00",X"00",X"00",X"00",X"00",X"FF",X"22",X"22",
		X"34",X"22",X"22",X"00",X"00",X"00",X"00",X"00",X"FF",X"22",X"22",X"34",X"22",X"22",X"00",X"01",
		X"11",X"11",X"00",X"FF",X"22",X"22",X"22",X"22",X"99",X"11",X"11",X"99",X"12",X"10",X"FF",X"22",
		X"22",X"29",X"99",X"11",X"99",X"99",X"99",X"12",X"10",X"FF",X"22",X"29",X"91",X"11",X"77",X"77",
		X"77",X"77",X"12",X"10",X"FF",X"02",X"29",X"17",X"77",X"88",X"88",X"88",X"88",X"81",X"00",X"FF",
		X"00",X"09",X"88",X"88",X"22",X"22",X"22",X"22",X"00",X"00",X"FF",X"00",X"00",X"AA",X"A2",X"22",
		X"22",X"22",X"11",X"11",X"00",X"FF",X"00",X"00",X"AA",X"A2",X"29",X"91",X"11",X"19",X"12",X"10",
		X"FF",X"00",X"00",X"AA",X"99",X"99",X"11",X"99",X"99",X"12",X"10",X"FF",X"00",X"09",X"99",X"99",
		X"77",X"77",X"77",X"77",X"12",X"10",X"FF",X"00",X"09",X"88",X"88",X"88",X"88",X"88",X"88",X"81",
		X"00",X"FF",X"02",X"22",X"22",X"22",X"28",X"88",X"22",X"22",X"00",X"00",X"FF",X"22",X"22",X"14",
		X"22",X"22",X"52",X"22",X"22",X"BB",X"00",X"FF",X"22",X"22",X"14",X"22",X"22",X"52",X"22",X"22",
		X"BB",X"00",X"FF",X"22",X"22",X"22",X"22",X"22",X"52",X"22",X"22",X"02",X"00",X"FF",X"22",X"22",
		X"22",X"22",X"22",X"52",X"CC",X"22",X"A2",X"00",X"FF",X"22",X"29",X"11",X"92",X"22",X"52",X"C2",
		X"20",X"00",X"00",X"FF",X"02",X"22",X"22",X"22",X"25",X"52",X"22",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"05",X"55",X"55",X"22",X"20",X"00",X"00",X"00",X"FF",X"00",X"00",X"22",X"22",X"22",X"55",
		X"22",X"20",X"00",X"00",X"FF",X"00",X"02",X"22",X"22",X"22",X"25",X"02",X"20",X"00",X"00",X"FF",
		X"00",X"02",X"22",X"22",X"22",X"22",X"00",X"00",X"00",X"00",X"FF",X"00",X"02",X"29",X"11",X"92",
		X"20",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"22",X"22",X"22",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"02",X"22",X"22",X"20",X"66",X"61",
		X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"22",X"22",X"22",X"2A",X"66",X"61",X"66",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"22",X"23",X"42",X"2A",X"66",X"61",X"56",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"22",X"23",X"42",X"AA",X"22",X"21",X"56",X"60",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"22",X"22",X"22",X"AA",X"22",X"21",X"55",X"60",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"22",X"22",X"22",X"AA",X"66",X"61",X"55",X"62",X"22",X"22",X"25",X"02",X"20",X"FF",X"22",X"22",
		X"92",X"AA",X"66",X"61",X"55",X"56",X"66",X"60",X"22",X"21",X"12",X"FF",X"02",X"22",X"92",X"AA",
		X"66",X"61",X"55",X"55",X"55",X"66",X"02",X"21",X"12",X"FF",X"00",X"00",X"92",X"AA",X"66",X"61",
		X"88",X"8D",X"DD",X"56",X"02",X"02",X"20",X"FF",X"00",X"00",X"92",X"AA",X"66",X"61",X"88",X"8D",
		X"DD",X"56",X"02",X"00",X"00",X"FF",X"00",X"00",X"92",X"AA",X"22",X"21",X"88",X"8D",X"DD",X"56",
		X"02",X"02",X"20",X"FF",X"00",X"00",X"92",X"AA",X"22",X"21",X"88",X"8D",X"DD",X"56",X"02",X"21",
		X"12",X"FF",X"00",X"00",X"92",X"AA",X"66",X"61",X"88",X"88",X"88",X"56",X"02",X"21",X"12",X"FF",
		X"00",X"00",X"92",X"AA",X"66",X"61",X"88",X"8D",X"DD",X"56",X"02",X"02",X"20",X"FF",X"02",X"22",
		X"22",X"AA",X"66",X"61",X"88",X"8D",X"DD",X"56",X"02",X"00",X"00",X"FF",X"22",X"22",X"22",X"AA",
		X"99",X"91",X"C8",X"8D",X"DD",X"56",X"02",X"02",X"20",X"FF",X"22",X"23",X"42",X"22",X"99",X"99",
		X"1C",X"8D",X"DD",X"56",X"02",X"21",X"12",X"FF",X"22",X"23",X"42",X"22",X"22",X"29",X"91",X"78",
		X"88",X"66",X"22",X"21",X"12",X"FF",X"22",X"22",X"22",X"22",X"22",X"22",X"99",X"72",X"22",X"22",
		X"20",X"02",X"20",X"FF",X"22",X"22",X"22",X"22",X"22",X"22",X"99",X"66",X"66",X"66",X"00",X"00",
		X"00",X"FF",X"22",X"E1",X"1E",X"22",X"22",X"99",X"99",X"99",X"66",X"60",X"00",X"00",X"00",X"FF",
		X"02",X"22",X"22",X"22",X"22",X"22",X"22",X"99",X"60",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"02",X"22",X"22",X"22",X"22",X"29",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"02",X"2E",
		X"11",X"E2",X"29",X"99",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"22",X"22",X"22",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"99",X"16",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"02",X"22",
		X"29",X"99",X"16",X"60",X"00",X"00",X"22",X"20",X"22",X"FF",X"22",X"22",X"29",X"99",X"15",X"66",
		X"00",X"22",X"20",X"22",X"12",X"FF",X"22",X"34",X"29",X"92",X"15",X"56",X"62",X"29",X"99",X"22",
		X"12",X"FF",X"22",X"34",X"A2",X"22",X"15",X"55",X"56",X"99",X"99",X"20",X"20",X"FF",X"22",X"22",
		X"A2",X"99",X"15",X"55",X"55",X"95",X"59",X"26",X"00",X"FF",X"22",X"22",X"A9",X"99",X"15",X"55",
		X"55",X"5E",X"59",X"26",X"22",X"FF",X"22",X"22",X"A9",X"99",X"18",X"55",X"55",X"EE",X"59",X"22",
		X"12",X"FF",X"02",X"22",X"A9",X"99",X"18",X"88",X"55",X"EE",X"59",X"22",X"12",X"FF",X"00",X"00",
		X"A9",X"99",X"18",X"88",X"55",X"EE",X"59",X"26",X"20",X"FF",X"00",X"00",X"A9",X"92",X"18",X"88",
		X"55",X"E5",X"59",X"26",X"60",X"FF",X"00",X"00",X"A2",X"22",X"18",X"88",X"55",X"5E",X"59",X"26",
		X"22",X"FF",X"00",X"00",X"A2",X"99",X"18",X"88",X"55",X"EE",X"59",X"22",X"12",X"FF",X"00",X"00",
		X"A9",X"99",X"18",X"88",X"55",X"EE",X"59",X"22",X"12",X"FF",X"00",X"00",X"A9",X"99",X"18",X"88",
		X"55",X"EE",X"59",X"26",X"20",X"FF",X"02",X"22",X"A9",X"96",X"61",X"18",X"55",X"E5",X"22",X"26",
		X"60",X"FF",X"22",X"22",X"26",X"66",X"67",X"71",X"15",X"22",X"29",X"66",X"60",X"FF",X"22",X"34",
		X"22",X"22",X"22",X"66",X"62",X"29",X"99",X"99",X"60",X"FF",X"22",X"34",X"22",X"22",X"22",X"26",
		X"66",X"66",X"99",X"99",X"60",X"FF",X"22",X"22",X"22",X"22",X"22",X"26",X"66",X"66",X"66",X"96",
		X"00",X"FF",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"26",X"66",X"00",X"FF",X"22",X"E1",
		X"1E",X"22",X"22",X"22",X"22",X"22",X"22",X"60",X"00",X"FF",X"02",X"22",X"22",X"20",X"22",X"22",
		X"22",X"22",X"66",X"60",X"00",X"FF",X"00",X"00",X"00",X"00",X"22",X"E1",X"1E",X"22",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"02",X"22",X"22",X"20",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"02",X"22",X"22",X"20",X"00",X"66",X"60",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"22",X"22",X"22",X"22",X"0A",X"66",X"60",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"22",X"22",X"34",X"22",X"AA",X"66",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"22",X"22",X"34",X"2A",X"AA",X"22",X"29",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"22",X"22",X"22",X"2A",X"AA",X"22",X"29",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"22",X"22",
		X"22",X"2A",X"AA",X"66",X"69",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"22",X"22",X"92",X"2A",
		X"AA",X"66",X"69",X"22",X"20",X"00",X"00",X"00",X"00",X"FF",X"02",X"22",X"92",X"2A",X"AA",X"66",
		X"69",X"67",X"22",X"20",X"00",X"00",X"00",X"FF",X"00",X"05",X"95",X"5A",X"AA",X"66",X"69",X"55",
		X"67",X"22",X"20",X"22",X"00",X"FF",X"00",X"02",X"92",X"2A",X"AA",X"66",X"69",X"85",X"55",X"70",
		X"22",X"11",X"20",X"FF",X"00",X"02",X"92",X"2A",X"AA",X"22",X"29",X"DD",X"D5",X"70",X"22",X"11",
		X"20",X"FF",X"00",X"02",X"92",X"2A",X"AA",X"22",X"29",X"DD",X"D5",X"70",X"20",X"22",X"00",X"FF",
		X"00",X"02",X"92",X"2A",X"AA",X"66",X"69",X"DD",X"D5",X"70",X"20",X"00",X"00",X"FF",X"00",X"00",
		X"92",X"2A",X"AA",X"66",X"69",X"DD",X"D5",X"70",X"20",X"22",X"00",X"FF",X"02",X"22",X"22",X"2A",
		X"AA",X"66",X"69",X"88",X"85",X"70",X"22",X"11",X"20",X"FF",X"22",X"22",X"22",X"2A",X"A9",X"99",
		X"69",X"DD",X"D5",X"70",X"22",X"11",X"20",X"FF",X"22",X"22",X"34",X"29",X"99",X"99",X"69",X"DD",
		X"D5",X"70",X"20",X"22",X"00",X"FF",X"22",X"22",X"34",X"29",X"99",X"99",X"69",X"DD",X"D5",X"70",
		X"20",X"00",X"00",X"FF",X"22",X"22",X"22",X"22",X"22",X"29",X"69",X"DD",X"D5",X"70",X"20",X"22",
		X"00",X"FF",X"22",X"22",X"22",X"22",X"22",X"29",X"67",X"88",X"85",X"70",X"22",X"11",X"20",X"FF",
		X"22",X"E1",X"1E",X"22",X"22",X"99",X"97",X"22",X"22",X"22",X"22",X"11",X"20",X"FF",X"02",X"22",
		X"22",X"22",X"99",X"99",X"99",X"99",X"99",X"90",X"00",X"22",X"00",X"FF",X"00",X"02",X"22",X"22",
		X"99",X"99",X"99",X"99",X"90",X"00",X"00",X"00",X"00",X"FF",X"00",X"02",X"22",X"22",X"22",X"22",
		X"99",X"90",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"02",X"22",X"22",X"22",X"22",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"02",X"22",X"22",X"22",X"29",X"99",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"02",X"2E",X"11",X"E2",X"29",X"90",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"22",X"22",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"55",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"22",X"22",X"53",X"80",X"00",X"00",X"00",X"07",X"10",X"FF",
		X"00",X"02",X"22",X"22",X"C3",X"8C",X"00",X"00",X"00",X"17",X"70",X"FF",X"00",X"22",X"22",X"12",
		X"C5",X"55",X"50",X"00",X"C0",X"77",X"70",X"FF",X"02",X"22",X"21",X"22",X"55",X"55",X"50",X"05",
		X"5C",X"71",X"00",X"FF",X"02",X"B2",X"22",X"22",X"35",X"55",X"00",X"08",X"85",X"C0",X"00",X"FF",
		X"0B",X"BB",X"22",X"22",X"22",X"20",X"00",X"00",X"88",X"CC",X"00",X"FF",X"00",X"8B",X"B2",X"22",
		X"22",X"52",X"50",X"17",X"08",X"CC",X"00",X"FF",X"00",X"08",X"BC",X"C2",X"25",X"C5",X"50",X"71",
		X"18",X"C1",X"00",X"FF",X"00",X"00",X"B5",X"CC",X"5C",X"25",X"60",X"17",X"10",X"05",X"10",X"FF",
		X"00",X"00",X"00",X"5C",X"5C",X"55",X"60",X"07",X"00",X"00",X"51",X"FF",X"00",X"00",X"00",X"00",
		X"55",X"56",X"05",X"50",X"0C",X"C0",X"00",X"FF",X"00",X"00",X"00",X"00",X"65",X"56",X"55",X"CC",
		X"05",X"CC",X"00",X"FF",X"00",X"AE",X"EE",X"A0",X"05",X"60",X"33",X"5C",X"03",X"CC",X"00",X"FF",
		X"0E",X"EE",X"EE",X"EE",X"05",X"50",X"88",X"5C",X"33",X"C0",X"00",X"FF",X"A2",X"EE",X"EE",X"EE",
		X"A5",X"53",X"55",X"CC",X"3C",X"00",X"00",X"FF",X"E2",X"1E",X"EE",X"EE",X"E5",X"55",X"55",X"CC",
		X"30",X"07",X"00",X"FF",X"EE",X"E2",X"AA",X"AE",X"E5",X"C5",X"55",X"55",X"50",X"07",X"70",X"FF",
		X"EE",X"EA",X"98",X"9A",X"E0",X"5C",X"25",X"55",X"00",X"00",X"00",X"FF",X"AE",X"EA",X"88",X"9A",
		X"E2",X"22",X"22",X"27",X"00",X"00",X"00",X"FF",X"0E",X"EA",X"98",X"9A",X"0B",X"B2",X"22",X"77",
		X"00",X"00",X"00",X"FF",X"00",X"A2",X"AA",X"A0",X"08",X"BB",X"22",X"20",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"8B",X"22",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"05",X"53",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"0A",X"22",X"22",X"0C",X"C5",X"80",X"00",X"00",X"00",X"07",X"10",X"FF",X"00",
		X"21",X"12",X"2B",X"B3",X"3C",X"55",X"00",X"00",X"00",X"07",X"10",X"FF",X"0A",X"22",X"22",X"BB",
		X"B3",X"3C",X"C5",X"00",X"00",X"80",X"71",X"10",X"FF",X"02",X"22",X"22",X"BB",X"22",X"33",X"C5",
		X"00",X"05",X"58",X"71",X"00",X"FF",X"02",X"22",X"22",X"BB",X"22",X"23",X"C0",X"00",X"85",X"55",
		X"80",X"00",X"FF",X"02",X"22",X"22",X"B6",X"55",X"20",X"00",X"00",X"68",X"55",X"58",X"00",X"FF",
		X"0A",X"22",X"22",X"65",X"54",X"50",X"00",X"00",X"01",X"85",X"58",X"00",X"FF",X"00",X"22",X"26",
		X"55",X"44",X"45",X"00",X"00",X"07",X"18",X"80",X"00",X"FF",X"00",X"0A",X"26",X"54",X"44",X"55",
		X"00",X"00",X"00",X"71",X"64",X"40",X"FF",X"00",X"00",X"06",X"55",X"55",X"55",X"00",X"00",X"00",
		X"07",X"64",X"44",X"FF",X"00",X"00",X"00",X"65",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"54",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"50",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"5C",X"51",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"55",X"5C",X"61",X"00",X"FF",X"00",X"22",X"22",X"B0",X"00",X"00",X"00",X"00",
		X"55",X"16",X"60",X"00",X"FF",X"02",X"22",X"22",X"2B",X"00",X"00",X"00",X"05",X"56",X"36",X"00",
		X"00",X"FF",X"AA",X"B2",X"22",X"22",X"B5",X"C0",X"00",X"05",X"56",X"31",X"00",X"00",X"FF",X"BB",
		X"BB",X"21",X"12",X"2C",X"35",X"00",X"05",X"56",X"33",X"00",X"00",X"FF",X"22",X"BB",X"22",X"22",
		X"2C",X"33",X"30",X"22",X"55",X"63",X"00",X"77",X"FF",X"22",X"BB",X"22",X"22",X"25",X"C3",X"32",
		X"22",X"55",X"50",X"00",X"00",X"FF",X"22",X"BB",X"22",X"22",X"20",X"5C",X"52",X"22",X"27",X"70",
		X"00",X"00",X"FF",X"02",X"BB",X"22",X"22",X"00",X"00",X"0B",X"B2",X"27",X"20",X"00",X"00",X"FF",
		X"00",X"B2",X"22",X"20",X"00",X"00",X"0B",X"BB",X"22",X"20",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"BB",X"22",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"05",X"63",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"55",X"63",X"30",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"22",X"22",X"B0",X"55",X"63",X"30",X"00",X"00",X"00",X"01",
		X"00",X"00",X"FF",X"00",X"02",X"22",X"22",X"2B",X"55",X"56",X"33",X"00",X"00",X"00",X"07",X"10",
		X"00",X"FF",X"00",X"AA",X"B2",X"22",X"22",X"B5",X"55",X"63",X"00",X"00",X"05",X"80",X"71",X"00",
		X"FF",X"00",X"BB",X"BB",X"21",X"12",X"20",X"55",X"66",X"00",X"00",X"55",X"88",X"07",X"00",X"FF",
		X"00",X"22",X"BB",X"22",X"44",X"46",X"00",X"00",X"00",X"00",X"55",X"58",X"00",X"00",X"FF",X"00",
		X"22",X"BB",X"24",X"44",X"41",X"00",X"00",X"00",X"00",X"55",X"58",X"80",X"00",X"FF",X"00",X"22",
		X"BB",X"44",X"44",X"41",X"00",X"00",X"CC",X"00",X"05",X"71",X"80",X"00",X"FF",X"00",X"02",X"BB",
		X"44",X"46",X"10",X"00",X"00",X"5C",X"C0",X"00",X"71",X"00",X"00",X"FF",X"00",X"00",X"B2",X"44",
		X"66",X"00",X"00",X"00",X"05",X"C0",X"07",X"11",X"00",X"00",X"FF",X"00",X"00",X"06",X"44",X"10",
		X"00",X"00",X"00",X"00",X"00",X"07",X"10",X"00",X"00",X"FF",X"00",X"00",X"06",X"66",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"FF",X"00",X"00",X"00",X"65",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"CC",X"60",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"66",X"60",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"89",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"55",
		X"58",X"85",X"50",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"66",X"55",
		X"55",X"50",X"00",X"FF",X"00",X"A2",X"22",X"20",X"00",X"00",X"00",X"00",X"06",X"33",X"65",X"55",
		X"00",X"00",X"FF",X"02",X"11",X"22",X"BB",X"00",X"00",X"00",X"00",X"0C",X"33",X"36",X"50",X"00",
		X"00",X"FF",X"A2",X"22",X"2B",X"BB",X"20",X"00",X"00",X"00",X"0C",X"33",X"36",X"60",X"00",X"00",
		X"FF",X"22",X"22",X"2B",X"B2",X"22",X"5C",X"00",X"00",X"0C",X"33",X"33",X"60",X"00",X"00",X"FF",
		X"22",X"22",X"2B",X"B2",X"22",X"55",X"C0",X"00",X"00",X"C3",X"33",X"60",X"07",X"70",X"FF",X"22",
		X"22",X"2B",X"B2",X"22",X"33",X"5C",X"00",X"00",X"23",X"33",X"60",X"07",X"00",X"FF",X"A2",X"22",
		X"22",X"BB",X"2B",X"33",X"3C",X"00",X"02",X"22",X"27",X"70",X"00",X"00",X"FF",X"02",X"22",X"22",
		X"2B",X"B0",X"03",X"3C",X"00",X"02",X"22",X"22",X"22",X"00",X"00",X"FF",X"00",X"A2",X"22",X"22",
		X"00",X"00",X"00",X"00",X"02",X"2B",X"B2",X"22",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"02",X"BB",X"BB",X"22",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"2B",X"B2",X"20",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"50",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"05",X"5C",X"C5",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"05",X"33",X"CC",
		X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"AE",X"EE",X"A0",X"00",X"88",X"CC",
		X"50",X"00",X"00",X"00",X"01",X"70",X"00",X"FF",X"00",X"0E",X"EE",X"EE",X"EE",X"00",X"55",X"CC",
		X"50",X"00",X"00",X"00",X"07",X"11",X"00",X"FF",X"00",X"A2",X"EE",X"EE",X"EE",X"A0",X"05",X"55",
		X"00",X"00",X"00",X"05",X"61",X"71",X"00",X"FF",X"00",X"E2",X"1E",X"EE",X"EE",X"E0",X"00",X"00",
		X"00",X"00",X"00",X"55",X"56",X"70",X"00",X"FF",X"00",X"EE",X"E5",X"55",X"5E",X"E0",X"00",X"00",
		X"00",X"00",X"00",X"55",X"56",X"00",X"00",X"FF",X"00",X"EE",X"55",X"5C",X"25",X"E0",X"00",X"00",
		X"00",X"00",X"00",X"55",X"55",X"60",X"00",X"FF",X"00",X"AE",X"55",X"CC",X"55",X"E0",X"00",X"00",
		X"00",X"10",X"00",X"05",X"55",X"60",X"00",X"FF",X"00",X"0E",X"EA",X"5C",X"25",X"00",X"00",X"00",
		X"00",X"51",X"00",X"05",X"67",X"10",X"00",X"FF",X"00",X"00",X"A2",X"A5",X"55",X"00",X"00",X"00",
		X"00",X"05",X"10",X"00",X"17",X"70",X"00",X"FF",X"00",X"00",X"0C",X"C5",X"25",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"77",X"70",X"00",X"FF",X"00",X"00",X"0C",X"C5",X"50",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"71",X"00",X"00",X"FF",X"00",X"00",X"06",X"66",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"5C",X"C0",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"05",X"C0",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"55",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"55",X"50",X"05",X"5C",X"C0",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"55",X"55",X"05",X"CC",X"C0",X"00",X"FF",X"00",X"02",X"22",X"2B",X"00",X"00",X"00",X"00",
		X"00",X"55",X"38",X"5C",X"CC",X"C0",X"00",X"FF",X"00",X"22",X"22",X"22",X"20",X"00",X"00",X"00",
		X"00",X"55",X"38",X"55",X"CC",X"00",X"00",X"FF",X"02",X"22",X"21",X"22",X"2B",X"00",X"00",X"00",
		X"00",X"55",X"5C",X"C5",X"C0",X"00",X"00",X"FF",X"22",X"22",X"12",X"22",X"22",X"00",X"00",X"00",
		X"00",X"03",X"55",X"C5",X"00",X"00",X"00",X"FF",X"2B",X"22",X"22",X"22",X"22",X"55",X"00",X"00",
		X"00",X"00",X"35",X"C2",X"00",X"00",X"00",X"FF",X"BB",X"B2",X"22",X"22",X"22",X"CC",X"50",X"00",
		X"00",X"08",X"B2",X"22",X"20",X"00",X"70",X"FF",X"08",X"BB",X"22",X"22",X"22",X"CC",X"C0",X"00",
		X"00",X"BB",X"22",X"72",X"20",X"07",X"70",X"FF",X"00",X"8B",X"22",X"22",X"23",X"55",X"C0",X"00",
		X"00",X"B2",X"22",X"77",X"20",X"00",X"00",X"FF",X"00",X"0B",X"22",X"22",X"00",X"03",X"50",X"00",
		X"00",X"22",X"22",X"22",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"22",X"20",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"53",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"C3",X"8C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"22",X"22",X"B0",X"00",X"C5",X"55",
		X"50",X"00",X"00",X"00",X"00",X"07",X"10",X"FF",X"00",X"02",X"22",X"22",X"22",X"00",X"55",X"55",
		X"50",X"00",X"00",X"00",X"00",X"17",X"70",X"FF",X"00",X"22",X"22",X"12",X"22",X"B0",X"35",X"55",
		X"00",X"00",X"00",X"00",X"0C",X"77",X"70",X"FF",X"02",X"22",X"21",X"22",X"22",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"55",X"71",X"00",X"FF",X"02",X"B2",X"25",X"25",X"22",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"88",X"5C",X"00",X"FF",X"0B",X"BB",X"5C",X"55",X"22",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"8C",X"C0",X"FF",X"00",X"85",X"C2",X"56",X"22",X"20",X"00",X"00",
		X"00",X"64",X"40",X"00",X"00",X"8C",X"C0",X"FF",X"00",X"05",X"C5",X"56",X"22",X"00",X"00",X"00",
		X"00",X"64",X"44",X"00",X"00",X"17",X"C0",X"FF",X"00",X"05",X"55",X"62",X"20",X"00",X"00",X"00",
		X"00",X"06",X"54",X"00",X"00",X"71",X"10",X"FF",X"00",X"06",X"55",X"60",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"17",X"10",X"FF",X"00",X"00",X"56",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"FF",X"00",X"00",X"5C",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"05",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"05",X"10",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"51",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"CC",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"05",X"CC",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"05",X"50",X"03",X"CC",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"55",X"CC",X"33",X"C0",X"00",X"FF",X"00",X"AE",X"EE",X"A0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"33",X"5C",X"3C",X"00",X"00",X"FF",X"0E",X"EE",X"EE",X"EE",X"00",X"00",X"00",X"00",
		X"00",X"00",X"88",X"5C",X"C0",X"00",X"00",X"FF",X"A2",X"EE",X"EE",X"EE",X"A0",X"00",X"00",X"00",
		X"00",X"00",X"55",X"CC",X"00",X"00",X"00",X"FF",X"E2",X"1E",X"EE",X"EE",X"E0",X"00",X"00",X"00",
		X"00",X"00",X"55",X"CC",X"30",X"00",X"00",X"FF",X"EE",X"E2",X"AA",X"AE",X"E5",X"00",X"00",X"00",
		X"00",X"00",X"85",X"55",X"50",X"00",X"70",X"FF",X"EE",X"EA",X"98",X"9A",X"E5",X"30",X"00",X"00",
		X"00",X"02",X"B5",X"55",X"22",X"70",X"77",X"FF",X"AE",X"EA",X"88",X"9A",X"E5",X"53",X"50",X"00",
		X"00",X"02",X"22",X"22",X"27",X"70",X"00",X"FF",X"0E",X"EA",X"98",X"9A",X"5C",X"55",X"50",X"00",
		X"00",X"02",X"22",X"22",X"22",X"00",X"00",X"FF",X"00",X"A2",X"AA",X"A0",X"05",X"C5",X"00",X"00",
		X"00",X"00",X"22",X"22",X"20",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"22",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"05",
		X"53",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"C5",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"3C",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"0A",X"22",X"22",
		X"00",X"00",X"03",X"3C",X"C5",X"00",X"00",X"00",X"00",X"00",X"07",X"10",X"FF",X"00",X"21",X"12",
		X"2B",X"B0",X"00",X"00",X"33",X"C5",X"00",X"00",X"00",X"00",X"00",X"07",X"10",X"FF",X"0A",X"22",
		X"22",X"BB",X"B2",X"00",X"00",X"03",X"C0",X"00",X"00",X"00",X"00",X"08",X"71",X"10",X"FF",X"02",
		X"22",X"22",X"BB",X"22",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"71",X"00",X"FF",
		X"02",X"26",X"55",X"BB",X"22",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"55",X"58",X"00",
		X"FF",X"02",X"65",X"54",X"5B",X"22",X"20",X"00",X"00",X"00",X"00",X"0C",X"C0",X"06",X"85",X"55",
		X"80",X"FF",X"06",X"55",X"44",X"45",X"B2",X"B0",X"00",X"00",X"00",X"00",X"0C",X"C6",X"00",X"68",
		X"55",X"80",X"FF",X"06",X"54",X"44",X"55",X"BB",X"00",X"00",X"00",X"00",X"00",X"06",X"66",X"00",
		X"06",X"88",X"00",X"FF",X"06",X"55",X"55",X"55",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"FF",X"00",X"65",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"07",X"10",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"71",X"FF",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"FF",X"00",X"05",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"51",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"64",X"40",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"64",X"44",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"54",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"55",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"55",X"10",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"56",
		X"10",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"C5",
		X"66",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"55",
		X"C5",X"60",X"00",X"FF",X"00",X"22",X"22",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",
		X"51",X"01",X"10",X"00",X"FF",X"02",X"22",X"22",X"2B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"63",X"00",X"00",X"00",X"FF",X"AA",X"B2",X"22",X"22",X"B0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"55",X"63",X"00",X"00",X"00",X"FF",X"BB",X"BB",X"21",X"12",X"25",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"55",X"63",X"30",X"00",X"77",X"FF",X"22",X"BB",X"22",X"22",X"2C",X"35",X"00",X"00",
		X"00",X"00",X"02",X"25",X"56",X"3B",X"77",X"00",X"FF",X"22",X"BB",X"22",X"22",X"2C",X"33",X"30",
		X"00",X"00",X"00",X"02",X"25",X"55",X"8B",X"70",X"00",X"FF",X"22",X"BB",X"22",X"22",X"25",X"C3",
		X"30",X"00",X"00",X"00",X"02",X"22",X"B8",X"8B",X"00",X"00",X"FF",X"02",X"BB",X"22",X"22",X"00",
		X"5C",X"50",X"00",X"00",X"00",X"02",X"22",X"BB",X"B0",X"00",X"00",X"FF",X"00",X"B2",X"22",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"22",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"53",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"55",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"0A",X"22",X"22",X"00",X"00",X"03",X"30",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"07",X"10",X"FF",X"00",X"21",X"12",X"2B",X"B0",X"00",X"00",X"03",X"C5",X"00",X"00",X"00",
		X"00",X"00",X"07",X"10",X"FF",X"0A",X"22",X"22",X"0B",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"08",X"71",X"10",X"FF",X"02",X"22",X"22",X"BB",X"22",X"20",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"05",X"01",X"00",X"FF",X"02",X"26",X"55",X"BB",X"02",X"20",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"55",X"08",X"00",X"FF",X"02",X"65",X"50",X"5B",X"20",X"00",X"00",X"00",
		X"00",X"00",X"00",X"C0",X"06",X"05",X"55",X"80",X"FF",X"06",X"05",X"44",X"45",X"B2",X"B0",X"00",
		X"00",X"00",X"00",X"0C",X"06",X"00",X"68",X"05",X"80",X"FF",X"06",X"54",X"44",X"55",X"0B",X"00",
		X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"06",X"88",X"00",X"FF",X"06",X"50",X"05",X"05",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"00",X"65",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"71",X"FF",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"FF",X"00",
		X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",
		X"40",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"60",X"44",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"06",X"54",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"55",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"05",X"05",X"10",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"10",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"05",X"05",X"66",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"C0",X"60",X"00",X"FF",X"00",X"20",X"02",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"01",X"01",X"10",X"00",X"FF",X"00",X"02",X"22",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"63",X"00",X"00",X"00",X"FF",X"0A",X"B2",X"02",
		X"22",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"63",X"00",X"00",X"00",X"FF",X"0B",X"BB",
		X"21",X"12",X"25",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"60",X"30",X"00",X"70",X"FF",X"22",
		X"0B",X"22",X"02",X"0C",X"00",X"00",X"00",X"00",X"00",X"02",X"20",X"56",X"3B",X"70",X"00",X"FF",
		X"22",X"BB",X"22",X"20",X"2C",X"30",X"30",X"00",X"00",X"00",X"00",X"20",X"55",X"0B",X"70",X"00",
		X"FF",X"22",X"BB",X"22",X"22",X"25",X"C3",X"30",X"00",X"00",X"00",X"00",X"02",X"B8",X"8B",X"00",
		X"00",X"FF",X"02",X"BB",X"22",X"22",X"00",X"5C",X"50",X"00",X"00",X"00",X"00",X"02",X"BB",X"B0",
		X"00",X"00",X"FF",X"00",X"B2",X"22",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"22",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"50",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3C",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"0A",X"02",X"02",X"00",X"00",
		X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"FF",X"00",X"21",X"10",X"00",X"B0",
		X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"FF",X"0A",X"02",X"20",X"0B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"71",X"00",X"FF",X"00",X"20",X"20",
		X"B0",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"01",X"00",X"FF",X"02",X"26",
		X"00",X"B0",X"02",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"05",X"08",X"00",X"FF",X"00",
		X"65",X"50",X"5B",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"06",X"00",X"55",X"80",X"FF",
		X"06",X"05",X"04",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"08",X"05",X"80",
		X"FF",X"00",X"54",X"04",X"50",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"06",X"88",
		X"00",X"FF",X"06",X"50",X"05",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"FF",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"40",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"44",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"54",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"10",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"05",X"66",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"60",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"01",X"01",
		X"10",X"00",X"FF",X"00",X"02",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"60",
		X"00",X"00",X"00",X"FF",X"00",X"B2",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"63",X"00",X"00",X"00",X"FF",X"00",X"BB",X"20",X"12",X"25",X"00",X"00",X"00",X"00",X"00",X"00",
		X"50",X"60",X"30",X"00",X"70",X"FF",X"22",X"0B",X"22",X"02",X"0C",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"06",X"0B",X"70",X"00",X"FF",X"20",X"B0",X"20",X"20",X"20",X"30",X"00",X"00",X"00",
		X"00",X"00",X"20",X"55",X"0B",X"70",X"00",X"FF",X"02",X"BB",X"22",X"22",X"25",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"02",X"B8",X"80",X"00",X"00",X"FF",X"02",X"BB",X"02",X"02",X"00",X"50",X"00",
		X"00",X"00",X"00",X"00",X"02",X"0B",X"00",X"00",X"00",X"FF",X"00",X"02",X"20",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"02",X"02",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",
		X"FF",X"00",X"21",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"FF",X"0A",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"71",X"00",X"FF",X"00",X"00",X"20",X"B0",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"05",X"00",X"00",X"FF",X"02",X"26",X"00",X"B0",X"02",X"20",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"00",X"08",X"00",X"FF",X"00",X"05",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"06",X"00",X"50",X"80",X"FF",X"06",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"06",X"00",X"08",X"00",X"00",X"FF",X"00",X"04",X"04",X"00",X"0B",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"06",X"00",X"00",X"05",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"05",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"04",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"05",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"06",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"FF",X"00",X"00",X"20",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"FF",X"00",X"02",X"00",X"02",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"B0",X"00",X"00",X"05",
		X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"60",X"30",X"00",X"70",X"FF",X"20",X"00",X"02",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"FF",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"FF",X"00",X"B0",
		X"00",X"20",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"FF",
		X"00",X"02",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"70",X"00",X"FF",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"00",X"FF",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"07",X"10",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"50",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"50",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"50",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"03",X"00",X"07",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"05",X"50",X"55",X"00",X"00",X"FF",X"00",X"55",X"D5",X"D5",X"50",X"00",X"FF",X"05",X"DD",X"5D",
		X"D5",X"D5",X"00",X"FF",X"05",X"DD",X"5D",X"5D",X"D5",X"00",X"FF",X"55",X"55",X"DD",X"DD",X"DD",
		X"50",X"FF",X"5D",X"D5",X"55",X"DD",X"55",X"50",X"FF",X"5D",X"DD",X"5D",X"55",X"DD",X"50",X"FF",
		X"5D",X"DD",X"5D",X"D5",X"DD",X"50",X"FF",X"05",X"55",X"DD",X"DD",X"55",X"00",X"FF",X"00",X"5D",
		X"DD",X"DD",X"50",X"00",X"FF",X"00",X"55",X"D5",X"55",X"50",X"00",X"FF",X"00",X"05",X"50",X"55",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"05",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"05",X"00",X"00",X"05",X"5E",X"00",X"FF",X"E5",X"50",
		X"B5",X"5B",X"1B",X"55",X"00",X"00",X"FF",X"00",X"55",X"1B",X"B1",X"BB",X"BB",X"00",X"00",X"FF",
		X"00",X"0B",X"B1",X"11",X"11",X"1B",X"55",X"E0",X"FF",X"00",X"0B",X"11",X"51",X"11",X"1B",X"50",
		X"00",X"FF",X"00",X"00",X"15",X"11",X"11",X"15",X"B0",X"00",X"FF",X"00",X"0B",X"55",X"11",X"B1",
		X"1B",X"B0",X"00",X"FF",X"00",X"0B",X"15",X"11",X"51",X"1B",X"00",X"00",X"FF",X"00",X"0B",X"B1",
		X"15",X"1B",X"BB",X"00",X"00",X"FF",X"00",X"05",X"B1",X"B1",X"55",X"BB",X"00",X"00",X"FF",X"00",
		X"55",X"51",X"11",X"BB",X"B5",X"00",X"00",X"FF",X"00",X"50",X"00",X"00",X"00",X"05",X"50",X"00",
		X"FF",X"04",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"0E",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"E0",X"00",X"50",X"00",X"E0",X"00",X"E0",X"FF",X"00",X"05",
		X"50",X"55",X"05",X"00",X"05",X"00",X"FF",X"00",X"00",X"55",X"55",X"55",X"55",X"50",X"00",X"FF",
		X"E5",X"55",X"B4",X"BB",X"55",X"BD",X"50",X"00",X"FF",X"00",X"55",X"DB",X"D5",X"5B",X"11",X"50",
		X"0E",X"FF",X"00",X"05",X"D1",X"1D",X"5B",X"1B",X"55",X"50",X"FF",X"00",X"05",X"B4",X"D5",X"5E",
		X"DB",X"50",X"00",X"FF",X"0E",X"5B",X"D5",X"55",X"55",X"DD",X"50",X"00",X"FF",X"00",X"01",X"BD",
		X"DD",X"BB",X"DD",X"50",X"00",X"FF",X"00",X"54",X"D5",X"D1",X"DB",X"15",X"55",X"E0",X"FF",X"00",
		X"55",X"51",X"11",X"BD",X"BD",X"40",X"00",X"FF",X"00",X"55",X"1D",X"DD",X"DD",X"B5",X"50",X"00",
		X"FF",X"00",X"55",X"55",X"05",X"D4",X"55",X"50",X"00",X"FF",X"05",X"05",X"00",X"05",X"50",X"50",
		X"05",X"00",X"FF",X"E0",X"0E",X"00",X"05",X"00",X"50",X"00",X"E0",X"FF",X"00",X"00",X"00",X"0E",
		X"00",X"E0",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"E0",X"00",X"00",X"50",X"00",X"05",X"00",X"04",X"40",X"00",X"FF",X"00",X"05",
		X"00",X"05",X"DB",X"B5",X"55",X"00",X"55",X"00",X"00",X"FF",X"00",X"05",X"5B",X"5D",X"DB",X"55",
		X"5B",X"BB",X"55",X"00",X"00",X"FF",X"00",X"00",X"5B",X"55",X"55",X"5D",X"55",X"B5",X"55",X"00",
		X"00",X"FF",X"E0",X"0B",X"55",X"51",X"B1",X"BD",X"5D",X"55",X"00",X"00",X"00",X"FF",X"05",X"55",
		X"5D",X"51",X"B1",X"15",X"15",X"D5",X"B0",X"0E",X"00",X"FF",X"00",X"0D",X"DD",X"55",X"BB",X"1B",
		X"15",X"D5",X"55",X"50",X"00",X"FF",X"00",X"5B",X"B1",X"15",X"55",X"BB",X"55",X"D1",X"1B",X"00",
		X"00",X"FF",X"00",X"5D",X"DB",X"15",X"DD",X"D5",X"1D",X"D5",X"B5",X"50",X"00",X"FF",X"00",X"5D",
		X"D5",X"55",X"D5",X"5D",X"B5",X"D5",X"55",X"55",X"40",X"FF",X"05",X"05",X"DB",X"5D",X"D1",X"15",
		X"D5",X"D1",X"BB",X"00",X"00",X"FF",X"00",X"55",X"B5",X"15",X"D1",X"15",X"D5",X"55",X"B5",X"00",
		X"00",X"FF",X"00",X"5D",X"5B",X"15",X"DB",X"B5",X"B1",X"55",X"55",X"55",X"E0",X"FF",X"00",X"5D",
		X"DB",X"B5",X"D5",X"5B",X"15",X"5D",X"D5",X"00",X"00",X"FF",X"E5",X"BD",X"DD",X"51",X"11",X"5B",
		X"15",X"DD",X"50",X"00",X"00",X"FF",X"00",X"00",X"D5",X"BB",X"11",X"55",X"B5",X"D5",X"55",X"00",
		X"00",X"FF",X"00",X"05",X"5D",X"55",X"BB",X"B5",X"55",X"BB",X"05",X"50",X"00",X"FF",X"00",X"00",
		X"0B",X"D5",X"55",X"55",X"DD",X"D5",X"00",X"04",X"00",X"FF",X"00",X"00",X"05",X"5B",X"55",X"5B",
		X"5D",X"D5",X"50",X"00",X"00",X"FF",X"00",X"00",X"05",X"00",X"05",X"50",X"5D",X"05",X"50",X"00",
		X"00",X"FF",X"00",X"00",X"E0",X"00",X"05",X"00",X"50",X"00",X"0E",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"55",
		X"00",X"00",X"60",X"00",X"FF",X"60",X"00",X"55",X"55",X"50",X"00",X"00",X"00",X"FF",X"00",X"05",
		X"55",X"D5",X"DD",X"55",X"50",X"00",X"FF",X"00",X"05",X"00",X"51",X"0D",X"5D",X"55",X"00",X"FF",
		X"00",X"55",X"15",X"0D",X"05",X"D1",X"55",X"50",X"FF",X"05",X"55",X"1D",X"0D",X"55",X"DD",X"D5",
		X"50",X"FF",X"05",X"55",X"55",X"D5",X"05",X"D5",X"15",X"50",X"FF",X"55",X"5D",X"5D",X"05",X"D0",
		X"00",X"5D",X"00",X"FF",X"55",X"D0",X"05",X"D5",X"5D",X"55",X"00",X"55",X"FF",X"55",X"D5",X"55",
		X"D1",X"55",X"55",X"15",X"55",X"FF",X"00",X"D0",X"1D",X"15",X"D5",X"DD",X"DD",X"55",X"FF",X"05",
		X"55",X"1D",X"55",X"1D",X"1D",X"55",X"D0",X"FF",X"05",X"5D",X"55",X"05",X"D5",X"DD",X"55",X"50",
		X"FF",X"05",X"55",X"5D",X"01",X"50",X"51",X"D5",X"50",X"FF",X"00",X"55",X"55",X"D5",X"51",X"0D",
		X"55",X"00",X"FF",X"60",X"05",X"0D",X"01",X"55",X"55",X"55",X"00",X"FF",X"00",X"05",X"05",X"55",
		X"55",X"50",X"00",X"00",X"FF",X"00",X"00",X"00",X"55",X"55",X"00",X"60",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"D0",X"00",X"00",X"00",X"60",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"0D",X"DD",X"50",X"D0",X"50",X"00",X"FF",X"00",X"6D",X"11",X"10",X"D5",X"D5",X"00",X"FF",X"00",
		X"66",X"11",X"D0",X"5D",X"15",X"50",X"FF",X"00",X"D6",X"D1",X"DD",X"DD",X"DD",X"50",X"FF",X"00",
		X"00",X"D0",X"0D",X"6D",X"51",X"00",X"FF",X"0D",X"D5",X"D0",X"16",X"D1",X"11",X"00",X"FF",X"D6",
		X"11",X"5D",X"56",X"D1",X"11",X"00",X"FF",X"D1",X"1D",X"11",X"16",X"6D",X"51",X"55",X"FF",X"D6",
		X"1D",X"61",X"DD",X"D1",X"DD",X"D5",X"FF",X"06",X"1D",X"61",X"5D",X"D1",X"D5",X"5D",X"FF",X"0D",
		X"6D",X"D6",X"00",X"6D",X"11",X"55",X"FF",X"05",X"D6",X"DD",X"15",X"6D",X"11",X"10",X"FF",X"00",
		X"5D",X"51",X"50",X"6D",X"1D",X"50",X"FF",X"00",X"00",X"D0",X"D0",X"06",X"DD",X"00",X"FF",X"0D",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"FF",X"00",
		X"00",X"00",X"D0",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"0D",X"00",X"FF",X"D0",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"05",X"11",X"10",X"00",X"00",X"FF",X"00",X"06",X"61",X"D0",X"00",X"00",X"FF",
		X"00",X"06",X"5D",X"10",X"61",X"00",X"FF",X"00",X"00",X"01",X"05",X"66",X"10",X"FF",X"00",X"15",
		X"00",X"0D",X"5D",X"10",X"FF",X"06",X"DD",X"10",X"00",X"5D",X"00",X"FF",X"0D",X"6D",X"1D",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"DD",X"56",X"D1",X"00",X"FF",X"00",X"61",X"1D",X"55",X"1D",X"10",
		X"FF",X"05",X"DD",X"50",X"66",X"51",X"00",X"FF",X"00",X"6D",X"10",X"06",X"11",X"00",X"FF",X"00",
		X"01",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"0D",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"FF",X"00",X"06",X"0D",X"00",
		X"FF",X"00",X"6D",X"D0",X"D0",X"FF",X"00",X"0D",X"DD",X"60",X"FF",X"00",X"06",X"D0",X"04",X"FF",
		X"00",X"00",X"00",X"D0",X"FF",X"D6",X"D0",X"04",X"6D",X"FF",X"05",X"DD",X"00",X"DD",X"FF",X"00",
		X"D0",X"0D",X"D0",X"FF",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"22",X"22",X"20",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"02",X"22",X"22",
		X"22",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"22",X"22",X"22",X"22",X"C0",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"22",X"22",X"22",X"22",X"2C",X"00",X"00",X"FF",X"00",X"00",X"00",X"22",X"22",
		X"22",X"22",X"2C",X"00",X"00",X"FF",X"00",X"00",X"00",X"22",X"22",X"22",X"22",X"55",X"50",X"00",
		X"FF",X"02",X"22",X"22",X"22",X"22",X"22",X"24",X"55",X"55",X"00",X"FF",X"22",X"22",X"22",X"22",
		X"BB",X"33",X"25",X"55",X"55",X"00",X"FF",X"22",X"22",X"22",X"33",X"33",X"33",X"25",X"55",X"C5",
		X"50",X"FF",X"22",X"22",X"22",X"33",X"33",X"33",X"25",X"55",X"CC",X"50",X"FF",X"22",X"22",X"22",
		X"33",X"33",X"33",X"25",X"55",X"CC",X"50",X"FF",X"22",X"BB",X"B3",X"33",X"33",X"33",X"25",X"55",
		X"CC",X"50",X"FF",X"02",X"BB",X"33",X"33",X"33",X"33",X"25",X"55",X"CC",X"50",X"FF",X"00",X"00",
		X"33",X"33",X"22",X"22",X"25",X"55",X"C5",X"50",X"FF",X"00",X"00",X"33",X"32",X"22",X"22",X"22",
		X"55",X"55",X"50",X"FF",X"00",X"00",X"33",X"22",X"22",X"22",X"22",X"25",X"55",X"50",X"FF",X"00",
		X"00",X"33",X"22",X"22",X"22",X"22",X"25",X"55",X"50",X"FF",X"00",X"00",X"33",X"22",X"22",X"22",
		X"22",X"2C",X"55",X"00",X"FF",X"00",X"00",X"33",X"22",X"22",X"22",X"22",X"2C",X"55",X"00",X"FF",
		X"02",X"22",X"22",X"22",X"22",X"22",X"22",X"2C",X"50",X"00",X"FF",X"22",X"22",X"22",X"22",X"B8",
		X"88",X"B2",X"C5",X"00",X"00",X"FF",X"22",X"22",X"22",X"22",X"BB",X"BB",X"BC",X"00",X"00",X"00",
		X"FF",X"22",X"22",X"22",X"22",X"55",X"5C",X"C0",X"00",X"00",X"00",X"FF",X"22",X"22",X"22",X"22",
		X"55",X"00",X"00",X"00",X"00",X"00",X"FF",X"22",X"B8",X"8B",X"22",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"02",X"BB",X"BB",X"2C",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"01",X"00",X"00",X"22",X"22",X"20",X"00",X"FF",X"00",X"00",
		X"11",X"01",X"00",X"02",X"22",X"22",X"22",X"00",X"FF",X"00",X"01",X"E1",X"11",X"00",X"22",X"22",
		X"22",X"22",X"20",X"FF",X"00",X"EE",X"12",X"22",X"10",X"22",X"22",X"22",X"22",X"20",X"FF",X"0E",
		X"E1",X"22",X"22",X"20",X"22",X"22",X"22",X"22",X"20",X"FF",X"0D",X"E1",X"11",X"22",X"21",X"22",
		X"22",X"22",X"22",X"20",X"FF",X"0E",X"12",X"21",X"22",X"13",X"22",X"33",X"33",X"22",X"20",X"FF",
		X"11",X"11",X"22",X"22",X"23",X"33",X"33",X"33",X"32",X"00",X"FF",X"ED",X"11",X"22",X"33",X"33",
		X"33",X"33",X"33",X"35",X"00",X"FF",X"DE",X"13",X"E3",X"33",X"33",X"23",X"33",X"33",X"35",X"00",
		X"FF",X"01",X"E1",X"33",X"31",X"13",X"23",X"33",X"33",X"30",X"00",X"FF",X"00",X"13",X"33",X"33",
		X"23",X"23",X"33",X"33",X"30",X"00",X"FF",X"00",X"13",X"3E",X"33",X"23",X"23",X"33",X"33",X"30",
		X"00",X"FF",X"00",X"13",X"11",X"E3",X"23",X"33",X"22",X"22",X"20",X"00",X"FF",X"01",X"11",X"33",
		X"33",X"33",X"12",X"22",X"22",X"22",X"00",X"FF",X"00",X"D1",X"EE",X"33",X"13",X"12",X"22",X"22",
		X"22",X"20",X"FF",X"E1",X"11",X"22",X"21",X"33",X"22",X"22",X"22",X"22",X"20",X"FF",X"EE",X"22",
		X"22",X"22",X"23",X"22",X"22",X"22",X"22",X"20",X"FF",X"E1",X"12",X"22",X"22",X"23",X"22",X"22",
		X"22",X"22",X"20",X"FF",X"11",X"12",X"21",X"21",X"23",X"22",X"22",X"22",X"22",X"20",X"FF",X"E1",
		X"11",X"12",X"12",X"23",X"52",X"B8",X"88",X"B2",X"00",X"FF",X"EE",X"11",X"11",X"B2",X"25",X"55",
		X"BB",X"BB",X"B5",X"00",X"FF",X"E1",X"10",X"EB",X"B2",X"11",X"51",X"55",X"55",X"50",X"00",X"FF",
		X"0E",X"11",X"11",X"11",X"00",X"15",X"55",X"50",X"00",X"00",X"FF",X"0E",X"E1",X"E0",X"11",X"10",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"E1",X"11",X"E1",X"01",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"01",X"00",X"10",X"10",X"01",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"EE",X"00",X"01",X"11",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"0E",X"EE",X"10",X"11",X"11",X"10",X"01",X"00",X"10",X"01",
		X"00",X"00",X"FF",X"0E",X"EE",X"11",X"22",X"12",X"21",X"00",X"11",X"10",X"00",X"00",X"00",X"00",
		X"FF",X"E0",X"E0",X"12",X"22",X"22",X"22",X"10",X"00",X"01",X"10",X"00",X"00",X"00",X"FF",X"0E",
		X"E1",X"11",X"12",X"22",X"22",X"21",X"01",X"10",X"00",X"00",X"00",X"00",X"FF",X"00",X"E1",X"12",
		X"22",X"22",X"22",X"21",X"10",X"00",X"00",X"00",X"00",X"01",X"FF",X"0E",X"01",X"11",X"12",X"22",
		X"22",X"20",X"00",X"01",X"00",X"00",X"00",X"00",X"FF",X"00",X"EE",X"11",X"11",X"22",X"22",X"21",
		X"00",X"00",X"00",X"00",X"10",X"00",X"FF",X"EE",X"E1",X"11",X"13",X"32",X"22",X"21",X"11",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"0E",X"01",X"E1",X"33",X"33",X"32",X"11",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"0E",X"EE",X"11",X"13",X"11",X"31",X"00",X"00",X"00",X"01",X"10",X"00",X"00",
		X"FF",X"EE",X"0E",X"11",X"11",X"13",X"31",X"11",X"10",X"00",X"11",X"00",X"00",X"00",X"FF",X"0E",
		X"EE",X"1E",X"1E",X"E1",X"31",X"10",X"00",X"01",X"00",X"00",X"00",X"00",X"FF",X"0E",X"E1",X"1E",
		X"31",X"33",X"31",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"FF",X"00",X"E1",X"11",X"11",X"33",
		X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"EE",X"E1",X"11",X"12",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"0E",X"E1",X"EE",X"22",X"12",X"22",X"11",X"00",X"00",
		X"11",X"00",X"00",X"00",X"FF",X"0E",X"E1",X"11",X"21",X"22",X"22",X"20",X"11",X"10",X"00",X"01",
		X"00",X"00",X"FF",X"0E",X"E1",X"11",X"21",X"22",X"22",X"20",X"00",X"00",X"00",X"10",X"00",X"00",
		X"FF",X"0E",X"E1",X"E1",X"12",X"22",X"22",X"21",X"10",X"00",X"00",X"00",X"00",X"00",X"FF",X"0E",
		X"E1",X"11",X"12",X"22",X"22",X"20",X"01",X"00",X"00",X"10",X"00",X"00",X"FF",X"0E",X"EE",X"11",
		X"11",X"B1",X"22",X"21",X"00",X"00",X"00",X"01",X"00",X"00",X"FF",X"E0",X"EE",X"1E",X"BB",X"B1",
		X"B2",X"11",X"10",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"0E",X"11",X"1B",X"BB",X"B1",X"01",
		X"10",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"E0",X"11",X"11",X"11",X"00",X"01",X"01",X"10",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"01",X"11",X"11",X"11",X"11",X"10",X"00",X"10",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"EE",X"11",X"11",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"0E",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"10",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"01",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"0E",X"E1",X"01",X"10",X"00",X"00",X"00",X"FF",X"00",X"E1",X"11",
		X"11",X"E0",X"00",X"00",X"00",X"FF",X"0E",X"E1",X"11",X"0E",X"11",X"01",X"00",X"00",X"FF",X"0E",
		X"1D",X"D1",X"11",X"00",X"00",X"10",X"00",X"FF",X"EE",X"1D",X"1D",X"10",X"00",X"00",X"00",X"00",
		X"FF",X"EE",X"11",X"DD",X"E0",X"11",X"10",X"01",X"00",X"FF",X"EE",X"11",X"DD",X"11",X"10",X"00",
		X"11",X"00",X"FF",X"11",X"1D",X"1E",X"E1",X"10",X"00",X"00",X"00",X"FF",X"EE",X"11",X"11",X"EE",
		X"01",X"10",X"00",X"00",X"FF",X"11",X"11",X"DD",X"11",X"11",X"E1",X"00",X"11",X"FF",X"E1",X"DD",
		X"DE",X"11",X"00",X"00",X"01",X"00",X"FF",X"E1",X"11",X"1D",X"10",X"00",X"00",X"00",X"00",X"FF",
		X"E1",X"1D",X"D1",X"E1",X"11",X"01",X"00",X"00",X"FF",X"E1",X"11",X"D1",X"11",X"E1",X"EE",X"11",
		X"01",X"FF",X"1E",X"11",X"11",X"10",X"1E",X"E0",X"01",X"00",X"FF",X"EE",X"11",X"DE",X"11",X"01",
		X"00",X"00",X"00",X"FF",X"EE",X"1E",X"1D",X"11",X"00",X"01",X"01",X"00",X"FF",X"0E",X"11",X"11",
		X"E1",X"01",X"10",X"00",X"00",X"FF",X"0E",X"E1",X"D1",X"10",X"10",X"01",X"00",X"00",X"FF",X"00",
		X"E1",X"E1",X"01",X"10",X"00",X"00",X"00",X"FF",X"00",X"0E",X"EE",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"10",X"00",X"FF",X"00",
		X"00",X"10",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"01",X"00",X"00",X"FF",X"00",X"00",X"10",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"01",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"01",X"FF",X"00",X"01",X"00",X"00",X"00",X"00",X"FF",X"01",X"0E",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"E0",X"00",X"FF",X"00",X"0E",
		X"00",X"00",X"00",X"01",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"0E",X"00",X"01",
		X"00",X"00",X"FF",X"00",X"01",X"01",X"00",X"00",X"00",X"FF",X"10",X"0E",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"10",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"0D",
		X"00",X"00",X"00",X"10",X"00",X"FF",X"00",X"00",X"01",X"00",X"01",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"01",X"00",X"00",X"FF",X"00",X"00",X"10",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"09",X"00",X"00",X"00",X"00",X"00",X"FF",X"DE",X"90",X"00",X"00",X"00",X"00",X"FF",X"DD",X"E7",
		X"7E",X"D1",X"70",X"00",X"FF",X"DE",X"E1",X"77",X"EE",X"1E",X"10",X"FF",X"D7",X"77",X"EE",X"17",
		X"71",X"70",X"FF",X"DE",X"E7",X"1E",X"EE",X"1E",X"E0",X"FF",X"DD",X"7E",X"EE",X"1D",X"70",X"00",
		X"FF",X"D7",X"E0",X"00",X"00",X"00",X"00",X"FF",X"09",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"0D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"0E",X"E0",X"00",X"00",X"00",X"00",
		X"DE",X"11",X"00",X"FF",X"DE",X"EE",X"EE",X"D1",X"E0",X"1E",X"11",X"E1",X"10",X"FF",X"ED",X"E7",
		X"7E",X"77",X"EE",X"ED",X"11",X"11",X"11",X"FF",X"DE",X"E7",X"77",X"EE",X"D1",X"E1",X"1E",X"11",
		X"E1",X"FF",X"1E",X"77",X"EE",X"77",X"EE",X"1E",X"11",X"11",X"11",X"FF",X"DD",X"E7",X"7E",X"EE",
		X"E1",X"E1",X"E1",X"11",X"11",X"FF",X"EE",X"7E",X"EE",X"E1",X"D1",X"EE",X"11",X"11",X"11",X"FF",
		X"DE",X"EE",X"00",X"00",X"00",X"E1",X"E1",X"E1",X"10",X"FF",X"0D",X"E0",X"00",X"00",X"00",X"00",
		X"11",X"11",X"00",X"FF",X"0D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"E1",X"E1",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"11",X"11",X"11",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"E1",X"11",X"11",X"11",X"00",X"FF",X"00",X"E0",X"00",X"00",
		X"00",X"EE",X"E1",X"1E",X"11",X"11",X"11",X"10",X"FF",X"0E",X"EE",X"00",X"00",X"00",X"0E",X"EE",
		X"E1",X"11",X"E1",X"1E",X"E0",X"FF",X"ED",X"11",X"E0",X"00",X"00",X"EE",X"EE",X"11",X"11",X"11",
		X"11",X"11",X"FF",X"D1",X"EE",X"1E",X"1E",X"EE",X"EE",X"11",X"11",X"11",X"11",X"11",X"11",X"FF",
		X"ED",X"11",X"E1",X"EE",X"EE",X"E7",X"E7",X"71",X"1E",X"1E",X"11",X"10",X"FF",X"D1",X"E1",X"1E",
		X"EE",X"EE",X"7E",X"7E",X"EE",X"11",X"11",X"11",X"11",X"FF",X"EE",X"1E",X"E0",X"00",X"00",X"EE",
		X"11",X"11",X"11",X"11",X"EE",X"11",X"FF",X"0E",X"1E",X"00",X"00",X"00",X"0E",X"E1",X"11",X"11",
		X"11",X"11",X"10",X"FF",X"00",X"E0",X"00",X"00",X"00",X"EE",X"EE",X"E1",X"E1",X"11",X"11",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"E1",X"E1",X"11",X"10",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"EE",X"11",X"11",X"11",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"EE",X"10",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E1",X"10",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D1",X"11",X"10",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E1",X"1E",X"1E",X"11",X"11",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E1",X"11",X"1E",X"11",X"11",X"E0",X"00",X"FF",X"00",
		X"D0",X"00",X"00",X"00",X"00",X"00",X"0E",X"11",X"11",X"11",X"1E",X"11",X"00",X"FF",X"0D",X"ED",
		X"00",X"00",X"00",X"00",X"0E",X"11",X"11",X"1E",X"11",X"11",X"11",X"10",X"FF",X"DE",X"DE",X"D0",
		X"00",X"00",X"00",X"E1",X"11",X"11",X"11",X"11",X"11",X"11",X"10",X"FF",X"EE",X"1E",X"D0",X"00",
		X"00",X"0E",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"10",X"FF",X"DE",X"EE",X"EE",X"11",X"E1",
		X"EE",X"E1",X"11",X"11",X"11",X"11",X"11",X"11",X"10",X"FF",X"ED",X"E1",X"E1",X"E1",X"1E",X"11",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"00",X"FF",X"DE",X"EE",X"EE",X"1E",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"11",X"10",X"FF",X"EE",X"1E",X"D0",X"00",X"00",X"1E",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"10",X"FF",X"DE",X"ED",X"D0",X"00",X"00",X"00",X"E1",X"11",X"E1",
		X"11",X"11",X"11",X"11",X"00",X"FF",X"0D",X"ED",X"00",X"00",X"00",X"00",X"01",X"11",X"11",X"11",
		X"11",X"1E",X"10",X"00",X"FF",X"00",X"D0",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"11",X"1E",
		X"11",X"11",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"11",X"11",X"1E",X"11",
		X"10",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"10",X"E1",X"11",X"11",X"10",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"E1",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"E1",X"11",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"11",X"10",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"EE",X"EE",X"E0",X"00",X"E0",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"E1",X"EE",X"E0",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",
		X"11",X"EE",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"07",X"1E",X"70",X"E1",X"11",
		X"10",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"07",X"0E",X"71",X"11",X"11",X"E0",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"1E",X"E0",X"EE",X"1E",X"17",X"11",X"00",X"E0",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"E0",X"EE",X"11",X"11",X"7E",X"00",X"00",X"FF",X"00",X"DD",
		X"90",X"00",X"E0",X"E1",X"11",X"1E",X"11",X"11",X"E7",X"10",X"00",X"FF",X"09",X"DE",X"D9",X"00",
		X"00",X"00",X"EE",X"11",X"11",X"11",X"11",X"E0",X"00",X"FF",X"9D",X"DD",X"D9",X"90",X"D0",X"1E",
		X"E1",X"11",X"1E",X"11",X"77",X"E0",X"00",X"FF",X"9D",X"EE",X"ED",X"9D",X"77",X"EE",X"1E",X"11",
		X"11",X"11",X"11",X"10",X"00",X"FF",X"9D",X"DE",X"DE",X"DD",X"DD",X"0E",X"E7",X"11",X"11",X"11",
		X"1E",X"00",X"00",X"FF",X"9D",X"DD",X"ED",X"9D",X"D7",X"7E",X"77",X"11",X"1E",X"E1",X"10",X"00",
		X"00",X"FF",X"9D",X"ED",X"E9",X"90",X"E0",X"01",X"71",X"11",X"11",X"11",X"11",X"10",X"00",X"FF",
		X"09",X"DE",X"D9",X"00",X"00",X"77",X"11",X"11",X"11",X"11",X"7E",X"00",X"00",X"FF",X"00",X"DD",
		X"90",X"00",X"E0",X"70",X"EE",X"01",X"11",X"11",X"11",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"0E",X"17",X"11",X"1E",X"71",X"EE",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"11",
		X"01",X"11",X"11",X"71",X"01",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"70",
		X"11",X"11",X"00",X"0E",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"70",X"E7",X"E1",X"11",X"1E",
		X"10",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E1",X"11",X"1E",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"E0",X"00",X"00",X"E0",X"11",X"11",X"E0",X"0E",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"E1",X"E0",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"0E",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"E0",X"0E",X"10",X"00",X"E0",X"0E",X"00",X"00",X"FF",X"00",X"01",X"01",X"1E",X"11",X"10",
		X"00",X"00",X"00",X"FF",X"00",X"1E",X"10",X"10",X"01",X"11",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"01",X"10",X"00",X"00",X"FF",X"00",X"01",X"11",X"01",X"01",X"10",X"00",X"10",
		X"00",X"FF",X"00",X"01",X"01",X"1E",X"11",X"0E",X"01",X"00",X"00",X"FF",X"01",X"11",X"01",X"10",
		X"11",X"00",X"11",X"10",X"00",X"FF",X"00",X"00",X"E0",X"00",X"10",X"10",X"00",X"10",X"00",X"FF",
		X"E0",X"00",X"E0",X"00",X"00",X"01",X"10",X"00",X"00",X"FF",X"D0",X"00",X"00",X"E0",X"11",X"10",
		X"00",X"01",X"00",X"FF",X"01",X"01",X"11",X"10",X"00",X"10",X"11",X"00",X"00",X"FF",X"E0",X"00",
		X"E0",X"00",X"11",X"11",X"0E",X"10",X"00",X"FF",X"00",X"00",X"E0",X"11",X"11",X"E0",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"11",X"10",X"00",
		X"01",X"11",X"11",X"00",X"E0",X"FF",X"00",X"00",X"01",X"0E",X"00",X"E1",X"01",X"00",X"00",X"FF",
		X"00",X"01",X"01",X"11",X"11",X"10",X"01",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"10",X"01",
		X"10",X"00",X"00",X"FF",X"00",X"0E",X"01",X"00",X"10",X"01",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"11",X"10",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"FF",X"00",X"00",X"00",X"03",X"33",X"33",
		X"33",X"FF",X"00",X"00",X"00",X"03",X"33",X"33",X"33",X"FF",X"00",X"00",X"00",X"03",X"33",X"33",
		X"33",X"FF",X"00",X"00",X"00",X"00",X"33",X"33",X"30",X"FF",X"00",X"00",X"00",X"00",X"33",X"33",
		X"30",X"FF",X"00",X"00",X"00",X"00",X"33",X"33",X"30",X"FF",X"00",X"00",X"00",X"00",X"03",X"33",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"03",X"33",X"00",X"FF",X"00",X"00",X"00",X"00",X"03",X"33",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"30",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"22",X"22",X"20",X"00",X"FF",X"02",X"22",X"22",X"22",
		X"00",X"FF",X"22",X"22",X"22",X"22",X"20",X"FF",X"22",X"22",X"22",X"22",X"20",X"FF",X"22",X"12",
		X"22",X"22",X"20",X"FF",X"22",X"21",X"22",X"22",X"20",X"FF",X"22",X"22",X"22",X"BB",X"B0",X"FF",
		X"02",X"22",X"2B",X"B8",X"00",X"FF",X"00",X"22",X"BB",X"80",X"00",X"FF",X"00",X"02",X"2B",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"22",X"22",X"B0",X"00",X"FF",X"02",X"22",X"22",X"2B",X"00",X"FF",
		X"2B",X"B2",X"22",X"BB",X"20",X"FF",X"2B",X"BB",X"BB",X"B2",X"20",X"FF",X"22",X"BB",X"BB",X"22",
		X"20",X"FF",X"22",X"22",X"22",X"22",X"20",X"FF",X"21",X"22",X"22",X"22",X"20",X"FF",X"21",X"22",
		X"22",X"22",X"20",X"FF",X"02",X"22",X"22",X"22",X"00",X"FF",X"00",X"22",X"22",X"20",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"22",X"22",X"20",
		X"00",X"FF",X"02",X"22",X"22",X"22",X"00",X"FF",X"22",X"21",X"22",X"22",X"20",X"FF",X"22",X"21",
		X"22",X"22",X"20",X"FF",X"22",X"22",X"22",X"22",X"20",X"FF",X"22",X"2B",X"BB",X"BB",X"20",X"FF",
		X"22",X"BB",X"BB",X"BB",X"B0",X"FF",X"02",X"AB",X"22",X"22",X"00",X"FF",X"00",X"AB",X"22",X"20",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"2E",
		X"EE",X"E0",X"00",X"FF",X"0E",X"EE",X"EA",X"AA",X"00",X"FF",X"2E",X"EE",X"AC",X"CC",X"A0",X"FF",
		X"EE",X"EE",X"AC",X"CC",X"A0",X"FF",X"EE",X"EE",X"AC",X"CC",X"A0",X"FF",X"EE",X"EE",X"2A",X"AA",
		X"20",X"FF",X"2E",X"E1",X"EE",X"EE",X"20",X"FF",X"0E",X"22",X"EE",X"EE",X"00",X"FF",X"00",X"2E",
		X"EE",X"20",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"05",X"55",X"50",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"55",X"51",X"15",
		X"00",X"FF",X"00",X"00",X"00",X"05",X"04",X"55",X"55",X"11",X"50",X"FF",X"01",X"11",X"10",X"05",
		X"34",X"55",X"55",X"51",X"50",X"FF",X"11",X"00",X"11",X"15",X"04",X"55",X"55",X"55",X"50",X"FF",
		X"00",X"00",X"00",X"00",X"04",X"55",X"55",X"55",X"50",X"FF",X"00",X"00",X"00",X"00",X"00",X"55",
		X"55",X"55",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"05",X"55",X"50",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"FF",X"00",X"22",X"22",
		X"00",X"FF",X"02",X"2D",X"D2",X"20",X"FF",X"22",X"D1",X"1D",X"22",X"FF",X"22",X"2D",X"D2",X"22",
		X"FF",X"22",X"22",X"22",X"22",X"FF",X"22",X"22",X"27",X"22",X"FF",X"22",X"22",X"27",X"22",X"FF",
		X"02",X"22",X"22",X"20",X"FF",X"00",X"22",X"22",X"00",X"FF",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"02",X"22",X"22",X"AD",X"00",X"00",X"00",X"00",X"00",X"FF",X"22",X"21",X"22",
		X"AD",X"D0",X"00",X"00",X"00",X"00",X"FF",X"22",X"21",X"22",X"AD",X"DD",X"00",X"00",X"00",X"00",
		X"FF",X"22",X"22",X"22",X"44",X"44",X"44",X"40",X"00",X"00",X"FF",X"22",X"22",X"24",X"49",X"11",
		X"AA",X"A4",X"00",X"20",X"FF",X"22",X"77",X"24",X"11",X"28",X"1A",X"AA",X"40",X"20",X"FF",X"02",
		X"22",X"41",X"91",X"28",X"1A",X"AA",X"22",X"20",X"FF",X"00",X"00",X"17",X"71",X"28",X"1A",X"AA",
		X"A0",X"00",X"FF",X"00",X"09",X"77",X"88",X"11",X"AA",X"AA",X"A0",X"00",X"FF",X"00",X"09",X"88",
		X"44",X"AA",X"AA",X"AA",X"22",X"20",X"FF",X"00",X"08",X"44",X"44",X"4A",X"AA",X"AA",X"A0",X"20",
		X"FF",X"02",X"22",X"22",X"AD",X"44",X"85",X"5A",X"40",X"20",X"FF",X"22",X"21",X"22",X"AD",X"D4",
		X"48",X"54",X"00",X"00",X"FF",X"22",X"21",X"22",X"AD",X"D4",X"44",X"44",X"00",X"00",X"FF",X"22",
		X"22",X"22",X"2A",X"D4",X"44",X"40",X"00",X"00",X"FF",X"22",X"22",X"22",X"22",X"AA",X"AD",X"40",
		X"00",X"00",X"FF",X"22",X"61",X"62",X"22",X"AA",X"AD",X"D0",X"00",X"00",X"FF",X"02",X"22",X"22",
		X"22",X"AA",X"AD",X"D0",X"00",X"00",X"FF",X"00",X"00",X"00",X"22",X"22",X"2A",X"D0",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"22",X"22",X"22",X"A0",X"00",X"00",X"FF",X"00",X"00",X"00",X"22",X"61",
		X"62",X"20",X"00",X"00",X"FF",X"00",X"00",X"00",X"02",X"22",X"22",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"0D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"02",X"2D",X"DD",
		X"00",X"00",X"00",X"02",X"00",X"00",X"FF",X"22",X"2D",X"DD",X"D0",X"00",X"00",X"02",X"00",X"00",
		X"FF",X"22",X"2D",X"DD",X"4A",X"AA",X"A4",X"22",X"00",X"00",X"FF",X"22",X"22",X"21",X"11",X"AA",
		X"AA",X"24",X"00",X"00",X"FF",X"22",X"22",X"18",X"88",X"1A",X"AA",X"AA",X"40",X"00",X"FF",X"22",
		X"21",X"12",X"28",X"1A",X"AA",X"A2",X"A0",X"00",X"FF",X"02",X"19",X"12",X"28",X"1A",X"AA",X"22",
		X"A4",X"00",X"FF",X"00",X"99",X"71",X"11",X"AA",X"AA",X"22",X"A4",X"00",X"FF",X"09",X"97",X"78",
		X"8A",X"AA",X"AA",X"A2",X"A4",X"00",X"FF",X"09",X"78",X"88",X"44",X"AA",X"A5",X"AA",X"44",X"A0",
		X"FF",X"00",X"88",X"44",X"44",X"44",X"55",X"54",X"4A",X"A0",X"FF",X"02",X"2D",X"DD",X"44",X"44",
		X"44",X"44",X"4A",X"A0",X"FF",X"22",X"2D",X"DD",X"D2",X"24",X"D4",X"44",X"4A",X"A0",X"FF",X"22",
		X"2D",X"DD",X"D2",X"44",X"DD",X"D4",X"44",X"A0",X"FF",X"22",X"22",X"2D",X"D4",X"44",X"DD",X"DD",
		X"D4",X"A0",X"FF",X"22",X"22",X"22",X"24",X"44",X"DD",X"DD",X"D4",X"40",X"FF",X"22",X"61",X"62",
		X"24",X"22",X"22",X"2D",X"D4",X"00",X"FF",X"02",X"22",X"22",X"00",X"22",X"22",X"22",X"20",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"22",X"61",X"62",X"20",X"00",X"FF",X"00",X"00",X"00",X"00",X"02",
		X"22",X"22",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"AD",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"02",X"22",X"22",X"AD",X"00",X"00",X"00",X"00",X"00",X"FF",X"22",X"21",X"22",
		X"AD",X"D0",X"00",X"00",X"00",X"00",X"FF",X"22",X"21",X"22",X"AD",X"D0",X"00",X"00",X"00",X"00",
		X"FF",X"22",X"22",X"22",X"44",X"44",X"40",X"00",X"00",X"00",X"FF",X"22",X"22",X"24",X"44",X"4A",
		X"A4",X"40",X"00",X"00",X"FF",X"22",X"22",X"44",X"44",X"AA",X"AA",X"A4",X"00",X"00",X"FF",X"02",
		X"22",X"44",X"41",X"11",X"1A",X"AA",X"40",X"00",X"FF",X"00",X"00",X"41",X"19",X"91",X"21",X"AA",
		X"40",X"02",X"FF",X"00",X"01",X"11",X"99",X"91",X"21",X"AA",X"A0",X"02",X"FF",X"00",X"01",X"97",
		X"77",X"71",X"21",X"AA",X"A2",X"22",X"FF",X"00",X"08",X"88",X"AD",X"88",X"1A",X"AA",X"A0",X"00",
		X"FF",X"02",X"22",X"22",X"AD",X"AA",X"AA",X"AA",X"A0",X"00",X"FF",X"22",X"21",X"22",X"AD",X"DA",
		X"AA",X"AA",X"A2",X"22",X"FF",X"22",X"21",X"22",X"AD",X"DA",X"A5",X"55",X"40",X"02",X"FF",X"22",
		X"22",X"22",X"2A",X"D4",X"AA",X"54",X"40",X"02",X"FF",X"22",X"22",X"22",X"2A",X"D4",X"44",X"44",
		X"00",X"00",X"FF",X"22",X"61",X"62",X"24",X"44",X"D4",X"00",X"00",X"00",X"FF",X"02",X"22",X"22",
		X"AA",X"AA",X"D4",X"00",X"00",X"00",X"FF",X"00",X"02",X"22",X"AA",X"AA",X"DD",X"00",X"00",X"00",
		X"FF",X"00",X"02",X"22",X"22",X"AA",X"DD",X"00",X"00",X"00",X"FF",X"00",X"02",X"22",X"22",X"22",
		X"0D",X"00",X"00",X"00",X"FF",X"00",X"02",X"22",X"22",X"22",X"0D",X"00",X"00",X"00",X"FF",X"00",
		X"02",X"26",X"16",X"22",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"22",X"22",X"20",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"0E",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"0E",X"3E",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"0E",X"33",X"E0",X"00",X"00",X"00",X"00",X"FF",X"0E",X"EE",X"EE",X"E0",X"0E",X"33",X"3E",
		X"00",X"00",X"00",X"00",X"FF",X"EE",X"EE",X"EE",X"EE",X"0E",X"33",X"33",X"EE",X"00",X"00",X"00",
		X"FF",X"EE",X"EE",X"ED",X"EE",X"0E",X"33",X"33",X"33",X"E0",X"00",X"00",X"FF",X"EE",X"EE",X"EE",
		X"EE",X"EE",X"33",X"33",X"33",X"3E",X"00",X"00",X"FF",X"EE",X"EE",X"EE",X"EE",X"EE",X"33",X"33",
		X"33",X"33",X"E0",X"00",X"FF",X"EE",X"55",X"55",X"EE",X"EE",X"33",X"33",X"33",X"33",X"3E",X"00",
		X"FF",X"0E",X"52",X"B5",X"EE",X"EE",X"33",X"33",X"33",X"33",X"33",X"E0",X"FF",X"00",X"01",X"0E",
		X"EE",X"EE",X"33",X"33",X"33",X"33",X"D4",X"44",X"FF",X"00",X"01",X"0E",X"E5",X"5E",X"33",X"33",
		X"34",X"4D",X"D4",X"00",X"FF",X"00",X"01",X"80",X"E5",X"1E",X"33",X"44",X"DD",X"00",X"00",X"00",
		X"FF",X"00",X"01",X"28",X"00",X"14",X"4D",X"D0",X"00",X"00",X"00",X"00",X"FF",X"00",X"01",X"02",
		X"24",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"02",X"00",X"24",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"0E",X"EE",X"EE",X"E8",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"EE",X"EE",X"EE",X"EE",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"EE",X"EE",X"ED",
		X"EE",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"E0",X"00",X"00",X"00",X"00",
		X"FF",X"EE",X"9D",X"D9",X"EE",X"EE",X"DE",X"E0",X"00",X"00",X"00",X"00",X"FF",X"0E",X"EE",X"EE",
		X"EE",X"EE",X"EE",X"E0",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"0E",X"EE",X"EE",X"EE",X"E0",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"0E",X"E9",X"DD",X"9E",X"E0",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"EE",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"EE",
		X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"E3",X"33",X"3E",X"EE",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"0E",X"33",X"33",X"33",X"3E",X"EE",X"EE",X"00",X"00",X"00",X"FF",
		X"0E",X"E3",X"33",X"33",X"33",X"33",X"3E",X"EE",X"EE",X"40",X"FF",X"0E",X"EE",X"33",X"33",X"33",
		X"33",X"33",X"33",X"34",X"40",X"FF",X"0E",X"EE",X"E3",X"33",X"33",X"33",X"33",X"33",X"DD",X"00",
		X"FF",X"0E",X"EE",X"EE",X"33",X"33",X"33",X"33",X"34",X"D0",X"00",X"FF",X"0E",X"E5",X"5E",X"33",
		X"33",X"33",X"33",X"44",X"E0",X"00",X"FF",X"00",X"E5",X"1B",X"E3",X"33",X"33",X"3D",X"DE",X"E0",
		X"00",X"FF",X"00",X"00",X"80",X"0E",X"33",X"33",X"44",X"5E",X"E0",X"00",X"FF",X"00",X"00",X"20",
		X"0E",X"33",X"3D",X"4B",X"5E",X"00",X"00",X"FF",X"00",X"00",X"11",X"20",X"E3",X"4D",X"80",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"11",X"11",X"24",X"40",X"20",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"20",X"02",X"24",X"22",X"10",X"00",X"00",X"00",X"FF",X"00",X"00",X"10",X"00",X"00",X"21",X"10",
		X"00",X"00",X"00",X"FF",X"00",X"EE",X"EE",X"EE",X"00",X"00",X"20",X"00",X"00",X"00",X"FF",X"0E",
		X"EE",X"EE",X"EE",X"E0",X"00",X"10",X"00",X"00",X"00",X"FF",X"0E",X"EE",X"ED",X"EE",X"E0",X"EE",
		X"EE",X"EE",X"00",X"00",X"FF",X"0E",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"E0",X"00",X"FF",
		X"0E",X"EE",X"EE",X"EE",X"EE",X"EE",X"ED",X"EE",X"E0",X"00",X"FF",X"0E",X"E9",X"DD",X"9E",X"EE",
		X"EE",X"EE",X"EE",X"E0",X"00",X"FF",X"00",X"EE",X"EE",X"EE",X"0E",X"EE",X"EE",X"EE",X"E0",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"0E",X"E9",X"DD",X"9E",X"E0",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"EE",X"EE",X"EE",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0E",X"3E",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",
		X"3E",X"00",X"00",X"FF",X"0E",X"EE",X"EE",X"E0",X"00",X"00",X"E3",X"33",X"E0",X"00",X"FF",X"EE",
		X"EE",X"EE",X"EE",X"00",X"00",X"E3",X"33",X"E0",X"00",X"FF",X"EE",X"EE",X"ED",X"EE",X"00",X"0E",
		X"33",X"33",X"3E",X"00",X"FF",X"EE",X"EE",X"EE",X"EE",X"00",X"0E",X"33",X"33",X"3E",X"00",X"FF",
		X"EE",X"EE",X"EE",X"EE",X"E0",X"0E",X"33",X"33",X"3E",X"00",X"FF",X"EE",X"55",X"55",X"EE",X"EE",
		X"E3",X"33",X"33",X"33",X"E0",X"FF",X"0E",X"52",X"B5",X"ED",X"EE",X"E3",X"33",X"33",X"33",X"E0",
		X"FF",X"00",X"E1",X"EE",X"EE",X"EE",X"E3",X"33",X"33",X"33",X"E0",X"FF",X"00",X"E2",X"EE",X"EE",
		X"EE",X"33",X"33",X"33",X"33",X"3E",X"FF",X"00",X"E1",X"55",X"55",X"EE",X"33",X"33",X"33",X"33",
		X"3E",X"FF",X"00",X"02",X"52",X"B5",X"EE",X"33",X"33",X"33",X"33",X"3E",X"FF",X"00",X"01",X"44",
		X"44",X"DD",X"44",X"DD",X"44",X"DD",X"44",X"FF",X"00",X"02",X"21",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"0E",X"EE",X"EE",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"EE",X"EE",
		X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"EE",X"EE",X"ED",X"EE",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"EE",X"EE",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"EE",
		X"EE",X"EE",X"EE",X"E0",X"00",X"00",X"00",X"00",X"00",X"FF",X"EE",X"9D",X"D9",X"EE",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"0E",X"EE",X"EE",X"ED",X"EE",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"EE",X"EE",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"EE",X"EE",X"EE",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"EE",X"9D",X"D9",X"EE",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"0E",X"EE",X"EE",X"E0",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"02",
		X"22",X"22",X"88",X"EE",X"D0",X"00",X"00",X"00",X"00",X"00",X"FF",X"22",X"22",X"28",X"82",X"22",
		X"D0",X"00",X"00",X"00",X"00",X"00",X"FF",X"22",X"21",X"28",X"81",X"D2",X"DD",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"22",X"22",X"58",X"82",X"22",X"DD",X"00",X"00",X"00",X"00",X"00",X"FF",X"22",
		X"22",X"58",X"81",X"D2",X"DD",X"D0",X"00",X"00",X"00",X"00",X"FF",X"22",X"25",X"58",X"82",X"22",
		X"D2",X"D2",X"22",X"22",X"0A",X"B0",X"FF",X"02",X"25",X"58",X"81",X"D2",X"D2",X"2D",X"DD",X"02",
		X"2A",X"B0",X"FF",X"00",X"05",X"58",X"82",X"22",X"D2",X"22",X"2D",X"D0",X"2A",X"B0",X"FF",X"00",
		X"05",X"58",X"81",X"D2",X"D2",X"22",X"22",X"D0",X"2A",X"B0",X"FF",X"00",X"05",X"58",X"82",X"22",
		X"D4",X"44",X"42",X"D0",X"2A",X"B0",X"FF",X"00",X"05",X"58",X"81",X"D2",X"D4",X"44",X"42",X"D2",
		X"27",X"60",X"FF",X"00",X"05",X"58",X"82",X"22",X"D4",X"44",X"42",X"D0",X"07",X"60",X"FF",X"00",
		X"05",X"58",X"81",X"D2",X"D4",X"44",X"42",X"D2",X"27",X"60",X"FF",X"02",X"22",X"28",X"82",X"22",
		X"D4",X"44",X"42",X"D0",X"27",X"60",X"FF",X"22",X"22",X"28",X"81",X"D2",X"D4",X"44",X"42",X"D0",
		X"2A",X"B0",X"FF",X"22",X"21",X"22",X"88",X"EE",X"D4",X"44",X"42",X"D0",X"2A",X"B0",X"FF",X"22",
		X"22",X"22",X"22",X"2D",X"DD",X"44",X"42",X"D0",X"2A",X"B0",X"FF",X"22",X"22",X"22",X"22",X"22",
		X"DD",X"D4",X"4D",X"D2",X"2A",X"B0",X"FF",X"22",X"E1",X"1E",X"22",X"DD",X"DD",X"D2",X"22",X"22",
		X"0A",X"B0",X"FF",X"02",X"22",X"22",X"22",X"22",X"22",X"2D",X"DD",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"02",X"22",X"22",X"22",X"22",X"DD",X"00",X"00",X"00",X"FF",X"00",X"00",X"02",X"22",X"22",
		X"22",X"2D",X"D0",X"00",X"00",X"00",X"FF",X"00",X"00",X"02",X"2E",X"11",X"E2",X"20",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"22",X"22",X"22",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"02",X"22",X"28",X"8E",X"ED",X"00",X"00",X"00",X"2A",X"B0",X"FF",X"22",X"22",X"82",X"D2",
		X"DD",X"D0",X"00",X"22",X"2A",X"B0",X"FF",X"22",X"12",X"81",X"22",X"D2",X"DD",X"02",X"20",X"0A",
		X"B0",X"FF",X"22",X"22",X"82",X"22",X"D2",X"2D",X"DD",X"DD",X"0A",X"B0",X"FF",X"22",X"22",X"82",
		X"D2",X"D2",X"22",X"2D",X"DD",X"DA",X"B0",X"FF",X"22",X"25",X"81",X"22",X"D2",X"22",X"22",X"28",
		X"27",X"60",X"FF",X"02",X"25",X"82",X"22",X"D4",X"42",X"22",X"22",X"27",X"60",X"FF",X"00",X"05",
		X"82",X"D2",X"D4",X"44",X"42",X"22",X"D7",X"60",X"FF",X"00",X"05",X"81",X"22",X"D4",X"44",X"42",
		X"22",X"D7",X"60",X"FF",X"00",X"05",X"82",X"22",X"D4",X"44",X"42",X"22",X"2A",X"B0",X"FF",X"00",
		X"05",X"82",X"D2",X"D4",X"44",X"42",X"22",X"2A",X"B0",X"FF",X"00",X"05",X"81",X"22",X"D4",X"44",
		X"42",X"22",X"DA",X"B0",X"FF",X"00",X"05",X"82",X"22",X"D4",X"44",X"42",X"22",X"DA",X"B0",X"FF",
		X"02",X"22",X"82",X"D2",X"D4",X"44",X"42",X"22",X"DA",X"B0",X"FF",X"22",X"22",X"81",X"22",X"DD",
		X"D4",X"42",X"22",X"22",X"D0",X"FF",X"22",X"12",X"28",X"88",X"EE",X"DD",X"D2",X"22",X"2D",X"D0",
		X"FF",X"22",X"22",X"22",X"EE",X"EE",X"EE",X"ED",X"DD",X"DD",X"D0",X"FF",X"22",X"22",X"22",X"22",
		X"22",X"EE",X"EE",X"EE",X"EE",X"00",X"FF",X"22",X"E1",X"1E",X"22",X"22",X"22",X"22",X"22",X"EE",
		X"00",X"FF",X"02",X"22",X"22",X"22",X"22",X"22",X"22",X"2E",X"E0",X"00",X"FF",X"00",X"00",X"00",
		X"02",X"2E",X"11",X"E2",X"20",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"22",X"22",X"22",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"02",X"22",X"25",X"88",X"EE",X"D0",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"22",X"22",X"25",X"88",X"22",X"20",X"00",X"00",X"00",X"00",X"00",X"FF",X"22",X"21",
		X"55",X"88",X"1D",X"20",X"00",X"00",X"00",X"00",X"00",X"FF",X"22",X"22",X"55",X"88",X"22",X"2D",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"22",X"22",X"55",X"88",X"1D",X"2D",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"22",X"25",X"55",X"88",X"22",X"2D",X"D2",X"22",X"00",X"00",X"00",X"FF",X"02",X"25",
		X"55",X"88",X"1D",X"2D",X"2D",X"D2",X"22",X"0A",X"B0",X"FF",X"00",X"05",X"55",X"88",X"22",X"2D",
		X"22",X"2D",X"D2",X"2A",X"B0",X"FF",X"00",X"05",X"55",X"88",X"1D",X"2D",X"22",X"22",X"D0",X"2A",
		X"B0",X"FF",X"00",X"05",X"55",X"88",X"22",X"2D",X"44",X"44",X"D0",X"2A",X"B0",X"FF",X"00",X"05",
		X"55",X"88",X"1D",X"2D",X"44",X"44",X"D0",X"2A",X"B0",X"FF",X"00",X"05",X"55",X"88",X"22",X"2D",
		X"44",X"44",X"D2",X"27",X"60",X"FF",X"00",X"05",X"55",X"88",X"1D",X"2D",X"44",X"44",X"D0",X"07",
		X"60",X"FF",X"02",X"22",X"55",X"88",X"22",X"2D",X"44",X"44",X"D2",X"27",X"60",X"FF",X"22",X"22",
		X"25",X"88",X"1D",X"2D",X"44",X"44",X"D0",X"27",X"60",X"FF",X"22",X"21",X"22",X"EE",X"EE",X"DD",
		X"44",X"44",X"D0",X"2A",X"B0",X"FF",X"22",X"22",X"22",X"2E",X"EE",X"DD",X"44",X"44",X"D0",X"2A",
		X"B0",X"FF",X"22",X"22",X"22",X"22",X"2E",X"ED",X"D4",X"4D",X"D0",X"2A",X"B0",X"FF",X"22",X"E1",
		X"1E",X"22",X"2E",X"ED",X"DD",X"DD",X"D2",X"2A",X"B0",X"FF",X"02",X"22",X"22",X"22",X"EE",X"EE",
		X"D2",X"22",X"22",X"0A",X"B0",X"FF",X"00",X"02",X"22",X"2E",X"EE",X"EE",X"ED",X"D0",X"00",X"00",
		X"00",X"FF",X"00",X"02",X"22",X"2E",X"EE",X"EE",X"ED",X"00",X"00",X"00",X"00",X"FF",X"00",X"02",
		X"22",X"22",X"22",X"22",X"D0",X"00",X"00",X"00",X"00",X"FF",X"00",X"02",X"22",X"22",X"22",X"2D",
		X"D0",X"00",X"00",X"00",X"00",X"FF",X"00",X"02",X"2E",X"11",X"E2",X"20",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"22",X"22",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"02",X"22",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"22",X"22",X"22",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"22",X"22",X"12",X"20",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"22",X"22",X"12",X"22",X"22",X"00",X"00",X"00",X"00",X"00",X"FF",X"22",X"22",X"22",X"22",
		X"22",X"20",X"00",X"00",X"00",X"00",X"FF",X"26",X"9A",X"92",X"22",X"12",X"20",X"00",X"00",X"00",
		X"00",X"FF",X"26",X"A1",X"AA",X"92",X"22",X"22",X"22",X"00",X"00",X"00",X"FF",X"06",X"22",X"1A",
		X"AA",X"AA",X"AA",X"11",X"AA",X"00",X"00",X"FF",X"06",X"22",X"1A",X"A8",X"88",X"88",X"91",X"AA",
		X"00",X"00",X"FF",X"06",X"22",X"1A",X"A8",X"83",X"33",X"38",X"81",X"00",X"00",X"FF",X"06",X"22",
		X"1A",X"A8",X"83",X"77",X"78",X"81",X"18",X"00",X"FF",X"06",X"A1",X"1A",X"A8",X"83",X"77",X"78",
		X"81",X"18",X"80",X"FF",X"06",X"68",X"AA",X"A8",X"83",X"77",X"78",X"81",X"18",X"80",X"FF",X"00",
		X"66",X"89",X"A8",X"88",X"88",X"88",X"81",X"18",X"80",X"FF",X"02",X"22",X"26",X"8A",X"BB",X"BB",
		X"66",X"81",X"18",X"80",X"FF",X"22",X"22",X"22",X"68",X"AB",X"BB",X"BB",X"44",X"46",X"80",X"FF",
		X"22",X"22",X"12",X"28",X"AA",X"8B",X"B4",X"44",X"BB",X"60",X"FF",X"22",X"22",X"12",X"22",X"8A",
		X"AA",X"44",X"4B",X"BB",X"00",X"FF",X"22",X"22",X"22",X"22",X"69",X"AA",X"14",X"BB",X"B0",X"00",
		X"FF",X"22",X"22",X"22",X"22",X"26",X"9A",X"11",X"AA",X"00",X"00",X"FF",X"22",X"5E",X"52",X"22",
		X"12",X"68",X"11",X"AA",X"00",X"00",X"FF",X"02",X"22",X"22",X"22",X"22",X"26",X"81",X"AA",X"00",
		X"00",X"FF",X"00",X"00",X"22",X"22",X"22",X"22",X"68",X"AA",X"00",X"00",X"FF",X"00",X"00",X"22",
		X"5E",X"52",X"22",X"26",X"88",X"00",X"00",X"FF",X"00",X"00",X"02",X"22",X"22",X"22",X"22",X"20",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"22",X"22",X"22",X"20",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"22",X"5E",X"52",X"20",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"02",X"22",X"22",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"02",X"22",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"22",X"22",X"22",
		X"22",X"22",X"20",X"00",X"00",X"00",X"FF",X"22",X"21",X"22",X"22",X"22",X"22",X"22",X"22",X"00",
		X"FF",X"22",X"21",X"22",X"22",X"12",X"B9",X"11",X"1A",X"A0",X"FF",X"22",X"2B",X"B9",X"99",X"AA",
		X"AA",X"11",X"1A",X"A0",X"FF",X"28",X"AA",X"AA",X"AA",X"AA",X"98",X"84",X"4A",X"A0",X"FF",X"B1",
		X"AA",X"AA",X"88",X"33",X"33",X"88",X"11",X"88",X"FF",X"22",X"1A",X"AA",X"88",X"33",X"77",X"88",
		X"11",X"88",X"FF",X"22",X"1A",X"AA",X"88",X"33",X"77",X"88",X"11",X"88",X"FF",X"22",X"1A",X"AA",
		X"88",X"33",X"77",X"88",X"11",X"88",X"FF",X"22",X"1A",X"AA",X"88",X"88",X"88",X"88",X"11",X"88",
		X"FF",X"B1",X"1A",X"AA",X"88",X"66",X"6B",X"BB",X"44",X"68",X"FF",X"B9",X"AA",X"AA",X"A9",X"66",
		X"BB",X"B4",X"44",X"BB",X"FF",X"0B",X"88",X"AA",X"AA",X"AA",X"AA",X"44",X"4B",X"BB",X"FF",X"02",
		X"22",X"28",X"8A",X"AA",X"AA",X"11",X"1B",X"B0",X"FF",X"22",X"22",X"22",X"22",X"AA",X"AA",X"11",
		X"1A",X"A0",X"FF",X"22",X"21",X"22",X"22",X"22",X"AA",X"11",X"1A",X"A0",X"FF",X"22",X"21",X"22",
		X"22",X"22",X"2A",X"11",X"1A",X"A0",X"FF",X"22",X"22",X"22",X"22",X"12",X"22",X"41",X"1A",X"A0",
		X"FF",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"4A",X"A0",X"FF",X"22",X"5E",X"52",X"22",X"22",
		X"22",X"22",X"22",X"20",X"FF",X"02",X"22",X"22",X"25",X"E5",X"22",X"22",X"22",X"20",X"FF",X"00",
		X"00",X"00",X"22",X"22",X"22",X"5E",X"52",X"20",X"FF",X"00",X"00",X"00",X"00",X"00",X"02",X"22",
		X"22",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"02",X"22",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"22",X"22",X"22",X"20",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"22",X"22",X"12",X"20",X"00",X"00",X"00",X"00",X"00",X"FF",X"22",
		X"22",X"22",X"20",X"00",X"00",X"00",X"00",X"00",X"FF",X"22",X"6A",X"A2",X"22",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"2B",X"91",X"AA",X"22",X"20",X"00",X"00",X"00",X"00",X"FF",X"2B",X"22",X"1A",
		X"A2",X"20",X"00",X"00",X"00",X"00",X"FF",X"0B",X"22",X"1A",X"AA",X"20",X"00",X"00",X"00",X"00",
		X"FF",X"0B",X"22",X"1A",X"AA",X"A2",X"00",X"00",X"00",X"00",X"FF",X"0B",X"22",X"1A",X"A8",X"88",
		X"89",X"00",X"00",X"00",X"FF",X"0B",X"91",X"1A",X"A8",X"83",X"33",X"89",X"00",X"00",X"FF",X"0B",
		X"6A",X"AA",X"A8",X"87",X"73",X"38",X"90",X"00",X"FF",X"0B",X"B8",X"AA",X"A8",X"87",X"77",X"38",
		X"84",X"00",X"FF",X"00",X"B6",X"8A",X"A8",X"87",X"77",X"38",X"81",X"40",X"FF",X"02",X"22",X"28",
		X"A8",X"88",X"97",X"38",X"81",X"19",X"FF",X"22",X"22",X"22",X"AA",X"BB",X"66",X"88",X"81",X"18",
		X"FF",X"22",X"22",X"12",X"8A",X"AB",X"BB",X"B6",X"81",X"18",X"FF",X"22",X"22",X"12",X"28",X"AA",
		X"BB",X"BB",X"B4",X"18",X"FF",X"22",X"22",X"22",X"28",X"AA",X"6B",X"B4",X"44",X"48",X"FF",X"22",
		X"22",X"22",X"22",X"8A",X"A4",X"44",X"44",X"BB",X"FF",X"22",X"5E",X"52",X"22",X"8A",X"A1",X"44",
		X"BB",X"BB",X"FF",X"02",X"22",X"22",X"22",X"28",X"A1",X"1B",X"BB",X"00",X"FF",X"00",X"22",X"22",
		X"22",X"28",X"A1",X"1A",X"00",X"00",X"FF",X"00",X"22",X"22",X"22",X"22",X"81",X"1A",X"00",X"00",
		X"FF",X"00",X"22",X"5E",X"52",X"22",X"81",X"1A",X"00",X"00",X"FF",X"00",X"02",X"22",X"22",X"22",
		X"28",X"1A",X"00",X"00",X"FF",X"00",X"00",X"22",X"22",X"22",X"28",X"8A",X"00",X"00",X"FF",X"00",
		X"00",X"22",X"22",X"22",X"20",X"88",X"00",X"00",X"FF",X"00",X"00",X"22",X"5E",X"52",X"20",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"02",X"22",X"22",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"DD",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"DD",X"DD",X"EE",X"DD",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"DD",X"DD",X"EE",X"DD",X"1D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"DD",X"DD",X"66",X"66",X"11",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"6D",X"DD",X"62",X"22",X"61",X"1D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"66",X"DD",X"62",X"AA",X"21",X"11",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"06",
		X"DD",X"EE",X"DD",X"21",X"11",X"1D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"06",X"DD",
		X"EE",X"DD",X"DD",X"11",X"11",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"06",X"DD",X"EE",
		X"DD",X"12",X"D1",X"11",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"D6",X"DD",X"EE",X"DD",
		X"12",X"2D",X"11",X"10",X"08",X"D0",X"00",X"00",X"00",X"00",X"FF",X"DD",X"DD",X"EE",X"DD",X"17",
		X"66",X"66",X"66",X"28",X"D1",X"EE",X"EE",X"D0",X"00",X"FF",X"DD",X"DD",X"66",X"66",X"17",X"66",
		X"66",X"66",X"28",X"D1",X"1E",X"EE",X"DD",X"00",X"FF",X"DD",X"DD",X"62",X"22",X"61",X"8E",X"EE",
		X"EE",X"E2",X"5D",X"11",X"8E",X"D1",X"D0",X"FF",X"DD",X"DD",X"62",X"AA",X"21",X"D8",X"EE",X"EE",
		X"22",X"55",X"D1",X"18",X"D1",X"10",X"FF",X"DD",X"DD",X"EE",X"DD",X"21",X"1D",X"55",X"00",X"00",
		X"55",X"5D",X"18",X"D1",X"10",X"FF",X"6E",X"DD",X"EE",X"DD",X"D1",X"11",X"D5",X"00",X"00",X"66",
		X"55",X"D8",X"D1",X"10",X"FF",X"06",X"8E",X"EE",X"EE",X"11",X"11",X"1D",X"00",X"00",X"66",X"88",
		X"8E",X"D1",X"10",X"FF",X"00",X"66",X"66",X"68",X"81",X"11",X"11",X"D0",X"00",X"66",X"EE",X"EE",
		X"D1",X"10",X"FF",X"00",X"06",X"66",X"66",X"66",X"D1",X"11",X"10",X"00",X"66",X"EE",X"EE",X"D1",
		X"10",X"FF",X"00",X"02",X"22",X"22",X"26",X"6D",X"11",X"10",X"00",X"66",X"55",X"55",X"5D",X"10",
		X"FF",X"00",X"02",X"22",X"22",X"22",X"66",X"D1",X"10",X"00",X"65",X"50",X"00",X"55",X"D0",X"FF",
		X"00",X"02",X"22",X"22",X"22",X"26",X"6D",X"10",X"00",X"55",X"20",X"00",X"25",X"50",X"FF",X"00",
		X"02",X"2A",X"99",X"A2",X"22",X"66",X"10",X"00",X"55",X"20",X"00",X"25",X"50",X"FF",X"00",X"00",
		X"22",X"22",X"22",X"22",X"26",X"D0",X"00",X"05",X"50",X"00",X"55",X"00",X"FF",X"00",X"00",X"00",
		X"22",X"A9",X"9A",X"22",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"02",
		X"22",X"22",X"20",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"D0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"DD",X"D0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"DD",X"DD",X"EE",X"DD",X"D0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"DD",X"DD",X"EE",X"DD",X"1D",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"DD",X"DD",X"66",X"66",X"11",X"D0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"6D",X"DD",X"62",X"22",X"61",X"1D",
		X"00",X"00",X"00",X"00",X"00",X"08",X"DD",X"D0",X"00",X"FF",X"66",X"DD",X"62",X"AA",X"21",X"11",
		X"D0",X"00",X"00",X"00",X"00",X"88",X"DD",X"D1",X"00",X"FF",X"06",X"DD",X"EE",X"DD",X"21",X"11",
		X"1D",X"00",X"8D",X"10",X"08",X"88",X"DD",X"D1",X"E0",X"FF",X"06",X"DD",X"EE",X"DD",X"DD",X"11",
		X"11",X"82",X"8D",X"11",X"18",X"66",X"DD",X"D1",X"10",X"FF",X"06",X"DD",X"EE",X"DD",X"E2",X"D1",
		X"86",X"62",X"8D",X"11",X"11",X"E6",X"DD",X"D1",X"10",X"FF",X"D6",X"DD",X"EE",X"DD",X"E2",X"86",
		X"66",X"82",X"55",X"5D",X"11",X"E6",X"DD",X"D1",X"10",X"FF",X"DD",X"DD",X"EE",X"DD",X"E6",X"66",
		X"8E",X"EE",X"25",X"55",X"5D",X"E6",X"DD",X"D1",X"10",X"FF",X"DD",X"DD",X"66",X"66",X"D6",X"6E",
		X"EE",X"E0",X"00",X"00",X"55",X"68",X"DD",X"D1",X"10",X"FF",X"DD",X"DD",X"62",X"22",X"61",X"8E",
		X"E2",X"D0",X"00",X"00",X"08",X"88",X"EE",X"E1",X"10",X"FF",X"DD",X"DD",X"62",X"AA",X"21",X"D8",
		X"55",X"00",X"00",X"00",X"08",X"85",X"55",X"5D",X"10",X"FF",X"DD",X"DD",X"EE",X"DD",X"21",X"1D",
		X"55",X"00",X"00",X"00",X"08",X"55",X"00",X"55",X"D0",X"FF",X"6E",X"DD",X"EE",X"DD",X"D1",X"1D",
		X"D5",X"00",X"00",X"00",X"05",X"5E",X"00",X"05",X"80",X"FF",X"06",X"8E",X"EE",X"EE",X"11",X"1D",
		X"DD",X"00",X"00",X"00",X"05",X"EE",X"00",X"00",X"50",X"FF",X"00",X"66",X"66",X"68",X"81",X"11",
		X"DD",X"E0",X"00",X"00",X"05",X"EE",X"00",X"00",X"50",X"FF",X"00",X"06",X"66",X"66",X"66",X"D1",
		X"1D",X"E0",X"00",X"00",X"05",X"5E",X"00",X"00",X"00",X"FF",X"00",X"02",X"22",X"22",X"26",X"6D",
		X"11",X"E0",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"FF",X"00",X"02",X"22",X"22",X"22",X"66",
		X"D1",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"02",X"22",X"22",X"22",X"26",
		X"6D",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"02",X"2A",X"99",X"A2",X"22",
		X"66",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"22",X"22",X"22",X"22",
		X"26",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"22",X"A9",X"9A",
		X"22",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"02",X"22",X"22",
		X"20",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"D1",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",
		X"D1",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"88",X"D1",X"FF",
		X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"88",X"D1",X"FF",X"DD",X"D0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"88",X"D1",X"FF",X"DD",X"DD",X"EE",X"DD",
		X"D0",X"00",X"00",X"00",X"00",X"00",X"08",X"88",X"D1",X"FF",X"DD",X"DD",X"EE",X"DD",X"1D",X"00",
		X"00",X"00",X"00",X"00",X"08",X"88",X"D1",X"FF",X"DD",X"DD",X"66",X"66",X"11",X"D0",X"00",X"0D",
		X"DD",X"DD",X"68",X"88",X"D1",X"FF",X"6D",X"DD",X"62",X"22",X"61",X"1D",X"00",X"2D",X"DD",X"DD",
		X"68",X"88",X"D1",X"FF",X"66",X"DD",X"62",X"AA",X"2D",X"11",X"D6",X"2E",X"EE",X"EE",X"68",X"85",
		X"55",X"FF",X"06",X"DD",X"EE",X"DE",X"2E",X"D1",X"66",X"22",X"55",X"55",X"58",X"55",X"EE",X"FF",
		X"06",X"DD",X"EE",X"EE",X"EE",X"E6",X"66",X"E2",X"00",X"00",X"05",X"5D",X"EE",X"FF",X"06",X"DD",
		X"EE",X"EE",X"E2",X"66",X"6E",X"EE",X"00",X"00",X"05",X"DD",X"EE",X"FF",X"D6",X"DD",X"EE",X"EE",
		X"E6",X"66",X"EE",X"E0",X"00",X"00",X"05",X"DD",X"EE",X"FF",X"DD",X"DD",X"EE",X"DE",X"E6",X"6E",
		X"EE",X"10",X"00",X"00",X"05",X"DD",X"EE",X"FF",X"DD",X"DD",X"66",X"66",X"E6",X"EE",X"ED",X"10",
		X"00",X"00",X"05",X"5D",X"EE",X"FF",X"DD",X"DD",X"62",X"22",X"6E",X"8E",X"22",X"D0",X"00",X"00",
		X"00",X"55",X"EE",X"FF",X"DD",X"DD",X"62",X"AA",X"2E",X"E5",X"55",X"00",X"00",X"00",X"00",X"05",
		X"55",X"FF",X"DD",X"DD",X"EE",X"DD",X"2D",X"EE",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"6E",X"DD",X"EE",X"DD",X"D1",X"DE",X"D5",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"06",X"8E",
		X"EE",X"EE",X"11",X"1D",X"DD",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"66",X"66",X"68",
		X"81",X"11",X"D1",X"D0",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"06",X"66",X"66",X"66",X"D1",
		X"11",X"10",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"02",X"22",X"22",X"26",X"6D",X"11",X"10",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"02",X"22",X"22",X"22",X"66",X"D1",X"10",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"02",X"22",X"22",X"22",X"26",X"6D",X"10",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"02",X"2A",X"99",X"A2",X"22",X"66",X"10",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"22",X"22",X"22",X"22",X"26",X"D0",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"22",X"A9",X"9A",X"22",X"D0",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"02",
		X"22",X"22",X"20",X"D0",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"EE",X"EE",X"DD",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"DD",X"DD",X"EE",X"EE",X"ED",X"DD",X"D0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"DD",X"DD",X"E5",X"55",X"5E",X"DD",X"DD",X"DD",
		X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"DD",X"DD",X"E6",X"62",X"22",X"DD",X"DD",X"DD",
		X"D1",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"DD",X"DD",X"E6",X"6A",X"A2",X"DD",X"DD",X"DD",
		X"D1",X"10",X"00",X"00",X"00",X"00",X"00",X"FF",X"DD",X"DD",X"EE",X"EE",X"EE",X"DD",X"DD",X"DD",
		X"D1",X"1D",X"00",X"00",X"00",X"00",X"00",X"FF",X"66",X"DD",X"EE",X"EE",X"DD",X"D8",X"8E",X"DD",
		X"D1",X"1D",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"DD",X"EE",X"EE",X"DD",X"D2",X"22",X"8E",
		X"D1",X"1D",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"DD",X"EE",X"EE",X"DD",X"D2",X"22",X"22",
		X"81",X"18",X"D0",X"00",X"00",X"00",X"00",X"FF",X"00",X"DD",X"EE",X"EE",X"ED",X"D5",X"66",X"66",
		X"66",X"28",X"D1",X"EE",X"EE",X"D0",X"00",X"FF",X"00",X"DD",X"E5",X"55",X"5E",X"D5",X"66",X"66",
		X"66",X"28",X"D1",X"1E",X"EE",X"DD",X"00",X"FF",X"DD",X"DD",X"E6",X"62",X"22",X"DD",X"D8",X"88",
		X"EE",X"E2",X"5D",X"11",X"8E",X"D1",X"D0",X"FF",X"DD",X"DD",X"E6",X"6A",X"A2",X"DD",X"DD",X"DD",
		X"8E",X"22",X"55",X"D1",X"18",X"D1",X"10",X"FF",X"DD",X"DD",X"EE",X"EE",X"EE",X"DD",X"DD",X"DD",
		X"D5",X"E8",X"55",X"5D",X"18",X"D1",X"10",X"FF",X"DD",X"DD",X"EE",X"EE",X"DD",X"DD",X"DD",X"DD",
		X"D1",X"E8",X"66",X"55",X"D8",X"D1",X"10",X"FF",X"DD",X"DD",X"EE",X"EE",X"DD",X"DD",X"DD",X"DD",
		X"D1",X"DE",X"66",X"88",X"8E",X"D1",X"10",X"FF",X"DD",X"DD",X"E8",X"88",X"88",X"ED",X"DD",X"DD",
		X"D1",X"DE",X"66",X"EE",X"EE",X"D1",X"10",X"FF",X"88",X"88",X"66",X"66",X"66",X"66",X"8E",X"DD",
		X"D1",X"1D",X"66",X"EE",X"EE",X"D1",X"10",X"FF",X"00",X"00",X"86",X"22",X"22",X"26",X"66",X"66",
		X"E1",X"1D",X"66",X"55",X"55",X"5D",X"10",X"FF",X"00",X"00",X"02",X"22",X"22",X"22",X"22",X"66",
		X"66",X"1D",X"65",X"50",X"00",X"55",X"D0",X"FF",X"00",X"00",X"02",X"2A",X"99",X"A2",X"22",X"22",
		X"26",X"6D",X"55",X"20",X"00",X"25",X"50",X"FF",X"00",X"00",X"00",X"22",X"22",X"22",X"A9",X"9A",
		X"22",X"60",X"55",X"20",X"00",X"25",X"50",X"FF",X"00",X"00",X"00",X"00",X"00",X"02",X"22",X"22",
		X"20",X"00",X"05",X"50",X"00",X"55",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"EE",X"EE",X"DD",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"DD",X"DD",X"EE",X"EE",X"ED",X"DD",
		X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"DD",X"DD",X"E5",X"55",X"5E",
		X"DD",X"DD",X"DD",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"DD",X"DD",X"E6",X"62",
		X"22",X"DD",X"DD",X"DD",X"D1",X"00",X"00",X"00",X"08",X"DD",X"D0",X"00",X"FF",X"DD",X"DD",X"E6",
		X"6A",X"A2",X"DD",X"DD",X"DD",X"D1",X"10",X"00",X"00",X"88",X"DD",X"D1",X"00",X"FF",X"DD",X"DD",
		X"EE",X"EE",X"EE",X"DD",X"DD",X"DD",X"D1",X"8D",X"10",X"08",X"88",X"DD",X"D1",X"E0",X"FF",X"66",
		X"DD",X"EE",X"EE",X"DD",X"D8",X"8E",X"DD",X"62",X"8D",X"11",X"18",X"66",X"DD",X"D1",X"10",X"FF",
		X"00",X"DD",X"EE",X"EE",X"DD",X"D2",X"22",X"66",X"62",X"8D",X"11",X"11",X"E6",X"DD",X"D1",X"10",
		X"FF",X"00",X"DD",X"EE",X"EE",X"DD",X"D2",X"66",X"66",X"82",X"55",X"5D",X"11",X"E6",X"DD",X"D1",
		X"10",X"FF",X"00",X"DD",X"EE",X"EE",X"ED",X"D5",X"66",X"6E",X"EE",X"25",X"55",X"5D",X"E6",X"DD",
		X"D1",X"10",X"FF",X"00",X"DD",X"E5",X"55",X"5E",X"D5",X"6E",X"EE",X"E2",X"28",X"00",X"55",X"68",
		X"DD",X"D1",X"10",X"FF",X"DD",X"DD",X"E6",X"62",X"22",X"DD",X"D8",X"85",X"55",X"58",X"00",X"08",
		X"88",X"EE",X"E1",X"10",X"FF",X"DD",X"DD",X"E6",X"6A",X"A2",X"DD",X"DD",X"DD",X"55",X"58",X"00",
		X"08",X"85",X"55",X"5D",X"10",X"FF",X"DD",X"DD",X"EE",X"EE",X"EE",X"DD",X"DD",X"DD",X"D5",X"58",
		X"00",X"08",X"55",X"00",X"55",X"D0",X"FF",X"DD",X"DD",X"EE",X"EE",X"DD",X"DD",X"DD",X"DD",X"DE",
		X"58",X"00",X"05",X"5E",X"00",X"05",X"80",X"FF",X"DD",X"DD",X"EE",X"EE",X"DD",X"DD",X"DD",X"DD",
		X"DE",X"E8",X"00",X"05",X"EE",X"00",X"00",X"50",X"FF",X"DD",X"DD",X"E8",X"88",X"88",X"ED",X"DD",
		X"DD",X"DD",X"EE",X"00",X"05",X"EE",X"00",X"00",X"50",X"FF",X"88",X"88",X"66",X"66",X"66",X"66",
		X"8E",X"DD",X"D1",X"DE",X"00",X"05",X"5E",X"00",X"00",X"00",X"FF",X"00",X"00",X"86",X"22",X"22",
		X"26",X"66",X"66",X"E1",X"1D",X"00",X"00",X"55",X"00",X"00",X"00",X"FF",X"00",X"00",X"02",X"22",
		X"22",X"22",X"22",X"66",X"66",X"1D",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"02",
		X"2A",X"99",X"A2",X"22",X"22",X"26",X"6D",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"22",X"22",X"22",X"A9",X"9A",X"22",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"02",X"22",X"22",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"D1",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"D1",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"88",X"D1",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"88",X"D1",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"88",X"D1",X"FF",X"00",X"00",X"EE",X"EE",X"DD",X"00",
		X"00",X"00",X"00",X"00",X"00",X"08",X"88",X"D1",X"FF",X"DD",X"DD",X"EE",X"EE",X"ED",X"DD",X"D0",
		X"00",X"00",X"00",X"00",X"08",X"88",X"D1",X"FF",X"DD",X"DD",X"E5",X"55",X"5E",X"DD",X"DD",X"DD",
		X"DD",X"DD",X"DD",X"68",X"88",X"D1",X"FF",X"DD",X"DD",X"E6",X"62",X"22",X"EE",X"ED",X"DD",X"2D",
		X"DD",X"DD",X"68",X"88",X"D1",X"FF",X"DD",X"DD",X"E6",X"6A",X"A2",X"EE",X"EE",X"E6",X"2E",X"EE",
		X"EE",X"68",X"85",X"55",X"FF",X"DD",X"DD",X"EE",X"EE",X"EE",X"EE",X"EE",X"66",X"22",X"55",X"55",
		X"58",X"55",X"EE",X"FF",X"66",X"DD",X"EE",X"EE",X"DE",X"E8",X"86",X"66",X"E2",X"1D",X"00",X"05",
		X"5D",X"EE",X"FF",X"00",X"DD",X"EE",X"EE",X"DE",X"E2",X"66",X"6E",X"EE",X"1D",X"00",X"05",X"DD",
		X"EE",X"FF",X"00",X"DD",X"EE",X"EE",X"DE",X"E5",X"66",X"EE",X"ED",X"1D",X"00",X"05",X"DD",X"EE",
		X"FF",X"00",X"DD",X"EE",X"EE",X"EE",X"E5",X"6E",X"EE",X"26",X"1D",X"00",X"05",X"DD",X"EE",X"FF",
		X"00",X"DD",X"E5",X"55",X"5E",X"E5",X"8E",X"E2",X"22",X"2D",X"00",X"05",X"5D",X"EE",X"FF",X"DD",
		X"DD",X"E6",X"62",X"22",X"EE",X"E8",X"55",X"55",X"5D",X"00",X"00",X"55",X"EE",X"FF",X"DD",X"DD",
		X"E6",X"6A",X"A2",X"EE",X"EE",X"EE",X"55",X"5D",X"00",X"00",X"05",X"55",X"FF",X"DD",X"DD",X"EE",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"E5",X"5D",X"00",X"00",X"00",X"00",X"FF",X"DD",X"DD",X"EE",X"EE",
		X"DD",X"DE",X"EE",X"EE",X"EE",X"5D",X"00",X"00",X"00",X"00",X"FF",X"DD",X"DD",X"EE",X"EE",X"DD",
		X"DD",X"DD",X"EE",X"EE",X"DD",X"00",X"00",X"00",X"00",X"FF",X"DD",X"DD",X"E8",X"88",X"88",X"ED",
		X"DD",X"DD",X"EE",X"1D",X"00",X"00",X"00",X"00",X"FF",X"88",X"88",X"66",X"66",X"66",X"66",X"8E",
		X"DD",X"DD",X"1D",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"86",X"22",X"22",X"26",X"66",X"66",
		X"E1",X"1D",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"02",X"22",X"22",X"22",X"22",X"66",X"66",
		X"1D",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"02",X"2A",X"99",X"A2",X"22",X"22",X"26",X"6D",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"22",X"22",X"22",X"A9",X"9A",X"22",X"60",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"02",X"22",X"22",X"20",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"1E",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"1E",X"E1",X"D0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"1E",X"E1",X"11",X"D0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"1E",X"E6",X"61",X"11",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"2E",X"E2",X"22",X"E1",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"2E",X"E2",X"AA",X"21",X"ED",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"2E",X"E1",X"E2",X"21",X"ED",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"2E",X"E1",
		X"11",X"81",X"ED",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"2E",X"E1",X"11",X"11",
		X"ED",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"1E",X"E1",X"11",X"11",X"2D",X"D0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"1E",X"E1",X"11",X"11",X"2E",X"DD",X"00",X"00",
		X"8D",X"00",X"00",X"00",X"00",X"FF",X"1E",X"E6",X"61",X"11",X"56",X"66",X"66",X"62",X"8D",X"1E",
		X"EE",X"ED",X"00",X"FF",X"1E",X"E2",X"22",X"E1",X"56",X"66",X"66",X"62",X"8D",X"11",X"EE",X"ED",
		X"D0",X"FF",X"1E",X"E2",X"AA",X"21",X"E8",X"EE",X"EE",X"EE",X"25",X"D1",X"18",X"ED",X"1D",X"FF",
		X"6E",X"E1",X"E2",X"21",X"E8",X"EE",X"EE",X"E2",X"25",X"5D",X"11",X"8D",X"11",X"FF",X"6E",X"E1",
		X"11",X"81",X"EE",X"28",X"00",X"00",X"05",X"55",X"D1",X"8D",X"11",X"FF",X"66",X"E1",X"11",X"11",
		X"ED",X"22",X"00",X"00",X"06",X"65",X"5D",X"8D",X"11",X"FF",X"06",X"66",X"61",X"11",X"ED",X"E2",
		X"00",X"00",X"06",X"68",X"88",X"ED",X"11",X"FF",X"00",X"66",X"66",X"61",X"ED",X"E2",X"00",X"00",
		X"06",X"6E",X"EE",X"ED",X"11",X"FF",X"02",X"22",X"26",X"66",X"ED",X"E2",X"00",X"00",X"06",X"6E",
		X"EE",X"ED",X"11",X"FF",X"02",X"22",X"22",X"26",X"6D",X"D8",X"00",X"00",X"06",X"65",X"55",X"55",
		X"D1",X"FF",X"02",X"22",X"22",X"22",X"66",X"D8",X"00",X"00",X"06",X"55",X"00",X"05",X"5D",X"FF",
		X"02",X"22",X"22",X"22",X"66",X"D8",X"00",X"00",X"05",X"52",X"00",X"02",X"55",X"FF",X"02",X"22",
		X"22",X"22",X"26",X"6D",X"00",X"00",X"05",X"52",X"00",X"02",X"55",X"FF",X"02",X"2A",X"99",X"A2",
		X"26",X"6D",X"00",X"00",X"00",X"55",X"00",X"05",X"50",X"FF",X"00",X"22",X"22",X"22",X"22",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"22",X"A9",X"9A",X"22",X"60",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"02",X"22",X"22",X"26",X"60",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"1E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"1E",X"E1",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"1E",X"E1",X"11",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"1E",X"E6",X"61",X"11",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"2E",X"E2",X"22",X"E1",X"E0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"2E",X"E2",X"AA",X"21",X"ED",X"00",X"00",X"00",
		X"00",X"00",X"00",X"8D",X"DD",X"00",X"FF",X"2E",X"E1",X"E2",X"21",X"ED",X"00",X"00",X"00",X"00",
		X"00",X"08",X"8D",X"DD",X"10",X"FF",X"2E",X"E1",X"11",X"81",X"ED",X"D0",X"00",X"08",X"D1",X"00",
		X"88",X"8D",X"DD",X"1E",X"FF",X"2E",X"E1",X"11",X"11",X"ED",X"D0",X"08",X"28",X"D1",X"11",X"86",
		X"6D",X"DD",X"11",X"FF",X"1E",X"E1",X"11",X"11",X"2D",X"D8",X"66",X"28",X"D1",X"11",X"1E",X"6D",
		X"DD",X"11",X"FF",X"1E",X"E1",X"11",X"11",X"28",X"66",X"68",X"25",X"55",X"D1",X"1E",X"6D",X"DD",
		X"11",X"FF",X"1E",X"E6",X"61",X"11",X"56",X"68",X"EE",X"E2",X"55",X"55",X"DE",X"6D",X"DD",X"11",
		X"FF",X"1E",X"E2",X"22",X"E1",X"56",X"EE",X"EE",X"00",X"00",X"05",X"56",X"8D",X"DD",X"11",X"FF",
		X"1E",X"E2",X"AA",X"21",X"E8",X"EE",X"00",X"00",X"00",X"00",X"88",X"8E",X"EE",X"11",X"FF",X"8E",
		X"E1",X"E2",X"21",X"E8",X"28",X"00",X"00",X"00",X"00",X"88",X"55",X"55",X"D1",X"FF",X"6E",X"E1",
		X"11",X"81",X"EE",X"28",X"00",X"00",X"00",X"00",X"85",X"50",X"05",X"5D",X"FF",X"66",X"E1",X"11",
		X"11",X"EE",X"22",X"00",X"00",X"00",X"00",X"55",X"E0",X"00",X"58",X"FF",X"06",X"66",X"61",X"11",
		X"ED",X"82",X"00",X"00",X"00",X"00",X"5E",X"E0",X"00",X"05",X"FF",X"00",X"66",X"66",X"61",X"ED",
		X"82",X"00",X"00",X"00",X"00",X"5E",X"E0",X"00",X"05",X"FF",X"02",X"22",X"26",X"66",X"ED",X"82",
		X"00",X"00",X"00",X"00",X"55",X"E0",X"00",X"00",X"FF",X"02",X"22",X"22",X"26",X"6D",X"E8",X"00",
		X"00",X"00",X"00",X"05",X"50",X"00",X"00",X"FF",X"02",X"22",X"22",X"22",X"66",X"D8",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"02",X"22",X"22",X"22",X"66",X"DE",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"02",X"22",X"22",X"22",X"26",X"6D",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"02",X"2A",X"99",X"A2",X"26",X"6D",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"22",X"22",X"22",X"22",X"60",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"22",X"A9",X"9A",X"22",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"02",X"22",X"22",X"26",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"D1",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"D1",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"88",X"D1",X"FF",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"88",X"D1",X"FF",X"1E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",
		X"88",X"D1",X"FF",X"1E",X"E1",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"88",X"D1",
		X"FF",X"1E",X"E1",X"11",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"88",X"D1",X"FF",X"1E",
		X"E6",X"61",X"11",X"E0",X"00",X"00",X"0D",X"DD",X"DD",X"68",X"88",X"D1",X"FF",X"2E",X"E2",X"22",
		X"E1",X"E0",X"00",X"00",X"2D",X"DD",X"DD",X"68",X"88",X"D1",X"FF",X"2E",X"E2",X"AA",X"21",X"ED",
		X"00",X"06",X"2E",X"EE",X"EE",X"68",X"85",X"55",X"FF",X"2E",X"E1",X"E2",X"21",X"ED",X"00",X"66",
		X"22",X"55",X"55",X"58",X"55",X"EE",X"FF",X"2E",X"E1",X"11",X"81",X"ED",X"D6",X"66",X"E2",X"00",
		X"00",X"05",X"5D",X"EE",X"FF",X"2E",X"E1",X"11",X"EE",X"EE",X"66",X"6E",X"EE",X"00",X"00",X"05",
		X"DD",X"EE",X"FF",X"1E",X"E1",X"11",X"EE",X"26",X"66",X"EE",X"E0",X"00",X"00",X"05",X"DD",X"EE",
		X"FF",X"1E",X"E1",X"11",X"EE",X"56",X"6E",X"EE",X"00",X"00",X"00",X"05",X"DD",X"EE",X"FF",X"1E",
		X"E6",X"61",X"1E",X"56",X"EE",X"E0",X"00",X"00",X"00",X"05",X"5D",X"EE",X"FF",X"1E",X"E2",X"22",
		X"E1",X"5E",X"EE",X"00",X"00",X"00",X"00",X"00",X"55",X"EE",X"FF",X"1E",X"E2",X"AA",X"21",X"E8",
		X"ED",X"00",X"00",X"00",X"00",X"00",X"05",X"55",X"FF",X"8E",X"E1",X"E2",X"21",X"E8",X"2D",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"6E",X"E1",X"11",X"81",X"E8",X"2E",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"66",X"E1",X"11",X"11",X"E8",X"22",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"06",X"66",X"61",X"11",X"E8",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"66",X"66",X"61",X"EE",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"02",
		X"22",X"26",X"66",X"ED",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"02",X"22",X"22",
		X"26",X"6D",X"ED",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"02",X"22",X"22",X"22",X"66",
		X"DD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"02",X"22",X"22",X"22",X"66",X"DD",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"02",X"22",X"22",X"22",X"26",X"6D",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"02",X"2A",X"99",X"A2",X"26",X"6D",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"22",X"22",X"22",X"22",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"22",X"A9",X"9A",X"22",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"02",X"22",X"22",X"26",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"11",X"10",X"00",X"FF",X"00",X"01",
		X"B1",X"EE",X"11",X"00",X"FF",X"09",X"B1",X"CB",X"EE",X"19",X"10",X"FF",X"0E",X"9C",X"CC",X"BE",
		X"C9",X"91",X"FF",X"E9",X"9C",X"CC",X"CC",X"C9",X"99",X"FF",X"99",X"EC",X"E9",X"99",X"C9",X"99",
		X"FF",X"78",X"CE",X"EE",X"99",X"3C",X"EE",X"FF",X"67",X"77",X"EE",X"EE",X"37",X"E7",X"FF",X"66",
		X"67",X"EE",X"E8",X"67",X"50",X"FF",X"55",X"62",X"7E",X"86",X"66",X"50",X"FF",X"05",X"52",X"27",
		X"26",X"55",X"00",X"FF",X"00",X"55",X"26",X"55",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"56",X"67",X"EE",X"00",X"00",X"FF",X"05",X"56",X"6E",X"EE",X"B3",X"00",X"FF",X"55",X"66",
		X"7C",X"EE",X"BB",X"00",X"FF",X"52",X"27",X"77",X"CC",X"CB",X"90",X"FF",X"22",X"77",X"77",X"7C",
		X"B1",X"30",X"FF",X"67",X"77",X"77",X"7C",X"B9",X"90",X"FF",X"52",X"87",X"77",X"EC",X"99",X"99",
		X"FF",X"56",X"68",X"7E",X"EC",X"BB",X"BB",X"FF",X"05",X"66",X"33",X"CC",X"C1",X"1B",X"FF",X"05",
		X"67",X"7C",X"99",X"B1",X"B0",X"FF",X"00",X"55",X"EE",X"99",X"B1",X"00",X"FF",X"00",X"00",X"7E",
		X"9B",X"10",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"77",X"26",X"55",X"00",X"00",X"FF",
		X"07",X"62",X"27",X"66",X"55",X"00",X"FF",X"46",X"62",X"7E",X"86",X"66",X"50",X"FF",X"66",X"6E",
		X"EE",X"E8",X"66",X"50",X"FF",X"44",X"6E",X"EE",X"EE",X"36",X"65",X"FF",X"EE",X"CE",X"EE",X"EE",
		X"3C",X"C6",X"FF",X"EE",X"EC",X"EE",X"EE",X"C9",X"99",X"FF",X"EE",X"EC",X"C9",X"9C",X"C9",X"99",
		X"FF",X"0E",X"EC",X"B9",X"9B",X"99",X"91",X"FF",X"0E",X"E1",X"99",X"99",X"19",X"10",X"FF",X"00",
		X"01",X"B1",X"BB",X"11",X"00",X"FF",X"00",X"00",X"00",X"11",X"10",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"0E",X"EC",X"75",X"50",
		X"00",X"FF",X"00",X"EE",X"CC",X"C2",X"25",X"00",X"FF",X"01",X"CC",X"C4",X"77",X"86",X"60",X"FF",
		X"03",X"CC",X"47",X"77",X"78",X"55",X"FF",X"3B",X"9C",X"47",X"77",X"75",X"55",X"FF",X"BB",X"BC",
		X"C1",X"77",X"72",X"65",X"FF",X"9B",X"BE",X"9C",X"97",X"26",X"66",X"FF",X"99",X"99",X"9C",X"78",
		X"66",X"65",X"FF",X"B9",X"9C",X"C7",X"77",X"76",X"50",X"FF",X"39",X"9C",X"77",X"77",X"86",X"50",
		X"FF",X"03",X"39",X"47",X"78",X"65",X"50",X"FF",X"00",X"09",X"44",X"46",X"55",X"00",X"FF",X"00",
		X"00",X"47",X"65",X"50",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"01",X"99",X"E7",X"00",
		X"00",X"FF",X"00",X"19",X"99",X"EE",X"55",X"00",X"FF",X"01",X"99",X"99",X"C7",X"76",X"50",X"FF",
		X"11",X"1C",X"4C",X"33",X"66",X"50",X"FF",X"19",X"BB",X"CB",X"EE",X"86",X"65",X"FF",X"1B",X"99",
		X"9E",X"EE",X"E8",X"25",X"FF",X"01",X"99",X"CE",X"EE",X"EE",X"76",X"FF",X"0B",X"B9",X"CE",X"EE",
		X"E7",X"22",X"FF",X"01",X"1C",X"9C",X"EE",X"E2",X"25",X"FF",X"00",X"EE",X"EE",X"C7",X"66",X"55",
		X"FF",X"00",X"EE",X"EE",X"E6",X"65",X"50",X"FF",X"00",X"00",X"EE",X"76",X"65",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"DD",X"E0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"DD",X"DD",X"EE",X"DD",X"D0",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"DD",X"DD",X"EE",X"DD",X"1D",X"00",X"00",X"00",X"00",X"00",X"FF",X"DD",X"DD",X"66",
		X"66",X"11",X"D0",X"00",X"00",X"00",X"00",X"FF",X"6D",X"DD",X"62",X"22",X"61",X"1D",X"00",X"00",
		X"00",X"00",X"FF",X"66",X"DD",X"62",X"AA",X"21",X"11",X"D0",X"00",X"00",X"00",X"FF",X"06",X"DD",
		X"EE",X"DD",X"21",X"EE",X"ED",X"00",X"00",X"00",X"FF",X"06",X"DD",X"EE",X"DD",X"D1",X"EE",X"EE",
		X"D0",X"00",X"00",X"FF",X"06",X"DD",X"EE",X"DD",X"11",X"EE",X"EE",X"DD",X"00",X"00",X"FF",X"D6",
		X"DD",X"EE",X"DD",X"11",X"EE",X"EE",X"DD",X"B0",X"00",X"FF",X"DD",X"DD",X"EE",X"DD",X"11",X"EE",
		X"EE",X"DD",X"B1",X"00",X"FF",X"DD",X"DD",X"66",X"66",X"11",X"EE",X"EE",X"DD",X"B1",X"10",X"FF",
		X"DD",X"DD",X"62",X"22",X"61",X"88",X"8E",X"DD",X"B1",X"10",X"FF",X"DD",X"DD",X"62",X"AA",X"21",
		X"58",X"88",X"8D",X"B1",X"10",X"FF",X"DD",X"DD",X"EE",X"DD",X"21",X"15",X"88",X"88",X"B1",X"10",
		X"FF",X"6E",X"DD",X"EE",X"DD",X"D1",X"11",X"53",X"33",X"3D",X"10",X"FF",X"06",X"8E",X"EE",X"EE",
		X"11",X"11",X"13",X"88",X"88",X"D0",X"FF",X"00",X"66",X"66",X"68",X"81",X"11",X"1B",X"58",X"88",
		X"80",X"FF",X"00",X"06",X"66",X"66",X"66",X"D1",X"1B",X"11",X"00",X"00",X"FF",X"00",X"02",X"22",
		X"22",X"26",X"6D",X"1B",X"11",X"00",X"00",X"FF",X"00",X"02",X"22",X"22",X"22",X"66",X"DB",X"11",
		X"00",X"00",X"FF",X"00",X"02",X"22",X"22",X"22",X"23",X"33",X"11",X"00",X"00",X"FF",X"00",X"02",
		X"2A",X"99",X"A2",X"22",X"66",X"D1",X"00",X"00",X"FF",X"00",X"00",X"22",X"22",X"22",X"22",X"28",
		X"8D",X"00",X"00",X"FF",X"00",X"00",X"00",X"22",X"A9",X"9A",X"22",X"8D",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"02",X"22",X"22",X"20",X"0D",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"EE",X"EE",X"DD",X"E0",X"00",X"00",X"00",X"00",X"FF",X"DD",X"DD",X"EE",X"EE",X"DD",
		X"DD",X"DD",X"00",X"00",X"00",X"FF",X"DD",X"DD",X"EE",X"EE",X"ED",X"DD",X"DD",X"AB",X"D0",X"00",
		X"FF",X"DD",X"DD",X"55",X"55",X"ED",X"DD",X"DD",X"AB",X"DD",X"00",X"FF",X"DD",X"DD",X"66",X"22",
		X"2D",X"DE",X"ED",X"AB",X"DD",X"10",X"FF",X"DD",X"DD",X"66",X"AA",X"2D",X"EE",X"ED",X"11",X"BD",
		X"D1",X"FF",X"66",X"DD",X"EE",X"EE",X"DD",X"EE",X"ED",X"11",X"BB",X"11",X"FF",X"00",X"DD",X"EE",
		X"EE",X"DD",X"EE",X"ED",X"11",X"BB",X"11",X"FF",X"00",X"DD",X"EE",X"EE",X"DD",X"EE",X"ED",X"11",
		X"BB",X"11",X"FF",X"00",X"DD",X"EE",X"EE",X"DD",X"EE",X"ED",X"D1",X"BB",X"11",X"FF",X"00",X"DD",
		X"EE",X"EE",X"ED",X"E8",X"66",X"66",X"BB",X"11",X"FF",X"DD",X"DD",X"55",X"55",X"ED",X"E6",X"66",
		X"6A",X"A6",X"61",X"FF",X"DD",X"DD",X"66",X"22",X"2D",X"DD",X"DD",X"AA",X"66",X"61",X"FF",X"DD",
		X"DD",X"66",X"AA",X"2D",X"DD",X"DD",X"AB",X"E6",X"11",X"FF",X"DD",X"DD",X"EE",X"EE",X"ED",X"DD",
		X"DD",X"AB",X"DD",X"11",X"FF",X"DD",X"DD",X"EE",X"EE",X"DD",X"DD",X"DD",X"AB",X"DD",X"11",X"FF",
		X"DD",X"DD",X"E8",X"88",X"88",X"ED",X"DD",X"AB",X"DD",X"11",X"FF",X"88",X"88",X"66",X"66",X"66",
		X"66",X"8E",X"AB",X"DD",X"11",X"FF",X"00",X"00",X"86",X"22",X"22",X"26",X"6A",X"B6",X"ED",X"11",
		X"FF",X"00",X"00",X"02",X"22",X"22",X"22",X"22",X"66",X"66",X"11",X"FF",X"00",X"00",X"02",X"2A",
		X"99",X"A2",X"22",X"22",X"26",X"61",X"FF",X"00",X"00",X"00",X"22",X"22",X"22",X"A9",X"9A",X"22",
		X"60",X"FF",X"00",X"00",X"00",X"00",X"00",X"02",X"22",X"22",X"20",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"1E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"1E",X"E1",X"D0",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"1E",X"E1",X"11",X"D0",X"00",X"00",X"00",X"00",X"FF",X"1E",X"66",
		X"11",X"11",X"E0",X"00",X"00",X"00",X"FF",X"2E",X"22",X"2E",X"11",X"E0",X"00",X"00",X"00",X"FF",
		X"2E",X"2A",X"A2",X"11",X"ED",X"00",X"00",X"00",X"FF",X"2E",X"EE",X"22",X"11",X"ED",X"00",X"00",
		X"00",X"FF",X"2E",X"E1",X"18",X"11",X"ED",X"D0",X"00",X"00",X"FF",X"2E",X"E1",X"11",X"11",X"E1",
		X"11",X"00",X"00",X"FF",X"1E",X"E1",X"11",X"11",X"E1",X"11",X"E0",X"00",X"FF",X"1E",X"66",X"11",
		X"11",X"E1",X"11",X"DA",X"00",X"FF",X"1E",X"22",X"2E",X"11",X"E1",X"11",X"DB",X"00",X"FF",X"1E",
		X"2A",X"A2",X"11",X"E1",X"11",X"DB",X"E0",X"FF",X"1E",X"EE",X"22",X"11",X"E1",X"11",X"DB",X"E0",
		X"FF",X"6E",X"E1",X"18",X"11",X"E8",X"88",X"DB",X"E0",X"FF",X"6E",X"E1",X"11",X"11",X"E5",X"88",
		X"8B",X"E0",X"FF",X"66",X"E1",X"11",X"11",X"EE",X"6A",X"AA",X"E0",X"FF",X"06",X"66",X"61",X"11",
		X"ED",X"AA",X"88",X"E0",X"FF",X"00",X"66",X"66",X"61",X"ED",X"B5",X"88",X"80",X"FF",X"02",X"22",
		X"26",X"66",X"ED",X"BE",X"00",X"00",X"FF",X"02",X"22",X"22",X"26",X"6D",X"BE",X"00",X"00",X"FF",
		X"02",X"22",X"22",X"22",X"66",X"BE",X"00",X"00",X"FF",X"02",X"22",X"22",X"22",X"66",X"BE",X"00",
		X"00",X"FF",X"02",X"22",X"22",X"22",X"2B",X"BE",X"00",X"00",X"FF",X"02",X"2A",X"99",X"A2",X"26",
		X"6E",X"00",X"00",X"FF",X"00",X"22",X"22",X"22",X"22",X"6E",X"00",X"00",X"FF",X"00",X"22",X"A9",
		X"9A",X"22",X"60",X"00",X"00",X"FF",X"00",X"02",X"22",X"22",X"29",X"60",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"06",X"D0",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"06",X"D0",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"06",X"D0",X"00",X"00",X"FF",X"02",X"22",X"22",X"00",X"06",X"DD",X"00",X"00",X"FF",X"22",X"22",
		X"22",X"20",X"06",X"DD",X"00",X"00",X"FF",X"22",X"22",X"22",X"21",X"11",X"11",X"00",X"00",X"FF",
		X"22",X"22",X"22",X"21",X"22",X"11",X"10",X"00",X"FF",X"22",X"69",X"62",X"21",X"82",X"11",X"11",
		X"00",X"FF",X"02",X"29",X"22",X"01",X"88",X"11",X"11",X"10",X"FF",X"00",X"09",X"90",X"01",X"11",
		X"11",X"11",X"11",X"FF",X"00",X"09",X"99",X"07",X"66",X"66",X"11",X"11",X"FF",X"00",X"09",X"09",
		X"91",X"11",X"11",X"6E",X"11",X"FF",X"00",X"09",X"09",X"91",X"22",X"11",X"16",X"81",X"FF",X"00",
		X"09",X"99",X"01",X"82",X"11",X"11",X"00",X"FF",X"00",X"09",X"90",X"01",X"88",X"11",X"11",X"10",
		X"FF",X"02",X"22",X"22",X"01",X"11",X"11",X"11",X"11",X"FF",X"22",X"22",X"22",X"27",X"66",X"66",
		X"11",X"11",X"FF",X"22",X"22",X"22",X"29",X"06",X"DD",X"6E",X"11",X"FF",X"22",X"22",X"22",X"22",
		X"26",X"DD",X"D6",X"81",X"FF",X"22",X"E1",X"E2",X"22",X"26",X"DD",X"D0",X"00",X"FF",X"02",X"22",
		X"22",X"22",X"26",X"DD",X"00",X"00",X"FF",X"00",X"00",X"22",X"22",X"26",X"DD",X"00",X"00",X"FF",
		X"00",X"00",X"22",X"E1",X"E6",X"DD",X"00",X"00",X"FF",X"00",X"00",X"02",X"22",X"26",X"D0",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"06",X"D0",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"6E",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"6E",X"E0",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"6E",X"E0",X"00",X"00",X"FF",X"02",X"22",X"22",X"00",X"6E",X"EE",X"00",X"00",
		X"FF",X"22",X"22",X"22",X"20",X"6E",X"EE",X"00",X"00",X"FF",X"22",X"22",X"22",X"DD",X"D1",X"EE",
		X"00",X"00",X"FF",X"22",X"22",X"22",X"D2",X"D1",X"11",X"10",X"00",X"FF",X"22",X"69",X"62",X"D2",
		X"D1",X"11",X"11",X"10",X"FF",X"02",X"29",X"22",X"D2",X"D1",X"11",X"11",X"10",X"FF",X"00",X"09",
		X"90",X"DD",X"D1",X"11",X"11",X"10",X"FF",X"00",X"09",X"90",X"76",X"66",X"8E",X"11",X"10",X"FF",
		X"00",X"09",X"99",X"DD",X"D1",X"90",X"00",X"00",X"FF",X"00",X"09",X"99",X"D2",X"D1",X"11",X"10",
		X"00",X"FF",X"00",X"09",X"90",X"D2",X"D1",X"11",X"11",X"10",X"FF",X"00",X"09",X"90",X"D8",X"D1",
		X"11",X"11",X"10",X"FF",X"02",X"22",X"22",X"DD",X"D1",X"11",X"11",X"10",X"FF",X"22",X"22",X"22",
		X"26",X"6E",X"EE",X"11",X"10",X"FF",X"22",X"22",X"22",X"22",X"6E",X"EE",X"20",X"00",X"FF",X"22",
		X"22",X"22",X"22",X"6E",X"EE",X"20",X"00",X"FF",X"22",X"E1",X"E2",X"22",X"6E",X"EE",X"20",X"00",
		X"FF",X"02",X"22",X"22",X"22",X"6E",X"E2",X"20",X"00",X"FF",X"00",X"00",X"00",X"02",X"6E",X"E2",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"6E",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"6D",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"6D",X"00",X"00",X"FF",
		X"02",X"22",X"22",X"00",X"00",X"6D",X"00",X"00",X"FF",X"22",X"22",X"22",X"20",X"00",X"6D",X"D0",
		X"00",X"FF",X"22",X"22",X"22",X"20",X"00",X"6D",X"D0",X"00",X"FF",X"22",X"22",X"22",X"22",X"11",
		X"11",X"10",X"00",X"FF",X"22",X"69",X"62",X"22",X"12",X"22",X"10",X"00",X"FF",X"02",X"29",X"22",
		X"22",X"18",X"22",X"1E",X"00",X"FF",X"00",X"29",X"92",X"29",X"18",X"82",X"11",X"00",X"FF",X"00",
		X"29",X"99",X"29",X"11",X"11",X"11",X"00",X"FF",X"00",X"29",X"29",X"99",X"76",X"66",X"E1",X"10",
		X"FF",X"00",X"09",X"29",X"99",X"11",X"11",X"11",X"10",X"FF",X"00",X"09",X"99",X"99",X"12",X"22",
		X"11",X"10",X"FF",X"00",X"09",X"90",X"99",X"18",X"22",X"1E",X"10",X"FF",X"02",X"22",X"22",X"90",
		X"18",X"82",X"11",X"00",X"FF",X"22",X"22",X"22",X"20",X"11",X"11",X"11",X"00",X"FF",X"22",X"22",
		X"22",X"20",X"76",X"66",X"11",X"10",X"FF",X"22",X"22",X"22",X"22",X"06",X"66",X"61",X"10",X"FF",
		X"22",X"E1",X"E2",X"22",X"20",X"6D",X"6E",X"10",X"FF",X"02",X"22",X"22",X"22",X"20",X"6D",X"D8",
		X"10",X"FF",X"00",X"22",X"22",X"22",X"20",X"6D",X"D0",X"00",X"FF",X"00",X"22",X"22",X"22",X"20",
		X"6D",X"D0",X"00",X"FF",X"00",X"22",X"E1",X"E2",X"20",X"6D",X"D0",X"00",X"FF",X"00",X"02",X"22",
		X"22",X"00",X"6D",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"6D",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"08",X"88",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"77",X"A8",X"88",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"74",X"47",X"AA",X"88",X"80",X"FF",X"00",X"00",X"07",X"44",X"74",X"47",
		X"A8",X"88",X"81",X"FF",X"00",X"74",X"44",X"44",X"74",X"47",X"A8",X"88",X"88",X"FF",X"74",X"44",
		X"44",X"44",X"74",X"48",X"88",X"88",X"88",X"FF",X"77",X"44",X"44",X"47",X"74",X"88",X"88",X"88",
		X"88",X"FF",X"00",X"77",X"77",X"47",X"74",X"88",X"88",X"8A",X"88",X"FF",X"00",X"00",X"07",X"77",
		X"74",X"78",X"8A",X"A8",X"80",X"FF",X"00",X"00",X"00",X"00",X"74",X"78",X"88",X"A8",X"80",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"77",X"88",X"88",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"08",
		X"80",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"9C",X"CC",X"C0",X"00",X"00",X"00",X"FF",X"09",X"CC",
		X"CC",X"CC",X"00",X"00",X"00",X"FF",X"9C",X"CC",X"CE",X"44",X"9D",X"EE",X"00",X"FF",X"9C",X"CC",
		X"EB",X"B9",X"DE",X"CC",X"E0",X"FF",X"9C",X"CE",X"BB",X"99",X"DC",X"CC",X"C0",X"FF",X"9C",X"CE",
		X"BB",X"99",X"DC",X"CC",X"C0",X"FF",X"9C",X"CE",X"BB",X"99",X"DC",X"CC",X"C0",X"FF",X"9C",X"CE",
		X"47",X"99",X"DC",X"CC",X"C0",X"FF",X"9C",X"EB",X"B3",X"99",X"DC",X"CC",X"C0",X"FF",X"9C",X"BB",
		X"33",X"49",X"DE",X"CC",X"E0",X"FF",X"9C",X"BB",X"B4",X"B5",X"9D",X"EE",X"00",X"FF",X"09",X"EB",
		X"47",X"B3",X"00",X"00",X"00",X"FF",X"00",X"9E",X"74",X"B3",X"40",X"00",X"00",X"FF",X"00",X"07",
		X"74",X"4B",X"40",X"00",X"00",X"FF",X"00",X"44",X"00",X"77",X"00",X"00",X"00",X"FF",X"04",X"B0",
		X"00",X"44",X"00",X"00",X"00",X"FF",X"0B",X"B0",X"04",X"BB",X"00",X"00",X"00",X"FF",X"04",X"40",
		X"0B",X"B0",X"00",X"00",X"00",X"FF",X"00",X"40",X"0B",X"B0",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"04",X"BB",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"AA",
		X"11",X"00",X"00",X"00",X"00",X"FF",X"0A",X"A8",X"88",X"11",X"00",X"00",X"80",X"FF",X"AA",X"88",
		X"88",X"81",X"10",X"08",X"88",X"FF",X"AA",X"38",X"33",X"38",X"12",X"A8",X"8A",X"FF",X"AA",X"38",
		X"38",X"38",X"12",X"AA",X"A0",X"FF",X"A3",X"33",X"33",X"33",X"82",X"D8",X"88",X"FF",X"AA",X"38",
		X"38",X"38",X"82",X"28",X"80",X"FF",X"A3",X"33",X"33",X"33",X"82",X"00",X"00",X"FF",X"AA",X"38",
		X"38",X"38",X"80",X"20",X"00",X"FF",X"AA",X"33",X"38",X"38",X"20",X"02",X"00",X"FF",X"0A",X"AA",
		X"88",X"88",X"02",X"02",X"00",X"FF",X"00",X"AA",X"AA",X"00",X"20",X"20",X"00",X"FF",X"00",X"00",
		X"00",X"02",X"20",X"00",X"00",X"FF",X"00",X"00",X"22",X"22",X"00",X"00",X"00",X"FF",X"00",X"02",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"02",X"22",X"22",X"00",X"FF",X"00",X"22",X"21",X"11",X"20",X"FF",
		X"02",X"21",X"11",X"11",X"22",X"FF",X"02",X"21",X"22",X"22",X"22",X"FF",X"22",X"22",X"22",X"22",
		X"62",X"FF",X"22",X"22",X"22",X"26",X"62",X"FF",X"22",X"22",X"22",X"26",X"62",X"FF",X"22",X"22",
		X"21",X"22",X"62",X"FF",X"22",X"22",X"21",X"12",X"22",X"FF",X"02",X"22",X"21",X"11",X"12",X"FF",
		X"02",X"22",X"22",X"11",X"22",X"FF",X"00",X"22",X"11",X"12",X"20",X"FF",X"00",X"02",X"22",X"22",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"02",X"22",X"22",X"25",X"88",X"8D",X"00",X"00",X"00",X"FF",X"22",X"22",X"22",X"25",
		X"82",X"8D",X"DD",X"00",X"00",X"FF",X"22",X"21",X"22",X"55",X"8C",X"8D",X"DD",X"D0",X"00",X"FF",
		X"22",X"21",X"25",X"55",X"8C",X"8D",X"D2",X"DD",X"D0",X"FF",X"22",X"22",X"25",X"55",X"82",X"8D",
		X"D2",X"22",X"DD",X"FF",X"22",X"22",X"55",X"55",X"88",X"8D",X"D9",X"92",X"2D",X"FF",X"22",X"22",
		X"55",X"55",X"53",X"8D",X"D9",X"99",X"2D",X"FF",X"02",X"22",X"55",X"52",X"22",X"8D",X"D9",X"99",
		X"2D",X"FF",X"00",X"02",X"55",X"22",X"22",X"8D",X"DD",X"99",X"2D",X"FF",X"00",X"02",X"55",X"25",
		X"53",X"8D",X"DD",X"DD",X"2D",X"FF",X"00",X"02",X"55",X"55",X"88",X"8D",X"D2",X"DD",X"DD",X"FF",
		X"00",X"02",X"55",X"55",X"82",X"8D",X"D2",X"22",X"DD",X"FF",X"00",X"02",X"55",X"55",X"8C",X"8D",
		X"D9",X"92",X"2D",X"FF",X"00",X"02",X"55",X"55",X"8C",X"8D",X"D9",X"99",X"2D",X"FF",X"02",X"22",
		X"22",X"55",X"82",X"8D",X"D9",X"99",X"2D",X"FF",X"22",X"22",X"22",X"55",X"88",X"8D",X"DD",X"99",
		X"2D",X"FF",X"22",X"21",X"22",X"22",X"55",X"58",X"DD",X"DD",X"2D",X"FF",X"22",X"21",X"22",X"22",
		X"25",X"55",X"55",X"8D",X"DD",X"FF",X"22",X"22",X"22",X"22",X"22",X"55",X"55",X"55",X"8D",X"FF",
		X"22",X"22",X"22",X"22",X"25",X"55",X"55",X"55",X"58",X"FF",X"22",X"D1",X"1D",X"22",X"55",X"55",
		X"56",X"65",X"58",X"FF",X"02",X"22",X"22",X"22",X"22",X"22",X"56",X"55",X"80",X"FF",X"00",X"00",
		X"02",X"22",X"22",X"22",X"25",X"80",X"00",X"FF",X"00",X"00",X"02",X"2D",X"11",X"D2",X"58",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"22",X"22",X"22",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"88",
		X"EE",X"E8",X"00",X"00",X"00",X"00",X"FF",X"02",X"22",X"25",X"28",X"EE",X"EE",X"EE",X"80",X"00",
		X"00",X"FF",X"22",X"12",X"55",X"C8",X"EE",X"22",X"2E",X"EE",X"E0",X"00",X"FF",X"22",X"15",X"55",
		X"C8",X"EE",X"99",X"42",X"2E",X"DE",X"00",X"FF",X"22",X"25",X"55",X"28",X"EE",X"99",X"99",X"4E",
		X"DD",X"E0",X"FF",X"22",X"25",X"55",X"88",X"EE",X"99",X"99",X"4E",X"DD",X"E0",X"FF",X"22",X"25",
		X"55",X"38",X"EE",X"99",X"99",X"4E",X"DD",X"D0",X"FF",X"22",X"55",X"52",X"28",X"EE",X"EE",X"E9",
		X"4E",X"DD",X"D0",X"FF",X"02",X"55",X"22",X"28",X"EE",X"EE",X"EE",X"EE",X"DD",X"D0",X"FF",X"00",
		X"55",X"25",X"38",X"EE",X"22",X"2E",X"EE",X"DD",X"D0",X"FF",X"00",X"55",X"55",X"88",X"EE",X"99",
		X"42",X"2E",X"DD",X"D0",X"FF",X"00",X"55",X"55",X"28",X"EE",X"99",X"99",X"4E",X"DD",X"D0",X"FF",
		X"00",X"55",X"55",X"C8",X"EE",X"99",X"99",X"4E",X"DD",X"D0",X"FF",X"00",X"55",X"55",X"C8",X"EE",
		X"99",X"99",X"4E",X"DD",X"D0",X"FF",X"00",X"55",X"55",X"28",X"EE",X"EE",X"E9",X"4E",X"DD",X"D0",
		X"FF",X"02",X"25",X"55",X"88",X"8E",X"EE",X"EE",X"EE",X"DD",X"D0",X"FF",X"22",X"25",X"55",X"55",
		X"55",X"55",X"8E",X"EE",X"DD",X"D0",X"FF",X"22",X"12",X"22",X"22",X"55",X"55",X"55",X"55",X"ED",
		X"D0",X"FF",X"22",X"12",X"22",X"22",X"25",X"55",X"55",X"55",X"5E",X"D0",X"FF",X"22",X"22",X"22",
		X"22",X"22",X"55",X"55",X"66",X"55",X"E0",X"FF",X"22",X"22",X"22",X"22",X"25",X"55",X"55",X"56",
		X"55",X"80",X"FF",X"22",X"E1",X"1E",X"22",X"22",X"22",X"22",X"25",X"55",X"00",X"FF",X"02",X"22",
		X"22",X"20",X"22",X"22",X"22",X"22",X"50",X"00",X"FF",X"00",X"00",X"00",X"00",X"22",X"22",X"22",
		X"22",X"20",X"00",X"FF",X"00",X"00",X"00",X"00",X"02",X"2E",X"11",X"E2",X"20",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"22",X"22",X"22",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"02",X"22",X"22",X"20",X"05",X"88",X"80",
		X"00",X"00",X"FF",X"22",X"22",X"22",X"22",X"55",X"82",X"8D",X"00",X"00",X"FF",X"22",X"21",X"22",
		X"25",X"55",X"8C",X"81",X"00",X"00",X"FF",X"22",X"21",X"22",X"55",X"55",X"8C",X"81",X"D0",X"00",
		X"FF",X"22",X"22",X"22",X"55",X"55",X"82",X"81",X"10",X"00",X"FF",X"22",X"22",X"25",X"55",X"55",
		X"88",X"81",X"2D",X"00",X"FF",X"22",X"22",X"25",X"55",X"55",X"53",X"81",X"2D",X"00",X"FF",X"02",
		X"22",X"25",X"55",X"52",X"22",X"81",X"92",X"E0",X"FF",X"00",X"00",X"25",X"55",X"22",X"22",X"81",
		X"92",X"D0",X"FF",X"00",X"00",X"25",X"55",X"25",X"53",X"81",X"92",X"D0",X"FF",X"00",X"00",X"25",
		X"55",X"55",X"88",X"81",X"12",X"D0",X"FF",X"00",X"00",X"25",X"55",X"55",X"82",X"81",X"2D",X"D0",
		X"FF",X"00",X"00",X"25",X"55",X"55",X"8C",X"81",X"2D",X"D0",X"FF",X"00",X"00",X"25",X"55",X"55",
		X"8C",X"81",X"92",X"D0",X"FF",X"02",X"22",X"22",X"25",X"55",X"82",X"81",X"92",X"D0",X"FF",X"22",
		X"22",X"22",X"25",X"55",X"88",X"8D",X"92",X"D0",X"FF",X"22",X"21",X"22",X"22",X"55",X"55",X"58",
		X"12",X"D0",X"FF",X"22",X"21",X"22",X"22",X"25",X"55",X"55",X"D2",X"D0",X"FF",X"22",X"22",X"22",
		X"22",X"22",X"55",X"55",X"8D",X"D0",X"FF",X"22",X"22",X"22",X"22",X"22",X"55",X"55",X"5D",X"D0",
		X"FF",X"22",X"D1",X"1D",X"22",X"25",X"55",X"55",X"58",X"D0",X"FF",X"02",X"22",X"22",X"22",X"55",
		X"55",X"55",X"55",X"E0",X"FF",X"00",X"02",X"22",X"55",X"55",X"55",X"56",X"55",X"80",X"FF",X"00",
		X"02",X"22",X"22",X"55",X"55",X"66",X"55",X"00",X"FF",X"00",X"02",X"22",X"22",X"22",X"55",X"55",
		X"50",X"00",X"FF",X"00",X"02",X"22",X"22",X"22",X"25",X"50",X"00",X"00",X"FF",X"00",X"02",X"2E",
		X"11",X"E2",X"25",X"00",X"00",X"00",X"FF",X"00",X"00",X"22",X"22",X"22",X"50",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"09",X"44",X"00",X"00",X"00",X"00",X"FF",X"00",X"94",X"5B",X"50",X"00",
		X"00",X"00",X"FF",X"00",X"94",X"B8",X"B0",X"00",X"00",X"00",X"FF",X"00",X"94",X"B8",X"B0",X"00",
		X"00",X"00",X"FF",X"00",X"94",X"5B",X"50",X"00",X"00",X"00",X"FF",X"00",X"09",X"44",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"0D",X"D0",X"00",X"00",X"00",X"FF",X"09",X"44",X"00",X"D0",X"00",
		X"00",X"00",X"FF",X"94",X"5B",X"50",X"DD",X"00",X"00",X"00",X"FF",X"94",X"B8",X"B0",X"0D",X"DD",
		X"00",X"00",X"FF",X"94",X"B8",X"B0",X"00",X"0D",X"DD",X"D0",X"FF",X"94",X"5B",X"5D",X"00",X"DD",
		X"DD",X"D0",X"FF",X"09",X"44",X"0D",X"DD",X"D0",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"0C",
		X"E0",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"CC",X"E0",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"CE",X"EE",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"CE",X"8E",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"15",X"EE",X"8E",X"00",X"00",X"00",X"00",X"00",X"FF",X"05",X"EE",X"EE",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"01",X"EE",X"EE",X"00",X"07",X"00",X"00",X"00",X"FF",X"05",X"EB",X"EC",
		X"00",X"07",X"70",X"00",X"00",X"FF",X"05",X"EB",X"CC",X"11",X"16",X"22",X"16",X"00",X"FF",X"15",
		X"EB",X"B1",X"11",X"16",X"11",X"16",X"60",X"FF",X"05",X"EE",X"C1",X"B1",X"66",X"66",X"66",X"60",
		X"FF",X"15",X"EE",X"C1",X"BB",X"B6",X"66",X"66",X"60",X"FF",X"01",X"EB",X"C6",X"6B",X"B6",X"66",
		X"66",X"60",X"FF",X"15",X"EB",X"B6",X"66",X"66",X"66",X"66",X"00",X"FF",X"15",X"EB",X"EE",X"66",
		X"66",X"66",X"60",X"00",X"FF",X"01",X"EE",X"EE",X"00",X"77",X"00",X"00",X"00",X"FF",X"05",X"CE",
		X"EE",X"00",X"07",X"00",X"00",X"00",X"FF",X"01",X"5E",X"E0",X"00",X"07",X"00",X"00",X"00",X"FF",
		X"01",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"01",X"01",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"10",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"0C",X"E0",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"CC",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"CE",X"EE",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"CE",
		X"8E",X"00",X"00",X"00",X"00",X"00",X"FF",X"05",X"EE",X"8E",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"15",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"FF",X"05",X"EE",X"EE",X"00",X"07",X"00",X"00",
		X"00",X"FF",X"05",X"EB",X"EC",X"00",X"07",X"70",X"00",X"00",X"FF",X"11",X"EB",X"CC",X"11",X"16",
		X"22",X"16",X"00",X"FF",X"05",X"EB",X"B1",X"11",X"16",X"11",X"16",X"60",X"FF",X"05",X"EE",X"C1",
		X"B1",X"66",X"66",X"66",X"60",X"FF",X"15",X"EE",X"C1",X"BB",X"B6",X"66",X"66",X"60",X"FF",X"05",
		X"EB",X"C6",X"6B",X"B6",X"66",X"66",X"60",X"FF",X"15",X"EB",X"B6",X"66",X"66",X"66",X"66",X"00",
		X"FF",X"15",X"EB",X"EE",X"66",X"66",X"66",X"60",X"00",X"FF",X"01",X"EE",X"EE",X"07",X"70",X"00",
		X"00",X"00",X"FF",X"05",X"CE",X"EE",X"07",X"00",X"00",X"00",X"00",X"FF",X"01",X"5E",X"E0",X"07",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"FF",X"01",X"01",
		X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"01",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"10",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"DD",X"DD",X"FF",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"FF",X"DD",X"5D",X"DD",X"CD",
		X"DD",X"DD",X"DD",X"DD",X"FF",X"DD",X"55",X"DC",X"ED",X"DD",X"DD",X"DD",X"DD",X"FF",X"DD",X"55",
		X"DE",X"ED",X"DD",X"DD",X"DD",X"DD",X"FF",X"DD",X"55",X"CE",X"EC",X"DD",X"DD",X"DD",X"DD",X"FF",
		X"D5",X"55",X"EE",X"EE",X"DD",X"DD",X"DD",X"DD",X"FF",X"D5",X"5C",X"EE",X"EE",X"DD",X"DD",X"DD",
		X"DD",X"FF",X"D5",X"5E",X"EE",X"EE",X"DD",X"DD",X"DD",X"DD",X"FF",X"D5",X"5E",X"EE",X"EE",X"DD",
		X"7D",X"DD",X"DD",X"FF",X"D5",X"CE",X"BE",X"EE",X"DD",X"77",X"DD",X"DD",X"FF",X"D5",X"EE",X"BC",
		X"C1",X"11",X"62",X"21",X"6D",X"FF",X"DD",X"EE",X"BB",X"11",X"11",X"61",X"11",X"66",X"FF",X"D1",
		X"EE",X"CC",X"11",X"16",X"66",X"66",X"66",X"FF",X"DD",X"EE",X"BC",X"11",X"B7",X"66",X"66",X"66",
		X"FF",X"1D",X"EE",X"BB",X"66",X"77",X"66",X"66",X"66",X"FF",X"1D",X"EE",X"BE",X"66",X"67",X"77",
		X"66",X"6D",X"FF",X"DD",X"EE",X"EE",X"D6",X"66",X"66",X"66",X"DD",X"FF",X"11",X"CE",X"ED",X"DD",
		X"DD",X"77",X"DD",X"DD",X"FF",X"D1",X"CC",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"FF",X"DD",X"DD",
		X"1D",X"DD",X"DD",X"DD",X"DD",X"DD",X"FF",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"FF",
		X"D1",X"DD",X"D1",X"DD",X"DD",X"DD",X"DD",X"DD",X"FF",X"DD",X"1D",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"DD",X"FF",X"DD",X"D1",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"FF",X"D1",X"DD",X"DD",X"DD",X"DD",
		X"DD",X"DD",X"DD",X"FF",X"DD",X"1D",X"1D",X"DD",X"DD",X"DD",X"DD",X"DD",X"FF",X"1D",X"1D",X"DD",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"FF",X"DD",X"D1",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"FF",X"DD",
		X"1D",X"D1",X"DD",X"DD",X"DD",X"DD",X"DD",X"FF",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"FF",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"FF",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"DD",X"DD",X"FF",X"DD",X"D1",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"FF",X"DD",X"DD",X"DD",X"DD",
		X"DD",X"DD",X"DD",X"DD",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"BB",X"CC",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"0C",X"BB",X"CC",X"BB",X"C0",X"00",X"00",
		X"FF",X"00",X"00",X"0B",X"CC",X"BB",X"CC",X"BB",X"C0",X"00",X"00",X"FF",X"00",X"00",X"00",X"BB",
		X"CC",X"BB",X"CC",X"BB",X"00",X"00",X"FF",X"0E",X"EE",X"EE",X"EB",X"CC",X"BB",X"CC",X"BB",X"00",
		X"00",X"FF",X"EE",X"EE",X"EE",X"EC",X"BB",X"CC",X"BB",X"CC",X"B0",X"00",X"FF",X"EE",X"EE",X"ED",
		X"EE",X"BB",X"CC",X"BB",X"CC",X"B0",X"00",X"FF",X"EE",X"EE",X"EE",X"EE",X"CC",X"BB",X"CC",X"BB",
		X"CC",X"00",X"FF",X"EE",X"EE",X"EE",X"EE",X"EC",X"BB",X"CC",X"BB",X"CC",X"00",X"FF",X"EE",X"55",
		X"55",X"EE",X"EB",X"CC",X"BB",X"CC",X"BB",X"C0",X"FF",X"0E",X"57",X"75",X"EE",X"EE",X"CC",X"BB",
		X"CC",X"BB",X"C0",X"FF",X"00",X"07",X"0E",X"EE",X"EE",X"BB",X"CC",X"BB",X"CC",X"77",X"FF",X"00",
		X"07",X"0E",X"E5",X"55",X"5B",X"CC",X"B7",X"77",X"70",X"FF",X"00",X"07",X"70",X"E5",X"44",X"5C",
		X"77",X"77",X"00",X"00",X"FF",X"00",X"07",X"77",X"00",X"47",X"77",X"70",X"00",X"00",X"00",X"FF",
		X"00",X"07",X"07",X"47",X"77",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"07",X"00",X"47",X"40",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"0E",X"EE",X"EE",X"E4",X"40",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"EE",X"EE",X"EE",X"EE",X"40",X"00",X"00",X"00",X"00",X"00",X"FF",X"EE",X"EE",X"ED",X"EE",
		X"40",X"00",X"00",X"00",X"00",X"00",X"FF",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"00",X"00",X"00",
		X"00",X"FF",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"E0",X"00",X"00",X"00",X"FF",X"EE",X"9D",X"D9",
		X"EE",X"EE",X"DE",X"E0",X"00",X"00",X"00",X"FF",X"0E",X"EE",X"EE",X"EE",X"EE",X"EE",X"E0",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"0E",X"EE",X"EE",X"EE",X"E0",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"0E",X"E9",X"DD",X"9E",X"E0",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"EE",X"EE",X"EE",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"0B",X"BC",X"C0",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"CB",
		X"BC",X"CB",X"B0",X"00",X"00",X"00",X"FF",X"00",X"0B",X"BC",X"CB",X"BC",X"CB",X"B0",X"00",X"00",
		X"FF",X"00",X"CB",X"BC",X"CB",X"BC",X"CB",X"BC",X"C0",X"00",X"FF",X"0B",X"BC",X"CB",X"BC",X"CB",
		X"BC",X"CB",X"BC",X"C7",X"FF",X"0B",X"BC",X"CB",X"BC",X"CB",X"BC",X"CB",X"BC",X"77",X"FF",X"EE",
		X"EB",X"BC",X"CB",X"BC",X"CB",X"BC",X"C7",X"70",X"FF",X"EE",X"EE",X"EC",X"CB",X"BC",X"CB",X"BC",
		X"77",X"00",X"FF",X"EE",X"55",X"5E",X"EC",X"CB",X"BC",X"C7",X"7E",X"00",X"FF",X"0E",X"57",X"7E",
		X"00",X"0B",X"BC",X"77",X"EE",X"00",X"FF",X"00",X"07",X"00",X"00",X"0E",X"E7",X"75",X"EE",X"00",
		X"FF",X"00",X"07",X"00",X"00",X"00",X"77",X"45",X"E0",X"00",X"FF",X"00",X"07",X"77",X"00",X"07",
		X"77",X"00",X"00",X"00",X"FF",X"00",X"07",X"77",X"77",X"77",X"07",X"00",X"00",X"00",X"FF",X"00",
		X"07",X"00",X"77",X"77",X"77",X"00",X"00",X"00",X"FF",X"00",X"07",X"00",X"00",X"07",X"77",X"00",
		X"00",X"00",X"FF",X"0E",X"EE",X"EE",X"E0",X"00",X"07",X"00",X"00",X"00",X"FF",X"EE",X"EE",X"EE",
		X"EE",X"00",X"07",X"00",X"00",X"00",X"FF",X"EE",X"EE",X"DE",X"EE",X"0E",X"EE",X"EE",X"E0",X"00",
		X"FF",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"00",X"FF",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"EE",X"DE",X"EE",X"00",X"FF",X"EE",X"9D",X"D9",X"EE",X"EE",X"EE",X"EE",X"EE",X"00",X"FF",X"0E",
		X"EE",X"EE",X"E0",X"EE",X"EE",X"EE",X"EE",X"00",X"FF",X"00",X"00",X"00",X"00",X"EE",X"9D",X"D9",
		X"EE",X"00",X"FF",X"00",X"00",X"00",X"00",X"0E",X"EE",X"EE",X"E0",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"0B",X"BC",X"CB",X"BC",X"C0",X"FF",X"00",X"00",X"00",X"00",X"00",X"0B",X"BC",X"CB",
		X"BC",X"C0",X"FF",X"00",X"00",X"00",X"00",X"00",X"0C",X"CB",X"BC",X"CB",X"B0",X"FF",X"0E",X"EE",
		X"EE",X"E0",X"00",X"0C",X"CB",X"BC",X"CB",X"B0",X"FF",X"EE",X"EE",X"EE",X"EE",X"00",X"0B",X"BC",
		X"CB",X"BC",X"C0",X"FF",X"EE",X"EE",X"ED",X"EE",X"00",X"0B",X"BC",X"CB",X"BC",X"C0",X"FF",X"EE",
		X"EE",X"EE",X"EE",X"00",X"0C",X"CB",X"BC",X"CB",X"B0",X"FF",X"EE",X"EE",X"EE",X"EE",X"E0",X"0C",
		X"CB",X"BC",X"CB",X"B0",X"FF",X"EE",X"55",X"55",X"EE",X"EE",X"0B",X"BC",X"CB",X"BC",X"C0",X"FF",
		X"0E",X"57",X"75",X"ED",X"EE",X"0B",X"BC",X"CB",X"BC",X"C0",X"FF",X"00",X"E7",X"EE",X"EE",X"EE",
		X"0C",X"CB",X"BC",X"CB",X"B0",X"FF",X"00",X"E7",X"EE",X"EE",X"EE",X"0C",X"CB",X"BC",X"CB",X"B0",
		X"FF",X"00",X"E7",X"55",X"55",X"EE",X"0B",X"BC",X"CB",X"BC",X"C0",X"FF",X"00",X"07",X"54",X"45",
		X"EE",X"0B",X"BC",X"CB",X"BC",X"C0",X"FF",X"00",X"07",X"77",X"77",X"77",X"77",X"77",X"77",X"77",
		X"70",X"FF",X"00",X"07",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"0E",X"EE",X"EE",
		X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"EE",X"EE",X"EE",X"EE",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"EE",X"EE",X"ED",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"EE",X"EE",
		X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"EE",X"EE",X"EE",X"EE",X"E0",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"EE",X"9D",X"D9",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"FF",X"0E",
		X"EE",X"EE",X"ED",X"EE",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"EE",X"EE",X"EE",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"EE",X"EE",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"EE",X"9D",X"D9",X"EE",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"0E",X"EE",X"EE",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"08",X"76",X"60",X"00",X"FF",X"00",X"87",X"66",
		X"66",X"00",X"FF",X"00",X"87",X"68",X"86",X"00",X"FF",X"08",X"76",X"99",X"88",X"60",X"FF",X"08",
		X"76",X"E9",X"98",X"60",X"FF",X"08",X"76",X"EE",X"98",X"60",X"FF",X"87",X"6E",X"EE",X"98",X"86",
		X"FF",X"87",X"6E",X"EE",X"99",X"86",X"FF",X"87",X"6E",X"EE",X"E9",X"86",X"FF",X"87",X"6E",X"EE",
		X"E9",X"86",X"FF",X"87",X"6E",X"EE",X"E9",X"86",X"FF",X"87",X"6E",X"EE",X"E9",X"86",X"FF",X"87",
		X"6E",X"EE",X"E9",X"86",X"FF",X"87",X"6E",X"EE",X"E9",X"86",X"FF",X"87",X"6E",X"EE",X"99",X"86",
		X"FF",X"87",X"6E",X"EE",X"98",X"86",X"FF",X"08",X"76",X"EE",X"98",X"60",X"FF",X"08",X"76",X"E9",
		X"98",X"60",X"FF",X"08",X"76",X"99",X"88",X"60",X"FF",X"00",X"87",X"68",X"86",X"00",X"FF",X"00",
		X"87",X"66",X"66",X"00",X"FF",X"00",X"08",X"76",X"60",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"08",X"76",X"60",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"87",X"66",X"66",X"00",X"00",X"00",X"00",X"FF",X"00",X"87",X"68",X"86",
		X"00",X"00",X"00",X"00",X"FF",X"08",X"76",X"99",X"88",X"60",X"00",X"00",X"00",X"FF",X"08",X"76",
		X"E9",X"98",X"60",X"00",X"00",X"00",X"FF",X"08",X"76",X"EE",X"98",X"60",X"00",X"00",X"00",X"FF",
		X"87",X"6E",X"54",X"32",X"86",X"00",X"00",X"00",X"FF",X"87",X"65",X"43",X"21",X"16",X"00",X"00",
		X"00",X"FF",X"87",X"65",X"42",X"23",X"31",X"DC",X"BB",X"A0",X"FF",X"87",X"65",X"3E",X"1E",X"31",
		X"00",X"00",X"00",X"FF",X"87",X"65",X"42",X"22",X"22",X"00",X"00",X"00",X"FF",X"87",X"65",X"42",
		X"22",X"22",X"00",X"00",X"00",X"FF",X"87",X"65",X"4E",X"2E",X"32",X"00",X"00",X"00",X"FF",X"87",
		X"65",X"44",X"33",X"32",X"DC",X"BB",X"A0",X"FF",X"87",X"65",X"54",X"43",X"26",X"00",X"00",X"00",
		X"FF",X"87",X"6E",X"55",X"44",X"86",X"00",X"00",X"00",X"FF",X"08",X"76",X"EE",X"98",X"60",X"00",
		X"00",X"00",X"FF",X"08",X"76",X"E9",X"98",X"60",X"00",X"00",X"00",X"FF",X"08",X"76",X"99",X"88",
		X"60",X"00",X"00",X"00",X"FF",X"00",X"87",X"68",X"86",X"00",X"00",X"00",X"00",X"FF",X"00",X"87",
		X"66",X"66",X"00",X"00",X"00",X"00",X"FF",X"00",X"08",X"76",X"60",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"08",X"76",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"87",X"66",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"87",X"68",
		X"86",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"08",X"76",X"99",X"88",X"60",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"08",X"76",X"E9",X"98",X"60",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"08",X"76",X"EE",X"98",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"87",X"6E",X"EE",
		X"98",X"86",X"05",X"43",X"20",X"00",X"00",X"00",X"FF",X"87",X"6E",X"EE",X"99",X"86",X"54",X"32",
		X"11",X"00",X"00",X"00",X"FF",X"87",X"64",X"23",X"23",X"2E",X"54",X"22",X"22",X"1D",X"CB",X"BA",
		X"FF",X"87",X"65",X"34",X"34",X"3E",X"53",X"E1",X"2E",X"10",X"00",X"00",X"FF",X"87",X"65",X"35",
		X"34",X"3E",X"54",X"22",X"22",X"20",X"00",X"00",X"FF",X"87",X"65",X"35",X"35",X"3E",X"54",X"22",
		X"22",X"20",X"00",X"00",X"FF",X"87",X"65",X"35",X"35",X"3E",X"54",X"E2",X"3E",X"20",X"00",X"00",
		X"FF",X"87",X"6E",X"4E",X"4E",X"4E",X"54",X"43",X"33",X"2D",X"CB",X"BA",X"FF",X"87",X"6E",X"EE",
		X"99",X"86",X"55",X"44",X"32",X"00",X"00",X"00",X"FF",X"87",X"6E",X"EE",X"98",X"86",X"05",X"54",
		X"40",X"00",X"00",X"00",X"FF",X"08",X"76",X"EE",X"98",X"60",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"08",X"76",X"E9",X"98",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"08",X"76",X"99",
		X"88",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"87",X"68",X"86",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"87",X"66",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"08",X"76",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"05",X"55",X"50",X"00",X"02",X"30",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"35",X"50",X"00",X"00",X"03",X"55",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"33",X"55",X"00",X"00",X"00",X"55",X"D0",X"0D",X"00",X"00",X"00",X"FF",X"00",X"00",X"05",
		X"0E",X"DD",X"E5",X"5D",X"DD",X"00",X"D0",X"00",X"00",X"FF",X"00",X"00",X"05",X"DD",X"DC",X"DD",
		X"DB",X"BC",X"CD",X"D0",X"00",X"00",X"FF",X"00",X"00",X"5D",X"DC",X"CC",X"BB",X"BC",X"CD",X"BB",
		X"CD",X"0D",X"00",X"FF",X"00",X"0E",X"ED",X"CC",X"BC",X"CB",X"CC",X"65",X"BC",X"CD",X"CD",X"00",
		X"FF",X"00",X"0E",X"DD",X"CB",X"AB",X"CC",X"CD",X"E5",X"DB",X"CC",X"D0",X"00",X"FF",X"00",X"ED",
		X"DC",X"BA",X"AA",X"BC",X"CD",X"EA",X"BB",X"BD",X"DD",X"00",X"FF",X"00",X"ED",X"CB",X"AA",X"BB",
		X"CC",X"3C",X"DD",X"BB",X"CC",X"CD",X"D0",X"FF",X"00",X"DC",X"CB",X"AB",X"BC",X"CC",X"3C",X"DB",
		X"BB",X"CC",X"CD",X"00",X"FF",X"00",X"ED",X"CD",X"BC",X"CC",X"CC",X"CD",X"EA",X"DB",X"BC",X"CC",
		X"D0",X"FF",X"03",X"EE",X"DD",X"DB",X"CC",X"CC",X"CD",X"E5",X"ED",X"CC",X"DD",X"0D",X"FF",X"35",
		X"53",X"33",X"DB",X"CC",X"BC",X"CC",X"65",X"EE",X"DC",X"D0",X"00",X"FF",X"55",X"ED",X"DB",X"BC",
		X"CC",X"CB",X"CC",X"CD",X"C4",X"2D",X"0D",X"00",X"FF",X"55",X"0E",X"DB",X"CD",X"DD",X"DD",X"BB",
		X"DE",X"41",X"4E",X"00",X"00",X"FF",X"55",X"0D",X"DC",X"DD",X"00",X"E5",X"5D",X"EE",X"24",X"20",
		X"00",X"00",X"FF",X"05",X"00",X"DC",X"D0",X"00",X"00",X"55",X"0E",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"ED",X"00",X"00",X"03",X"55",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"0E",
		X"D0",X"00",X"02",X"30",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"23",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"05",X"00",
		X"00",X"00",X"35",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"55",X"00",X"00",X"00",X"00",
		X"55",X"00",X"D0",X"0D",X"00",X"00",X"00",X"FF",X"55",X"00",X"00",X"0E",X"DD",X"E5",X"DD",X"DD",
		X"00",X"D0",X"00",X"00",X"FF",X"35",X"50",X"0E",X"DD",X"DC",X"DD",X"DB",X"BC",X"CD",X"D0",X"00",
		X"00",X"FF",X"35",X"33",X"33",X"DC",X"CC",X"BB",X"BC",X"CD",X"BB",X"CD",X"0D",X"00",X"FF",X"03",
		X"0E",X"ED",X"CC",X"BC",X"CB",X"CC",X"65",X"BC",X"CD",X"CD",X"00",X"FF",X"00",X"0E",X"DD",X"CB",
		X"AB",X"CC",X"CD",X"E5",X"DB",X"CC",X"D0",X"00",X"FF",X"00",X"ED",X"DC",X"BA",X"AA",X"BC",X"3D",
		X"EA",X"BB",X"BD",X"DD",X"00",X"FF",X"00",X"ED",X"CB",X"AA",X"BB",X"CC",X"3C",X"DD",X"BB",X"CC",
		X"CD",X"D0",X"FF",X"00",X"DC",X"CB",X"AB",X"BC",X"CC",X"3C",X"DB",X"BB",X"CC",X"CD",X"00",X"FF",
		X"00",X"ED",X"CD",X"BC",X"CC",X"CC",X"3D",X"EA",X"DB",X"BC",X"CC",X"D0",X"FF",X"03",X"EE",X"DD",
		X"DB",X"CC",X"CC",X"CD",X"E5",X"ED",X"CC",X"DD",X"0D",X"FF",X"35",X"33",X"33",X"DB",X"CC",X"BC",
		X"CC",X"65",X"EE",X"DC",X"D0",X"00",X"FF",X"35",X"5D",X"DB",X"BC",X"CC",X"CB",X"CC",X"CD",X"C4",
		X"2D",X"0D",X"00",X"FF",X"55",X"0E",X"DB",X"CD",X"DD",X"DD",X"BB",X"DE",X"41",X"4E",X"00",X"00",
		X"FF",X"55",X"0D",X"DC",X"DD",X"00",X"E5",X"ED",X"EE",X"24",X"20",X"00",X"00",X"FF",X"05",X"00",
		X"DC",X"D0",X"00",X"55",X"00",X"0E",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"ED",X"00",X"35",
		X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"0E",X"D0",X"23",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"05",X"00",X"00",X"00",X"35",X"50",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"55",X"00",X"00",X"00",X"00",X"33",X"00",X"D0",X"00",X"00",
		X"00",X"00",X"FF",X"55",X"00",X"00",X"0E",X"DD",X"E3",X"CD",X"DC",X"00",X"D0",X"00",X"00",X"FF",
		X"35",X"50",X"0E",X"DD",X"DD",X"DD",X"AA",X"AA",X"CD",X"D0",X"00",X"00",X"FF",X"35",X"33",X"33",
		X"DC",X"DD",X"BA",X"69",X"6A",X"1B",X"DD",X"0D",X"00",X"FF",X"03",X"0E",X"ED",X"CC",X"DB",X"AA",
		X"99",X"99",X"11",X"BD",X"CD",X"00",X"FF",X"00",X"0E",X"DD",X"CC",X"DB",X"A6",X"69",X"66",X"A1",
		X"BC",X"D0",X"00",X"FF",X"00",X"ED",X"DB",X"BB",X"DB",X"A9",X"99",X"99",X"A1",X"BC",X"DD",X"00",
		X"FF",X"00",X"ED",X"BB",X"BC",X"DB",X"A6",X"69",X"66",X"A1",X"BC",X"CD",X"D0",X"FF",X"00",X"DC",
		X"BB",X"CB",X"CB",X"A9",X"99",X"99",X"A1",X"BC",X"DD",X"00",X"FF",X"00",X"ED",X"CD",X"BC",X"CB",
		X"A6",X"69",X"66",X"A1",X"BC",X"CC",X"D0",X"FF",X"03",X"EE",X"DD",X"DB",X"DB",X"A9",X"99",X"99",
		X"A1",X"BD",X"DD",X"0D",X"FF",X"35",X"33",X"33",X"DB",X"DB",X"AA",X"69",X"66",X"11",X"BD",X"D0",
		X"00",X"FF",X"35",X"5D",X"CB",X"BC",X"CD",X"BA",X"A9",X"9A",X"1C",X"22",X"0D",X"00",X"FF",X"55",
		X"0E",X"DB",X"CD",X"DD",X"DD",X"AA",X"AA",X"D2",X"12",X"00",X"00",X"FF",X"55",X"0D",X"DC",X"DD",
		X"00",X"E3",X"ED",X"EE",X"02",X"20",X"00",X"00",X"FF",X"05",X"00",X"DC",X"D0",X"00",X"33",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"ED",X"00",X"55",X"50",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"0E",X"D0",X"25",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"05",X"00",X"00",X"00",X"35",X"50",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"55",X"00",X"00",X"00",X"00",X"33",X"00",X"D0",X"00",X"00",X"00",X"00",X"FF",X"55",X"00",
		X"00",X"0E",X"DD",X"E3",X"CD",X"DC",X"00",X"D0",X"00",X"00",X"FF",X"35",X"50",X"0E",X"DD",X"DD",
		X"DD",X"AA",X"AA",X"CD",X"D0",X"00",X"00",X"FF",X"35",X"33",X"33",X"DC",X"DD",X"BA",X"69",X"6A",
		X"1B",X"DD",X"0D",X"00",X"FF",X"03",X"0E",X"ED",X"CC",X"DB",X"AA",X"99",X"99",X"11",X"BD",X"CD",
		X"00",X"FF",X"00",X"0E",X"DD",X"CC",X"DB",X"A6",X"99",X"96",X"A1",X"BC",X"D0",X"00",X"FF",X"00",
		X"ED",X"DB",X"BB",X"DB",X"A9",X"99",X"99",X"A1",X"BC",X"DD",X"00",X"FF",X"00",X"ED",X"BB",X"BC",
		X"DB",X"A6",X"99",X"96",X"A1",X"BC",X"CD",X"D0",X"FF",X"00",X"DC",X"BB",X"CB",X"CB",X"A9",X"99",
		X"99",X"A1",X"BC",X"DD",X"00",X"FF",X"00",X"ED",X"CD",X"BC",X"CB",X"A6",X"99",X"96",X"A1",X"BC",
		X"CC",X"D0",X"FF",X"03",X"EE",X"DD",X"DB",X"DB",X"A9",X"99",X"99",X"A1",X"BD",X"DD",X"0D",X"FF",
		X"35",X"33",X"33",X"DB",X"DB",X"AA",X"69",X"96",X"11",X"BD",X"D0",X"00",X"FF",X"35",X"5D",X"CB",
		X"BC",X"CD",X"BA",X"A9",X"9A",X"1C",X"22",X"0D",X"00",X"FF",X"55",X"0E",X"DB",X"CD",X"DD",X"DD",
		X"AA",X"AA",X"D2",X"12",X"00",X"00",X"FF",X"55",X"0D",X"DC",X"DD",X"00",X"E3",X"ED",X"EE",X"02",
		X"20",X"00",X"00",X"FF",X"05",X"00",X"DC",X"D0",X"00",X"33",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"ED",X"00",X"55",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"0E",X"D0",X"25",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"0E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"10",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"20",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"30",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"40",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"50",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"60",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"70",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"80",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"90",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
