library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

-- bass.wav    e:RIFF n:1 sr:11025 br:11025 al:1 bps:8 lg:  2005 start:    44(x   2C) stop:  2050(x  802)
-- congal.wav  e:RIFF n:1 sr:11025 br:11025 al:1 bps:8 lg:  2003 start:  2094(x  82E) stop:  4098(x 1002)
-- congah.wav  e:RIFF n:1 sr:11025 br:11025 al:1 bps:8 lg:  1970 start:  4142(x 102E) stop:  6112(x 17E0)
-- rim.wav     e:RIFF n:1 sr:11025 br:11025 al:1 bps:8 lg:   373 start:  6156(x 180C) stop:  6530(x 1982)
-- gorilla.wav e:RIFF n:1 sr:11025 br:11025 al:1 bps:8 lg:  4991 start:  6574(x 19AE) stop: 11566(x 2D2E)

entity congo_samples is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of congo_samples is
	type rom is array(0 to  11565) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"52",X"49",X"46",X"46",X"FA",X"07",X"00",X"00",X"57",X"41",X"56",X"45",X"66",X"6D",X"74",X"20",
		X"10",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"11",X"2B",X"00",X"00",X"11",X"2B",X"00",X"00",
		X"01",X"00",X"08",X"00",X"64",X"61",X"74",X"61",X"D5",X"07",X"00",X"00",X"80",X"7E",X"80",X"7F",
		X"81",X"7F",X"7F",X"80",X"81",X"7E",X"81",X"7F",X"7E",X"7F",X"81",X"80",X"7D",X"7F",X"7D",X"80",
		X"79",X"85",X"36",X"00",X"10",X"0A",X"10",X"0E",X"15",X"12",X"15",X"19",X"1D",X"20",X"1F",X"22",
		X"23",X"25",X"28",X"27",X"2C",X"2D",X"30",X"31",X"32",X"36",X"37",X"3A",X"3B",X"43",X"4B",X"50",
		X"56",X"5C",X"64",X"6C",X"73",X"7B",X"82",X"8B",X"92",X"9A",X"A3",X"AA",X"B2",X"B9",X"C0",X"C7",
		X"CE",X"D5",X"DB",X"E1",X"E7",X"EB",X"F1",X"F0",X"ED",X"EC",X"E9",X"E7",X"E5",X"E3",X"E1",X"DF",
		X"DC",X"DA",X"D9",X"D6",X"D4",X"D3",X"D1",X"CF",X"CE",X"CC",X"CB",X"C9",X"C7",X"C6",X"C4",X"C3",
		X"C1",X"C0",X"BE",X"BD",X"BB",X"BA",X"B8",X"B8",X"B6",X"B5",X"B4",X"B3",X"B2",X"B0",X"B0",X"AE",
		X"AD",X"AC",X"AB",X"AA",X"A9",X"A8",X"A7",X"A6",X"A5",X"A4",X"A4",X"A3",X"A2",X"A1",X"A0",X"9F",
		X"9F",X"9E",X"9D",X"9C",X"9B",X"9A",X"98",X"97",X"95",X"94",X"92",X"90",X"8F",X"8D",X"8B",X"89",
		X"87",X"85",X"83",X"80",X"7E",X"7C",X"7A",X"77",X"75",X"73",X"70",X"6E",X"6C",X"69",X"67",X"65",
		X"62",X"60",X"5E",X"5C",X"59",X"57",X"55",X"53",X"51",X"50",X"4E",X"4C",X"4A",X"49",X"47",X"46",
		X"44",X"43",X"42",X"41",X"40",X"3F",X"3E",X"3E",X"3D",X"3C",X"3C",X"3B",X"3B",X"3B",X"3B",X"3B",
		X"3B",X"3C",X"3C",X"3D",X"3D",X"3E",X"3F",X"40",X"41",X"42",X"43",X"44",X"45",X"47",X"49",X"4A",
		X"4C",X"4E",X"4F",X"51",X"53",X"55",X"57",X"59",X"5B",X"5E",X"60",X"62",X"64",X"67",X"69",X"6C",
		X"6E",X"70",X"73",X"75",X"78",X"7A",X"7C",X"7F",X"81",X"83",X"85",X"88",X"8A",X"8C",X"8E",X"90",
		X"92",X"94",X"96",X"98",X"9A",X"9C",X"9E",X"9F",X"A1",X"A2",X"A3",X"A5",X"A6",X"A7",X"A8",X"A9",
		X"AA",X"AB",X"AC",X"AC",X"AD",X"AD",X"AE",X"AE",X"AE",X"AE",X"AE",X"AE",X"AE",X"AE",X"AD",X"AD",
		X"AC",X"AC",X"AB",X"AB",X"AA",X"A9",X"A8",X"A7",X"A6",X"A4",X"A3",X"A2",X"A1",X"9F",X"9E",X"9C",
		X"9B",X"99",X"98",X"96",X"94",X"92",X"90",X"8F",X"8D",X"8B",X"89",X"87",X"85",X"83",X"81",X"7F",
		X"7D",X"7B",X"7A",X"78",X"76",X"74",X"72",X"70",X"6F",X"6D",X"6B",X"6A",X"68",X"66",X"65",X"63",
		X"62",X"61",X"5F",X"5E",X"5D",X"5C",X"5B",X"5A",X"59",X"58",X"57",X"57",X"56",X"55",X"55",X"55",
		X"54",X"54",X"54",X"54",X"54",X"54",X"54",X"54",X"54",X"55",X"55",X"56",X"56",X"57",X"57",X"58",
		X"59",X"5A",X"5B",X"5C",X"5D",X"5E",X"5F",X"61",X"62",X"63",X"65",X"66",X"67",X"69",X"6B",X"6C",
		X"6E",X"6F",X"71",X"72",X"74",X"76",X"77",X"79",X"7B",X"7D",X"7E",X"80",X"82",X"83",X"85",X"87",
		X"88",X"8A",X"8B",X"8D",X"8E",X"90",X"91",X"93",X"94",X"95",X"97",X"98",X"99",X"9A",X"9B",X"9C",
		X"9D",X"9E",X"9F",X"A0",X"A1",X"A1",X"A2",X"A2",X"A3",X"A3",X"A4",X"A4",X"A4",X"A4",X"A4",X"A4",
		X"A4",X"A4",X"A4",X"A3",X"A3",X"A3",X"A2",X"A2",X"A1",X"A1",X"A0",X"9F",X"9E",X"9D",X"9C",X"9B",
		X"9A",X"99",X"98",X"97",X"96",X"95",X"93",X"92",X"91",X"90",X"8E",X"8D",X"8B",X"8A",X"89",X"87",
		X"85",X"84",X"83",X"81",X"80",X"7E",X"7D",X"7B",X"7A",X"78",X"77",X"76",X"74",X"73",X"72",X"70",
		X"6F",X"6E",X"6D",X"6C",X"6A",X"6A",X"69",X"68",X"67",X"66",X"65",X"64",X"64",X"63",X"62",X"62",
		X"61",X"61",X"60",X"60",X"60",X"60",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"60",X"60",X"60",X"61",
		X"61",X"61",X"62",X"62",X"63",X"64",X"64",X"65",X"66",X"67",X"68",X"69",X"69",X"6A",X"6B",X"6C",
		X"6E",X"6F",X"70",X"71",X"72",X"73",X"74",X"76",X"77",X"78",X"79",X"7A",X"7C",X"7D",X"7E",X"7F",
		X"81",X"82",X"83",X"84",X"85",X"87",X"88",X"89",X"8A",X"8B",X"8C",X"8D",X"8E",X"8F",X"90",X"91",
		X"92",X"93",X"93",X"94",X"95",X"96",X"96",X"97",X"97",X"98",X"98",X"99",X"99",X"99",X"9A",X"9A",
		X"9A",X"9B",X"9B",X"9A",X"9B",X"9A",X"9A",X"9A",X"9A",X"9A",X"99",X"99",X"99",X"98",X"98",X"97",
		X"97",X"96",X"95",X"95",X"94",X"93",X"93",X"92",X"91",X"90",X"8F",X"8E",X"8D",X"8D",X"8B",X"8A",
		X"8A",X"88",X"87",X"86",X"85",X"84",X"83",X"82",X"81",X"80",X"7F",X"7E",X"7D",X"7C",X"7B",X"7A",
		X"79",X"78",X"77",X"76",X"75",X"74",X"73",X"72",X"71",X"70",X"6F",X"6F",X"6E",X"6D",X"6D",X"6C",
		X"6B",X"6B",X"6A",X"6A",X"69",X"69",X"69",X"68",X"68",X"68",X"68",X"68",X"67",X"68",X"67",X"68",
		X"68",X"68",X"68",X"68",X"68",X"68",X"69",X"69",X"69",X"6A",X"6B",X"6B",X"6C",X"6C",X"6D",X"6D",
		X"6E",X"6F",X"6F",X"70",X"71",X"72",X"72",X"73",X"74",X"75",X"76",X"77",X"78",X"79",X"7A",X"7B",
		X"7C",X"7D",X"7D",X"7E",X"7F",X"80",X"81",X"82",X"83",X"84",X"85",X"86",X"87",X"87",X"88",X"89",
		X"8A",X"8B",X"8B",X"8C",X"8D",X"8D",X"8E",X"8F",X"8F",X"90",X"90",X"91",X"91",X"92",X"92",X"92",
		X"92",X"93",X"93",X"93",X"93",X"93",X"94",X"94",X"94",X"94",X"94",X"93",X"93",X"93",X"93",X"93",
		X"92",X"92",X"92",X"91",X"91",X"91",X"90",X"90",X"8F",X"8F",X"8E",X"8D",X"8D",X"8C",X"8B",X"8B",
		X"8A",X"89",X"89",X"88",X"87",X"86",X"86",X"85",X"84",X"83",X"82",X"82",X"81",X"80",X"7F",X"7E",
		X"7E",X"7D",X"7C",X"7B",X"7B",X"7A",X"79",X"78",X"78",X"77",X"76",X"76",X"75",X"75",X"74",X"74",
		X"73",X"73",X"72",X"72",X"71",X"71",X"70",X"70",X"70",X"70",X"6F",X"6F",X"6F",X"6F",X"6E",X"6E",
		X"6E",X"6E",X"6E",X"6E",X"6E",X"6E",X"6E",X"6F",X"6F",X"6F",X"6F",X"6F",X"70",X"70",X"70",X"70",
		X"71",X"71",X"72",X"72",X"73",X"73",X"74",X"74",X"75",X"75",X"76",X"76",X"77",X"78",X"78",X"79",
		X"79",X"7A",X"7B",X"7B",X"7C",X"7D",X"7D",X"7E",X"7F",X"7F",X"80",X"81",X"81",X"82",X"83",X"83",
		X"84",X"84",X"85",X"86",X"86",X"87",X"87",X"88",X"88",X"89",X"89",X"8A",X"8A",X"8B",X"8B",X"8C",
		X"8C",X"8C",X"8D",X"8D",X"8D",X"8E",X"8E",X"8E",X"8E",X"8E",X"8E",X"8E",X"8F",X"8F",X"8F",X"8E",
		X"8E",X"8E",X"8E",X"8E",X"8E",X"8E",X"8E",X"8D",X"8D",X"8D",X"8D",X"8C",X"8C",X"8C",X"8B",X"8B",
		X"8A",X"8A",X"89",X"89",X"88",X"88",X"87",X"87",X"86",X"85",X"85",X"84",X"84",X"83",X"83",X"82",
		X"81",X"81",X"80",X"80",X"7F",X"7E",X"7E",X"7D",X"7D",X"7C",X"7C",X"7B",X"7A",X"7A",X"79",X"79",
		X"78",X"78",X"77",X"77",X"76",X"76",X"76",X"75",X"75",X"75",X"74",X"74",X"74",X"73",X"73",X"73",
		X"73",X"72",X"72",X"72",X"72",X"72",X"72",X"72",X"72",X"72",X"72",X"72",X"73",X"73",X"73",X"73",
		X"73",X"73",X"74",X"74",X"74",X"75",X"75",X"75",X"76",X"76",X"76",X"77",X"77",X"78",X"78",X"78",
		X"79",X"79",X"7A",X"7A",X"7B",X"7B",X"7C",X"7C",X"7D",X"7D",X"7E",X"7E",X"7F",X"7F",X"80",X"80",
		X"81",X"81",X"82",X"82",X"83",X"83",X"84",X"84",X"84",X"85",X"85",X"86",X"86",X"86",X"87",X"87",
		X"87",X"88",X"88",X"88",X"88",X"89",X"89",X"89",X"89",X"89",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",
		X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",X"89",X"89",X"89",X"89",X"88",
		X"88",X"88",X"88",X"87",X"87",X"87",X"87",X"86",X"86",X"86",X"85",X"85",X"84",X"84",X"84",X"83",
		X"83",X"82",X"82",X"82",X"81",X"81",X"80",X"80",X"80",X"7F",X"7F",X"7E",X"7E",X"7E",X"7D",X"7D",
		X"7C",X"7C",X"7C",X"7B",X"7B",X"7A",X"7A",X"7A",X"79",X"79",X"79",X"78",X"78",X"78",X"78",X"77",
		X"77",X"77",X"77",X"76",X"76",X"76",X"76",X"76",X"76",X"76",X"75",X"75",X"75",X"75",X"75",X"76",
		X"75",X"76",X"76",X"76",X"76",X"76",X"76",X"76",X"76",X"77",X"77",X"77",X"77",X"78",X"78",X"78",
		X"79",X"79",X"79",X"7A",X"7A",X"7A",X"7A",X"7B",X"7B",X"7C",X"7C",X"7C",X"7D",X"7D",X"7D",X"7E",
		X"7E",X"7F",X"7F",X"80",X"80",X"80",X"81",X"81",X"82",X"82",X"82",X"83",X"83",X"83",X"84",X"84",
		X"84",X"85",X"85",X"85",X"85",X"86",X"86",X"86",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"87",X"87",X"87",X"87",
		X"87",X"87",X"87",X"86",X"86",X"86",X"86",X"86",X"85",X"85",X"85",X"85",X"84",X"84",X"84",X"83",
		X"83",X"83",X"82",X"82",X"82",X"82",X"81",X"81",X"81",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7E",
		X"7E",X"7E",X"7D",X"7D",X"7D",X"7C",X"7C",X"7C",X"7C",X"7B",X"7B",X"7B",X"7B",X"7B",X"7A",X"7A",
		X"7A",X"7A",X"7A",X"7A",X"79",X"79",X"79",X"79",X"79",X"79",X"79",X"79",X"79",X"79",X"79",X"79",
		X"79",X"79",X"79",X"79",X"79",X"79",X"79",X"79",X"79",X"79",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",
		X"7A",X"7A",X"7A",X"7B",X"7B",X"7B",X"7B",X"7B",X"7C",X"7C",X"7C",X"7C",X"7D",X"7D",X"7D",X"7D",
		X"7E",X"7E",X"7E",X"7E",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"81",X"81",X"81",X"81",
		X"81",X"82",X"82",X"82",X"82",X"83",X"83",X"83",X"83",X"83",X"83",X"84",X"84",X"84",X"84",X"84",
		X"84",X"84",X"84",X"85",X"85",X"85",X"85",X"85",X"85",X"85",X"85",X"85",X"85",X"85",X"85",X"85",
		X"85",X"85",X"85",X"85",X"85",X"85",X"85",X"85",X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"84",
		X"83",X"83",X"83",X"83",X"83",X"83",X"82",X"82",X"82",X"82",X"81",X"81",X"81",X"81",X"80",X"80",
		X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7E",X"7E",X"7E",X"7E",X"7E",X"7D",X"7D",X"7D",X"7D",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7A",
		X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",
		X"7A",X"7A",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7C",X"7C",X"7C",X"7C",X"7C",X"7D",X"7D",
		X"7D",X"7D",X"7D",X"7E",X"7E",X"7E",X"7E",X"7E",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",
		X"80",X"81",X"81",X"81",X"81",X"81",X"81",X"82",X"82",X"82",X"82",X"82",X"82",X"83",X"83",X"83",
		X"83",X"83",X"83",X"83",X"83",X"83",X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"84",
		X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"83",X"83",X"83",X"83",X"83",X"83",
		X"83",X"83",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"81",X"81",X"81",X"81",X"81",X"81",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7E",X"7E",X"7E",
		X"7E",X"7E",X"7E",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7D",X"7D",X"7D",
		X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"83",X"83",X"83",
		X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",
		X"83",X"83",X"83",X"83",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",
		X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",
		X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7E",X"7E",X"7E",X"7E",
		X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"82",X"81",X"81",X"81",X"81",X"81",X"81",
		X"82",X"81",X"81",X"82",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7D",X"7E",X"7E",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7E",
		X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"7E",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7E",X"7E",X"7E",X"7E",
		X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"7E",X"7E",X"7E",X"7E",X"7E",X"7F",X"80",X"7F",X"80",X"7F",X"80",X"7F",X"7F",X"7F",X"80",X"7F",
		X"80",X"00",X"52",X"49",X"46",X"46",X"F8",X"07",X"00",X"00",X"57",X"41",X"56",X"45",X"66",X"6D",
		X"74",X"20",X"10",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"11",X"2B",X"00",X"00",X"11",X"2B",
		X"00",X"00",X"01",X"00",X"08",X"00",X"64",X"61",X"74",X"61",X"D3",X"07",X"00",X"00",X"80",X"80",
		X"80",X"80",X"81",X"80",X"81",X"80",X"81",X"80",X"81",X"7F",X"81",X"7F",X"81",X"7F",X"81",X"7F",
		X"81",X"7F",X"81",X"7E",X"81",X"7B",X"23",X"13",X"1B",X"18",X"1E",X"1B",X"21",X"1E",X"23",X"22",
		X"26",X"26",X"29",X"29",X"2D",X"3C",X"57",X"79",X"A1",X"CE",X"DB",X"D7",X"D7",X"D4",X"D3",X"D1",
		X"D0",X"CE",X"CD",X"CB",X"C9",X"C8",X"C7",X"C5",X"C4",X"C3",X"C1",X"C0",X"BF",X"BD",X"BC",X"BB",
		X"BA",X"B9",X"B8",X"B7",X"B6",X"B4",X"B3",X"B2",X"B1",X"B0",X"AF",X"AE",X"AD",X"AC",X"AC",X"AB",
		X"AA",X"A9",X"A8",X"A7",X"A6",X"A6",X"A4",X"A1",X"9C",X"96",X"8E",X"85",X"7B",X"70",X"65",X"5A",
		X"4F",X"45",X"3A",X"31",X"29",X"22",X"1D",X"19",X"17",X"16",X"17",X"1A",X"1E",X"25",X"2C",X"35",
		X"3F",X"4A",X"55",X"61",X"6D",X"79",X"85",X"90",X"9B",X"A4",X"AC",X"B3",X"B9",X"BC",X"BC",X"BA",
		X"B9",X"B7",X"B4",X"AF",X"A9",X"A1",X"99",X"90",X"87",X"7D",X"73",X"6A",X"60",X"58",X"50",X"49",
		X"43",X"3E",X"3B",X"38",X"38",X"38",X"3A",X"3E",X"43",X"49",X"50",X"58",X"61",X"6A",X"74",X"7E",
		X"87",X"91",X"99",X"A2",X"A9",X"AF",X"B4",X"B8",X"BB",X"BD",X"BD",X"BB",X"B9",X"B5",X"B0",X"AA",
		X"A3",X"9B",X"93",X"8A",X"81",X"78",X"70",X"67",X"5F",X"58",X"52",X"4D",X"49",X"46",X"44",X"44",
		X"45",X"47",X"4A",X"4F",X"54",X"5B",X"62",X"6A",X"72",X"7A",X"83",X"8B",X"93",X"9B",X"A2",X"A8",
		X"AE",X"B2",X"B5",X"B7",X"B8",X"B7",X"B6",X"B3",X"AF",X"AB",X"A5",X"9E",X"97",X"90",X"88",X"80",
		X"78",X"70",X"69",X"62",X"5C",X"57",X"52",X"4F",X"4D",X"4B",X"4B",X"4C",X"4F",X"52",X"56",X"5B",
		X"61",X"68",X"6F",X"76",X"7E",X"86",X"8D",X"94",X"9B",X"A1",X"A6",X"AB",X"AE",X"B1",X"B2",X"B2",
		X"B2",X"B0",X"AD",X"AA",X"A5",X"A0",X"9A",X"93",X"8C",X"85",X"7E",X"77",X"70",X"6A",X"64",X"5E",
		X"5A",X"56",X"53",X"52",X"51",X"51",X"52",X"54",X"57",X"5C",X"60",X"66",X"6C",X"72",X"79",X"80",
		X"86",X"8D",X"93",X"99",X"9E",X"A3",X"A7",X"A9",X"AB",X"AC",X"AC",X"AB",X"A9",X"A7",X"A3",X"9F",
		X"9A",X"95",X"8F",X"88",X"82",X"7C",X"75",X"6F",X"6A",X"64",X"60",X"5C",X"59",X"57",X"56",X"55",
		X"56",X"57",X"59",X"5C",X"60",X"65",X"6A",X"6F",X"75",X"7B",X"81",X"87",X"8D",X"93",X"98",X"9C",
		X"A0",X"A3",X"A6",X"A8",X"A8",X"A8",X"A7",X"A5",X"A3",X"9F",X"9B",X"96",X"91",X"8C",X"86",X"81",
		X"7B",X"75",X"70",X"6B",X"66",X"62",X"5F",X"5D",X"5B",X"5A",X"5A",X"5A",X"5C",X"5E",X"61",X"65",
		X"69",X"6E",X"73",X"78",X"7D",X"83",X"88",X"8D",X"92",X"96",X"9A",X"9D",X"A0",X"A2",X"A3",X"A4",
		X"A3",X"A2",X"A0",X"9E",X"9B",X"97",X"92",X"8E",X"89",X"84",X"7E",X"79",X"74",X"6F",X"6B",X"67",
		X"64",X"61",X"5F",X"5E",X"5D",X"5D",X"5E",X"5F",X"62",X"65",X"68",X"6C",X"70",X"75",X"7A",X"7F",
		X"84",X"88",X"8D",X"91",X"95",X"99",X"9B",X"9D",X"9F",X"A0",X"A0",X"9F",X"9E",X"9D",X"9A",X"97",
		X"94",X"90",X"8C",X"87",X"82",X"7E",X"79",X"75",X"70",X"6D",X"69",X"66",X"64",X"62",X"61",X"61",
		X"61",X"62",X"63",X"66",X"68",X"6B",X"6F",X"73",X"77",X"7C",X"80",X"85",X"89",X"8D",X"90",X"94",
		X"97",X"99",X"9B",X"9C",X"9C",X"9C",X"9C",X"9A",X"99",X"96",X"94",X"91",X"8D",X"89",X"85",X"80",
		X"7C",X"78",X"74",X"70",X"6D",X"6A",X"68",X"66",X"64",X"63",X"63",X"63",X"64",X"66",X"68",X"6B",
		X"6E",X"71",X"75",X"79",X"7D",X"81",X"85",X"89",X"8C",X"90",X"93",X"95",X"97",X"98",X"99",X"9A",
		X"9A",X"99",X"98",X"96",X"94",X"91",X"8E",X"8B",X"87",X"84",X"80",X"7C",X"78",X"75",X"71",X"6F",
		X"6C",X"6A",X"68",X"67",X"67",X"66",X"67",X"68",X"69",X"6C",X"6E",X"71",X"74",X"77",X"7B",X"7E",
		X"82",X"86",X"89",X"8C",X"8F",X"92",X"94",X"95",X"97",X"97",X"98",X"97",X"96",X"95",X"93",X"91",
		X"8F",X"8C",X"89",X"85",X"82",X"7F",X"7B",X"78",X"75",X"72",X"6F",X"6D",X"6B",X"6A",X"69",X"68",
		X"68",X"69",X"6A",X"6B",X"6D",X"70",X"72",X"75",X"78",X"7C",X"7F",X"82",X"86",X"89",X"8B",X"8E",
		X"90",X"92",X"93",X"95",X"95",X"95",X"95",X"94",X"93",X"91",X"8F",X"8D",X"8A",X"87",X"84",X"81",
		X"7E",X"7B",X"78",X"75",X"73",X"70",X"6F",X"6D",X"6C",X"6B",X"6A",X"6B",X"6B",X"6D",X"6E",X"70",
		X"72",X"75",X"78",X"7A",X"7D",X"80",X"83",X"86",X"89",X"8B",X"8E",X"90",X"91",X"92",X"93",X"93",
		X"93",X"93",X"92",X"91",X"8F",X"8D",X"8B",X"88",X"86",X"83",X"80",X"7D",X"7A",X"78",X"75",X"73",
		X"71",X"6F",X"6E",X"6D",X"6C",X"6C",X"6C",X"6D",X"6E",X"70",X"71",X"73",X"76",X"78",X"7B",X"7E",
		X"80",X"83",X"86",X"88",X"8B",X"8C",X"8E",X"8F",X"90",X"91",X"91",X"91",X"91",X"90",X"8E",X"8D",
		X"8B",X"89",X"87",X"84",X"82",X"7F",X"7D",X"7A",X"78",X"76",X"74",X"72",X"71",X"70",X"6F",X"6E",
		X"6E",X"6F",X"6F",X"70",X"72",X"74",X"76",X"78",X"7A",X"7D",X"7F",X"82",X"84",X"86",X"89",X"8B",
		X"8C",X"8E",X"8F",X"90",X"90",X"90",X"90",X"8F",X"8E",X"8D",X"8C",X"8A",X"88",X"86",X"84",X"81",
		X"7F",X"7C",X"7A",X"78",X"76",X"74",X"73",X"71",X"70",X"70",X"70",X"70",X"70",X"71",X"72",X"73",
		X"75",X"77",X"79",X"7B",X"7D",X"7F",X"82",X"84",X"86",X"88",X"8A",X"8B",X"8C",X"8D",X"8E",X"8E",
		X"8E",X"8E",X"8D",X"8C",X"8B",X"8A",X"88",X"87",X"85",X"83",X"80",X"7E",X"7C",X"7A",X"78",X"76",
		X"75",X"73",X"72",X"71",X"71",X"71",X"71",X"72",X"72",X"74",X"75",X"76",X"78",X"7A",X"7C",X"7E",
		X"80",X"82",X"85",X"86",X"88",X"8A",X"8B",X"8C",X"8D",X"8D",X"8E",X"8D",X"8D",X"8D",X"8C",X"8A",
		X"89",X"87",X"86",X"84",X"82",X"80",X"7E",X"7C",X"7A",X"78",X"77",X"75",X"74",X"73",X"72",X"72",
		X"72",X"72",X"73",X"73",X"75",X"76",X"77",X"79",X"7B",X"7D",X"7E",X"80",X"82",X"84",X"86",X"87",
		X"89",X"8A",X"8B",X"8B",X"8C",X"8C",X"8C",X"8B",X"8B",X"8A",X"89",X"87",X"86",X"84",X"83",X"81",
		X"7F",X"7D",X"7C",X"7A",X"78",X"77",X"76",X"74",X"74",X"73",X"73",X"73",X"73",X"74",X"75",X"76",
		X"77",X"79",X"7A",X"7C",X"7E",X"7F",X"81",X"83",X"84",X"86",X"88",X"89",X"8A",X"8B",X"8B",X"8B",
		X"8B",X"8B",X"8B",X"8A",X"89",X"88",X"87",X"86",X"84",X"82",X"81",X"7F",X"7E",X"7C",X"7A",X"79",
		X"78",X"76",X"75",X"75",X"74",X"74",X"74",X"75",X"75",X"76",X"77",X"78",X"79",X"7B",X"7D",X"7E",
		X"80",X"81",X"83",X"84",X"86",X"87",X"88",X"89",X"89",X"8A",X"8A",X"8A",X"8A",X"89",X"89",X"88",
		X"87",X"86",X"84",X"83",X"81",X"80",X"7E",X"7D",X"7B",X"7A",X"79",X"78",X"77",X"76",X"75",X"75",
		X"75",X"75",X"76",X"76",X"77",X"78",X"79",X"7A",X"7C",X"7D",X"7F",X"80",X"82",X"83",X"85",X"86",
		X"87",X"88",X"88",X"89",X"89",X"89",X"89",X"89",X"89",X"88",X"87",X"86",X"85",X"84",X"82",X"81",
		X"80",X"7E",X"7D",X"7C",X"7A",X"79",X"78",X"78",X"77",X"77",X"76",X"76",X"77",X"77",X"78",X"78",
		X"79",X"7A",X"7B",X"7D",X"7E",X"7F",X"80",X"82",X"83",X"84",X"85",X"86",X"87",X"87",X"88",X"88",
		X"88",X"88",X"87",X"87",X"86",X"86",X"84",X"84",X"82",X"81",X"80",X"7F",X"7E",X"7C",X"7B",X"7A",
		X"79",X"78",X"78",X"77",X"77",X"77",X"77",X"77",X"78",X"78",X"79",X"7A",X"7B",X"7C",X"7D",X"7E",
		X"7F",X"80",X"82",X"83",X"84",X"85",X"86",X"86",X"87",X"87",X"87",X"87",X"87",X"87",X"86",X"86",
		X"85",X"84",X"83",X"82",X"81",X"80",X"7F",X"7E",X"7D",X"7C",X"7B",X"7A",X"7A",X"79",X"79",X"78",
		X"78",X"79",X"79",X"79",X"7A",X"7A",X"7B",X"7C",X"7D",X"7E",X"7F",X"80",X"81",X"82",X"83",X"84",
		X"84",X"85",X"86",X"86",X"86",X"86",X"86",X"86",X"86",X"85",X"85",X"84",X"83",X"82",X"82",X"80",
		X"7F",X"7E",X"7D",X"7D",X"7C",X"7B",X"7A",X"7A",X"79",X"79",X"79",X"79",X"79",X"79",X"7A",X"7A",
		X"7B",X"7B",X"7C",X"7D",X"7E",X"7F",X"80",X"81",X"82",X"82",X"83",X"84",X"84",X"85",X"85",X"86",
		X"86",X"86",X"85",X"85",X"85",X"84",X"84",X"83",X"82",X"81",X"80",X"80",X"7F",X"7E",X"7D",X"7C",
		X"7C",X"7B",X"7B",X"7A",X"7A",X"7A",X"7A",X"7A",X"7B",X"7B",X"7B",X"7C",X"7D",X"7D",X"7E",X"7F",
		X"80",X"80",X"81",X"82",X"82",X"83",X"84",X"84",X"84",X"85",X"85",X"85",X"85",X"85",X"84",X"84",
		X"83",X"83",X"82",X"81",X"80",X"80",X"7F",X"7E",X"7D",X"7D",X"7C",X"7C",X"7B",X"7B",X"7A",X"7A",
		X"7A",X"7A",X"7A",X"7B",X"7B",X"7B",X"7C",X"7D",X"7D",X"7E",X"7F",X"7F",X"80",X"81",X"81",X"82",
		X"82",X"83",X"83",X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"83",X"83",X"82",X"82",X"81",X"80",
		X"80",X"7F",X"7E",X"7E",X"7D",X"7D",X"7C",X"7C",X"7C",X"7B",X"7B",X"7B",X"7B",X"7C",X"7C",X"7C",
		X"7D",X"7D",X"7E",X"7E",X"7F",X"7F",X"80",X"81",X"81",X"82",X"82",X"83",X"83",X"83",X"84",X"84",
		X"84",X"84",X"84",X"83",X"83",X"83",X"82",X"82",X"81",X"81",X"80",X"80",X"7F",X"7E",X"7E",X"7D",
		X"7D",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7D",X"7D",X"7E",X"7E",X"7F",
		X"7F",X"80",X"80",X"81",X"81",X"82",X"82",X"82",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"82",
		X"82",X"82",X"81",X"81",X"80",X"80",X"7F",X"7F",X"7E",X"7E",X"7E",X"7D",X"7D",X"7D",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7D",X"7D",X"7D",X"7E",X"7E",X"7E",X"7F",X"7F",X"80",X"80",X"81",X"81",X"82",
		X"82",X"82",X"82",X"83",X"83",X"83",X"83",X"83",X"83",X"82",X"82",X"82",X"81",X"81",X"81",X"80",
		X"80",X"7F",X"7F",X"7F",X"7E",X"7E",X"7D",X"7D",X"7D",X"7C",X"7C",X"7C",X"7C",X"7D",X"7D",X"7D",
		X"7D",X"7D",X"7E",X"7E",X"7E",X"7F",X"7F",X"80",X"80",X"81",X"81",X"81",X"81",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"81",X"81",X"81",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7E",X"7E",
		X"7E",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7E",X"7E",X"7E",X"7E",X"7F",X"7F",
		X"7F",X"80",X"80",X"81",X"81",X"81",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"81",X"81",X"81",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"7D",X"7E",X"7E",X"7D",X"7E",X"7E",X"7E",X"7E",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"80",X"80",X"80",X"80",
		X"7F",X"7F",X"7F",X"7F",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7D",X"7E",X"7E",X"7E",X"7E",
		X"7E",X"7E",X"7E",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"81",X"81",X"81",X"81",X"81",X"81",X"82",
		X"82",X"82",X"82",X"81",X"81",X"81",X"81",X"81",X"81",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",
		X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"80",X"80",X"80",X"80",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"80",X"80",X"80",
		X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"7E",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"81",X"81",X"81",X"81",X"81",X"81",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7E",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"00",X"52",X"49",X"46",X"46",X"D6",X"07",X"00",X"00",X"57",X"41",X"56",X"45",X"66",X"6D",
		X"74",X"20",X"10",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"11",X"2B",X"00",X"00",X"11",X"2B",
		X"00",X"00",X"01",X"00",X"08",X"00",X"64",X"61",X"74",X"61",X"B2",X"07",X"00",X"00",X"81",X"83",
		X"80",X"80",X"7E",X"7F",X"80",X"7F",X"81",X"81",X"81",X"82",X"83",X"7F",X"83",X"7D",X"84",X"7B",
		X"8B",X"44",X"01",X"12",X"09",X"13",X"0F",X"14",X"10",X"12",X"16",X"18",X"1B",X"21",X"22",X"24",
		X"2B",X"4D",X"7A",X"B7",X"E9",X"E5",X"E6",X"E2",X"E1",X"DE",X"DB",X"DB",X"D8",X"D4",X"D4",X"D2",
		X"D4",X"CE",X"C9",X"CC",X"C9",X"C6",X"C9",X"C9",X"C1",X"C0",X"C0",X"BF",X"BE",X"BB",X"B9",X"B9",
		X"B9",X"B8",X"B4",X"B3",X"B4",X"B3",X"B1",X"B1",X"B0",X"AE",X"AD",X"AC",X"AC",X"AB",X"AA",X"A9",
		X"A8",X"A6",X"A4",X"A1",X"99",X"8F",X"84",X"76",X"68",X"59",X"4A",X"3A",X"2C",X"20",X"15",X"0D",
		X"07",X"04",X"03",X"05",X"09",X"11",X"1B",X"28",X"36",X"46",X"56",X"67",X"78",X"88",X"97",X"A5",
		X"B0",X"BA",X"C0",X"C0",X"BE",X"BC",X"B9",X"B4",X"AC",X"A2",X"96",X"89",X"7C",X"6E",X"61",X"54",
		X"48",X"3E",X"35",X"2F",X"2A",X"28",X"28",X"2B",X"30",X"37",X"41",X"4C",X"58",X"65",X"73",X"81",
		X"8E",X"9A",X"A6",X"B0",X"B8",X"BF",X"C3",X"C5",X"C4",X"C2",X"BD",X"B6",X"AD",X"A3",X"98",X"8B",
		X"7F",X"73",X"67",X"5B",X"51",X"49",X"41",X"3C",X"39",X"38",X"39",X"3D",X"42",X"49",X"52",X"5D",
		X"68",X"74",X"80",X"8C",X"98",X"A2",X"AC",X"B4",X"BB",X"BF",X"C2",X"C2",X"C0",X"BD",X"B8",X"B0",
		X"A7",X"9D",X"92",X"86",X"7B",X"6F",X"64",X"5B",X"52",X"4A",X"45",X"41",X"3F",X"3F",X"41",X"45",
		X"4B",X"53",X"5C",X"66",X"71",X"7C",X"88",X"93",X"9D",X"A6",X"AE",X"B4",X"B9",X"BC",X"BD",X"BC",
		X"B9",X"B5",X"AF",X"A7",X"9E",X"94",X"8A",X"7F",X"74",X"6A",X"60",X"58",X"51",X"4B",X"47",X"45",
		X"44",X"46",X"49",X"4E",X"55",X"5D",X"66",X"70",X"7A",X"84",X"8F",X"98",X"A1",X"A9",X"AF",X"B4",
		X"B8",X"B9",X"B9",X"B7",X"B3",X"AE",X"A7",X"A0",X"97",X"8D",X"83",X"79",X"70",X"67",X"5F",X"58",
		X"52",X"4E",X"4B",X"4A",X"4A",X"4C",X"50",X"56",X"5C",X"64",X"6D",X"76",X"7F",X"89",X"92",X"9A",
		X"A2",X"A8",X"AD",X"B1",X"B3",X"B3",X"B2",X"AF",X"AB",X"A6",X"9F",X"97",X"8E",X"85",X"7C",X"73",
		X"6B",X"63",X"5C",X"56",X"51",X"4E",X"4D",X"4D",X"4E",X"51",X"56",X"5B",X"62",X"6A",X"73",X"7B",
		X"84",X"8C",X"94",X"9C",X"A2",X"A7",X"AB",X"AD",X"AF",X"AE",X"AC",X"AA",X"A5",X"A0",X"99",X"91",
		X"89",X"81",X"79",X"71",X"69",X"62",X"5C",X"57",X"54",X"52",X"51",X"51",X"54",X"57",X"5C",X"62",
		X"69",X"70",X"78",X"80",X"89",X"90",X"97",X"9E",X"A3",X"A7",X"AA",X"AC",X"AC",X"AA",X"A8",X"A5",
		X"A0",X"99",X"93",X"8B",X"84",X"7C",X"74",X"6D",X"66",X"60",X"5C",X"58",X"56",X"54",X"54",X"56",
		X"59",X"5D",X"62",X"68",X"6F",X"76",X"7D",X"85",X"8C",X"93",X"98",X"9E",X"A2",X"A5",X"A7",X"A8",
		X"A7",X"A5",X"A2",X"9E",X"99",X"93",X"8C",X"85",X"7E",X"77",X"70",X"6A",X"65",X"60",X"5C",X"59",
		X"58",X"57",X"58",X"5B",X"5E",X"62",X"68",X"6E",X"74",X"7B",X"82",X"89",X"90",X"95",X"9B",X"9F",
		X"A2",X"A4",X"A6",X"A6",X"A4",X"A2",X"9F",X"9B",X"95",X"90",X"89",X"83",X"7C",X"75",X"6F",X"6A",
		X"65",X"61",X"5E",X"5C",X"5B",X"5B",X"5D",X"5F",X"63",X"68",X"6D",X"73",X"79",X"7F",X"85",X"8C",
		X"91",X"96",X"9B",X"9E",X"A0",X"A2",X"A2",X"A2",X"A0",X"9D",X"9A",X"95",X"90",X"8A",X"84",X"7E",
		X"78",X"72",X"6C",X"68",X"64",X"61",X"5F",X"5D",X"5D",X"5E",X"60",X"62",X"66",X"6B",X"70",X"76",
		X"7C",X"82",X"88",X"8D",X"92",X"96",X"9A",X"9D",X"9E",X"A0",X"9F",X"9E",X"9C",X"99",X"96",X"91",
		X"8C",X"86",X"81",X"7B",X"75",X"70",X"6C",X"67",X"64",X"62",X"60",X"5F",X"60",X"61",X"63",X"67",
		X"6B",X"70",X"75",X"7A",X"80",X"85",X"8B",X"90",X"94",X"98",X"9B",X"9D",X"9E",X"9E",X"9D",X"9C",
		X"9A",X"96",X"92",X"8D",X"88",X"83",X"7E",X"78",X"73",X"6F",X"6A",X"67",X"65",X"63",X"62",X"62",
		X"62",X"65",X"68",X"6B",X"6F",X"74",X"79",X"7E",X"83",X"88",X"8D",X"91",X"94",X"97",X"99",X"9B",
		X"9B",X"9A",X"99",X"97",X"95",X"91",X"8D",X"88",X"83",X"7E",X"79",X"74",X"70",X"6C",X"69",X"66",
		X"64",X"63",X"63",X"64",X"65",X"68",X"6B",X"6F",X"73",X"78",X"7D",X"82",X"87",X"8B",X"90",X"93",
		X"97",X"98",X"9A",X"9B",X"9A",X"9A",X"98",X"96",X"93",X"8F",X"8B",X"86",X"81",X"7C",X"78",X"74",
		X"70",X"6C",X"6A",X"68",X"66",X"65",X"66",X"67",X"69",X"6C",X"6F",X"73",X"77",X"7C",X"81",X"85",
		X"89",X"8E",X"91",X"94",X"97",X"98",X"99",X"99",X"99",X"97",X"95",X"93",X"90",X"8B",X"87",X"83",
		X"7E",X"79",X"75",X"71",X"6D",X"6B",X"69",X"67",X"66",X"66",X"67",X"68",X"6B",X"6E",X"71",X"75",
		X"79",X"7E",X"82",X"86",X"8A",X"8E",X"91",X"94",X"96",X"96",X"97",X"97",X"96",X"94",X"92",X"8F",
		X"8B",X"88",X"83",X"7F",X"7B",X"77",X"73",X"70",X"6D",X"6B",X"69",X"68",X"67",X"68",X"69",X"6B",
		X"6E",X"71",X"74",X"78",X"7D",X"81",X"85",X"89",X"8C",X"90",X"92",X"95",X"96",X"97",X"97",X"96",
		X"95",X"92",X"90",X"8D",X"8A",X"86",X"82",X"7E",X"7A",X"76",X"73",X"70",X"6D",X"6B",X"6A",X"69",
		X"69",X"6A",X"6B",X"6D",X"70",X"73",X"77",X"7B",X"7F",X"83",X"86",X"8A",X"8D",X"90",X"92",X"94",
		X"95",X"95",X"94",X"93",X"92",X"90",X"8D",X"8A",X"87",X"83",X"7F",X"7B",X"77",X"74",X"71",X"6E",
		X"6C",X"6B",X"6A",X"69",X"6A",X"6B",X"6D",X"6F",X"72",X"75",X"79",X"7D",X"81",X"84",X"88",X"8B",
		X"8E",X"90",X"92",X"94",X"94",X"94",X"93",X"92",X"90",X"8E",X"8C",X"88",X"85",X"82",X"7E",X"7A",
		X"77",X"74",X"72",X"6F",X"6E",X"6D",X"6C",X"6C",X"6D",X"6F",X"70",X"73",X"76",X"79",X"7D",X"80",
		X"84",X"87",X"8A",X"8D",X"8F",X"91",X"93",X"93",X"93",X"93",X"92",X"90",X"8E",X"8C",X"89",X"86",
		X"82",X"7F",X"7C",X"78",X"75",X"73",X"70",X"6E",X"6D",X"6C",X"6C",X"6D",X"6E",X"70",X"72",X"75",
		X"78",X"7B",X"7E",X"81",X"84",X"88",X"8A",X"8D",X"8E",X"90",X"91",X"91",X"91",X"90",X"8F",X"8D",
		X"8B",X"89",X"86",X"83",X"80",X"7C",X"79",X"76",X"74",X"72",X"70",X"6E",X"6E",X"6D",X"6D",X"6E",
		X"70",X"72",X"74",X"77",X"7A",X"7D",X"80",X"83",X"86",X"89",X"8C",X"8E",X"8F",X"91",X"91",X"91",
		X"91",X"90",X"8E",X"8D",X"8A",X"88",X"85",X"82",X"7F",X"7C",X"79",X"76",X"74",X"72",X"70",X"6F",
		X"6E",X"6E",X"6F",X"70",X"71",X"74",X"76",X"79",X"7C",X"7F",X"82",X"85",X"88",X"8A",X"8C",X"8E",
		X"8F",X"90",X"90",X"90",X"8F",X"8E",X"8C",X"8A",X"88",X"86",X"83",X"80",X"7D",X"7A",X"77",X"75",
		X"73",X"71",X"70",X"6F",X"6E",X"6F",X"6F",X"71",X"73",X"74",X"77",X"7A",X"7D",X"7F",X"82",X"85",
		X"88",X"8A",X"8C",X"8D",X"8E",X"8F",X"8F",X"8E",X"8D",X"8C",X"8B",X"89",X"87",X"84",X"81",X"7F",
		X"7C",X"79",X"77",X"75",X"74",X"72",X"71",X"70",X"71",X"71",X"73",X"74",X"76",X"78",X"7B",X"7D",
		X"80",X"83",X"85",X"88",X"8A",X"8C",X"8D",X"8E",X"8F",X"8F",X"8F",X"8E",X"8D",X"8B",X"8A",X"88",
		X"85",X"83",X"80",X"7D",X"7B",X"78",X"76",X"74",X"73",X"72",X"71",X"70",X"71",X"71",X"73",X"74",
		X"76",X"79",X"7B",X"7E",X"80",X"83",X"86",X"88",X"8A",X"8C",X"8D",X"8E",X"8E",X"8E",X"8D",X"8C",
		X"8B",X"89",X"87",X"85",X"82",X"80",X"7D",X"7B",X"78",X"76",X"74",X"72",X"71",X"70",X"70",X"70",
		X"71",X"72",X"73",X"75",X"77",X"7A",X"7D",X"7F",X"82",X"84",X"87",X"89",X"8B",X"8C",X"8E",X"8E",
		X"8E",X"8E",X"8D",X"8C",X"8B",X"89",X"87",X"85",X"82",X"80",X"7D",X"7A",X"78",X"76",X"74",X"73",
		X"71",X"71",X"71",X"71",X"72",X"73",X"75",X"77",X"79",X"7C",X"7E",X"81",X"84",X"86",X"89",X"8A",
		X"8C",X"8D",X"8E",X"8E",X"8E",X"8E",X"8C",X"8B",X"89",X"88",X"85",X"83",X"80",X"7E",X"7B",X"79",
		X"76",X"75",X"73",X"71",X"70",X"70",X"70",X"71",X"72",X"74",X"76",X"78",X"7A",X"7D",X"7F",X"82",
		X"84",X"86",X"88",X"8A",X"8B",X"8C",X"8D",X"8D",X"8D",X"8C",X"8B",X"8A",X"88",X"86",X"84",X"82",
		X"7F",X"7D",X"7A",X"78",X"76",X"75",X"73",X"72",X"72",X"72",X"72",X"73",X"74",X"76",X"78",X"7A",
		X"7D",X"7F",X"81",X"84",X"86",X"88",X"8A",X"8B",X"8D",X"8D",X"8E",X"8E",X"8D",X"8C",X"8B",X"89",
		X"88",X"86",X"84",X"82",X"7F",X"7D",X"7A",X"78",X"77",X"75",X"74",X"73",X"73",X"73",X"73",X"74",
		X"75",X"77",X"79",X"7B",X"7D",X"80",X"82",X"84",X"86",X"88",X"89",X"8A",X"8B",X"8C",X"8C",X"8C",
		X"8B",X"8A",X"88",X"87",X"85",X"83",X"81",X"7F",X"7D",X"7A",X"78",X"76",X"75",X"73",X"72",X"72",
		X"72",X"72",X"73",X"74",X"76",X"78",X"7A",X"7C",X"7E",X"81",X"83",X"85",X"87",X"89",X"8A",X"8B",
		X"8C",X"8C",X"8C",X"8B",X"8B",X"89",X"88",X"86",X"84",X"82",X"80",X"7E",X"7C",X"7A",X"78",X"76",
		X"75",X"74",X"73",X"73",X"73",X"74",X"75",X"76",X"78",X"7A",X"7C",X"7E",X"80",X"83",X"85",X"87",
		X"88",X"8A",X"8B",X"8C",X"8C",X"8C",X"8C",X"8B",X"8A",X"88",X"86",X"85",X"83",X"81",X"7E",X"7C",
		X"7A",X"78",X"77",X"75",X"74",X"73",X"73",X"73",X"73",X"74",X"75",X"77",X"79",X"7B",X"7D",X"7F",
		X"81",X"83",X"85",X"87",X"88",X"89",X"8A",X"8B",X"8B",X"8A",X"8A",X"89",X"88",X"86",X"85",X"83",
		X"81",X"80",X"7D",X"7C",X"7A",X"78",X"77",X"75",X"74",X"74",X"74",X"74",X"75",X"76",X"77",X"79",
		X"7B",X"7D",X"7F",X"81",X"83",X"85",X"87",X"88",X"8A",X"8B",X"8B",X"8B",X"8B",X"8B",X"8A",X"89",
		X"88",X"87",X"85",X"83",X"81",X"80",X"7E",X"7C",X"7A",X"78",X"77",X"76",X"75",X"75",X"75",X"75",
		X"76",X"77",X"78",X"7A",X"7C",X"7E",X"80",X"82",X"84",X"85",X"87",X"88",X"89",X"8A",X"8B",X"8B",
		X"8B",X"8A",X"89",X"88",X"86",X"85",X"83",X"81",X"7F",X"7D",X"7B",X"7A",X"78",X"77",X"75",X"74",
		X"74",X"74",X"74",X"75",X"76",X"77",X"78",X"7A",X"7C",X"7E",X"80",X"82",X"84",X"85",X"86",X"88",
		X"89",X"89",X"8A",X"8A",X"89",X"89",X"88",X"86",X"85",X"84",X"82",X"80",X"7E",X"7D",X"7B",X"79",
		X"78",X"77",X"76",X"75",X"75",X"75",X"76",X"77",X"78",X"79",X"7B",X"7C",X"7E",X"80",X"82",X"83",
		X"85",X"87",X"88",X"89",X"89",X"8A",X"8A",X"8A",X"89",X"89",X"87",X"86",X"85",X"83",X"81",X"7F",
		X"7E",X"7C",X"7B",X"79",X"78",X"76",X"76",X"75",X"76",X"76",X"76",X"77",X"78",X"7A",X"7B",X"7D",
		X"7E",X"80",X"82",X"83",X"85",X"86",X"87",X"88",X"88",X"89",X"88",X"88",X"87",X"86",X"85",X"84",
		X"83",X"81",X"7F",X"7E",X"7C",X"7B",X"7A",X"78",X"77",X"77",X"77",X"76",X"76",X"77",X"77",X"79",
		X"7A",X"7B",X"7D",X"7E",X"80",X"82",X"83",X"85",X"86",X"87",X"88",X"88",X"89",X"89",X"88",X"88",
		X"87",X"86",X"85",X"84",X"82",X"81",X"80",X"7E",X"7D",X"7B",X"7A",X"79",X"79",X"78",X"78",X"78",
		X"78",X"79",X"7A",X"7B",X"7C",X"7D",X"7F",X"80",X"81",X"83",X"84",X"85",X"86",X"87",X"87",X"88",
		X"88",X"87",X"87",X"86",X"85",X"84",X"83",X"82",X"81",X"7F",X"7E",X"7D",X"7B",X"7A",X"79",X"79",
		X"78",X"78",X"78",X"78",X"79",X"79",X"7A",X"7B",X"7C",X"7D",X"7E",X"7F",X"81",X"82",X"83",X"84",
		X"85",X"86",X"86",X"86",X"86",X"86",X"85",X"85",X"84",X"83",X"82",X"81",X"80",X"7E",X"7D",X"7C",
		X"7B",X"7A",X"7A",X"79",X"79",X"79",X"79",X"79",X"7A",X"7A",X"7B",X"7C",X"7E",X"7F",X"80",X"81",
		X"82",X"83",X"84",X"85",X"86",X"86",X"87",X"87",X"86",X"86",X"85",X"85",X"84",X"83",X"82",X"81",
		X"80",X"7F",X"7D",X"7C",X"7B",X"7A",X"7A",X"7A",X"79",X"79",X"7A",X"7A",X"7B",X"7B",X"7C",X"7D",
		X"7E",X"7F",X"80",X"81",X"82",X"83",X"84",X"84",X"85",X"85",X"85",X"85",X"85",X"84",X"84",X"83",
		X"82",X"81",X"80",X"7F",X"7E",X"7D",X"7C",X"7B",X"7B",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7B",
		X"7B",X"7C",X"7D",X"7E",X"7F",X"80",X"81",X"82",X"82",X"83",X"84",X"84",X"85",X"85",X"85",X"85",
		X"85",X"84",X"84",X"83",X"82",X"81",X"80",X"7F",X"7F",X"7E",X"7D",X"7C",X"7C",X"7B",X"7B",X"7B",
		X"7B",X"7B",X"7C",X"7C",X"7D",X"7E",X"7F",X"80",X"80",X"81",X"82",X"83",X"83",X"84",X"84",X"85",
		X"85",X"85",X"85",X"85",X"84",X"83",X"83",X"82",X"81",X"80",X"80",X"7F",X"7E",X"7D",X"7C",X"7C",
		X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7C",X"7C",X"7D",X"7E",X"7F",X"7F",X"80",X"81",X"82",
		X"82",X"83",X"83",X"83",X"84",X"83",X"83",X"83",X"83",X"82",X"81",X"81",X"80",X"7F",X"7E",X"7E",
		X"7D",X"7C",X"7C",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7C",X"7C",X"7D",X"7D",X"7E",X"7F",X"80",
		X"81",X"81",X"82",X"82",X"83",X"83",X"84",X"84",X"84",X"84",X"83",X"83",X"83",X"82",X"81",X"81",
		X"80",X"80",X"7F",X"7E",X"7E",X"7D",X"7D",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7D",X"7D",X"7E",
		X"7E",X"7F",X"80",X"80",X"81",X"81",X"82",X"82",X"83",X"83",X"83",X"83",X"83",X"83",X"82",X"82",
		X"82",X"81",X"80",X"7F",X"7F",X"7E",X"7E",X"7D",X"7D",X"7C",X"7C",X"7C",X"7B",X"7C",X"7C",X"7C",
		X"7C",X"7D",X"7D",X"7E",X"7E",X"7F",X"7F",X"80",X"81",X"81",X"82",X"82",X"82",X"82",X"83",X"82",
		X"82",X"82",X"82",X"82",X"81",X"81",X"80",X"80",X"7F",X"7F",X"7E",X"7E",X"7E",X"7D",X"7D",X"7D",
		X"7D",X"7D",X"7D",X"7E",X"7E",X"7E",X"7F",X"7F",X"80",X"80",X"81",X"82",X"82",X"82",X"83",X"83",
		X"83",X"83",X"83",X"83",X"83",X"82",X"82",X"82",X"81",X"81",X"80",X"7F",X"7F",X"7F",X"7E",X"7E",
		X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7E",X"7E",X"7E",X"7F",X"7F",X"80",X"80",X"81",
		X"81",X"81",X"81",X"82",X"81",X"80",X"80",X"80",X"80",X"80",X"7F",X"80",X"7F",X"7F",X"7F",X"7F",
		X"52",X"49",X"46",X"46",X"9A",X"01",X"00",X"00",X"57",X"41",X"56",X"45",X"66",X"6D",X"74",X"20",
		X"10",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"11",X"2B",X"00",X"00",X"11",X"2B",X"00",X"00",
		X"01",X"00",X"08",X"00",X"64",X"61",X"74",X"61",X"75",X"01",X"00",X"00",X"7F",X"80",X"82",X"69",
		X"00",X"4B",X"F9",X"F6",X"F7",X"F3",X"E8",X"AB",X"59",X"12",X"07",X"06",X"25",X"78",X"C7",X"F6",
		X"F3",X"E0",X"A7",X"66",X"2D",X"12",X"17",X"42",X"7D",X"B8",X"DE",X"E4",X"CB",X"98",X"5F",X"31",
		X"1E",X"28",X"52",X"87",X"B9",X"D5",X"D6",X"BB",X"8C",X"5A",X"36",X"28",X"38",X"5F",X"8F",X"B8",
		X"CD",X"C9",X"AE",X"83",X"57",X"3A",X"32",X"44",X"6A",X"94",X"B6",X"C5",X"BE",X"A3",X"7B",X"56",
		X"3F",X"3B",X"4F",X"72",X"98",X"B4",X"BE",X"B4",X"99",X"75",X"56",X"43",X"44",X"59",X"79",X"9B",
		X"B2",X"B7",X"AC",X"92",X"71",X"56",X"48",X"4B",X"61",X"80",X"9D",X"B0",X"B2",X"A5",X"8C",X"6E",
		X"58",X"4C",X"52",X"68",X"84",X"9E",X"AD",X"AC",X"9F",X"87",X"6C",X"59",X"51",X"59",X"6E",X"88",
		X"9F",X"AA",X"A8",X"9A",X"83",X"6B",X"5A",X"54",X"5F",X"73",X"8B",X"9F",X"A8",X"A3",X"95",X"80",
		X"6A",X"5C",X"58",X"63",X"77",X"8E",X"9E",X"A5",X"A0",X"91",X"7D",X"69",X"5D",X"5B",X"68",X"7B",
		X"8F",X"9E",X"A2",X"9B",X"8D",X"7A",X"69",X"5E",X"5E",X"6B",X"7E",X"91",X"9D",X"A0",X"98",X"8A",
		X"78",X"68",X"5F",X"61",X"6E",X"80",X"91",X"9C",X"9D",X"94",X"87",X"76",X"68",X"60",X"64",X"71",
		X"82",X"92",X"9B",X"9B",X"92",X"85",X"75",X"68",X"62",X"68",X"75",X"85",X"92",X"9A",X"98",X"8F",
		X"82",X"75",X"69",X"64",X"6B",X"77",X"86",X"93",X"99",X"96",X"8D",X"80",X"74",X"69",X"67",X"6E",
		X"7A",X"88",X"93",X"97",X"94",X"8A",X"7E",X"72",X"6A",X"6A",X"72",X"7D",X"89",X"92",X"94",X"90",
		X"87",X"7C",X"72",X"6D",X"6E",X"75",X"7F",X"8A",X"90",X"91",X"8D",X"84",X"7A",X"72",X"6F",X"71",
		X"78",X"81",X"89",X"8E",X"8E",X"89",X"82",X"79",X"73",X"71",X"74",X"7A",X"82",X"88",X"8C",X"8B",
		X"86",X"80",X"79",X"74",X"74",X"77",X"7C",X"83",X"88",X"8A",X"88",X"84",X"7E",X"79",X"76",X"76",
		X"79",X"7E",X"84",X"87",X"89",X"87",X"82",X"7D",X"79",X"77",X"78",X"7B",X"7F",X"84",X"86",X"87",
		X"85",X"81",X"7D",X"7A",X"79",X"7A",X"7D",X"80",X"84",X"86",X"86",X"84",X"81",X"7D",X"7B",X"7A",
		X"7B",X"7E",X"81",X"84",X"85",X"85",X"83",X"80",X"7D",X"7B",X"7B",X"7C",X"7F",X"81",X"83",X"84",
		X"83",X"82",X"7F",X"7D",X"7B",X"7B",X"7D",X"7F",X"81",X"83",X"83",X"82",X"81",X"7E",X"7D",X"7C",
		X"7C",X"7D",X"7F",X"81",X"82",X"82",X"81",X"80",X"7E",X"7D",X"7C",X"7D",X"7E",X"7F",X"81",X"82",
		X"82",X"81",X"7F",X"7E",X"7D",X"7C",X"7D",X"7E",X"80",X"81",X"82",X"81",X"81",X"7F",X"7E",X"7D",
		X"7E",X"00",X"52",X"49",X"46",X"46",X"A4",X"13",X"00",X"00",X"57",X"41",X"56",X"45",X"66",X"6D",
		X"74",X"20",X"10",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"11",X"2B",X"00",X"00",X"11",X"2B",
		X"00",X"00",X"01",X"00",X"08",X"00",X"64",X"61",X"74",X"61",X"7F",X"13",X"00",X"00",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"82",X"84",X"88",X"8F",X"98",X"A3",
		X"B0",X"BB",X"C1",X"C3",X"BE",X"B4",X"A5",X"94",X"80",X"6C",X"57",X"43",X"31",X"22",X"1E",X"23",
		X"2E",X"3F",X"53",X"6A",X"80",X"98",X"AD",X"C0",X"CB",X"CA",X"C4",X"B8",X"A8",X"95",X"81",X"6F",
		X"67",X"67",X"6C",X"76",X"83",X"92",X"A1",X"AE",X"B1",X"AD",X"A3",X"95",X"85",X"73",X"61",X"51",
		X"4A",X"4C",X"54",X"61",X"70",X"82",X"95",X"A6",X"B4",X"B7",X"B2",X"A9",X"9A",X"89",X"77",X"64",
		X"52",X"46",X"43",X"49",X"54",X"63",X"74",X"87",X"99",X"A8",X"AC",X"A9",X"A1",X"94",X"84",X"73",
		X"61",X"51",X"49",X"4B",X"53",X"60",X"70",X"82",X"94",X"A6",X"B7",X"C1",X"C1",X"B9",X"AD",X"9C",
		X"89",X"76",X"62",X"4F",X"3C",X"2B",X"1C",X"13",X"15",X"20",X"31",X"45",X"5C",X"75",X"8D",X"A5",
		X"BB",X"D0",X"E2",X"F2",X"FC",X"FD",X"FC",X"F0",X"DD",X"C6",X"AC",X"91",X"77",X"5D",X"46",X"30",
		X"1D",X"0C",X"02",X"03",X"02",X"0C",X"21",X"39",X"53",X"6E",X"88",X"A1",X"B8",X"CD",X"E0",X"EF",
		X"FB",X"FB",X"F3",X"E3",X"D0",X"B8",X"9F",X"85",X"6B",X"54",X"3D",X"28",X"17",X"0E",X"11",X"1C",
		X"2D",X"41",X"58",X"71",X"89",X"A0",X"B6",X"C8",X"D2",X"D1",X"C9",X"BC",X"AA",X"96",X"81",X"72",
		X"6C",X"6D",X"73",X"7D",X"89",X"98",X"A7",X"B4",X"BC",X"B9",X"B1",X"A4",X"93",X"7F",X"6C",X"58",
		X"45",X"3A",X"3A",X"41",X"4D",X"5D",X"6F",X"81",X"92",X"99",X"98",X"93",X"88",X"7B",X"6C",X"5B",
		X"4C",X"46",X"49",X"52",X"5F",X"6F",X"82",X"94",X"A6",X"B1",X"B1",X"AB",X"A0",X"91",X"80",X"6E",
		X"5B",X"4C",X"46",X"49",X"52",X"60",X"71",X"83",X"95",X"A5",X"AB",X"A8",X"A1",X"94",X"85",X"74",
		X"62",X"52",X"41",X"31",X"22",X"19",X"1A",X"24",X"35",X"49",X"60",X"79",X"91",X"A9",X"BF",X"D2",
		X"DF",X"E1",X"DA",X"CD",X"BC",X"A6",X"90",X"7A",X"64",X"4F",X"3C",X"2C",X"24",X"28",X"32",X"42",
		X"56",X"6D",X"84",X"9B",X"B2",X"C6",X"D9",X"E9",X"F8",X"FE",X"FD",X"FE",X"F7",X"E4",X"CC",X"B2",
		X"97",X"7C",X"62",X"4B",X"34",X"21",X"0F",X"04",X"03",X"0B",X"1B",X"2F",X"47",X"61",X"7A",X"93",
		X"AC",X"C2",X"D6",X"E6",X"F4",X"F8",X"F0",X"E2",X"CF",X"B8",X"9F",X"86",X"6D",X"56",X"49",X"46",
		X"4A",X"55",X"63",X"73",X"84",X"95",X"A0",X"A0",X"9C",X"92",X"83",X"73",X"62",X"50",X"3E",X"2E",
		X"20",X"14",X"12",X"1A",X"28",X"3B",X"52",X"69",X"81",X"99",X"AF",X"C3",X"D2",X"D5",X"D0",X"C5",
		X"B6",X"A1",X"8C",X"76",X"60",X"4C",X"39",X"29",X"23",X"27",X"32",X"43",X"57",X"6D",X"85",X"9B",
		X"B2",X"C6",X"D9",X"E8",X"F5",X"FA",X"F3",X"E6",X"D2",X"BD",X"A4",X"8B",X"71",X"5C",X"51",X"4F",
		X"54",X"5E",X"6C",X"7A",X"89",X"8F",X"8E",X"88",X"7D",X"70",X"61",X"52",X"4A",X"4B",X"52",X"5E",
		X"6E",X"7F",X"92",X"A4",X"B4",X"C0",X"C1",X"BA",X"AF",X"9E",X"8B",X"76",X"62",X"4F",X"45",X"44",
		X"4B",X"56",X"65",X"76",X"89",X"9C",X"AC",X"B6",X"B5",X"AE",X"A2",X"92",X"7F",X"6B",X"58",X"46",
		X"34",X"24",X"15",X"09",X"04",X"0A",X"18",X"2B",X"43",X"5D",X"77",X"90",X"A8",X"BF",X"D4",X"E6",
		X"F6",X"FC",X"FC",X"FC",X"F2",X"DD",X"C6",X"AC",X"92",X"78",X"5E",X"47",X"31",X"1E",X"12",X"11",
		X"19",X"27",X"3A",X"51",X"69",X"81",X"99",X"AF",X"C5",X"D6",X"E5",X"EF",X"EC",X"E0",X"D0",X"BC",
		X"A4",X"8D",X"74",X"5D",X"47",X"32",X"1F",X"0F",X"06",X"08",X"14",X"24",X"3A",X"52",X"6C",X"85",
		X"9E",X"B5",X"CA",X"DC",X"ED",X"FA",X"FD",X"FC",X"FD",X"F8",X"E5",X"CD",X"B2",X"96",X"7B",X"60",
		X"48",X"31",X"1C",X"0A",X"02",X"03",X"02",X"08",X"1B",X"32",X"4C",X"66",X"80",X"9A",X"B1",X"C7",
		X"DA",X"EA",X"F6",X"F6",X"ED",X"DE",X"CA",X"B2",X"98",X"7F",X"65",X"4E",X"38",X"24",X"12",X"05",
		X"03",X"03",X"08",X"1B",X"31",X"4A",X"64",X"7F",X"97",X"AF",X"C4",X"D6",X"E2",X"E1",X"D9",X"CB",
		X"B9",X"A3",X"8D",X"76",X"5F",X"4A",X"35",X"26",X"22",X"27",X"33",X"45",X"59",X"6F",X"86",X"9D",
		X"B2",X"C7",X"D9",X"E8",X"F3",X"F6",X"ED",X"DE",X"CA",X"B3",X"99",X"81",X"68",X"50",X"3A",X"26",
		X"14",X"05",X"02",X"03",X"0B",X"1E",X"34",X"4D",X"67",X"81",X"9A",X"B3",X"CA",X"DD",X"EF",X"FC",
		X"FE",X"FD",X"FE",X"F6",X"E2",X"C9",X"AE",X"93",X"78",X"5F",X"4D",X"46",X"47",X"4E",X"5A",X"69",
		X"7B",X"8B",X"98",X"9B",X"97",X"8F",X"82",X"73",X"63",X"52",X"42",X"39",X"39",X"41",X"4E",X"5E",
		X"70",X"82",X"93",X"9C",X"9B",X"96",X"8B",X"7E",X"6E",X"5E",X"4D",X"3D",X"2E",X"20",X"17",X"1A",
		X"24",X"34",X"49",X"60",X"78",X"90",X"A8",X"BE",X"D2",X"E4",X"F4",X"FD",X"FD",X"FD",X"F8",X"E6",
		X"CF",X"B5",X"9A",X"7F",X"65",X"4D",X"36",X"22",X"14",X"11",X"17",X"25",X"37",X"4C",X"64",X"7C",
		X"93",X"A8",X"B8",X"BC",X"B8",X"B0",X"A2",X"91",X"7F",X"6C",X"5C",X"56",X"58",X"60",X"6C",X"7B",
		X"8C",X"9D",X"AE",X"BE",X"CB",X"CE",X"C7",X"BC",X"AC",X"98",X"83",X"6E",X"59",X"4E",X"4B",X"50",
		X"5B",X"69",X"79",X"8C",X"9D",X"AD",X"B7",X"B5",X"AE",X"A2",X"92",X"80",X"6D",X"5A",X"48",X"40",
		X"40",X"47",X"54",X"65",X"77",X"8A",X"9C",X"AC",X"B2",X"AF",X"A7",X"99",X"89",X"77",X"64",X"52",
		X"40",X"2F",X"1F",X"12",X"07",X"05",X"0D",X"1D",X"31",X"49",X"63",X"7E",X"98",X"B0",X"C7",X"DB",
		X"ED",X"FA",X"FD",X"FC",X"FC",X"F3",X"DE",X"C7",X"AC",X"92",X"77",X"5E",X"47",X"32",X"1F",X"10",
		X"0D",X"14",X"21",X"34",X"4A",X"62",X"7B",X"94",X"AC",X"C1",X"D5",X"E5",X"F2",X"F8",X"F2",X"E5",
		X"D1",X"BB",X"A1",X"88",X"6F",X"57",X"41",X"2C",X"1A",X"09",X"02",X"02",X"06",X"18",X"2D",X"46",
		X"61",X"7C",X"96",X"AE",X"C4",X"D8",X"E9",X"F8",X"FE",X"FC",X"FD",X"F2",X"DE",X"C6",X"AB",X"8F",
		X"75",X"5B",X"43",X"2D",X"1A",X"09",X"02",X"02",X"05",X"14",X"29",X"41",X"5B",X"75",X"8F",X"A7",
		X"BE",X"D3",X"E4",X"F4",X"FD",X"FC",X"FB",X"EF",X"DB",X"C3",X"A9",X"8E",X"74",X"5A",X"42",X"2B",
		X"18",X"08",X"02",X"03",X"0E",X"20",X"36",X"4E",X"68",X"82",X"9B",X"B3",X"C8",X"DB",X"E9",X"F6",
		X"F9",X"F1",X"E2",X"CE",X"B8",X"9D",X"84",X"6B",X"53",X"3C",X"27",X"15",X"06",X"01",X"04",X"10",
		X"23",X"39",X"52",X"6C",X"86",X"A0",X"B7",X"CD",X"E0",X"EF",X"FB",X"FD",X"F4",X"E4",X"D0",X"B8",
		X"9E",X"83",X"69",X"51",X"3A",X"26",X"13",X"05",X"02",X"02",X"0A",X"1D",X"33",X"4C",X"65",X"80",
		X"9A",X"B2",X"C8",X"DC",X"ED",X"FA",X"FE",X"FC",X"FC",X"F4",X"DF",X"C7",X"AD",X"91",X"77",X"5D",
		X"45",X"37",X"34",X"38",X"43",X"52",X"64",X"77",X"8A",X"99",X"9F",X"9D",X"95",X"89",X"7A",X"69",
		X"57",X"45",X"35",X"25",X"17",X"0A",X"04",X"08",X"15",X"28",X"3E",X"57",X"71",X"8B",X"A4",X"BB",
		X"D1",X"E3",X"F3",X"FD",X"FD",X"FD",X"FD",X"F0",X"DA",X"C1",X"A5",X"8A",X"6E",X"55",X"3D",X"28",
		X"15",X"08",X"06",X"0F",X"1E",X"32",X"49",X"61",X"7B",X"94",X"AB",X"C1",X"D5",X"E4",X"F1",X"F6",
		X"EF",X"E1",X"CE",X"B7",X"9E",X"85",X"6B",X"53",X"3C",X"28",X"16",X"0A",X"0A",X"13",X"22",X"35",
		X"4C",X"64",X"7D",X"96",X"AE",X"C3",X"D7",X"E6",X"F2",X"F6",X"EF",X"E0",X"CC",X"B6",X"9C",X"83",
		X"6A",X"52",X"40",X"38",X"39",X"42",X"4F",X"60",X"72",X"83",X"91",X"95",X"93",X"8B",X"7E",X"70",
		X"60",X"50",X"46",X"45",X"4C",X"58",X"67",X"79",X"8D",X"A0",X"B1",X"C0",X"C6",X"C2",X"B8",X"AA",
		X"98",X"84",X"70",X"5C",X"4B",X"43",X"45",X"4C",X"59",X"69",X"7B",X"8E",X"9F",X"AD",X"B0",X"AB",
		X"A2",X"93",X"83",X"71",X"5E",X"4C",X"42",X"42",X"48",X"55",X"66",X"77",X"8B",X"9D",X"AD",X"B3",
		X"B1",X"A9",X"9C",X"8B",X"7A",X"67",X"56",X"4E",X"4F",X"57",X"63",X"72",X"84",X"96",X"A8",X"BA",
		X"CA",X"DA",X"E8",X"F5",X"FD",X"FE",X"FE",X"FE",X"FD",X"FD",X"FC",X"FC",X"F8",X"E3",X"C8",X"AA",
		X"8B",X"6D",X"51",X"36",X"1E",X"09",X"03",X"04",X"03",X"03",X"0F",X"25",X"3C",X"56",X"6F",X"88",
		X"9F",X"B4",X"C6",X"D6",X"E4",X"F0",X"F9",X"FE",X"FD",X"FE",X"FE",X"FD",X"EE",X"D5",X"BB",X"9C",
		X"7D",X"60",X"43",X"28",X"10",X"02",X"03",X"02",X"02",X"01",X"01",X"01",X"01",X"01",X"03",X"01",
		X"09",X"28",X"48",X"68",X"86",X"A3",X"BD",X"D3",X"E6",X"F7",X"FE",X"FD",X"FE",X"FD",X"FE",X"FD",
		X"FD",X"FC",X"FD",X"FA",X"E4",X"C6",X"A6",X"86",X"68",X"4A",X"30",X"17",X"05",X"02",X"03",X"02",
		X"02",X"01",X"01",X"00",X"01",X"00",X"06",X"22",X"42",X"62",X"82",X"9F",X"BA",X"D1",X"E6",X"F8",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FD",X"FE",X"F8",X"E0",X"C0",X"A0",X"81",X"63",X"47",
		X"2E",X"16",X"05",X"02",X"02",X"01",X"02",X"01",X"02",X"01",X"03",X"02",X"08",X"23",X"44",X"63",
		X"83",X"A0",X"BC",X"D4",X"EB",X"FB",X"FE",X"FE",X"FE",X"FE",X"FE",X"FD",X"FE",X"FD",X"FD",X"F9",
		X"E0",X"BF",X"A0",X"81",X"65",X"4A",X"31",X"1B",X"08",X"02",X"03",X"03",X"03",X"02",X"02",X"03",
		X"02",X"10",X"2E",X"4C",X"6B",X"89",X"A6",X"C1",X"D9",X"EF",X"FD",X"FD",X"FD",X"FD",X"FE",X"FD",
		X"FD",X"FD",X"FD",X"FC",X"FD",X"ED",X"CE",X"AE",X"8F",X"70",X"54",X"3B",X"24",X"0F",X"03",X"03",
		X"03",X"03",X"03",X"03",X"03",X"03",X"02",X"0F",X"2D",X"4B",X"6B",X"8A",X"A8",X"C3",X"DB",X"F1",
		X"FD",X"FC",X"FD",X"FD",X"FD",X"FC",X"FC",X"FB",X"E7",X"CA",X"AD",X"90",X"73",X"58",X"41",X"2B",
		X"17",X"07",X"02",X"02",X"03",X"02",X"03",X"02",X"08",X"22",X"3E",X"5D",X"7C",X"99",X"B5",X"CF",
		X"E6",X"F9",X"FD",X"FC",X"FC",X"FB",X"FC",X"FB",X"FC",X"FC",X"FD",X"FC",X"FD",X"EE",X"CE",X"AE",
		X"8F",X"71",X"55",X"3B",X"24",X"10",X"03",X"02",X"02",X"02",X"03",X"03",X"04",X"02",X"07",X"21",
		X"40",X"5F",X"7F",X"9C",X"B9",X"D2",X"EA",X"FB",X"FF",X"FE",X"FF",X"FE",X"FE",X"FD",X"FD",X"FD",
		X"FD",X"FC",X"FD",X"F8",X"DC",X"BB",X"9C",X"7D",X"5F",X"44",X"2D",X"17",X"06",X"03",X"02",X"02",
		X"02",X"02",X"02",X"02",X"01",X"05",X"1E",X"3E",X"5E",X"7E",X"9C",X"B8",X"D1",X"E8",X"F9",X"FD",
		X"FC",X"FC",X"FC",X"FC",X"FD",X"F5",X"DB",X"BF",X"A2",X"86",X"6B",X"52",X"3C",X"27",X"15",X"06",
		X"01",X"01",X"01",X"01",X"02",X"02",X"05",X"1B",X"39",X"57",X"76",X"94",X"B1",X"CC",X"E4",X"F9",
		X"FE",X"FD",X"FF",X"FE",X"FF",X"FE",X"FE",X"FE",X"FE",X"FD",X"FD",X"FC",X"FC",X"EB",X"C8",X"A8",
		X"88",X"6A",X"4E",X"36",X"20",X"0C",X"02",X"02",X"01",X"02",X"01",X"02",X"01",X"0F",X"2C",X"49",
		X"68",X"86",X"A2",X"BC",X"D4",X"EA",X"FA",X"FD",X"FD",X"FE",X"FD",X"FF",X"F9",X"E2",X"C6",X"AA",
		X"8E",X"72",X"58",X"40",X"2A",X"18",X"07",X"01",X"01",X"01",X"02",X"02",X"08",X"1E",X"3A",X"57",
		X"76",X"93",X"B0",X"C9",X"E0",X"F5",X"FE",X"FD",X"FD",X"FD",X"FD",X"FC",X"FD",X"F8",X"E0",X"C3",
		X"A5",X"88",X"6E",X"54",X"3D",X"28",X"16",X"07",X"02",X"03",X"03",X"03",X"02",X"02",X"02",X"07",
		X"20",X"3F",X"5E",X"7D",X"9B",X"B9",X"D3",X"EB",X"FB",X"FD",X"FC",X"FD",X"FC",X"FD",X"FC",X"FC",
		X"FC",X"FC",X"FC",X"FD",X"F5",X"D6",X"B5",X"95",X"76",X"5A",X"40",X"2A",X"16",X"06",X"01",X"03",
		X"02",X"03",X"02",X"03",X"02",X"06",X"20",X"3F",X"5E",X"7E",X"9B",X"B7",X"D0",X"E7",X"F9",X"FC",
		X"FC",X"FB",X"FB",X"FC",X"FD",X"F6",X"DE",X"C1",X"A4",X"89",X"6E",X"55",X"3E",X"29",X"18",X"08",
		X"02",X"02",X"02",X"02",X"02",X"02",X"03",X"14",X"31",X"4F",X"6E",X"8D",X"AA",X"C6",X"DF",X"F5",
		X"FE",X"FD",X"FD",X"FC",X"FD",X"FD",X"FD",X"FC",X"FD",X"FC",X"FE",X"FD",X"FD",X"EE",X"CC",X"AC",
		X"8C",X"6D",X"51",X"38",X"22",X"0E",X"02",X"02",X"02",X"02",X"02",X"02",X"01",X"02",X"01",X"11",
		X"31",X"50",X"6F",X"8D",X"AB",X"C6",X"DE",X"F3",X"FD",X"FB",X"FC",X"FD",X"FD",X"FD",X"FC",X"FC",
		X"FC",X"FB",X"FD",X"EE",X"CD",X"AD",X"8E",X"70",X"54",X"3A",X"23",X"0F",X"03",X"02",X"02",X"03",
		X"02",X"03",X"02",X"03",X"02",X"0F",X"2E",X"4D",X"6C",X"8B",X"A9",X"C4",X"DC",X"F2",X"FE",X"FE",
		X"FE",X"FE",X"FE",X"FE",X"FF",X"F5",X"D9",X"BB",X"9E",X"82",X"67",X"4F",X"37",X"24",X"12",X"04",
		X"01",X"02",X"02",X"03",X"02",X"09",X"21",X"3D",X"5B",X"79",X"97",X"B3",X"CC",X"E2",X"F6",X"FE",
		X"FD",X"FF",X"FE",X"FF",X"FE",X"FE",X"FE",X"FE",X"FD",X"FE",X"ED",X"CC",X"AD",X"8E",X"6F",X"53",
		X"3A",X"23",X"0F",X"02",X"02",X"01",X"02",X"02",X"03",X"02",X"03",X"02",X"0D",X"2B",X"49",X"69",
		X"88",X"A6",X"C1",X"D9",X"F0",X"FD",X"FE",X"FD",X"FC",X"FD",X"FD",X"FE",X"FD",X"FD",X"FC",X"FC",
		X"FA",X"E3",X"C1",X"A2",X"83",X"65",X"4A",X"31",X"1B",X"08",X"01",X"01",X"01",X"03",X"02",X"03",
		X"02",X"04",X"03",X"09",X"23",X"41",X"61",X"81",X"9F",X"BB",X"D4",X"EB",X"FB",X"FD",X"FD",X"FD",
		X"FD",X"FC",X"FC",X"FA",X"E5",X"C8",X"AB",X"8E",X"73",X"59",X"43",X"2D",X"1B",X"0B",X"03",X"03",
		X"02",X"03",X"04",X"15",X"2F",X"4A",X"67",X"84",X"A1",X"BB",X"D3",X"E9",X"FA",X"FE",X"FE",X"FD",
		X"FE",X"FD",X"FC",X"FC",X"EC",X"CE",X"B2",X"95",X"7A",X"5F",X"48",X"32",X"20",X"0E",X"03",X"02",
		X"02",X"02",X"01",X"02",X"03",X"16",X"33",X"50",X"6F",X"8D",X"A9",X"C3",X"DC",X"F2",X"FD",X"FC",
		X"FE",X"FE",X"FF",X"FE",X"FE",X"FD",X"FD",X"FC",X"FC",X"EE",X"CE",X"AF",X"90",X"73",X"58",X"3F",
		X"29",X"15",X"05",X"02",X"02",X"01",X"01",X"00",X"01",X"02",X"02",X"14",X"33",X"51",X"71",X"8F",
		X"AC",X"C6",X"DE",X"F4",X"FE",X"FD",X"FE",X"FE",X"FE",X"FE",X"FE",X"FA",X"E3",X"C5",X"A8",X"8B",
		X"6F",X"55",X"3E",X"29",X"17",X"07",X"01",X"03",X"02",X"02",X"01",X"0A",X"23",X"3E",X"5C",X"79",
		X"96",X"B1",X"CB",X"E2",X"F6",X"FD",X"FC",X"FC",X"FD",X"FD",X"FD",X"FA",X"E6",X"CA",X"AE",X"92",
		X"77",X"5C",X"44",X"2F",X"1D",X"0D",X"03",X"02",X"02",X"02",X"02",X"05",X"19",X"34",X"50",X"6E",
		X"8C",X"A8",X"C2",X"D9",X"EF",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FD",X"FD",X"FD",X"FD",X"FE",
		X"F5",X"D7",X"B7",X"98",X"79",X"5C",X"43",X"2C",X"18",X"06",X"02",X"03",X"02",X"02",X"02",X"01",
		X"02",X"01",X"06",X"20",X"3E",X"5D",X"7C",X"9A",X"B6",X"CF",X"E5",X"F8",X"FE",X"FD",X"FE",X"FD",
		X"FD",X"FD",X"FC",X"FC",X"FC",X"FC",X"F5",X"DB",X"BB",X"9D",X"7E",X"61",X"47",X"2F",X"1A",X"07",
		X"01",X"02",X"01",X"02",X"01",X"00",X"00",X"00",X"01",X"14",X"34",X"53",X"73",X"91",X"AD",X"C6",
		X"DD",X"F2",X"FD",X"FD",X"FD",X"FD",X"FE",X"FE",X"FE",X"FE",X"FD",X"FD",X"F9",X"E0",X"BF",X"A0",
		X"81",X"63",X"48",X"31",X"1C",X"08",X"01",X"02",X"02",X"03",X"03",X"03",X"02",X"03",X"17",X"35",
		X"53",X"72",X"8F",X"AB",X"C5",X"DB",X"EF",X"FC",X"FD",X"FC",X"FC",X"FB",X"FC",X"F2",X"D9",X"BF",
		X"A3",X"87",X"6D",X"54",X"3D",X"28",X"16",X"07",X"00",X"02",X"02",X"02",X"02",X"0B",X"23",X"3E",
		X"5B",X"77",X"94",X"AE",X"C7",X"DC",X"F0",X"FC",X"FD",X"FE",X"FE",X"FE",X"FE",X"FD",X"FD",X"FD",
		X"FC",X"E8",X"C9",X"AB",X"8D",X"70",X"54",X"3B",X"25",X"11",X"02",X"01",X"01",X"01",X"02",X"02",
		X"02",X"02",X"02",X"03",X"18",X"36",X"55",X"74",X"92",X"AE",X"C9",X"E0",X"F4",X"FE",X"FD",X"FE",
		X"FD",X"FD",X"FD",X"FD",X"FE",X"FD",X"FE",X"F2",X"D4",X"B5",X"96",X"79",X"5D",X"44",X"2D",X"19",
		X"07",X"01",X"02",X"02",X"03",X"02",X"03",X"01",X"0C",X"28",X"45",X"62",X"7F",X"9B",X"B5",X"CD",
		X"E2",X"F5",X"FD",X"FC",X"FC",X"FC",X"FC",X"FC",X"F1",X"D7",X"BC",X"A0",X"85",X"6B",X"53",X"3D",
		X"29",X"1B",X"18",X"1D",X"2A",X"3C",X"51",X"68",X"80",X"97",X"AE",X"C2",X"D5",X"E5",X"F1",X"F9",
		X"F6",X"EB",X"D9",X"C5",X"AD",X"95",X"7D",X"65",X"4F",X"3A",X"27",X"16",X"08",X"02",X"05",X"0F",
		X"20",X"36",X"4F",X"68",X"81",X"99",X"B1",X"C6",X"D9",X"EA",X"F8",X"FD",X"FC",X"FC",X"F7",X"E4",
		X"CE",X"B4",X"9A",X"80",X"67",X"50",X"3A",X"26",X"15",X"06",X"01",X"02",X"02",X"02",X"01",X"02",
		X"01",X"10",X"2B",X"47",X"65",X"82",X"9E",X"B8",X"D1",X"E5",X"F8",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"FD",X"FB",X"E7",X"CB",X"B0",X"93",X"78",X"5F",X"47",X"32",X"20",X"10",X"04",X"01",X"02",X"02",
		X"02",X"02",X"0D",X"27",X"41",X"5E",X"7A",X"95",X"AE",X"C7",X"DC",X"F0",X"FC",X"FD",X"FD",X"FD",
		X"FE",X"FD",X"FE",X"F6",X"DD",X"C2",X"A5",X"8A",X"70",X"58",X"42",X"2D",X"1B",X"0C",X"02",X"02",
		X"02",X"02",X"0A",X"1F",X"37",X"52",X"6E",X"88",X"A2",X"BA",X"D0",X"E3",X"F4",X"FD",X"FD",X"FD",
		X"FC",X"FD",X"F4",X"DC",X"C3",X"A8",X"8F",X"74",X"5D",X"46",X"32",X"20",X"14",X"11",X"18",X"25",
		X"37",X"4D",X"64",X"7C",X"93",X"A9",X"BD",X"D0",X"DF",X"EC",X"ED",X"E5",X"D7",X"C6",X"B1",X"9A",
		X"84",X"6D",X"57",X"43",X"31",X"21",X"1A",X"1D",X"28",X"37",X"4B",X"61",X"77",X"8E",X"A3",X"B8",
		X"CB",X"DC",X"E9",X"F4",X"FB",X"F6",X"EA",X"D9",X"C4",X"AC",X"94",X"7B",X"64",X"4E",X"3B",X"29",
		X"19",X"0C",X"04",X"04",X"04",X"04",X"03",X"08",X"1D",X"35",X"4F",X"6A",X"85",X"9F",X"B7",X"CE",
		X"E0",X"F2",X"FC",X"FC",X"FD",X"FD",X"FD",X"F1",X"DA",X"C2",X"A8",X"8F",X"75",X"5E",X"48",X"34",
		X"24",X"1B",X"1D",X"26",X"35",X"48",X"5D",X"73",X"89",X"9E",X"B3",X"C5",X"D7",X"E4",X"EF",X"F3",
		X"EC",X"DD",X"CC",X"B7",X"A0",X"89",X"71",X"5C",X"47",X"34",X"23",X"15",X"09",X"02",X"02",X"02",
		X"03",X"03",X"02",X"09",X"1E",X"37",X"52",X"6D",X"88",X"A2",X"B9",X"D0",X"E2",X"F4",X"FD",X"FD",
		X"FE",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"F8",X"E3",X"C6",X"AA",X"8D",X"72",X"59",X"42",X"2D",
		X"1C",X"0C",X"02",X"02",X"01",X"02",X"02",X"03",X"03",X"07",X"1B",X"35",X"50",X"6B",X"86",X"A0",
		X"B7",X"CD",X"DF",X"EF",X"FA",X"FD",X"FD",X"FE",X"FD",X"FE",X"FD",X"FE",X"F9",X"E3",X"C9",X"AC",
		X"91",X"77",X"5E",X"47",X"32",X"1F",X"0F",X"03",X"01",X"01",X"08",X"19",X"2D",X"45",X"5C",X"75",
		X"8C",X"A2",X"B6",X"C8",X"D7",X"E2",X"E5",X"DF",X"D2",X"C2",X"AE",X"98",X"83",X"6D",X"59",X"46",
		X"35",X"25",X"18",X"0D",X"09",X"0F",X"1B",X"2D",X"41",X"57",X"6E",X"84",X"9B",X"B0",X"C3",X"D4",
		X"E3",X"EE",X"F8",X"FC",X"F6",X"EA",X"D7",X"C3",X"AC",X"94",X"7C",X"65",X"50",X"3D",X"2D",X"1E",
		X"12",X"0D",X"11",X"1C",X"2C",X"40",X"55",X"6B",X"82",X"97",X"AA",X"BA",X"BF",X"BC",X"B5",X"AA",
		X"9A",X"8A",X"79",X"68",X"57",X"48",X"3A",X"31",X"30",X"36",X"42",X"53",X"65",X"78",X"8C",X"A0",
		X"B3",X"C4",X"D3",X"E1",X"EB",X"F3",X"F6",X"F0",X"E3",X"D1",X"BD",X"A6",X"90",X"79",X"63",X"4F",
		X"3E",X"2D",X"20",X"14",X"0A",X"03",X"01",X"01",X"01",X"02",X"0C",X"1F",X"35",X"4E",X"67",X"80",
		X"98",X"AE",X"C3",X"D5",X"E5",X"F2",X"FC",X"FD",X"FD",X"FD",X"FE",X"F8",X"E4",X"CF",X"B7",X"9E",
		X"86",X"6F",X"5A",X"47",X"36",X"27",X"1E",X"1F",X"27",X"34",X"45",X"58",X"6D",X"81",X"95",X"A8",
		X"BA",X"C9",X"D7",X"E2",X"EA",X"EC",X"E4",X"D7",X"C6",X"B3",X"9D",X"88",X"73",X"5F",X"4D",X"3C",
		X"2E",X"22",X"1E",X"22",X"2C",X"3A",X"4C",X"5E",X"72",X"85",X"99",X"AB",X"BB",X"CA",X"D6",X"DF",
		X"DF",X"D7",X"CA",X"BA",X"A7",X"93",X"7F",X"6C",X"59",X"48",X"38",X"2B",X"21",X"1F",X"25",X"31",
		X"40",X"52",X"65",X"79",X"8C",X"9E",X"AF",X"BF",X"CD",X"D8",X"DF",X"DD",X"D4",X"C6",X"B5",X"A2",
		X"8E",X"7A",X"67",X"55",X"45",X"36",X"29",X"1E",X"19",X"1D",X"27",X"35",X"47",X"5A",X"6E",X"81",
		X"95",X"A6",X"B5",X"BE",X"BF",X"BA",X"B0",X"A3",X"94",X"85",X"74",X"65",X"56",X"48",X"3F",X"3D",
		X"41",X"4A",X"57",X"67",X"77",X"88",X"99",X"A9",X"B7",X"C5",X"D1",X"DA",X"DF",X"DB",X"D1",X"C3",
		X"B2",X"9F",X"8C",X"79",X"67",X"56",X"46",X"39",X"2D",X"23",X"1F",X"22",X"2C",X"39",X"4A",X"5C",
		X"6F",X"82",X"94",X"A6",X"B6",X"C4",X"D0",X"DA",X"E1",X"E0",X"D8",X"CB",X"BB",X"A8",X"94",X"81",
		X"6E",X"5D",X"4D",X"3F",X"32",X"29",X"28",X"2E",X"38",X"46",X"56",X"68",X"79",X"8A",X"9B",X"AB",
		X"B9",X"C4",X"CD",X"CE",X"C8",X"BE",X"B0",X"A0",X"8F",X"7E",X"6D",X"5D",X"4E",X"41",X"35",X"2B",
		X"29",X"2D",X"36",X"44",X"53",X"65",X"76",X"88",X"98",X"A8",X"B7",X"C4",X"CE",X"D6",X"D7",X"D0",
		X"C4",X"B6",X"A6",X"94",X"82",X"71",X"61",X"51",X"44",X"38",X"2F",X"2E",X"34",X"3E",X"4B",X"5A",
		X"6A",X"7B",X"8C",X"9B",X"AA",X"B7",X"C3",X"CC",X"D3",X"D2",X"CB",X"C0",X"B2",X"A1",X"90",X"7F",
		X"6E",X"5E",X"50",X"43",X"37",X"2D",X"24",X"1E",X"18",X"14",X"13",X"18",X"23",X"32",X"43",X"56",
		X"69",X"7C",X"8F",X"A1",X"B1",X"BF",X"CC",X"D6",X"DE",X"E6",X"EC",X"EF",X"F1",X"F1",X"EB",X"DE",
		X"CD",X"BB",X"A7",X"93",X"7F",X"6C",X"5B",X"4C",X"3E",X"32",X"28",X"23",X"25",X"2C",X"38",X"46",
		X"56",X"66",X"77",X"88",X"97",X"A5",X"B2",X"BC",X"C3",X"C1",X"BB",X"B1",X"A4",X"96",X"86",X"77",
		X"68",X"5A",X"4D",X"42",X"38",X"30",X"29",X"23",X"1F",X"1C",X"1E",X"26",X"33",X"42",X"54",X"66",
		X"78",X"89",X"9A",X"A9",X"B6",X"C3",X"CD",X"D5",X"DA",X"D9",X"D1",X"C6",X"B8",X"A9",X"98",X"88",
		X"78",X"69",X"5B",X"4F",X"45",X"41",X"43",X"49",X"53",X"5F",X"6D",X"7A",X"88",X"96",X"A2",X"AE",
		X"B8",X"C1",X"C7",X"CA",X"C5",X"BD",X"B1",X"A4",X"94",X"85",X"75",X"67",X"5A",X"4E",X"43",X"3A",
		X"36",X"38",X"3F",X"49",X"56",X"63",X"72",X"80",X"8E",X"9B",X"A6",X"B2",X"BA",X"C2",X"C5",X"C1",
		X"BA",X"AF",X"A2",X"94",X"85",X"77",X"69",X"5C",X"50",X"46",X"3D",X"36",X"34",X"38",X"3F",X"4A",
		X"57",X"65",X"73",X"81",X"8F",X"9C",X"A8",X"B2",X"BB",X"C2",X"C6",X"C4",X"BC",X"B2",X"A6",X"98",
		X"89",X"7B",X"6D",X"61",X"55",X"4B",X"42",X"3C",X"3D",X"42",X"4B",X"56",X"62",X"70",X"7D",X"8A",
		X"96",X"A1",X"AC",X"B4",X"BA",X"BC",X"B8",X"B0",X"A6",X"9B",X"8D",X"80",X"73",X"67",X"5C",X"51",
		X"48",X"41",X"3E",X"41",X"48",X"52",X"5D",X"6A",X"77",X"83",X"8F",X"9B",X"A5",X"AE",X"B5",X"BB",
		X"BD",X"BA",X"B2",X"A8",X"9D",X"90",X"83",X"76",X"6A",X"5E",X"54",X"4B",X"43",X"3D",X"3C",X"41",
		X"48",X"52",X"5E",X"6A",X"77",X"83",X"8F",X"99",X"A2",X"A5",X"A3",X"9E",X"97",X"8E",X"85",X"7B",
		X"71",X"67",X"5E",X"56",X"4F",X"4D",X"4F",X"55",X"5D",X"67",X"72",X"7D",X"88",X"93",X"9D",X"A5",
		X"AE",X"B4",X"BA",X"BB",X"B6",X"AF",X"A6",X"9B",X"8F",X"83",X"77",X"6C",X"61",X"58",X"4F",X"48",
		X"45",X"46",X"4C",X"54",X"5E",X"69",X"74",X"80",X"8B",X"95",X"9F",X"A7",X"AF",X"B4",X"B9",X"B8",
		X"B3",X"AB",X"A1",X"96",X"8A",X"7E",X"73",X"68",X"5E",X"56",X"4E",X"47",X"44",X"46",X"4B",X"53",
		X"5C",X"67",X"72",X"7E",X"88",X"93",X"9C",X"A4",X"AB",X"B1",X"B4",X"B2",X"AD",X"A5",X"9C",X"91",
		X"86",X"7B",X"70",X"66",X"5D",X"55",X"4E",X"48",X"45",X"46",X"4B",X"53",X"5D",X"67",X"72",X"7D",
		X"88",X"92",X"9B",X"A3",X"AA",X"B0",X"B4",X"B7",X"B5",X"AF",X"A7",X"9E",X"93",X"87",X"7C",X"72",
		X"68",X"5F",X"57",X"50",X"4A",X"45",X"43",X"45",X"4B",X"52",X"5C",X"66",X"71",X"7C",X"86",X"90",
		X"99",X"A0",X"A7",X"AD",X"B1",X"B3",X"B0",X"AB",X"A3",X"9A",X"8F",X"85",X"7A",X"71",X"67",X"5F",
		X"58",X"51",X"4E",X"4F",X"53",X"5A",X"62",X"6B",X"74",X"7E",X"87",X"8F",X"97",X"9E",X"A4",X"A9",
		X"AC",X"AC",X"A8",X"A2",X"9A",X"91",X"87",X"7D",X"74",X"6B",X"63",X"5C",X"55",X"51",X"50",X"54",
		X"59",X"60",X"69",X"71",X"7A",X"82",X"8A",X"8F",X"90",X"8E",X"8B",X"86",X"80",X"7A",X"73",X"6D",
		X"67",X"61",X"5E",X"5F",X"62",X"67",X"6E",X"75",X"7C",X"84",X"8B",X"92",X"98",X"9E",X"A2",X"A6",
		X"A7",X"A4",X"9E",X"98",X"90",X"87",X"7F",X"77",X"6F",X"68",X"61",X"5B",X"59",X"5A",X"5E",X"63",
		X"6A",X"71",X"79",X"80",X"87",X"8E",X"92",X"92",X"90",X"8D",X"88",X"82",X"7C",X"76",X"70",X"6A",
		X"64",X"5F",X"5C",X"5C",X"5F",X"64",X"6A",X"71",X"79",X"80",X"88",X"8F",X"95",X"9B",X"9F",X"A4",
		X"A7",X"A9",X"A8",X"A4",X"9F",X"98",X"90",X"87",X"7F",X"77",X"6F",X"68",X"62",X"5C",X"58",X"54",
		X"54",X"56",X"5B",X"62",X"69",X"71",X"79",X"81",X"88",X"8F",X"95",X"9A",X"9E",X"A1",X"A1",X"9E",
		X"99",X"93",X"8C",X"85",X"7D",X"76",X"6F",X"69",X"63",X"5F",X"5C",X"5C",X"5F",X"64",X"6A",X"70",
		X"77",X"7E",X"85",X"8B",X"91",X"96",X"9A",X"9D",X"A0",X"9F",X"9C",X"97",X"92",X"8B",X"84",X"7C",
		X"75",X"6F",X"69",X"63",X"5F",X"5B",X"58",X"59",X"5B",X"60",X"66",X"6D",X"74",X"7B",X"82",X"88",
		X"8E",X"93",X"98",X"9C",X"9F",X"A0",X"9F",X"9B",X"96",X"90",X"89",X"82",X"7B",X"74",X"6E",X"68",
		X"63",X"5F",X"5D",X"5E",X"61",X"65",X"6B",X"71",X"77",X"7E",X"83",X"89",X"8C",X"8D",X"8C",X"89",
		X"86",X"81",X"7D",X"78",X"73",X"6F",X"6A",X"66",X"63",X"62",X"64",X"67",X"6B",X"71",X"77",X"7C",
		X"82",X"88",X"8D",X"92",X"96",X"99",X"9B",X"9D",X"9C",X"99",X"94",X"8F",X"89",X"83",X"7D",X"77",
		X"71",X"6C",X"68",X"64",X"61",X"61",X"63",X"67",X"6C",X"71",X"77",X"7C",X"82",X"87",X"8C",X"91",
		X"94",X"97",X"9A",X"9B",X"99",X"96",X"92",X"8D",X"87",X"81",X"7B",X"76",X"70",X"6B",X"67",X"63",
		X"60",X"5E",X"5F",X"62",X"66",X"6C",X"71",X"77",X"7D",X"82",X"88",X"8C",X"90",X"94",X"97",X"98",
		X"98",X"96",X"92",X"8E",X"89",X"84",X"7E",X"79",X"74",X"70",X"6B",X"68",X"64",X"62",X"61",X"62",
		X"65",X"69",X"6E",X"74",X"79",X"7E",X"83",X"88",X"8C",X"90",X"93",X"96",X"98",X"98",X"95",X"92",
		X"8E",X"89",X"84",X"7F",X"7A",X"75",X"71",X"6D",X"69",X"66",X"66",X"67",X"6A",X"6D",X"72",X"76",
		X"7B",X"80",X"84",X"88",X"8C",X"8F",X"92",X"94",X"95",X"95",X"92",X"8F",X"8B",X"87",X"82",X"7D",
		X"79",X"74",X"70",X"6C",X"69",X"66",X"65",X"66",X"69",X"6C",X"70",X"75",X"79",X"7E",X"82",X"86",
		X"8A",X"8D",X"8F",X"91",X"93",X"92",X"8F",X"8C",X"89",X"84",X"80",X"7B",X"77",X"73",X"70",X"6C",
		X"6A",X"67",X"66",X"67",X"69",X"6D",X"70",X"75",X"79",X"7D",X"82",X"86",X"89",X"8C",X"8E",X"90",
		X"91",X"90",X"8D",X"8A",X"87",X"83",X"7F",X"7B",X"77",X"73",X"70",X"6D",X"6B",X"6B",X"6C",X"6E",
		X"71",X"75",X"78",X"7C",X"80",X"84",X"87",X"8A",X"8C",X"8E",X"8F",X"8E",X"8C",X"89",X"86",X"82",
		X"7F",X"7B",X"77",X"74",X"71",X"6E",X"6D",X"6E",X"70",X"72",X"75",X"78",X"7C",X"7F",X"82",X"84",
		X"84",X"84",X"82",X"80",X"7E",X"7B",X"79",X"76",X"74",X"72",X"70",X"6E",X"6D",X"6D",X"6F",X"72",
		X"75",X"78",X"7C",X"80",X"83",X"86",X"89",X"8C",X"8E",X"90",X"91",X"92",X"91",X"8F",X"8D",X"89",
		X"86",X"82",X"7E",X"7B",X"78",X"74",X"72",X"6F",X"6E",X"6E",X"6F",X"71",X"74",X"77",X"7A",X"7E",
		X"81",X"84",X"86",X"89",X"8B",X"8D",X"8D",X"8D",X"8B",X"89",X"86",X"83",X"80",X"7D",X"7A",X"77",
		X"74",X"71",X"6F",X"6D",X"6D",X"6E",X"70",X"72",X"75",X"78",X"7C",X"7F",X"82",X"85",X"87",X"89",
		X"8B",X"8C",X"8C",X"8B",X"89",X"87",X"84",X"81",X"7E",X"7B",X"78",X"76",X"73",X"71",X"70",X"70",
		X"71",X"73",X"75",X"78",X"7B",X"7E",X"80",X"83",X"85",X"87",X"89",X"8A",X"8B",X"8A",X"89",X"87",
		X"85",X"82",X"7F",X"7D",X"7A",X"77",X"75",X"72",X"71",X"6F",X"6E",X"6F",X"71",X"73",X"76",X"79",
		X"7C",X"7E",X"81",X"84",X"86",X"88",X"8A",X"8B",X"8B",X"8B",X"89",X"87",X"85",X"82",X"80",X"7D",
		X"7A",X"78",X"75",X"73",X"72",X"71",X"71",X"72",X"74",X"76",X"79",X"7B",X"7E",X"80",X"83",X"84",
		X"85",X"84",X"83",X"82",X"80",X"7E",X"7C",X"7A",X"78",X"77",X"75",X"74",X"75",X"76",X"78",X"79",
		X"7C",X"7E",X"80",X"82",X"84",X"85",X"87",X"88",X"89",X"89",X"89",X"88",X"86",X"84",X"82",X"7F",
		X"7D",X"7B",X"78",X"76",X"75",X"73",X"72",X"72",X"73",X"74",X"76",X"78",X"7B",X"7D",X"7F",X"81",
		X"83",X"85",X"86",X"87",X"88",X"88",X"87",X"86",X"84",X"82",X"80",X"7E",X"7C",X"7A",X"78",X"76",
		X"75",X"74",X"73",X"74",X"75",X"77",X"79",X"7B",X"7D",X"7F",X"81",X"83",X"84",X"85",X"86",X"87",
		X"86",X"85",X"83",X"81",X"7F",X"7D",X"7B",X"79",X"78",X"76",X"75",X"74",X"73",X"73",X"74",X"75",
		X"77",X"79",X"7B",X"7D",X"7F",X"81",X"82",X"84",X"85",X"86",X"87",X"86",X"86",X"84",X"83",X"81",
		X"7F",X"7D",X"7B",X"79",X"78",X"76",X"75",X"75",X"75",X"76",X"77",X"79",X"7B",X"7D",X"7E",X"80",
		X"82",X"83",X"84",X"85",X"86",X"86",X"85",X"84",X"83",X"81",X"7F",X"7E",X"7C",X"7A",X"78",X"77",
		X"76",X"75",X"74",X"74",X"74",X"75",X"77",X"79",X"7B",X"7C",X"7E",X"80",X"82",X"83",X"84",X"85",
		X"86",X"86",X"85",X"84",X"83",X"81",X"80",X"7E",X"7C",X"7B",X"79",X"78",X"77",X"76",X"76",X"76",
		X"77",X"79",X"7A",X"7C",X"7E",X"7F",X"81",X"82",X"83",X"84",X"85",X"84",X"84",X"83",X"82",X"80",
		X"7F",X"7D",X"7C",X"7A",X"79",X"78",X"77",X"76",X"76",X"77",X"78",X"79",X"7A",X"7C",X"7E",X"7F",
		X"80",X"82",X"83",X"84",X"84",X"85",X"85",X"85",X"84",X"83",X"82",X"80",X"7F",X"7D",X"7C",X"7A",
		X"79",X"78",X"77",X"77",X"77",X"78",X"79",X"7A",X"7B",X"7D",X"7E",X"80",X"81",X"82",X"83",X"84",
		X"84",X"84",X"84",X"83",X"82",X"81",X"7F",X"7E",X"7D",X"7B",X"7A",X"79",X"78",X"77",X"77",X"77",
		X"78",X"79",X"7A",X"7C",X"7D",X"7E",X"7F",X"81",X"82",X"82",X"83",X"84",X"84",X"83",X"82",X"82",
		X"80",X"7F",X"7E",X"7D",X"7B",X"7A",X"79",X"78",X"77",X"77",X"77",X"78",X"79",X"7A",X"7B",X"7C",
		X"7D",X"7F",X"80",X"81",X"82",X"82",X"83",X"83",X"82",X"82",X"81",X"80",X"7E",X"7D",X"7C",X"7B",
		X"7A",X"79",X"78",X"78",X"78",X"78",X"79",X"7A",X"7B",X"7D",X"7E",X"7F",X"80",X"81",X"82",X"82",
		X"83",X"83",X"83",X"82",X"81",X"80",X"7F",X"7E",X"7D",X"7C",X"7B",X"7A",X"79",X"78",X"78",X"78",
		X"78",X"79",X"7A",X"7B",X"7C",X"7D",X"7E",X"7F",X"80",X"81",X"82",X"82",X"83",X"83",X"82",X"82",
		X"81",X"80",X"7F",X"7E",X"7D",X"7C",X"7B",X"7A",X"79",X"78",X"78",X"79",X"79",X"7A",X"7B",X"7C",
		X"7D",X"7E",X"7F",X"80",X"80",X"80",X"80",X"7F",X"7E",X"7E",X"7D",X"7C",X"7B",X"7B",X"7A",X"79",
		X"79",X"79",X"7A",X"7A",X"7B",X"7C",X"7D",X"7E",X"7F",X"80",X"80",X"81",X"82",X"82",X"82",X"83",
		X"82",X"82",X"81",X"80",X"7F",X"7E",X"7D",X"7C",X"7B",X"7B",X"7A",X"79",X"79",X"79",X"79",X"7A",
		X"7B",X"7C",X"7D",X"7E",X"7E",X"7F",X"80",X"81",X"81",X"81",X"80",X"80",X"7F",X"7E",X"7E",X"7D",
		X"7C",X"7C",X"7B",X"7B",X"7B",X"7B",X"7C",X"7C",X"7D",X"7E",X"7E",X"7F",X"80",X"80",X"80",X"80",
		X"7F",X"7F",X"7E",X"7E",X"7D",X"7C",X"7C",X"7B",X"7B",X"7B",X"7B",X"7B",X"7C",X"7C",X"7D",X"7E",
		X"7E",X"7F",X"80",X"80",X"81",X"81",X"80",X"80",X"7F",X"7E",X"7E",X"7D",X"7C",X"7C",X"7B",X"7A",
		X"7A",X"7A",X"7A",X"7A",X"7B",X"7C",X"7C",X"7D",X"7E",X"7F",X"7F",X"80",X"80",X"81",X"81",X"81",
		X"81",X"81",X"80",X"80",X"7F",X"7E",X"7E",X"7D",X"7C",X"7B",X"7B",X"7A",X"7A",X"7A",X"7A",X"7B",
		X"7C",X"7C",X"7D",X"7E",X"7E",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7E",X"7D",X"7D",X"7C",X"7C",
		X"7B",X"7B",X"7B",X"7B",X"7C",X"7C",X"7D",X"7D",X"7E",X"7E",X"7F",X"7F",X"80",X"80",X"81",X"81",
		X"81",X"81",X"80",X"80",X"7F",X"7E",X"7E",X"7D",X"7C",X"7C",X"7B",X"7B",X"7A",X"7A",X"7A",X"7A",
		X"7B",X"7C",X"7C",X"7D",X"7D",X"7E",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",
		X"7E",X"7E",X"7D",X"7D",X"7C",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7C",X"7C",X"7D",X"7D",X"7E",
		X"7F",X"7F",X"7F",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7E",X"7E",X"7D",X"7D",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7D",X"7D",X"7D",X"7E",X"7E",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"7F",X"7F",X"7E",X"7D",X"7D",X"7C",X"7C",X"7C",X"7B",X"7B",X"7B",X"7B",X"7B",X"7C",X"7C",
		X"7D",X"7D",X"7E",X"7E",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"7F",X"7F",X"7E",X"7E",X"7E",X"7D",
		X"7D",X"7C",X"7C",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7C",X"7C",X"7D",X"7D",X"7E",X"7E",X"7F",
		X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7E",X"7E",X"7D",X"7D",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7D",X"7D",X"7E",X"7E",X"7E",X"7F",X"7F",X"7E",X"7E",X"7E",X"7E",
		X"7D",X"7D",X"7D",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7D",X"7D",X"7D",X"7E",X"7E",X"7E",
		X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7E",X"7E",X"7D",X"7D",X"7C",X"7C",
		X"7C",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7C",X"7C",X"7D",X"7D",X"7E",X"7E",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7E",X"7E",X"7E",X"7D",X"7D",X"7D",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7D",X"7D",X"7D",X"7E",X"7E",X"7E",X"7F",X"7F",X"7F",X"7F",X"7F",X"7E",X"7E",X"7E",X"7D",
		X"7D",X"7D",X"7D",X"7C",X"7C",X"7C",X"7D",X"7D",X"7D",X"7D",X"7E",X"7E",X"7E",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7E",X"7E",X"7E",X"7E",X"7D",X"7D",X"7D",X"7C",X"7C",X"7C",X"7C",X"7D",X"7D",X"7D",
		X"7D",X"7E",X"7E",X"7E",X"7E",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7E",X"7E",X"7E",X"7D",
		X"7D",X"7D",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7D",X"7D",X"7D",X"7E",X"7E",
		X"7E",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7E",X"7E",X"7E",X"7D",X"7D",X"7D",X"7D",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7D",X"7D",X"7D",X"7E",X"7E",X"7E",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7E",X"7E",X"7E",X"7D",X"7D",X"7D",X"7D",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7D",X"7D",X"7D",X"7D",X"7E",X"7E",X"7E",X"7E",X"7E",X"7F",X"7F",X"7F",X"7F",X"7E",
		X"7E",X"7E",X"7E",X"7D",X"7D",X"7D",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7D",X"7D",X"7D",
		X"7D",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",
		X"7D",X"7D",X"7D",X"7D",X"7E",X"7E",X"7E",X"7E",X"7E",X"7F",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7E",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
