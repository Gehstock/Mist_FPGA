library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity tapper_bg_bits_1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of tapper_bg_bits_1 is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"03",X"BB",X"0B",X"FF",X"2B",X"FF",X"2B",X"FF",X"0B",X"FF",X"03",X"FF",X"00",X"FC",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",
		X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",
		X"55",X"00",X"54",X"00",X"54",X"00",X"50",X"00",X"50",X"00",X"40",X"00",X"40",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"5A",X"AA",X"5A",X"AA",X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"00",
		X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"00",X"70",X"00",X"AA",X"AA",X"5A",X"AA",X"50",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"00",X"00",
		X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"AA",X"3C",X"2A",X"3F",X"02",X"3F",X"F0",X"3F",X"FC",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"50",X"55",X"00",X"54",X"00",X"52",X"80",X"50",X"20",
		X"54",X"00",X"50",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"15",X"55",X"05",X"55",X"05",X"55",X"01",X"55",X"01",X"55",X"00",X"55",X"00",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"08",X"40",X"08",X"40",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"03",X"3C",X"0F",X"3F",X"3F",X"3F",X"FF",
		X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"15",
		X"40",X"20",X"52",X"80",X"54",X"00",X"55",X"00",X"55",X"50",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",
		X"55",X"56",X"55",X"56",X"55",X"56",X"55",X"56",X"55",X"56",X"55",X"56",X"55",X"56",X"55",X"56",
		X"55",X"56",X"55",X"56",X"55",X"56",X"55",X"56",X"55",X"56",X"55",X"56",X"55",X"55",X"55",X"55",
		X"55",X"56",X"55",X"56",X"55",X"5A",X"55",X"5B",X"55",X"5B",X"55",X"6B",X"55",X"6B",X"55",X"6B",
		X"55",X"AB",X"55",X"AB",X"55",X"AB",X"56",X"AB",X"56",X"AB",X"56",X"AB",X"5A",X"AB",X"5A",X"AB",
		X"5A",X"AB",X"6A",X"AB",X"6A",X"AB",X"6A",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",
		X"02",X"A8",X"30",X"A8",X"3C",X"20",X"3F",X"00",X"3F",X"C0",X"3F",X"FC",X"3F",X"FF",X"3F",X"FF",
		X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",
		X"3F",X"FF",X"3F",X"FF",X"00",X"00",X"A9",X"50",X"A9",X"70",X"A5",X"AA",X"A5",X"50",X"A5",X"50",
		X"95",X"55",X"95",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"56",X"55",X"56",X"55",X"56",X"55",X"56",X"95",X"56",X"95",X"56",X"95",X"56",X"95",X"56",
		X"05",X"50",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"05",X"50",X"00",X"00",
		X"05",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"05",X"50",X"00",X"00",
		X"05",X"50",X"14",X"54",X"00",X"14",X"00",X"50",X"01",X"40",X"05",X"00",X"15",X"54",X"00",X"00",
		X"05",X"50",X"14",X"14",X"00",X"14",X"01",X"50",X"00",X"14",X"14",X"14",X"05",X"50",X"00",X"00",
		X"01",X"14",X"05",X"14",X"04",X"14",X"14",X"14",X"15",X"54",X"00",X"14",X"00",X"14",X"00",X"00",
		X"15",X"54",X"14",X"00",X"15",X"50",X"00",X"14",X"00",X"14",X"15",X"54",X"15",X"50",X"00",X"00",
		X"01",X"50",X"05",X"04",X"14",X"00",X"15",X"50",X"14",X"14",X"14",X"14",X"05",X"50",X"00",X"00",
		X"15",X"54",X"10",X"14",X"00",X"50",X"01",X"40",X"05",X"40",X"05",X"00",X"05",X"00",X"00",X"00",
		X"05",X"50",X"14",X"14",X"14",X"14",X"05",X"50",X"14",X"14",X"14",X"14",X"05",X"50",X"00",X"00",
		X"05",X"50",X"14",X"14",X"14",X"14",X"05",X"54",X"00",X"14",X"00",X"14",X"00",X"14",X"00",X"00",
		X"15",X"50",X"40",X"04",X"45",X"44",X"44",X"04",X"45",X"44",X"40",X"04",X"15",X"50",X"00",X"00",
		X"FF",X"FF",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"05",X"50",X"14",X"14",X"14",X"14",X"15",X"54",X"14",X"14",X"14",X"14",X"14",X"14",X"00",X"00",
		X"15",X"50",X"14",X"14",X"14",X"14",X"15",X"50",X"14",X"14",X"14",X"14",X"15",X"50",X"00",X"00",
		X"05",X"50",X"14",X"14",X"14",X"00",X"14",X"00",X"14",X"00",X"14",X"04",X"05",X"50",X"00",X"00",
		X"15",X"50",X"14",X"14",X"14",X"04",X"14",X"04",X"14",X"04",X"14",X"14",X"15",X"50",X"00",X"00",
		X"15",X"54",X"14",X"00",X"14",X"00",X"15",X"40",X"14",X"00",X"14",X"00",X"15",X"54",X"00",X"00",
		X"15",X"54",X"14",X"00",X"14",X"00",X"15",X"40",X"14",X"00",X"14",X"00",X"14",X"00",X"00",X"00",
		X"05",X"54",X"14",X"00",X"14",X"00",X"14",X"54",X"14",X"04",X"15",X"54",X"05",X"44",X"00",X"00",
		X"14",X"14",X"14",X"14",X"14",X"14",X"15",X"54",X"14",X"14",X"14",X"14",X"14",X"14",X"00",X"00",
		X"05",X"50",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"05",X"50",X"00",X"00",
		X"05",X"54",X"00",X"50",X"00",X"50",X"00",X"50",X"14",X"50",X"15",X"50",X"05",X"40",X"00",X"00",
		X"14",X"04",X"14",X"14",X"14",X"50",X"15",X"50",X"14",X"14",X"14",X"04",X"14",X"04",X"00",X"00",
		X"14",X"00",X"14",X"00",X"14",X"00",X"14",X"00",X"14",X"00",X"14",X"04",X"15",X"54",X"00",X"00",
		X"14",X"14",X"14",X"14",X"11",X"44",X"11",X"44",X"10",X"04",X"10",X"04",X"10",X"04",X"00",X"00",
		X"14",X"04",X"15",X"04",X"15",X"04",X"11",X"44",X"10",X"44",X"10",X"54",X"10",X"14",X"00",X"00",
		X"05",X"50",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"05",X"50",X"00",X"00",
		X"15",X"50",X"14",X"14",X"14",X"04",X"15",X"54",X"14",X"00",X"14",X"00",X"14",X"00",X"00",X"00",
		X"05",X"50",X"14",X"14",X"10",X"04",X"10",X"04",X"10",X"44",X"14",X"50",X"05",X"54",X"00",X"00",
		X"15",X"50",X"14",X"14",X"14",X"04",X"15",X"54",X"14",X"10",X"14",X"14",X"14",X"04",X"00",X"00",
		X"05",X"54",X"14",X"04",X"14",X"00",X"15",X"54",X"00",X"14",X"10",X"14",X"15",X"50",X"00",X"00",
		X"15",X"54",X"15",X"54",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"00",X"00",
		X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"05",X"50",X"00",X"00",
		X"10",X"04",X"10",X"04",X"14",X"14",X"04",X"10",X"05",X"50",X"01",X"40",X"01",X"40",X"00",X"00",
		X"10",X"04",X"10",X"04",X"10",X"04",X"11",X"44",X"11",X"44",X"15",X"54",X"04",X"10",X"00",X"00",
		X"10",X"04",X"14",X"14",X"05",X"50",X"01",X"40",X"05",X"50",X"14",X"14",X"10",X"04",X"00",X"00",
		X"10",X"04",X"10",X"04",X"14",X"14",X"05",X"50",X"01",X"40",X"01",X"40",X"01",X"40",X"00",X"00",
		X"15",X"54",X"10",X"14",X"00",X"50",X"01",X"40",X"05",X"00",X"14",X"04",X"15",X"54",X"00",X"00",
		X"95",X"56",X"95",X"56",X"95",X"56",X"95",X"56",X"95",X"56",X"95",X"56",X"95",X"55",X"01",X"55",
		X"30",X"55",X"3C",X"15",X"3F",X"01",X"3F",X"F0",X"3F",X"FC",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",
		X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",
		X"C0",X"00",X"C0",X"00",X"CA",X"AA",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",
		X"C0",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"00",X"00",X"00",X"00",
		X"30",X"AA",X"3C",X"2A",X"3F",X"02",X"3F",X"F0",X"3F",X"FC",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"15",X"55",X"15",X"55",X"15",X"55",X"15",X"55",
		X"15",X"55",X"15",X"55",X"15",X"55",X"15",X"55",X"15",X"55",X"15",X"55",X"15",X"55",X"15",X"55",
		X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",
		X"FE",X"AA",X"FF",X"EA",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"EA",X"AA",X"FE",X"AA",X"FF",X"EA",X"FF",X"FE",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"EA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AB",X"AA",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"BF",X"AF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AF",X"AB",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"BF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AE",X"AA",X"FE",
		X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"D5",X"55",X"DF",X"FF",X"D7",X"D7",X"F7",X"DD",X"F7",X"DD",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"DF",X"FF",X"F7",X"FF",X"F7",X"FF",
		X"FE",X"AA",X"FF",X"EA",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FD",X"57",X"FD",X"FD",X"FD",X"7D",
		X"AA",X"AA",X"AA",X"AF",X"AB",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"D7",X"FF",X"7D",X"FF",X"7D",X"FF",
		X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",
		X"F7",X"D7",X"F7",X"FF",X"F7",X"D7",X"F7",X"D5",X"F7",X"DD",X"F7",X"DD",X"F7",X"D5",X"D7",X"D7",
		X"D7",X"FF",X"5D",X"75",X"DF",X"DF",X"F7",X"D7",X"F7",X"D7",X"F7",X"D7",X"F7",X"D7",X"D7",X"DF",
		X"FF",X"7D",X"F5",X"7D",X"5F",X"FF",X"7D",X"7D",X"7D",X"FD",X"7D",X"FD",X"7D",X"7D",X"7D",X"7D",
		X"FF",X"FF",X"5D",X"5D",X"F7",X"F7",X"DD",X"DD",X"F7",X"F7",X"F7",X"77",X"7F",X"7F",X"7D",X"7D",
		X"FF",X"FF",X"5D",X"57",X"F7",X"FD",X"DF",X"5F",X"DF",X"5F",X"5F",X"FF",X"5F",X"55",X"DF",X"5F",
		X"D7",X"FF",X"5D",X"D5",X"FD",X"7F",X"7D",X"F5",X"7D",X"F5",X"7D",X"7F",X"7D",X"57",X"7D",X"D7",
		X"FF",X"FF",X"7D",X"57",X"D7",X"FD",X"DF",X"5F",X"5F",X"5F",X"5F",X"FF",X"DF",X"55",X"DF",X"5F",
		X"D7",X"7E",X"5D",X"DE",X"FF",X"DE",X"7D",X"DE",X"7D",X"7E",X"7D",X"FE",X"7D",X"FE",X"7D",X"DE",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"EA",X"AA",
		X"DF",X"FF",X"D5",X"55",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"75",X"F7",X"FD",X"5D",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",
		X"DF",X"FF",X"55",X"55",X"FF",X"FF",X"FF",X"FA",X"FF",X"A9",X"FA",X"95",X"A9",X"5A",X"95",X"AA",
		X"7D",X"7D",X"D7",X"D5",X"FF",X"FF",X"AF",X"FF",X"6A",X"FF",X"56",X"AB",X"A5",X"5A",X"AA",X"95",
		X"D7",X"FD",X"F5",X"57",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AF",X"FF",X"6A",X"BF",
		X"FF",X"FF",X"55",X"D5",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"57",X"FD",X"75",X"57",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"76",X"55",X"DE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AB",
		X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",X"A9",X"FA",X"95",X"A9",X"5A",X"96",X"AA",
		X"FF",X"A9",X"FA",X"95",X"A9",X"5A",X"95",X"AA",X"5A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"55",X"AA",X"A9",X"56",X"AA",X"A5",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"AB",X"FF",X"5A",X"AF",X"95",X"6A",X"AA",X"55",X"AA",X"A9",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"FF",X"AA",X"FF",X"56",X"AB",X"A5",X"5A",X"AA",X"95",
		X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"AF",X"FE",X"6A",X"BE",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"55",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"5A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FF",X"AB",X"EA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",
		X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",
		X"55",X"55",X"55",X"55",X"55",X"57",X"55",X"5F",X"55",X"5E",X"55",X"7E",X"55",X"FA",X"55",X"EA",
		X"FA",X"95",X"EA",X"55",X"E9",X"55",X"A9",X"55",X"A5",X"55",X"95",X"55",X"95",X"55",X"55",X"55",
		X"55",X"EE",X"55",X"EE",X"55",X"EE",X"55",X"EE",X"55",X"EE",X"55",X"EE",X"55",X"6E",X"55",X"6E",
		X"AF",X"EE",X"BF",X"EE",X"BF",X"EE",X"FF",X"EE",X"D7",X"EE",X"57",X"EE",X"55",X"EE",X"55",X"EE",
		X"55",X"5E",X"55",X"7E",X"55",X"FA",X"55",X"EA",X"57",X"EB",X"5F",X"AB",X"5E",X"AF",X"7E",X"95",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"57",X"55",X"5F",
		X"57",X"EE",X"5F",X"AE",X"5E",X"AE",X"7E",X"AE",X"FA",X"AE",X"EA",X"EE",X"EB",X"EE",X"AB",X"EE",
		X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"5E",X"55",X"5E",X"55",X"7E",X"55",X"FE",X"55",X"EE",
		X"57",X"E9",X"5F",X"A9",X"5E",X"A5",X"7E",X"95",X"FA",X"95",X"EA",X"55",X"E9",X"55",X"A9",X"55",
		X"55",X"55",X"55",X"57",X"55",X"D7",X"57",X"5D",X"57",X"5D",X"5D",X"DD",X"5D",X"DD",X"5D",X"5D",
		X"55",X"6E",X"55",X"6E",X"55",X"6E",X"55",X"6E",X"55",X"6E",X"55",X"6E",X"55",X"6E",X"55",X"6E",
		X"55",X"6E",X"55",X"6E",X"55",X"6E",X"55",X"6E",X"55",X"6E",X"55",X"6E",X"55",X"6E",X"55",X"6E",
		X"57",X"55",X"5D",X"55",X"DD",X"D5",X"5D",X"D5",X"5D",X"55",X"DD",X"55",X"DD",X"55",X"D5",X"55",
		X"A5",X"55",X"95",X"55",X"95",X"55",X"55",X"57",X"55",X"57",X"55",X"5D",X"55",X"5D",X"55",X"5D",
		X"55",X"5E",X"55",X"7E",X"55",X"FA",X"55",X"EA",X"57",X"E9",X"5F",X"A9",X"5E",X"A5",X"7E",X"95",
		X"FA",X"95",X"EA",X"55",X"E9",X"55",X"E9",X"55",X"E9",X"55",X"E9",X"55",X"E9",X"55",X"E9",X"55",
		X"55",X"5D",X"55",X"DD",X"57",X"5D",X"57",X"5D",X"5D",X"DD",X"5D",X"DD",X"5D",X"DD",X"5D",X"55",
		X"55",X"55",X"55",X"55",X"D5",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"BE",X"55",X"BA",X"56",X"F9",X"56",X"E9",X"5B",X"E5",X"5B",X"A5",X"6F",X"95",X"6E",X"95",
		X"BE",X"55",X"BA",X"55",X"F9",X"55",X"E9",X"55",X"E5",X"55",X"A5",X"55",X"95",X"55",X"95",X"55",
		X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"56",X"55",X"5B",X"55",X"5B",X"55",X"6F",X"55",X"6E",
		X"57",X"55",X"5D",X"D5",X"DD",X"D5",X"DD",X"55",X"5D",X"55",X"5D",X"55",X"5D",X"55",X"55",X"55",
		X"E9",X"55",X"E9",X"55",X"E9",X"55",X"E9",X"55",X"E9",X"57",X"E9",X"57",X"E9",X"5D",X"E9",X"5D",
		X"E9",X"5D",X"E9",X"5D",X"E9",X"55",X"E9",X"55",X"E9",X"55",X"E9",X"55",X"E9",X"55",X"E9",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"BE",X"55",X"BA",X"56",X"F9",X"56",X"E9",X"5B",X"E5",X"5B",X"A5",X"6F",X"95",X"6E",X"95",
		X"BE",X"55",X"BA",X"55",X"F9",X"55",X"E9",X"55",X"E5",X"55",X"A5",X"55",X"95",X"55",X"95",X"55",
		X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"56",X"55",X"5B",X"55",X"7B",X"55",X"EF",X"55",X"EE",
		X"E9",X"55",X"EB",X"55",X"EB",X"55",X"EB",X"55",X"EB",X"55",X"EB",X"55",X"EB",X"55",X"EB",X"D5",
		X"EB",X"D5",X"EB",X"D5",X"EB",X"D5",X"EB",X"F5",X"EB",X"F5",X"EB",X"FF",X"EB",X"FF",X"EB",X"FF",
		X"EB",X"FF",X"EB",X"FF",X"EB",X"FE",X"EB",X"FE",X"EB",X"FB",X"EB",X"FB",X"EB",X"EF",X"EB",X"EE",
		X"EB",X"BE",X"EB",X"BA",X"EA",X"F9",X"EA",X"E9",X"EB",X"E5",X"EB",X"A5",X"EF",X"95",X"EE",X"95",
		X"EE",X"55",X"EA",X"55",X"E9",X"55",X"E9",X"55",X"E5",X"55",X"E5",X"55",X"D5",X"55",X"D5",X"55",
		X"BE",X"55",X"BA",X"55",X"F9",X"55",X"E9",X"55",X"E5",X"55",X"A5",X"55",X"95",X"55",X"95",X"55",
		X"57",X"BE",X"5F",X"BA",X"7E",X"F9",X"7E",X"E9",X"FB",X"E5",X"FB",X"A5",X"EF",X"95",X"EE",X"95",
		X"02",X"EA",X"02",X"EA",X"02",X"EA",X"02",X"EA",X"02",X"EA",X"02",X"EA",X"02",X"EA",X"02",X"EA",
		X"02",X"FA",X"02",X"EA",X"02",X"EA",X"02",X"EA",X"02",X"EA",X"02",X"EA",X"02",X"EA",X"02",X"EA",
		X"00",X"0B",X"00",X"2B",X"00",X"2F",X"00",X"2E",X"00",X"AE",X"00",X"BE",X"00",X"BA",X"02",X"BA",
		X"C0",X"00",X"C0",X"00",X"C0",X"00",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"0A",X"00",X"0B",
		X"AE",X"AB",X"BE",X"AB",X"BA",X"AB",X"BA",X"AB",X"FA",X"AB",X"EA",X"AB",X"EA",X"AB",X"EA",X"AB",
		X"02",X"FB",X"02",X"EB",X"0A",X"EB",X"0B",X"EB",X"0B",X"AB",X"2B",X"AB",X"2F",X"AB",X"2E",X"AB",
		X"00",X"0B",X"00",X"2B",X"00",X"2F",X"00",X"2F",X"00",X"AF",X"00",X"BB",X"00",X"BB",X"02",X"BB",
		X"FF",X"00",X"FC",X"00",X"FC",X"00",X"FC",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"C0",X"00",
		X"00",X"FF",X"03",X"FC",X"03",X"FC",X"03",X"FC",X"0F",X"F0",X"0F",X"F0",X"0F",X"F0",X"3F",X"C0",
		X"00",X"00",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"3F",
		X"C0",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"03",X"00",X"03",
		X"3F",X"C0",X"3F",X"C0",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FC",X"00",X"FC",X"00",X"FC",X"00",
		X"00",X"3F",X"00",X"3F",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"03",X"FC",X"03",X"FC",X"03",X"FC",
		X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"3F",X"00",X"3F",X"00",X"3F",X"00",X"FF",X"00",X"FF",
		X"F0",X"00",X"F0",X"00",X"F0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"F0",X"0F",X"F0",X"0F",X"F0",X"3F",X"C0",X"3F",X"C0",X"3F",X"C0",X"FF",X"00",X"FF",X"00",
		X"02",X"EA",X"02",X"EA",X"02",X"EA",X"02",X"EA",X"02",X"EA",X"02",X"EA",X"02",X"EA",X"02",X"EB",
		X"02",X"EB",X"02",X"EB",X"02",X"EF",X"02",X"EC",X"02",X"AC",X"02",X"BC",X"02",X"B0",X"56",X"B0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AC",X"00",X"BC",X"00",X"B0",X"00",X"B0",X"00",X"F0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",
		X"AA",X"F0",X"AA",X"C0",X"AA",X"C0",X"AB",X"C0",X"AB",X"00",X"AB",X"00",X"AF",X"00",X"AC",X"00",
		X"AA",X"AB",X"AA",X"AB",X"AA",X"AF",X"AA",X"AC",X"AA",X"AC",X"AA",X"BC",X"AA",X"B0",X"AA",X"B0",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"35",X"00",X"5F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"54",X"00",
		X"01",X"5F",X"05",X"FF",X"07",X"FF",X"17",X"FF",X"17",X"FF",X"5F",X"FF",X"5F",X"FF",X"5F",X"FF",
		X"F5",X"40",X"FD",X"50",X"FD",X"50",X"FF",X"54",X"FF",X"D4",X"FF",X"D5",X"FF",X"D5",X"FF",X"D5",
		X"FF",X"D5",X"FF",X"D5",X"FF",X"D5",X"FF",X"D4",X"FF",X"54",X"FF",X"50",X"FD",X"50",X"F5",X"40",
		X"5F",X"FF",X"5F",X"FF",X"5F",X"FF",X"1F",X"FF",X"17",X"FF",X"07",X"FF",X"05",X"FF",X"01",X"7F",
		X"00",X"7F",X"00",X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"5F",X"05",X"FF",X"07",X"FF",X"17",X"FF",X"17",X"FF",X"5F",X"FF",X"5F",X"FF",X"5F",X"FF",
		X"01",X"5F",X"05",X"FF",X"07",X"FF",X"17",X"FF",X"17",X"FF",X"5F",X"FF",X"5F",X"FF",X"5F",X"FF",
		X"F5",X"7F",X"FD",X"5F",X"FD",X"5F",X"FF",X"57",X"FF",X"D7",X"FF",X"D5",X"FF",X"D5",X"FF",X"D5",
		X"F5",X"40",X"FD",X"50",X"FD",X"50",X"FF",X"54",X"FF",X"D4",X"FF",X"D5",X"FF",X"D5",X"FF",X"D5",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"54",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"F5",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"5F",X"00",X"57",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"35",X"00",X"FF",
		X"F5",X"55",X"D5",X"55",X"55",X"54",X"55",X"50",X"55",X"40",X"54",X"00",X"90",X"00",X"40",X"00",
		X"00",X"00",X"40",X"00",X"55",X"00",X"55",X"50",X"D5",X"54",X"F5",X"55",X"F5",X"55",X"F5",X"55",
		X"55",X"50",X"FF",X"55",X"FF",X"F5",X"FF",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"55",X"55",X"55",X"55",X"55",X"AA",X"AA",X"56",X"66",
		X"5F",X"FF",X"57",X"FF",X"15",X"7F",X"05",X"57",X"01",X"55",X"00",X"15",X"00",X"0A",X"00",X"01",
		X"00",X"03",X"00",X"FF",X"0F",X"FF",X"3F",X"FF",X"FF",X"FF",X"7F",X"FF",X"7F",X"FF",X"5F",X"FF",
		X"55",X"99",X"16",X"64",X"05",X"90",X"05",X"60",X"05",X"90",X"05",X"60",X"05",X"90",X"05",X"60",
		X"02",X"C0",X"02",X"FF",X"0F",X"FF",X"3F",X"FF",X"FF",X"FF",X"7F",X"FF",X"7F",X"FF",X"5F",X"FF",
		X"5F",X"FF",X"57",X"FF",X"15",X"7F",X"05",X"57",X"01",X"55",X"02",X"D5",X"02",X"EA",X"02",X"C1",
		X"02",X"C0",X"02",X"C0",X"55",X"C0",X"55",X"50",X"D5",X"54",X"F5",X"55",X"F5",X"55",X"F5",X"55",
		X"F5",X"55",X"D5",X"55",X"55",X"54",X"55",X"50",X"55",X"40",X"56",X"C0",X"92",X"C0",X"62",X"C0",
		X"55",X"99",X"15",X"64",X"05",X"90",X"05",X"60",X"05",X"90",X"55",X"55",X"FF",X"FF",X"55",X"55",
		X"02",X"C0",X"02",X"C0",X"02",X"C0",X"02",X"C0",X"03",X"C0",X"55",X"55",X"FF",X"FF",X"55",X"55",
		X"02",X"C0",X"02",X"C0",X"02",X"C0",X"02",X"C0",X"03",X"C0",X"15",X"55",X"BF",X"FF",X"15",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"FF",X"FF",X"55",X"55",
		X"95",X"55",X"95",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"54",X"55",X"54",X"55",X"50",
		X"55",X"50",X"55",X"54",X"55",X"54",X"55",X"55",X"55",X"55",X"95",X"55",X"95",X"55",X"95",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"6A",X"AA",X"6A",X"AA",X"6A",X"AA",X"55",X"55",X"55",X"55",X"15",X"55",X"15",X"55",X"05",X"55",
		X"05",X"55",X"15",X"55",X"15",X"55",X"55",X"55",X"55",X"55",X"6A",X"AA",X"6A",X"AA",X"6A",X"AA",
		X"D5",X"55",X"D5",X"55",X"D5",X"55",X"55",X"55",X"55",X"55",X"55",X"54",X"55",X"54",X"55",X"50",
		X"55",X"50",X"55",X"54",X"55",X"54",X"55",X"55",X"55",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"7F",X"FF",X"7F",X"FF",X"7F",X"FF",X"55",X"55",X"55",X"55",X"15",X"55",X"15",X"55",X"05",X"55",
		X"05",X"55",X"15",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"7F",X"FF",X"7F",X"FF",X"7F",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"5F",X"F5",
		X"03",X"C0",X"03",X"C0",X"02",X"C0",X"02",X"C0",X"02",X"C0",X"02",X"C0",X"02",X"C0",X"02",X"C0",
		X"02",X"C0",X"02",X"C0",X"02",X"C0",X"02",X"C0",X"02",X"C0",X"02",X"C0",X"02",X"C0",X"02",X"C0",
		X"02",X"C0",X"02",X"C0",X"02",X"C0",X"02",X"C0",X"02",X"C0",X"02",X"C0",X"02",X"C0",X"03",X"C0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"5F",X"F5",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"FF",X"0F",X"FF",X"0F",X"FF",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"F0",X"FF",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"C0",X"FC",X"00",X"F0",X"00",X"F0",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"BF",X"AA",X"AF",
		X"D5",X"5F",X"F5",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"9F",X"AA",X"9F",X"AA",X"9F",X"AA",X"9F",X"AA",X"9F",X"AA",X"9F",X"AA",X"9F",X"AA",X"9F",
		X"FD",X"5A",X"FF",X"D5",X"FF",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"5A",X"AA",X"D5",X"AA",X"FD",X"5A",X"FF",X"D5",X"FF",X"FD",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"5A",X"AA",X"D5",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"95",X"A5",X"5F",X"57",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A9",X"AA",X"55",X"95",X"7F",X"5F",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A5",
		X"A9",X"57",X"55",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",
		X"FD",X"5A",X"FF",X"D5",X"FF",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"5A",X"AA",X"D5",X"AA",X"FD",X"5A",X"FF",X"D5",X"FF",X"FD",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"5A",X"AA",X"D5",X"A5",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A9",X"AA",X"55",X"95",X"7F",X"5F",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"95",X"A5",X"5F",X"57",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"A9",X"57",X"55",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"9F",X"AA",X"9F",X"AA",X"9F",X"AA",X"9F",X"AA",X"9F",X"AA",X"9F",X"AA",X"9F",X"AA",X"9F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"7F",X"FF",X"5F",X"FF",X"DF",X"FF",X"DF",X"FF",X"DF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"55",X"FF",X"FD",X"7F",X"FF",X"7F",X"FD",X"7F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"FD",X"FF",X"FF",X"FF",X"FF",
		X"FD",X"57",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"7F",X"FF",X"7F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"FF",X"DF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",
		X"FF",X"DF",X"FF",X"DF",X"FF",X"DF",X"FF",X"DF",X"FF",X"DF",X"FF",X"DF",X"FF",X"DF",X"FF",X"DF",
		X"FD",X"FD",X"FF",X"FF",X"FF",X"F7",X"FF",X"FD",X"55",X"FD",X"FD",X"7F",X"FF",X"5F",X"FF",X"DF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"7F",X"D7",X"7F",X"F7",X"7F",X"F7",X"7F",X"F7",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FD",X"FF",X"F7",X"F5",X"F7",X"DD",X"F7",X"FF",
		X"7F",X"FF",X"7F",X"FF",X"7F",X"FF",X"7D",X"FF",X"FD",X"7D",X"FF",X"5F",X"7F",X"DF",X"7F",X"D7",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"F7",X"D7",X"D5",X"F7",X"FD",X"DF",X"F7",X"DF",X"F7",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"FF",X"7F",X"F7",X"7F",X"FD",X"FF",X"FD",X"FF",X"DD",X"F5",
		X"FF",X"DF",X"FF",X"F7",X"FF",X"F5",X"FF",X"DF",X"5F",X"D7",X"D7",X"F7",X"FF",X"F7",X"57",X"F7",
		X"FF",X"FF",X"7F",X"FF",X"FD",X"FD",X"F7",X"FF",X"F7",X"D7",X"F7",X"F5",X"F7",X"FD",X"FD",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FD",X"FF",X"FD",X"FD",X"F7",X"FF",X"77",X"FF",X"F7",X"D5",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"5F",X"7F",X"5F",X"5F",X"DF",X"FF",X"DF",X"5F",X"DF",
		X"FF",X"FD",X"FF",X"FD",X"7F",X"FD",X"FF",X"FD",X"DF",X"FD",X"5F",X"FD",X"D5",X"FD",X"FF",X"FD",
		X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",X"FD",X"FD",X"7D",X"7D",X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",
		X"F7",X"DF",X"DF",X"DF",X"FD",X"5F",X"F7",X"7F",X"5F",X"55",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F7",X"FF",X"F7",X"FF",X"F5",X"FF",X"7D",X"7F",X"FF",X"55",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FD",X"57",X"F7",X"F7",X"F7",X"FF",X"F7",X"7F",X"55",X"55",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FD",X"F7",X"F7",X"F7",X"FF",X"77",X"FD",X"DF",X"57",X"D5",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FD",X"FF",X"7D",X"FF",X"FD",X"7F",X"FF",X"5F",X"FF",X"D5",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FD",X"FF",X"FD",X"7F",X"7F",X"7D",X"57",X"57",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"F7",X"FF",X"F5",X"FF",X"FD",X"DF",X"FD",X"55",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F7",X"FD",X"F7",X"FD",X"F5",X"FF",X"FD",X"7F",X"5F",X"55",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"F7",X"7F",X"7F",X"7F",X"FF",X"5F",X"FD",X"D5",X"55",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"5F",X"FD",X"7F",X"FD",X"FF",X"FF",X"FD",X"FF",X"F7",X"55",X"5F",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"DF",X"FF",X"DF",X"FF",X"5F",X"FF",X"7F",X"FF",X"7F",X"FF",X"55",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"D5",X"FD",X"5A",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"D5",X"7F",X"5A",X"55",X"AA",X"A9",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"57",X"FF",X"A5",X"5F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"9F",X"AA",X"9F",X"AA",X"9F",X"AA",X"9F",X"AA",X"9F",X"AA",X"9D",X"AA",X"95",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FD",X"FF",X"D5",X"FD",X"5A",X"D5",X"AA",X"5A",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"D5",X"AA",X"5A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"D5",X"FD",X"5A",
		X"FF",X"FF",X"FF",X"FD",X"FF",X"D5",X"FD",X"5A",X"D5",X"AA",X"5A",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"D5",X"AA",X"5A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"95",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"7F",X"FF",X"55",X"FF",X"A9",X"57",X"AA",X"A5",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"5F",X"FF",X"95",X"7F",X"AA",X"55",X"AA",X"A9",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"57",X"FF",X"A5",X"5F",
		X"AA",X"95",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"7F",X"FF",X"55",X"FF",X"A9",X"57",X"AA",X"A5",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"5F",X"FF",X"95",X"7F",X"AA",X"55",X"AA",X"A9",X"AA",X"AA",
		X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",X"57",X"FD",X"A5",X"5D",
		X"AA",X"95",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"55",X"95",X"7D",X"5F",X"FD",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A5",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"95",X"AA",X"9D",X"AA",X"9F",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"5A",X"AA",X"D5",X"AA",
		X"55",X"54",X"55",X"50",X"55",X"40",X"55",X"00",X"54",X"00",X"50",X"00",X"40",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"56",X"AA",X"56",X"AA",X"56",X"AA",
		X"54",X"00",X"54",X"00",X"54",X"00",X"54",X"00",X"54",X"00",X"54",X"00",X"54",X"00",X"54",X"00",
		X"54",X"00",X"54",X"00",X"54",X"00",X"54",X"00",X"54",X"00",X"54",X"00",X"54",X"00",X"54",X"00",
		X"58",X"00",X"6C",X"00",X"BC",X"00",X"F8",X"00",X"6A",X"AA",X"7F",X"FF",X"56",X"AA",X"56",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"AA",X"AA",X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"55",X"54",X"55",X"54",X"55",X"50",X"55",X"50",X"55",X"40",X"55",X"40",X"55",X"00",X"55",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"54",X"00",X"54",X"00",X"50",X"00",X"50",X"00",X"40",X"00",X"40",X"00",X"00",X"00",X"00",X"00",
		X"D5",X"54",X"D5",X"54",X"F5",X"50",X"F5",X"50",X"FD",X"40",X"FD",X"40",X"FF",X"00",X"FF",X"00",
		X"FF",X"C0",X"FF",X"C0",X"FF",X"F0",X"FF",X"F0",X"FF",X"FC",X"FF",X"FC",X"BF",X"FF",X"BF",X"FF",
		X"AF",X"FF",X"2F",X"FF",X"2B",X"FF",X"0B",X"FF",X"0A",X"FF",X"02",X"FF",X"02",X"BF",X"00",X"BF",
		X"C0",X"00",X"C0",X"00",X"F0",X"00",X"F0",X"00",X"FC",X"00",X"FC",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"AF",X"00",X"2F",X"00",X"2B",X"00",X"0B",X"00",X"0A",X"00",X"02",X"00",X"02",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"FB",X"AF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",X"FF",X"FF",X"FB",X"BF",X"AB",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",X"FF",X"FF",X"FF",X"AB",X"BF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"EA",X"AF",X"EA",X"AF",X"AA",X"BF",X"AA",X"FF",X"AA",X"FF",X"AB",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"6A",X"6A",X"A9",X"59",X"65",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FD",X"FF",X"F5",X"FF",X"F5",X"FF",X"D5",X"FD",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"7F",X"FF",X"7F",X"FF",X"5F",X"FF",X"55",X"FF",X"55",X"5F",X"55",X"5F",X"55",X"5F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"EA",X"AF",X"EA",X"AF",X"FA",X"AB",X"FE",X"AB",X"FE",X"AB",X"FF",X"AB",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"BF",
		X"FF",X"FF",X"FF",X"FE",X"FF",X"FA",X"FF",X"FA",X"FF",X"FA",X"FF",X"FA",X"FF",X"FA",X"FF",X"FE",
		X"EA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FF",X"AA",X"FF",X"AB",X"FF",X"AB",X"FF",X"A7",X"FA",
		X"AA",X"AB",X"AA",X"AA",X"AA",X"AA",X"EA",X"AA",X"FA",X"AA",X"FE",X"AA",X"FE",X"AA",X"BE",X"65",
		X"FF",X"FF",X"FF",X"FF",X"BF",X"FF",X"AF",X"FF",X"AF",X"FF",X"AF",X"FF",X"6F",X"FF",X"AF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"F5",X"FF",X"D5",X"FF",X"D5",X"FF",X"D5",X"FF",X"D5",
		X"FF",X"55",X"55",X"55",X"55",X"5F",X"55",X"7F",X"55",X"FF",X"55",X"FF",X"57",X"FF",X"57",X"FF",
		X"55",X"55",X"55",X"55",X"F5",X"55",X"FD",X"55",X"FD",X"55",X"FD",X"55",X"FD",X"55",X"FD",X"55",
		X"57",X"FF",X"57",X"FF",X"57",X"FF",X"57",X"FF",X"57",X"FF",X"57",X"FF",X"57",X"FF",X"57",X"FF",
		X"FF",X"D5",X"FF",X"D5",X"FF",X"D5",X"FF",X"D5",X"FF",X"D5",X"FF",X"F5",X"FF",X"F5",X"FF",X"FD",
		X"57",X"FF",X"55",X"FF",X"55",X"FF",X"55",X"7F",X"55",X"5F",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FD",X"55",X"FD",X"55",X"FD",X"55",X"F5",X"55",X"D5",X"55",X"55",X"55",X"7D",X"55",X"FD",X"55",
		X"57",X"FF",X"57",X"FF",X"57",X"FF",X"57",X"FF",X"55",X"57",X"55",X"57",X"55",X"57",X"55",X"57",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F5",X"5F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"FE",X"BF",X"FA",X"BF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AF",X"FF",X"AA",X"BF",
		X"AA",X"AF",X"AA",X"AB",X"AA",X"AB",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"E5",X"96",
		X"AA",X"AA",X"AA",X"AA",X"AF",X"AA",X"FF",X"FA",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"BA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AB",X"AA",X"AF",X"AA",X"AF",X"96",X"AF",
		X"FF",X"FF",X"FA",X"AA",X"FA",X"AA",X"FA",X"AA",X"FF",X"AA",X"FF",X"EA",X"FF",X"F9",X"FF",X"FA",
		X"FF",X"F5",X"FF",X"F5",X"FF",X"F5",X"FF",X"F5",X"FF",X"F5",X"FF",X"F5",X"FF",X"F5",X"FF",X"F5",
		X"55",X"6F",X"55",X"5F",X"55",X"5F",X"55",X"5F",X"55",X"5F",X"55",X"5F",X"55",X"5F",X"55",X"5F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"D5",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"57",X"55",X"5F",X"55",X"7F",X"57",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FD",X"FF",X"F5",X"5F",X"D5",X"55",X"55",X"55",X"55",X"55",X"45",X"FD",X"01",
		X"55",X"57",X"55",X"57",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"45",X"5F",X"50",X"5F",
		X"FF",X"F5",X"FF",X"F5",X"FF",X"F5",X"FF",X"F5",X"FF",X"F5",X"FF",X"F5",X"FF",X"F5",X"FF",X"F5",
		X"FF",X"F0",X"FF",X"F0",X"FF",X"F0",X"FF",X"F0",X"FF",X"F0",X"FF",X"F0",X"FF",X"C0",X"FF",X"C0",
		X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FA",X"FF",X"FA",X"FF",X"FA",X"FF",X"FF",X"FF",X"FF",X"BF",X"FF",X"BF",X"FF",
		X"7F",X"FF",X"7F",X"FF",X"7F",X"FF",X"7F",X"FF",X"7F",X"FF",X"7F",X"FF",X"7F",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"E9",X"AA",X"FA",X"9A",X"FA",X"95",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"FF",X"BF",X"FA",X"BF",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"AF",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"FF",
		X"AF",X"FF",X"AB",X"FF",X"AB",X"FF",X"AA",X"FF",X"AA",X"FF",X"AA",X"FF",X"9A",X"BF",X"6A",X"BF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FA",X"AA",X"FE",X"AA",X"FF",X"AA",X"FF",X"AA",X"FF",X"E9",
		X"BA",X"AA",X"AA",X"AA",X"AA",X"AF",X"AA",X"FF",X"AB",X"FF",X"AF",X"FF",X"AF",X"FF",X"AF",X"FF",
		X"F6",X"55",X"F5",X"55",X"F5",X"55",X"F5",X"55",X"F5",X"55",X"F5",X"55",X"F5",X"55",X"F5",X"55",
		X"5F",X"FF",X"5F",X"FF",X"5F",X"FF",X"5F",X"FF",X"5F",X"FF",X"5F",X"FF",X"5F",X"FF",X"5F",X"FF",
		X"FF",X"D5",X"FF",X"D5",X"FF",X"D5",X"FF",X"D5",X"FF",X"D5",X"FF",X"D5",X"FF",X"55",X"FF",X"55",
		X"55",X"7F",X"55",X"7F",X"55",X"7F",X"55",X"7F",X"55",X"7F",X"55",X"7F",X"55",X"7F",X"55",X"FF",
		X"55",X"FF",X"55",X"FF",X"55",X"FF",X"57",X"FF",X"5F",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"55",X"FD",X"55",X"F5",X"55",X"D5",X"55",X"55",X"55",X"51",X"55",X"55",X"57",X"41",X"FF",
		X"5F",X"FF",X"57",X"FF",X"55",X"FF",X"55",X"5F",X"55",X"55",X"55",X"55",X"5F",X"55",X"1F",X"FD",
		X"F5",X"55",X"F5",X"55",X"F5",X"55",X"F5",X"55",X"F5",X"55",X"F4",X"55",X"F5",X"55",X"F5",X"45",
		X"F1",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"C0",X"00",X"C0",X"00",
		X"0F",X"FF",X"0F",X"FF",X"0F",X"FF",X"0F",X"FF",X"0F",X"FF",X"0F",X"FF",X"0F",X"FF",X"0F",X"FF",
		X"FF",X"FA",X"FF",X"EA",X"FF",X"AA",X"FE",X"AA",X"FE",X"AA",X"FA",X"AA",X"FA",X"A9",X"FA",X"5A",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"FF",X"AB",X"FF",X"AF",X"FF",X"AF",X"FF",X"AF",X"FF",X"6F",X"FF",
		X"AA",X"AF",X"AA",X"AB",X"AA",X"AB",X"EA",X"AA",X"FA",X"AA",X"F9",X"AA",X"FA",X"5A",X"FA",X"56",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AB",X"FF",X"AA",X"AF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"5F",X"FF",X"5F",X"FF",X"5F",X"FF",X"5F",X"FF",X"5F",X"FF",
		X"F5",X"55",X"F5",X"55",X"F5",X"55",X"F5",X"55",X"F5",X"55",X"F5",X"55",X"F5",X"55",X"F5",X"55",
		X"F5",X"55",X"F5",X"55",X"FD",X"55",X"FD",X"55",X"FD",X"55",X"FF",X"55",X"FF",X"D5",X"FF",X"F5",
		X"5F",X"FF",X"57",X"FF",X"57",X"FF",X"55",X"FF",X"55",X"5F",X"55",X"55",X"51",X"55",X"55",X"45",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"D5",X"FD",X"55",X"55",X"55",X"55",X"57",X"55",X"1F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"D4",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"5F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"BF",X"FF",X"BF",X"FF",X"BF",X"FF",
		X"5F",X"FF",X"5F",X"FF",X"5F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"FF",X"5F",X"FF",X"5F",X"FF",X"5F",X"FF",X"7F",X"FF",X"FF",X"F5",X"FF",X"F5",X"FF",X"F5",
		X"FD",X"55",X"FD",X"55",X"FD",X"55",X"F5",X"55",X"D5",X"55",X"55",X"55",X"51",X"55",X"05",X"55",
		X"FD",X"55",X"FD",X"55",X"FD",X"55",X"FD",X"55",X"FD",X"55",X"FD",X"55",X"FD",X"55",X"FD",X"55",
		X"FF",X"FA",X"FF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FA",X"AA",X"FE",X"AA",X"FE",X"59",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EB",X"FF",X"AB",X"FA",
		X"AB",X"AA",X"AA",X"AA",X"AA",X"BF",X"AA",X"FF",X"AB",X"FE",X"AB",X"FE",X"9B",X"FF",X"6B",X"FF",
		X"57",X"FF",X"57",X"FF",X"57",X"FF",X"57",X"FF",X"57",X"FF",X"57",X"FF",X"57",X"FF",X"57",X"FF",
		X"57",X"FF",X"57",X"FF",X"57",X"FF",X"57",X"FF",X"55",X"FF",X"55",X"57",X"41",X"57",X"01",X"57",
		X"AA",X"AF",X"AA",X"AB",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"6B",X"A5",X"AB",
		X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",
		X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7D",X"FD",X"7D",
		X"FD",X"7D",X"FD",X"75",X"FD",X"75",X"FD",X"75",X"FD",X"55",X"FD",X"55",X"FD",X"55",X"FD",X"55",
		X"FD",X"55",X"FD",X"55",X"FD",X"55",X"FD",X"55",X"FD",X"55",X"F5",X"55",X"F5",X"55",X"F5",X"55",
		X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"7D",X"7F",
		X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"6F",X"FD",X"6F",
		X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7D",X"FD",X"7D",
		X"D5",X"55",X"D5",X"55",X"D5",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"7D",X"7F",X"7D",X"7F",X"5D",X"7F",X"5D",X"7F",X"5D",X"7F",X"55",X"7F",X"55",X"7F",X"55",X"7F",
		X"FD",X"6F",X"FD",X"6F",X"FD",X"6E",X"FD",X"6E",X"FD",X"6E",X"FD",X"AE",X"FD",X"BB",X"FD",X"BB",
		X"FD",X"7D",X"FD",X"75",X"FD",X"75",X"FD",X"75",X"FD",X"55",X"BD",X"55",X"BD",X"55",X"BD",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"7F",X"55",X"7F",X"55",X"7F",X"55",X"7F",X"55",X"7F",X"55",X"7F",X"55",X"5F",X"55",X"5F",
		X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FC",X"3F",X"F3",X"0F",X"FF",X"CF",X"FF",X"CF",
		X"FE",X"BB",X"FE",X"EB",X"FE",X"EB",X"FA",X"EB",X"FB",X"AB",X"FB",X"AB",X"EB",X"AB",X"EE",X"AB",
		X"BD",X"55",X"BD",X"55",X"BD",X"5F",X"BF",X"7F",X"BD",X"7F",X"BD",X"FD",X"B5",X"F6",X"97",X"F6",
		X"55",X"55",X"55",X"55",X"55",X"55",X"F5",X"55",X"FF",X"55",X"7F",X"F5",X"97",X"FD",X"A9",X"FD",
		X"AA",X"A1",X"AA",X"85",X"AA",X"85",X"AA",X"15",X"AF",X"14",X"AC",X"54",X"A8",X"5B",X"A1",X"52",
		X"4A",X"AA",X"52",X"AA",X"54",X"AA",X"05",X"2A",X"BD",X"4A",X"EF",X"52",X"AA",X"D4",X"AF",X"D4",
		X"55",X"5A",X"55",X"6A",X"55",X"6B",X"F5",X"5A",X"FF",X"55",X"7F",X"F5",X"97",X"FD",X"A5",X"FD",
		X"55",X"5F",X"55",X"57",X"55",X"57",X"55",X"57",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"C3",X"FF",X"C0",X"F3",X"00",X"FC",X"30",X"FD",X"70",X"FD",X"70",X"FD",X"70",X"FD",X"70",
		X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7E",X"FD",X"7E",X"FD",X"7E",X"FD",X"7A",
		X"EE",X"AB",X"AE",X"AB",X"BA",X"AB",X"BA",X"AF",X"BA",X"AD",X"EA",X"AD",X"EA",X"A5",X"56",X"A7",
		X"97",X"DA",X"9F",X"DA",X"5F",X"D6",X"7F",X"F5",X"7D",X"7F",X"FD",X"97",X"F5",X"A5",X"F6",X"AA",
		X"A9",X"F5",X"A5",X"F5",X"A7",X"D5",X"97",X"D5",X"5F",X"55",X"FF",X"55",X"7D",X"55",X"7D",X"55",
		X"85",X"5B",X"85",X"54",X"95",X"15",X"94",X"05",X"94",X"F1",X"93",X"FE",X"8F",X"FE",X"8F",X"FF",
		X"EB",X"D4",X"BE",X"D2",X"3F",X"52",X"41",X"4A",X"55",X"2A",X"54",X"AA",X"A4",X"AA",X"12",X"AA",
		X"7D",X"70",X"7D",X"70",X"5D",X"70",X"5D",X"70",X"5D",X"70",X"55",X"70",X"55",X"70",X"55",X"70",
		X"FD",X"79",X"FD",X"77",X"FD",X"5F",X"FD",X"7E",X"FD",X"FA",X"F7",X"EA",X"DF",X"AA",X"DF",X"5A",
		X"F5",X"00",X"FD",X"40",X"BF",X"50",X"AF",X"D4",X"AB",X"F5",X"AA",X"FD",X"AA",X"BF",X"AA",X"9F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"50",X"00",X"D4",X"00",
		X"00",X"55",X"00",X"15",X"00",X"15",X"00",X"05",X"00",X"05",X"00",X"01",X"00",X"01",X"00",X"00",
		X"55",X"70",X"55",X"70",X"55",X"70",X"55",X"70",X"55",X"70",X"55",X"A0",X"5A",X"B0",X"6A",X"BF",
		X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"AD",X"7F",X"EA",X"7F",X"EA",X"BF",
		X"DF",X"D6",X"F7",X"F5",X"FD",X"FD",X"FD",X"7F",X"FD",X"DF",X"FD",X"F7",X"FD",X"79",X"FD",X"7B",
		X"AA",X"70",X"A9",X"F0",X"57",X"FA",X"5F",X"EA",X"FF",X"AA",X"FD",X"AA",X"FD",X"6A",X"7F",X"5A",
		X"F5",X"00",X"BD",X"7F",X"BF",X"5F",X"AF",X"D7",X"AB",X"F5",X"AA",X"FD",X"AA",X"7F",X"A9",X"7F",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"6A",X"AA",X"5A",X"AA",X"D0",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"A9",X"AA",X"A5",X"00",X"05",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",X"00",X"00",
		X"5A",X"AA",X"55",X"AA",X"55",X"55",X"55",X"55",X"55",X"55",X"57",X"55",X"57",X"D5",X"57",X"F7",
		X"AA",X"7F",X"A5",X"7F",X"55",X"5F",X"55",X"5F",X"55",X"5F",X"75",X"5F",X"F5",X"5F",X"F5",X"5F",
		X"FD",X"7B",X"FD",X"7B",X"FD",X"7B",X"FD",X"7B",X"FD",X"7B",X"FD",X"7B",X"FD",X"7B",X"FD",X"7B",
		X"5F",X"D6",X"57",X"F5",X"51",X"FD",X"50",X"7F",X"50",X"1F",X"50",X"07",X"50",X"01",X"50",X"00",
		X"A5",X"FF",X"97",X"FF",X"5F",X"FD",X"7F",X"F4",X"FF",X"D0",X"FF",X"40",X"FD",X"00",X"74",X"00",
		X"E0",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"5B",X"56",X"AA",
		X"57",X"FF",X"57",X"F7",X"57",X"D5",X"57",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"D5",X"55",
		X"F5",X"5F",X"F5",X"5F",X"F5",X"5F",X"75",X"5F",X"55",X"5F",X"55",X"5F",X"55",X"7F",X"55",X"7F",
		X"5F",X"FF",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"DF",X"FF",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"F5",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"5A",X"EB",X"55",X"AA",X"55",X"57",X"55",X"5A",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"A5",X"55",X"A9",X"55",X"AA",X"AA",X"AB",X"AA",X"56",X"AB",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"FF",X"5A",X"7F",X"AA",X"7F",X"AE",X"BF",X"A9",X"7F",X"55",X"7F",X"55",X"5F",X"55",X"5F",
		X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"FF",X"FD",X"FF",
		X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",
		X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"7F",
		X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",
		X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",
		X"FF",X"7F",X"FF",X"7F",X"FF",X"7F",X"FE",X"7F",X"FF",X"7F",X"FF",X"7F",X"FF",X"7F",X"FF",X"7F",
		X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",
		X"FF",X"FF",X"FF",X"EB",X"FF",X"B0",X"FF",X"C0",X"FF",X"B0",X"FF",X"EB",X"F7",X"F5",X"F5",X"57",
		X"FD",X"7F",X"0D",X"7F",X"31",X"7F",X"01",X"7F",X"01",X"7F",X"0D",X"7F",X"FD",X"7F",X"FD",X"7F",
		X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"FF",X"FD",X"FF",
		X"FF",X"6F",X"FF",X"7F",X"FB",X"7F",X"FA",X"7F",X"EB",X"6F",X"EF",X"6F",X"BF",X"AF",X"BE",X"BF",
		X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",
		X"F5",X"57",X"FD",X"5F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",
		X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",X"FF",X"FA",X"FF",X"FE",X"FF",X"FE",X"FF",X"EE",
		X"AB",X"7F",X"EE",X"BF",X"AE",X"BF",X"EE",X"6F",X"EA",X"7F",X"EF",X"6F",X"AE",X"BF",X"AA",X"7F",
		X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",
		X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",
		X"FF",X"EA",X"FF",X"AA",X"FF",X"AA",X"FF",X"EA",X"FF",X"FA",X"FF",X"BA",X"FE",X"AA",X"FF",X"AA",
		X"AA",X"7F",X"AB",X"7F",X"AA",X"BF",X"AA",X"BF",X"AB",X"BF",X"AA",X"6F",X"AA",X"7F",X"AA",X"BF",
		X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"FF",X"FD",X"FF",
		X"FF",X"AA",X"FE",X"AA",X"FA",X"BA",X"FE",X"EA",X"FF",X"EA",X"FF",X"AA",X"FE",X"BA",X"FE",X"EA",
		X"AA",X"7F",X"AE",X"BF",X"AB",X"6F",X"AA",X"7F",X"AA",X"BF",X"AF",X"7F",X"AA",X"7F",X"BB",X"7F",
		X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",X"FF",X"EB",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"57",X"55",X"5F",X"55",X"5F",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"D5",X"55",X"F5",X"55",X"F5",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"AB",X"56",X"BF",X"5A",X"FF",X"5B",X"FF",X"5B",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"F5",X"55",X"FD",X"55",X"FF",X"55",X"FF",X"55",X"C0",X"0F",
		X"55",X"5F",X"5D",X"5F",X"5F",X"5F",X"5F",X"7F",X"5F",X"FF",X"5F",X"FF",X"7F",X"F5",X"FF",X"15",
		X"F5",X"55",X"F5",X"55",X"F5",X"55",X"F5",X"55",X"F5",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"57",X"D5",X"5F",X"F5",X"5F",X"F5",X"5F",X"FD",X"5F",X"FD",X"5F",X"FF",
		X"6F",X"C0",X"6F",X"00",X"6F",X"00",X"7C",X"03",X"7C",X"3F",X"7F",X"FF",X"FF",X"F0",X"FF",X"00",
		X"00",X"03",X"00",X"03",X"00",X"00",X"00",X"03",X"C0",X"F3",X"03",X"EC",X"03",X"FC",X"00",X"F0",
		X"F1",X"55",X"05",X"55",X"15",X"55",X"C5",X"55",X"B5",X"55",X"F5",X"55",X"C5",X"55",X"01",X"55",
		X"57",X"FF",X"55",X"FD",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"EF",X"00",X"6B",X"C0",X"5B",X"C0",X"5A",X"F0",X"56",X"FC",X"56",X"BF",X"55",X"AF",X"55",X"6A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"0C",X"00",X"CC",X"C0",X"8C",X"C0",
		X"00",X"55",X"00",X"15",X"00",X"05",X"00",X"01",X"08",X"80",X"08",X"80",X"08",X"80",X"00",X"00",
		X"4C",X"C5",X"4F",X"C5",X"53",X"15",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"01",X"40",X"05",X"50",X"15",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",X"FF",X"EB",X"FE",X"EF",X"FE",X"AF",X"FF",X"AF",X"FF",X"EF",
		X"FF",X"FB",X"FF",X"AB",X"FE",X"AF",X"FF",X"EA",X"FF",X"AB",X"FE",X"AF",X"FF",X"AB",X"FB",X"EA",
		X"AA",X"FF",X"AB",X"FF",X"EF",X"FF",X"EB",X"FF",X"EF",X"FF",X"AF",X"FF",X"AF",X"FF",X"AB",X"FF",
		X"FF",X"EA",X"FE",X"AA",X"FF",X"AB",X"FE",X"AF",X"FE",X"AB",X"FA",X"AB",X"FE",X"AB",X"FA",X"AB",
		X"FA",X"AA",X"FA",X"AB",X"FA",X"EB",X"FF",X"EA",X"FF",X"EA",X"FF",X"AE",X"FB",X"AF",X"FA",X"AB",
		X"BF",X"FF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"FF",X"FF",X"7F",X"FF",X"7F",X"FF",X"7F",
		X"FA",X"AB",X"FE",X"AB",X"FF",X"AB",X"FE",X"AF",X"FA",X"BF",X"FA",X"AF",X"FA",X"BF",X"FA",X"AF",
		X"FE",X"BF",X"FF",X"BF",X"FF",X"AF",X"FF",X"BF",X"FE",X"BF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",
		X"FE",X"AF",X"FE",X"AB",X"FF",X"AB",X"FF",X"AF",X"FF",X"AF",X"FE",X"AB",X"FA",X"EB",X"FA",X"EB",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",
		X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"7F",X"FF",X"7F",
		X"FB",X"EF",X"FF",X"AF",X"FF",X"BF",X"FE",X"BF",X"FF",X"BF",X"FF",X"EF",X"FF",X"AF",X"FF",X"BB",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"A9",X"AA",X"9A",X"AA",X"5A",X"A6",X"56",X"A5",X"76",X"A7",X"76",
		X"95",X"5A",X"A6",X"5A",X"AA",X"9A",X"AA",X"9A",X"AA",X"5A",X"A6",X"7A",X"AA",X"9A",X"AA",X"AA",
		X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"55",
		X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"FD",X"7F",X"5D",X"7F",
		X"F5",X"55",X"F5",X"55",X"F5",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"55",X"55",X"AA",X"A9",
		X"55",X"7F",X"55",X"7F",X"55",X"7F",X"55",X"7F",X"55",X"7F",X"75",X"7F",X"65",X"7F",X"75",X"7F",
		X"AA",X"A9",X"AA",X"A9",X"AA",X"A9",X"AA",X"A9",X"AA",X"A9",X"AA",X"A9",X"AA",X"A9",X"AA",X"A9",
		X"E5",X"7F",X"B5",X"7F",X"E5",X"7F",X"B5",X"7F",X"E5",X"7F",X"B5",X"7F",X"E5",X"7F",X"95",X"7F",
		X"AA",X"A9",X"AA",X"A9",X"AA",X"A9",X"AA",X"A9",X"AA",X"A9",X"AA",X"A9",X"AA",X"A9",X"AA",X"A9",
		X"D5",X"7F",X"95",X"7F",X"5D",X"7F",X"5D",X"7F",X"5D",X"7F",X"7D",X"7F",X"7D",X"7F",X"7D",X"7F",
		X"55",X"55",X"40",X"00",X"4F",X"33",X"4C",X"33",X"4C",X"33",X"4C",X"33",X"4F",X"3F",X"55",X"55",
		X"55",X"55",X"00",X"00",X"3C",X"FC",X"30",X"30",X"3C",X"30",X"0C",X"30",X"3C",X"30",X"55",X"55",
		X"55",X"55",X"00",X"00",X"FC",X"C3",X"CC",X"FF",X"CC",X"FF",X"CC",X"C3",X"FC",X"C3",X"55",X"55",
		X"55",X"55",X"00",X"00",X"3C",X"FC",X"30",X"CC",X"3C",X"FC",X"30",X"CC",X"3C",X"CC",X"55",X"55",
		X"55",X"55",X"01",X"00",X"F1",X"00",X"C1",X"00",X"F1",X"00",X"31",X"00",X"F1",X"00",X"55",X"55",
		X"55",X"55",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"55",X"55",
		X"55",X"55",X"01",X"00",X"F1",X"3C",X"C1",X"0C",X"F1",X"0C",X"31",X"0C",X"F1",X"3F",X"55",X"55",
		X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",
		X"55",X"55",X"00",X"00",X"0F",X"F0",X"0C",X"30",X"0C",X"30",X"0C",X"30",X"0F",X"F0",X"55",X"55",
		X"55",X"55",X"00",X"00",X"03",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"03",X"F0",X"55",X"55",
		X"55",X"55",X"00",X"00",X"0F",X"F0",X"00",X"30",X"0F",X"F0",X"0C",X"00",X"0F",X"F0",X"55",X"55",
		X"55",X"55",X"00",X"00",X"0F",X"F0",X"00",X"30",X"0F",X"F0",X"00",X"30",X"0F",X"F0",X"55",X"55",
		X"55",X"55",X"00",X"00",X"0C",X"C0",X"0C",X"C0",X"0F",X"F0",X"00",X"C0",X"00",X"C0",X"55",X"55",
		X"55",X"55",X"00",X"00",X"0F",X"F0",X"0C",X"00",X"0F",X"F0",X"00",X"30",X"0F",X"F0",X"55",X"55",
		X"55",X"55",X"00",X"00",X"0F",X"F0",X"0C",X"00",X"0F",X"F0",X"0C",X"30",X"0F",X"F0",X"55",X"55",
		X"55",X"55",X"00",X"00",X"0F",X"F0",X"00",X"30",X"00",X"F0",X"00",X"C0",X"00",X"C0",X"55",X"55",
		X"55",X"55",X"00",X"00",X"0F",X"F0",X"0C",X"30",X"0F",X"F0",X"0C",X"30",X"0F",X"F0",X"55",X"55",
		X"55",X"55",X"00",X"00",X"0F",X"F0",X"0C",X"30",X"0F",X"F0",X"00",X"30",X"00",X"30",X"55",X"55",
		X"55",X"55",X"00",X"01",X"3F",X"C1",X"30",X"C1",X"30",X"C1",X"30",X"C1",X"3F",X"C1",X"55",X"55",
		X"55",X"55",X"00",X"01",X"0F",X"01",X"03",X"01",X"03",X"01",X"03",X"01",X"0F",X"C1",X"55",X"55",
		X"55",X"55",X"00",X"01",X"3F",X"C1",X"00",X"C1",X"3F",X"C1",X"30",X"01",X"3F",X"C1",X"55",X"55",
		X"55",X"55",X"00",X"01",X"3F",X"C1",X"00",X"C1",X"3F",X"C1",X"00",X"C1",X"3F",X"C1",X"55",X"55",
		X"55",X"55",X"00",X"01",X"33",X"01",X"33",X"01",X"3F",X"C1",X"03",X"01",X"03",X"01",X"55",X"55",
		X"55",X"55",X"00",X"01",X"3F",X"C1",X"30",X"01",X"3F",X"C1",X"00",X"C1",X"3F",X"C1",X"55",X"55",
		X"55",X"55",X"00",X"01",X"3F",X"C1",X"30",X"01",X"3F",X"C1",X"30",X"C1",X"3F",X"C1",X"55",X"55",
		X"55",X"55",X"00",X"01",X"3F",X"C1",X"00",X"C1",X"03",X"C1",X"03",X"01",X"03",X"01",X"55",X"55",
		X"55",X"55",X"00",X"01",X"3F",X"C1",X"30",X"C1",X"3F",X"C1",X"30",X"C1",X"3F",X"C1",X"55",X"55",
		X"55",X"55",X"00",X"01",X"3F",X"C1",X"30",X"C1",X"3F",X"C1",X"00",X"C1",X"00",X"C1",X"55",X"55",
		X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",
		X"BE",X"AA",X"AB",X"EA",X"AA",X"BE",X"AA",X"AB",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"EA",X"AA",X"BE",X"AA",X"AB",X"EA",X"AA",X"BE",X"AA",X"AB",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"EA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AB",X"AA",X"FE",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"BF",X"AF",X"EA",X"FA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AF",X"AB",X"FA",X"FE",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"BF",X"AE",X"EA",X"AE",X"AA",X"AE",X"AA",X"AE",X"AA",X"AE",X"AA",X"AE",X"AA",X"AE",X"AA",X"AE",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AE",X"AA",X"FE",
		X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"95",X"55",X"9F",X"FF",X"97",X"D7",X"A7",X"D9",X"A7",X"D9",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"6A",X"AA",X"DA",X"AA",X"F6",X"AA",X"F6",X"AA",
		X"BE",X"AA",X"AB",X"EA",X"AA",X"BE",X"AA",X"AB",X"AA",X"AA",X"A9",X"56",X"A9",X"FD",X"A9",X"BD",
		X"AA",X"AA",X"AA",X"AF",X"AB",X"FA",X"FE",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"BF",X"AA",X"EA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"96",X"AA",X"7D",X"AA",X"7D",X"AA",
		X"AA",X"AE",X"AA",X"AE",X"AA",X"AE",X"AA",X"AE",X"AA",X"AE",X"AA",X"AE",X"AA",X"AE",X"AA",X"AE",
		X"A7",X"D7",X"A7",X"FF",X"A7",X"D7",X"A7",X"D9",X"A7",X"D9",X"A7",X"D9",X"A7",X"D5",X"97",X"D7",
		X"D6",X"AA",X"59",X"65",X"DF",X"DF",X"FB",X"E7",X"F7",X"E7",X"F7",X"E7",X"F7",X"D7",X"D7",X"DF",
		X"AA",X"7D",X"A5",X"7D",X"5F",X"FF",X"7D",X"7D",X"7D",X"BD",X"7D",X"BD",X"7D",X"7D",X"7D",X"7D",
		X"AA",X"AA",X"59",X"59",X"F7",X"F7",X"D9",X"D9",X"F7",X"F7",X"F7",X"77",X"7F",X"7F",X"7D",X"7D",
		X"AA",X"AA",X"59",X"56",X"F7",X"FD",X"DF",X"AF",X"DF",X"5F",X"5F",X"FF",X"5F",X"A5",X"9F",X"5F",
		X"96",X"AA",X"5E",X"95",X"FD",X"7F",X"BD",X"FA",X"7D",X"F5",X"7D",X"BF",X"7D",X"6B",X"7D",X"D7",
		X"AA",X"AA",X"69",X"56",X"D7",X"FD",X"DF",X"AF",X"9F",X"5F",X"5F",X"FF",X"DF",X"A9",X"DF",X"5F",
		X"96",X"6E",X"5D",X"DE",X"FF",X"DE",X"7E",X"DE",X"7D",X"AE",X"7D",X"AE",X"7D",X"AE",X"7D",X"9E",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"EA",X"AA",
		X"9F",X"FF",X"95",X"55",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"65",X"F7",X"A9",X"59",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AF",X"AA",X"FA",
		X"DF",X"FF",X"65",X"55",X"AA",X"AF",X"AA",X"FA",X"AF",X"AA",X"FA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"7E",X"7D",X"96",X"96",X"FA",X"AA",X"AF",X"AA",X"AA",X"FE",X"AA",X"AB",X"AA",X"AA",X"AA",X"AA",
		X"97",X"FD",X"A5",X"56",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FA",X"AA",X"AF",X"EA",X"AA",X"BF",
		X"FF",X"FF",X"55",X"95",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"57",X"FD",X"65",X"56",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"76",X"55",X"9E",X"AA",X"AE",X"AA",X"AE",X"AA",X"AE",X"AA",X"AE",X"AA",X"AE",X"AA",X"AE",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AB",
		X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AF",X"AA",X"FA",X"AF",X"AA",X"BA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AF",X"AA",X"FA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FE",X"AA",X"AB",X"FA",X"AA",X"AF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"EA",X"AA",X"BF",X"AA",X"AA",X"FE",X"AA",X"AB",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AE",X"AA",X"AE",X"AA",X"AE",X"AA",X"AE",X"AA",X"AE",X"FA",X"AE",X"AF",X"EE",X"AA",X"BE",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"57",X"FF",X"57",X"FF",X"55",X"FF",X"55",X"7F",X"55",X"57",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FD",X"FF",X"FF",X"FF",X"FD",X"FF",X"FD",X"F5",X"F5",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"AA",X"55",X"FF",X"55",X"FF",X"55",X"FF",X"55",X"FF",X"55",X"FD",X"55",
		X"6A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"57",
		X"55",X"55",X"55",X"5F",X"55",X"FF",X"57",X"FF",X"5F",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"F5",X"FF",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"55",X"55",X"55",X"D5",X"55",X"FD",X"55",X"FF",X"55",X"FF",X"D5",X"FF",X"F5",X"FF",X"FD",
		X"55",X"55",X"AA",X"A5",X"FF",X"F5",X"FF",X"F5",X"FF",X"F5",X"FF",X"D5",X"FF",X"D5",X"FF",X"D6",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"AA",X"AA",
		X"6A",X"A8",X"1A",X"20",X"06",X"A0",X"06",X"20",X"06",X"A0",X"55",X"55",X"FF",X"FF",X"55",X"55",
		X"55",X"5F",X"55",X"7F",X"55",X"FF",X"57",X"FF",X"55",X"5F",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"57",X"FF",X"55",X"5F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"55",X"D5",X"55",
		X"57",X"FF",X"5F",X"FF",X"5F",X"FF",X"5F",X"FF",X"7F",X"FF",X"7F",X"FF",X"7F",X"FF",X"FF",X"FF",
		X"FF",X"57",X"FF",X"5F",X"FF",X"5F",X"FD",X"5F",X"FD",X"7F",X"FD",X"7F",X"F5",X"7F",X"F5",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",X"FF",X"F5",X"FF",X"F5",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"6A",X"AA",X"7F",X"FF",X"FF",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"A5",X"55",X"F5",X"55",X"F5",X"55",
		X"6A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"FF",X"FF",X"55",X"55",
		X"AA",X"AA",X"AA",X"AF",X"AA",X"FF",X"AB",X"FF",X"AF",X"FF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"FA",X"AA",X"FE",X"AA",X"FF",X"AA",X"FF",X"EA",X"FF",X"FA",X"FF",X"FE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",
		X"F5",X"AF",X"D5",X"AA",X"D6",X"AA",X"D6",X"AA",X"56",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",
		X"FF",X"F5",X"FF",X"D5",X"AF",X"D7",X"AA",X"D7",X"AA",X"A7",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AF",X"FF",X"AA",X"7D",
		X"F5",X"55",X"D5",X"55",X"D5",X"55",X"D6",X"AA",X"57",X"FF",X"5F",X"FF",X"5F",X"FF",X"7F",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"AA",X"55",X"FF",X"55",X"FF",X"55",X"FF",X"55",X"FD",X"55",
		X"2A",X"AA",X"2A",X"AA",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"02",X"AA",X"02",X"AA",X"02",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"0F",X"00",X"0F",X"00",X"15",X"00",X"15",
		X"AA",X"AF",X"AA",X"BF",X"AA",X"FF",X"AB",X"FF",X"AA",X"BF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AB",X"FF",X"AA",X"AF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"AA",X"EA",X"AA",
		X"FF",X"FD",X"FF",X"FD",X"FF",X"F5",X"FF",X"F5",X"FF",X"F5",X"FF",X"D5",X"FF",X"D6",X"FF",X"D6",
		X"6A",X"AA",X"6A",X"AA",X"6A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"2A",X"AA",
		X"AA",X"AD",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"7F",X"FF",X"7F",X"FF",X"AF",X"FF",X"AA",X"FF",X"AA",X"AB",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FD",X"55",X"FD",X"6A",X"F5",X"7F",X"F5",X"FF",X"F5",X"FF",X"D5",X"FF",X"D7",X"FF",X"D7",X"FF",
		X"55",X"55",X"AA",X"A5",X"FF",X"F5",X"FF",X"F5",X"FF",X"F5",X"FF",X"D5",X"FF",X"D5",X"FF",X"D5",
		X"AA",X"20",X"AA",X"20",X"AA",X"28",X"AA",X"08",X"AA",X"08",X"AA",X"0A",X"AA",X"02",X"AA",X"16",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"0A",X"FE",X"2A",X"BF",X"95",X"A5",
		X"00",X"0A",X"00",X"02",X"00",X"22",X"00",X"22",X"00",X"20",X"FA",X"20",X"BE",X"A0",X"67",X"E0",
		X"00",X"05",X"00",X"01",X"00",X"21",X"00",X"21",X"00",X"20",X"3C",X"20",X"7F",X"20",X"77",X"70",
		X"57",X"FF",X"5F",X"FF",X"5F",X"FF",X"5F",X"FF",X"7F",X"FF",X"7F",X"FF",X"7F",X"FF",X"FF",X"FF",
		X"FF",X"56",X"FF",X"5A",X"FF",X"5F",X"FD",X"5F",X"FD",X"7F",X"F5",X"7F",X"F5",X"7F",X"F5",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FA",X"AA",X"FF",X"AA",X"FF",X"FA",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"57",X"FF",X"5F",X"FF",X"5F",X"FF",X"5F",X"FF",X"7F",X"FF",X"7F",X"FF",X"7F",X"FF",X"FF",X"FF",
		X"FF",X"56",X"FF",X"56",X"FF",X"56",X"FD",X"56",X"FD",X"5A",X"FD",X"5A",X"F5",X"5A",X"F5",X"6A",
		X"AA",X"55",X"AA",X"A5",X"A5",X"65",X"A5",X"69",X"95",X"59",X"95",X"59",X"95",X"59",X"95",X"59",
		X"00",X"D5",X"01",X"FF",X"01",X"5F",X"0A",X"95",X"15",X"65",X"55",X"59",X"00",X"00",X"00",X"00",
		X"69",X"E0",X"5A",X"50",X"56",X"90",X"95",X"94",X"9D",X"94",X"7D",X"A4",X"FD",X"66",X"FD",X"66",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",
		X"F5",X"FF",X"D5",X"FF",X"D7",X"FF",X"D6",X"AA",X"57",X"FF",X"5F",X"FF",X"5F",X"FF",X"5F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"7F",X"FF",X"7F",X"FF",X"7F",X"FF",X"7F",X"FD",X"7F",
		X"FF",X"AA",X"FF",X"FA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FA",X"AA",X"FF",X"AA",X"FF",X"FA",X"FF",X"FE",X"FF",X"FE",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",
		X"F5",X"6A",X"D5",X"AA",X"D5",X"AA",X"D5",X"AA",X"56",X"AA",X"56",X"AA",X"56",X"AA",X"5A",X"AA",
		X"95",X"59",X"95",X"59",X"95",X"59",X"95",X"59",X"A5",X"69",X"A5",X"65",X"A9",X"A5",X"AA",X"55",
		X"5F",X"FF",X"5F",X"F7",X"5F",X"D5",X"52",X"01",X"62",X"01",X"02",X"81",X"00",X"80",X"00",X"80",
		X"FD",X"66",X"FD",X"66",X"FD",X"6F",X"7D",X"F7",X"FE",X"DF",X"7B",X"D3",X"6B",X"FF",X"BE",X"BF",
		X"00",X"AA",X"80",X"AA",X"80",X"AA",X"C0",X"2A",X"30",X"2A",X"30",X"2A",X"F0",X"0A",X"FC",X"0A",
		X"FD",X"7F",X"FD",X"6A",X"F5",X"7F",X"F5",X"FF",X"F5",X"FF",X"D5",X"FF",X"D7",X"FF",X"D7",X"FF",
		X"FF",X"FF",X"AA",X"A7",X"FF",X"F7",X"FF",X"F7",X"FF",X"F7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D6",
		X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"AA",X"AA",
		X"AA",X"BF",X"AA",X"F0",X"AA",X"FF",X"AB",X"C0",X"AB",X"FF",X"AF",X"00",X"AF",X"FF",X"7F",X"FF",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"AA",X"03",X"EA",X"FF",X"EA",X"00",X"FA",X"FF",X"FA",X"00",X"3E",X"FF",X"FE",X"FF",X"FF",
		X"AA",X"A0",X"AA",X"A0",X"AA",X"A0",X"AA",X"A8",X"AA",X"A8",X"AA",X"A8",X"AA",X"AA",X"AA",X"AA",
		X"00",X"A0",X"00",X"20",X"00",X"20",X"00",X"2A",X"00",X"20",X"00",X"20",X"00",X"20",X"00",X"20",
		X"AB",X"C3",X"00",X"00",X"00",X"00",X"AA",X"AA",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"AC",X"0A",X"00",X"02",X"00",X"02",X"AA",X"A2",X"80",X"82",X"80",X"82",X"80",X"82",X"80",X"82",
		X"57",X"FF",X"5F",X"FF",X"5F",X"FF",X"5F",X"FF",X"7F",X"FF",X"7F",X"FF",X"7F",X"FF",X"FF",X"FF",
		X"FF",X"57",X"FF",X"5F",X"FF",X"5F",X"FD",X"5F",X"FD",X"7F",X"FD",X"7F",X"F5",X"7F",X"F5",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",X"FF",X"F5",X"FF",X"F5",
		X"6A",X"AA",X"40",X"00",X"40",X"00",X"40",X"00",X"6A",X"AA",X"60",X"2A",X"7F",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"D0",X"00",X"D0",X"00",
		X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"A8",X"2A",X"08",X"20",X"08",X"20",
		X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"A0",X"0A",X"20",X"0A",X"08",X"0A",
		X"05",X"50",X"3D",X"55",X"FD",X"55",X"F5",X"5F",X"D5",X"57",X"55",X"57",X"55",X"57",X"5F",X"FF",
		X"00",X"20",X"80",X"20",X"80",X"20",X"80",X"20",X"A0",X"20",X"A0",X"20",X"A0",X"20",X"A8",X"20",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"8A",X"82",X"AA",X"8A",X"FF",X"AF",X"FF",X"BF",X"C0",
		X"80",X"82",X"80",X"82",X"80",X"82",X"A8",X"82",X"AA",X"82",X"FA",X"A2",X"FF",X"A2",X"0F",X"EB",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",
		X"F5",X"FF",X"D5",X"FF",X"D7",X"FF",X"D7",X"FF",X"57",X"FF",X"5F",X"FF",X"5F",X"FF",X"5F",X"FF",
		X"FF",X"F5",X"FF",X"D5",X"FF",X"D7",X"FF",X"D7",X"FF",X"57",X"FF",X"5F",X"FF",X"5F",X"FD",X"5F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",X"FF",X"F5",
		X"D0",X"00",X"50",X"00",X"52",X"AA",X"5A",X"AA",X"58",X"AA",X"5A",X"AA",X"6A",X"AA",X"6A",X"AA",
		X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"0A",X"00",X"0A",X"A8",X"0A",X"A8",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"AA",
		X"A5",X"69",X"65",X"5A",X"65",X"56",X"69",X"56",X"5D",X"55",X"5F",X"55",X"5F",X"D5",X"5F",X"F7",
		X"A8",X"20",X"A8",X"20",X"AA",X"20",X"AA",X"20",X"AA",X"20",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"BC",X"0A",X"FC",X"AA",X"F0",X"A0",X"F2",X"80",X"F2",X"80",X"F2",X"80",X"F0",X"A0",X"FC",X"AA",
		X"80",X"EF",X"A8",X"FF",X"A8",X"FF",X"2B",X"FF",X"2A",X"3F",X"2A",X"3A",X"A8",X"3A",X"A8",X"FA",
		X"FF",X"FD",X"FF",X"FD",X"FF",X"F5",X"FF",X"F5",X"FF",X"F5",X"FF",X"D5",X"FF",X"D7",X"FF",X"D7",
		X"7F",X"FF",X"7F",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FD",X"7F",X"FD",X"7F",X"F5",X"7F",X"F5",X"FF",X"F5",X"FF",X"D5",X"FF",X"D7",X"FF",X"D7",X"FF",
		X"FF",X"F5",X"FF",X"F5",X"FF",X"D5",X"FF",X"D5",X"FF",X"D6",X"FF",X"56",X"FF",X"56",X"FF",X"5A",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AB",
		X"BC",X"20",X"BF",X"20",X"AF",X"28",X"AA",X"08",X"AA",X"08",X"AA",X"0A",X"AA",X"02",X"AA",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"FF",X"00",X"CF",X"69",X"56",
		X"FF",X"FD",X"FF",X"FD",X"FF",X"F5",X"FF",X"F5",X"FF",X"F5",X"FF",X"D5",X"FF",X"D7",X"FF",X"D7",
		X"FF",X"57",X"FF",X"5F",X"FF",X"5F",X"FD",X"5F",X"FD",X"7F",X"FD",X"7F",X"F5",X"7F",X"F5",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",X"FF",X"F5",X"FF",X"F5",
		X"7F",X"FF",X"7F",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F5",X"FF",X"D5",X"FF",X"D7",X"FF",X"D7",X"FF",X"57",X"FF",X"5F",X"FF",X"5F",X"FF",X"5F",X"FF",
		X"FF",X"F5",X"FF",X"D5",X"FF",X"D7",X"FF",X"D7",X"FF",X"57",X"FF",X"5F",X"FF",X"5F",X"FD",X"5F",
		X"55",X"50",X"FF",X"55",X"FF",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"55",X"55",X"55",X"55",X"55",X"AA",X"AA",X"AA",X"AA",
		X"00",X"03",X"00",X"FF",X"0F",X"FF",X"3F",X"FF",X"FF",X"FF",X"7F",X"FF",X"7F",X"FF",X"5F",X"FF",
		X"7F",X"FF",X"57",X"FF",X"15",X"7F",X"05",X"57",X"01",X"55",X"00",X"15",X"00",X"0A",X"00",X"01",
		X"00",X"00",X"00",X"00",X"55",X"00",X"D5",X"50",X"F5",X"54",X"F5",X"55",X"F5",X"55",X"F5",X"55",
		X"F5",X"55",X"D5",X"55",X"55",X"54",X"55",X"50",X"55",X"40",X"54",X"00",X"80",X"00",X"80",X"00",
		X"02",X"C0",X"02",X"AA",X"0A",X"AA",X"0F",X"AA",X"3E",X"AA",X"7E",X"AA",X"6A",X"AA",X"5A",X"AA",
		X"5A",X"AA",X"56",X"AA",X"15",X"6A",X"05",X"56",X"01",X"55",X"02",X"D5",X"02",X"C0",X"02",X"C0",
		X"02",X"C0",X"02",X"C0",X"55",X"C0",X"55",X"50",X"95",X"54",X"A5",X"55",X"A5",X"55",X"A5",X"55",
		X"A5",X"55",X"95",X"55",X"55",X"54",X"55",X"50",X"55",X"40",X"56",X"C0",X"02",X"C0",X"02",X"C0",
		X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"57",X"55",X"5F",X"55",X"FF",X"55",X"FF",
		X"FD",X"5A",X"FD",X"5A",X"FD",X"6A",X"F5",X"6A",X"F5",X"6A",X"F5",X"AA",X"D5",X"AA",X"D5",X"AA",
		X"D6",X"AA",X"56",X"AA",X"56",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"6A",X"AA",X"6A",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",X"FF",X"F5",
		X"FF",X"F5",X"FF",X"F5",X"FF",X"D5",X"FF",X"D5",X"FF",X"D6",X"FF",X"56",X"FF",X"56",X"FF",X"5A",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"5F",X"55",X"F7",X"F5",X"FD",X"F5",X"FF",X"FD",
		X"57",X"FF",X"5F",X"FF",X"5F",X"FF",X"5F",X"FF",X"7F",X"FF",X"7F",X"FF",X"7F",X"FF",X"FF",X"FF",
		X"FF",X"57",X"FF",X"5F",X"FF",X"5F",X"FD",X"5F",X"FD",X"7F",X"FD",X"7F",X"F5",X"7F",X"F5",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",X"FF",X"F5",X"FF",X"F5",
		X"57",X"FF",X"5F",X"FF",X"5F",X"FF",X"5F",X"FF",X"7F",X"FF",X"7F",X"FF",X"7F",X"FF",X"FF",X"FF",
		X"FF",X"F5",X"FF",X"D5",X"FF",X"D7",X"FF",X"D7",X"FF",X"57",X"FF",X"5F",X"FF",X"5F",X"FD",X"5F",
		X"FD",X"7F",X"FD",X"7F",X"F5",X"7F",X"F5",X"FF",X"F5",X"FF",X"D5",X"FF",X"D7",X"FF",X"D7",X"FF",
		X"AA",X"AA",X"EA",X"AA",X"FA",X"AA",X"FE",X"AA",X"FA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FD",X"7F",X"FD",X"7F",X"F5",X"7F",X"F5",X"FF",X"F5",X"FF",X"D5",X"FF",X"D7",X"FF",X"D7",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",X"FF",X"F5",X"FF",X"F5",
		X"F5",X"FF",X"D5",X"FF",X"D7",X"FF",X"D7",X"FF",X"57",X"FF",X"5F",X"FF",X"5F",X"FF",X"5F",X"FF",
		X"7F",X"FF",X"7F",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FD",X"FF",X"FD",X"FF",X"F5",X"FF",X"F5",X"FF",X"F5",X"FF",X"D5",X"FF",X"D7",X"FF",X"D7",
		X"56",X"95",X"56",X"95",X"56",X"95",X"56",X"95",X"56",X"95",X"56",X"95",X"56",X"95",X"16",X"95",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",
		X"FF",X"F5",X"FF",X"D5",X"FF",X"D7",X"FF",X"D7",X"FF",X"57",X"FF",X"5F",X"FF",X"5F",X"FD",X"5F",
		X"FD",X"7F",X"FD",X"7F",X"F5",X"7F",X"F5",X"FF",X"F5",X"FF",X"D5",X"FF",X"D7",X"FF",X"D7",X"FF",
		X"7F",X"FF",X"7F",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FD",X"7F",X"FD",X"7F",X"F5",X"7F",X"F5",X"FF",X"F5",X"FF",X"D5",X"FF",X"D7",X"FF",X"D7",X"FF",
		X"FF",X"F5",X"FF",X"D5",X"FF",X"D7",X"FF",X"D7",X"FF",X"57",X"FF",X"5F",X"FF",X"5F",X"FD",X"5F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",X"FF",X"F5",X"FF",X"F5",
		X"FD",X"55",X"FD",X"6A",X"F5",X"7F",X"F5",X"FF",X"F5",X"FF",X"D5",X"FF",X"D7",X"FF",X"D7",X"FF",
		X"D5",X"55",X"D5",X"55",X"D6",X"AA",X"57",X"FF",X"5F",X"FF",X"5F",X"FF",X"5F",X"FF",X"7F",X"FF",
		X"7F",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"55",X"D5",X"55",X"F5",X"55",X"FD",X"55",X"F5",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"15",X"55",X"55",X"55",X"55",X"F5",X"55",X"75",X"55",X"75",X"55",X"D7",X"75",X"FF",X"FF",
		X"55",X"FD",X"55",X"7F",X"55",X"5F",X"7D",X"57",X"5D",X"55",X"5D",X"55",X"FD",X"55",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"55",X"55",X"FF",X"FD",X"FF",X"FF",X"FF",X"FF",X"55",X"5F",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"5F",
		X"55",X"5F",X"95",X"7F",X"A5",X"FF",X"97",X"FF",X"5F",X"FF",X"FF",X"FF",X"55",X"55",X"DA",X"AA",
		X"DA",X"AA",X"F5",X"6A",X"55",X"5A",X"55",X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"55",X"55",X"AF",X"FF",X"56",X"BF",X"01",X"6B",X"00",X"16",
		X"55",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"F5",X"55",X"56",X"AB",X"AA",X"BB",X"AA",X"BA",X"A9",X"AA",X"A5",X"55",X"55",X"55",X"55",
		X"55",X"FF",X"A9",X"55",X"6A",X"7A",X"6A",X"BB",X"5A",X"AB",X"56",X"AA",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"55",X"55",X"55",X"55",X"55",X"56",X"02",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"3D",X"03",X"FF",X"3F",X"FF",X"FF",X"FF",
		X"55",X"5A",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"D5",X"7D",X"5F",X"F5",X"FF",X"55",X"F5",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"FD",X"55",X"5F",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"5F",X"FF",X"DF",X"7F",X"FF",X"55",X"7F",X"FF",
		X"AA",X"9F",X"5A",X"9F",X"56",X"5F",X"56",X"75",X"55",X"FD",X"55",X"7F",X"55",X"57",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"57",X"55",X"7F",X"55",X"F5",X"56",X"7F",X"56",X"5F",X"5A",X"9F",
		X"55",X"FF",X"7F",X"FF",X"FF",X"55",X"DF",X"7F",X"5F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"55",X"7F",X"FF",X"7D",X"FF",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"56",X"F5",X"56",X"FF",X"56",X"FF",X"F5",X"57",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"95",X"55",X"A5",X"55",X"A5",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"BF",X"55",X"6F",X"FF",X"1B",X"FF",X"06",X"FF",X"01",X"BF",X"00",X"65",X"00",X"15",X"00",X"01",
		X"00",X"21",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"DF",X"00",X"FF",X"00",X"FC",X"00",X"F0",X"00",X"70",X"00",X"40",X"00",X"40",X"00",X"F0",X"03",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"05",X"55",X"FD",X"55",X"FF",X"FF",X"DF",X"F0",X"7F",X"F0",X"FF",X"C0",X"7F",X"C0",
		X"00",X"00",X"55",X"40",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"0F",X"C0",X"33",X"C0",X"0F",X"54",X"3F",X"50",X"0C",X"C0",X"00",X"C0",X"00",X"F0",X"00",
		X"50",X"00",X"FC",X"00",X"FC",X"00",X"FF",X"00",X"FF",X"00",X"7F",X"C0",X"55",X"54",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"0C",X"00",
		X"F0",X"00",X"FC",X"F0",X"FF",X"0F",X"F0",X"F0",X"3C",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
