library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_P2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_P2 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"F2",X"A5",X"8F",X"10",X"0D",X"A9",X"00",X"38",X"E5",X"D2",X"85",X"D2",X"A9",X"00",X"E5",X"D3",
		X"85",X"D3",X"60",X"BD",X"00",X"00",X"A9",X"00",X"85",X"D3",X"A5",X"8F",X"38",X"E9",X"07",X"AA",
		X"29",X"07",X"85",X"8F",X"8A",X"29",X"F8",X"0A",X"26",X"D3",X"0A",X"26",X"D3",X"85",X"D2",X"A5",
		X"8E",X"38",X"E9",X"06",X"AA",X"29",X"07",X"85",X"8E",X"8A",X"4A",X"4A",X"4A",X"18",X"65",X"D2",
		X"85",X"D2",X"A9",X"08",X"65",X"D3",X"85",X"D3",X"A4",X"8C",X"A2",X"00",X"A1",X"D2",X"29",X"3F",
		X"C9",X"1B",X"90",X"31",X"E9",X"1B",X"AA",X"BD",X"CF",X"3B",X"4A",X"4A",X"4A",X"4A",X"C5",X"8F",
		X"F0",X"02",X"B0",X"21",X"BD",X"CF",X"3B",X"29",X"0F",X"C5",X"8F",X"90",X"18",X"BD",X"AA",X"3B",
		X"4A",X"4A",X"4A",X"4A",X"C5",X"8E",X"F0",X"02",X"B0",X"0B",X"BD",X"AA",X"3B",X"29",X"0F",X"C5",
		X"8E",X"90",X"02",X"38",X"60",X"18",X"60",X"A5",X"80",X"29",X"F8",X"C9",X"C0",X"90",X"02",X"29",
		X"78",X"95",X"99",X"95",X"C4",X"A5",X"80",X"C9",X"D8",X"90",X"03",X"38",X"E9",X"28",X"C9",X"38",
		X"B0",X"03",X"18",X"69",X"38",X"95",X"B8",X"2A",X"2A",X"2A",X"2A",X"C9",X"C8",X"90",X"03",X"38",
		X"E9",X"38",X"C9",X"28",X"B0",X"03",X"18",X"69",X"28",X"95",X"B9",X"C9",X"70",X"B0",X"12",X"C9",
		X"28",X"90",X"0E",X"B5",X"B8",X"C9",X"7A",X"B0",X"08",X"C9",X"43",X"90",X"04",X"69",X"50",X"95",
		X"B8",X"B5",X"B9",X"C9",X"BC",X"B0",X"12",X"C9",X"79",X"90",X"0E",X"B5",X"B8",X"C9",X"C4",X"B0",
		X"08",X"C9",X"8B",X"90",X"04",X"E9",X"50",X"95",X"B8",X"86",X"D2",X"20",X"BA",X"32",X"A6",X"D2",
		X"B5",X"A0",X"29",X"F7",X"95",X"A0",X"29",X"06",X"F0",X"0A",X"A5",X"80",X"18",X"69",X"10",X"85",
		X"80",X"4C",X"87",X"30",X"60",X"B9",X"B8",X"00",X"95",X"90",X"B9",X"B9",X"00",X"95",X"98",X"60",
		X"A0",X"0A",X"A5",X"80",X"6A",X"90",X"02",X"A0",X"06",X"A2",X"06",X"20",X"05",X"31",X"B9",X"C4",
		X"00",X"95",X"99",X"88",X"88",X"A2",X"04",X"20",X"05",X"31",X"B9",X"C4",X"00",X"95",X"99",X"A2",
		X"02",X"A0",X"02",X"20",X"05",X"31",X"A2",X"00",X"A0",X"00",X"20",X"05",X"31",X"60",X"A2",X"0A",
		X"A9",X"F9",X"95",X"C4",X"A9",X"00",X"95",X"A0",X"CA",X"CA",X"E0",X"02",X"D0",X"F2",X"A2",X"02",
		X"20",X"87",X"30",X"A5",X"80",X"18",X"69",X"20",X"85",X"80",X"B5",X"A0",X"29",X"F1",X"95",X"A0",
		X"CA",X"CA",X"10",X"EC",X"A9",X"00",X"85",X"95",X"8D",X"80",X"08",X"8D",X"81",X"08",X"60",X"AD",
		X"82",X"08",X"48",X"20",X"40",X"3C",X"68",X"8D",X"82",X"08",X"20",X"BC",X"38",X"BD",X"62",X"3B",
		X"85",X"8E",X"BD",X"63",X"3B",X"85",X"8F",X"A0",X"1F",X"B1",X"8E",X"09",X"C0",X"99",X"00",X"08",
		X"88",X"10",X"F6",X"A2",X"75",X"8A",X"4A",X"A8",X"BD",X"74",X"3A",X"85",X"8D",X"CA",X"BD",X"74",
		X"3A",X"85",X"8C",X"B9",X"39",X"3A",X"A0",X"00",X"91",X"8C",X"CA",X"10",X"E8",X"A0",X"1D",X"A9",
		X"1B",X"BE",X"EA",X"3A",X"9D",X"00",X"08",X"BE",X"08",X"3B",X"9D",X"80",X"08",X"BE",X"26",X"3B",
		X"9D",X"00",X"0A",X"BE",X"44",X"3B",X"9D",X"00",X"0B",X"88",X"10",X"E5",X"60",X"A5",X"C5",X"4A",
		X"4A",X"4A",X"4A",X"09",X"70",X"8D",X"23",X"08",X"29",X"3F",X"09",X"80",X"8D",X"3B",X"08",X"AD",
		X"C5",X"00",X"29",X"0F",X"09",X"70",X"8D",X"24",X"08",X"29",X"3F",X"09",X"80",X"8D",X"3C",X"08",
		X"A5",X"C7",X"4A",X"4A",X"4A",X"4A",X"09",X"70",X"8D",X"39",X"08",X"29",X"3F",X"09",X"80",X"8D",
		X"25",X"08",X"A5",X"C7",X"29",X"0F",X"09",X"70",X"8D",X"3A",X"08",X"29",X"3F",X"09",X"80",X"8D",
		X"26",X"08",X"A5",X"82",X"20",X"7B",X"32",X"8E",X"68",X"0B",X"8D",X"67",X"0B",X"A5",X"83",X"20",
		X"7B",X"32",X"8E",X"65",X"0B",X"C9",X"F0",X"D0",X"02",X"A9",X"00",X"8D",X"64",X"0B",X"A9",X"EC",
		X"8D",X"66",X"0B",X"A2",X"04",X"A5",X"83",X"D0",X"2E",X"A5",X"82",X"F0",X"2A",X"C9",X"16",X"B0",
		X"26",X"A5",X"61",X"6A",X"B0",X"21",X"A5",X"63",X"29",X"02",X"D0",X"1B",X"A5",X"80",X"29",X"10",
		X"F0",X"15",X"BD",X"44",X"0B",X"29",X"3F",X"9D",X"44",X"0B",X"BD",X"64",X"0B",X"29",X"3F",X"9D",
		X"64",X"0B",X"CA",X"10",X"ED",X"30",X"13",X"BD",X"44",X"0B",X"09",X"C0",X"9D",X"44",X"0B",X"BD",
		X"64",X"0B",X"09",X"C0",X"9D",X"64",X"0B",X"CA",X"10",X"ED",X"60",X"A8",X"09",X"F0",X"AA",X"98",
		X"4A",X"4A",X"4A",X"4A",X"09",X"F0",X"60",X"A2",X"04",X"A5",X"80",X"29",X"18",X"F0",X"19",X"A9",
		X"9B",X"9D",X"C0",X"0A",X"A9",X"5B",X"9D",X"DB",X"0A",X"A9",X"5B",X"9D",X"BB",X"0A",X"A9",X"9B",
		X"9D",X"A0",X"0A",X"CA",X"10",X"E9",X"30",X"11",X"A9",X"1B",X"9D",X"C0",X"0A",X"9D",X"DB",X"0A",
		X"9D",X"A0",X"0A",X"9D",X"BB",X"0A",X"CA",X"10",X"F1",X"60",X"A2",X"0A",X"B5",X"A0",X"29",X"F9",
		X"95",X"A0",X"CA",X"CA",X"10",X"F6",X"A2",X"02",X"A0",X"00",X"B5",X"B8",X"38",X"F9",X"B8",X"00",
		X"10",X"06",X"C9",X"F8",X"B0",X"06",X"90",X"2A",X"C9",X"09",X"B0",X"26",X"B5",X"B9",X"38",X"F9",
		X"B9",X"00",X"10",X"06",X"C9",X"F8",X"B0",X"06",X"90",X"18",X"C9",X"09",X"B0",X"14",X"B5",X"A0",
		X"09",X"02",X"95",X"A0",X"B9",X"A0",X"00",X"09",X"02",X"99",X"A0",X"00",X"A5",X"CF",X"09",X"01",
		X"85",X"CF",X"A2",X"0A",X"20",X"2D",X"33",X"A2",X"06",X"20",X"2D",X"33",X"A0",X"02",X"A2",X"04",
		X"20",X"2D",X"33",X"A2",X"08",X"20",X"2D",X"33",X"A0",X"06",X"20",X"DA",X"33",X"A0",X"0A",X"20",
		X"DA",X"33",X"A2",X"04",X"20",X"DA",X"33",X"A0",X"06",X"20",X"DA",X"33",X"60",X"86",X"8D",X"84",
		X"8C",X"B5",X"C4",X"C9",X"C1",X"90",X"01",X"60",X"4A",X"4A",X"4A",X"A8",X"B9",X"25",X"34",X"18",
		X"75",X"B9",X"85",X"8E",X"B9",X"3D",X"34",X"18",X"75",X"B8",X"85",X"8F",X"20",X"B3",X"33",X"90",
		X"28",X"A6",X"8D",X"B5",X"C4",X"4A",X"4A",X"4A",X"A8",X"38",X"A9",X"00",X"F9",X"25",X"34",X"18",
		X"75",X"B9",X"85",X"8E",X"38",X"A9",X"00",X"F9",X"3D",X"34",X"18",X"75",X"B8",X"85",X"8F",X"20",
		X"B3",X"33",X"90",X"05",X"A6",X"8D",X"A4",X"8C",X"60",X"A6",X"8D",X"A4",X"8C",X"B5",X"A0",X"09",
		X"02",X"95",X"A0",X"B9",X"A0",X"00",X"09",X"04",X"99",X"A0",X"00",X"A9",X"3F",X"8D",X"80",X"08",
		X"A5",X"E4",X"D0",X"04",X"A5",X"CF",X"10",X"13",X"F8",X"A9",X"01",X"C0",X"02",X"18",X"F0",X"06",
		X"65",X"C7",X"85",X"C7",X"D0",X"04",X"65",X"C5",X"85",X"C5",X"D8",X"A9",X"20",X"99",X"A1",X"00",
		X"95",X"A1",X"60",X"A6",X"8C",X"B5",X"C4",X"4A",X"4A",X"4A",X"A8",X"B5",X"B8",X"38",X"E5",X"8F",
		X"B0",X"04",X"49",X"FF",X"69",X"01",X"D9",X"6D",X"34",X"B0",X"0E",X"B5",X"B9",X"38",X"E5",X"8E",
		X"B0",X"04",X"49",X"FF",X"69",X"01",X"D9",X"55",X"34",X"60",X"A9",X"C0",X"D5",X"C4",X"90",X"05",
		X"D9",X"C4",X"00",X"B0",X"01",X"60",X"B5",X"B8",X"38",X"F9",X"B8",X"00",X"10",X"06",X"C9",X"FC",
		X"B0",X"06",X"90",X"F1",X"C9",X"05",X"B0",X"ED",X"B5",X"B9",X"38",X"F9",X"B9",X"00",X"10",X"06",
		X"C9",X"FC",X"B0",X"06",X"90",X"DF",X"C9",X"05",X"B0",X"DB",X"B5",X"A0",X"09",X"04",X"95",X"A0",
		X"B9",X"A0",X"00",X"09",X"04",X"99",X"A0",X"00",X"A9",X"3F",X"8D",X"81",X"08",X"A9",X"20",X"99",
		X"A1",X"00",X"95",X"A1",X"60",X"FE",X"FE",X"FE",X"FE",X"FF",X"FF",X"00",X"01",X"01",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"01",X"01",X"00",X"FF",X"FF",X"FE",X"FE",X"FE",X"00",X"01",X"01",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"01",X"01",X"00",X"FF",X"FF",X"FE",X"FE",X"FE",X"FE",
		X"FE",X"FE",X"FE",X"FF",X"FF",X"08",X"08",X"08",X"07",X"05",X"05",X"03",X"05",X"06",X"06",X"07",
		X"08",X"08",X"08",X"07",X"06",X"06",X"05",X"03",X"04",X"05",X"07",X"08",X"08",X"03",X"04",X"05",
		X"07",X"08",X"08",X"08",X"08",X"08",X"07",X"05",X"04",X"03",X"05",X"06",X"06",X"07",X"08",X"08",
		X"08",X"07",X"06",X"06",X"05",X"1B",X"00",X"00",X"00",X"00",X"00",X"00",X"85",X"40",X"A5",X"E4",
		X"D0",X"07",X"A5",X"CF",X"30",X"03",X"4C",X"3A",X"35",X"A5",X"80",X"29",X"03",X"D0",X"08",X"A5",
		X"95",X"29",X"0F",X"F0",X"02",X"C6",X"95",X"AD",X"80",X"08",X"F0",X"09",X"A5",X"80",X"29",X"01",
		X"D0",X"03",X"CE",X"80",X"08",X"AD",X"81",X"08",X"F0",X"09",X"A5",X"80",X"29",X"00",X"D0",X"03",
		X"CE",X"81",X"08",X"AD",X"80",X"08",X"C9",X"10",X"B0",X"55",X"A0",X"00",X"A5",X"CF",X"10",X"2A",
		X"A5",X"E4",X"D0",X"26",X"A5",X"CF",X"6A",X"90",X"21",X"A5",X"AC",X"45",X"AD",X"45",X"AE",X"45",
		X"AF",X"45",X"80",X"45",X"84",X"45",X"85",X"45",X"86",X"45",X"87",X"45",X"C9",X"45",X"CB",X"2A",
		X"2A",X"2A",X"2A",X"C9",X"60",X"B0",X"02",X"69",X"60",X"A8",X"AD",X"81",X"08",X"0A",X"0A",X"84",
		X"8C",X"18",X"65",X"8C",X"90",X"02",X"A9",X"F0",X"A8",X"C9",X"10",X"B0",X"05",X"AD",X"80",X"08",
		X"D0",X"0D",X"A9",X"00",X"8D",X"80",X"08",X"85",X"6A",X"85",X"69",X"98",X"4C",X"28",X"35",X"85",
		X"6B",X"85",X"68",X"AD",X"80",X"08",X"0A",X"0A",X"29",X"F0",X"85",X"8C",X"A5",X"95",X"29",X"0F",
		X"05",X"8C",X"85",X"95",X"A5",X"CF",X"29",X"FE",X"85",X"CF",X"A2",X"02",X"A5",X"80",X"29",X"0F",
		X"D0",X"08",X"BD",X"40",X"08",X"F0",X"03",X"DE",X"40",X"08",X"A5",X"80",X"29",X"07",X"D0",X"08",
		X"BD",X"41",X"08",X"F0",X"03",X"DE",X"41",X"08",X"A5",X"80",X"29",X"01",X"D0",X"08",X"BD",X"61",
		X"08",X"F0",X"03",X"DE",X"61",X"08",X"B5",X"A0",X"29",X"0E",X"F0",X"0D",X"B5",X"90",X"95",X"D5",
		X"B5",X"98",X"95",X"D6",X"A9",X"3F",X"9D",X"61",X"08",X"CA",X"CA",X"10",X"BF",X"A5",X"CF",X"30",
		X"14",X"A5",X"80",X"D0",X"10",X"CE",X"82",X"08",X"10",X"0B",X"A9",X"1F",X"8D",X"82",X"08",X"20",
		X"3E",X"31",X"20",X"6F",X"31",X"A5",X"24",X"30",X"FC",X"60",X"A2",X"00",X"A5",X"CF",X"10",X"23",
		X"A5",X"C5",X"C0",X"02",X"F0",X"02",X"A5",X"C7",X"38",X"F8",X"F9",X"C5",X"00",X"D8",X"90",X"15",
		X"C9",X"02",X"90",X"10",X"C9",X"04",X"90",X"0B",X"C9",X"06",X"90",X"06",X"C9",X"08",X"90",X"01",
		X"E8",X"E8",X"E8",X"E8",X"E8",X"60",X"86",X"8C",X"A5",X"90",X"38",X"E5",X"92",X"B0",X"04",X"49",
		X"FF",X"69",X"01",X"C9",X"80",X"B0",X"0F",X"85",X"D1",X"A5",X"98",X"38",X"E5",X"9A",X"B0",X"04",
		X"49",X"FF",X"69",X"01",X"C9",X"80",X"B0",X"3B",X"18",X"65",X"D1",X"6A",X"85",X"D0",X"20",X"9A",
		X"35",X"A5",X"D0",X"C9",X"10",X"90",X"2F",X"C9",X"18",X"90",X"12",X"C9",X"20",X"90",X"14",X"C9",
		X"30",X"90",X"16",X"C9",X"40",X"90",X"18",X"E0",X"00",X"F0",X"1B",X"D0",X"16",X"E0",X"05",X"90",
		X"15",X"B0",X"10",X"E0",X"04",X"90",X"0F",X"B0",X"0A",X"E0",X"03",X"90",X"09",X"B0",X"04",X"E0",
		X"02",X"90",X"03",X"18",X"90",X"01",X"38",X"A6",X"8C",X"60",X"A2",X"02",X"B5",X"21",X"30",X"35",
		X"A5",X"E4",X"D0",X"04",X"A5",X"CF",X"30",X"2D",X"A5",X"63",X"29",X"02",X"D0",X"0A",X"A5",X"83",
		X"D0",X"15",X"A5",X"82",X"D0",X"11",X"F0",X"1D",X"B5",X"A0",X"30",X"19",X"A5",X"61",X"6A",X"B0",
		X"06",X"A5",X"97",X"F0",X"10",X"C6",X"97",X"A5",X"CF",X"30",X"04",X"09",X"C0",X"85",X"CF",X"B5",
		X"A0",X"09",X"80",X"95",X"A0",X"CA",X"CA",X"10",X"C3",X"A5",X"A0",X"10",X"08",X"A5",X"A2",X"10",
		X"04",X"A9",X"00",X"85",X"E4",X"A5",X"80",X"29",X"0F",X"F0",X"01",X"60",X"85",X"61",X"85",X"63",
		X"A9",X"00",X"85",X"8C",X"24",X"CF",X"10",X"04",X"A5",X"E4",X"F0",X"3C",X"A5",X"61",X"6A",X"B0",
		X"06",X"A5",X"63",X"29",X"02",X"D0",X"3C",X"A5",X"8C",X"09",X"C0",X"85",X"8C",X"A5",X"80",X"29",
		X"10",X"F0",X"20",X"A5",X"83",X"D0",X"04",X"A5",X"82",X"F0",X"1D",X"A5",X"8C",X"24",X"A0",X"10",
		X"04",X"09",X"04",X"D0",X"02",X"09",X"10",X"24",X"A2",X"10",X"04",X"09",X"08",X"D0",X"02",X"09",
		X"20",X"85",X"8C",X"A5",X"61",X"6A",X"90",X"03",X"4C",X"33",X"37",X"A5",X"8C",X"09",X"03",X"85",
		X"8C",X"D0",X"60",X"A5",X"97",X"D0",X"04",X"A5",X"CF",X"10",X"10",X"A5",X"8C",X"24",X"A0",X"30",
		X"02",X"09",X"40",X"24",X"A2",X"30",X"02",X"09",X"80",X"85",X"8C",X"A5",X"97",X"C9",X"02",X"B0",
		X"18",X"C9",X"01",X"D0",X"04",X"A5",X"CF",X"30",X"10",X"A5",X"8C",X"24",X"A0",X"30",X"02",X"09",
		X"01",X"24",X"A2",X"30",X"02",X"09",X"02",X"85",X"8C",X"A5",X"80",X"29",X"10",X"F0",X"24",X"A5",
		X"8C",X"24",X"A0",X"10",X"02",X"09",X"04",X"24",X"A2",X"10",X"02",X"09",X"08",X"85",X"8C",X"A5",
		X"97",X"F0",X"10",X"A5",X"8C",X"24",X"A0",X"30",X"02",X"09",X"10",X"24",X"A2",X"30",X"02",X"09",
		X"20",X"85",X"8C",X"A5",X"8C",X"29",X"C0",X"85",X"8D",X"20",X"BC",X"38",X"A5",X"61",X"6A",X"90",
		X"03",X"4C",X"DD",X"37",X"A5",X"63",X"29",X"02",X"D0",X"50",X"20",X"AB",X"38",X"BD",X"0C",X"3C",
		X"29",X"0F",X"09",X"30",X"05",X"8D",X"8D",X"CC",X"09",X"BD",X"0C",X"3C",X"4A",X"4A",X"4A",X"4A",
		X"09",X"30",X"05",X"8D",X"8D",X"CB",X"09",X"A9",X"2C",X"05",X"8D",X"8D",X"CA",X"09",X"BD",X"0D",
		X"3C",X"09",X"30",X"05",X"8D",X"8D",X"C9",X"09",X"A9",X"00",X"8D",X"CD",X"09",X"20",X"BC",X"38",
		X"BD",X"D3",X"38",X"85",X"8E",X"BD",X"D4",X"38",X"85",X"8F",X"A0",X"09",X"B1",X"8E",X"29",X"3F",
		X"05",X"8D",X"99",X"CE",X"09",X"88",X"10",X"F4",X"30",X"43",X"BD",X"F3",X"38",X"85",X"8E",X"BD",
		X"F4",X"38",X"85",X"8F",X"A0",X"12",X"98",X"DD",X"BD",X"39",X"D0",X"01",X"88",X"C9",X"11",X"D0",
		X"0E",X"E0",X"00",X"D0",X"0A",X"A5",X"97",X"C9",X"01",X"D0",X"04",X"99",X"C7",X"09",X"88",X"B1",
		X"8E",X"29",X"3F",X"05",X"8D",X"99",X"C7",X"09",X"88",X"10",X"DB",X"BC",X"BD",X"39",X"A9",X"04",
		X"C5",X"97",X"90",X"02",X"A5",X"97",X"09",X"30",X"05",X"8D",X"99",X"C7",X"09",X"A5",X"8C",X"0A",
		X"0A",X"29",X"C0",X"85",X"8D",X"10",X"02",X"85",X"62",X"24",X"8D",X"50",X"02",X"85",X"60",X"A5",
		X"A0",X"10",X"02",X"85",X"60",X"A5",X"A2",X"10",X"02",X"85",X"62",X"BD",X"DB",X"38",X"85",X"8E");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
