library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity loc_snd_rom is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of loc_snd_rom is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"21",X"00",X"20",X"06",X"00",X"C3",X"6A",X"01",X"32",X"00",X"50",X"3A",X"00",X"40",X"C9",X"FF",
		X"32",X"00",X"70",X"3A",X"00",X"60",X"C9",X"FF",X"78",X"CF",X"79",X"32",X"00",X"40",X"C9",X"FF",
		X"78",X"D7",X"79",X"32",X"00",X"60",X"C9",X"FF",X"87",X"85",X"6F",X"7C",X"CE",X"00",X"67",X"7E",
		X"23",X"66",X"6F",X"E9",X"FF",X"FF",X"FF",X"FF",X"D9",X"08",X"CD",X"40",X"00",X"08",X"D9",X"C9",
		X"3E",X"0E",X"CF",X"B7",X"28",X"0D",X"57",X"CB",X"BF",X"FE",X"2D",X"D0",X"CB",X"7A",X"28",X"29",
		X"C3",X"70",X"00",X"21",X"00",X"20",X"06",X"0C",X"AF",X"77",X"23",X"10",X"FC",X"C9",X"21",X"00",
		X"20",X"06",X"06",X"0E",X"07",X"BE",X"28",X"05",X"23",X"23",X"10",X"F9",X"41",X"79",X"90",X"C9",
		X"CD",X"5E",X"00",X"C8",X"AF",X"77",X"23",X"77",X"C9",X"32",X"17",X"20",X"CD",X"5E",X"00",X"28",
		X"04",X"23",X"36",X"00",X"C9",X"AF",X"CD",X"5E",X"00",X"28",X"08",X"3A",X"17",X"20",X"77",X"23",
		X"36",X"00",X"C9",X"CD",X"EF",X"00",X"CD",X"1A",X"01",X"B7",X"28",X"2D",X"3A",X"15",X"20",X"B7",
		X"28",X"1F",X"3A",X"16",X"20",X"21",X"06",X"20",X"CD",X"DE",X"00",X"CD",X"E6",X"00",X"57",X"3A",
		X"15",X"20",X"21",X"00",X"20",X"CD",X"DE",X"00",X"CD",X"E6",X"00",X"BA",X"F2",X"C1",X"00",X"18",
		X"08",X"3A",X"16",X"20",X"21",X"06",X"20",X"18",X"06",X"3A",X"15",X"20",X"21",X"00",X"20",X"B7",
		X"C8",X"3D",X"87",X"4F",X"06",X"00",X"09",X"3A",X"17",X"20",X"77",X"23",X"70",X"C9",X"3D",X"87",
		X"4F",X"06",X"00",X"09",X"7E",X"C9",X"21",X"F6",X"0C",X"06",X"00",X"4F",X"09",X"7E",X"C9",X"3A",
		X"00",X"20",X"CD",X"E6",X"00",X"32",X"11",X"20",X"3A",X"02",X"20",X"CD",X"E6",X"00",X"32",X"12",
		X"20",X"3A",X"04",X"20",X"CD",X"E6",X"00",X"32",X"13",X"20",X"3A",X"17",X"20",X"CD",X"E6",X"00",
		X"32",X"14",X"20",X"CD",X"45",X"01",X"32",X"15",X"20",X"C9",X"3A",X"06",X"20",X"CD",X"E6",X"00",
		X"32",X"11",X"20",X"3A",X"08",X"20",X"CD",X"E6",X"00",X"32",X"12",X"20",X"3A",X"0A",X"20",X"CD",
		X"E6",X"00",X"32",X"13",X"20",X"3A",X"17",X"20",X"CD",X"E6",X"00",X"32",X"14",X"20",X"CD",X"45",
		X"01",X"32",X"16",X"20",X"C9",X"21",X"11",X"20",X"3A",X"14",X"20",X"06",X"03",X"4F",X"7E",X"B9",
		X"F2",X"54",X"01",X"4F",X"23",X"10",X"F7",X"79",X"06",X"03",X"0E",X"01",X"21",X"11",X"20",X"BE",
		X"28",X"06",X"0C",X"23",X"10",X"F9",X"0E",X"00",X"79",X"C9",X"70",X"23",X"7C",X"FE",X"24",X"20",
		X"F9",X"F9",X"ED",X"56",X"21",X"00",X"30",X"22",X"0C",X"20",X"77",X"01",X"3F",X"07",X"DF",X"E7",
		X"32",X"0E",X"20",X"32",X"0F",X"20",X"CD",X"7C",X"02",X"CD",X"80",X"02",X"CD",X"84",X"02",X"CD",
		X"8A",X"02",X"CD",X"8E",X"02",X"CD",X"92",X"02",X"FB",X"3E",X"0F",X"CF",X"E6",X"40",X"20",X"F9",
		X"3E",X"0F",X"CF",X"E6",X"40",X"28",X"F9",X"F3",X"3E",X"01",X"32",X"10",X"20",X"3A",X"01",X"20",
		X"B7",X"3A",X"00",X"20",X"CA",X"BC",X"01",X"CD",X"64",X"02",X"18",X"03",X"CD",X"4A",X"02",X"FB",
		X"00",X"00",X"F3",X"3E",X"02",X"32",X"10",X"20",X"3A",X"03",X"20",X"B7",X"3A",X"02",X"20",X"CA",
		X"D7",X"01",X"CD",X"64",X"02",X"18",X"03",X"CD",X"4A",X"02",X"FB",X"00",X"00",X"F3",X"3E",X"03",
		X"32",X"10",X"20",X"3A",X"05",X"20",X"B7",X"3A",X"04",X"20",X"CA",X"F2",X"01",X"CD",X"64",X"02",
		X"18",X"03",X"CD",X"4A",X"02",X"FB",X"00",X"00",X"F3",X"3E",X"04",X"32",X"10",X"20",X"3A",X"07",
		X"20",X"B7",X"3A",X"06",X"20",X"CA",X"0D",X"02",X"CD",X"64",X"02",X"18",X"03",X"CD",X"4A",X"02",
		X"FB",X"00",X"00",X"F3",X"3E",X"05",X"32",X"10",X"20",X"3A",X"09",X"20",X"B7",X"3A",X"08",X"20",
		X"CA",X"28",X"02",X"CD",X"64",X"02",X"18",X"03",X"CD",X"4A",X"02",X"FB",X"00",X"00",X"F3",X"3E",
		X"06",X"32",X"10",X"20",X"3A",X"0B",X"20",X"B7",X"3A",X"0A",X"20",X"CA",X"44",X"02",X"CD",X"64",
		X"02",X"C3",X"98",X"01",X"CD",X"4A",X"02",X"C3",X"98",X"01",X"21",X"23",X"0D",X"EF",X"B7",X"20",
		X"1B",X"E5",X"21",X"01",X"20",X"3A",X"10",X"20",X"3D",X"87",X"D5",X"5F",X"16",X"00",X"19",X"D1",
		X"36",X"01",X"E1",X"C9",X"B7",X"C8",X"21",X"7D",X"0D",X"EF",X"B7",X"C8",X"21",X"00",X"20",X"3A",
		X"10",X"20",X"3D",X"4F",X"06",X"00",X"09",X"09",X"70",X"23",X"70",X"C9",X"06",X"08",X"18",X"06",
		X"06",X"09",X"18",X"02",X"06",X"0A",X"0E",X"00",X"DF",X"C9",X"06",X"08",X"18",X"06",X"06",X"09",
		X"18",X"02",X"06",X"0A",X"0E",X"00",X"E7",X"C9",X"3A",X"10",X"20",X"3D",X"21",X"A2",X"02",X"EF",
		X"AF",X"C9",X"AE",X"02",X"B7",X"02",X"C0",X"02",X"C9",X"02",X"D2",X"02",X"DB",X"02",X"CD",X"7C",
		X"02",X"0E",X"09",X"CD",X"E4",X"02",X"C9",X"CD",X"80",X"02",X"0E",X"12",X"CD",X"E4",X"02",X"C9",
		X"CD",X"84",X"02",X"0E",X"24",X"CD",X"E4",X"02",X"C9",X"CD",X"8A",X"02",X"0E",X"09",X"CD",X"F0",
		X"02",X"C9",X"CD",X"8E",X"02",X"0E",X"12",X"CD",X"F0",X"02",X"C9",X"CD",X"92",X"02",X"0E",X"24",
		X"CD",X"F0",X"02",X"C9",X"3A",X"0E",X"20",X"B1",X"32",X"0E",X"20",X"06",X"07",X"4F",X"DF",X"C9",
		X"3A",X"0F",X"20",X"B1",X"32",X"0F",X"20",X"06",X"07",X"4F",X"E7",X"C9",X"06",X"06",X"3A",X"10",
		X"20",X"FE",X"04",X"FA",X"08",X"03",X"E7",X"C9",X"DF",X"C9",X"3A",X"0E",X"20",X"A0",X"B1",X"32",
		X"0E",X"20",X"4F",X"06",X"07",X"DF",X"C9",X"3A",X"0F",X"20",X"A0",X"B1",X"32",X"0F",X"20",X"4F",
		X"06",X"07",X"E7",X"C9",X"3A",X"10",X"20",X"3D",X"21",X"2D",X"03",X"EF",X"C9",X"39",X"03",X"40",
		X"03",X"47",X"03",X"4E",X"03",X"55",X"03",X"5C",X"03",X"01",X"08",X"FE",X"CD",X"0A",X"03",X"C9",
		X"01",X"10",X"FD",X"CD",X"0A",X"03",X"C9",X"01",X"20",X"FB",X"CD",X"0A",X"03",X"C9",X"01",X"08",
		X"FE",X"CD",X"17",X"03",X"C9",X"01",X"10",X"FD",X"CD",X"17",X"03",X"C9",X"01",X"20",X"FB",X"CD",
		X"17",X"03",X"C9",X"3A",X"10",X"20",X"3D",X"21",X"6C",X"03",X"EF",X"C9",X"78",X"03",X"7F",X"03",
		X"86",X"03",X"8D",X"03",X"94",X"03",X"9B",X"03",X"01",X"01",X"F7",X"CD",X"0A",X"03",X"C9",X"01",
		X"02",X"EF",X"CD",X"0A",X"03",X"C9",X"01",X"04",X"DF",X"CD",X"0A",X"03",X"C9",X"01",X"01",X"F7",
		X"CD",X"17",X"03",X"C9",X"01",X"02",X"EF",X"CD",X"17",X"03",X"C9",X"01",X"04",X"DF",X"CD",X"17",
		X"03",X"C9",X"3A",X"10",X"20",X"3D",X"21",X"AB",X"03",X"EF",X"C9",X"B7",X"03",X"BE",X"03",X"C5",
		X"03",X"CC",X"03",X"D3",X"03",X"DA",X"03",X"01",X"00",X"F6",X"CD",X"0A",X"03",X"C9",X"01",X"00",
		X"ED",X"CD",X"0A",X"03",X"C9",X"01",X"00",X"DB",X"CD",X"0A",X"03",X"C9",X"01",X"00",X"F6",X"CD",
		X"17",X"03",X"C9",X"01",X"00",X"ED",X"CD",X"17",X"03",X"C9",X"01",X"00",X"DB",X"CD",X"17",X"03",
		X"C9",X"3A",X"10",X"20",X"FE",X"04",X"30",X"05",X"C6",X"07",X"47",X"DF",X"C9",X"C6",X"04",X"47",
		X"E7",X"C9",X"3A",X"10",X"20",X"FE",X"04",X"30",X"09",X"3D",X"87",X"47",X"4D",X"DF",X"4C",X"04",
		X"DF",X"C9",X"D6",X"04",X"87",X"47",X"4D",X"E7",X"4C",X"04",X"E7",X"C9",X"FE",X"04",X"D0",X"F5",
		X"CD",X"5C",X"04",X"F1",X"B7",X"20",X"02",X"77",X"C9",X"21",X"2C",X"04",X"87",X"87",X"4F",X"87",
		X"81",X"4F",X"06",X"00",X"09",X"3A",X"10",X"20",X"3D",X"EF",X"77",X"C9",X"7F",X"04",X"84",X"04",
		X"89",X"04",X"8E",X"04",X"93",X"04",X"98",X"04",X"9D",X"04",X"A2",X"04",X"A7",X"04",X"AC",X"04",
		X"B1",X"04",X"B6",X"04",X"BB",X"04",X"C0",X"04",X"C5",X"04",X"CA",X"04",X"CF",X"04",X"D4",X"04",
		X"D9",X"04",X"DE",X"04",X"E3",X"04",X"E8",X"04",X"ED",X"04",X"F2",X"04",X"21",X"2C",X"04",X"3A",
		X"10",X"20",X"3D",X"EF",X"C9",X"2A",X"0C",X"20",X"7B",X"A5",X"6F",X"7A",X"A4",X"67",X"22",X"0C",
		X"20",X"C9",X"2A",X"0C",X"20",X"7B",X"B5",X"6F",X"7A",X"B4",X"67",X"22",X"0C",X"20",X"C9",X"11",
		X"3F",X"FF",X"18",X"E1",X"11",X"FF",X"FC",X"18",X"DC",X"11",X"FF",X"F3",X"18",X"D7",X"11",X"FC",
		X"FF",X"18",X"D2",X"11",X"F3",X"FF",X"18",X"CD",X"11",X"CF",X"FF",X"18",X"C8",X"11",X"80",X"00",
		X"18",X"D0",X"11",X"00",X"02",X"18",X"CB",X"11",X"00",X"08",X"18",X"C6",X"11",X"02",X"00",X"18",
		X"C1",X"11",X"08",X"00",X"18",X"BC",X"11",X"20",X"00",X"18",X"B7",X"11",X"40",X"00",X"18",X"B2",
		X"11",X"00",X"01",X"18",X"AD",X"11",X"00",X"04",X"18",X"A8",X"11",X"01",X"00",X"18",X"A3",X"11",
		X"04",X"00",X"18",X"9E",X"11",X"10",X"00",X"18",X"99",X"11",X"C0",X"00",X"18",X"94",X"11",X"00",
		X"03",X"18",X"8F",X"11",X"00",X"0C",X"18",X"8A",X"11",X"03",X"00",X"18",X"85",X"11",X"0C",X"00",
		X"18",X"80",X"11",X"30",X"00",X"C3",X"72",X"04",X"DD",X"7E",X"00",X"32",X"37",X"20",X"FE",X"FF",
		X"C8",X"CD",X"06",X"05",X"AF",X"C9",X"DD",X"35",X"01",X"C0",X"3A",X"32",X"20",X"DD",X"77",X"01",
		X"DD",X"CB",X"00",X"46",X"C2",X"29",X"05",X"DD",X"7E",X"07",X"D6",X"01",X"FA",X"29",X"05",X"DD",
		X"77",X"07",X"32",X"34",X"20",X"4F",X"CD",X"E1",X"03",X"DD",X"35",X"00",X"C0",X"DD",X"6E",X"02",
		X"DD",X"66",X"03",X"7E",X"47",X"E6",X"1F",X"CA",X"C1",X"05",X"FE",X"1F",X"C2",X"D8",X"05",X"23",
		X"DD",X"75",X"02",X"DD",X"74",X"03",X"78",X"E6",X"E0",X"0F",X"0F",X"0F",X"0F",X"4F",X"06",X"00",
		X"21",X"59",X"05",X"09",X"5E",X"23",X"56",X"EB",X"E9",X"69",X"05",X"87",X"05",X"9D",X"05",X"B7",
		X"05",X"B7",X"05",X"B7",X"05",X"B7",X"05",X"B7",X"05",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"4E",
		X"CB",X"21",X"06",X"00",X"21",X"11",X"06",X"09",X"5E",X"23",X"56",X"ED",X"53",X"30",X"20",X"DD",
		X"73",X"04",X"DD",X"72",X"05",X"18",X"20",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"4E",X"06",X"00",
		X"21",X"A9",X"06",X"09",X"7E",X"32",X"32",X"20",X"DD",X"77",X"01",X"18",X"0A",X"DD",X"6E",X"02",
		X"DD",X"66",X"03",X"7E",X"DD",X"77",X"06",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"23",X"DD",X"75",
		X"02",X"DD",X"74",X"03",X"C3",X"2D",X"05",X"0E",X"00",X"CD",X"E1",X"03",X"DD",X"36",X"00",X"FF",
		X"C9",X"CD",X"C6",X"05",X"18",X"3D",X"78",X"E6",X"E0",X"07",X"07",X"07",X"47",X"3E",X"01",X"18",
		X"01",X"07",X"10",X"FD",X"DD",X"77",X"00",X"C9",X"C5",X"CD",X"C6",X"05",X"C1",X"78",X"E6",X"1F",
		X"3D",X"07",X"4F",X"06",X"00",X"DD",X"6E",X"04",X"DD",X"66",X"05",X"09",X"5E",X"23",X"56",X"EB",
		X"22",X"35",X"20",X"CD",X"F2",X"03",X"DD",X"4E",X"06",X"79",X"DD",X"77",X"07",X"32",X"34",X"20",
		X"CD",X"E1",X"03",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"23",X"DD",X"75",X"02",X"DD",X"74",X"03",
		X"C9",X"31",X"06",X"35",X"06",X"39",X"06",X"3D",X"06",X"41",X"06",X"45",X"06",X"49",X"06",X"4D",
		X"06",X"51",X"06",X"55",X"06",X"59",X"06",X"5D",X"06",X"61",X"06",X"65",X"06",X"69",X"06",X"6D",
		X"06",X"6B",X"08",X"F2",X"07",X"80",X"07",X"14",X"07",X"AE",X"06",X"4E",X"06",X"F3",X"05",X"9E",
		X"05",X"4E",X"05",X"01",X"05",X"B9",X"04",X"76",X"04",X"36",X"04",X"F9",X"03",X"C0",X"03",X"8A",
		X"03",X"57",X"03",X"27",X"03",X"FA",X"02",X"CF",X"02",X"A7",X"02",X"81",X"02",X"5D",X"02",X"3B",
		X"02",X"1B",X"02",X"FD",X"01",X"E0",X"01",X"C5",X"01",X"AC",X"01",X"94",X"01",X"7D",X"01",X"68",
		X"01",X"53",X"01",X"40",X"01",X"2E",X"01",X"1D",X"01",X"0D",X"01",X"FE",X"00",X"F0",X"00",X"E3",
		X"00",X"D6",X"00",X"CA",X"00",X"BE",X"00",X"B4",X"00",X"AA",X"00",X"A0",X"00",X"97",X"00",X"8F",
		X"00",X"87",X"00",X"7F",X"00",X"78",X"00",X"71",X"00",X"6B",X"00",X"65",X"00",X"5F",X"00",X"5A",
		X"00",X"55",X"00",X"50",X"00",X"4C",X"00",X"47",X"00",X"46",X"3F",X"38",X"31",X"2B",X"26",X"21",
		X"1C",X"18",X"15",X"12",X"0F",X"0D",X"0C",X"0B",X"0A",X"AF",X"32",X"37",X"20",X"21",X"EF",X"06",
		X"11",X"18",X"20",X"01",X"18",X"00",X"ED",X"B0",X"3A",X"33",X"20",X"07",X"4F",X"07",X"81",X"4F",
		X"06",X"00",X"21",X"07",X"0E",X"09",X"11",X"1A",X"20",X"CD",X"E5",X"06",X"11",X"22",X"20",X"CD",
		X"E5",X"06",X"11",X"2A",X"20",X"7E",X"12",X"CD",X"EC",X"06",X"7E",X"12",X"23",X"13",X"C9",X"01",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"1E",X"C3",X"4F",X"07",X"3E",X"1D",X"C3",X"4F",
		X"07",X"3E",X"1C",X"C3",X"4F",X"07",X"3E",X"1B",X"C3",X"4F",X"07",X"3E",X"1A",X"C3",X"4F",X"07",
		X"3E",X"19",X"C3",X"4F",X"07",X"3E",X"18",X"C3",X"4F",X"07",X"3E",X"17",X"C3",X"4F",X"07",X"3E",
		X"16",X"C3",X"4F",X"07",X"3E",X"15",X"C3",X"4F",X"07",X"3E",X"14",X"C3",X"4F",X"07",X"3E",X"13",
		X"C3",X"4F",X"07",X"3E",X"12",X"C3",X"4F",X"07",X"3E",X"11",X"C3",X"4F",X"07",X"3E",X"10",X"32",
		X"49",X"20",X"3E",X"FF",X"C9",X"3E",X"01",X"CD",X"0C",X"04",X"CD",X"24",X"03",X"21",X"00",X"05",
		X"22",X"3B",X"20",X"CD",X"F2",X"03",X"3E",X"0A",X"32",X"3A",X"20",X"4F",X"CD",X"E1",X"03",X"3E",
		X"40",X"32",X"38",X"20",X"3E",X"F0",X"32",X"39",X"20",X"AF",X"32",X"3D",X"20",X"C9",X"21",X"3D",
		X"20",X"35",X"7E",X"E6",X"01",X"20",X"36",X"21",X"38",X"20",X"35",X"7E",X"57",X"20",X"0A",X"36",
		X"40",X"21",X"3A",X"20",X"35",X"4E",X"CD",X"E1",X"03",X"2A",X"3B",X"20",X"CB",X"62",X"3A",X"39",
		X"20",X"06",X"FF",X"20",X"05",X"04",X"ED",X"44",X"CB",X"3F",X"4F",X"09",X"22",X"3B",X"20",X"CD",
		X"F2",X"03",X"7A",X"E6",X"1F",X"20",X"06",X"21",X"39",X"20",X"34",X"28",X"02",X"AF",X"C9",X"3D",
		X"C9",X"3E",X"01",X"CD",X"0C",X"04",X"CD",X"24",X"03",X"21",X"60",X"00",X"22",X"40",X"20",X"CD",
		X"F2",X"03",X"3E",X"0C",X"32",X"3F",X"20",X"4F",X"CD",X"E1",X"03",X"3E",X"20",X"32",X"3E",X"20",
		X"AF",X"C9",X"3A",X"3D",X"20",X"E6",X"01",X"C8",X"21",X"3E",X"20",X"35",X"28",X"17",X"7E",X"2A",
		X"40",X"20",X"FE",X"18",X"01",X"E8",X"FF",X"38",X"03",X"01",X"08",X"00",X"09",X"22",X"40",X"20",
		X"CD",X"F2",X"03",X"AF",X"C9",X"36",X"20",X"21",X"60",X"00",X"22",X"40",X"20",X"CD",X"F2",X"03",
		X"21",X"3F",X"20",X"35",X"28",X"06",X"4E",X"CD",X"E1",X"03",X"AF",X"C9",X"3D",X"C9",X"3E",X"01",
		X"CD",X"0C",X"04",X"CD",X"24",X"03",X"21",X"00",X"01",X"22",X"45",X"20",X"CD",X"F2",X"03",X"0E",
		X"0C",X"CD",X"E1",X"03",X"AF",X"32",X"42",X"20",X"32",X"43",X"20",X"C9",X"3A",X"3D",X"20",X"E6",
		X"01",X"C8",X"21",X"43",X"20",X"35",X"7E",X"28",X"21",X"57",X"FE",X"DC",X"28",X"2A",X"38",X"30",
		X"FE",X"E8",X"28",X"18",X"2A",X"45",X"20",X"3A",X"42",X"20",X"C6",X"9D",X"32",X"42",X"20",X"AA",
		X"AD",X"6F",X"22",X"45",X"20",X"CD",X"F2",X"03",X"AF",X"C9",X"3D",X"C9",X"3E",X"0F",X"32",X"44",
		X"20",X"4F",X"CD",X"E1",X"03",X"C3",X"54",X"08",X"3E",X"02",X"CD",X"0C",X"04",X"C3",X"54",X"08",
		X"E6",X"0F",X"20",X"D0",X"23",X"35",X"4E",X"CD",X"E1",X"03",X"C3",X"54",X"08",X"3E",X"02",X"CD",
		X"0C",X"04",X"CD",X"63",X"03",X"3E",X"01",X"32",X"47",X"20",X"3E",X"0B",X"32",X"4A",X"20",X"4F",
		X"CD",X"E1",X"03",X"AF",X"32",X"48",X"20",X"32",X"4B",X"20",X"C9",X"21",X"4B",X"20",X"35",X"7E",
		X"E6",X"01",X"C8",X"21",X"47",X"20",X"35",X"20",X"2D",X"3A",X"49",X"20",X"CB",X"3F",X"CB",X"3F",
		X"77",X"21",X"48",X"20",X"35",X"7E",X"E6",X"1F",X"16",X"0B",X"28",X"12",X"16",X"F2",X"FE",X"18",
		X"28",X"0C",X"3A",X"4A",X"20",X"57",X"CB",X"56",X"3E",X"FF",X"28",X"02",X"ED",X"44",X"82",X"32",
		X"4A",X"20",X"4F",X"CD",X"E1",X"03",X"3A",X"49",X"20",X"4F",X"CD",X"FC",X"02",X"AF",X"C9",X"3E",
		X"01",X"CD",X"0C",X"04",X"CD",X"24",X"03",X"0E",X"0A",X"CD",X"E1",X"03",X"21",X"00",X"00",X"CD",
		X"F2",X"03",X"3E",X"0F",X"32",X"4C",X"20",X"32",X"4D",X"20",X"AF",X"C9",X"21",X"4C",X"20",X"35",
		X"7E",X"E6",X"0F",X"21",X"4D",X"20",X"20",X"03",X"35",X"28",X"E1",X"BE",X"21",X"F0",X"00",X"38",
		X"02",X"2E",X"00",X"CD",X"F2",X"03",X"AF",X"C9",X"3E",X"03",X"CD",X"0C",X"04",X"CD",X"24",X"03",
		X"0E",X"0B",X"CD",X"E1",X"03",X"21",X"FF",X"02",X"7D",X"32",X"4E",X"20",X"32",X"4F",X"20",X"CD",
		X"F2",X"03",X"3E",X"08",X"32",X"50",X"20",X"AF",X"32",X"51",X"20",X"C9",X"21",X"51",X"20",X"35",
		X"7E",X"E6",X"03",X"20",X"19",X"21",X"50",X"20",X"3A",X"4F",X"20",X"57",X"B7",X"3A",X"4E",X"20",
		X"28",X"0E",X"96",X"38",X"0F",X"32",X"4E",X"20",X"6F",X"26",X"02",X"CD",X"F2",X"03",X"AF",X"C9",
		X"86",X"C3",X"63",X"09",X"7A",X"2F",X"32",X"4F",X"20",X"7E",X"3C",X"FE",X"3E",X"30",X"EF",X"77",
		X"AF",X"C9",X"3E",X"01",X"CD",X"0C",X"04",X"CD",X"24",X"03",X"0E",X"00",X"CD",X"E1",X"03",X"3E",
		X"03",X"21",X"56",X"20",X"77",X"2C",X"77",X"21",X"A0",X"00",X"22",X"54",X"20",X"3E",X"0A",X"32",
		X"53",X"20",X"3E",X"58",X"32",X"52",X"20",X"AF",X"C9",X"21",X"56",X"20",X"35",X"7E",X"2C",X"A6",
		X"20",X"28",X"21",X"52",X"20",X"35",X"28",X"DF",X"7E",X"57",X"E6",X"0F",X"20",X"09",X"21",X"53",
		X"20",X"35",X"35",X"4E",X"CD",X"E1",X"03",X"2A",X"54",X"20",X"CB",X"42",X"3E",X"0C",X"28",X"02",
		X"ED",X"44",X"85",X"6F",X"22",X"54",X"20",X"CD",X"F2",X"03",X"AF",X"C9",X"3E",X"01",X"32",X"57",
		X"20",X"3E",X"FF",X"C9",X"3E",X"01",X"CD",X"0C",X"04",X"CD",X"24",X"03",X"21",X"00",X"00",X"22",
		X"5C",X"20",X"CD",X"F2",X"03",X"3E",X"0F",X"32",X"5A",X"20",X"4F",X"CD",X"E1",X"03",X"3E",X"02",
		X"32",X"59",X"20",X"AF",X"32",X"58",X"20",X"32",X"5B",X"20",X"32",X"5E",X"20",X"C9",X"21",X"5E",
		X"20",X"35",X"7E",X"E6",X"01",X"C8",X"21",X"58",X"20",X"35",X"7E",X"57",X"20",X"04",X"2C",X"35",
		X"28",X"28",X"E6",X"1F",X"20",X"08",X"21",X"5A",X"20",X"35",X"4E",X"CD",X"E1",X"03",X"2A",X"5C",
		X"20",X"3A",X"5B",X"20",X"C6",X"C5",X"32",X"5B",X"20",X"AA",X"AD",X"6F",X"67",X"1F",X"38",X"02",
		X"26",X"01",X"22",X"5C",X"20",X"CD",X"F2",X"03",X"AF",X"C9",X"3D",X"C9",X"AF",X"CD",X"0C",X"04",
		X"CD",X"24",X"03",X"21",X"20",X"00",X"22",X"61",X"20",X"CD",X"F2",X"03",X"0E",X"09",X"CD",X"E1",
		X"03",X"3E",X"20",X"32",X"5F",X"20",X"3E",X"1E",X"32",X"60",X"20",X"AF",X"C9",X"3A",X"5E",X"20",
		X"E6",X"01",X"20",X"1C",X"21",X"5F",X"20",X"35",X"7E",X"28",X"17",X"2C",X"BE",X"38",X"11",X"0E",
		X"00",X"28",X"18",X"2A",X"61",X"20",X"01",X"0C",X"00",X"09",X"22",X"61",X"20",X"CD",X"F2",X"03",
		X"AF",X"C9",X"36",X"20",X"2C",X"35",X"35",X"28",X"07",X"0E",X"09",X"CD",X"E1",X"03",X"AF",X"C9",
		X"3D",X"C9",X"3E",X"01",X"CD",X"0C",X"04",X"CD",X"24",X"03",X"21",X"20",X"00",X"CD",X"F2",X"03",
		X"3E",X"08",X"32",X"64",X"20",X"4F",X"CD",X"E1",X"03",X"3E",X"01",X"32",X"65",X"20",X"AF",X"32",
		X"63",X"20",X"C9",X"21",X"63",X"20",X"35",X"7E",X"E6",X"3F",X"4F",X"28",X"19",X"FE",X"0C",X"20",
		X"18",X"21",X"65",X"20",X"3A",X"64",X"20",X"86",X"28",X"11",X"32",X"64",X"20",X"FE",X"0F",X"4F",
		X"20",X"04",X"7E",X"ED",X"44",X"77",X"CD",X"E1",X"03",X"AF",X"C9",X"3D",X"C9",X"3E",X"01",X"CD",
		X"0C",X"04",X"CD",X"24",X"03",X"21",X"00",X"01",X"CD",X"F2",X"03",X"3E",X"E0",X"32",X"67",X"20",
		X"32",X"69",X"20",X"32",X"66",X"20",X"3E",X"0C",X"32",X"68",X"20",X"4F",X"CD",X"E1",X"03",X"AF",
		X"C9",X"21",X"69",X"20",X"35",X"7E",X"E6",X"01",X"C8",X"21",X"67",X"20",X"35",X"7E",X"28",X"2B",
		X"57",X"E6",X"07",X"20",X"13",X"7A",X"FE",X"60",X"28",X"DC",X"FE",X"80",X"28",X"D8",X"FE",X"C0",
		X"28",X"D4",X"2C",X"35",X"4E",X"CD",X"E1",X"03",X"3A",X"66",X"20",X"C6",X"9B",X"32",X"66",X"20",
		X"AA",X"6F",X"17",X"9F",X"3C",X"67",X"CD",X"F2",X"03",X"AF",X"C9",X"3D",X"C9",X"3E",X"01",X"CD",
		X"0C",X"04",X"CD",X"24",X"03",X"21",X"50",X"01",X"CD",X"F2",X"03",X"3E",X"07",X"32",X"6C",X"20",
		X"4F",X"CD",X"E1",X"03",X"3E",X"80",X"32",X"6A",X"20",X"AF",X"32",X"6B",X"20",X"32",X"6D",X"20",
		X"C9",X"21",X"6D",X"20",X"35",X"7E",X"E6",X"01",X"C8",X"21",X"6B",X"20",X"35",X"7E",X"28",X"2F",
		X"FE",X"C0",X"38",X"17",X"E6",X"07",X"20",X"13",X"3A",X"6A",X"20",X"D6",X"0A",X"32",X"6A",X"20",
		X"3A",X"6C",X"20",X"3C",X"32",X"6C",X"20",X"4F",X"CD",X"E1",X"03",X"7E",X"E6",X"03",X"07",X"07",
		X"07",X"07",X"57",X"3A",X"6A",X"20",X"92",X"6F",X"26",X"01",X"CD",X"F2",X"03",X"AF",X"C9",X"3D",
		X"C9",X"3E",X"01",X"CD",X"0C",X"04",X"CD",X"24",X"03",X"21",X"38",X"01",X"CD",X"F2",X"03",X"3E",
		X"04",X"32",X"70",X"20",X"4F",X"CD",X"E1",X"03",X"3E",X"68",X"32",X"6E",X"20",X"AF",X"32",X"6F",
		X"20",X"32",X"71",X"20",X"C9",X"21",X"71",X"20",X"35",X"7E",X"E6",X"01",X"C8",X"21",X"6F",X"20",
		X"35",X"7E",X"28",X"2F",X"FE",X"C0",X"38",X"17",X"E6",X"07",X"20",X"13",X"3A",X"6E",X"20",X"D6",
		X"0A",X"32",X"6E",X"20",X"3A",X"70",X"20",X"3C",X"32",X"70",X"20",X"4F",X"CD",X"E1",X"03",X"7E",
		X"E6",X"03",X"07",X"07",X"07",X"07",X"57",X"3A",X"6E",X"20",X"92",X"6F",X"26",X"01",X"CD",X"F2",
		X"03",X"AF",X"C9",X"3D",X"C9",X"3E",X"00",X"CD",X"0C",X"04",X"CD",X"24",X"03",X"21",X"00",X"00",
		X"22",X"75",X"20",X"CD",X"F2",X"03",X"AF",X"32",X"74",X"20",X"4F",X"CD",X"E1",X"03",X"AF",X"32",
		X"72",X"20",X"32",X"73",X"20",X"32",X"77",X"20",X"C9",X"21",X"77",X"20",X"35",X"7E",X"E6",X"01",
		X"C8",X"21",X"73",X"20",X"35",X"7E",X"28",X"29",X"57",X"FE",X"D0",X"28",X"3A",X"38",X"51",X"FE",
		X"E0",X"28",X"20",X"38",X"25",X"2C",X"34",X"4E",X"CD",X"E1",X"03",X"2A",X"75",X"20",X"3A",X"72",
		X"20",X"C6",X"9D",X"32",X"72",X"20",X"AA",X"AD",X"6F",X"22",X"75",X"20",X"CD",X"F2",X"03",X"AF",
		X"C9",X"3D",X"C9",X"21",X"10",X"00",X"CD",X"F2",X"03",X"7A",X"E6",X"02",X"0E",X"00",X"28",X"02",
		X"0E",X"0F",X"CD",X"E1",X"03",X"AF",X"C9",X"3E",X"01",X"CD",X"0C",X"04",X"21",X"70",X"00",X"22",
		X"75",X"20",X"CD",X"F2",X"03",X"3E",X"05",X"32",X"74",X"20",X"4F",X"CD",X"E1",X"03",X"AF",X"C9",
		X"E6",X"3F",X"20",X"06",X"2C",X"35",X"4E",X"CD",X"E1",X"03",X"2A",X"75",X"20",X"CB",X"52",X"3E",
		X"01",X"28",X"02",X"ED",X"44",X"85",X"6F",X"CD",X"F2",X"03",X"AF",X"C9",X"3E",X"01",X"CD",X"0C",
		X"04",X"CD",X"24",X"03",X"21",X"00",X"01",X"CD",X"F2",X"03",X"3E",X"0F",X"32",X"79",X"20",X"4F",
		X"CD",X"E1",X"03",X"AF",X"32",X"78",X"20",X"C9",X"21",X"78",X"20",X"35",X"7E",X"E6",X"3F",X"FE",
		X"0C",X"0E",X"00",X"28",X"0A",X"B7",X"20",X"0A",X"21",X"79",X"20",X"35",X"28",X"06",X"4E",X"CD",
		X"E1",X"03",X"AF",X"C9",X"3D",X"C9",X"00",X"10",X"0F",X"0E",X"0D",X"0C",X"0B",X"0A",X"09",X"08",
		X"07",X"06",X"05",X"04",X"03",X"02",X"01",X"2C",X"2B",X"2A",X"29",X"28",X"27",X"26",X"25",X"24",
		X"23",X"22",X"21",X"20",X"1F",X"1E",X"1D",X"1C",X"1B",X"1A",X"19",X"18",X"17",X"16",X"15",X"14",
		X"13",X"12",X"11",X"98",X"02",X"55",X"07",X"C1",X"07",X"1E",X"08",X"8D",X"08",X"EF",X"08",X"28",
		X"09",X"82",X"09",X"DC",X"09",X"E4",X"09",X"4C",X"0A",X"A2",X"0A",X"ED",X"0A",X"4D",X"0B",X"B1",
		X"0B",X"15",X"0C",X"BC",X"0C",X"B9",X"0D",X"D0",X"0D",X"D0",X"0D",X"D0",X"0D",X"BE",X"0D",X"D0",
		X"0D",X"D0",X"0D",X"C3",X"0D",X"D0",X"0D",X"D0",X"0D",X"C8",X"0D",X"D0",X"0D",X"D0",X"0D",X"07",
		X"07",X"0C",X"07",X"11",X"07",X"16",X"07",X"1B",X"07",X"20",X"07",X"25",X"07",X"2A",X"07",X"2F",
		X"07",X"34",X"07",X"39",X"07",X"3E",X"07",X"43",X"07",X"48",X"07",X"4D",X"07",X"00",X"00",X"7E",
		X"07",X"E2",X"07",X"3C",X"08",X"AB",X"08",X"0C",X"09",X"4C",X"09",X"A9",X"09",X"00",X"00",X"0E",
		X"0A",X"6D",X"0A",X"C3",X"0A",X"11",X"0B",X"71",X"0B",X"D5",X"0B",X"39",X"0C",X"D8",X"0C",X"D9",
		X"0D",X"EE",X"0D",X"E0",X"0D",X"E7",X"0D",X"D9",X"0D",X"E0",X"0D",X"E7",X"0D",X"D9",X"0D",X"E0",
		X"0D",X"E7",X"0D",X"D9",X"0D",X"E0",X"0D",X"E7",X"0D",X"3E",X"00",X"C3",X"CA",X"0D",X"3E",X"01",
		X"C3",X"CA",X"0D",X"3E",X"02",X"C3",X"CA",X"0D",X"3E",X"03",X"32",X"33",X"20",X"CD",X"B9",X"06",
		X"AF",X"CD",X"0C",X"04",X"CD",X"24",X"03",X"AF",X"C9",X"DD",X"21",X"18",X"20",X"C3",X"F8",X"04",
		X"DD",X"21",X"20",X"20",X"C3",X"F8",X"04",X"DD",X"21",X"28",X"20",X"C3",X"F8",X"04",X"3A",X"37",
		X"20",X"FE",X"FF",X"C8",X"3A",X"34",X"20",X"4F",X"CD",X"E1",X"03",X"2A",X"35",X"20",X"CB",X"3C",
		X"CB",X"1D",X"CD",X"F2",X"03",X"AF",X"C9",X"1F",X"0E",X"3D",X"0E",X"72",X"0E",X"87",X"0E",X"B3",
		X"0E",X"DD",X"0E",X"F2",X"0E",X"21",X"0F",X"4E",X"0F",X"62",X"0F",X"AC",X"0F",X"CF",X"0F",X"1F",
		X"0F",X"5F",X"09",X"3F",X"0A",X"A6",X"80",X"81",X"86",X"60",X"61",X"86",X"60",X"68",X"3F",X"0B",
		X"CA",X"C6",X"3F",X"0C",X"AB",X"80",X"8B",X"A6",X"A8",X"3F",X"0D",X"EA",X"FF",X"1F",X"03",X"5F",
		X"07",X"80",X"76",X"76",X"80",X"76",X"76",X"80",X"76",X"76",X"80",X"76",X"76",X"80",X"76",X"76",
		X"80",X"76",X"76",X"80",X"76",X"76",X"80",X"76",X"76",X"80",X"77",X"77",X"80",X"77",X"77",X"80",
		X"77",X"77",X"80",X"77",X"77",X"80",X"76",X"76",X"80",X"76",X"76",X"80",X"76",X"76",X"80",X"76",
		X"76",X"FF",X"1F",X"03",X"5F",X"08",X"A6",X"A1",X"A6",X"A1",X"A6",X"A1",X"A6",X"AA",X"AB",X"A6",
		X"AB",X"AB",X"A6",X"A5",X"A3",X"A1",X"FF",X"1F",X"0E",X"3F",X"03",X"5F",X"09",X"38",X"38",X"38",
		X"38",X"78",X"3A",X"5A",X"38",X"3A",X"5A",X"3D",X"38",X"38",X"38",X"38",X"78",X"36",X"56",X"35",
		X"36",X"56",X"38",X"35",X"35",X"35",X"35",X"75",X"33",X"53",X"31",X"33",X"53",X"35",X"71",X"71",
		X"71",X"60",X"FF",X"1F",X"0E",X"5F",X"09",X"35",X"35",X"35",X"35",X"75",X"36",X"56",X"35",X"36",
		X"56",X"3A",X"35",X"35",X"35",X"35",X"75",X"33",X"53",X"31",X"33",X"53",X"35",X"31",X"31",X"31",
		X"31",X"71",X"30",X"50",X"2E",X"30",X"50",X"31",X"6E",X"6E",X"6E",X"60",X"FF",X"1F",X"08",X"5F",
		X"09",X"69",X"69",X"6A",X"6A",X"69",X"69",X"67",X"67",X"65",X"65",X"67",X"67",X"65",X"65",X"65",
		X"60",X"FF",X"1F",X"0E",X"3F",X"0B",X"5F",X"09",X"8E",X"6E",X"6E",X"8E",X"6E",X"6E",X"90",X"70",
		X"70",X"90",X"70",X"70",X"8E",X"6E",X"6E",X"8E",X"6E",X"6E",X"90",X"70",X"70",X"90",X"70",X"70",
		X"92",X"72",X"72",X"93",X"73",X"73",X"B2",X"B0",X"8E",X"6E",X"6E",X"6E",X"72",X"6E",X"72",X"AE",
		X"FF",X"1F",X"0E",X"5F",X"09",X"92",X"72",X"72",X"92",X"72",X"72",X"93",X"73",X"73",X"93",X"73",
		X"73",X"92",X"72",X"72",X"92",X"72",X"72",X"93",X"73",X"73",X"93",X"73",X"73",X"95",X"75",X"75",
		X"97",X"77",X"77",X"B5",X"B3",X"92",X"72",X"72",X"72",X"75",X"72",X"75",X"B2",X"FF",X"1F",X"02",
		X"5F",X"08",X"AE",X"A0",X"B0",X"A0",X"AE",X"A0",X"B0",X"A0",X"B2",X"B3",X"B2",X"B0",X"B2",X"B2",
		X"B2",X"FF",X"1F",X"0E",X"5F",X"09",X"3F",X"0B",X"69",X"66",X"82",X"82",X"62",X"64",X"66",X"67",
		X"89",X"89",X"89",X"86",X"3F",X"0A",X"8B",X"8B",X"8B",X"60",X"69",X"8B",X"60",X"69",X"6B",X"6D",
		X"6E",X"70",X"3F",X"09",X"92",X"1F",X"08",X"89",X"89",X"1F",X"0E",X"6E",X"69",X"3F",X"08",X"8E",
		X"1F",X"08",X"89",X"89",X"1F",X"0E",X"69",X"66",X"3F",X"07",X"89",X"1F",X"08",X"89",X"89",X"1F",
		X"0E",X"64",X"66",X"3F",X"06",X"82",X"1F",X"08",X"89",X"89",X"A0",X"FF",X"1F",X"08",X"5F",X"08",
		X"80",X"82",X"89",X"89",X"89",X"82",X"89",X"89",X"89",X"82",X"8B",X"8B",X"8B",X"82",X"8B",X"8B",
		X"8B",X"80",X"86",X"86",X"A0",X"86",X"86",X"A0",X"87",X"87",X"A0",X"86",X"86",X"A0",X"FF",X"1F",
		X"08",X"5F",X"08",X"A0",X"86",X"86",X"86",X"80",X"86",X"86",X"86",X"80",X"87",X"87",X"87",X"80",
		X"87",X"87",X"87",X"80",X"82",X"82",X"A0",X"82",X"82",X"A0",X"81",X"81",X"A0",X"82",X"82",X"A0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
