library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity swimmer_sound_rom is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of swimmer_sound_rom is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"31",X"00",X"24",X"F3",X"ED",X"56",X"C3",X"F5",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"08",X"D9",X"2A",X"D8",X"20",X"3A",X"00",X"30",
		X"77",X"23",X"22",X"D8",X"20",X"21",X"D0",X"20",X"CB",X"D6",X"D9",X"08",X"FB",X"ED",X"4D",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F5",X"D5",X"E5",X"21",X"D0",X"20",X"CB",X"C6",X"CB",X"4E",
		X"28",X"0F",X"ED",X"5B",X"D5",X"20",X"1B",X"ED",X"53",X"D5",X"20",X"7A",X"B3",X"20",X"02",X"CB",
		X"8E",X"E1",X"D1",X"F1",X"32",X"00",X"40",X"ED",X"45",X"F5",X"C5",X"3E",X"11",X"42",X"4B",X"11",
		X"00",X"00",X"EB",X"B7",X"ED",X"42",X"3F",X"38",X"02",X"09",X"B7",X"EB",X"ED",X"6A",X"EB",X"ED",
		X"6A",X"3D",X"20",X"EF",X"CB",X"3C",X"CB",X"1D",X"EB",X"C1",X"F1",X"C9",X"F5",X"C5",X"D5",X"4D",
		X"44",X"21",X"00",X"00",X"7B",X"B2",X"28",X"0D",X"CB",X"3A",X"CB",X"1B",X"30",X"01",X"09",X"CB",
		X"21",X"CB",X"10",X"18",X"EF",X"D1",X"C1",X"F1",X"C9",X"FD",X"E1",X"21",X"00",X"20",X"06",X"04",
		X"36",X"00",X"2C",X"20",X"FB",X"24",X"10",X"F8",X"32",X"00",X"40",X"21",X"00",X"23",X"22",X"D8",
		X"20",X"21",X"00",X"08",X"22",X"09",X"20",X"21",X"02",X"09",X"22",X"29",X"20",X"21",X"04",X"0A",
		X"22",X"49",X"20",X"FD",X"E9",X"CD",X"C9",X"00",X"FB",X"21",X"D0",X"20",X"CB",X"56",X"E5",X"C4",
		X"1A",X"01",X"E1",X"CB",X"46",X"28",X"F5",X"CB",X"86",X"CB",X"66",X"E5",X"C4",X"C7",X"01",X"E1",
		X"CB",X"76",X"C4",X"92",X"03",X"CD",X"15",X"07",X"18",X"DF",X"F3",X"ED",X"5B",X"D8",X"20",X"4B",
		X"1D",X"ED",X"53",X"D8",X"20",X"20",X"02",X"CB",X"96",X"11",X"00",X"23",X"1A",X"21",X"01",X"23",
		X"06",X"00",X"ED",X"B0",X"4F",X"E6",X"E0",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"5F",
		X"50",X"21",X"4B",X"01",X"19",X"5E",X"23",X"56",X"EB",X"FB",X"E9",X"5B",X"01",X"66",X"01",X"79",
		X"01",X"82",X"01",X"AD",X"01",X"89",X"01",X"9B",X"01",X"00",X"00",X"C9",X"79",X"E6",X"0F",X"C6",
		X"10",X"21",X"D0",X"20",X"18",X"59",X"79",X"E6",X"1F",X"6F",X"60",X"06",X"04",X"29",X"10",X"FD",
		X"22",X"D5",X"20",X"21",X"D0",X"20",X"CB",X"CE",X"C9",X"79",X"E6",X"1F",X"21",X"D4",X"20",X"86",
		X"77",X"C9",X"79",X"E6",X"1F",X"ED",X"44",X"18",X"F3",X"AF",X"32",X"00",X"20",X"32",X"20",X"20",
		X"32",X"40",X"20",X"21",X"D0",X"20",X"CB",X"A6",X"CB",X"AE",X"C9",X"AF",X"32",X"60",X"20",X"32",
		X"70",X"20",X"32",X"80",X"20",X"21",X"D0",X"20",X"CB",X"B6",X"CB",X"BE",X"C9",X"79",X"E6",X"0F",
		X"21",X"D0",X"20",X"CB",X"61",X"20",X"08",X"32",X"D1",X"20",X"CB",X"E6",X"CB",X"EE",X"C9",X"32",
		X"D2",X"20",X"CB",X"F6",X"CB",X"FE",X"C9",X"CB",X"4E",X"C0",X"CB",X"6E",X"C2",X"55",X"03",X"DD",
		X"21",X"00",X"20",X"DD",X"7E",X"00",X"87",X"C4",X"F1",X"01",X"DD",X"21",X"20",X"20",X"DD",X"7E",
		X"00",X"87",X"C4",X"F1",X"01",X"DD",X"21",X"40",X"20",X"DD",X"7E",X"00",X"87",X"C4",X"F1",X"01",
		X"C9",X"5F",X"16",X"00",X"21",X"FD",X"01",X"19",X"5E",X"23",X"56",X"EB",X"E9",X"00",X"00",X"05",
		X"02",X"42",X"02",X"56",X"02",X"DD",X"35",X"01",X"20",X"20",X"DD",X"7E",X"02",X"DD",X"35",X"02",
		X"B7",X"20",X"17",X"CD",X"6C",X"02",X"DD",X"5E",X"01",X"DD",X"56",X"02",X"DD",X"66",X"0F",X"2E",
		X"00",X"CD",X"89",X"00",X"DD",X"75",X"0D",X"DD",X"74",X"0E",X"DD",X"6E",X"0B",X"DD",X"66",X"0C",
		X"DD",X"5E",X"0D",X"DD",X"56",X"0E",X"B7",X"ED",X"52",X"DD",X"75",X"0B",X"DD",X"74",X"0C",X"C3",
		X"37",X"03",X"DD",X"35",X"01",X"20",X"0C",X"DD",X"7E",X"02",X"DD",X"35",X"02",X"B7",X"20",X"03",
		X"CD",X"6C",X"02",X"C3",X"37",X"03",X"DD",X"35",X"01",X"C0",X"DD",X"7E",X"02",X"DD",X"35",X"02",
		X"B7",X"C0",X"DD",X"7E",X"12",X"DD",X"77",X"00",X"CD",X"6C",X"02",X"C9",X"DD",X"6E",X"03",X"DD",
		X"66",X"04",X"7E",X"FE",X"FF",X"28",X"50",X"FE",X"64",X"CA",X"15",X"03",X"E5",X"87",X"5F",X"16",
		X"00",X"21",X"94",X"07",X"19",X"5E",X"23",X"56",X"E1",X"DD",X"73",X"07",X"DD",X"72",X"08",X"23",
		X"4E",X"23",X"DD",X"75",X"03",X"DD",X"74",X"04",X"26",X"00",X"69",X"3A",X"D4",X"20",X"47",X"3A",
		X"D3",X"20",X"80",X"54",X"CB",X"7F",X"20",X"16",X"3C",X"5F",X"CD",X"AC",X"00",X"DD",X"75",X"01",
		X"DD",X"74",X"02",X"DD",X"7E",X"0F",X"DD",X"77",X"0C",X"DD",X"36",X"0B",X"00",X"C9",X"ED",X"44",
		X"3C",X"5F",X"CD",X"89",X"00",X"18",X"E6",X"DD",X"6E",X"05",X"DD",X"66",X"06",X"7E",X"DD",X"77",
		X"00",X"B7",X"20",X"01",X"C9",X"FE",X"FF",X"20",X"1E",X"DD",X"36",X"0B",X"00",X"DD",X"36",X"0C",
		X"00",X"DD",X"36",X"07",X"00",X"DD",X"36",X"08",X"00",X"DD",X"6E",X"10",X"DD",X"66",X"11",X"DD",
		X"75",X"05",X"DD",X"74",X"06",X"18",X"D0",X"23",X"7E",X"32",X"D3",X"20",X"23",X"7E",X"DD",X"77",
		X"0F",X"23",X"5E",X"23",X"56",X"23",X"DD",X"73",X"03",X"DD",X"72",X"04",X"DD",X"75",X"05",X"DD",
		X"74",X"06",X"C3",X"6C",X"02",X"DD",X"36",X"07",X"00",X"DD",X"36",X"08",X"00",X"DD",X"36",X"0B",
		X"00",X"DD",X"36",X"0C",X"00",X"E5",X"CD",X"37",X"03",X"E1",X"DD",X"7E",X"00",X"DD",X"77",X"12",
		X"DD",X"36",X"00",X"03",X"C3",X"8F",X"02",X"06",X"00",X"DD",X"4E",X"09",X"21",X"A0",X"20",X"09",
		X"DD",X"5E",X"07",X"DD",X"56",X"08",X"73",X"23",X"72",X"DD",X"4E",X"0A",X"21",X"A0",X"20",X"09",
		X"DD",X"7E",X"0C",X"77",X"C9",X"CB",X"AE",X"AF",X"32",X"D4",X"20",X"3A",X"D1",X"20",X"87",X"5F",
		X"16",X"00",X"21",X"70",X"09",X"19",X"5E",X"23",X"56",X"EB",X"DD",X"21",X"00",X"20",X"CD",X"7C",
		X"03",X"DD",X"21",X"20",X"20",X"CD",X"7C",X"03",X"DD",X"21",X"40",X"20",X"5E",X"23",X"56",X"23",
		X"E5",X"DD",X"73",X"05",X"DD",X"72",X"06",X"DD",X"73",X"10",X"DD",X"72",X"11",X"CD",X"C7",X"02",
		X"E1",X"C9",X"CB",X"7E",X"28",X"03",X"CD",X"AF",X"03",X"DD",X"21",X"60",X"20",X"CD",X"BC",X"05",
		X"DD",X"21",X"70",X"20",X"CD",X"BC",X"05",X"DD",X"21",X"80",X"20",X"CD",X"BC",X"05",X"C9",X"CB",
		X"BE",X"3A",X"D2",X"20",X"87",X"5F",X"16",X"00",X"21",X"CC",X"03",X"19",X"5E",X"23",X"56",X"EB",
		X"5E",X"23",X"56",X"23",X"7E",X"4F",X"23",X"06",X"00",X"ED",X"B0",X"C9",X"0C",X"04",X"24",X"04",
		X"42",X"04",X"5A",X"04",X"8F",X"04",X"A1",X"04",X"C5",X"04",X"E3",X"04",X"FB",X"04",X"13",X"05",
		X"31",X"05",X"49",X"05",X"67",X"05",X"8B",X"05",X"98",X"05",X"A4",X"05",X"00",X"10",X"00",X"11",
		X"00",X"12",X"00",X"13",X"00",X"14",X"00",X"15",X"00",X"16",X"00",X"17",X"00",X"18",X"00",X"19",
		X"00",X"1A",X"00",X"1B",X"00",X"1C",X"00",X"1D",X"00",X"1E",X"00",X"1F",X"70",X"20",X"0F",X"01",
		X"00",X"F0",X"04",X"00",X"01",X"02",X"09",X"20",X"00",X"FE",X"FF",X"1D",X"04",X"10",X"00",X"00",
		X"00",X"10",X"00",X"00",X"70",X"20",X"0F",X"01",X"00",X"F0",X"00",X"39",X"00",X"02",X"09",X"10",
		X"02",X"FF",X"FF",X"35",X"04",X"30",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"FF",X"00",X"01",
		X"00",X"00",X"70",X"20",X"0F",X"01",X"00",X"FF",X"00",X"70",X"00",X"02",X"09",X"02",X"00",X"FF",
		X"00",X"53",X"04",X"80",X"00",X"FF",X"00",X"C0",X"FF",X"00",X"60",X"20",X"1F",X"01",X"00",X"00",
		X"00",X"30",X"00",X"00",X"08",X"40",X"00",X"00",X"00",X"7B",X"04",X"00",X"00",X"01",X"03",X"F0",
		X"00",X"40",X"00",X"02",X"09",X"40",X"FE",X"00",X"00",X"8E",X"04",X"01",X"00",X"F0",X"00",X"00",
		X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"FF",X"00",X"FF",X"FF",X"00",X"00",X"60",
		X"20",X"0F",X"01",X"00",X"FF",X"00",X"C0",X"00",X"00",X"08",X"10",X"FA",X"03",X"00",X"A0",X"04",
		X"00",X"60",X"20",X"0F",X"01",X"0F",X"F0",X"00",X"E0",X"00",X"00",X"08",X"10",X"00",X"00",X"00",
		X"B2",X"04",X"0F",X"0F",X"F0",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"80",X"00",
		X"FF",X"00",X"FF",X"03",X"00",X"60",X"20",X"0F",X"01",X"00",X"F0",X"00",X"3E",X"00",X"00",X"08",
		X"30",X"FC",X"01",X"00",X"D6",X"04",X"30",X"00",X"04",X"00",X"01",X"00",X"40",X"00",X"FF",X"00",
		X"01",X"00",X"00",X"60",X"20",X"0F",X"01",X"00",X"F0",X"00",X"F0",X"00",X"00",X"08",X"1F",X"F8",
		X"00",X"00",X"F4",X"04",X"10",X"00",X"F8",X"00",X"FC",X"FF",X"00",X"80",X"20",X"0F",X"01",X"00",
		X"00",X"00",X"29",X"00",X"04",X"0A",X"00",X"00",X"00",X"00",X"0C",X"05",X"FF",X"00",X"FA",X"00",
		X"00",X"00",X"00",X"80",X"20",X"0F",X"01",X"00",X"80",X"00",X"00",X"02",X"04",X"0A",X"00",X"00",
		X"00",X"00",X"24",X"05",X"3F",X"00",X"04",X"00",X"F8",X"FF",X"1F",X"00",X"FC",X"00",X"F0",X"FF",
		X"00",X"80",X"20",X"0F",X"01",X"00",X"00",X"00",X"3E",X"00",X"04",X"0A",X"00",X"00",X"00",X"00",
		X"42",X"05",X"7F",X"00",X"FE",X"00",X"00",X"00",X"00",X"70",X"20",X"0F",X"01",X"00",X"80",X"00",
		X"00",X"00",X"02",X"09",X"00",X"00",X"00",X"00",X"5A",X"05",X"3F",X"0F",X"02",X"00",X"00",X"00",
		X"3F",X"01",X"FE",X"00",X"00",X"00",X"00",X"80",X"20",X"0F",X"01",X"00",X"80",X"00",X"80",X"00",
		X"04",X"0A",X"12",X"07",X"FF",X"FF",X"78",X"05",X"0F",X"00",X"F0",X"00",X"FF",X"FF",X"20",X"00",
		X"07",X"00",X"FF",X"FF",X"08",X"00",X"E8",X"00",X"FF",X"FF",X"00",X"70",X"20",X"0F",X"03",X"00",
		X"F0",X"00",X"00",X"00",X"02",X"09",X"01",X"09",X"70",X"20",X"0F",X"02",X"00",X"00",X"00",X"00",
		X"00",X"02",X"09",X"0A",X"70",X"20",X"0F",X"01",X"00",X"00",X"00",X"29",X"00",X"02",X"09",X"00",
		X"00",X"00",X"00",X"B5",X"05",X"1F",X"00",X"FC",X"00",X"00",X"00",X"00",X"DD",X"7E",X"00",X"87",
		X"C8",X"5F",X"16",X"00",X"21",X"D1",X"05",X"19",X"5E",X"23",X"56",X"EB",X"11",X"A4",X"06",X"D5",
		X"E9",X"00",X"00",X"F3",X"05",X"68",X"06",X"84",X"06",X"F3",X"05",X"F3",X"05",X"F3",X"05",X"F3",
		X"05",X"F3",X"05",X"F3",X"05",X"F3",X"05",X"F3",X"05",X"F3",X"05",X"F3",X"05",X"F3",X"05",X"F3",
		X"05",X"F3",X"05",X"DD",X"E5",X"DD",X"7E",X"08",X"A7",X"20",X"46",X"DD",X"6E",X"0C",X"DD",X"66",
		X"0D",X"7E",X"A7",X"20",X"07",X"AF",X"DD",X"77",X"00",X"DD",X"E1",X"C9",X"DD",X"77",X"08",X"23",
		X"7E",X"23",X"DD",X"77",X"01",X"E6",X"10",X"28",X"12",X"DD",X"E5",X"D1",X"13",X"13",X"01",X"04",
		X"00",X"ED",X"B0",X"DD",X"75",X"0C",X"DD",X"74",X"0D",X"18",X"DE",X"7E",X"DD",X"77",X"09",X"23",
		X"23",X"7E",X"DD",X"77",X"0A",X"23",X"7E",X"DD",X"77",X"0B",X"23",X"DD",X"75",X"0C",X"DD",X"74",
		X"0D",X"DD",X"35",X"08",X"DD",X"CB",X"01",X"66",X"20",X"09",X"DD",X"7E",X"02",X"DD",X"86",X"09",
		X"DD",X"77",X"02",X"DD",X"5E",X"04",X"DD",X"56",X"05",X"DD",X"6E",X"0A",X"DD",X"66",X"0B",X"19",
		X"DD",X"75",X"04",X"DD",X"74",X"05",X"18",X"A1",X"DD",X"7E",X"02",X"D6",X"10",X"DD",X"77",X"02",
		X"D0",X"DD",X"35",X"08",X"20",X"05",X"DD",X"36",X"00",X"00",X"C9",X"ED",X"5F",X"F6",X"10",X"27",
		X"DD",X"77",X"04",X"C9",X"DD",X"35",X"08",X"C0",X"DD",X"35",X"09",X"20",X"05",X"DD",X"36",X"00",
		X"00",X"C9",X"DD",X"36",X"08",X"0F",X"DD",X"36",X"04",X"35",X"DD",X"CB",X"09",X"46",X"C8",X"DD",
		X"36",X"04",X"30",X"C9",X"DD",X"CB",X"01",X"46",X"28",X"09",X"DD",X"7E",X"01",X"E6",X"0E",X"87",
		X"32",X"C6",X"20",X"DD",X"CB",X"01",X"66",X"28",X"30",X"DD",X"CB",X"01",X"A6",X"DD",X"7E",X"01",
		X"21",X"BB",X"20",X"36",X"FF",X"E6",X"E0",X"07",X"07",X"07",X"5F",X"16",X"00",X"21",X"0D",X"07",
		X"19",X"7E",X"32",X"CD",X"20",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"22",X"CB",X"20",X"DD",X"5E",
		X"07",X"21",X"C0",X"20",X"19",X"36",X"10",X"18",X"13",X"DD",X"7E",X"02",X"E6",X"F0",X"0F",X"0F",
		X"0F",X"0F",X"DD",X"5E",X"07",X"16",X"00",X"21",X"C0",X"20",X"19",X"77",X"DD",X"5E",X"06",X"21",
		X"C0",X"20",X"19",X"DD",X"5E",X"04",X"DD",X"56",X"05",X"73",X"23",X"72",X"C9",X"00",X"04",X"08",
		X"09",X"0A",X"0B",X"0C",X"0D",X"0E",X"3F",X"3A",X"D0",X"20",X"CB",X"4F",X"20",X"18",X"3A",X"00",
		X"20",X"B7",X"28",X"02",X"CB",X"81",X"3A",X"20",X"20",X"B7",X"28",X"02",X"CB",X"89",X"3A",X"40",
		X"20",X"B7",X"28",X"02",X"CB",X"91",X"79",X"32",X"A7",X"20",X"21",X"90",X"20",X"11",X"A0",X"20",
		X"0E",X"01",X"CD",X"7E",X"07",X"0E",X"3F",X"AF",X"2A",X"60",X"20",X"BD",X"28",X"08",X"CB",X"81",
		X"CB",X"44",X"28",X"02",X"CB",X"99",X"2A",X"70",X"20",X"BD",X"28",X"08",X"CB",X"89",X"CB",X"44",
		X"28",X"02",X"CB",X"A1",X"2A",X"80",X"20",X"BD",X"28",X"08",X"CB",X"91",X"CB",X"44",X"28",X"02",
		X"CB",X"A9",X"79",X"32",X"C7",X"20",X"21",X"B0",X"20",X"11",X"C0",X"20",X"0E",X"81",X"06",X"0E",
		X"1A",X"BE",X"28",X"0B",X"77",X"3E",X"0E",X"90",X"ED",X"79",X"0D",X"7E",X"ED",X"79",X"0C",X"23",
		X"13",X"10",X"ED",X"C9",X"5D",X"0D",X"9C",X"0C",X"E7",X"0B",X"3C",X"0B",X"9B",X"0A",X"02",X"0A",
		X"73",X"09",X"EB",X"08",X"6B",X"08",X"F2",X"07",X"80",X"07",X"14",X"07",X"AE",X"06",X"4E",X"06",
		X"F4",X"05",X"9E",X"05",X"4D",X"05",X"01",X"05",X"B9",X"04",X"75",X"04",X"35",X"04",X"F9",X"03",
		X"C0",X"03",X"8A",X"03",X"57",X"03",X"27",X"03",X"FA",X"02",X"CF",X"02",X"A7",X"02",X"81",X"02",
		X"5D",X"02",X"3B",X"02",X"1B",X"02",X"FC",X"01",X"E0",X"01",X"C5",X"01",X"AC",X"01",X"94",X"01",
		X"7D",X"01",X"68",X"01",X"53",X"01",X"40",X"01",X"2E",X"01",X"1D",X"01",X"0D",X"01",X"FE",X"00",
		X"F0",X"00",X"E2",X"00",X"D6",X"00",X"CA",X"00",X"BE",X"00",X"B4",X"00",X"AA",X"00",X"A0",X"00",
		X"97",X"00",X"8F",X"00",X"87",X"00",X"7F",X"00",X"78",X"00",X"71",X"00",X"6B",X"00",X"65",X"00",
		X"5F",X"00",X"5A",X"00",X"55",X"00",X"50",X"00",X"4C",X"00",X"47",X"00",X"43",X"00",X"40",X"00",
		X"3C",X"00",X"39",X"00",X"35",X"00",X"32",X"00",X"30",X"00",X"2D",X"00",X"2A",X"00",X"28",X"00",
		X"26",X"00",X"24",X"00",X"22",X"00",X"20",X"00",X"1E",X"00",X"1C",X"00",X"1B",X"00",X"19",X"00",
		X"18",X"00",X"16",X"00",X"15",X"00",X"14",X"00",X"13",X"00",X"12",X"00",X"11",X"00",X"10",X"00",
		X"0F",X"00",X"0E",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"4D",X"6F",X"6E",X"69",X"74",X"65",X"72",X"20",X"62",X"79",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"4D",X"2E",X"49",X"73",X"68",X"69",X"7A",X"75",X"6B",X"61",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"53",X"6F",X"75",X"6E",X"64",X"20",X"62",X"79",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"4D",X"2E",X"49",X"73",X"68",X"69",X"7A",X"75",X"6B",X"61",X"20",X"20",
		X"20",X"20",X"20",X"20",X"52",X"2E",X"4B",X"61",X"77",X"61",X"6D",X"6F",X"74",X"6F",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"48",X"61",X"72",X"64",X"20",X"77",X"65",X"72",X"65",X"20",X"62",X"79",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"59",X"2E",X"4B",X"6F",X"74",X"6F",X"79",X"6F",X"72",X"69",X"20",X"20",
		X"20",X"20",X"20",X"20",X"4D",X"2E",X"59",X"6F",X"6E",X"65",X"64",X"61",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"44",X"65",X"62",X"75",X"67",X"20",X"62",X"79",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"4D",X"2E",X"54",X"73",X"75",X"6A",X"69",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"4D",X"75",X"73",X"69",X"63",X"20",X"62",X"79",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"52",X"2E",X"4E",X"69",X"73",X"68",X"69",X"7A",X"61",X"77",X"61",X"20",
		X"90",X"09",X"C2",X"09",X"94",X"0B",X"DD",X"0B",X"25",X"0C",X"9D",X"0C",X"BA",X"0C",X"D1",X"0C",
		X"61",X"0D",X"C4",X"0D",X"EA",X"0D",X"2E",X"0E",X"61",X"0C",X"8B",X"0E",X"8B",X"0E",X"8B",X"0E",
		X"96",X"09",X"9C",X"09",X"96",X"09",X"01",X"02",X"0F",X"A2",X"09",X"00",X"01",X"02",X"0F",X"AB",
		X"09",X"00",X"35",X"10",X"30",X"24",X"35",X"08",X"39",X"18",X"FF",X"64",X"10",X"0C",X"08",X"0C",
		X"04",X"0C",X"04",X"0C",X"08",X"0C",X"08",X"15",X"08",X"15",X"04",X"15",X"04",X"15",X"08",X"15",
		X"08",X"FF",X"C8",X"09",X"58",X"0A",X"13",X"0B",X"01",X"02",X"0F",X"00",X"0A",X"01",X"02",X"0F",
		X"00",X"0A",X"01",X"02",X"0F",X"0D",X"0A",X"01",X"02",X"0F",X"1A",X"0A",X"01",X"02",X"0F",X"00",
		X"0A",X"01",X"02",X"0F",X"00",X"0A",X"01",X"02",X"0F",X"0D",X"0A",X"01",X"02",X"0F",X"27",X"0A",
		X"01",X"02",X"0F",X"34",X"0A",X"01",X"02",X"0F",X"34",X"0A",X"01",X"02",X"0F",X"55",X"0A",X"FF",
		X"2B",X"08",X"2D",X"10",X"30",X"08",X"34",X"08",X"30",X"10",X"64",X"08",X"FF",X"32",X"08",X"32",
		X"10",X"32",X"08",X"32",X"08",X"32",X"10",X"30",X"08",X"FF",X"2F",X"08",X"2F",X"08",X"2D",X"08",
		X"2D",X"08",X"2B",X"10",X"64",X"10",X"FF",X"2F",X"08",X"2F",X"08",X"2D",X"08",X"2F",X"08",X"30",
		X"10",X"64",X"10",X"FF",X"34",X"08",X"34",X"08",X"30",X"08",X"30",X"08",X"2B",X"08",X"2B",X"08",
		X"30",X"08",X"34",X"08",X"32",X"08",X"32",X"08",X"2F",X"08",X"2F",X"08",X"2B",X"08",X"2B",X"08",
		X"2F",X"08",X"32",X"08",X"FF",X"30",X"40",X"FF",X"02",X"02",X"0C",X"90",X"0A",X"02",X"02",X"0C",
		X"90",X"0A",X"02",X"02",X"0C",X"9B",X"0A",X"02",X"02",X"0C",X"AC",X"0A",X"02",X"02",X"0C",X"90",
		X"0A",X"02",X"02",X"0C",X"90",X"0A",X"02",X"02",X"0C",X"9B",X"0A",X"02",X"02",X"0C",X"BF",X"0A",
		X"02",X"02",X"0C",X"CC",X"0A",X"02",X"02",X"0C",X"FD",X"0A",X"02",X"02",X"0C",X"06",X"0B",X"FF",
		X"48",X"20",X"64",X"08",X"43",X"08",X"45",X"08",X"47",X"08",X"FF",X"4A",X"08",X"48",X"08",X"47",
		X"08",X"45",X"08",X"4A",X"08",X"48",X"08",X"47",X"08",X"45",X"08",X"FF",X"47",X"08",X"45",X"08",
		X"47",X"08",X"45",X"08",X"43",X"04",X"64",X"04",X"43",X"08",X"45",X"08",X"47",X"08",X"FF",X"43",
		X"08",X"43",X"08",X"45",X"08",X"47",X"08",X"48",X"10",X"64",X"10",X"FF",X"4D",X"08",X"4C",X"08",
		X"4A",X"08",X"48",X"08",X"47",X"08",X"47",X"08",X"48",X"08",X"4A",X"08",X"4C",X"08",X"4A",X"08",
		X"48",X"08",X"47",X"08",X"45",X"08",X"45",X"08",X"47",X"08",X"48",X"08",X"4A",X"08",X"48",X"08",
		X"47",X"08",X"45",X"08",X"43",X"08",X"43",X"08",X"45",X"08",X"47",X"08",X"FF",X"48",X"10",X"43",
		X"10",X"48",X"10",X"64",X"10",X"FF",X"48",X"10",X"43",X"10",X"48",X"08",X"43",X"08",X"45",X"08",
		X"47",X"08",X"FF",X"01",X"02",X"0F",X"55",X"0B",X"01",X"02",X"0F",X"55",X"0B",X"01",X"02",X"0F",
		X"5E",X"0B",X"01",X"02",X"0F",X"67",X"0B",X"01",X"02",X"0F",X"55",X"0B",X"01",X"02",X"0F",X"55",
		X"0B",X"01",X"02",X"0F",X"5E",X"0B",X"01",X"02",X"0F",X"70",X"0B",X"01",X"02",X"0F",X"79",X"0B",
		X"01",X"02",X"0F",X"82",X"0B",X"01",X"02",X"0F",X"79",X"0B",X"01",X"02",X"0F",X"8B",X"0B",X"01",
		X"02",X"0F",X"55",X"0B",X"FF",X"18",X"10",X"13",X"10",X"18",X"10",X"64",X"10",X"FF",X"1A",X"10",
		X"15",X"10",X"1A",X"10",X"15",X"10",X"FF",X"13",X"10",X"15",X"10",X"13",X"10",X"64",X"10",X"FF",
		X"13",X"10",X"15",X"10",X"18",X"10",X"64",X"10",X"FF",X"1C",X"10",X"18",X"10",X"1C",X"10",X"18",
		X"10",X"FF",X"1A",X"10",X"17",X"10",X"1A",X"10",X"17",X"10",X"FF",X"1A",X"10",X"17",X"10",X"13",
		X"10",X"1A",X"10",X"FF",X"9A",X"0B",X"A0",X"0B",X"A6",X"0B",X"01",X"10",X"0F",X"AC",X"0B",X"FF",
		X"02",X"10",X"0C",X"C5",X"0B",X"FF",X"01",X"10",X"0F",X"D4",X"0B",X"FF",X"34",X"02",X"34",X"01",
		X"34",X"01",X"37",X"02",X"37",X"01",X"37",X"01",X"34",X"02",X"34",X"01",X"34",X"01",X"30",X"02",
		X"30",X"01",X"30",X"01",X"FF",X"18",X"02",X"1A",X"02",X"1C",X"02",X"1A",X"02",X"18",X"04",X"11",
		X"02",X"13",X"02",X"FF",X"58",X"04",X"58",X"04",X"58",X"04",X"58",X"04",X"FF",X"E3",X"0B",X"E9",
		X"0B",X"E3",X"0B",X"01",X"02",X"0F",X"EF",X"0B",X"00",X"01",X"02",X"0F",X"14",X"0C",X"00",X"24",
		X"08",X"24",X"08",X"24",X"08",X"28",X"10",X"24",X"08",X"28",X"08",X"28",X"08",X"28",X"08",X"2B",
		X"10",X"28",X"08",X"2B",X"08",X"2B",X"08",X"2F",X"10",X"23",X"08",X"28",X"08",X"28",X"08",X"28",
		X"08",X"2B",X"18",X"FF",X"64",X"18",X"0C",X"08",X"64",X"28",X"10",X"08",X"64",X"28",X"13",X"08",
		X"64",X"28",X"0C",X"08",X"FF",X"2B",X"0C",X"40",X"0C",X"2B",X"0C",X"02",X"02",X"0A",X"46",X"0C",
		X"02",X"02",X"0A",X"46",X"0C",X"02",X"02",X"0A",X"4F",X"0C",X"02",X"02",X"0A",X"4F",X"0C",X"FF",
		X"01",X"02",X"0F",X"58",X"0C",X"FF",X"35",X"08",X"34",X"08",X"35",X"08",X"34",X"08",X"FF",X"35",
		X"08",X"35",X"08",X"39",X"08",X"3B",X"08",X"FF",X"11",X"08",X"10",X"08",X"11",X"08",X"10",X"08",
		X"FF",X"67",X"0C",X"6D",X"0C",X"67",X"0C",X"01",X"02",X"0F",X"73",X"0C",X"00",X"01",X"02",X"0F",
		X"88",X"0C",X"00",X"30",X"08",X"30",X"08",X"30",X"08",X"34",X"08",X"34",X"08",X"34",X"08",X"35",
		X"08",X"35",X"08",X"35",X"08",X"37",X"18",X"FF",X"00",X"08",X"00",X"08",X"00",X"08",X"04",X"08",
		X"04",X"08",X"04",X"08",X"05",X"08",X"05",X"08",X"05",X"08",X"07",X"18",X"FF",X"A3",X"0C",X"A3",
		X"0C",X"A3",X"0C",X"01",X"04",X"0F",X"A9",X"0C",X"00",X"3C",X"04",X"39",X"04",X"3C",X"04",X"39",
		X"04",X"3C",X"04",X"39",X"04",X"3C",X"04",X"39",X"04",X"FF",X"C0",X"0C",X"C0",X"0C",X"C0",X"0C",
		X"01",X"04",X"0F",X"C6",X"0C",X"00",X"3C",X"08",X"37",X"08",X"34",X"08",X"37",X"08",X"30",X"08",
		X"FF",X"D7",X"0C",X"DD",X"0C",X"D7",X"0C",X"01",X"04",X"0F",X"E3",X"0C",X"00",X"01",X"04",X"0F",
		X"22",X"0D",X"00",X"35",X"08",X"30",X"08",X"35",X"08",X"30",X"08",X"35",X"08",X"30",X"08",X"35",
		X"08",X"30",X"08",X"32",X"08",X"2D",X"08",X"32",X"08",X"2D",X"08",X"32",X"08",X"2D",X"08",X"32",
		X"08",X"2D",X"08",X"34",X"08",X"30",X"08",X"34",X"08",X"30",X"08",X"34",X"08",X"30",X"08",X"34",
		X"08",X"30",X"08",X"35",X"08",X"30",X"08",X"35",X"08",X"30",X"08",X"35",X"07",X"30",X"08",X"35",
		X"10",X"FF",X"1D",X"08",X"18",X"08",X"1D",X"08",X"18",X"08",X"1D",X"08",X"18",X"08",X"1D",X"08",
		X"18",X"08",X"1A",X"08",X"15",X"08",X"1A",X"08",X"15",X"08",X"1A",X"08",X"15",X"08",X"1A",X"08",
		X"15",X"08",X"1C",X"08",X"18",X"08",X"1C",X"08",X"18",X"08",X"1C",X"08",X"18",X"08",X"1C",X"08",
		X"18",X"08",X"1D",X"08",X"18",X"08",X"1D",X"08",X"18",X"08",X"1D",X"07",X"18",X"08",X"1D",X"10",
		X"FF",X"67",X"0D",X"77",X"0D",X"67",X"0D",X"01",X"02",X"0F",X"7D",X"0D",X"01",X"02",X"0F",X"7D",
		X"0D",X"01",X"02",X"0F",X"88",X"0D",X"00",X"01",X"02",X"0F",X"A5",X"0D",X"00",X"30",X"08",X"2D",
		X"08",X"29",X"08",X"2D",X"08",X"2D",X"08",X"FF",X"30",X"08",X"30",X"08",X"32",X"08",X"32",X"08",
		X"30",X"08",X"30",X"08",X"2E",X"08",X"2E",X"08",X"2D",X"08",X"2D",X"08",X"2E",X"08",X"2E",X"08",
		X"30",X"10",X"30",X"08",X"FF",X"18",X"08",X"64",X"08",X"11",X"08",X"64",X"08",X"18",X"08",X"64",
		X"08",X"11",X"08",X"64",X"08",X"18",X"10",X"16",X"10",X"15",X"10",X"13",X"10",X"15",X"10",X"13",
		X"10",X"11",X"18",X"FF",X"CA",X"0D",X"D0",X"0D",X"CA",X"0D",X"01",X"02",X"0F",X"D6",X"0D",X"00",
		X"01",X"02",X"0F",X"DF",X"0D",X"00",X"30",X"10",X"2B",X"10",X"30",X"10",X"24",X"08",X"FF",X"0C",
		X"08",X"0C",X"08",X"13",X"08",X"10",X"08",X"0C",X"10",X"FF",X"F0",X"0D",X"F6",X"0D",X"F0",X"0D",
		X"01",X"02",X"0F",X"FC",X"0D",X"FF",X"01",X"02",X"0F",X"1D",X"0E",X"FF",X"43",X"04",X"40",X"04",
		X"43",X"04",X"40",X"04",X"43",X"04",X"40",X"04",X"43",X"04",X"40",X"04",X"41",X"04",X"3E",X"04",
		X"41",X"04",X"3E",X"04",X"41",X"04",X"3E",X"04",X"41",X"04",X"3E",X"04",X"FF",X"18",X"08",X"18",
		X"08",X"18",X"08",X"18",X"08",X"13",X"08",X"13",X"08",X"13",X"08",X"13",X"08",X"FF",X"34",X"0E",
		X"3A",X"0E",X"34",X"0E",X"01",X"02",X"0F",X"40",X"0E",X"FF",X"01",X"02",X"0F",X"61",X"0E",X"FF",
		X"39",X"10",X"39",X"10",X"39",X"10",X"35",X"10",X"30",X"10",X"30",X"10",X"35",X"10",X"39",X"10",
		X"37",X"10",X"37",X"10",X"37",X"10",X"34",X"10",X"30",X"10",X"30",X"10",X"34",X"10",X"37",X"10",
		X"FF",X"64",X"10",X"15",X"10",X"64",X"10",X"15",X"10",X"64",X"10",X"11",X"10",X"64",X"10",X"11",
		X"10",X"64",X"10",X"13",X"10",X"64",X"10",X"13",X"10",X"64",X"10",X"10",X"10",X"64",X"10",X"10",
		X"10",X"FF",X"03",X"00",X"00",X"88",X"0E",X"00",X"00",X"01",X"FF",X"91",X"0E",X"91",X"0E",X"91",
		X"0E",X"01",X"08",X"0F",X"D8",X"0E",X"01",X"08",X"0F",X"D8",X"0E",X"02",X"08",X"0F",X"20",X"0F",
		X"02",X"08",X"0F",X"27",X"0F",X"02",X"08",X"0F",X"20",X"0F",X"02",X"08",X"0F",X"27",X"0F",X"01",
		X"08",X"0F",X"2E",X"0F",X"02",X"08",X"0F",X"F5",X"0E",X"02",X"08",X"0F",X"F5",X"0E",X"01",X"08",
		X"0F",X"12",X"0F",X"01",X"08",X"0F",X"19",X"0F",X"01",X"08",X"0F",X"12",X"0F",X"01",X"08",X"0F",
		X"19",X"0F",X"02",X"08",X"0F",X"3B",X"0F",X"00",X"18",X"04",X"1D",X"04",X"1D",X"04",X"1F",X"04",
		X"1F",X"04",X"21",X"08",X"22",X"04",X"24",X"04",X"22",X"04",X"21",X"04",X"21",X"04",X"1F",X"04",
		X"1F",X"04",X"1D",X"08",X"FF",X"30",X"04",X"35",X"04",X"35",X"04",X"37",X"04",X"37",X"04",X"39",
		X"08",X"3A",X"04",X"3C",X"04",X"3A",X"04",X"39",X"04",X"39",X"04",X"37",X"04",X"37",X"04",X"35",
		X"08",X"FF",X"24",X"04",X"22",X"04",X"21",X"08",X"FF",X"22",X"04",X"21",X"04",X"1F",X"08",X"FF",
		X"3C",X"04",X"3A",X"04",X"39",X"08",X"FF",X"3A",X"04",X"39",X"04",X"37",X"08",X"FF",X"24",X"04",
		X"21",X"04",X"1D",X"04",X"1F",X"04",X"1F",X"04",X"1D",X"10",X"FF",X"3C",X"04",X"39",X"04",X"35",
		X"04",X"37",X"04",X"37",X"04",X"35",X"10",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"53",X"57",X"49",X"4D",X"4D",X"45",X"52",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"43",X"6F",X"70",X"79",X"20",X"72",X"69",X"67",X"68",X"74",X"20",X"31",X"39",X"38",X"32",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"54",X"45",X"48",X"4B",X"41",X"4E",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"49",X"6E",X"74",X"65",X"72",X"6E",X"61",X"74",X"69",X"6F",X"6E",X"61",X"6C",
		X"20",X"20",X"20",X"20",X"43",X"6F",X"72",X"70",X"72",X"61",X"74",X"69",X"6F",X"6E",X"20",X"20",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
