library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity cmd_prg_rom is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of cmd_prg_rom is
	type rom is array(0 to  20479) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"C3",X"A0",X"00",X"2A",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"31",X"39",X"38",X"33",X"2E",X"30",X"39",X"20",X"20",X"20",X"20",X"42",X"59",X"20",
		X"20",X"45",X"4C",X"53",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"2A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3A",X"00",X"A1",X"CB",X"5F",X"C0",X"3E",X"03",X"32",X"E4",X"9B",X"C9",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F5",X"AF",X"32",X"81",X"A1",X"C5",X"D5",X"E5",X"DD",X"E5",
		X"FD",X"E5",X"00",X"00",X"00",X"CD",X"5F",X"11",X"CD",X"C2",X"11",X"CD",X"88",X"0B",X"CD",X"56",
		X"0F",X"CD",X"BD",X"0F",X"CD",X"EC",X"0A",X"3E",X"00",X"32",X"80",X"A0",X"FD",X"E1",X"DD",X"E1",
		X"E1",X"D1",X"C1",X"3E",X"01",X"32",X"81",X"A1",X"F1",X"ED",X"45",X"00",X"00",X"00",X"00",X"00",
		X"AF",X"32",X"81",X"A1",X"3E",X"01",X"32",X"83",X"A1",X"ED",X"47",X"AF",X"21",X"00",X"98",X"11",
		X"01",X"98",X"01",X"FF",X"07",X"77",X"ED",X"B0",X"31",X"FF",X"9F",X"CD",X"01",X"07",X"CD",X"DB",
		X"0A",X"21",X"FF",X"FF",X"22",X"F0",X"9B",X"AF",X"32",X"E6",X"9B",X"AF",X"32",X"F2",X"9B",X"32",
		X"F3",X"9B",X"CD",X"02",X"06",X"3A",X"F4",X"9B",X"2F",X"47",X"3A",X"F5",X"9B",X"2F",X"A0",X"CA",
		X"C6",X"01",X"3A",X"F6",X"9B",X"A7",X"C2",X"0D",X"01",X"3A",X"F7",X"9B",X"47",X"3A",X"F8",X"9B",
		X"B0",X"CA",X"CB",X"00",X"2A",X"F0",X"9B",X"7C",X"B5",X"CA",X"3F",X"01",X"2B",X"22",X"F0",X"9B",
		X"CD",X"CE",X"01",X"CD",X"33",X"01",X"AF",X"32",X"F9",X"9B",X"C3",X"E2",X"00",X"CD",X"B5",X"10",
		X"CD",X"F2",X"12",X"CD",X"3F",X"02",X"AF",X"32",X"F9",X"9B",X"3A",X"F2",X"9B",X"A7",X"C2",X"6A",
		X"01",X"3A",X"F6",X"9B",X"FE",X"02",X"DA",X"13",X"01",X"3A",X"F3",X"9B",X"A7",X"C2",X"78",X"01",
		X"C3",X"13",X"01",X"3A",X"F9",X"9B",X"A7",X"C8",X"CD",X"B5",X"10",X"CD",X"F2",X"12",X"C9",X"3A",
		X"FA",X"9B",X"A7",X"C2",X"56",X"01",X"3E",X"FF",X"32",X"FA",X"9B",X"3A",X"F7",X"9B",X"47",X"3A",
		X"F8",X"9B",X"80",X"C3",X"C7",X"00",X"3A",X"F7",X"9B",X"47",X"3A",X"F8",X"9B",X"80",X"47",X"B8",
		X"CA",X"CB",X"00",X"AF",X"32",X"FA",X"9B",X"C3",X"C1",X"00",X"AF",X"32",X"E3",X"9B",X"3A",X"F6",
		X"9B",X"3D",X"32",X"F6",X"9B",X"C3",X"85",X"01",X"3E",X"FF",X"32",X"E3",X"9B",X"3A",X"F6",X"9B",
		X"D6",X"02",X"32",X"F6",X"9B",X"AF",X"32",X"F2",X"9B",X"32",X"F3",X"9B",X"CD",X"16",X"07",X"CD",
		X"3E",X"04",X"CD",X"3D",X"0C",X"3A",X"EE",X"9B",X"47",X"3A",X"EF",X"9B",X"A0",X"CA",X"8F",X"01",
		X"AF",X"32",X"FC",X"9B",X"32",X"6C",X"9C",X"32",X"83",X"A1",X"32",X"54",X"9A",X"3E",X"FF",X"32",
		X"FB",X"9B",X"CD",X"F2",X"12",X"AF",X"32",X"5D",X"9A",X"CD",X"2B",X"37",X"3A",X"6C",X"9C",X"A7",
		X"CA",X"B9",X"01",X"C3",X"C1",X"00",X"3E",X"FF",X"32",X"F6",X"9B",X"C3",X"1A",X"01",X"3A",X"F6",
		X"9B",X"A7",X"C0",X"CD",X"36",X"04",X"21",X"C2",X"3B",X"CD",X"84",X"10",X"3A",X"F7",X"9B",X"A7",
		X"C2",X"EB",X"01",X"3A",X"F8",X"9B",X"A7",X"C2",X"28",X"02",X"C9",X"3A",X"F4",X"9B",X"4F",X"06",
		X"00",X"CB",X"21",X"DD",X"21",X"77",X"3C",X"DD",X"09",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"11",
		X"E3",X"01",X"D5",X"ED",X"5B",X"59",X"9A",X"01",X"FF",X"03",X"7B",X"A1",X"4F",X"7A",X"A0",X"B1",
		X"CC",X"84",X"10",X"E5",X"EB",X"11",X"00",X"02",X"19",X"EB",X"E1",X"01",X"FF",X"03",X"7B",X"A1",
		X"4F",X"7A",X"A0",X"B1",X"CA",X"DD",X"0F",X"C9",X"3A",X"F5",X"9B",X"4F",X"06",X"00",X"CB",X"21",
		X"DD",X"21",X"26",X"3D",X"DD",X"09",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"C3",X"03",X"02",X"CD",
		X"36",X"04",X"21",X"85",X"3C",X"CD",X"DD",X"0F",X"21",X"D6",X"3B",X"CD",X"DD",X"0F",X"21",X"C2",
		X"3B",X"CD",X"DD",X"0F",X"3A",X"F6",X"9B",X"FE",X"02",X"DA",X"65",X"02",X"21",X"B0",X"3B",X"22",
		X"85",X"9C",X"C3",X"6B",X"02",X"21",X"9F",X"3B",X"22",X"85",X"9C",X"2A",X"59",X"9A",X"01",X"FF",
		X"03",X"79",X"A5",X"4F",X"78",X"A4",X"B1",X"CA",X"8B",X"02",X"01",X"00",X"02",X"09",X"01",X"FF",
		X"03",X"79",X"A5",X"4F",X"78",X"A4",X"B1",X"CA",X"98",X"02",X"C9",X"21",X"8A",X"3B",X"CD",X"84",
		X"10",X"2A",X"85",X"9C",X"CD",X"84",X"10",X"C9",X"2A",X"85",X"9C",X"CD",X"DD",X"0F",X"C9",X"3A",
		X"F4",X"9B",X"FE",X"00",X"CA",X"E7",X"02",X"FE",X"01",X"CA",X"2F",X"03",X"FE",X"02",X"CA",X"5F",
		X"03",X"FE",X"03",X"CA",X"77",X"03",X"FE",X"04",X"CA",X"FF",X"02",X"FE",X"05",X"CA",X"17",X"03",
		X"C3",X"47",X"03",X"3A",X"F5",X"9B",X"FE",X"00",X"CA",X"8F",X"03",X"FE",X"01",X"CA",X"D6",X"03",
		X"FE",X"02",X"CA",X"06",X"04",X"FE",X"03",X"CA",X"1E",X"04",X"FE",X"04",X"CA",X"A6",X"03",X"FE",
		X"05",X"CA",X"BE",X"03",X"C3",X"EE",X"03",X"3A",X"F7",X"9B",X"C6",X"01",X"32",X"F7",X"9B",X"FE",
		X"01",X"C0",X"3A",X"F6",X"9B",X"C6",X"01",X"32",X"F6",X"9B",X"AF",X"32",X"F7",X"9B",X"C9",X"3A",
		X"F7",X"9B",X"C6",X"01",X"32",X"F7",X"9B",X"FE",X"01",X"C0",X"3A",X"F6",X"9B",X"C6",X"02",X"32",
		X"F6",X"9B",X"AF",X"32",X"F7",X"9B",X"C9",X"3A",X"F7",X"9B",X"C6",X"01",X"32",X"F7",X"9B",X"FE",
		X"01",X"C0",X"3A",X"F6",X"9B",X"C6",X"03",X"32",X"F6",X"9B",X"AF",X"32",X"F7",X"9B",X"C9",X"3A",
		X"F7",X"9B",X"C6",X"01",X"32",X"F7",X"9B",X"FE",X"02",X"C0",X"3A",X"F6",X"9B",X"C6",X"01",X"32",
		X"F6",X"9B",X"AF",X"32",X"F7",X"9B",X"C9",X"3A",X"F7",X"9B",X"C6",X"01",X"32",X"F7",X"9B",X"FE",
		X"02",X"C0",X"3A",X"F6",X"9B",X"C6",X"03",X"32",X"F6",X"9B",X"AF",X"32",X"F7",X"9B",X"C9",X"3A",
		X"F7",X"9B",X"C6",X"01",X"32",X"F7",X"9B",X"FE",X"03",X"C0",X"3A",X"F6",X"9B",X"C6",X"01",X"32",
		X"F6",X"9B",X"AF",X"32",X"F7",X"9B",X"C9",X"3A",X"F7",X"9B",X"C6",X"01",X"32",X"F7",X"9B",X"FE",
		X"04",X"C0",X"3A",X"F6",X"9B",X"C6",X"01",X"32",X"F6",X"9B",X"AF",X"32",X"F7",X"9B",X"C9",X"3A",
		X"F8",X"9B",X"C6",X"01",X"32",X"F8",X"9B",X"FE",X"01",X"C0",X"3A",X"F6",X"9B",X"3C",X"32",X"F6",
		X"9B",X"AF",X"32",X"F8",X"9B",X"C9",X"3A",X"F8",X"9B",X"C6",X"01",X"32",X"F8",X"9B",X"FE",X"01",
		X"C0",X"3A",X"F6",X"9B",X"C6",X"02",X"32",X"F6",X"9B",X"AF",X"32",X"F8",X"9B",X"C9",X"3A",X"F8",
		X"9B",X"C6",X"01",X"32",X"F8",X"9B",X"FE",X"01",X"C0",X"3A",X"F6",X"9B",X"C6",X"03",X"32",X"F6",
		X"9B",X"AF",X"32",X"F8",X"9B",X"C9",X"3A",X"F8",X"9B",X"C6",X"01",X"32",X"F8",X"9B",X"FE",X"02",
		X"C0",X"3A",X"F6",X"9B",X"C6",X"01",X"32",X"F6",X"9B",X"AF",X"32",X"F8",X"9B",X"C9",X"3A",X"F8",
		X"9B",X"C6",X"01",X"32",X"F8",X"9B",X"FE",X"02",X"C0",X"3A",X"F6",X"9B",X"C6",X"03",X"32",X"F6",
		X"9B",X"AF",X"32",X"F8",X"9B",X"C9",X"3A",X"F8",X"9B",X"C6",X"01",X"32",X"F8",X"9B",X"FE",X"03",
		X"C0",X"3A",X"F6",X"9B",X"C6",X"01",X"32",X"F6",X"9B",X"AF",X"32",X"F8",X"9B",X"C9",X"3A",X"F8",
		X"9B",X"C6",X"01",X"32",X"F8",X"9B",X"FE",X"04",X"C0",X"3A",X"F6",X"9B",X"C6",X"01",X"32",X"F6",
		X"9B",X"AF",X"32",X"F8",X"9B",X"C9",X"2A",X"59",X"9A",X"23",X"22",X"59",X"9A",X"C9",X"3A",X"66",
		X"9A",X"FE",X"0F",X"CA",X"55",X"04",X"FE",X"1F",X"CA",X"EE",X"04",X"CD",X"DB",X"0A",X"CD",X"8F",
		X"07",X"CD",X"DB",X"0A",X"C9",X"CD",X"F2",X"12",X"3A",X"5D",X"9A",X"A7",X"C2",X"7E",X"04",X"3A",
		X"8F",X"9C",X"A7",X"3E",X"00",X"32",X"8F",X"9C",X"C2",X"E1",X"04",X"3A",X"90",X"9C",X"A7",X"3E",
		X"00",X"32",X"90",X"9C",X"C2",X"BB",X"04",X"DD",X"21",X"67",X"9A",X"C3",X"9A",X"04",X"3A",X"91",
		X"9C",X"A7",X"3E",X"00",X"32",X"91",X"9C",X"C2",X"E7",X"04",X"3A",X"92",X"9C",X"A7",X"3E",X"00",
		X"32",X"92",X"9C",X"C2",X"BB",X"04",X"DD",X"21",X"25",X"9B",X"DD",X"7E",X"00",X"32",X"8B",X"9C",
		X"DD",X"7E",X"01",X"32",X"53",X"9A",X"DD",X"E5",X"E1",X"23",X"23",X"11",X"40",X"9A",X"01",X"11",
		X"00",X"ED",X"B0",X"11",X"50",X"99",X"01",X"A0",X"00",X"ED",X"B0",X"CD",X"1E",X"14",X"CD",X"D1",
		X"12",X"CD",X"09",X"14",X"CD",X"B3",X"12",X"CD",X"F7",X"0F",X"CD",X"2B",X"11",X"CD",X"5C",X"0E",
		X"CD",X"E1",X"0A",X"3E",X"1F",X"32",X"66",X"9A",X"3E",X"03",X"CD",X"09",X"11",X"CD",X"E1",X"0A",
		X"C9",X"CD",X"A3",X"12",X"C3",X"BB",X"04",X"AF",X"32",X"8B",X"9C",X"C3",X"E1",X"04",X"CD",X"6E",
		X"15",X"CD",X"D0",X"20",X"CD",X"B7",X"21",X"CD",X"3B",X"24",X"CD",X"CF",X"25",X"CD",X"0B",X"28",
		X"CD",X"AD",X"19",X"CD",X"0A",X"05",X"CD",X"12",X"05",X"C9",X"3A",X"59",X"9A",X"3C",X"32",X"59",
		X"9A",X"C9",X"3A",X"51",X"9A",X"A7",X"CA",X"2D",X"05",X"3E",X"00",X"32",X"66",X"9A",X"32",X"51",
		X"9A",X"32",X"8C",X"9C",X"CD",X"DB",X"0A",X"3E",X"08",X"CD",X"09",X"11",X"C9",X"3A",X"8B",X"9C",
		X"FE",X"10",X"D8",X"DD",X"21",X"50",X"99",X"01",X"20",X"00",X"16",X"05",X"3E",X"00",X"DD",X"B6",
		X"00",X"DD",X"09",X"15",X"C2",X"3E",X"05",X"A7",X"C0",X"AF",X"32",X"8B",X"9C",X"3E",X"06",X"CD",
		X"09",X"11",X"CD",X"AA",X"05",X"CD",X"98",X"05",X"3A",X"40",X"9A",X"3C",X"32",X"40",X"9A",X"FE",
		X"04",X"D2",X"8E",X"05",X"CD",X"0D",X"13",X"21",X"41",X"9A",X"11",X"42",X"9A",X"01",X"10",X"00",
		X"36",X"00",X"ED",X"B0",X"3E",X"0F",X"32",X"66",X"9A",X"3A",X"5D",X"9A",X"A7",X"C2",X"86",X"05",
		X"3E",X"FF",X"32",X"90",X"9C",X"C9",X"3E",X"FF",X"32",X"92",X"9C",X"C9",X"04",X"C9",X"AF",X"32",
		X"40",X"9A",X"CD",X"D6",X"10",X"C3",X"64",X"05",X"3A",X"53",X"9A",X"3C",X"FE",X"04",X"D2",X"A5",
		X"05",X"32",X"53",X"9A",X"C9",X"AF",X"32",X"53",X"9A",X"C9",X"CD",X"B5",X"10",X"CD",X"F2",X"12",
		X"21",X"B0",X"44",X"CD",X"84",X"10",X"21",X"B9",X"44",X"CD",X"84",X"10",X"16",X"03",X"CD",X"51",
		X"36",X"21",X"41",X"9A",X"0E",X"08",X"06",X"00",X"7E",X"A7",X"CC",X"8C",X"05",X"23",X"23",X"0D",
		X"C2",X"C8",X"05",X"78",X"32",X"2B",X"86",X"4F",X"06",X"00",X"DD",X"21",X"C3",X"44",X"CB",X"21",
		X"CB",X"10",X"DD",X"09",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"22",X"5B",X"9A",X"DD",X"21",X"11",
		X"45",X"DD",X"09",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"CD",X"84",X"10",X"3E",X"08",X"CD",X"09",
		X"11",X"C9",X"3A",X"E6",X"9B",X"A7",X"CA",X"5D",X"06",X"FE",X"0F",X"CA",X"92",X"06",X"CD",X"3E",
		X"04",X"CD",X"21",X"06",X"3A",X"EE",X"9B",X"A7",X"C8",X"CD",X"CA",X"06",X"AF",X"32",X"E6",X"9B",
		X"C9",X"3A",X"59",X"9A",X"E6",X"1F",X"C0",X"2A",X"E7",X"9B",X"23",X"22",X"E7",X"9B",X"E5",X"01",
		X"A0",X"00",X"A7",X"ED",X"42",X"E1",X"D2",X"56",X"06",X"CB",X"3C",X"CB",X"1D",X"CB",X"3C",X"CB",
		X"1D",X"01",X"D9",X"44",X"09",X"7E",X"32",X"54",X"9A",X"CB",X"45",X"C8",X"AF",X"32",X"55",X"9A",
		X"3E",X"FF",X"32",X"56",X"9A",X"C9",X"21",X"00",X"00",X"22",X"E7",X"9B",X"C9",X"CD",X"B5",X"10",
		X"CD",X"F2",X"12",X"CD",X"5C",X"0B",X"CD",X"DB",X"0A",X"AF",X"32",X"5D",X"9A",X"32",X"E3",X"9B",
		X"32",X"EE",X"9B",X"3E",X"00",X"32",X"E4",X"9B",X"3E",X"0F",X"32",X"E6",X"9B",X"21",X"00",X"00",
		X"22",X"E7",X"9B",X"22",X"87",X"9C",X"3E",X"01",X"32",X"EA",X"9B",X"32",X"52",X"9A",X"CD",X"A3",
		X"12",X"C9",X"CD",X"E4",X"06",X"CD",X"0A",X"05",X"2A",X"E7",X"9B",X"01",X"FA",X"00",X"A7",X"ED",
		X"42",X"D8",X"3E",X"08",X"CD",X"09",X"11",X"3E",X"FF",X"32",X"E6",X"9B",X"3E",X"0F",X"32",X"66",
		X"9A",X"3E",X"FF",X"32",X"8F",X"9C",X"AF",X"32",X"90",X"9C",X"32",X"EE",X"9B",X"2F",X"32",X"EF",
		X"9B",X"3E",X"01",X"32",X"52",X"9A",X"CD",X"F2",X"12",X"C9",X"3A",X"E9",X"9B",X"FE",X"03",X"D2",
		X"D7",X"06",X"3C",X"32",X"E9",X"9B",X"C9",X"AF",X"32",X"E9",X"9B",X"CD",X"A5",X"3A",X"3E",X"08",
		X"CD",X"09",X"11",X"C9",X"3A",X"59",X"9A",X"E6",X"7F",X"C0",X"CD",X"63",X"08",X"CD",X"9D",X"08",
		X"CD",X"16",X"09",X"CD",X"83",X"0A",X"CD",X"B1",X"0A",X"2A",X"E7",X"9B",X"23",X"22",X"E7",X"9B",
		X"C9",X"CD",X"B5",X"10",X"CD",X"F2",X"12",X"CD",X"0D",X"13",X"CD",X"6B",X"12",X"CD",X"D9",X"11",
		X"3E",X"01",X"32",X"81",X"A1",X"C9",X"CD",X"B5",X"10",X"CD",X"FB",X"10",X"CD",X"07",X"0F",X"CD",
		X"F2",X"12",X"CD",X"0D",X"13",X"CD",X"F7",X"0F",X"CD",X"A3",X"12",X"21",X"00",X"00",X"22",X"5B",
		X"9A",X"3E",X"0F",X"32",X"66",X"9A",X"3E",X"01",X"32",X"EA",X"9B",X"32",X"EB",X"9B",X"32",X"52",
		X"9A",X"CD",X"D5",X"0C",X"AF",X"32",X"EC",X"9B",X"32",X"ED",X"9B",X"32",X"51",X"9A",X"32",X"53",
		X"9A",X"32",X"E6",X"9B",X"32",X"8B",X"9C",X"32",X"8C",X"9C",X"CD",X"B3",X"12",X"3A",X"E3",X"9B",
		X"A7",X"C2",X"77",X"07",X"AF",X"3A",X"5D",X"9A",X"32",X"90",X"9C",X"2F",X"32",X"EF",X"9B",X"32",
		X"8F",X"9C",X"AF",X"32",X"EE",X"9B",X"C9",X"AF",X"32",X"5D",X"9A",X"32",X"EF",X"9B",X"32",X"90",
		X"9C",X"32",X"92",X"9C",X"3E",X"FF",X"32",X"91",X"9C",X"32",X"8F",X"9C",X"C3",X"72",X"07",X"CD",
		X"37",X"08",X"CD",X"0D",X"13",X"CD",X"F2",X"12",X"3A",X"E3",X"9B",X"A7",X"C2",X"BE",X"07",X"3A",
		X"E4",X"9B",X"A7",X"CA",X"B0",X"07",X"3D",X"32",X"E4",X"9B",X"3E",X"0F",X"32",X"66",X"9A",X"C9",
		X"CD",X"51",X"11",X"3E",X"08",X"CD",X"09",X"11",X"3E",X"FF",X"32",X"EE",X"9B",X"C9",X"3A",X"5D",
		X"9A",X"A7",X"C2",X"FE",X"07",X"3A",X"E4",X"9B",X"A7",X"CA",X"E1",X"07",X"3D",X"32",X"E4",X"9B",
		X"3A",X"EF",X"9B",X"A7",X"CA",X"F3",X"07",X"AF",X"32",X"5D",X"9A",X"3E",X"0F",X"32",X"66",X"9A",
		X"C9",X"CD",X"43",X"11",X"3E",X"08",X"CD",X"09",X"11",X"3E",X"FF",X"32",X"EE",X"9B",X"3A",X"EF",
		X"9B",X"A7",X"C0",X"3E",X"FF",X"32",X"5D",X"9A",X"3E",X"0F",X"32",X"66",X"9A",X"C9",X"3A",X"E5",
		X"9B",X"A7",X"CA",X"1B",X"08",X"3D",X"32",X"E5",X"9B",X"3A",X"EE",X"9B",X"A7",X"CA",X"2D",X"08",
		X"3E",X"FF",X"32",X"5D",X"9A",X"3E",X"0F",X"32",X"66",X"9A",X"C9",X"CD",X"4A",X"11",X"3E",X"08",
		X"CD",X"09",X"11",X"3E",X"FF",X"32",X"EF",X"9B",X"3A",X"EE",X"9B",X"A7",X"C0",X"AF",X"32",X"5D",
		X"9A",X"3E",X"0F",X"32",X"66",X"9A",X"C9",X"3A",X"5D",X"9A",X"A7",X"C2",X"44",X"08",X"11",X"67",
		X"9A",X"C3",X"47",X"08",X"11",X"25",X"9B",X"3A",X"8B",X"9C",X"12",X"21",X"53",X"9A",X"13",X"7E",
		X"12",X"13",X"21",X"40",X"9A",X"01",X"11",X"00",X"ED",X"B0",X"21",X"50",X"99",X"01",X"A0",X"00",
		X"ED",X"B0",X"C9",X"3A",X"87",X"9C",X"A7",X"C0",X"DD",X"21",X"B3",X"40",X"ED",X"4B",X"E7",X"9B",
		X"CB",X"21",X"CB",X"10",X"DD",X"09",X"DD",X"7E",X"00",X"FE",X"FF",X"CA",X"97",X"08",X"FE",X"F0",
		X"CA",X"8D",X"08",X"DD",X"56",X"00",X"DD",X"5E",X"01",X"CD",X"9C",X"33",X"C9",X"DD",X"56",X"00",
		X"DD",X"5E",X"01",X"CD",X"B0",X"33",X"C9",X"3E",X"FF",X"32",X"87",X"9C",X"C9",X"2A",X"E7",X"9B",
		X"01",X"28",X"00",X"A7",X"ED",X"42",X"D8",X"DD",X"21",X"E7",X"42",X"0E",X"07",X"DD",X"5E",X"00",
		X"DD",X"56",X"01",X"A7",X"ED",X"52",X"CA",X"C4",X"08",X"DD",X"23",X"DD",X"23",X"DD",X"23",X"0D",
		X"C2",X"AD",X"08",X"C9",X"DD",X"4E",X"02",X"06",X"00",X"CB",X"21",X"CB",X"10",X"DD",X"21",X"FC",
		X"42",X"DD",X"09",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"E5",X"E5",X"E5",X"E5",X"FD",X"E1",X"DD",
		X"E1",X"0E",X"0C",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"FD",X"7E",X"18",X"77",X"DD",X"23",X"DD",
		X"23",X"FD",X"23",X"0D",X"C2",X"E3",X"08",X"DD",X"E1",X"FD",X"E1",X"11",X"00",X"08",X"0E",X"0C",
		X"DD",X"6E",X"00",X"DD",X"66",X"01",X"19",X"FD",X"7E",X"24",X"77",X"DD",X"23",X"DD",X"23",X"FD",
		X"23",X"0D",X"C2",X"00",X"09",X"C9",X"3A",X"88",X"9C",X"A7",X"C0",X"2A",X"E7",X"9B",X"01",X"64",
		X"00",X"A7",X"ED",X"42",X"D8",X"01",X"24",X"43",X"CB",X"25",X"CB",X"14",X"09",X"E5",X"DD",X"E1",
		X"DD",X"7E",X"00",X"FE",X"FF",X"CA",X"7D",X"0A",X"57",X"DD",X"5E",X"01",X"F5",X"CD",X"82",X"34",
		X"F1",X"32",X"63",X"9A",X"47",X"3A",X"62",X"9A",X"4F",X"3E",X"01",X"32",X"62",X"9A",X"78",X"FE",
		X"40",X"CA",X"84",X"09",X"FE",X"60",X"CA",X"A3",X"09",X"FE",X"70",X"CA",X"C2",X"09",X"FE",X"90",
		X"CA",X"E1",X"09",X"FE",X"A0",X"CA",X"39",X"0A",X"FE",X"B0",X"CA",X"45",X"0A",X"FE",X"C0",X"CA",
		X"51",X"0A",X"FE",X"F0",X"D2",X"7C",X"09",X"79",X"32",X"62",X"9A",X"C9",X"DD",X"5E",X"01",X"57",
		X"CD",X"B0",X"33",X"C9",X"21",X"6B",X"45",X"CD",X"84",X"10",X"16",X"28",X"1E",X"88",X"26",X"8B",
		X"2E",X"10",X"3E",X"00",X"CD",X"62",X"32",X"DD",X"21",X"97",X"41",X"FD",X"21",X"BB",X"41",X"CD",
		X"5D",X"0A",X"C9",X"21",X"82",X"45",X"CD",X"84",X"10",X"16",X"28",X"1E",X"A0",X"26",X"AF",X"2E",
		X"13",X"3E",X"01",X"CD",X"62",X"32",X"DD",X"21",X"C7",X"41",X"FD",X"21",X"EB",X"41",X"CD",X"5D",
		X"0A",X"C9",X"21",X"93",X"45",X"CD",X"84",X"10",X"16",X"28",X"1E",X"B8",X"26",X"67",X"2E",X"12",
		X"3E",X"02",X"CD",X"62",X"32",X"DD",X"21",X"F7",X"41",X"FD",X"21",X"1B",X"42",X"CD",X"5D",X"0A",
		X"C9",X"21",X"A4",X"45",X"CD",X"84",X"10",X"CD",X"F6",X"09",X"DD",X"21",X"27",X"42",X"FD",X"21",
		X"4B",X"42",X"CD",X"5D",X"0A",X"C9",X"FD",X"21",X"67",X"84",X"DD",X"21",X"BC",X"4C",X"DD",X"E5",
		X"11",X"04",X"00",X"3E",X"06",X"DD",X"4E",X"00",X"FD",X"71",X"00",X"DD",X"4E",X"01",X"FD",X"71",
		X"20",X"DD",X"4E",X"02",X"FD",X"71",X"40",X"DD",X"4E",X"03",X"FD",X"71",X"60",X"DD",X"19",X"FD",
		X"2B",X"3D",X"C8",X"FE",X"03",X"C2",X"05",X"0A",X"DD",X"E1",X"11",X"0C",X"00",X"DD",X"19",X"11",
		X"04",X"00",X"FD",X"21",X"67",X"8C",X"C3",X"05",X"0A",X"DD",X"21",X"B7",X"42",X"FD",X"21",X"DB",
		X"42",X"CD",X"5D",X"0A",X"C9",X"DD",X"21",X"57",X"42",X"FD",X"21",X"7B",X"42",X"CD",X"5D",X"0A",
		X"C9",X"DD",X"21",X"87",X"42",X"FD",X"21",X"AB",X"42",X"CD",X"5D",X"0A",X"C9",X"11",X"00",X"08",
		X"06",X"04",X"0E",X"0C",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"FD",X"7E",X"00",X"E6",X"F0",X"80",
		X"19",X"77",X"DD",X"23",X"DD",X"23",X"FD",X"23",X"0D",X"C2",X"64",X"0A",X"C9",X"3E",X"FF",X"32",
		X"88",X"9C",X"C9",X"2A",X"E7",X"9B",X"01",X"64",X"00",X"A7",X"ED",X"42",X"C0",X"21",X"23",X"85",
		X"FD",X"21",X"23",X"8D",X"DD",X"21",X"0A",X"43",X"0E",X"0D",X"11",X"20",X"00",X"DD",X"7E",X"00",
		X"77",X"DD",X"7E",X"0D",X"FD",X"77",X"00",X"DD",X"23",X"FD",X"19",X"19",X"0D",X"C2",X"9D",X"0A",
		X"C9",X"3A",X"62",X"9A",X"A7",X"C8",X"4F",X"3C",X"32",X"62",X"9A",X"06",X"00",X"21",X"B5",X"45",
		X"09",X"7E",X"FE",X"50",X"D2",X"D6",X"0A",X"5F",X"3A",X"63",X"9A",X"57",X"26",X"08",X"2E",X"00",
		X"3E",X"00",X"CD",X"0E",X"32",X"C9",X"AF",X"32",X"62",X"9A",X"C9",X"21",X"17",X"9C",X"CB",X"C6",
		X"C9",X"3A",X"E6",X"9B",X"A7",X"C0",X"21",X"17",X"9C",X"CB",X"CE",X"C9",X"3A",X"E6",X"9B",X"A7",
		X"C4",X"36",X"0B",X"3A",X"17",X"9C",X"47",X"3E",X"00",X"32",X"17",X"9C",X"CB",X"40",X"C2",X"4E",
		X"0B",X"CB",X"48",X"C2",X"49",X"0B",X"3A",X"16",X"9C",X"CB",X"47",X"C2",X"53",X"0B",X"3A",X"16",
		X"9C",X"47",X"CB",X"F8",X"CB",X"80",X"CD",X"3C",X"0B",X"AF",X"32",X"16",X"9C",X"78",X"32",X"00",
		X"A1",X"3E",X"01",X"32",X"80",X"A1",X"00",X"00",X"00",X"AF",X"32",X"80",X"A1",X"00",X"00",X"00",
		X"3E",X"01",X"32",X"80",X"A1",X"C9",X"3E",X"00",X"32",X"16",X"9C",X"C9",X"3A",X"15",X"9C",X"A7",
		X"3E",X"00",X"32",X"15",X"9C",X"C8",X"CB",X"C0",X"C9",X"3E",X"02",X"C3",X"1E",X"0B",X"3E",X"01",
		X"C3",X"1E",X"0B",X"AF",X"32",X"16",X"9C",X"3E",X"04",X"C3",X"1E",X"0B",X"DD",X"21",X"CD",X"45",
		X"FD",X"21",X"00",X"00",X"0E",X"30",X"3E",X"00",X"DD",X"86",X"00",X"FD",X"86",X"00",X"DD",X"23",
		X"FD",X"23",X"0D",X"C2",X"68",X"0B",X"FE",X"F3",X"C8",X"21",X"CD",X"45",X"CD",X"84",X"10",X"21",
		X"DD",X"45",X"CD",X"84",X"10",X"C3",X"79",X"0B",X"3A",X"E6",X"9B",X"A7",X"C0",X"3A",X"56",X"9A",
		X"32",X"55",X"9A",X"3A",X"58",X"9A",X"32",X"57",X"9A",X"AF",X"32",X"56",X"9A",X"32",X"58",X"9A",
		X"32",X"54",X"9A",X"3A",X"E3",X"9B",X"A7",X"CA",X"DE",X"0B",X"3A",X"00",X"9C",X"A7",X"C2",X"DE",
		X"0B",X"3A",X"5D",X"9A",X"A7",X"CA",X"DE",X"0B",X"3A",X"80",X"A0",X"CB",X"5F",X"CC",X"37",X"0C",
		X"CD",X"13",X"0C",X"3A",X"00",X"A0",X"CB",X"47",X"CA",X"1F",X"0C",X"3A",X"80",X"A0",X"CB",X"4F",
		X"CA",X"25",X"0C",X"CB",X"6F",X"CA",X"2B",X"0C",X"CB",X"67",X"CA",X"31",X"0C",X"C9",X"3A",X"00",
		X"A0",X"CB",X"5F",X"CC",X"37",X"0C",X"CD",X"07",X"0C",X"3A",X"80",X"A0",X"CB",X"47",X"CA",X"1F",
		X"0C",X"3A",X"00",X"A0",X"CB",X"6F",X"CA",X"31",X"0C",X"CB",X"67",X"CA",X"2B",X"0C",X"3A",X"00",
		X"A1",X"CB",X"7F",X"CA",X"25",X"0C",X"C9",X"3A",X"00",X"A1",X"CB",X"77",X"C0",X"3E",X"FF",X"32",
		X"58",X"9A",X"C9",X"3A",X"80",X"A0",X"CB",X"57",X"C0",X"3E",X"FF",X"32",X"58",X"9A",X"C9",X"3E",
		X"10",X"32",X"54",X"9A",X"C9",X"3E",X"20",X"32",X"54",X"9A",X"C9",X"3E",X"02",X"32",X"54",X"9A",
		X"C9",X"3E",X"01",X"32",X"54",X"9A",X"C9",X"3E",X"FF",X"32",X"56",X"9A",X"C9",X"CD",X"5B",X"0C",
		X"CD",X"32",X"0D",X"CD",X"BE",X"0D",X"3A",X"5D",X"9A",X"A7",X"C2",X"54",X"0C",X"3A",X"EA",X"9B",
		X"32",X"52",X"9A",X"C9",X"3A",X"EB",X"9B",X"32",X"52",X"9A",X"C9",X"3A",X"5D",X"9A",X"A7",X"C2",
		X"6D",X"0C",X"DD",X"21",X"0D",X"9C",X"FD",X"21",X"01",X"9C",X"C3",X"78",X"0C",X"DD",X"21",X"10",
		X"9C",X"FD",X"21",X"07",X"9C",X"C3",X"78",X"0C",X"3A",X"FD",X"9B",X"A7",X"C2",X"D5",X"0C",X"2A",
		X"5B",X"9A",X"7C",X"B5",X"C8",X"DD",X"7E",X"02",X"85",X"27",X"DD",X"77",X"02",X"DD",X"7E",X"01",
		X"8C",X"27",X"DD",X"77",X"01",X"06",X"00",X"DD",X"7E",X"00",X"88",X"27",X"DD",X"77",X"00",X"21",
		X"00",X"00",X"22",X"5B",X"9A",X"DD",X"E5",X"E1",X"AF",X"ED",X"6F",X"FD",X"77",X"00",X"ED",X"67",
		X"7E",X"E6",X"0F",X"FD",X"77",X"01",X"23",X"ED",X"6F",X"FD",X"77",X"02",X"ED",X"67",X"7E",X"E6",
		X"0F",X"FD",X"77",X"03",X"23",X"ED",X"6F",X"FD",X"77",X"04",X"ED",X"67",X"7E",X"E6",X"0F",X"FD",
		X"77",X"05",X"CD",X"D1",X"0E",X"3A",X"5D",X"9A",X"A7",X"C2",X"E6",X"0C",X"21",X"66",X"80",X"FD",
		X"21",X"01",X"9C",X"C3",X"ED",X"0C",X"21",X"E6",X"82",X"FD",X"21",X"07",X"9C",X"11",X"20",X"00",
		X"06",X"06",X"FD",X"7E",X"00",X"77",X"19",X"FD",X"23",X"05",X"C2",X"F2",X"0C",X"3A",X"52",X"9A",
		X"CB",X"47",X"CA",X"1C",X"0D",X"11",X"00",X"08",X"19",X"11",X"E0",X"FF",X"19",X"06",X"06",X"36",
		X"00",X"19",X"05",X"C2",X"0F",X"0D",X"19",X"AF",X"32",X"FD",X"9B",X"C9",X"11",X"00",X"08",X"19",
		X"11",X"E0",X"FF",X"19",X"06",X"06",X"36",X"10",X"19",X"05",X"C2",X"26",X"0D",X"AF",X"32",X"FD",
		X"9B",X"C9",X"3A",X"E3",X"9B",X"A7",X"C8",X"3A",X"5D",X"9A",X"A7",X"C2",X"81",X"0D",X"DD",X"21",
		X"67",X"80",X"FD",X"21",X"E7",X"82",X"01",X"01",X"02",X"3A",X"59",X"9A",X"5F",X"E6",X"3F",X"CA",
		X"8F",X"0D",X"7B",X"C6",X"20",X"E6",X"3F",X"C0",X"DD",X"71",X"00",X"DD",X"36",X"20",X"1E",X"DD",
		X"36",X"40",X"19",X"01",X"00",X"08",X"DD",X"09",X"06",X"03",X"3A",X"52",X"9A",X"CB",X"47",X"CC",
		X"7C",X"0D",X"DD",X"70",X"00",X"DD",X"70",X"20",X"DD",X"70",X"40",X"C9",X"3E",X"FF",X"CB",X"E0",
		X"C9",X"DD",X"21",X"E7",X"82",X"FD",X"21",X"67",X"80",X"01",X"02",X"01",X"C3",X"49",X"0D",X"3E",
		X"7F",X"DD",X"77",X"00",X"DD",X"77",X"20",X"DD",X"77",X"40",X"FD",X"70",X"00",X"FD",X"36",X"20",
		X"1E",X"FD",X"36",X"40",X"19",X"01",X"00",X"08",X"FD",X"09",X"06",X"03",X"3A",X"52",X"9A",X"CB",
		X"47",X"CC",X"7C",X"0D",X"FD",X"70",X"00",X"FD",X"70",X"20",X"FD",X"70",X"40",X"C9",X"DD",X"21",
		X"0D",X"9C",X"FD",X"21",X"10",X"9C",X"DD",X"7E",X"00",X"FD",X"BE",X"00",X"DA",X"0E",X"0E",X"C2",
		X"E7",X"0D",X"DD",X"7E",X"01",X"FD",X"BE",X"01",X"DA",X"0E",X"0E",X"C2",X"E7",X"0D",X"DD",X"7E",
		X"02",X"FD",X"BE",X"02",X"DA",X"0E",X"0E",X"DD",X"21",X"0D",X"9C",X"FD",X"21",X"73",X"9C",X"DD",
		X"7E",X"00",X"FD",X"BE",X"00",X"D8",X"C2",X"19",X"0E",X"DD",X"7E",X"01",X"FD",X"BE",X"01",X"D8",
		X"C2",X"19",X"0E",X"DD",X"7E",X"02",X"FD",X"BE",X"02",X"D8",X"C8",X"C3",X"19",X"0E",X"DD",X"21",
		X"10",X"9C",X"FD",X"21",X"73",X"9C",X"C3",X"EF",X"0D",X"DD",X"7E",X"00",X"DD",X"46",X"01",X"DD",
		X"4E",X"02",X"FD",X"77",X"00",X"FD",X"70",X"01",X"FD",X"71",X"02",X"FD",X"E5",X"E1",X"DD",X"21",
		X"6D",X"9C",X"AF",X"ED",X"6F",X"DD",X"77",X"00",X"ED",X"67",X"7E",X"E6",X"0F",X"DD",X"77",X"01",
		X"23",X"ED",X"6F",X"DD",X"77",X"02",X"ED",X"67",X"7E",X"E6",X"0F",X"DD",X"77",X"03",X"23",X"ED",
		X"6F",X"DD",X"77",X"04",X"ED",X"67",X"7E",X"E6",X"0F",X"DD",X"77",X"05",X"3A",X"E3",X"9B",X"A7",
		X"C2",X"6D",X"0E",X"21",X"87",X"81",X"DD",X"21",X"6D",X"9C",X"C3",X"77",X"0E",X"21",X"87",X"81",
		X"DD",X"21",X"6D",X"9C",X"C3",X"77",X"0E",X"11",X"20",X"00",X"E5",X"36",X"11",X"19",X"36",X"12",
		X"19",X"36",X"4D",X"19",X"36",X"1C",X"19",X"36",X"0C",X"19",X"36",X"18",X"19",X"36",X"1B",X"19",
		X"36",X"0E",X"19",X"E1",X"E5",X"2B",X"19",X"0E",X"06",X"DD",X"7E",X"00",X"77",X"19",X"DD",X"23",
		X"0D",X"C2",X"99",X"0E",X"E1",X"01",X"00",X"08",X"09",X"E5",X"0E",X"08",X"06",X"08",X"3A",X"52",
		X"9A",X"CB",X"47",X"CC",X"7C",X"0D",X"70",X"19",X"0D",X"C2",X"B6",X"0E",X"0E",X"07",X"E1",X"2B",
		X"06",X"00",X"3A",X"52",X"9A",X"CB",X"47",X"CC",X"7C",X"0D",X"70",X"19",X"0D",X"C2",X"CA",X"0E",
		X"C9",X"3A",X"5D",X"9A",X"A7",X"C2",X"E1",X"0E",X"11",X"EC",X"9B",X"21",X"E4",X"9B",X"C3",X"EA",
		X"0E",X"11",X"ED",X"9B",X"21",X"E5",X"9B",X"C3",X"EA",X"0E",X"1A",X"A7",X"C0",X"FD",X"7E",X"00",
		X"A7",X"C2",X"FD",X"0E",X"3A",X"FE",X"9B",X"47",X"FD",X"7E",X"01",X"B8",X"D8",X"7E",X"3C",X"77",
		X"3E",X"FF",X"12",X"CD",X"F7",X"0F",X"C9",X"3A",X"FF",X"9B",X"E6",X"03",X"47",X"3A",X"E3",X"9B",
		X"A7",X"C2",X"19",X"0F",X"0E",X"00",X"C3",X"1B",X"0F",X"0E",X"FF",X"78",X"FE",X"00",X"CA",X"2E",
		X"0F",X"FE",X"01",X"CA",X"38",X"0F",X"FE",X"02",X"CA",X"42",X"0F",X"C3",X"4C",X"0F",X"3E",X"02",
		X"32",X"E4",X"9B",X"A1",X"32",X"E5",X"9B",X"C9",X"3E",X"03",X"32",X"E4",X"9B",X"A1",X"32",X"E5",
		X"9B",X"C9",X"3E",X"04",X"32",X"E4",X"9B",X"A1",X"32",X"E5",X"9B",X"C9",X"3E",X"05",X"32",X"E4",
		X"9B",X"A1",X"32",X"E5",X"9B",X"C9",X"21",X"80",X"86",X"11",X"20",X"00",X"0E",X"08",X"FD",X"21",
		X"4B",X"3D",X"FD",X"7E",X"00",X"77",X"19",X"FD",X"23",X"0D",X"C2",X"62",X"0F",X"21",X"80",X"8E",
		X"3E",X"00",X"0E",X"0A",X"77",X"19",X"0D",X"C2",X"74",X"0F",X"3A",X"F6",X"9B",X"FE",X"64",X"D2",
		X"A7",X"0F",X"A7",X"CA",X"B4",X"0F",X"47",X"0E",X"01",X"AF",X"81",X"27",X"05",X"C2",X"8A",X"0F",
		X"FD",X"21",X"60",X"87",X"47",X"E6",X"0F",X"FD",X"77",X"20",X"78",X"CB",X"3F",X"CB",X"3F",X"CB",
		X"3F",X"CB",X"3F",X"FD",X"77",X"00",X"C9",X"FD",X"21",X"60",X"87",X"3E",X"28",X"FD",X"77",X"00",
		X"FD",X"77",X"20",X"C9",X"FD",X"21",X"60",X"87",X"AF",X"FD",X"77",X"20",X"C9",X"3A",X"E3",X"9B",
		X"A7",X"CA",X"D7",X"0F",X"3A",X"00",X"9C",X"A7",X"C2",X"D7",X"0F",X"3A",X"5D",X"9A",X"A7",X"CA",
		X"D7",X"0F",X"AF",X"32",X"83",X"A1",X"C9",X"3E",X"01",X"32",X"83",X"A1",X"C9",X"E5",X"DD",X"E1",
		X"D9",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"DD",X"4E",X"00",X"11",X"20",X"00",X"3E",X"FF",X"77",
		X"19",X"0D",X"C2",X"EF",X"0F",X"D9",X"C9",X"3A",X"5D",X"9A",X"A7",X"C2",X"04",X"10",X"21",X"E4",
		X"9B",X"C3",X"07",X"10",X"21",X"E5",X"9B",X"7E",X"A7",X"CA",X"4E",X"10",X"F5",X"CD",X"4E",X"10",
		X"DD",X"21",X"41",X"84",X"11",X"40",X"00",X"F1",X"FE",X"08",X"D0",X"4F",X"DD",X"36",X"00",X"7C",
		X"DD",X"36",X"FF",X"7B",X"DD",X"36",X"20",X"7E",X"DD",X"36",X"1F",X"7D",X"DD",X"E5",X"D5",X"11",
		X"00",X"08",X"DD",X"19",X"DD",X"36",X"00",X"1C",X"DD",X"36",X"FF",X"1C",X"DD",X"36",X"20",X"1C",
		X"DD",X"36",X"1F",X"1C",X"D1",X"DD",X"E1",X"DD",X"19",X"0D",X"C2",X"1C",X"10",X"C9",X"21",X"41",
		X"84",X"11",X"20",X"00",X"3E",X"7A",X"0E",X"10",X"77",X"19",X"0D",X"C2",X"58",X"10",X"21",X"40",
		X"84",X"0E",X"10",X"77",X"19",X"0D",X"C2",X"63",X"10",X"21",X"41",X"8C",X"3E",X"00",X"0E",X"10",
		X"77",X"19",X"0D",X"C2",X"70",X"10",X"21",X"40",X"8C",X"0E",X"10",X"3E",X"00",X"77",X"19",X"0D",
		X"C2",X"7D",X"10",X"C9",X"E5",X"DD",X"E1",X"D9",X"DD",X"46",X"00",X"DD",X"4E",X"01",X"DD",X"6E",
		X"02",X"DD",X"66",X"03",X"E5",X"C5",X"11",X"20",X"00",X"DD",X"7E",X"04",X"77",X"19",X"DD",X"23",
		X"05",X"C2",X"99",X"10",X"C1",X"E1",X"11",X"00",X"08",X"19",X"11",X"20",X"00",X"71",X"19",X"05",
		X"C2",X"AD",X"10",X"D9",X"C9",X"21",X"40",X"80",X"0E",X"FF",X"11",X"80",X"07",X"71",X"23",X"1B",
		X"7A",X"B3",X"C2",X"BD",X"10",X"21",X"40",X"88",X"0E",X"00",X"11",X"80",X"07",X"71",X"23",X"1B",
		X"7A",X"B3",X"C2",X"CD",X"10",X"C9",X"CD",X"E0",X"10",X"21",X"00",X"50",X"22",X"5B",X"9A",X"C9",
		X"3A",X"5D",X"9A",X"A7",X"C2",X"F1",X"10",X"3A",X"EA",X"9B",X"C6",X"01",X"27",X"32",X"EA",X"9B",
		X"C9",X"3A",X"EB",X"9B",X"C6",X"01",X"27",X"32",X"EB",X"9B",X"C9",X"21",X"01",X"9C",X"11",X"02",
		X"9C",X"01",X"12",X"00",X"AF",X"77",X"ED",X"B0",X"C9",X"06",X"FF",X"0E",X"FF",X"0D",X"C2",X"0D",
		X"11",X"05",X"C2",X"0B",X"11",X"3D",X"C2",X"09",X"11",X"C9",X"21",X"00",X"80",X"01",X"FF",X"07",
		X"16",X"FF",X"72",X"23",X"0B",X"78",X"B1",X"C2",X"22",X"11",X"C9",X"3A",X"5D",X"9A",X"F5",X"AF",
		X"32",X"5D",X"9A",X"CD",X"D5",X"0C",X"3E",X"FF",X"32",X"5D",X"9A",X"CD",X"D5",X"0C",X"F1",X"32",
		X"5D",X"9A",X"C9",X"21",X"6A",X"3D",X"CD",X"84",X"10",X"C9",X"21",X"7E",X"3D",X"CD",X"84",X"10",
		X"C9",X"21",X"92",X"3D",X"CD",X"84",X"10",X"C9",X"21",X"9F",X"3D",X"CD",X"84",X"10",X"C9",X"3A",
		X"00",X"A0",X"CB",X"7F",X"3E",X"00",X"28",X"14",X"3A",X"13",X"9C",X"A7",X"CA",X"80",X"11",X"32",
		X"15",X"9C",X"2F",X"32",X"13",X"9C",X"CD",X"9F",X"02",X"C3",X"80",X"11",X"2F",X"32",X"13",X"9C",
		X"3A",X"00",X"A0",X"CB",X"77",X"3E",X"00",X"28",X"14",X"3A",X"14",X"9C",X"A7",X"CA",X"A1",X"11",
		X"32",X"15",X"9C",X"2F",X"32",X"14",X"9C",X"CD",X"C3",X"02",X"C3",X"A1",X"11",X"2F",X"32",X"14",
		X"9C",X"3A",X"00",X"A0",X"CB",X"67",X"C3",X"BD",X"11",X"3A",X"19",X"9C",X"A7",X"C0",X"2F",X"32",
		X"19",X"9C",X"32",X"15",X"9C",X"3A",X"F6",X"9B",X"3C",X"32",X"F6",X"9B",X"C9",X"AF",X"32",X"19",
		X"9C",X"C9",X"3A",X"80",X"A0",X"CB",X"7F",X"CA",X"D3",X"11",X"CB",X"77",X"C0",X"3E",X"FF",X"32",
		X"F3",X"9B",X"C9",X"3E",X"FF",X"32",X"F2",X"9B",X"C9",X"3A",X"80",X"A1",X"2F",X"32",X"FF",X"9B",
		X"5F",X"3A",X"00",X"A1",X"2F",X"57",X"CD",X"F3",X"11",X"CD",X"23",X"12",X"CD",X"48",X"12",X"CD",
		X"59",X"12",X"C9",X"7B",X"CB",X"3F",X"CB",X"3F",X"E6",X"07",X"21",X"F4",X"9B",X"FE",X"00",X"CA",
		X"2C",X"12",X"FE",X"01",X"CA",X"30",X"12",X"FE",X"02",X"CA",X"34",X"12",X"FE",X"03",X"CA",X"38",
		X"12",X"FE",X"04",X"CA",X"3C",X"12",X"FE",X"05",X"CA",X"40",X"12",X"FE",X"06",X"CA",X"44",X"12",
		X"36",X"FF",X"C9",X"21",X"F5",X"9B",X"7A",X"E6",X"07",X"C3",X"FD",X"11",X"3E",X"00",X"77",X"C9",
		X"3E",X"01",X"77",X"C9",X"3E",X"02",X"77",X"C9",X"3E",X"03",X"77",X"C9",X"3E",X"04",X"77",X"C9",
		X"3E",X"05",X"77",X"C9",X"3E",X"06",X"77",X"C9",X"7B",X"CB",X"7F",X"C2",X"53",X"12",X"AF",X"32",
		X"00",X"9C",X"C9",X"3E",X"FF",X"32",X"00",X"9C",X"C9",X"7B",X"CB",X"5F",X"C2",X"65",X"12",X"3E",
		X"03",X"32",X"FE",X"9B",X"C9",X"3E",X"05",X"32",X"FE",X"9B",X"C9",X"21",X"BC",X"3D",X"11",X"1A",
		X"9C",X"01",X"10",X"00",X"ED",X"B0",X"21",X"CC",X"3D",X"11",X"2A",X"9C",X"01",X"10",X"00",X"ED",
		X"B0",X"21",X"DC",X"3D",X"11",X"3A",X"9C",X"01",X"10",X"00",X"ED",X"B0",X"21",X"EC",X"3D",X"11",
		X"4A",X"9C",X"01",X"10",X"00",X"ED",X"B0",X"21",X"FC",X"3D",X"11",X"5A",X"9C",X"01",X"10",X"00",
		X"ED",X"B0",X"C9",X"21",X"37",X"3F",X"11",X"40",X"9A",X"01",X"11",X"00",X"ED",X"B0",X"AF",X"32",
		X"53",X"9A",X"C9",X"DD",X"21",X"20",X"9A",X"DD",X"36",X"03",X"80",X"DD",X"36",X"04",X"80",X"DD",
		X"36",X"00",X"FF",X"16",X"80",X"1E",X"E8",X"26",X"D3",X"2E",X"1A",X"3E",X"00",X"CD",X"62",X"32",
		X"C9",X"DD",X"21",X"40",X"9A",X"0E",X"08",X"06",X"01",X"50",X"C5",X"DD",X"7E",X"01",X"A7",X"F5",
		X"CC",X"51",X"36",X"F1",X"C4",X"A6",X"36",X"C1",X"DD",X"23",X"DD",X"23",X"04",X"0D",X"C2",X"D9",
		X"12",X"C9",X"21",X"00",X"80",X"0E",X"40",X"06",X"FF",X"70",X"23",X"0D",X"C2",X"F9",X"12",X"21",
		X"00",X"88",X"0E",X"40",X"06",X"FF",X"70",X"23",X"0D",X"C2",X"06",X"13",X"C9",X"21",X"00",X"98",
		X"11",X"01",X"98",X"01",X"3F",X"02",X"36",X"00",X"ED",X"B0",X"DD",X"21",X"00",X"98",X"FD",X"21",
		X"3B",X"3E",X"0E",X"09",X"11",X"10",X"00",X"CD",X"C3",X"13",X"DD",X"19",X"FD",X"23",X"FD",X"23",
		X"FD",X"23",X"0D",X"C2",X"27",X"13",X"DD",X"21",X"90",X"98",X"FD",X"21",X"56",X"3E",X"0E",X"02",
		X"11",X"10",X"00",X"CD",X"C3",X"13",X"DD",X"19",X"FD",X"23",X"FD",X"23",X"FD",X"23",X"0D",X"C2",
		X"43",X"13",X"DD",X"21",X"B0",X"98",X"FD",X"21",X"68",X"3E",X"0E",X"05",X"11",X"20",X"00",X"CD",
		X"E9",X"13",X"DD",X"19",X"FD",X"23",X"FD",X"23",X"FD",X"23",X"0D",X"C2",X"5F",X"13",X"DD",X"21",
		X"50",X"99",X"FD",X"21",X"86",X"3E",X"0E",X"05",X"11",X"20",X"00",X"CD",X"F6",X"13",X"DD",X"19",
		X"FD",X"23",X"FD",X"23",X"FD",X"23",X"0D",X"C2",X"7B",X"13",X"DD",X"21",X"F0",X"99",X"FD",X"21",
		X"5C",X"3E",X"0E",X"03",X"11",X"10",X"00",X"CD",X"E9",X"13",X"DD",X"19",X"FD",X"23",X"FD",X"23",
		X"FD",X"23",X"0D",X"C2",X"97",X"13",X"DD",X"21",X"20",X"9A",X"FD",X"21",X"65",X"3E",X"0E",X"01",
		X"11",X"20",X"00",X"CD",X"E9",X"13",X"DD",X"19",X"FD",X"23",X"FD",X"23",X"FD",X"23",X"0D",X"C2",
		X"B3",X"13",X"C9",X"FD",X"7E",X"00",X"DD",X"77",X"01",X"FD",X"7E",X"01",X"DD",X"77",X"02",X"FD",
		X"7E",X"02",X"DD",X"77",X"0E",X"C9",X"FD",X"7E",X"00",X"DD",X"77",X"01",X"FD",X"7E",X"01",X"DD",
		X"77",X"02",X"FD",X"7E",X"02",X"DD",X"77",X"03",X"C9",X"FD",X"7E",X"00",X"DD",X"77",X"01",X"FD",
		X"7E",X"01",X"DD",X"77",X"02",X"C9",X"FD",X"7E",X"00",X"DD",X"77",X"01",X"FD",X"7E",X"01",X"DD",
		X"77",X"02",X"FD",X"7E",X"02",X"DD",X"77",X"1F",X"C9",X"DD",X"21",X"50",X"99",X"01",X"20",X"00",
		X"16",X"05",X"1E",X"00",X"DD",X"73",X"07",X"DD",X"09",X"15",X"C2",X"14",X"14",X"C9",X"3A",X"52",
		X"9A",X"CB",X"47",X"CA",X"14",X"15",X"21",X"44",X"80",X"06",X"7F",X"0E",X"00",X"11",X"64",X"03",
		X"70",X"23",X"1B",X"7B",X"B2",X"C2",X"30",X"14",X"21",X"44",X"88",X"11",X"64",X"03",X"71",X"23",
		X"1B",X"7B",X"B2",X"C2",X"3E",X"14",X"DD",X"21",X"40",X"84",X"06",X"7A",X"0E",X"00",X"26",X"0B",
		X"11",X"20",X"00",X"CD",X"B9",X"14",X"DD",X"21",X"40",X"8C",X"41",X"26",X"0B",X"11",X"20",X"00",
		X"CD",X"B9",X"14",X"DD",X"21",X"4B",X"84",X"06",X"7F",X"26",X"11",X"11",X"20",X"00",X"CD",X"B9",
		X"14",X"DD",X"21",X"4B",X"8C",X"26",X"11",X"06",X"00",X"CD",X"B9",X"14",X"DD",X"21",X"95",X"3E",
		X"FD",X"21",X"CB",X"3E",X"0E",X"36",X"FD",X"6E",X"00",X"FD",X"66",X"01",X"DD",X"7E",X"00",X"77",
		X"FD",X"23",X"FD",X"23",X"DD",X"23",X"0D",X"C2",X"86",X"14",X"DD",X"21",X"CB",X"3E",X"0E",X"36",
		X"11",X"00",X"08",X"06",X"01",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"19",X"70",X"DD",X"23",X"DD",
		X"23",X"0D",X"C2",X"A5",X"14",X"CD",X"CF",X"14",X"C9",X"DD",X"E5",X"FD",X"E1",X"2E",X"1C",X"FD",
		X"70",X"00",X"FD",X"19",X"2D",X"C2",X"BF",X"14",X"DD",X"23",X"25",X"C2",X"B9",X"14",X"C9",X"DD",
		X"21",X"67",X"80",X"DD",X"36",X"00",X"01",X"DD",X"36",X"20",X"1E",X"DD",X"36",X"40",X"19",X"DD",
		X"21",X"E7",X"82",X"DD",X"36",X"00",X"02",X"DD",X"36",X"20",X"1E",X"DD",X"36",X"40",X"19",X"06",
		X"03",X"3A",X"52",X"9A",X"CB",X"47",X"CC",X"7C",X"0D",X"DD",X"21",X"67",X"88",X"FD",X"21",X"E7",
		X"8A",X"DD",X"70",X"00",X"DD",X"70",X"20",X"DD",X"70",X"40",X"FD",X"70",X"00",X"FD",X"70",X"20",
		X"FD",X"70",X"40",X"C9",X"21",X"44",X"80",X"06",X"7F",X"0E",X"10",X"11",X"64",X"03",X"70",X"23",
		X"1B",X"7B",X"B2",X"C2",X"1E",X"15",X"21",X"44",X"88",X"11",X"64",X"03",X"71",X"23",X"1B",X"7B",
		X"B2",X"C2",X"2C",X"15",X"DD",X"21",X"40",X"84",X"06",X"7A",X"0E",X"00",X"26",X"0B",X"11",X"20",
		X"00",X"CD",X"B9",X"14",X"DD",X"21",X"40",X"8C",X"41",X"26",X"0B",X"11",X"20",X"00",X"CD",X"B9",
		X"14",X"DD",X"21",X"4B",X"84",X"06",X"7F",X"26",X"11",X"11",X"20",X"00",X"CD",X"B9",X"14",X"DD",
		X"21",X"4B",X"8C",X"26",X"11",X"06",X"10",X"CD",X"B9",X"14",X"CD",X"CF",X"14",X"C9",X"DD",X"21",
		X"20",X"9A",X"CD",X"A1",X"15",X"CD",X"65",X"16",X"CD",X"D7",X"16",X"DD",X"7E",X"00",X"A7",X"C8",
		X"DD",X"7E",X"05",X"A7",X"C0",X"CD",X"7F",X"17",X"DD",X"7E",X"06",X"A7",X"C0",X"CD",X"4B",X"18",
		X"CD",X"8A",X"18",X"3A",X"59",X"9A",X"DD",X"86",X"02",X"DD",X"A6",X"01",X"C0",X"CD",X"D5",X"18",
		X"C9",X"DD",X"7E",X"05",X"A7",X"C2",X"F4",X"15",X"0E",X"0B",X"FD",X"21",X"00",X"98",X"CD",X"C4",
		X"15",X"11",X"10",X"00",X"FD",X"19",X"0D",X"C2",X"AE",X"15",X"DD",X"7E",X"05",X"A7",X"C8",X"DD",
		X"36",X"06",X"3F",X"C9",X"FD",X"7E",X"00",X"A7",X"C8",X"21",X"E4",X"45",X"FD",X"46",X"04",X"3E",
		X"E8",X"96",X"B8",X"D0",X"23",X"3E",X"E8",X"86",X"B8",X"D8",X"23",X"FD",X"46",X"03",X"DD",X"7E",
		X"03",X"57",X"96",X"B8",X"D0",X"23",X"7A",X"86",X"B8",X"D8",X"DD",X"36",X"05",X"FF",X"21",X"16",
		X"9C",X"CB",X"C6",X"C9",X"3A",X"59",X"9A",X"DD",X"86",X"02",X"DD",X"A6",X"01",X"C0",X"21",X"16",
		X"9C",X"CB",X"C6",X"DD",X"7E",X"06",X"FE",X"30",X"CA",X"50",X"16",X"D2",X"1B",X"16",X"FE",X"20",
		X"CA",X"57",X"16",X"FE",X"10",X"CA",X"5E",X"16",X"C3",X"1F",X"16",X"DD",X"36",X"0F",X"E3",X"DD",
		X"56",X"03",X"1E",X"E8",X"DD",X"66",X"0F",X"2E",X"19",X"3E",X"00",X"CD",X"62",X"32",X"DD",X"35",
		X"06",X"C0",X"3E",X"FF",X"32",X"51",X"9A",X"DD",X"36",X"05",X"00",X"DD",X"36",X"00",X"00",X"DD",
		X"36",X"07",X"00",X"DD",X"36",X"09",X"00",X"DD",X"36",X"0F",X"D3",X"DD",X"36",X"12",X"00",X"C9",
		X"DD",X"36",X"0F",X"E7",X"C3",X"1F",X"16",X"DD",X"36",X"0F",X"EB",X"C3",X"1F",X"16",X"DD",X"36",
		X"0F",X"EF",X"C3",X"1F",X"16",X"DD",X"7E",X"07",X"A7",X"C8",X"3A",X"59",X"9A",X"E6",X"01",X"C0",
		X"DD",X"7E",X"08",X"D6",X"02",X"DD",X"77",X"08",X"06",X"05",X"CD",X"8A",X"16",X"DD",X"7E",X"08",
		X"C6",X"08",X"06",X"06",X"CD",X"8A",X"16",X"C3",X"97",X"16",X"DD",X"56",X"1E",X"5F",X"26",X"0B",
		X"2E",X"00",X"78",X"CD",X"0E",X"32",X"C9",X"FD",X"21",X"25",X"46",X"06",X"00",X"0E",X"06",X"DD",
		X"66",X"1E",X"DD",X"6E",X"08",X"CD",X"B7",X"16",X"78",X"A7",X"C2",X"C8",X"16",X"0D",X"C8",X"11",
		X"03",X"00",X"FD",X"19",X"C3",X"A5",X"16",X"7D",X"FD",X"BE",X"00",X"D0",X"7C",X"FD",X"BE",X"01",
		X"D8",X"FD",X"BE",X"02",X"D0",X"06",X"FF",X"C9",X"DD",X"36",X"07",X"00",X"3E",X"05",X"CD",X"5D",
		X"18",X"3E",X"06",X"CD",X"5D",X"18",X"C9",X"DD",X"7E",X"09",X"A7",X"C8",X"3A",X"59",X"9A",X"E6",
		X"01",X"C0",X"DD",X"7E",X"1D",X"A7",X"C2",X"5F",X"17",X"DD",X"7E",X"0C",X"A7",X"C2",X"01",X"17",
		X"DD",X"7E",X"0B",X"DD",X"BE",X"11",X"DA",X"01",X"17",X"D6",X"02",X"DD",X"77",X"0B",X"C3",X"37",
		X"17",X"DD",X"66",X"0E",X"DD",X"6E",X"0D",X"E5",X"FD",X"E1",X"DD",X"7E",X"0C",X"A7",X"CA",X"22",
		X"17",X"11",X"02",X"00",X"FD",X"19",X"3D",X"C2",X"11",X"17",X"FD",X"7E",X"00",X"FE",X"80",X"CA",
		X"47",X"17",X"DD",X"7E",X"0B",X"FD",X"86",X"00",X"DD",X"77",X"0B",X"FD",X"7E",X"01",X"DD",X"86",
		X"0A",X"DD",X"77",X"0A",X"DD",X"34",X"0C",X"DD",X"56",X"0A",X"DD",X"5E",X"0B",X"26",X"0C",X"2E",
		X"00",X"3E",X"04",X"CD",X"0E",X"32",X"C9",X"DD",X"36",X"1D",X"FF",X"DD",X"36",X"0C",X"03",X"DD",
		X"56",X"0A",X"DD",X"5E",X"0B",X"26",X"0A",X"2E",X"00",X"3E",X"04",X"CD",X"0E",X"32",X"C9",X"DD",
		X"35",X"0C",X"C0",X"DD",X"36",X"09",X"00",X"DD",X"36",X"1D",X"00",X"16",X"08",X"DD",X"72",X"0A",
		X"1E",X"10",X"DD",X"73",X"0B",X"26",X"0F",X"2E",X"00",X"3E",X"04",X"CD",X"0E",X"32",X"C9",X"DD",
		X"7E",X"06",X"FE",X"FF",X"C0",X"3A",X"59",X"9A",X"DD",X"86",X"02",X"DD",X"A6",X"01",X"C0",X"FD",
		X"21",X"CE",X"4F",X"06",X"00",X"DD",X"7E",X"12",X"D6",X"03",X"A7",X"CA",X"A6",X"17",X"FD",X"23",
		X"FD",X"23",X"3D",X"C2",X"9E",X"17",X"FD",X"6E",X"00",X"FD",X"66",X"01",X"E5",X"FD",X"E1",X"FD",
		X"6E",X"0D",X"FD",X"66",X"0E",X"FD",X"7E",X"0C",X"A7",X"CA",X"C4",X"17",X"11",X"04",X"00",X"19",
		X"3D",X"C2",X"BC",X"17",X"7E",X"FE",X"80",X"CA",X"1B",X"18",X"FD",X"86",X"04",X"FD",X"77",X"04",
		X"5F",X"23",X"7E",X"FD",X"86",X"03",X"FD",X"77",X"03",X"57",X"23",X"46",X"23",X"4E",X"C5",X"E1",
		X"FD",X"74",X"0F",X"DD",X"7E",X"12",X"CD",X"62",X"32",X"FD",X"34",X"0C",X"FD",X"7E",X"0B",X"FE",
		X"10",X"C2",X"00",X"18",X"DD",X"7E",X"03",X"D6",X"03",X"FD",X"BE",X"03",X"D0",X"C3",X"09",X"18",
		X"DD",X"7E",X"03",X"C6",X"03",X"FD",X"BE",X"03",X"D8",X"DD",X"7E",X"03",X"D6",X"02",X"57",X"1E",
		X"DE",X"26",X"09",X"2E",X"00",X"3E",X"06",X"CD",X"0E",X"32",X"C9",X"DD",X"36",X"06",X"3F",X"DD",
		X"36",X"05",X"FF",X"21",X"16",X"9C",X"CB",X"C6",X"16",X"F8",X"1E",X"F0",X"26",X"FF",X"FD",X"74",
		X"0F",X"2E",X"0F",X"DD",X"7E",X"12",X"CD",X"62",X"32",X"3E",X"06",X"CD",X"5D",X"18",X"FD",X"36",
		X"05",X"FF",X"FD",X"36",X"06",X"1E",X"FD",X"36",X"1E",X"00",X"C9",X"DD",X"7E",X"07",X"A7",X"C0",
		X"3E",X"05",X"CD",X"5D",X"18",X"3E",X"06",X"CD",X"5D",X"18",X"C3",X"6C",X"18",X"16",X"08",X"1E",
		X"10",X"DD",X"73",X"08",X"26",X"0F",X"2E",X"00",X"CD",X"0E",X"32",X"C9",X"3A",X"57",X"9A",X"A7",
		X"C0",X"3A",X"58",X"9A",X"A7",X"C8",X"DD",X"36",X"07",X"FF",X"DD",X"36",X"08",X"DA",X"DD",X"7E",
		X"03",X"DD",X"77",X"1E",X"21",X"16",X"9C",X"CB",X"D6",X"C9",X"DD",X"7E",X"09",X"A7",X"C0",X"16",
		X"08",X"1E",X"10",X"DD",X"73",X"0B",X"26",X"0F",X"2E",X"00",X"3E",X"04",X"CD",X"0E",X"32",X"3A",
		X"55",X"9A",X"A7",X"C0",X"3A",X"56",X"9A",X"A7",X"C8",X"DD",X"36",X"09",X"FF",X"DD",X"7E",X"03",
		X"DD",X"77",X"0A",X"C6",X"10",X"DD",X"77",X"10",X"DD",X"7E",X"04",X"DD",X"77",X"11",X"DD",X"36",
		X"0B",X"DA",X"DD",X"36",X"0C",X"00",X"21",X"FC",X"45",X"DD",X"75",X"0D",X"DD",X"74",X"0E",X"21",
		X"16",X"9C",X"CB",X"CE",X"C9",X"3A",X"54",X"9A",X"CB",X"47",X"C2",X"E9",X"18",X"CB",X"4F",X"C2",
		X"03",X"19",X"DD",X"36",X"0F",X"D3",X"C3",X"2F",X"19",X"DD",X"7E",X"03",X"C6",X"01",X"FE",X"DE",
		X"D2",X"FC",X"18",X"DD",X"77",X"03",X"CD",X"1D",X"19",X"C3",X"2F",X"19",X"DD",X"36",X"03",X"DE",
		X"C3",X"2F",X"19",X"DD",X"7E",X"03",X"D6",X"01",X"FE",X"1C",X"DA",X"16",X"19",X"DD",X"77",X"03",
		X"CD",X"1D",X"19",X"C3",X"2F",X"19",X"DD",X"36",X"03",X"1C",X"C3",X"2F",X"19",X"DD",X"7E",X"0F",
		X"FE",X"D3",X"CA",X"2A",X"19",X"DD",X"36",X"0F",X"D3",X"C9",X"DD",X"36",X"0F",X"D7",X"C9",X"DD",
		X"56",X"03",X"1E",X"E8",X"DD",X"66",X"0F",X"2E",X"1A",X"3E",X"00",X"CD",X"62",X"32",X"3A",X"54",
		X"9A",X"CB",X"67",X"C2",X"4E",X"19",X"CB",X"6F",X"C2",X"65",X"19",X"C3",X"7C",X"19",X"DD",X"7E",
		X"04",X"D6",X"01",X"FE",X"22",X"DA",X"5E",X"19",X"DD",X"77",X"04",X"C3",X"7C",X"19",X"DD",X"36",
		X"04",X"22",X"C3",X"7C",X"19",X"DD",X"7E",X"04",X"C6",X"01",X"FE",X"96",X"D2",X"75",X"19",X"DD",
		X"77",X"04",X"C3",X"7C",X"19",X"DD",X"36",X"04",X"96",X"C3",X"7C",X"19",X"DD",X"7E",X"03",X"C6",
		X"10",X"57",X"DD",X"5E",X"04",X"CD",X"B5",X"31",X"C9",X"DD",X"21",X"B0",X"98",X"CD",X"B4",X"19",
		X"DD",X"21",X"D0",X"98",X"CD",X"B4",X"19",X"DD",X"21",X"F0",X"98",X"CD",X"B4",X"19",X"DD",X"21",
		X"10",X"99",X"CD",X"B4",X"19",X"DD",X"21",X"30",X"99",X"CD",X"B4",X"19",X"C9",X"CD",X"89",X"19",
		X"CD",X"77",X"1F",X"C9",X"CD",X"CD",X"19",X"DD",X"7E",X"00",X"A7",X"C8",X"CD",X"43",X"1A",X"3A",
		X"59",X"9A",X"DD",X"86",X"02",X"DD",X"A6",X"01",X"C0",X"CD",X"25",X"1B",X"C9",X"DD",X"7E",X"07",
		X"A7",X"C8",X"DD",X"6E",X"08",X"DD",X"66",X"09",X"E5",X"FD",X"E1",X"FD",X"7E",X"00",X"A7",X"C8",
		X"3A",X"59",X"9A",X"FD",X"86",X"02",X"FD",X"A6",X"01",X"C0",X"FD",X"7E",X"04",X"C6",X"08",X"FD",
		X"77",X"04",X"FE",X"F0",X"D2",X"04",X"1A",X"DD",X"7E",X"12",X"A7",X"C2",X"15",X"1A",X"3E",X"FF",
		X"CD",X"21",X"1A",X"C9",X"AF",X"CD",X"21",X"1A",X"FD",X"E5",X"E1",X"3E",X"0D",X"CD",X"70",X"20",
		X"DD",X"36",X"07",X"00",X"C9",X"FD",X"7E",X"03",X"FD",X"86",X"08",X"FD",X"77",X"03",X"C3",X"FE",
		X"19",X"A7",X"CA",X"36",X"1A",X"FD",X"7E",X"0E",X"FD",X"56",X"03",X"FD",X"5E",X"04",X"26",X"0D",
		X"2E",X"00",X"CD",X"0E",X"32",X"C9",X"FD",X"7E",X"0E",X"11",X"F0",X"08",X"21",X"FF",X"FF",X"CD",
		X"0E",X"32",X"C9",X"DD",X"7E",X"05",X"A7",X"C2",X"96",X"1A",X"CD",X"6E",X"31",X"A7",X"C8",X"FD",
		X"21",X"20",X"9A",X"DD",X"7E",X"03",X"C6",X"06",X"FD",X"96",X"0A",X"DA",X"64",X"1A",X"FE",X"10",
		X"D0",X"C3",X"67",X"1A",X"FE",X"10",X"D0",X"DD",X"7E",X"04",X"C6",X"00",X"FD",X"96",X"0B",X"DA",
		X"78",X"1A",X"FE",X"10",X"D0",X"C3",X"7D",X"1A",X"ED",X"44",X"FE",X"10",X"D0",X"DD",X"36",X"05",
		X"FF",X"DD",X"36",X"06",X"30",X"21",X"16",X"9C",X"CB",X"DE",X"3E",X"00",X"32",X"29",X"9A",X"CD",
		X"60",X"20",X"CD",X"80",X"20",X"C9",X"DD",X"7E",X"06",X"A7",X"CA",X"E3",X"1A",X"FE",X"10",X"CA",
		X"A7",X"1A",X"3D",X"DD",X"77",X"06",X"C9",X"DD",X"7E",X"11",X"A7",X"C2",X"C5",X"1A",X"DD",X"56",
		X"03",X"DD",X"5E",X"04",X"CD",X"A6",X"33",X"DD",X"7E",X"06",X"3D",X"DD",X"77",X"06",X"21",X"50",
		X"00",X"22",X"5B",X"9A",X"C9",X"DD",X"56",X"03",X"DD",X"5E",X"04",X"26",X"EF",X"2E",X"19",X"DD",
		X"7E",X"1F",X"CD",X"62",X"32",X"DD",X"35",X"06",X"DD",X"36",X"0C",X"40",X"21",X"00",X"02",X"22",
		X"5B",X"9A",X"C9",X"DD",X"7E",X"11",X"A7",X"C2",X"00",X"1B",X"C3",X"91",X"1B",X"DD",X"56",X"03",
		X"DD",X"5E",X"04",X"21",X"F0",X"08",X"DD",X"7E",X"1F",X"CD",X"62",X"32",X"CD",X"09",X"1F",X"C9",
		X"DD",X"7E",X"0C",X"A7",X"CA",X"ED",X"1A",X"FE",X"20",X"CA",X"11",X"1B",X"3D",X"DD",X"77",X"0C",
		X"C9",X"DD",X"56",X"03",X"DD",X"5E",X"04",X"26",X"F3",X"2E",X"10",X"DD",X"7E",X"1F",X"CD",X"62",
		X"32",X"DD",X"35",X"0C",X"C9",X"DD",X"7E",X"05",X"A7",X"C0",X"CD",X"3E",X"1B",X"DD",X"7E",X"11",
		X"A7",X"C2",X"48",X"1B",X"CD",X"66",X"1B",X"CD",X"9E",X"1B",X"CD",X"14",X"1C",X"C9",X"3A",X"8B",
		X"9C",X"FE",X"0E",X"D8",X"CD",X"80",X"20",X"C9",X"DD",X"7E",X"12",X"A7",X"C2",X"59",X"1B",X"CD",
		X"53",X"1D",X"CD",X"14",X"1C",X"CD",X"70",X"1C",X"C9",X"CD",X"E7",X"1D",X"CD",X"47",X"1F",X"CD",
		X"14",X"1C",X"CD",X"62",X"1E",X"C9",X"DD",X"7E",X"03",X"C6",X"02",X"DD",X"77",X"03",X"FE",X"F0",
		X"D2",X"8E",X"1B",X"DD",X"7E",X"12",X"A7",X"C2",X"84",X"1B",X"DD",X"56",X"03",X"DD",X"5E",X"04",
		X"CD",X"BC",X"33",X"C9",X"DD",X"56",X"03",X"DD",X"5E",X"04",X"CD",X"82",X"34",X"C9",X"CD",X"57",
		X"20",X"DD",X"56",X"03",X"DD",X"5E",X"04",X"CD",X"B0",X"33",X"CD",X"09",X"1F",X"C9",X"FD",X"21",
		X"B0",X"98",X"0E",X"05",X"11",X"20",X"00",X"3A",X"53",X"9A",X"06",X"06",X"FE",X"02",X"DA",X"B3",
		X"1B",X"06",X"08",X"FD",X"7E",X"00",X"A7",X"C4",X"FE",X"1B",X"FD",X"19",X"0D",X"C2",X"B3",X"1B",
		X"78",X"A7",X"C8",X"3A",X"23",X"9A",X"DD",X"96",X"03",X"D8",X"FE",X"10",X"D0",X"DD",X"36",X"0B",
		X"00",X"DD",X"36",X"14",X"01",X"DD",X"56",X"03",X"DD",X"5E",X"04",X"C5",X"CD",X"B0",X"33",X"C1",
		X"DD",X"36",X"11",X"FF",X"CB",X"48",X"C2",X"F4",X"1B",X"CB",X"50",X"C2",X"F9",X"1B",X"3E",X"03",
		X"DD",X"77",X"1F",X"C9",X"DD",X"36",X"1F",X"01",X"C9",X"DD",X"36",X"1F",X"02",X"C9",X"FD",X"7E",
		X"1F",X"FE",X"01",X"CA",X"0E",X"1C",X"FE",X"02",X"CA",X"11",X"1C",X"CB",X"98",X"C9",X"CB",X"88",
		X"C9",X"CB",X"90",X"C9",X"3A",X"59",X"9A",X"DD",X"86",X"02",X"DD",X"46",X"01",X"CB",X"20",X"CB",
		X"C0",X"A0",X"C0",X"DD",X"7E",X"13",X"3C",X"DD",X"77",X"13",X"FE",X"60",X"D8",X"DD",X"36",X"13",
		X"00",X"16",X"09",X"FD",X"21",X"00",X"98",X"01",X"10",X"00",X"FD",X"7E",X"00",X"A7",X"CA",X"48",
		X"1C",X"FD",X"09",X"15",X"C2",X"3A",X"1C",X"C9",X"FD",X"36",X"00",X"FF",X"DD",X"7E",X"03",X"DD",
		X"46",X"04",X"FD",X"77",X"03",X"FD",X"70",X"04",X"FD",X"36",X"06",X"00",X"FD",X"36",X"05",X"00",
		X"FD",X"77",X"08",X"FD",X"36",X"09",X"E8",X"FD",X"36",X"0A",X"00",X"FD",X"36",X"07",X"02",X"C9",
		X"DD",X"4E",X"0D",X"DD",X"46",X"0E",X"CB",X"21",X"CB",X"10",X"CB",X"21",X"CB",X"10",X"DD",X"5E",
		X"14",X"FD",X"21",X"A3",X"40",X"16",X"00",X"CB",X"23",X"CB",X"12",X"FD",X"19",X"FD",X"5E",X"00",
		X"FD",X"56",X"01",X"D5",X"FD",X"E1",X"FD",X"09",X"FD",X"7E",X"00",X"FE",X"80",X"CA",X"E5",X"1C",
		X"DD",X"86",X"03",X"DD",X"77",X"03",X"57",X"FD",X"7E",X"01",X"DD",X"86",X"04",X"DD",X"77",X"04",
		X"5F",X"FD",X"66",X"02",X"FD",X"6E",X"03",X"DD",X"7E",X"1F",X"CD",X"62",X"32",X"DD",X"7E",X"03",
		X"FE",X"F0",X"D2",X"F4",X"1E",X"FE",X"10",X"DA",X"F4",X"1E",X"DD",X"7E",X"04",X"FE",X"10",X"DA",
		X"F4",X"1E",X"FE",X"F0",X"D2",X"F4",X"1E",X"DD",X"6E",X"0D",X"DD",X"66",X"0E",X"23",X"DD",X"75",
		X"0D",X"DD",X"74",X"0E",X"C9",X"3E",X"01",X"DD",X"46",X"0A",X"DD",X"34",X"0A",X"B8",X"DA",X"10",
		X"1D",X"FD",X"46",X"01",X"ED",X"5F",X"CB",X"47",X"CA",X"44",X"1D",X"78",X"CB",X"3F",X"CB",X"3F",
		X"CB",X"3F",X"CB",X"3F",X"DD",X"77",X"14",X"DD",X"36",X"0D",X"00",X"DD",X"36",X"0E",X"00",X"C9",
		X"DD",X"7E",X"14",X"FE",X"00",X"CA",X"2A",X"1D",X"FE",X"04",X"CA",X"37",X"1D",X"FE",X"06",X"CA",
		X"2A",X"1D",X"FE",X"07",X"CA",X"37",X"1D",X"C3",X"F1",X"1C",X"DD",X"36",X"14",X"06",X"DD",X"36",
		X"0D",X"00",X"DD",X"36",X"0E",X"00",X"C9",X"DD",X"36",X"14",X"07",X"DD",X"36",X"0D",X"00",X"DD",
		X"36",X"0E",X"00",X"C9",X"78",X"E6",X"0F",X"DD",X"77",X"14",X"DD",X"36",X"0D",X"00",X"DD",X"36",
		X"0E",X"00",X"C9",X"DD",X"7E",X"14",X"FE",X"03",X"CA",X"61",X"1D",X"FE",X"01",X"CA",X"61",X"1D",
		X"C9",X"DD",X"7E",X"0D",X"FE",X"05",X"C0",X"3A",X"23",X"9A",X"DD",X"96",X"03",X"DA",X"76",X"1D",
		X"FE",X"20",X"D0",X"C3",X"31",X"1C",X"ED",X"44",X"FE",X"20",X"D0",X"C3",X"31",X"1C",X"FD",X"21",
		X"00",X"98",X"01",X"10",X"00",X"2E",X"09",X"FD",X"7E",X"00",X"A7",X"CA",X"95",X"1D",X"FD",X"09",
		X"2D",X"C2",X"87",X"1D",X"C9",X"FD",X"36",X"00",X"FF",X"DD",X"36",X"07",X"FF",X"DD",X"7E",X"03",
		X"FD",X"77",X"03",X"DD",X"7E",X"04",X"FD",X"77",X"04",X"FD",X"36",X"05",X"00",X"FD",X"36",X"06",
		X"00",X"FD",X"36",X"07",X"01",X"FD",X"E5",X"E1",X"DD",X"75",X"08",X"DD",X"74",X"09",X"3E",X"E8",
		X"FD",X"77",X"09",X"3A",X"23",X"9A",X"DD",X"96",X"03",X"DA",X"D8",X"1D",X"CB",X"3F",X"CB",X"3F",
		X"CB",X"3F",X"CB",X"3F",X"FD",X"77",X"08",X"C9",X"ED",X"44",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",
		X"CB",X"3F",X"2F",X"FD",X"77",X"08",X"C9",X"DD",X"7E",X"0B",X"E6",X"F0",X"C2",X"32",X"1E",X"3A",
		X"52",X"9A",X"DD",X"BE",X"0A",X"D8",X"3A",X"23",X"9A",X"47",X"DD",X"7E",X"0B",X"E6",X"0F",X"C2",
		X"1A",X"1E",X"DD",X"7E",X"03",X"90",X"D8",X"FE",X"20",X"D8",X"DD",X"36",X"0B",X"F0",X"DD",X"36",
		X"0C",X"08",X"DD",X"34",X"0A",X"DD",X"36",X"16",X"00",X"C9",X"78",X"DD",X"96",X"03",X"D8",X"FE",
		X"20",X"D8",X"DD",X"36",X"0B",X"FF",X"DD",X"36",X"0C",X"08",X"DD",X"34",X"0A",X"DD",X"36",X"16",
		X"00",X"C9",X"CD",X"57",X"1E",X"DD",X"56",X"03",X"DD",X"5E",X"04",X"26",X"BF",X"2E",X"11",X"DD",
		X"7E",X"1F",X"CD",X"62",X"32",X"DD",X"7E",X"0C",X"3D",X"DD",X"77",X"0C",X"C0",X"DD",X"7E",X"0B",
		X"2F",X"E6",X"0F",X"DD",X"77",X"0B",X"C9",X"DD",X"7E",X"04",X"3C",X"FE",X"90",X"D0",X"DD",X"77",
		X"04",X"C9",X"DD",X"7E",X"0B",X"E6",X"F0",X"C0",X"DD",X"7E",X"07",X"A7",X"C2",X"CF",X"1E",X"DD",
		X"34",X"0C",X"DD",X"7E",X"0B",X"E6",X"0F",X"C2",X"8D",X"1E",X"CD",X"B0",X"1E",X"DD",X"7E",X"03",
		X"C6",X"02",X"DD",X"77",X"03",X"FE",X"F0",X"D2",X"F4",X"1E",X"C3",X"A0",X"1E",X"CD",X"C2",X"1E",
		X"DD",X"7E",X"03",X"D6",X"02",X"DD",X"77",X"03",X"FE",X"10",X"DA",X"F4",X"1E",X"C3",X"A0",X"1E",
		X"DD",X"56",X"03",X"DD",X"5E",X"04",X"DD",X"7E",X"1F",X"CD",X"62",X"32",X"DD",X"34",X"0C",X"C9",
		X"DD",X"7E",X"0C",X"CB",X"47",X"CA",X"BD",X"1E",X"26",X"BB",X"2E",X"11",X"C9",X"26",X"B7",X"2E",
		X"11",X"C9",X"DD",X"7E",X"0C",X"CB",X"47",X"CA",X"EF",X"1E",X"26",X"C7",X"2E",X"11",X"C9",X"DD",
		X"7E",X"0B",X"E6",X"0F",X"C2",X"E8",X"1E",X"26",X"CB",X"2E",X"11",X"DD",X"56",X"03",X"DD",X"5E",
		X"04",X"DD",X"7E",X"1F",X"CD",X"62",X"32",X"C9",X"26",X"CF",X"2E",X"11",X"C3",X"DB",X"1E",X"26",
		X"C3",X"2E",X"11",X"C9",X"16",X"08",X"1E",X"FF",X"26",X"FF",X"2E",X"FF",X"DD",X"7E",X"1F",X"CD",
		X"62",X"32",X"CD",X"09",X"1F",X"CD",X"57",X"20",X"C9",X"DD",X"46",X"07",X"DD",X"4E",X"08",X"DD",
		X"56",X"09",X"DD",X"5E",X"12",X"DD",X"E5",X"E1",X"23",X"23",X"23",X"3E",X"1D",X"36",X"00",X"23",
		X"3D",X"C2",X"1D",X"1F",X"DD",X"36",X"00",X"00",X"DD",X"70",X"07",X"DD",X"71",X"08",X"DD",X"72",
		X"09",X"DD",X"73",X"12",X"C9",X"DD",X"7E",X"07",X"A7",X"C8",X"DD",X"6E",X"08",X"DD",X"66",X"09",
		X"E5",X"FD",X"E1",X"CD",X"04",X"1A",X"C9",X"DD",X"7E",X"07",X"A7",X"C0",X"DD",X"7E",X"16",X"3C",
		X"DD",X"77",X"16",X"FE",X"04",X"D0",X"DD",X"7E",X"0B",X"47",X"E6",X"F0",X"C0",X"78",X"E6",X"0F",
		X"CA",X"6D",X"1F",X"3A",X"23",X"9A",X"DD",X"BE",X"03",X"D0",X"C3",X"7E",X"1D",X"3A",X"23",X"9A",
		X"DD",X"BE",X"03",X"D8",X"C3",X"7E",X"1D",X"3A",X"59",X"9A",X"E6",X"3F",X"C0",X"3A",X"89",X"9C",
		X"FE",X"08",X"D2",X"8A",X"1F",X"3C",X"32",X"89",X"9C",X"C9",X"AF",X"32",X"89",X"9C",X"3A",X"8B",
		X"9C",X"47",X"3A",X"8C",X"9C",X"4F",X"CD",X"C5",X"1F",X"90",X"D8",X"C8",X"91",X"C8",X"D8",X"3A",
		X"8A",X"9C",X"FE",X"09",X"D2",X"B8",X"1F",X"4F",X"3C",X"32",X"8A",X"9C",X"06",X"00",X"21",X"4F",
		X"3F",X"09",X"5E",X"16",X"10",X"C3",X"D0",X"1F",X"AF",X"32",X"8A",X"9C",X"3A",X"4F",X"3F",X"5F",
		X"16",X"10",X"C3",X"D0",X"1F",X"3A",X"FF",X"9B",X"CB",X"77",X"3E",X"10",X"C8",X"3E",X"18",X"C9",
		X"3A",X"53",X"9A",X"FE",X"00",X"CA",X"E5",X"1F",X"FE",X"01",X"CA",X"0F",X"20",X"FE",X"02",X"CA",
		X"14",X"20",X"C3",X"39",X"20",X"26",X"00",X"DD",X"21",X"B0",X"98",X"01",X"20",X"00",X"2E",X"05",
		X"DD",X"7E",X"00",X"A7",X"CA",X"FE",X"1F",X"DD",X"09",X"2D",X"C2",X"F0",X"1F",X"C9",X"DD",X"36",
		X"00",X"FF",X"DD",X"72",X"03",X"DD",X"73",X"04",X"DD",X"74",X"12",X"CD",X"4F",X"20",X"C9",X"26",
		X"FF",X"C3",X"E7",X"1F",X"DD",X"21",X"F0",X"99",X"01",X"10",X"00",X"2E",X"03",X"DD",X"7E",X"00",
		X"A7",X"CA",X"2B",X"20",X"DD",X"09",X"2D",X"C2",X"1D",X"20",X"C9",X"DD",X"36",X"00",X"FF",X"DD",
		X"72",X"03",X"DD",X"73",X"04",X"CD",X"4F",X"20",X"C9",X"ED",X"5F",X"E6",X"03",X"FE",X"00",X"CA",
		X"E5",X"1F",X"FE",X"01",X"CA",X"0F",X"20",X"FE",X"02",X"CA",X"14",X"20",X"C3",X"14",X"20",X"3A",
		X"8C",X"9C",X"3C",X"32",X"8C",X"9C",X"C9",X"3A",X"8C",X"9C",X"3D",X"F8",X"32",X"8C",X"9C",X"C9",
		X"3A",X"8B",X"9C",X"3C",X"32",X"8B",X"9C",X"3A",X"8C",X"9C",X"3D",X"F8",X"32",X"8C",X"9C",X"C9",
		X"36",X"00",X"23",X"23",X"23",X"0E",X"00",X"D6",X"03",X"71",X"23",X"3D",X"C2",X"79",X"20",X"C9",
		X"3A",X"53",X"9A",X"FE",X"02",X"D2",X"9F",X"20",X"FD",X"21",X"50",X"99",X"01",X"20",X"00",X"1E",
		X"05",X"FD",X"7E",X"00",X"A7",X"CA",X"AB",X"20",X"FD",X"09",X"1D",X"C2",X"91",X"20",X"C9",X"FD",
		X"21",X"70",X"99",X"01",X"20",X"00",X"1E",X"04",X"C3",X"91",X"20",X"FD",X"36",X"00",X"FF",X"DD",
		X"7E",X"03",X"FD",X"77",X"03",X"DD",X"7E",X"04",X"FD",X"77",X"04",X"AF",X"FD",X"77",X"05",X"FD",
		X"77",X"06",X"FD",X"77",X"0C",X"FD",X"77",X"17",X"FD",X"77",X"18",X"FD",X"36",X"1E",X"00",X"C9",
		X"DD",X"21",X"F0",X"97",X"11",X"10",X"00",X"DD",X"19",X"DD",X"E5",X"E1",X"01",X"90",X"98",X"ED",
		X"42",X"C8",X"CD",X"E8",X"20",X"C3",X"D4",X"20",X"DD",X"7E",X"00",X"A7",X"C8",X"DD",X"7E",X"07",
		X"FE",X"02",X"C0",X"CD",X"11",X"21",X"DD",X"7E",X"05",X"A7",X"C0",X"DD",X"7E",X"00",X"A7",X"C8",
		X"3A",X"59",X"9A",X"DD",X"86",X"02",X"DD",X"A6",X"01",X"C0",X"CD",X"1D",X"21",X"CD",X"58",X"21",
		X"C9",X"DD",X"E5",X"FD",X"E1",X"DD",X"7E",X"05",X"A7",X"C2",X"3F",X"31",X"C9",X"DD",X"7E",X"04",
		X"FE",X"D4",X"D0",X"C6",X"02",X"DD",X"77",X"04",X"5F",X"DD",X"56",X"03",X"26",X"0D",X"2E",X"00",
		X"DD",X"7E",X"0E",X"CD",X"0E",X"32",X"DD",X"7E",X"04",X"FE",X"D4",X"D8",X"DD",X"7E",X"03",X"FE",
		X"80",X"D2",X"4A",X"21",X"21",X"4D",X"46",X"C3",X"4D",X"21",X"21",X"37",X"46",X"DD",X"75",X"0B",
		X"DD",X"74",X"0C",X"DD",X"36",X"0A",X"00",X"C9",X"DD",X"7E",X"04",X"FE",X"D4",X"D8",X"FE",X"E9",
		X"DA",X"7C",X"21",X"DD",X"36",X"05",X"FF",X"DD",X"56",X"03",X"DD",X"5E",X"04",X"26",X"0A",X"2E",
		X"00",X"DD",X"7E",X"0E",X"CD",X"0E",X"32",X"DD",X"36",X"06",X"08",X"C9",X"DD",X"66",X"0C",X"DD",
		X"6E",X"0B",X"E5",X"FD",X"E1",X"DD",X"7E",X"0A",X"A7",X"CA",X"95",X"21",X"11",X"02",X"00",X"FD",
		X"19",X"3D",X"C2",X"8C",X"21",X"FD",X"7E",X"01",X"DD",X"86",X"03",X"DD",X"77",X"03",X"57",X"FD",
		X"7E",X"00",X"DD",X"86",X"04",X"DD",X"77",X"04",X"5F",X"26",X"0D",X"2E",X"00",X"DD",X"7E",X"0E",
		X"CD",X"0E",X"32",X"DD",X"34",X"0A",X"C9",X"DD",X"21",X"E0",X"99",X"11",X"10",X"00",X"DD",X"19",
		X"DD",X"E5",X"E1",X"01",X"20",X"9A",X"ED",X"42",X"C8",X"CD",X"CF",X"21",X"C3",X"BB",X"21",X"DD",
		X"7E",X"00",X"A7",X"C8",X"CD",X"F1",X"21",X"3A",X"59",X"9A",X"DD",X"86",X"02",X"DD",X"A6",X"01",
		X"C0",X"CD",X"69",X"22",X"CD",X"99",X"22",X"CD",X"22",X"23",X"CD",X"91",X"23",X"CD",X"18",X"24",
		X"C9",X"DD",X"7E",X"05",X"A7",X"C2",X"49",X"22",X"CD",X"6E",X"31",X"A7",X"C8",X"21",X"EC",X"45",
		X"FD",X"21",X"20",X"9A",X"DD",X"7E",X"04",X"47",X"96",X"FD",X"BE",X"11",X"D0",X"23",X"78",X"86",
		X"FD",X"BE",X"11",X"D8",X"23",X"DD",X"7E",X"03",X"47",X"96",X"FD",X"BE",X"10",X"D0",X"23",X"78",
		X"86",X"FD",X"BE",X"10",X"D8",X"DD",X"36",X"05",X"FF",X"DD",X"36",X"06",X"07",X"FD",X"36",X"09",
		X"00",X"21",X"50",X"00",X"22",X"5B",X"9A",X"CD",X"60",X"20",X"DD",X"56",X"03",X"DD",X"5E",X"04",
		X"CD",X"A6",X"33",X"21",X"16",X"9C",X"CB",X"DE",X"C9",X"3A",X"59",X"9A",X"DD",X"86",X"02",X"DD",
		X"A6",X"01",X"C0",X"DD",X"35",X"06",X"C0",X"DD",X"36",X"00",X"00",X"DD",X"36",X"05",X"00",X"DD",
		X"56",X"03",X"DD",X"5E",X"04",X"CD",X"B0",X"33",X"C9",X"DD",X"7E",X"05",X"A7",X"C0",X"DD",X"7E",
		X"00",X"A7",X"C8",X"DD",X"7E",X"03",X"C6",X"02",X"FE",X"FC",X"D2",X"88",X"22",X"DD",X"77",X"03",
		X"57",X"DD",X"5E",X"04",X"CD",X"9C",X"33",X"C9",X"DD",X"36",X"00",X"00",X"DD",X"56",X"03",X"DD",
		X"5E",X"04",X"CD",X"B0",X"33",X"CD",X"57",X"20",X"C9",X"DD",X"7E",X"08",X"A7",X"C2",X"E7",X"22",
		X"DD",X"7E",X"05",X"A7",X"C0",X"FD",X"21",X"F0",X"97",X"11",X"10",X"00",X"0E",X"08",X"FD",X"19",
		X"FD",X"7E",X"00",X"A7",X"CA",X"BC",X"22",X"0D",X"C2",X"AE",X"22",X"C9",X"FD",X"36",X"00",X"FF",
		X"FD",X"36",X"07",X"08",X"FD",X"36",X"05",X"00",X"FD",X"36",X"06",X"00",X"DD",X"7E",X"03",X"FD",
		X"77",X"03",X"DD",X"7E",X"04",X"C6",X"0A",X"FD",X"77",X"04",X"DD",X"34",X"08",X"FD",X"E5",X"E1",
		X"DD",X"74",X"0A",X"DD",X"75",X"09",X"C9",X"DD",X"34",X"08",X"DD",X"7E",X"08",X"FE",X"1E",X"CA",
		X"18",X"23",X"FE",X"06",X"CA",X"1D",X"23",X"D0",X"DD",X"66",X"0A",X"DD",X"6E",X"09",X"E5",X"FD",
		X"E1",X"FD",X"7E",X"04",X"C6",X"02",X"FD",X"77",X"04",X"5F",X"FD",X"56",X"03",X"26",X"0B",X"2E",
		X"00",X"FD",X"7E",X"0E",X"CD",X"0E",X"32",X"C9",X"DD",X"36",X"08",X"00",X"C9",X"DD",X"36",X"07",
		X"FF",X"C9",X"DD",X"7E",X"07",X"A7",X"C8",X"FD",X"21",X"80",X"98",X"11",X"10",X"00",X"0E",X"02",
		X"FD",X"19",X"FD",X"7E",X"00",X"A7",X"CA",X"3E",X"23",X"0D",X"C2",X"30",X"23",X"C9",X"FD",X"E5",
		X"D1",X"DD",X"66",X"0A",X"DD",X"6E",X"09",X"E5",X"FD",X"E1",X"FD",X"46",X"03",X"FD",X"4E",X"04",
		X"FD",X"36",X"00",X"00",X"FD",X"36",X"07",X"00",X"D5",X"FD",X"E1",X"FD",X"36",X"00",X"FF",X"FD",
		X"70",X"03",X"FD",X"71",X"04",X"FD",X"36",X"05",X"00",X"FD",X"21",X"20",X"9A",X"FD",X"7E",X"03",
		X"D5",X"FD",X"E1",X"FD",X"77",X"08",X"DD",X"36",X"07",X"00",X"E5",X"FD",X"E1",X"16",X"08",X"1E",
		X"08",X"26",X"00",X"2E",X"00",X"FD",X"7E",X"0E",X"CD",X"0E",X"32",X"21",X"16",X"9C",X"CB",X"E6",
		X"C9",X"DD",X"7E",X"07",X"A7",X"C8",X"3A",X"53",X"9A",X"FE",X"03",X"C2",X"A7",X"23",X"FD",X"21",
		X"50",X"99",X"0E",X"04",X"C3",X"AD",X"23",X"FD",X"21",X"30",X"99",X"0E",X"05",X"11",X"20",X"00",
		X"3A",X"52",X"9A",X"FE",X"03",X"D2",X"B9",X"23",X"0D",X"FD",X"19",X"FD",X"7E",X"00",X"A7",X"CA",
		X"C7",X"23",X"0D",X"C2",X"B9",X"23",X"C9",X"FD",X"E5",X"D1",X"DD",X"66",X"0A",X"DD",X"6E",X"09",
		X"E5",X"FD",X"E1",X"FD",X"46",X"03",X"FD",X"4E",X"04",X"FD",X"36",X"00",X"00",X"D5",X"FD",X"E1",
		X"FD",X"36",X"00",X"FF",X"FD",X"70",X"03",X"FD",X"71",X"04",X"FD",X"36",X"05",X"00",X"FD",X"36",
		X"06",X"00",X"FD",X"36",X"0C",X"00",X"FD",X"36",X"17",X"00",X"FD",X"36",X"18",X"00",X"FD",X"36",
		X"1E",X"00",X"DD",X"36",X"07",X"00",X"E5",X"FD",X"E1",X"16",X"08",X"1E",X"08",X"26",X"00",X"2E",
		X"00",X"FD",X"7E",X"0E",X"CD",X"0E",X"32",X"C9",X"DD",X"7E",X"07",X"A7",X"C8",X"DD",X"66",X"0A",
		X"DD",X"6E",X"09",X"E5",X"FD",X"E1",X"FD",X"36",X"05",X"00",X"FD",X"36",X"06",X"00",X"FD",X"36",
		X"0A",X"00",X"FD",X"36",X"07",X"02",X"DD",X"36",X"07",X"00",X"C9",X"DD",X"21",X"80",X"98",X"11",
		X"10",X"00",X"DD",X"19",X"DD",X"E5",X"E1",X"01",X"B0",X"98",X"ED",X"42",X"C8",X"CD",X"53",X"24",
		X"C3",X"3F",X"24",X"DD",X"7E",X"00",X"A7",X"C8",X"CD",X"76",X"24",X"DD",X"7E",X"05",X"A7",X"C0",
		X"3A",X"59",X"9A",X"DD",X"86",X"02",X"DD",X"A6",X"01",X"C0",X"DD",X"7E",X"00",X"A7",X"C8",X"CD",
		X"2D",X"25",X"CD",X"41",X"25",X"C9",X"DD",X"7E",X"05",X"A7",X"C2",X"E6",X"24",X"FD",X"21",X"20",
		X"9A",X"CD",X"6E",X"31",X"A7",X"CA",X"A2",X"24",X"21",X"E8",X"45",X"FD",X"56",X"10",X"FD",X"5E",
		X"11",X"CD",X"BA",X"24",X"DD",X"7E",X"05",X"A7",X"CA",X"A2",X"24",X"FD",X"36",X"09",X"00",X"C3",
		X"D7",X"24",X"21",X"E8",X"45",X"FD",X"56",X"1E",X"FD",X"5E",X"08",X"CD",X"BA",X"24",X"DD",X"7E",
		X"05",X"A7",X"C8",X"FD",X"36",X"07",X"00",X"C3",X"D7",X"24",X"DD",X"7E",X"04",X"96",X"BB",X"D0",
		X"23",X"DD",X"7E",X"04",X"86",X"BB",X"D8",X"23",X"DD",X"7E",X"03",X"96",X"BA",X"D0",X"23",X"86",
		X"BA",X"D8",X"DD",X"36",X"05",X"FF",X"C9",X"DD",X"36",X"06",X"04",X"DD",X"36",X"07",X"05",X"21",
		X"00",X"02",X"22",X"5B",X"9A",X"C9",X"3A",X"59",X"9A",X"DD",X"86",X"02",X"DD",X"A6",X"01",X"C0",
		X"DD",X"7E",X"06",X"A7",X"CA",X"02",X"25",X"26",X"EB",X"2E",X"19",X"CD",X"20",X"25",X"DD",X"35",
		X"06",X"C9",X"26",X"F3",X"2E",X"12",X"CD",X"20",X"25",X"DD",X"35",X"07",X"C0",X"DD",X"36",X"00",
		X"00",X"26",X"FF",X"2E",X"0F",X"16",X"08",X"1E",X"10",X"DD",X"7E",X"0E",X"CD",X"62",X"32",X"C9",
		X"DD",X"56",X"03",X"DD",X"5E",X"04",X"DD",X"7E",X"0E",X"CD",X"62",X"32",X"C9",X"DD",X"7E",X"04",
		X"FE",X"70",X"D8",X"FE",X"A8",X"D0",X"FD",X"21",X"20",X"9A",X"FD",X"7E",X"03",X"DD",X"77",X"08",
		X"C9",X"DD",X"7E",X"03",X"FE",X"10",X"DA",X"58",X"25",X"FE",X"F0",X"D2",X"58",X"25",X"DD",X"7E",
		X"04",X"C6",X"02",X"FE",X"E8",X"DA",X"75",X"25",X"DD",X"36",X"00",X"00",X"DD",X"36",X"05",X"00",
		X"26",X"FF",X"2E",X"0F",X"16",X"08",X"DD",X"72",X"03",X"1E",X"10",X"DD",X"73",X"04",X"DD",X"7E",
		X"0E",X"CD",X"62",X"32",X"C9",X"DD",X"77",X"04",X"3E",X"E8",X"DD",X"96",X"04",X"47",X"CB",X"28",
		X"DD",X"7E",X"08",X"DD",X"BE",X"03",X"CA",X"AA",X"25",X"DD",X"96",X"03",X"CB",X"7F",X"C2",X"9E",
		X"25",X"B8",X"DA",X"98",X"25",X"DD",X"34",X"03",X"DD",X"34",X"03",X"C3",X"AA",X"25",X"ED",X"44",
		X"B8",X"DA",X"A7",X"25",X"DD",X"35",X"03",X"DD",X"35",X"03",X"DD",X"7E",X"0F",X"FE",X"DB",X"CA",
		X"B9",X"25",X"DD",X"36",X"0F",X"DB",X"C3",X"BD",X"25",X"DD",X"36",X"0F",X"DF",X"DD",X"56",X"03",
		X"DD",X"5E",X"04",X"DD",X"66",X"0F",X"2E",X"14",X"DD",X"7E",X"0E",X"CD",X"62",X"32",X"C9",X"DD",
		X"21",X"30",X"99",X"11",X"20",X"00",X"DD",X"19",X"DD",X"E5",X"E1",X"01",X"F0",X"99",X"ED",X"42",
		X"C8",X"CD",X"E7",X"25",X"C3",X"D3",X"25",X"DD",X"7E",X"1E",X"FE",X"00",X"C0",X"DD",X"7E",X"00",
		X"A7",X"C8",X"DD",X"36",X"01",X"0F",X"CD",X"1A",X"26",X"CD",X"4B",X"26",X"DD",X"7E",X"05",X"A7",
		X"C0",X"3A",X"59",X"9A",X"DD",X"86",X"02",X"DD",X"A6",X"01",X"C0",X"DD",X"7E",X"00",X"A7",X"C8",
		X"DD",X"34",X"06",X"CD",X"C7",X"26",X"CD",X"9F",X"27",X"C9",X"DD",X"7E",X"04",X"FE",X"60",X"D8",
		X"DD",X"7E",X"17",X"A7",X"C0",X"FD",X"21",X"30",X"99",X"11",X"20",X"00",X"0E",X"05",X"FD",X"19",
		X"0D",X"CA",X"42",X"26",X"FD",X"7E",X"00",X"A7",X"CA",X"2E",X"26",X"FD",X"36",X"0A",X"FF",X"C3",
		X"2E",X"26",X"DD",X"36",X"0A",X"00",X"DD",X"36",X"17",X"FF",X"C9",X"DD",X"7E",X"05",X"A7",X"C2",
		X"98",X"26",X"CD",X"6E",X"31",X"A7",X"C8",X"FD",X"21",X"20",X"9A",X"21",X"F0",X"45",X"DD",X"7E",
		X"04",X"96",X"FD",X"BE",X"11",X"D0",X"23",X"DD",X"7E",X"04",X"86",X"FD",X"BE",X"11",X"D8",X"23",
		X"DD",X"7E",X"03",X"96",X"FD",X"BE",X"10",X"D0",X"23",X"DD",X"7E",X"03",X"86",X"FD",X"BE",X"10",
		X"D8",X"DD",X"36",X"05",X"FF",X"FD",X"36",X"09",X"00",X"21",X"00",X"03",X"22",X"5B",X"9A",X"DD",
		X"36",X"06",X"04",X"DD",X"36",X"0F",X"F7",X"C9",X"3A",X"59",X"9A",X"DD",X"86",X"02",X"DD",X"A6",
		X"01",X"C0",X"DD",X"56",X"03",X"DD",X"5E",X"04",X"DD",X"66",X"0F",X"2E",X"12",X"DD",X"7E",X"1F",
		X"CD",X"62",X"32",X"DD",X"35",X"06",X"C0",X"DD",X"36",X"00",X"00",X"CD",X"F6",X"2F",X"DD",X"36",
		X"17",X"00",X"DD",X"36",X"18",X"00",X"C9",X"DD",X"66",X"0E",X"DD",X"6E",X"0D",X"E5",X"FD",X"E1",
		X"DD",X"7E",X"0C",X"A7",X"CA",X"0C",X"27",X"11",X"04",X"00",X"FD",X"19",X"3D",X"C2",X"DA",X"26",
		X"FD",X"7E",X"00",X"FE",X"80",X"CA",X"0C",X"27",X"DD",X"7E",X"03",X"FD",X"86",X"01",X"DD",X"77",
		X"03",X"57",X"DD",X"7E",X"04",X"FD",X"86",X"00",X"DD",X"77",X"04",X"5F",X"FD",X"66",X"02",X"FD",
		X"6E",X"03",X"DD",X"7E",X"1F",X"CD",X"62",X"32",X"DD",X"34",X"0C",X"C9",X"DD",X"7E",X"18",X"A7",
		X"CA",X"3A",X"27",X"21",X"63",X"46",X"C3",X"94",X"27",X"ED",X"5F",X"E6",X"7F",X"47",X"3A",X"59",
		X"9A",X"80",X"47",X"3A",X"52",X"9A",X"17",X"17",X"4F",X"3E",X"3F",X"91",X"B8",X"DA",X"3A",X"27",
		X"21",X"63",X"46",X"DD",X"36",X"18",X"FF",X"C3",X"94",X"27",X"21",X"E9",X"46",X"DD",X"7E",X"03",
		X"BE",X"DA",X"58",X"27",X"23",X"BE",X"DA",X"6C",X"27",X"23",X"BE",X"DA",X"80",X"27",X"23",X"3E",
		X"FF",X"BE",X"CA",X"58",X"27",X"C3",X"3D",X"27",X"DD",X"7E",X"06",X"FE",X"08",X"D2",X"66",X"27",
		X"21",X"63",X"46",X"C3",X"94",X"27",X"21",X"8E",X"46",X"C3",X"94",X"27",X"DD",X"7E",X"06",X"FE",
		X"08",X"D2",X"7A",X"27",X"21",X"7C",X"46",X"C3",X"94",X"27",X"21",X"AF",X"46",X"C3",X"94",X"27",
		X"DD",X"7E",X"06",X"FE",X"08",X"D2",X"8E",X"27",X"21",X"85",X"46",X"C3",X"94",X"27",X"21",X"CC",
		X"46",X"C3",X"94",X"27",X"DD",X"74",X"0E",X"DD",X"75",X"0D",X"DD",X"36",X"0C",X"01",X"C9",X"DD",
		X"7E",X"04",X"FE",X"A0",X"D8",X"DD",X"7E",X"18",X"A7",X"C2",X"E6",X"27",X"DD",X"36",X"01",X"0F",
		X"DD",X"56",X"03",X"1E",X"A0",X"DD",X"73",X"04",X"DD",X"36",X"06",X"00",X"DD",X"36",X"09",X"00",
		X"DD",X"36",X"0B",X"00",X"DD",X"36",X"0C",X"00",X"26",X"83",X"DD",X"74",X"0F",X"DD",X"36",X"15",
		X"00",X"DD",X"36",X"17",X"00",X"DD",X"36",X"18",X"00",X"DD",X"36",X"1E",X"FF",X"2E",X"12",X"DD",
		X"7E",X"1F",X"CD",X"62",X"32",X"C9",X"16",X"08",X"DD",X"72",X"03",X"1E",X"10",X"DD",X"73",X"04",
		X"26",X"FF",X"2E",X"0F",X"DD",X"7E",X"1F",X"CD",X"62",X"32",X"DD",X"36",X"00",X"00",X"DD",X"36",
		X"17",X"00",X"DD",X"36",X"18",X"00",X"DD",X"36",X"06",X"00",X"C9",X"3A",X"59",X"9A",X"E6",X"0F",
		X"C2",X"1F",X"28",X"3A",X"6D",X"99",X"3D",X"C2",X"1C",X"28",X"3E",X"8F",X"32",X"6D",X"99",X"DD",
		X"21",X"30",X"99",X"11",X"20",X"00",X"DD",X"19",X"DD",X"E5",X"E1",X"01",X"F0",X"99",X"ED",X"42",
		X"C8",X"CD",X"37",X"28",X"C3",X"23",X"28",X"CD",X"91",X"28",X"DD",X"7E",X"00",X"A7",X"C8",X"DD",
		X"7E",X"1E",X"FE",X"FF",X"C0",X"3A",X"26",X"9A",X"A7",X"C0",X"3A",X"25",X"9A",X"A7",X"C0",X"CD",
		X"AB",X"29",X"DD",X"7E",X"05",X"A7",X"C0",X"3A",X"6D",X"99",X"FE",X"8F",X"C2",X"63",X"28",X"DD",
		X"36",X"0A",X"FF",X"3A",X"59",X"9A",X"DD",X"86",X"02",X"DD",X"A6",X"01",X"C0",X"DD",X"7E",X"00",
		X"A7",X"C8",X"DD",X"7E",X"09",X"FE",X"00",X"CA",X"89",X"28",X"FE",X"20",X"CA",X"8D",X"28",X"CD",
		X"0A",X"2B",X"CD",X"65",X"2C",X"CD",X"FB",X"2C",X"C9",X"CD",X"78",X"2A",X"C9",X"CD",X"40",X"2E",
		X"C9",X"DD",X"7E",X"11",X"A7",X"C2",X"6F",X"29",X"DD",X"7E",X"07",X"A7",X"C8",X"DD",X"66",X"14",
		X"DD",X"6E",X"13",X"E5",X"FD",X"E1",X"FD",X"7E",X"05",X"A7",X"CA",X"BA",X"28",X"CD",X"3F",X"31",
		X"FD",X"7E",X"00",X"A7",X"C0",X"DD",X"36",X"07",X"00",X"C9",X"3A",X"59",X"9A",X"DD",X"86",X"02",
		X"E6",X"07",X"C0",X"FD",X"66",X"0C",X"FD",X"6E",X"0B",X"FD",X"7E",X"0A",X"A7",X"CA",X"DC",X"28",
		X"23",X"23",X"3D",X"C2",X"D0",X"28",X"7E",X"FE",X"80",X"CA",X"FD",X"28",X"FD",X"7E",X"04",X"86",
		X"FD",X"77",X"04",X"5F",X"23",X"FD",X"7E",X"03",X"86",X"FD",X"77",X"03",X"57",X"26",X"0B",X"2E",
		X"00",X"FD",X"7E",X"0E",X"CD",X"0E",X"32",X"FD",X"34",X"0A",X"C3",X"13",X"29",X"FD",X"7E",X"04",
		X"C6",X"03",X"FD",X"77",X"04",X"5F",X"FD",X"56",X"03",X"26",X"0B",X"2E",X"00",X"FD",X"7E",X"0E",
		X"CD",X"0E",X"32",X"FD",X"7E",X"04",X"FD",X"BE",X"09",X"D8",X"FD",X"7E",X"09",X"FE",X"E8",X"D2",
		X"56",X"29",X"21",X"40",X"9A",X"DD",X"5E",X"10",X"16",X"00",X"CB",X"23",X"1D",X"19",X"36",X"FF",
		X"DD",X"36",X"11",X"FF",X"DD",X"36",X"12",X"02",X"DD",X"56",X"10",X"CD",X"FB",X"36",X"FD",X"36",
		X"00",X"00",X"16",X"08",X"1E",X"10",X"26",X"00",X"2E",X"00",X"FD",X"7E",X"0E",X"CD",X"0E",X"32",
		X"21",X"16",X"9C",X"CB",X"DE",X"C9",X"FD",X"36",X"05",X"FF",X"FD",X"36",X"06",X"03",X"FD",X"56",
		X"03",X"FD",X"5E",X"04",X"26",X"0A",X"2E",X"00",X"FD",X"7E",X"0E",X"CD",X"0E",X"32",X"C9",X"DD",
		X"7E",X"11",X"FE",X"0F",X"CA",X"8A",X"29",X"DD",X"35",X"12",X"C0",X"DD",X"36",X"11",X"0F",X"DD",
		X"36",X"12",X"02",X"DD",X"56",X"10",X"CD",X"13",X"37",X"C9",X"DD",X"35",X"12",X"C0",X"DD",X"36",
		X"11",X"00",X"DD",X"56",X"10",X"CD",X"A6",X"36",X"21",X"40",X"9A",X"DD",X"5E",X"10",X"16",X"00",
		X"CB",X"23",X"1D",X"19",X"36",X"FF",X"DD",X"36",X"07",X"00",X"C9",X"DD",X"7E",X"05",X"A7",X"C2",
		X"0F",X"2A",X"DD",X"7E",X"09",X"FE",X"20",X"C2",X"2F",X"2A",X"3A",X"54",X"9A",X"A7",X"C8",X"DD",
		X"7E",X"04",X"FE",X"E6",X"D8",X"FD",X"21",X"20",X"9A",X"FD",X"7E",X"03",X"D6",X"10",X"DD",X"BE",
		X"03",X"D0",X"FD",X"7E",X"03",X"C6",X"10",X"DD",X"BE",X"03",X"D8",X"DD",X"36",X"05",X"FF",X"DD",
		X"36",X"06",X"50",X"21",X"00",X"03",X"22",X"5B",X"9A",X"DD",X"56",X"03",X"DD",X"5E",X"04",X"DD",
		X"7E",X"0B",X"FE",X"10",X"CA",X"FC",X"29",X"26",X"77",X"C3",X"FE",X"29",X"26",X"6B",X"2E",X"12",
		X"DD",X"75",X"0F",X"DD",X"7E",X"1F",X"CD",X"62",X"32",X"21",X"16",X"9C",X"CB",X"EE",X"C9",X"DD",
		X"35",X"06",X"C0",X"DD",X"36",X"00",X"00",X"DD",X"36",X"1E",X"00",X"DD",X"36",X"05",X"00",X"DD",
		X"36",X"09",X"00",X"DD",X"36",X"0C",X"00",X"DD",X"36",X"15",X"00",X"CD",X"F6",X"2F",X"C9",X"21",
		X"F4",X"45",X"FD",X"21",X"20",X"9A",X"FD",X"7E",X"07",X"A7",X"C8",X"DD",X"7E",X"04",X"96",X"FD",
		X"BE",X"08",X"D0",X"23",X"DD",X"7E",X"04",X"86",X"FD",X"BE",X"08",X"D8",X"23",X"DD",X"7E",X"03",
		X"96",X"FD",X"BE",X"1E",X"D0",X"23",X"DD",X"7E",X"03",X"86",X"FD",X"BE",X"1E",X"D8",X"FD",X"36",
		X"07",X"00",X"DD",X"7E",X"09",X"FE",X"12",X"C2",X"DB",X"29",X"21",X"00",X"03",X"22",X"5B",X"9A",
		X"21",X"16",X"9C",X"CB",X"EE",X"C3",X"13",X"2A",X"DD",X"7E",X"07",X"A7",X"C0",X"FD",X"21",X"87",
		X"47",X"11",X"03",X"00",X"0E",X"00",X"DD",X"7E",X"03",X"FD",X"BE",X"01",X"D2",X"9B",X"2A",X"FD",
		X"19",X"0C",X"79",X"FE",X"03",X"CA",X"9B",X"2A",X"C3",X"86",X"2A",X"79",X"A7",X"CA",X"DE",X"2A",
		X"DD",X"71",X"10",X"21",X"40",X"9A",X"5F",X"16",X"00",X"CB",X"23",X"1D",X"19",X"7E",X"A7",X"C2",
		X"DE",X"2A",X"DD",X"36",X"0B",X"10",X"3A",X"40",X"9A",X"FE",X"00",X"C2",X"DA",X"2A",X"CD",X"0B",
		X"30",X"A7",X"CA",X"C8",X"2A",X"CD",X"2A",X"30",X"DD",X"36",X"09",X"10",X"21",X"E8",X"47",X"DD",
		X"74",X"0E",X"DD",X"75",X"0D",X"DD",X"36",X"0C",X"00",X"C9",X"CD",X"2A",X"30",X"C9",X"0C",X"DD",
		X"71",X"10",X"DD",X"36",X"09",X"10",X"DD",X"36",X"0B",X"20",X"DD",X"7E",X"10",X"FE",X"04",X"CA",
		X"F8",X"2A",X"21",X"C7",X"47",X"C3",X"FF",X"2A",X"21",X"09",X"48",X"DD",X"36",X"0B",X"10",X"DD",
		X"74",X"0E",X"DD",X"75",X"0D",X"DD",X"36",X"0C",X"00",X"C9",X"DD",X"7E",X"09",X"FE",X"10",X"C0",
		X"DD",X"7E",X"07",X"A7",X"C0",X"FD",X"21",X"6F",X"47",X"11",X"03",X"00",X"0E",X"08",X"DD",X"7E",
		X"04",X"FD",X"BE",X"00",X"D2",X"36",X"2B",X"DD",X"7E",X"03",X"FD",X"BE",X"01",X"D2",X"36",X"2B",
		X"FD",X"BE",X"02",X"D2",X"3F",X"2B",X"FD",X"19",X"0D",X"C2",X"1E",X"2B",X"C3",X"6A",X"2B",X"21",
		X"40",X"9A",X"7E",X"FE",X"00",X"CA",X"56",X"2B",X"DD",X"5E",X"10",X"16",X"00",X"CB",X"23",X"1D",
		X"19",X"7E",X"A7",X"CA",X"5D",X"2B",X"CD",X"0B",X"30",X"A7",X"CA",X"6A",X"2B",X"DD",X"7E",X"15",
		X"FE",X"03",X"D2",X"6A",X"2B",X"CD",X"2A",X"30",X"A7",X"C8",X"DD",X"66",X"0E",X"DD",X"6E",X"0D",
		X"E5",X"FD",X"E1",X"11",X"04",X"00",X"DD",X"7E",X"0C",X"A7",X"CA",X"92",X"2B",X"FD",X"19",X"3D",
		X"C2",X"7D",X"2B",X"FD",X"7E",X"00",X"FE",X"80",X"C2",X"92",X"2B",X"DD",X"36",X"0C",X"00",X"C3",
		X"6A",X"2B",X"DD",X"7E",X"03",X"FD",X"86",X"01",X"57",X"DD",X"77",X"03",X"DD",X"7E",X"04",X"FD",
		X"86",X"00",X"5F",X"DD",X"77",X"04",X"FD",X"66",X"02",X"DD",X"74",X"0F",X"FD",X"6E",X"03",X"DD",
		X"7E",X"1F",X"CD",X"62",X"32",X"21",X"16",X"9C",X"CB",X"F6",X"DD",X"34",X"0C",X"FD",X"21",X"87",
		X"47",X"11",X"03",X"00",X"DD",X"4E",X"10",X"0D",X"CA",X"D0",X"2B",X"FD",X"19",X"C3",X"C7",X"2B",
		X"DD",X"7E",X"03",X"FD",X"BE",X"01",X"D0",X"FD",X"BE",X"02",X"D8",X"3A",X"40",X"9A",X"FE",X"00",
		X"C2",X"16",X"2C",X"21",X"40",X"9A",X"DD",X"5E",X"10",X"16",X"00",X"CB",X"23",X"1D",X"19",X"7E",
		X"A7",X"C2",X"16",X"2C",X"DD",X"7E",X"10",X"FE",X"06",X"CA",X"10",X"2C",X"DD",X"7E",X"0B",X"FE",
		X"10",X"CA",X"0A",X"2C",X"21",X"E3",X"48",X"C3",X"56",X"2C",X"21",X"9A",X"48",X"C3",X"56",X"2C",
		X"21",X"2C",X"49",X"C3",X"56",X"2C",X"DD",X"7E",X"10",X"FE",X"06",X"CA",X"53",X"2C",X"ED",X"5F",
		X"47",X"3A",X"59",X"9A",X"80",X"DD",X"86",X"02",X"EA",X"3F",X"2C",X"DD",X"7E",X"0B",X"FE",X"10",
		X"CA",X"39",X"2C",X"21",X"87",X"49",X"C3",X"56",X"2C",X"21",X"72",X"49",X"C3",X"56",X"2C",X"DD",
		X"7E",X"0B",X"FE",X"10",X"CA",X"4D",X"2C",X"21",X"9C",X"49",X"C3",X"56",X"2C",X"21",X"AD",X"49",
		X"C3",X"56",X"2C",X"21",X"5D",X"49",X"DD",X"74",X"0E",X"DD",X"75",X"0D",X"DD",X"36",X"0C",X"00",
		X"DD",X"36",X"09",X"11",X"C9",X"DD",X"7E",X"09",X"FE",X"11",X"C0",X"DD",X"36",X"15",X"00",X"21",
		X"40",X"9A",X"DD",X"5E",X"10",X"16",X"00",X"CB",X"23",X"19",X"7E",X"A7",X"CA",X"83",X"2C",X"DD",
		X"36",X"0A",X"FF",X"DD",X"66",X"0E",X"DD",X"6E",X"0D",X"11",X"04",X"00",X"DD",X"7E",X"0C",X"A7",
		X"CA",X"98",X"2C",X"19",X"3D",X"C2",X"93",X"2C",X"DD",X"7E",X"04",X"86",X"DD",X"77",X"04",X"5F",
		X"23",X"DD",X"7E",X"03",X"86",X"DD",X"77",X"03",X"57",X"23",X"46",X"23",X"4E",X"DD",X"70",X"0F",
		X"23",X"7E",X"FE",X"80",X"CA",X"C3",X"2C",X"C5",X"E1",X"DD",X"7E",X"1F",X"CD",X"62",X"32",X"DD",
		X"34",X"0C",X"C9",X"CD",X"F6",X"2F",X"21",X"40",X"9A",X"7E",X"FE",X"00",X"C2",X"E5",X"2C",X"DD",
		X"5E",X"10",X"16",X"00",X"CB",X"23",X"1D",X"19",X"7E",X"A7",X"C2",X"E5",X"2C",X"36",X"FF",X"DD",
		X"56",X"10",X"CD",X"A6",X"36",X"DD",X"36",X"09",X"12",X"21",X"40",X"9A",X"DD",X"5E",X"10",X"16",
		X"00",X"CB",X"23",X"19",X"36",X"FF",X"DD",X"36",X"06",X"10",X"C9",X"DD",X"7E",X"09",X"FE",X"12",
		X"C0",X"DD",X"7E",X"0A",X"A7",X"C2",X"65",X"2D",X"DD",X"35",X"06",X"C0",X"DD",X"7E",X"07",X"A7",
		X"C0",X"CD",X"0B",X"30",X"A7",X"CA",X"2C",X"2D",X"DD",X"7E",X"15",X"FE",X"03",X"D2",X"2C",X"2D",
		X"CD",X"2A",X"30",X"A7",X"CA",X"2C",X"2D",X"DD",X"36",X"06",X"10",X"C9",X"DD",X"7E",X"0F",X"FE",
		X"FF",X"CA",X"3A",X"2D",X"CD",X"F6",X"2F",X"C3",X"60",X"2D",X"DD",X"7E",X"10",X"21",X"A3",X"47",
		X"11",X"04",X"00",X"19",X"3D",X"C2",X"43",X"2D",X"5E",X"DD",X"73",X"04",X"23",X"56",X"DD",X"72",
		X"03",X"23",X"46",X"DD",X"70",X"0F",X"23",X"4E",X"C5",X"E1",X"DD",X"7E",X"1F",X"CD",X"62",X"32",
		X"DD",X"36",X"06",X"10",X"C9",X"DD",X"36",X"15",X"00",X"DD",X"7E",X"10",X"FE",X"06",X"DA",X"8E",
		X"2D",X"5F",X"FE",X"08",X"CA",X"00",X"2E",X"ED",X"5F",X"E6",X"7F",X"EA",X"8E",X"2D",X"21",X"40",
		X"9A",X"16",X"00",X"CB",X"23",X"19",X"36",X"00",X"23",X"7E",X"A7",X"C2",X"00",X"2E",X"21",X"68",
		X"4A",X"DD",X"7E",X"10",X"3D",X"CA",X"9D",X"2D",X"23",X"23",X"C3",X"94",X"2D",X"7E",X"DD",X"77",
		X"04",X"23",X"7E",X"DD",X"77",X"03",X"DD",X"7E",X"10",X"FE",X"03",X"CA",X"C2",X"2D",X"FE",X"04",
		X"CA",X"CC",X"2D",X"FE",X"05",X"CA",X"D6",X"2D",X"21",X"C7",X"47",X"DD",X"36",X"0B",X"20",X"C3",
		X"DD",X"2D",X"21",X"09",X"48",X"DD",X"36",X"0B",X"10",X"C3",X"DD",X"2D",X"21",X"E8",X"47",X"DD",
		X"36",X"0B",X"10",X"C3",X"DD",X"2D",X"21",X"E8",X"47",X"DD",X"36",X"0B",X"10",X"DD",X"74",X"0E",
		X"DD",X"75",X"0D",X"DD",X"36",X"0C",X"00",X"DD",X"36",X"09",X"10",X"21",X"40",X"9A",X"16",X"00",
		X"DD",X"5E",X"10",X"CB",X"23",X"19",X"36",X"00",X"DD",X"34",X"10",X"DD",X"36",X"0A",X"00",X"C9",
		X"DD",X"7E",X"10",X"FE",X"08",X"CA",X"12",X"2E",X"21",X"BE",X"49",X"DD",X"36",X"0B",X"20",X"C3",
		X"19",X"2E",X"21",X"E2",X"49",X"DD",X"36",X"0B",X"10",X"DD",X"74",X"0E",X"DD",X"75",X"0D",X"21",
		X"68",X"4A",X"DD",X"7E",X"10",X"3D",X"CA",X"2E",X"2E",X"23",X"23",X"C3",X"25",X"2E",X"7E",X"DD",
		X"77",X"04",X"23",X"7E",X"DD",X"77",X"03",X"DD",X"36",X"0C",X"00",X"DD",X"36",X"09",X"20",X"C9",
		X"DD",X"7E",X"04",X"FE",X"E8",X"DA",X"7F",X"2F",X"DD",X"66",X"0E",X"DD",X"6E",X"0D",X"11",X"04",
		X"00",X"DD",X"7E",X"0C",X"A7",X"CA",X"5D",X"2E",X"19",X"3D",X"C2",X"58",X"2E",X"DD",X"7E",X"04",
		X"86",X"DD",X"77",X"04",X"5F",X"23",X"DD",X"7E",X"03",X"86",X"DD",X"77",X"03",X"57",X"23",X"46",
		X"DD",X"70",X"0F",X"23",X"4E",X"C5",X"E1",X"DD",X"7E",X"1F",X"CD",X"62",X"32",X"21",X"16",X"9C",
		X"CB",X"F6",X"DD",X"34",X"0C",X"DD",X"7E",X"0B",X"FE",X"10",X"CA",X"98",X"2E",X"3A",X"54",X"9A",
		X"CB",X"47",X"C2",X"FA",X"2E",X"C3",X"A3",X"2E",X"3A",X"54",X"9A",X"CB",X"4F",X"C2",X"FA",X"2E",
		X"C3",X"BB",X"2E",X"DD",X"7E",X"03",X"FD",X"21",X"20",X"9A",X"FD",X"BE",X"03",X"DA",X"31",X"2F",
		X"D6",X"14",X"FD",X"BE",X"03",X"D2",X"31",X"2F",X"C3",X"D0",X"2E",X"DD",X"7E",X"03",X"FD",X"21",
		X"20",X"9A",X"FD",X"BE",X"03",X"D2",X"31",X"2F",X"C6",X"14",X"FD",X"BE",X"03",X"DA",X"31",X"2F",
		X"DD",X"36",X"01",X"0F",X"FD",X"36",X"06",X"FF",X"DD",X"7E",X"0B",X"FE",X"10",X"CA",X"E6",X"2E",
		X"21",X"06",X"4A",X"C3",X"E9",X"2E",X"21",X"37",X"4A",X"DD",X"74",X"0E",X"DD",X"75",X"0D",X"DD",
		X"36",X"0C",X"00",X"DD",X"7E",X"1F",X"FD",X"77",X"12",X"C9",X"DD",X"7E",X"0B",X"FE",X"10",X"CA",
		X"0C",X"2F",X"DD",X"36",X"0B",X"10",X"21",X"E8",X"47",X"C3",X"13",X"2F",X"DD",X"36",X"0B",X"20",
		X"21",X"C7",X"47",X"DD",X"74",X"0E",X"DD",X"75",X"0D",X"DD",X"7E",X"01",X"FE",X"0F",X"CA",X"28",
		X"2F",X"DD",X"36",X"01",X"0F",X"C3",X"2C",X"2F",X"DD",X"36",X"01",X"03",X"DD",X"36",X"0C",X"00",
		X"C9",X"DD",X"7E",X"03",X"FE",X"E6",X"D2",X"6A",X"2F",X"FE",X"1B",X"DA",X"6A",X"2F",X"DD",X"66",
		X"0E",X"DD",X"6E",X"0D",X"11",X"04",X"00",X"DD",X"7E",X"0C",X"A7",X"C8",X"19",X"3D",X"C2",X"4C",
		X"2F",X"19",X"7E",X"FE",X"80",X"C0",X"DD",X"7E",X"0B",X"FE",X"10",X"CA",X"64",X"2F",X"21",X"C7",
		X"47",X"C3",X"74",X"2F",X"21",X"E8",X"47",X"C3",X"74",X"2F",X"3A",X"54",X"9A",X"A7",X"CA",X"FA",
		X"2E",X"21",X"91",X"48",X"DD",X"74",X"0E",X"DD",X"75",X"0D",X"DD",X"36",X"0C",X"00",X"C9",X"DD",
		X"66",X"0E",X"DD",X"6E",X"0D",X"E5",X"FD",X"E1",X"11",X"04",X"00",X"DD",X"7E",X"0C",X"A7",X"CA",
		X"98",X"2F",X"FD",X"19",X"3D",X"C2",X"92",X"2F",X"DD",X"7E",X"03",X"FD",X"86",X"01",X"57",X"DD",
		X"77",X"03",X"DD",X"7E",X"04",X"FD",X"86",X"00",X"5F",X"DD",X"77",X"04",X"FD",X"66",X"02",X"DD",
		X"74",X"0F",X"FD",X"6E",X"03",X"DD",X"7E",X"1F",X"CD",X"62",X"32",X"21",X"16",X"9C",X"CB",X"F6",
		X"DD",X"34",X"0C",X"DD",X"7E",X"04",X"FE",X"E8",X"D8",X"DD",X"7E",X"03",X"FD",X"21",X"20",X"9A",
		X"FD",X"BE",X"03",X"DA",X"E0",X"2F",X"DD",X"36",X"0B",X"20",X"21",X"C7",X"47",X"C3",X"E7",X"2F",
		X"DD",X"36",X"0B",X"10",X"21",X"E8",X"47",X"DD",X"74",X"0E",X"DD",X"75",X"0D",X"DD",X"36",X"0C",
		X"00",X"DD",X"36",X"01",X"03",X"C9",X"16",X"08",X"1E",X"10",X"DD",X"73",X"04",X"26",X"FF",X"DD",
		X"74",X"0F",X"2E",X"0F",X"DD",X"7E",X"1F",X"CD",X"62",X"32",X"C9",X"FD",X"21",X"20",X"9A",X"DD",
		X"7E",X"03",X"C6",X"20",X"FD",X"BE",X"03",X"DA",X"28",X"30",X"DD",X"7E",X"03",X"D6",X"20",X"FD",
		X"BE",X"03",X"D2",X"28",X"30",X"3E",X"FF",X"C9",X"AF",X"C9",X"FD",X"21",X"00",X"98",X"11",X"10",
		X"00",X"FD",X"7E",X"00",X"A7",X"CA",X"4A",X"30",X"FD",X"19",X"FD",X"E5",X"E1",X"01",X"90",X"98",
		X"ED",X"42",X"CA",X"48",X"30",X"C3",X"31",X"30",X"AF",X"C9",X"DD",X"34",X"15",X"FD",X"36",X"00",
		X"FF",X"FD",X"36",X"05",X"00",X"FD",X"36",X"06",X"00",X"FD",X"36",X"07",X"04",X"FD",X"36",X"0A",
		X"00",X"DD",X"36",X"07",X"FF",X"FD",X"E5",X"E1",X"DD",X"74",X"14",X"DD",X"75",X"13",X"DD",X"7E",
		X"09",X"FE",X"12",X"CA",X"E8",X"30",X"DD",X"56",X"03",X"DD",X"5E",X"04",X"26",X"67",X"2E",X"12",
		X"DD",X"7E",X"1F",X"CD",X"62",X"32",X"DD",X"7E",X"03",X"D6",X"04",X"FD",X"77",X"03",X"DD",X"7E",
		X"04",X"D6",X"06",X"FD",X"77",X"04",X"21",X"40",X"9A",X"7E",X"FE",X"00",X"CA",X"C2",X"30",X"DD",
		X"5E",X"10",X"16",X"00",X"CB",X"23",X"1D",X"19",X"7E",X"A7",X"C2",X"C2",X"30",X"DD",X"7E",X"10",
		X"21",X"9F",X"47",X"3D",X"CA",X"BB",X"30",X"23",X"C3",X"B3",X"30",X"7E",X"FD",X"77",X"09",X"C3",
		X"C6",X"30",X"FD",X"36",X"09",X"EB",X"DD",X"7E",X"10",X"FE",X"06",X"CA",X"DC",X"30",X"DD",X"7E",
		X"0B",X"FE",X"10",X"C2",X"E2",X"30",X"21",X"31",X"47",X"C3",X"36",X"31",X"21",X"58",X"47",X"C3",
		X"36",X"31",X"21",X"F3",X"46",X"C3",X"36",X"31",X"DD",X"7E",X"10",X"21",X"A3",X"47",X"11",X"04",
		X"00",X"19",X"3D",X"C2",X"F1",X"30",X"7E",X"DD",X"77",X"04",X"5F",X"D6",X"08",X"FD",X"77",X"04",
		X"23",X"56",X"DD",X"72",X"03",X"FD",X"72",X"03",X"FD",X"36",X"09",X"EB",X"2E",X"12",X"DD",X"7E",
		X"10",X"3D",X"CB",X"4F",X"CA",X"28",X"31",X"26",X"2B",X"DD",X"74",X"0F",X"DD",X"7E",X"1F",X"CD",
		X"62",X"32",X"21",X"58",X"47",X"C3",X"36",X"31",X"26",X"33",X"DD",X"74",X"0F",X"DD",X"7E",X"1F",
		X"CD",X"62",X"32",X"21",X"1A",X"47",X"FD",X"74",X"0C",X"FD",X"75",X"0B",X"3E",X"FF",X"C9",X"3A",
		X"59",X"9A",X"DD",X"86",X"02",X"DD",X"A6",X"01",X"C0",X"FD",X"35",X"06",X"C0",X"FD",X"36",X"00",
		X"00",X"FD",X"36",X"05",X"00",X"FD",X"36",X"06",X"00",X"FD",X"36",X"07",X"00",X"FD",X"36",X"0A",
		X"00",X"11",X"F0",X"08",X"21",X"FF",X"FF",X"FD",X"7E",X"0E",X"CD",X"0E",X"32",X"C9",X"3A",X"29",
		X"9A",X"A7",X"C8",X"3A",X"3D",X"9A",X"A7",X"C0",X"FD",X"E5",X"FD",X"21",X"20",X"9A",X"21",X"F8",
		X"45",X"FD",X"7E",X"11",X"96",X"FD",X"BE",X"0B",X"D2",X"B1",X"31",X"23",X"FD",X"7E",X"11",X"86",
		X"FD",X"BE",X"0B",X"DA",X"B1",X"31",X"23",X"FD",X"7E",X"10",X"96",X"FD",X"BE",X"0A",X"D2",X"B1",
		X"31",X"23",X"FD",X"7E",X"10",X"86",X"FD",X"BE",X"0A",X"DA",X"B1",X"31",X"3E",X"FF",X"FD",X"E1",
		X"C9",X"AF",X"FD",X"E1",X"C9",X"DD",X"E5",X"FD",X"E5",X"DD",X"21",X"3C",X"4C",X"FD",X"21",X"0C",
		X"4F",X"3A",X"5D",X"9A",X"47",X"3A",X"00",X"9C",X"90",X"FE",X"01",X"C2",X"D6",X"31",X"3E",X"00",
		X"92",X"57",X"3E",X"00",X"93",X"5F",X"0E",X"04",X"DD",X"6E",X"04",X"DD",X"66",X"05",X"FD",X"7E",
		X"00",X"CB",X"DF",X"77",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"FD",X"7E",X"01",X"82",X"77",X"DD",
		X"6E",X"02",X"DD",X"66",X"03",X"FD",X"7E",X"02",X"83",X"77",X"C5",X"01",X"04",X"00",X"DD",X"09",
		X"DD",X"09",X"FD",X"09",X"C1",X"0D",X"C2",X"D8",X"31",X"FD",X"E1",X"DD",X"E1",X"C9",X"DD",X"E5",
		X"FD",X"E5",X"DD",X"21",X"3C",X"4C",X"4F",X"06",X"00",X"CB",X"21",X"CB",X"10",X"CB",X"21",X"CB",
		X"10",X"CB",X"21",X"CB",X"10",X"DD",X"09",X"3A",X"5D",X"9A",X"47",X"3A",X"00",X"9C",X"90",X"FE",
		X"01",X"CA",X"37",X"32",X"C3",X"3F",X"32",X"3E",X"00",X"92",X"57",X"3E",X"00",X"93",X"5F",X"DD",
		X"4E",X"00",X"DD",X"46",X"01",X"7A",X"D6",X"02",X"02",X"DD",X"4E",X"02",X"DD",X"46",X"03",X"7B",
		X"D6",X"02",X"02",X"DD",X"4E",X"04",X"DD",X"46",X"05",X"CB",X"DC",X"7C",X"02",X"FD",X"E1",X"DD",
		X"E1",X"C9",X"DD",X"E5",X"FD",X"E5",X"DD",X"21",X"FC",X"4B",X"4F",X"06",X"00",X"CB",X"21",X"CB",
		X"10",X"CB",X"21",X"CB",X"10",X"CB",X"21",X"CB",X"10",X"DD",X"09",X"3A",X"5D",X"9A",X"47",X"3A",
		X"00",X"9C",X"90",X"FE",X"01",X"CA",X"8B",X"32",X"C3",X"97",X"32",X"3E",X"00",X"92",X"57",X"3E",
		X"00",X"93",X"5F",X"7C",X"EE",X"02",X"67",X"DD",X"4E",X"00",X"DD",X"46",X"01",X"7A",X"D6",X"08",
		X"02",X"DD",X"4E",X"02",X"DD",X"46",X"03",X"7B",X"D6",X"08",X"02",X"DD",X"4E",X"04",X"DD",X"46",
		X"05",X"7C",X"02",X"DD",X"4E",X"06",X"DD",X"46",X"07",X"7D",X"02",X"FD",X"E1",X"DD",X"E1",X"C9",
		X"DD",X"E5",X"FD",X"E5",X"DD",X"2A",X"60",X"9A",X"7A",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"FE",
		X"1C",X"D4",X"94",X"33",X"06",X"00",X"D6",X"02",X"DC",X"99",X"33",X"4F",X"FD",X"21",X"1B",X"84",
		X"CB",X"21",X"CB",X"10",X"CB",X"21",X"CB",X"10",X"CB",X"21",X"CB",X"10",X"CB",X"21",X"CB",X"10",
		X"CB",X"21",X"CB",X"10",X"FD",X"09",X"7B",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"D6",X"04",X"4F",
		X"06",X"00",X"A7",X"FD",X"E5",X"E1",X"ED",X"42",X"E5",X"FD",X"E1",X"7A",X"E6",X"07",X"CB",X"3F",
		X"4F",X"06",X"00",X"21",X"00",X"00",X"C5",X"E1",X"CB",X"21",X"CB",X"10",X"CB",X"21",X"CB",X"10",
		X"CB",X"21",X"CB",X"10",X"CB",X"25",X"CB",X"14",X"09",X"E5",X"C1",X"DD",X"56",X"00",X"DD",X"5E",
		X"01",X"DD",X"09",X"01",X"20",X"00",X"2E",X"05",X"FD",X"E5",X"DD",X"7E",X"02",X"FD",X"77",X"00",
		X"FD",X"09",X"DD",X"23",X"2D",X"C2",X"3A",X"33",X"FD",X"E1",X"FD",X"E5",X"FD",X"2B",X"2E",X"05",
		X"DD",X"7E",X"02",X"FD",X"77",X"00",X"FD",X"09",X"DD",X"23",X"2D",X"C2",X"50",X"33",X"3A",X"52",
		X"9A",X"CB",X"47",X"CC",X"92",X"33",X"7A",X"FD",X"E1",X"01",X"00",X"08",X"FD",X"09",X"01",X"20",
		X"00",X"FD",X"E5",X"2E",X"05",X"FD",X"77",X"00",X"FD",X"09",X"2D",X"C2",X"75",X"33",X"2E",X"05",
		X"FD",X"E1",X"FD",X"2B",X"FD",X"77",X"00",X"FD",X"09",X"2D",X"C2",X"84",X"33",X"FD",X"E1",X"DD",
		X"E1",X"C9",X"53",X"C9",X"3E",X"1C",X"16",X"E0",X"C9",X"3E",X"00",X"C9",X"21",X"1C",X"4F",X"22",
		X"60",X"9A",X"CD",X"C0",X"32",X"C9",X"21",X"7A",X"4F",X"22",X"60",X"9A",X"CD",X"C0",X"32",X"C9",
		X"21",X"A4",X"4F",X"22",X"60",X"9A",X"CD",X"C0",X"32",X"C9",X"53",X"C9",X"DD",X"E5",X"FD",X"E5",
		X"DD",X"21",X"46",X"4F",X"7A",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"06",X"00",X"D6",X"02",X"DC",
		X"99",X"33",X"4F",X"CB",X"21",X"CB",X"10",X"CB",X"21",X"CB",X"10",X"CB",X"21",X"CB",X"10",X"CB",
		X"21",X"CB",X"10",X"CB",X"21",X"CB",X"10",X"FD",X"21",X"1B",X"84",X"FD",X"09",X"7B",X"CB",X"3F",
		X"CB",X"3F",X"CB",X"3F",X"D6",X"04",X"06",X"00",X"4F",X"A7",X"FD",X"E5",X"E1",X"ED",X"42",X"E5",
		X"FD",X"E1",X"7A",X"E6",X"07",X"CB",X"3F",X"4F",X"06",X"00",X"C5",X"E1",X"CB",X"21",X"CB",X"10",
		X"CB",X"21",X"CB",X"10",X"CB",X"25",X"CB",X"14",X"09",X"E5",X"C1",X"DD",X"56",X"00",X"DD",X"5E",
		X"01",X"DD",X"09",X"01",X"20",X"00",X"2E",X"03",X"FD",X"E5",X"DD",X"7E",X"02",X"FD",X"77",X"00",
		X"FD",X"09",X"DD",X"23",X"2D",X"C2",X"2A",X"34",X"FD",X"E1",X"FD",X"E5",X"FD",X"2B",X"2E",X"03",
		X"DD",X"7E",X"02",X"FD",X"77",X"00",X"FD",X"09",X"DD",X"23",X"2D",X"C2",X"40",X"34",X"3A",X"52",
		X"9A",X"CB",X"47",X"CC",X"BA",X"33",X"7A",X"FD",X"E1",X"01",X"00",X"08",X"FD",X"09",X"01",X"20",
		X"00",X"FD",X"E5",X"2E",X"03",X"FD",X"77",X"00",X"FD",X"09",X"2D",X"C2",X"65",X"34",X"FD",X"E1",
		X"FD",X"2B",X"2E",X"03",X"FD",X"77",X"00",X"FD",X"09",X"2D",X"C2",X"74",X"34",X"FD",X"E1",X"DD",
		X"E1",X"C9",X"DD",X"E5",X"FD",X"E5",X"DD",X"21",X"60",X"4F",X"7A",X"CB",X"3F",X"CB",X"3F",X"CB",
		X"3F",X"06",X"00",X"D6",X"02",X"DC",X"99",X"33",X"4F",X"CB",X"21",X"CB",X"10",X"CB",X"21",X"CB",
		X"10",X"CB",X"21",X"CB",X"10",X"CB",X"21",X"CB",X"10",X"CB",X"21",X"CB",X"10",X"FD",X"21",X"1B",
		X"84",X"FD",X"09",X"7B",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"D6",X"04",X"06",X"00",X"4F",X"A7",
		X"FD",X"E5",X"E1",X"ED",X"42",X"E5",X"FD",X"E1",X"7A",X"E6",X"07",X"CB",X"3F",X"4F",X"06",X"00",
		X"C5",X"E1",X"CB",X"21",X"CB",X"10",X"CB",X"21",X"CB",X"10",X"CB",X"25",X"CB",X"14",X"09",X"E5",
		X"C1",X"DD",X"56",X"00",X"DD",X"5E",X"01",X"DD",X"09",X"01",X"20",X"00",X"2E",X"03",X"FD",X"E5",
		X"DD",X"7E",X"02",X"FD",X"77",X"00",X"FD",X"09",X"DD",X"23",X"2D",X"C2",X"F0",X"34",X"FD",X"E1",
		X"FD",X"E5",X"FD",X"2B",X"2E",X"03",X"DD",X"7E",X"02",X"FD",X"77",X"00",X"FD",X"09",X"DD",X"23",
		X"2D",X"C2",X"06",X"35",X"3A",X"52",X"9A",X"CB",X"47",X"CC",X"BA",X"33",X"7A",X"FD",X"E1",X"01",
		X"00",X"08",X"FD",X"09",X"01",X"20",X"00",X"FD",X"E5",X"2E",X"03",X"FD",X"77",X"00",X"FD",X"09",
		X"2D",X"C2",X"2B",X"35",X"FD",X"E1",X"FD",X"2B",X"2E",X"03",X"FD",X"77",X"00",X"FD",X"09",X"2D",
		X"C2",X"3A",X"35",X"FD",X"E1",X"DD",X"E1",X"C9",X"DD",X"E5",X"FD",X"E5",X"15",X"5A",X"CB",X"23",
		X"16",X"00",X"DD",X"21",X"FC",X"4E",X"DD",X"19",X"DD",X"5E",X"00",X"DD",X"56",X"01",X"3A",X"5E",
		X"9A",X"4F",X"06",X"00",X"C5",X"E1",X"CB",X"21",X"CB",X"10",X"CB",X"21",X"CB",X"10",X"CB",X"21",
		X"CB",X"10",X"CB",X"21",X"CB",X"10",X"CB",X"21",X"CB",X"10",X"CB",X"25",X"CB",X"14",X"CB",X"25",
		X"CB",X"14",X"09",X"E5",X"C1",X"DD",X"21",X"BC",X"4C",X"DD",X"09",X"01",X"20",X"00",X"D5",X"FD",
		X"E1",X"2E",X"04",X"DD",X"7E",X"00",X"FD",X"77",X"00",X"FD",X"09",X"DD",X"23",X"2D",X"C2",X"93",
		X"35",X"D5",X"FD",X"E1",X"FD",X"2B",X"2E",X"04",X"DD",X"7E",X"00",X"FD",X"77",X"00",X"FD",X"09",
		X"DD",X"23",X"2D",X"C2",X"A8",X"35",X"D5",X"FD",X"E1",X"FD",X"2B",X"FD",X"2B",X"2E",X"04",X"DD",
		X"7E",X"00",X"FD",X"77",X"00",X"FD",X"09",X"DD",X"23",X"2D",X"C2",X"BF",X"35",X"D5",X"FD",X"E1",
		X"FD",X"2B",X"FD",X"2B",X"FD",X"2B",X"3A",X"52",X"9A",X"CB",X"47",X"CC",X"4B",X"36",X"D5",X"FD",
		X"E1",X"01",X"00",X"08",X"FD",X"09",X"01",X"20",X"00",X"2E",X"04",X"DD",X"7E",X"00",X"FD",X"77",
		X"00",X"FD",X"09",X"DD",X"23",X"2D",X"C2",X"EB",X"35",X"D5",X"FD",X"E1",X"01",X"00",X"08",X"FD",
		X"2B",X"FD",X"09",X"01",X"20",X"00",X"2E",X"04",X"DD",X"7E",X"00",X"FD",X"77",X"00",X"FD",X"09",
		X"DD",X"23",X"2D",X"C2",X"08",X"36",X"D5",X"FD",X"E1",X"01",X"00",X"08",X"FD",X"2B",X"FD",X"2B",
		X"FD",X"09",X"01",X"20",X"00",X"2E",X"04",X"DD",X"7E",X"00",X"FD",X"77",X"00",X"FD",X"09",X"DD",
		X"23",X"2D",X"C2",X"27",X"36",X"D5",X"FD",X"E1",X"01",X"00",X"08",X"FD",X"2B",X"FD",X"2B",X"FD",
		X"2B",X"FD",X"09",X"01",X"20",X"00",X"FD",X"E1",X"DD",X"E1",X"C9",X"01",X"0C",X"00",X"DD",X"09",
		X"C9",X"3A",X"40",X"9A",X"FE",X"00",X"CA",X"76",X"36",X"FE",X"01",X"CA",X"8E",X"36",X"7A",X"FE",
		X"04",X"DA",X"6D",X"36",X"3E",X"05",X"32",X"5E",X"9A",X"CD",X"48",X"35",X"C9",X"3E",X"04",X"32",
		X"5E",X"9A",X"CD",X"48",X"35",X"C9",X"7A",X"FE",X"04",X"DA",X"85",X"36",X"3E",X"01",X"32",X"5E",
		X"9A",X"CD",X"48",X"35",X"C9",X"3E",X"00",X"32",X"5E",X"9A",X"CD",X"48",X"35",X"C9",X"7A",X"FE",
		X"04",X"DA",X"9D",X"36",X"3E",X"09",X"32",X"5E",X"9A",X"CD",X"48",X"35",X"C9",X"3E",X"08",X"32",
		X"5E",X"9A",X"CD",X"48",X"35",X"C9",X"3A",X"40",X"9A",X"FE",X"00",X"CA",X"CB",X"36",X"FE",X"01",
		X"CA",X"E3",X"36",X"7A",X"FE",X"04",X"DA",X"C2",X"36",X"3E",X"07",X"32",X"5E",X"9A",X"CD",X"48",
		X"35",X"C9",X"3E",X"06",X"32",X"5E",X"9A",X"CD",X"48",X"35",X"C9",X"7A",X"FE",X"04",X"DA",X"DA",
		X"36",X"3E",X"03",X"32",X"5E",X"9A",X"CD",X"48",X"35",X"C9",X"3E",X"02",X"32",X"5E",X"9A",X"CD",
		X"48",X"35",X"C9",X"7A",X"FE",X"04",X"DA",X"F2",X"36",X"3E",X"0B",X"32",X"5E",X"9A",X"CD",X"48",
		X"35",X"C9",X"3E",X"0A",X"32",X"5E",X"9A",X"CD",X"48",X"35",X"C9",X"7A",X"FE",X"04",X"DA",X"0A",
		X"37",X"3E",X"0D",X"32",X"5E",X"9A",X"CD",X"48",X"35",X"C9",X"3E",X"0C",X"32",X"5E",X"9A",X"CD",
		X"48",X"35",X"C9",X"7A",X"FE",X"04",X"DA",X"22",X"37",X"3E",X"0F",X"32",X"5E",X"9A",X"CD",X"48",
		X"35",X"C9",X"3E",X"0E",X"32",X"5E",X"9A",X"CD",X"48",X"35",X"C9",X"CD",X"55",X"37",X"3A",X"6A",
		X"9C",X"47",X"3A",X"6B",X"9C",X"B0",X"C0",X"3E",X"FF",X"32",X"6C",X"9C",X"AF",X"CD",X"B5",X"10",
		X"C9",X"3A",X"76",X"9C",X"3C",X"32",X"76",X"9C",X"06",X"0F",X"0E",X"26",X"0D",X"C2",X"4C",X"37",
		X"05",X"C2",X"4A",X"37",X"C9",X"CD",X"41",X"37",X"3A",X"FB",X"9B",X"A7",X"CA",X"5D",X"39",X"AF",
		X"32",X"FB",X"9B",X"32",X"6A",X"9C",X"32",X"6B",X"9C",X"32",X"84",X"9C",X"32",X"80",X"9C",X"32",
		X"7E",X"9C",X"21",X"70",X"00",X"22",X"82",X"9C",X"DD",X"21",X"01",X"9C",X"21",X"78",X"9C",X"11",
		X"6A",X"9C",X"CD",X"9F",X"37",X"DD",X"21",X"07",X"9C",X"21",X"7A",X"9C",X"11",X"6B",X"9C",X"CD",
		X"9F",X"37",X"3A",X"6A",X"9C",X"47",X"3A",X"6B",X"9C",X"B0",X"C8",X"CD",X"A5",X"3A",X"C9",X"FD",
		X"21",X"64",X"3B",X"CD",X"16",X"39",X"A7",X"C8",X"FD",X"21",X"5A",X"9C",X"CD",X"16",X"39",X"A7",
		X"C8",X"3E",X"FF",X"12",X"FD",X"21",X"4A",X"9C",X"CD",X"16",X"39",X"A7",X"CA",X"2F",X"38",X"FD",
		X"21",X"3A",X"9C",X"CD",X"16",X"39",X"A7",X"CA",X"65",X"38",X"FD",X"21",X"2A",X"9C",X"CD",X"16",
		X"39",X"A7",X"CA",X"9C",X"38",X"FD",X"21",X"1A",X"9C",X"CD",X"16",X"39",X"A7",X"CA",X"D9",X"38",
		X"FD",X"22",X"7C",X"9C",X"ED",X"4B",X"7C",X"9C",X"71",X"23",X"70",X"21",X"5A",X"9C",X"11",X"0F",
		X"00",X"19",X"EB",X"21",X"5A",X"9C",X"2B",X"01",X"3F",X"00",X"ED",X"B8",X"21",X"1A",X"9C",X"23",
		X"54",X"5D",X"2B",X"3E",X"FF",X"77",X"01",X"0F",X"00",X"ED",X"B0",X"11",X"1A",X"9C",X"DD",X"22",
		X"7C",X"9C",X"2A",X"7C",X"9C",X"01",X"06",X"00",X"ED",X"B0",X"2A",X"7C",X"9C",X"11",X"01",X"9C",
		X"A7",X"ED",X"52",X"C8",X"2A",X"78",X"9C",X"11",X"10",X"00",X"19",X"22",X"78",X"9C",X"C9",X"01",
		X"5A",X"9C",X"71",X"23",X"70",X"21",X"5A",X"9C",X"23",X"54",X"5D",X"2B",X"3E",X"FF",X"77",X"01",
		X"0F",X"00",X"ED",X"B0",X"DD",X"22",X"7C",X"9C",X"2A",X"7C",X"9C",X"11",X"5A",X"9C",X"01",X"06",
		X"00",X"ED",X"B0",X"3A",X"84",X"9C",X"A7",X"C2",X"60",X"38",X"3E",X"FF",X"32",X"84",X"9C",X"C9",
		X"AF",X"32",X"6A",X"9C",X"C9",X"01",X"4A",X"9C",X"71",X"23",X"70",X"21",X"4A",X"9C",X"11",X"5A",
		X"9C",X"01",X"0F",X"00",X"ED",X"B0",X"21",X"4A",X"9C",X"23",X"54",X"5D",X"2B",X"3E",X"FF",X"77",
		X"01",X"0F",X"00",X"ED",X"B0",X"DD",X"22",X"7C",X"9C",X"2A",X"7C",X"9C",X"11",X"4A",X"9C",X"01",
		X"06",X"00",X"ED",X"B0",X"DD",X"21",X"4A",X"9C",X"CD",X"40",X"3B",X"C9",X"01",X"3A",X"9C",X"71",
		X"23",X"70",X"21",X"5A",X"9C",X"11",X"0F",X"00",X"19",X"EB",X"21",X"5A",X"9C",X"2B",X"01",X"1F",
		X"00",X"ED",X"B8",X"21",X"3A",X"9C",X"23",X"54",X"5D",X"2B",X"01",X"0F",X"00",X"3E",X"FF",X"77",
		X"ED",X"B0",X"DD",X"22",X"7C",X"9C",X"2A",X"7C",X"9C",X"11",X"3A",X"9C",X"01",X"06",X"00",X"ED",
		X"B0",X"DD",X"21",X"3A",X"9C",X"CD",X"40",X"3B",X"C9",X"01",X"2A",X"9C",X"71",X"23",X"70",X"21",
		X"5A",X"9C",X"11",X"0F",X"00",X"19",X"EB",X"21",X"5A",X"9C",X"2B",X"01",X"2F",X"00",X"ED",X"B8",
		X"21",X"2A",X"9C",X"23",X"54",X"5D",X"2B",X"3E",X"FF",X"77",X"01",X"0F",X"00",X"ED",X"B0",X"DD",
		X"22",X"7C",X"9C",X"2A",X"7C",X"9C",X"11",X"2A",X"9C",X"01",X"06",X"00",X"ED",X"B0",X"DD",X"21",
		X"2A",X"9C",X"CD",X"40",X"3B",X"C9",X"DD",X"7E",X"00",X"FD",X"46",X"00",X"B8",X"DA",X"57",X"39",
		X"C2",X"5A",X"39",X"DD",X"7E",X"01",X"FD",X"46",X"01",X"B8",X"DA",X"57",X"39",X"C2",X"5A",X"39",
		X"DD",X"7E",X"02",X"FD",X"46",X"02",X"B8",X"DA",X"57",X"39",X"C2",X"5A",X"39",X"DD",X"7E",X"03",
		X"FD",X"46",X"03",X"B8",X"DA",X"57",X"39",X"C2",X"5A",X"39",X"DD",X"7E",X"04",X"FD",X"46",X"04",
		X"B8",X"DA",X"57",X"39",X"C2",X"5A",X"39",X"3E",X"00",X"C9",X"3E",X"FF",X"C9",X"DD",X"21",X"78",
		X"9C",X"CD",X"8D",X"0B",X"FD",X"21",X"6A",X"9C",X"3A",X"6A",X"9C",X"A7",X"C2",X"87",X"39",X"DD",
		X"21",X"7A",X"9C",X"3E",X"FF",X"32",X"5D",X"9A",X"CD",X"8D",X"0B",X"FD",X"21",X"6B",X"9C",X"3A",
		X"6B",X"9C",X"A7",X"C2",X"87",X"39",X"C9",X"3A",X"76",X"9C",X"E6",X"3F",X"C0",X"2A",X"82",X"9C",
		X"2B",X"22",X"82",X"9C",X"7D",X"44",X"B0",X"CA",X"29",X"3A",X"3A",X"54",X"9A",X"57",X"FE",X"01",
		X"CC",X"03",X"3A",X"7A",X"FE",X"02",X"CC",X"16",X"3A",X"CD",X"64",X"3A",X"3A",X"56",X"9A",X"A7",
		X"CA",X"FE",X"39",X"3A",X"93",X"9C",X"A7",X"C0",X"3E",X"FF",X"32",X"93",X"9C",X"3A",X"7E",X"9C",
		X"FE",X"1C",X"CA",X"29",X"3A",X"3A",X"7E",X"9C",X"FE",X"1B",X"CA",X"3D",X"3A",X"3A",X"80",X"9C",
		X"FE",X"03",X"C8",X"D0",X"6F",X"26",X"00",X"DD",X"4E",X"00",X"DD",X"46",X"01",X"09",X"22",X"7C",
		X"9C",X"DD",X"2A",X"7C",X"9C",X"3A",X"7E",X"9C",X"4F",X"06",X"00",X"21",X"6A",X"3B",X"09",X"7E",
		X"DD",X"77",X"06",X"3A",X"80",X"9C",X"3C",X"32",X"80",X"9C",X"CD",X"A5",X"3A",X"C9",X"AF",X"32",
		X"93",X"9C",X"C9",X"3A",X"7E",X"9C",X"FE",X"1C",X"CA",X"10",X"3A",X"3C",X"32",X"7E",X"9C",X"C9",
		X"3E",X"00",X"32",X"7E",X"9C",X"C9",X"3A",X"7E",X"9C",X"FE",X"00",X"CA",X"23",X"3A",X"3D",X"32",
		X"7E",X"9C",X"C9",X"3E",X"1C",X"32",X"7E",X"9C",X"C9",X"AF",X"FD",X"77",X"00",X"32",X"7E",X"9C",
		X"32",X"80",X"9C",X"21",X"70",X"00",X"22",X"82",X"9C",X"CD",X"A5",X"3A",X"C9",X"3A",X"80",X"9C",
		X"FE",X"00",X"CA",X"FA",X"39",X"4F",X"06",X"00",X"3D",X"32",X"80",X"9C",X"DD",X"6E",X"00",X"DD",
		X"66",X"01",X"09",X"22",X"7C",X"9C",X"DD",X"2A",X"7C",X"9C",X"DD",X"2B",X"3E",X"FF",X"DD",X"77",
		X"06",X"C3",X"FA",X"39",X"21",X"6A",X"3B",X"06",X"00",X"3A",X"7E",X"9C",X"FE",X"1B",X"CA",X"85",
		X"3A",X"FE",X"1C",X"CA",X"95",X"3A",X"4F",X"09",X"7E",X"32",X"F8",X"85",X"3E",X"FF",X"32",X"18",
		X"86",X"32",X"D8",X"85",X"C9",X"3E",X"1B",X"32",X"D8",X"85",X"3E",X"1E",X"32",X"F8",X"85",X"3E",
		X"0B",X"32",X"18",X"86",X"C9",X"3E",X"0E",X"32",X"D8",X"85",X"3E",X"17",X"32",X"F8",X"85",X"3E",
		X"0D",X"32",X"18",X"86",X"C9",X"00",X"CD",X"B5",X"10",X"3E",X"01",X"32",X"D5",X"84",X"3E",X"02",
		X"32",X"D3",X"84",X"3E",X"03",X"32",X"D1",X"84",X"3E",X"04",X"32",X"CF",X"84",X"3E",X"05",X"32",
		X"CD",X"84",X"DD",X"21",X"1A",X"9C",X"21",X"15",X"85",X"CD",X"F5",X"3A",X"DD",X"21",X"2A",X"9C",
		X"21",X"13",X"85",X"CD",X"F5",X"3A",X"DD",X"21",X"3A",X"9C",X"21",X"11",X"85",X"CD",X"F5",X"3A",
		X"DD",X"21",X"4A",X"9C",X"21",X"0F",X"85",X"CD",X"F5",X"3A",X"DD",X"21",X"5A",X"9C",X"21",X"0D",
		X"85",X"CD",X"F5",X"3A",X"C9",X"E5",X"06",X"06",X"11",X"20",X"00",X"DD",X"7E",X"00",X"77",X"DD",
		X"23",X"19",X"05",X"C2",X"FB",X"3A",X"06",X"06",X"11",X"00",X"08",X"19",X"11",X"E0",X"FF",X"19",
		X"3E",X"00",X"77",X"19",X"05",X"C2",X"12",X"3B",X"E1",X"11",X"20",X"01",X"19",X"06",X"0A",X"11",
		X"20",X"00",X"DD",X"7E",X"00",X"77",X"DD",X"23",X"19",X"05",X"C2",X"22",X"3B",X"06",X"0A",X"11",
		X"00",X"08",X"19",X"11",X"E0",X"FF",X"19",X"3E",X"01",X"77",X"19",X"05",X"C2",X"39",X"3B",X"C9",
		X"2A",X"7C",X"9C",X"11",X"01",X"9C",X"A7",X"ED",X"52",X"C8",X"2A",X"78",X"9C",X"DD",X"22",X"7C",
		X"9C",X"ED",X"5B",X"7C",X"9C",X"A7",X"ED",X"52",X"D8",X"2A",X"78",X"9C",X"11",X"10",X"00",X"19",
		X"22",X"78",X"9C",X"C9",X"00",X"00",X"03",X"00",X"00",X"00",X"0A",X"0B",X"0C",X"0D",X"0E",X"0F",
		X"10",X"11",X"12",X"13",X"14",X"15",X"16",X"17",X"18",X"19",X"1A",X"1B",X"1C",X"1D",X"1E",X"1F",
		X"20",X"21",X"22",X"23",X"4D",X"4D",X"FF",X"FF",X"FF",X"FF",X"11",X"02",X"13",X"85",X"19",X"1E",
		X"1C",X"11",X"FF",X"1C",X"1D",X"0A",X"1B",X"1D",X"FF",X"0B",X"1E",X"1D",X"1D",X"18",X"17",X"0D",
		X"02",X"50",X"85",X"01",X"FF",X"19",X"15",X"0A",X"22",X"0E",X"1B",X"FF",X"18",X"17",X"15",X"22",
		X"0E",X"02",X"50",X"85",X"01",X"FF",X"18",X"1B",X"FF",X"02",X"FF",X"19",X"15",X"0A",X"22",X"0E",
		X"1B",X"1C",X"10",X"01",X"51",X"85",X"19",X"15",X"0E",X"0A",X"1C",X"0E",X"FF",X"16",X"18",X"1B",
		X"0E",X"FF",X"0C",X"18",X"12",X"17",X"13",X"01",X"4C",X"85",X"0C",X"18",X"12",X"17",X"FF",X"0A",
		X"FF",X"FF",X"01",X"0C",X"18",X"12",X"17",X"FF",X"01",X"19",X"15",X"0A",X"22",X"13",X"01",X"4C",
		X"85",X"0C",X"18",X"12",X"17",X"FF",X"0A",X"FF",X"02",X"0C",X"18",X"12",X"17",X"1C",X"FF",X"01",
		X"19",X"15",X"0A",X"22",X"13",X"01",X"4C",X"85",X"0C",X"18",X"12",X"17",X"FF",X"0A",X"FF",X"03",
		X"0C",X"18",X"12",X"17",X"1C",X"FF",X"01",X"19",X"15",X"0A",X"22",X"13",X"01",X"4C",X"85",X"0C",
		X"18",X"12",X"17",X"FF",X"0A",X"FF",X"04",X"0C",X"18",X"12",X"17",X"1C",X"FF",X"01",X"19",X"15",
		X"0A",X"22",X"13",X"01",X"4C",X"85",X"0C",X"18",X"12",X"17",X"FF",X"0A",X"FF",X"FF",X"01",X"0C",
		X"18",X"12",X"17",X"FF",X"02",X"19",X"15",X"0A",X"22",X"13",X"01",X"4C",X"85",X"0C",X"18",X"12",
		X"17",X"FF",X"0A",X"FF",X"FF",X"01",X"0C",X"18",X"12",X"17",X"FF",X"03",X"19",X"15",X"0A",X"22",
		X"13",X"01",X"4C",X"85",X"0C",X"18",X"12",X"17",X"FF",X"0A",X"FF",X"02",X"0C",X"18",X"12",X"17",
		X"1C",X"FF",X"03",X"19",X"15",X"0A",X"22",X"D6",X"3B",X"ED",X"3B",X"04",X"3C",X"1B",X"3C",X"32",
		X"3C",X"49",X"3C",X"60",X"3C",X"13",X"01",X"4D",X"85",X"0C",X"18",X"12",X"17",X"FF",X"0B",X"FF",
		X"FF",X"01",X"0C",X"18",X"12",X"17",X"FF",X"01",X"19",X"15",X"0A",X"22",X"13",X"01",X"4D",X"85",
		X"0C",X"18",X"12",X"17",X"FF",X"0B",X"FF",X"02",X"0C",X"18",X"12",X"17",X"1C",X"FF",X"01",X"19",
		X"15",X"0A",X"22",X"13",X"01",X"4D",X"85",X"0C",X"18",X"12",X"17",X"FF",X"0B",X"FF",X"03",X"0C",
		X"18",X"12",X"17",X"1C",X"FF",X"01",X"19",X"15",X"0A",X"22",X"13",X"01",X"4D",X"85",X"0C",X"18",
		X"12",X"17",X"FF",X"0B",X"FF",X"04",X"0C",X"18",X"12",X"17",X"1C",X"FF",X"01",X"19",X"15",X"0A",
		X"22",X"13",X"01",X"4D",X"85",X"0C",X"18",X"12",X"17",X"FF",X"0B",X"FF",X"FF",X"01",X"0C",X"18",
		X"12",X"17",X"FF",X"02",X"19",X"15",X"0A",X"22",X"13",X"01",X"4D",X"85",X"0C",X"18",X"12",X"17",
		X"FF",X"0B",X"FF",X"FF",X"01",X"0C",X"18",X"12",X"17",X"FF",X"03",X"19",X"15",X"0A",X"22",X"13",
		X"01",X"4D",X"85",X"0C",X"18",X"12",X"17",X"FF",X"0B",X"FF",X"02",X"0C",X"18",X"12",X"17",X"1C",
		X"FF",X"03",X"19",X"15",X"0A",X"22",X"85",X"3C",X"9C",X"3C",X"B3",X"3C",X"CA",X"3C",X"E1",X"3C",
		X"F8",X"3C",X"0F",X"3D",X"09",X"01",X"50",X"85",X"10",X"0A",X"16",X"0E",X"FF",X"18",X"1F",X"0E",
		X"1B",X"0A",X"0A",X"0A",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0C",X"1B",X"0E",X"0D",X"12",
		X"1D",X"FF",X"00",X"0B",X"01",X"B5",X"85",X"12",X"17",X"1C",X"0E",X"1B",X"1D",X"FF",X"0C",X"18",
		X"12",X"17",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"34",X"85",X"FF",X"01",
		X"1E",X"19",X"FF",X"10",X"0A",X"16",X"0E",X"FF",X"18",X"1F",X"0E",X"1B",X"FF",X"FF",X"10",X"00",
		X"34",X"85",X"FF",X"02",X"1E",X"19",X"FF",X"10",X"0A",X"16",X"0E",X"FF",X"18",X"1F",X"0E",X"1B",
		X"FF",X"FF",X"09",X"00",X"74",X"85",X"10",X"0A",X"16",X"0E",X"FF",X"18",X"1F",X"0E",X"1B",X"05",
		X"00",X"B4",X"85",X"1C",X"1D",X"0A",X"1B",X"1D",X"10",X"00",X"4E",X"85",X"24",X"FF",X"01",X"09",
		X"08",X"03",X"FF",X"0F",X"0A",X"15",X"0C",X"18",X"17",X"FF",X"FF",X"FF",X"00",X"00",X"07",X"05",
		X"00",X"00",X"0F",X"0A",X"15",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"06",X"08",
		X"00",X"00",X"0E",X"15",X"1C",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"05",X"05",
		X"00",X"00",X"14",X"FF",X"22",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"03",X"09",
		X"00",X"00",X"1D",X"14",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"03",X"08",
		X"00",X"00",X"1D",X"1C",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0E",X"00",X"C9",X"96",
		X"0D",X"18",X"FF",X"17",X"18",X"1D",X"FF",X"1B",X"0E",X"20",X"1B",X"12",X"1D",X"0E",X"FF",X"FF",
		X"0B",X"00",X"6B",X"96",X"16",X"0E",X"16",X"18",X"1B",X"22",X"FF",X"0D",X"0A",X"1D",X"0A",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"03",X"00",X"30",X"96",X"0E",X"15",X"1C",X"0F",X"00",X"07",X"0F",X"01",
		X"08",X"0F",X"02",X"09",X"0F",X"03",X"0A",X"0F",X"04",X"0B",X"0F",X"05",X"0C",X"0F",X"06",X"0D",
		X"0F",X"07",X"0E",X"0F",X"08",X"0F",X"0F",X"09",X"01",X"0F",X"0A",X"02",X"0F",X"1A",X"00",X"0F",
		X"1B",X"00",X"0F",X"1E",X"00",X"03",X"1D",X"00",X"0F",X"0B",X"00",X"0F",X"0C",X"00",X"0F",X"0D",
		X"00",X"0F",X"0E",X"00",X"0F",X"0F",X"00",X"0F",X"10",X"03",X"0F",X"11",X"04",X"0F",X"12",X"05",
		X"0F",X"13",X"06",X"0F",X"14",X"07",X"0F",X"15",X"03",X"0F",X"16",X"04",X"0F",X"17",X"05",X"0F",
		X"18",X"06",X"0F",X"19",X"07",X"3D",X"3D",X"3D",X"3D",X"3D",X"3D",X"3D",X"3D",X"42",X"7A",X"7A",
		X"7A",X"7A",X"7A",X"7A",X"3A",X"43",X"7A",X"3A",X"37",X"41",X"3C",X"43",X"39",X"41",X"39",X"40",
		X"3F",X"3F",X"3E",X"3D",X"3D",X"38",X"3C",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"3B",X"37",X"7A",
		X"7A",X"7A",X"7A",X"3C",X"7A",X"7A",X"7A",X"3B",X"3A",X"37",X"39",X"4F",X"84",X"6F",X"84",X"8F",
		X"84",X"AF",X"84",X"CF",X"84",X"EF",X"84",X"0F",X"85",X"2F",X"85",X"4F",X"85",X"50",X"84",X"70",
		X"84",X"90",X"84",X"B0",X"84",X"D0",X"84",X"F0",X"84",X"10",X"85",X"30",X"85",X"51",X"84",X"71",
		X"84",X"91",X"84",X"B1",X"84",X"D1",X"84",X"F1",X"84",X"11",X"85",X"52",X"84",X"72",X"84",X"EF",
		X"86",X"0F",X"87",X"2F",X"87",X"4F",X"87",X"6F",X"87",X"8F",X"87",X"AF",X"87",X"F0",X"86",X"10",
		X"87",X"30",X"87",X"50",X"87",X"70",X"87",X"90",X"87",X"B0",X"87",X"11",X"87",X"31",X"87",X"51",
		X"87",X"71",X"87",X"91",X"87",X"B1",X"87",X"52",X"87",X"72",X"87",X"92",X"87",X"B2",X"87",X"73",
		X"87",X"93",X"87",X"B3",X"87",X"94",X"87",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",
		X"40",X"20",X"40",X"20",X"30",X"40",X"20",X"30",X"40",X"20",X"40",X"20",X"30",X"20",X"30",X"FE",
		X"00",X"93",X"10",X"FE",X"00",X"93",X"10",X"FE",X"10",X"93",X"10",X"FE",X"00",X"93",X"10",X"FE",
		X"00",X"93",X"10",X"FE",X"00",X"93",X"10",X"FE",X"00",X"93",X"10",X"FE",X"00",X"93",X"10",X"FE",
		X"00",X"93",X"10",X"FE",X"00",X"93",X"10",X"FE",X"00",X"93",X"10",X"FE",X"00",X"93",X"10",X"FE",
		X"00",X"93",X"10",X"FE",X"00",X"93",X"10",X"FE",X"00",X"93",X"10",X"FE",X"00",X"93",X"10",X"FE",
		X"00",X"93",X"10",X"FE",X"00",X"93",X"10",X"FE",X"00",X"93",X"10",X"FE",X"00",X"93",X"10",X"FE",
		X"00",X"93",X"10",X"FE",X"00",X"93",X"10",X"FE",X"00",X"93",X"10",X"FE",X"00",X"93",X"10",X"FE",
		X"00",X"93",X"10",X"FE",X"00",X"93",X"10",X"FE",X"00",X"93",X"10",X"FE",X"00",X"93",X"10",X"FE",
		X"00",X"93",X"10",X"FE",X"00",X"93",X"10",X"FE",X"00",X"93",X"10",X"FE",X"00",X"93",X"10",X"FE",
		X"00",X"93",X"10",X"FE",X"00",X"93",X"10",X"FE",X"00",X"93",X"10",X"FE",X"00",X"93",X"10",X"FE",
		X"00",X"93",X"10",X"FE",X"00",X"93",X"10",X"FE",X"00",X"93",X"10",X"FE",X"00",X"93",X"10",X"FE",
		X"00",X"93",X"10",X"80",X"62",X"02",X"00",X"8B",X"10",X"02",X"00",X"8B",X"10",X"02",X"00",X"8B",
		X"10",X"02",X"00",X"8B",X"10",X"02",X"00",X"8B",X"10",X"02",X"00",X"8B",X"10",X"02",X"00",X"8B",
		X"10",X"02",X"00",X"8B",X"10",X"02",X"00",X"8B",X"10",X"02",X"00",X"8B",X"10",X"02",X"00",X"8B",
		X"10",X"02",X"00",X"8B",X"10",X"02",X"00",X"8B",X"10",X"02",X"00",X"8B",X"10",X"02",X"00",X"8B",
		X"10",X"02",X"00",X"8B",X"10",X"02",X"00",X"8B",X"10",X"02",X"00",X"8B",X"10",X"02",X"00",X"8B",
		X"10",X"02",X"00",X"8B",X"10",X"02",X"00",X"8B",X"10",X"02",X"00",X"8B",X"10",X"02",X"00",X"8B",
		X"10",X"02",X"00",X"8B",X"10",X"02",X"00",X"8B",X"10",X"02",X"00",X"8B",X"10",X"02",X"00",X"8B",
		X"10",X"02",X"00",X"8B",X"10",X"02",X"00",X"8B",X"10",X"02",X"00",X"8B",X"10",X"02",X"00",X"8B",
		X"10",X"02",X"00",X"8B",X"10",X"02",X"00",X"8B",X"10",X"02",X"00",X"8B",X"10",X"02",X"00",X"8B",
		X"10",X"02",X"00",X"8B",X"10",X"02",X"00",X"8B",X"10",X"02",X"00",X"8B",X"10",X"02",X"00",X"8B",
		X"10",X"80",X"73",X"98",X"4B",X"78",X"4A",X"DC",X"4A",X"AA",X"4A",X"CA",X"4B",X"3A",X"4B",X"05",
		X"40",X"5F",X"3F",X"10",X"58",X"12",X"58",X"14",X"58",X"16",X"58",X"18",X"58",X"1A",X"58",X"1C",
		X"58",X"1E",X"58",X"20",X"58",X"22",X"58",X"24",X"58",X"26",X"58",X"28",X"58",X"2A",X"58",X"2C",
		X"58",X"2E",X"58",X"30",X"58",X"32",X"58",X"34",X"58",X"36",X"58",X"38",X"58",X"3A",X"58",X"3C",
		X"58",X"3E",X"58",X"40",X"58",X"42",X"58",X"44",X"58",X"46",X"58",X"48",X"58",X"4A",X"58",X"4C",
		X"58",X"4E",X"58",X"50",X"58",X"52",X"58",X"54",X"58",X"56",X"58",X"58",X"58",X"5A",X"58",X"5C",
		X"58",X"5E",X"58",X"60",X"58",X"62",X"58",X"64",X"58",X"66",X"58",X"68",X"58",X"6A",X"58",X"6C",
		X"58",X"6E",X"58",X"70",X"58",X"72",X"58",X"74",X"58",X"76",X"58",X"78",X"58",X"7A",X"58",X"7C",
		X"58",X"7E",X"58",X"80",X"58",X"82",X"58",X"84",X"58",X"86",X"58",X"88",X"58",X"8A",X"58",X"8C",
		X"58",X"8E",X"58",X"90",X"58",X"92",X"58",X"94",X"58",X"96",X"58",X"98",X"58",X"9A",X"58",X"9C",
		X"58",X"9E",X"58",X"A0",X"58",X"A2",X"58",X"A4",X"58",X"A6",X"58",X"A8",X"58",X"AA",X"58",X"AC",
		X"58",X"AE",X"58",X"B0",X"58",X"B2",X"58",X"B4",X"58",X"B6",X"58",X"B8",X"58",X"BA",X"58",X"BC",
		X"58",X"BE",X"58",X"C0",X"58",X"C2",X"58",X"C4",X"58",X"C6",X"58",X"C8",X"58",X"CA",X"58",X"CC",
		X"58",X"CE",X"58",X"D0",X"58",X"D2",X"58",X"D4",X"58",X"D6",X"58",X"D8",X"58",X"DA",X"58",X"DC",
		X"58",X"DE",X"58",X"E0",X"58",X"E2",X"58",X"E4",X"58",X"E6",X"58",X"E8",X"58",X"EA",X"58",X"EC",
		X"58",X"EE",X"58",X"F0",X"58",X"FF",X"FF",X"F5",X"84",X"F4",X"84",X"F3",X"84",X"F5",X"84",X"F4",
		X"84",X"F3",X"84",X"15",X"85",X"14",X"85",X"13",X"85",X"35",X"85",X"34",X"85",X"33",X"85",X"1F",
		X"20",X"21",X"1F",X"20",X"21",X"1C",X"1D",X"1E",X"19",X"1A",X"1B",X"4B",X"4B",X"4B",X"4B",X"4B",
		X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"55",X"85",X"54",X"85",X"53",X"85",X"55",X"85",X"54",
		X"85",X"53",X"85",X"55",X"85",X"54",X"85",X"53",X"85",X"75",X"85",X"74",X"85",X"73",X"85",X"16",
		X"17",X"18",X"16",X"17",X"18",X"16",X"17",X"18",X"13",X"14",X"15",X"4B",X"4B",X"4B",X"4B",X"4B",
		X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"95",X"85",X"94",X"85",X"93",X"85",X"95",X"85",X"94",
		X"85",X"93",X"85",X"B5",X"85",X"B4",X"85",X"B3",X"85",X"D5",X"85",X"D4",X"85",X"D3",X"85",X"10",
		X"11",X"12",X"10",X"11",X"12",X"0D",X"0E",X"0F",X"0A",X"0B",X"0C",X"4B",X"4B",X"4B",X"4B",X"4B",
		X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"F5",X"85",X"F4",X"85",X"F3",X"85",X"F5",X"85",X"F4",
		X"85",X"F3",X"85",X"F5",X"85",X"F4",X"85",X"F3",X"85",X"15",X"86",X"14",X"86",X"13",X"86",X"07",
		X"08",X"09",X"07",X"08",X"09",X"07",X"08",X"09",X"04",X"05",X"06",X"4B",X"4B",X"4B",X"4B",X"4B",
		X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"75",X"86",X"74",X"86",X"73",X"86",X"75",X"86",X"74",
		X"86",X"73",X"86",X"95",X"86",X"94",X"86",X"93",X"86",X"B5",X"86",X"B4",X"86",X"B3",X"86",X"FA",
		X"FB",X"FC",X"FA",X"FB",X"FC",X"F7",X"F8",X"F9",X"F4",X"F5",X"F6",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"D5",X"86",X"D4",X"86",X"D3",X"86",X"F5",X"86",X"F4",
		X"86",X"F3",X"86",X"15",X"87",X"14",X"87",X"13",X"87",X"35",X"87",X"34",X"87",X"33",X"87",X"F1",
		X"F2",X"F3",X"EE",X"EF",X"F0",X"EB",X"EC",X"ED",X"E8",X"E9",X"EA",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"35",X"86",X"34",X"86",X"33",X"86",X"35",X"86",X"34",
		X"86",X"33",X"86",X"35",X"86",X"34",X"86",X"33",X"86",X"55",X"86",X"54",X"86",X"53",X"86",X"01",
		X"02",X"03",X"01",X"02",X"03",X"01",X"02",X"03",X"FD",X"FE",X"00",X"4B",X"4B",X"4B",X"4B",X"4B",
		X"4B",X"4B",X"4B",X"4B",X"0B",X"0B",X"4B",X"08",X"00",X"00",X"0A",X"00",X"01",X"0C",X"00",X"02",
		X"0E",X"00",X"03",X"10",X"00",X"04",X"12",X"00",X"05",X"14",X"00",X"06",X"97",X"41",X"C7",X"41",
		X"F7",X"41",X"27",X"42",X"B7",X"42",X"57",X"42",X"87",X"42",X"24",X"FF",X"01",X"09",X"08",X"03",
		X"FF",X"2A",X"29",X"28",X"27",X"26",X"25",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"10",X"30",X"12",X"30",X"14",X"30",X"16",X"30",X"18",X"30",X"1A",X"30",
		X"1C",X"30",X"1E",X"30",X"20",X"30",X"22",X"30",X"24",X"30",X"26",X"30",X"28",X"30",X"2A",X"30",
		X"2C",X"30",X"2E",X"30",X"30",X"30",X"32",X"30",X"34",X"30",X"36",X"30",X"38",X"30",X"3A",X"30",
		X"3C",X"30",X"3E",X"30",X"40",X"30",X"42",X"30",X"44",X"30",X"46",X"30",X"48",X"30",X"4A",X"30",
		X"4C",X"30",X"4E",X"30",X"50",X"30",X"52",X"30",X"54",X"30",X"56",X"30",X"58",X"30",X"5A",X"30",
		X"5C",X"30",X"5E",X"30",X"60",X"30",X"62",X"30",X"64",X"30",X"66",X"30",X"68",X"30",X"6A",X"30",
		X"6C",X"30",X"6E",X"30",X"70",X"30",X"72",X"30",X"74",X"30",X"76",X"30",X"78",X"30",X"7A",X"30",
		X"7C",X"30",X"7E",X"30",X"80",X"30",X"82",X"30",X"84",X"30",X"86",X"30",X"88",X"30",X"8A",X"30",
		X"8C",X"30",X"8E",X"30",X"90",X"30",X"92",X"30",X"94",X"30",X"96",X"30",X"98",X"30",X"9A",X"30",
		X"9C",X"30",X"9E",X"30",X"A0",X"30",X"A2",X"30",X"A4",X"30",X"A6",X"30",X"A8",X"30",X"AA",X"30",
		X"AC",X"30",X"AE",X"30",X"B0",X"30",X"B2",X"30",X"B4",X"30",X"B6",X"30",X"B8",X"30",X"BA",X"30",
		X"BC",X"30",X"BE",X"30",X"C0",X"30",X"C2",X"30",X"C4",X"30",X"C6",X"30",X"C8",X"30",X"CA",X"30",
		X"CC",X"30",X"CE",X"30",X"D0",X"30",X"D2",X"30",X"D4",X"30",X"D6",X"30",X"D8",X"30",X"DA",X"30",
		X"DC",X"30",X"DE",X"30",X"E0",X"30",X"E2",X"30",X"E4",X"30",X"E6",X"30",X"E8",X"30",X"EA",X"30",
		X"EC",X"30",X"EE",X"30",X"F0",X"30",X"F8",X"30",X"FF",X"FF",X"FF",X"FF",X"01",X"01",X"34",X"31",
		X"2E",X"2B",X"7F",X"35",X"32",X"2F",X"2C",X"7F",X"34",X"31",X"2E",X"2B",X"7F",X"35",X"32",X"2F",
		X"2C",X"7F",X"34",X"31",X"2E",X"2B",X"7F",X"35",X"32",X"2F",X"2C",X"7F",X"34",X"31",X"2E",X"2B",
		X"7F",X"35",X"32",X"2F",X"2C",X"7F",X"01",X"01",X"36",X"33",X"30",X"2D",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"36",X"33",X"30",X"2D",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"36",X"33",X"30",X"2D",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"36",X"33",X"30",X"2D",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"A0",X"E0",X"A0",X"D8",X"A0",X"D0",X"A0",X"C8",X"A0",X"C0",X"A0",X"B8",X"A0",X"B0",X"A0",X"A8",
		X"A0",X"A0",X"A0",X"98",X"A0",X"90",X"A0",X"88",X"A0",X"80",X"A0",X"80",X"A0",X"80",X"A0",X"80",
		X"A0",X"80",X"A0",X"80",X"A0",X"80",X"A0",X"80",X"A0",X"80",X"A0",X"80",X"A0",X"80",X"A0",X"80",
		X"A0",X"80",X"A0",X"80",X"A0",X"80",X"A0",X"80",X"A0",X"80",X"A0",X"80",X"A0",X"80",X"A0",X"80",
		X"A0",X"80",X"A0",X"80",X"A0",X"80",X"A0",X"80",X"A0",X"80",X"A0",X"80",X"A0",X"80",X"A0",X"80",
		X"05",X"00",X"91",X"85",X"0B",X"18",X"17",X"1E",X"1C",X"06",X"00",X"6B",X"85",X"05",X"00",X"00",
		X"FF",X"4C",X"FF",X"00",X"00",X"00",X"05",X"00",X"10",X"00",X"15",X"00",X"20",X"00",X"25",X"00",
		X"30",X"00",X"35",X"00",X"40",X"00",X"45",X"00",X"50",X"10",X"10",X"20",X"01",X"02",X"02",X"02",
		X"00",X"10",X"01",X"01",X"01",X"02",X"02",X"10",X"20",X"00",X"00",X"20",X"20",X"10",X"10",X"10",
		X"01",X"01",X"01",X"02",X"02",X"02",X"10",X"10",X"10",X"20",X"20",X"01",X"01",X"20",X"10",X"20",
		X"20",X"10",X"01",X"01",X"02",X"02",X"02",X"10",X"10",X"10",X"10",X"10",X"01",X"01",X"02",X"02",
		X"00",X"23",X"45",X"2B",X"45",X"33",X"45",X"3B",X"45",X"43",X"45",X"4B",X"45",X"53",X"45",X"5B",
		X"45",X"63",X"45",X"04",X"01",X"51",X"86",X"00",X"00",X"00",X"00",X"04",X"01",X"51",X"86",X"FF",
		X"05",X"00",X"00",X"04",X"01",X"51",X"86",X"01",X"00",X"00",X"00",X"04",X"01",X"51",X"86",X"01",
		X"05",X"00",X"00",X"04",X"01",X"51",X"86",X"02",X"00",X"00",X"00",X"04",X"01",X"51",X"86",X"02",
		X"05",X"00",X"00",X"04",X"01",X"51",X"86",X"03",X"00",X"00",X"00",X"04",X"01",X"51",X"86",X"03",
		X"05",X"00",X"00",X"04",X"01",X"51",X"86",X"04",X"00",X"00",X"00",X"13",X"02",X"0F",X"85",X"4D",
		X"4D",X"4D",X"FF",X"05",X"00",X"FF",X"18",X"1B",X"FF",X"02",X"00",X"00",X"FF",X"19",X"18",X"12",
		X"17",X"1D",X"0D",X"02",X"0C",X"85",X"4D",X"4D",X"4D",X"FF",X"02",X"00",X"00",X"FF",X"19",X"18",
		X"12",X"17",X"1D",X"0D",X"02",X"09",X"85",X"4D",X"4D",X"4D",X"FF",X"03",X"00",X"00",X"FF",X"19",
		X"18",X"12",X"17",X"1D",X"0D",X"02",X"06",X"85",X"4D",X"4D",X"4D",X"FF",X"05",X"00",X"00",X"FF",
		X"19",X"18",X"12",X"17",X"1D",X"30",X"32",X"34",X"36",X"38",X"3A",X"3C",X"3E",X"40",X"42",X"44",
		X"46",X"48",X"4A",X"4C",X"4E",X"50",X"52",X"54",X"56",X"58",X"5A",X"5C",X"5E",X"0C",X"03",X"54",
		X"85",X"0D",X"18",X"17",X"1D",X"FF",X"1B",X"0E",X"20",X"1B",X"12",X"1D",X"0E",X"03",X"03",X"0D",
		X"86",X"0E",X"15",X"1C",X"07",X"08",X"09",X"09",X"0A",X"08",X"0A",X"0B",X"09",X"0A",X"11",X"13",
		X"06",X"07",X"07",X"07",X"06",X"04",X"08",X"08",X"03",X"05",X"04",X"04",X"FE",X"01",X"FE",X"00",
		X"FE",X"01",X"FE",X"00",X"FE",X"01",X"FE",X"01",X"FE",X"01",X"FF",X"02",X"00",X"02",X"01",X"02",
		X"02",X"01",X"02",X"01",X"02",X"01",X"02",X"00",X"02",X"01",X"02",X"00",X"02",X"01",X"02",X"01",
		X"01",X"00",X"00",X"00",X"80",X"9C",X"10",X"F0",X"B4",X"4E",X"62",X"B4",X"9E",X"B2",X"CC",X"20",
		X"32",X"CC",X"76",X"8B",X"CC",X"CE",X"E0",X"01",X"FD",X"03",X"FF",X"02",X"03",X"01",X"FD",X"03",
		X"FF",X"02",X"03",X"01",X"FD",X"03",X"FF",X"02",X"03",X"01",X"FD",X"03",X"FF",X"01",X"03",X"03",
		X"01",X"02",X"FD",X"01",X"03",X"03",X"01",X"02",X"FD",X"01",X"03",X"03",X"01",X"02",X"FD",X"01",
		X"03",X"03",X"01",X"02",X"FF",X"A7",X"13",X"02",X"00",X"A7",X"13",X"02",X"01",X"A7",X"13",X"02",
		X"01",X"A7",X"13",X"02",X"00",X"A7",X"13",X"02",X"FF",X"A7",X"13",X"80",X"02",X"FE",X"A7",X"13",
		X"02",X"00",X"A7",X"13",X"80",X"02",X"02",X"A7",X"13",X"02",X"00",X"A7",X"13",X"80",X"02",X"00",
		X"AF",X"13",X"02",X"00",X"AF",X"13",X"02",X"00",X"B3",X"13",X"02",X"00",X"B3",X"13",X"02",X"00",
		X"AF",X"13",X"02",X"00",X"AF",X"13",X"02",X"00",X"AB",X"13",X"02",X"00",X"AB",X"13",X"80",X"02",
		X"FE",X"B3",X"13",X"02",X"FE",X"B3",X"13",X"02",X"FF",X"B3",X"13",X"02",X"FF",X"AF",X"13",X"02",
		X"FF",X"B3",X"13",X"02",X"FE",X"B3",X"13",X"02",X"FE",X"B3",X"13",X"80",X"02",X"02",X"AB",X"13",
		X"02",X"02",X"AB",X"13",X"02",X"01",X"AB",X"13",X"02",X"01",X"AF",X"13",X"02",X"01",X"AB",X"13",
		X"02",X"02",X"AB",X"13",X"02",X"02",X"AB",X"13",X"80",X"18",X"30",X"50",X"60",X"80",X"A0",X"B0",
		X"D0",X"E9",X"FF",X"FD",X"00",X"FD",X"FF",X"FE",X"FE",X"FE",X"FD",X"FD",X"FE",X"FE",X"FD",X"FF",
		X"FD",X"00",X"FD",X"01",X"FD",X"01",X"FD",X"02",X"FD",X"02",X"FD",X"03",X"FE",X"02",X"FE",X"03",
		X"FE",X"03",X"FF",X"03",X"FF",X"03",X"FF",X"03",X"00",X"80",X"FE",X"00",X"FE",X"FF",X"FD",X"FF",
		X"FD",X"FF",X"FD",X"FE",X"FD",X"FE",X"00",X"FE",X"03",X"FE",X"03",X"FE",X"03",X"FF",X"03",X"FF",
		X"80",X"FD",X"00",X"FD",X"01",X"FE",X"02",X"FE",X"03",X"FD",X"02",X"FE",X"03",X"FF",X"03",X"00",
		X"03",X"01",X"03",X"01",X"03",X"02",X"03",X"02",X"03",X"03",X"02",X"02",X"02",X"03",X"02",X"03",
		X"01",X"03",X"01",X"03",X"01",X"03",X"00",X"80",X"FE",X"00",X"FE",X"01",X"FD",X"01",X"FD",X"01",
		X"FD",X"02",X"FD",X"02",X"00",X"02",X"03",X"02",X"03",X"02",X"03",X"01",X"03",X"01",X"80",X"A2",
		X"F0",X"E8",X"A2",X"B2",X"9E",X"A2",X"62",X"4E",X"BA",X"34",X"2C",X"BA",X"84",X"7C",X"BA",X"D2",
		X"CE",X"D2",X"A8",X"A4",X"D2",X"48",X"44",X"A2",X"E7",X"B9",X"A2",X"97",X"69",X"A2",X"47",X"19",
		X"BA",X"60",X"41",X"BA",X"B0",X"91",X"BA",X"E0",X"D0",X"D2",X"97",X"78",X"D2",X"3F",X"20",X"A4",
		X"A4",X"A4",X"BC",X"BC",X"D4",X"D4",X"D4",X"9C",X"C0",X"37",X"12",X"9C",X"70",X"37",X"12",X"9C",
		X"42",X"2F",X"12",X"B4",X"6A",X"2F",X"12",X"B4",X"98",X"37",X"12",X"CC",X"C8",X"37",X"12",X"CC",
		X"92",X"2F",X"12",X"CC",X"3A",X"2F",X"12",X"00",X"FE",X"4B",X"12",X"00",X"FE",X"4B",X"12",X"00",
		X"FE",X"4F",X"12",X"00",X"FE",X"4F",X"12",X"00",X"FE",X"53",X"12",X"00",X"FE",X"53",X"12",X"00",
		X"FE",X"4F",X"12",X"00",X"FE",X"4F",X"12",X"80",X"00",X"02",X"3F",X"12",X"00",X"02",X"3F",X"12",
		X"00",X"02",X"43",X"12",X"00",X"02",X"43",X"12",X"00",X"02",X"47",X"12",X"00",X"02",X"47",X"12",
		X"00",X"02",X"43",X"12",X"00",X"02",X"43",X"12",X"80",X"03",X"00",X"83",X"12",X"03",X"00",X"83",
		X"12",X"03",X"00",X"83",X"12",X"03",X"00",X"83",X"12",X"03",X"00",X"3F",X"12",X"02",X"02",X"3F",
		X"12",X"02",X"02",X"43",X"12",X"02",X"02",X"43",X"12",X"02",X"02",X"47",X"12",X"01",X"02",X"47",
		X"12",X"00",X"02",X"43",X"12",X"00",X"02",X"43",X"12",X"00",X"02",X"3F",X"12",X"00",X"02",X"3F",
		X"12",X"00",X"02",X"43",X"12",X"00",X"02",X"43",X"12",X"00",X"02",X"47",X"12",X"00",X"02",X"47",
		X"12",X"00",X"02",X"43",X"12",X"00",X"02",X"43",X"12",X"00",X"02",X"3F",X"12",X"00",X"02",X"3F",
		X"12",X"00",X"02",X"43",X"12",X"00",X"02",X"43",X"12",X"00",X"02",X"47",X"12",X"00",X"02",X"47",
		X"12",X"00",X"02",X"43",X"12",X"00",X"02",X"43",X"12",X"00",X"02",X"3F",X"12",X"00",X"02",X"3F",
		X"12",X"00",X"02",X"43",X"12",X"00",X"02",X"43",X"12",X"00",X"02",X"47",X"12",X"00",X"02",X"47",
		X"12",X"00",X"00",X"87",X"12",X"00",X"00",X"87",X"12",X"80",X"FD",X"01",X"57",X"12",X"FD",X"01",
		X"57",X"12",X"FD",X"01",X"57",X"12",X"FD",X"01",X"57",X"12",X"FE",X"02",X"57",X"12",X"FD",X"02",
		X"57",X"12",X"FE",X"03",X"57",X"12",X"FF",X"03",X"57",X"12",X"00",X"03",X"57",X"12",X"01",X"03",
		X"57",X"12",X"02",X"03",X"57",X"12",X"01",X"01",X"83",X"12",X"00",X"00",X"87",X"12",X"00",X"00",
		X"87",X"12",X"00",X"00",X"83",X"12",X"00",X"00",X"83",X"12",X"00",X"00",X"87",X"12",X"00",X"00",
		X"87",X"12",X"80",X"FD",X"FF",X"5B",X"12",X"FD",X"FF",X"5B",X"12",X"FD",X"FF",X"5B",X"12",X"FD",
		X"FF",X"5B",X"12",X"FE",X"FE",X"5B",X"12",X"FD",X"FE",X"5B",X"12",X"FE",X"FD",X"5B",X"12",X"FF",
		X"FD",X"5B",X"12",X"00",X"FD",X"5B",X"12",X"01",X"FD",X"5B",X"12",X"02",X"FD",X"5B",X"12",X"01",
		X"FF",X"83",X"12",X"00",X"00",X"87",X"12",X"00",X"00",X"87",X"12",X"00",X"00",X"83",X"12",X"00",
		X"00",X"83",X"12",X"00",X"00",X"87",X"12",X"00",X"00",X"87",X"12",X"80",X"00",X"02",X"57",X"12",
		X"01",X"03",X"57",X"12",X"03",X"02",X"57",X"12",X"03",X"01",X"57",X"12",X"01",X"00",X"83",X"12",
		X"00",X"00",X"87",X"12",X"00",X"00",X"87",X"12",X"00",X"00",X"87",X"12",X"00",X"00",X"83",X"12",
		X"00",X"00",X"83",X"12",X"00",X"00",X"87",X"12",X"00",X"00",X"87",X"12",X"80",X"00",X"02",X"57",
		X"12",X"01",X"03",X"57",X"12",X"03",X"02",X"57",X"12",X"03",X"02",X"57",X"12",X"00",X"00",X"87",
		X"12",X"80",X"00",X"00",X"6F",X"12",X"00",X"00",X"6F",X"12",X"00",X"06",X"73",X"12",X"00",X"00",
		X"73",X"12",X"00",X"00",X"73",X"12",X"80",X"00",X"00",X"7B",X"12",X"00",X"00",X"7B",X"12",X"00",
		X"FA",X"7F",X"12",X"00",X"00",X"7F",X"12",X"00",X"00",X"7F",X"12",X"80",X"00",X"00",X"77",X"12",
		X"00",X"00",X"7B",X"12",X"00",X"FA",X"7F",X"12",X"00",X"00",X"7F",X"12",X"80",X"00",X"00",X"6B",
		X"12",X"00",X"00",X"6F",X"12",X"00",X"06",X"73",X"12",X"00",X"00",X"73",X"12",X"80",X"03",X"FF",
		X"4B",X"12",X"03",X"FF",X"4B",X"12",X"03",X"FF",X"4F",X"12",X"03",X"FF",X"4F",X"12",X"03",X"FF",
		X"53",X"12",X"03",X"FF",X"53",X"12",X"03",X"FF",X"4F",X"12",X"03",X"FF",X"4F",X"12",X"01",X"FF",
		X"4B",X"12",X"03",X"01",X"3F",X"12",X"03",X"01",X"3F",X"12",X"03",X"01",X"43",X"12",X"03",X"01",
		X"43",X"12",X"03",X"01",X"47",X"12",X"03",X"01",X"47",X"12",X"03",X"01",X"43",X"12",X"03",X"01",
		X"43",X"12",X"01",X"01",X"3F",X"12",X"FD",X"FF",X"5B",X"12",X"FD",X"FF",X"5B",X"12",X"FD",X"FE",
		X"5B",X"12",X"FD",X"FE",X"5B",X"12",X"FD",X"FE",X"5B",X"12",X"FE",X"FD",X"5B",X"12",X"FE",X"FD",
		X"5B",X"12",X"FF",X"FD",X"5B",X"12",X"00",X"FD",X"5B",X"12",X"01",X"FD",X"5B",X"12",X"01",X"FD",
		X"5B",X"12",X"02",X"FE",X"5B",X"12",X"80",X"FD",X"01",X"57",X"12",X"FD",X"01",X"57",X"12",X"FD",
		X"02",X"57",X"12",X"FD",X"02",X"57",X"12",X"FD",X"02",X"57",X"12",X"FE",X"03",X"57",X"12",X"FE",
		X"03",X"57",X"12",X"FE",X"03",X"57",X"12",X"00",X"03",X"57",X"12",X"01",X"03",X"57",X"12",X"01",
		X"03",X"57",X"12",X"02",X"02",X"57",X"12",X"80",X"A0",X"B8",X"A0",X"68",X"A0",X"18",X"B8",X"70",
		X"B8",X"C0",X"D0",X"C0",X"D0",X"68",X"D0",X"40",X"03",X"10",X"8B",X"10",X"03",X"01",X"8B",X"10",
		X"03",X"01",X"8B",X"10",X"03",X"01",X"9F",X"10",X"03",X"02",X"9F",X"10",X"03",X"03",X"9F",X"10",
		X"02",X"03",X"9F",X"10",X"02",X"03",X"9F",X"10",X"01",X"03",X"8F",X"10",X"00",X"03",X"8F",X"10",
		X"01",X"02",X"8F",X"10",X"00",X"03",X"8F",X"10",X"80",X"22",X"FD",X"00",X"93",X"10",X"FD",X"01",
		X"93",X"10",X"FD",X"01",X"93",X"10",X"FD",X"01",X"A3",X"10",X"FD",X"02",X"A3",X"10",X"FE",X"03",
		X"A3",X"10",X"FE",X"03",X"A3",X"10",X"FE",X"03",X"A3",X"10",X"FF",X"03",X"8F",X"10",X"00",X"03",
		X"8F",X"10",X"FF",X"02",X"8F",X"10",X"00",X"02",X"8F",X"10",X"80",X"55",X"00",X"03",X"8F",X"10",
		X"FF",X"03",X"8F",X"10",X"FF",X"03",X"8F",X"10",X"FF",X"03",X"A3",X"10",X"FE",X"03",X"A3",X"10",
		X"FE",X"02",X"A3",X"10",X"FD",X"02",X"A3",X"10",X"FD",X"02",X"A3",X"10",X"FD",X"02",X"93",X"10",
		X"FD",X"00",X"93",X"10",X"FD",X"01",X"93",X"10",X"FD",X"00",X"93",X"10",X"FD",X"00",X"93",X"10",
		X"FD",X"FF",X"93",X"10",X"FD",X"FF",X"9B",X"10",X"FD",X"FE",X"9B",X"10",X"FD",X"FE",X"9B",X"10",
		X"FE",X"FD",X"9B",X"10",X"FE",X"FD",X"9B",X"10",X"FE",X"FD",X"8D",X"10",X"FF",X"FD",X"8D",X"10",
		X"FF",X"FD",X"8D",X"10",X"00",X"FD",X"8D",X"10",X"80",X"00",X"00",X"03",X"8F",X"10",X"01",X"03",
		X"8F",X"10",X"01",X"03",X"8F",X"10",X"01",X"03",X"9F",X"10",X"02",X"03",X"9F",X"10",X"02",X"02",
		X"9F",X"10",X"03",X"02",X"9F",X"10",X"03",X"02",X"9F",X"10",X"03",X"02",X"8B",X"10",X"03",X"00",
		X"8B",X"10",X"03",X"01",X"8B",X"10",X"03",X"00",X"8B",X"10",X"03",X"00",X"8B",X"10",X"03",X"FF",
		X"8B",X"10",X"03",X"FF",X"97",X"10",X"03",X"FE",X"97",X"10",X"03",X"FE",X"97",X"10",X"02",X"FD",
		X"97",X"10",X"02",X"FD",X"97",X"10",X"02",X"FD",X"8D",X"10",X"01",X"FD",X"8D",X"10",X"01",X"FD",
		X"8D",X"10",X"00",X"FD",X"8D",X"10",X"80",X"44",X"00",X"FD",X"8D",X"10",X"01",X"FD",X"8D",X"10",
		X"01",X"FD",X"8D",X"10",X"01",X"FD",X"97",X"10",X"02",X"FD",X"97",X"10",X"02",X"FE",X"97",X"10",
		X"02",X"FE",X"97",X"10",X"03",X"FE",X"97",X"10",X"03",X"FF",X"8B",X"10",X"03",X"FF",X"8B",X"10",
		X"03",X"FF",X"8B",X"10",X"03",X"00",X"8B",X"10",X"80",X"61",X"00",X"FD",X"8D",X"10",X"FF",X"FD",
		X"8D",X"10",X"FF",X"FD",X"8D",X"10",X"FF",X"FD",X"9B",X"10",X"FE",X"FD",X"9B",X"10",X"FE",X"FE",
		X"9B",X"10",X"FE",X"FE",X"9B",X"10",X"FD",X"FE",X"9B",X"10",X"FD",X"FF",X"93",X"10",X"FD",X"FF",
		X"93",X"10",X"FD",X"FF",X"93",X"10",X"FD",X"00",X"93",X"10",X"80",X"73",X"00",X"88",X"01",X"80",
		X"00",X"80",X"01",X"88",X"02",X"88",X"03",X"80",X"02",X"80",X"03",X"88",X"14",X"88",X"15",X"80",
		X"14",X"80",X"15",X"88",X"16",X"88",X"17",X"80",X"16",X"80",X"17",X"88",X"18",X"88",X"19",X"80",
		X"18",X"80",X"19",X"88",X"1A",X"88",X"1B",X"80",X"1A",X"80",X"1B",X"88",X"1C",X"88",X"1D",X"80",
		X"1C",X"80",X"1D",X"88",X"1E",X"88",X"1F",X"80",X"1E",X"80",X"1F",X"88",X"20",X"88",X"20",X"80",
		X"00",X"A0",X"62",X"9A",X"21",X"88",X"21",X"80",X"01",X"A0",X"62",X"9A",X"22",X"88",X"22",X"80",
		X"02",X"A0",X"62",X"9A",X"23",X"88",X"23",X"80",X"03",X"A0",X"62",X"9A",X"34",X"88",X"34",X"80",
		X"04",X"A0",X"62",X"9A",X"35",X"88",X"35",X"80",X"05",X"A0",X"62",X"9A",X"36",X"88",X"36",X"80",
		X"06",X"A0",X"62",X"9A",X"37",X"88",X"37",X"80",X"07",X"A0",X"62",X"9A",X"38",X"88",X"38",X"80",
		X"08",X"A0",X"62",X"9A",X"39",X"88",X"39",X"80",X"09",X"A0",X"62",X"9A",X"3A",X"88",X"3A",X"80",
		X"0A",X"A0",X"62",X"9A",X"3B",X"88",X"3B",X"80",X"0B",X"A0",X"62",X"9A",X"3C",X"88",X"3C",X"80",
		X"0C",X"A0",X"62",X"9A",X"3D",X"88",X"3D",X"80",X"0D",X"A0",X"62",X"9A",X"3E",X"88",X"3E",X"80",
		X"0E",X"A0",X"62",X"9A",X"3F",X"88",X"3F",X"80",X"0F",X"A0",X"62",X"9A",X"7F",X"7F",X"7F",X"7F",
		X"47",X"46",X"45",X"44",X"79",X"78",X"77",X"76",X"00",X"00",X"00",X"00",X"05",X"05",X"05",X"05",
		X"05",X"05",X"05",X"05",X"10",X"10",X"10",X"10",X"15",X"15",X"15",X"15",X"05",X"05",X"05",X"05",
		X"7A",X"7A",X"7A",X"7A",X"4A",X"46",X"45",X"49",X"79",X"78",X"77",X"76",X"00",X"00",X"00",X"00",
		X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"00",X"00",X"00",X"00",X"05",X"05",X"05",X"05",
		X"05",X"05",X"05",X"05",X"7F",X"7F",X"48",X"7F",X"47",X"46",X"45",X"44",X"7A",X"7A",X"7A",X"7A",
		X"00",X"00",X"01",X"00",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"10",X"10",X"11",X"10",
		X"15",X"05",X"05",X"15",X"05",X"05",X"05",X"05",X"7A",X"7A",X"4B",X"7A",X"4A",X"46",X"45",X"49",
		X"7A",X"7A",X"7A",X"7A",X"00",X"00",X"07",X"00",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",
		X"00",X"00",X"07",X"00",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"7F",X"51",X"4F",X"7F",
		X"53",X"52",X"50",X"4E",X"79",X"78",X"77",X"76",X"00",X"06",X"06",X"00",X"06",X"06",X"06",X"06",
		X"04",X"04",X"04",X"04",X"10",X"16",X"16",X"10",X"16",X"16",X"16",X"16",X"04",X"04",X"04",X"04",
		X"7A",X"5B",X"59",X"7A",X"5D",X"5C",X"5A",X"58",X"79",X"78",X"77",X"76",X"00",X"06",X"06",X"00",
		X"06",X"06",X"06",X"06",X"04",X"04",X"04",X"04",X"00",X"06",X"06",X"00",X"06",X"06",X"06",X"06",
		X"04",X"04",X"04",X"04",X"7F",X"7F",X"7F",X"7F",X"57",X"56",X"55",X"54",X"7A",X"7A",X"7A",X"7A",
		X"00",X"00",X"00",X"00",X"06",X"06",X"06",X"06",X"04",X"04",X"04",X"04",X"10",X"10",X"10",X"10",
		X"16",X"16",X"16",X"16",X"04",X"04",X"04",X"04",X"7A",X"7A",X"7A",X"7A",X"61",X"60",X"5F",X"5E",
		X"7A",X"7A",X"7A",X"7A",X"00",X"00",X"00",X"00",X"06",X"06",X"06",X"06",X"04",X"04",X"04",X"04",
		X"00",X"00",X"00",X"00",X"06",X"06",X"06",X"06",X"04",X"04",X"04",X"04",X"7F",X"65",X"63",X"7F",
		X"67",X"66",X"64",X"62",X"79",X"78",X"77",X"76",X"00",X"08",X"08",X"00",X"08",X"08",X"08",X"08",
		X"01",X"01",X"01",X"01",X"10",X"18",X"18",X"10",X"18",X"18",X"18",X"18",X"01",X"01",X"01",X"01",
		X"7A",X"6F",X"6D",X"7A",X"71",X"70",X"6E",X"6C",X"79",X"78",X"77",X"76",X"00",X"08",X"08",X"00",
		X"08",X"08",X"08",X"08",X"01",X"01",X"01",X"01",X"00",X"08",X"08",X"00",X"08",X"08",X"08",X"08",
		X"01",X"01",X"01",X"01",X"7F",X"7F",X"7F",X"7F",X"6B",X"6A",X"69",X"68",X"7A",X"7A",X"7A",X"7A",
		X"00",X"00",X"00",X"00",X"08",X"08",X"08",X"08",X"01",X"01",X"01",X"01",X"10",X"10",X"10",X"10",
		X"18",X"18",X"18",X"18",X"01",X"01",X"01",X"01",X"7A",X"7A",X"7A",X"7A",X"75",X"74",X"73",X"72",
		X"7A",X"7A",X"7A",X"7A",X"00",X"00",X"00",X"00",X"08",X"08",X"08",X"08",X"01",X"01",X"01",X"01",
		X"10",X"10",X"10",X"10",X"08",X"08",X"08",X"08",X"01",X"01",X"01",X"01",X"7F",X"D4",X"D2",X"7F",
		X"7F",X"D5",X"D3",X"7F",X"7A",X"7A",X"7A",X"7A",X"00",X"09",X"09",X"00",X"00",X"09",X"09",X"00",
		X"01",X"01",X"01",X"01",X"10",X"19",X"19",X"10",X"10",X"19",X"19",X"10",X"01",X"01",X"01",X"01",
		X"7A",X"D4",X"D2",X"7A",X"7A",X"D5",X"D3",X"7A",X"7A",X"7A",X"7A",X"7A",X"00",X"09",X"09",X"00",
		X"00",X"09",X"09",X"00",X"01",X"01",X"01",X"01",X"00",X"09",X"09",X"00",X"00",X"09",X"09",X"00",
		X"01",X"01",X"01",X"01",X"DC",X"DA",X"D8",X"D6",X"DD",X"DB",X"D9",X"D7",X"7A",X"7A",X"7A",X"7A",
		X"09",X"09",X"09",X"09",X"09",X"09",X"09",X"09",X"04",X"04",X"04",X"04",X"19",X"19",X"19",X"19",
		X"19",X"19",X"19",X"19",X"04",X"04",X"04",X"04",X"DC",X"DA",X"D8",X"D6",X"DD",X"DB",X"D9",X"D7",
		X"7A",X"7A",X"7A",X"7A",X"09",X"09",X"09",X"09",X"09",X"09",X"09",X"09",X"04",X"04",X"04",X"04",
		X"09",X"09",X"09",X"09",X"09",X"09",X"09",X"09",X"04",X"04",X"04",X"04",X"0D",X"87",X"CD",X"85",
		X"8D",X"84",X"2A",X"85",X"6A",X"86",X"27",X"87",X"C7",X"85",X"67",X"84",X"0F",X"FC",X"FC",X"00",
		X"0E",X"FC",X"00",X"00",X"0E",X"00",X"FC",X"00",X"0F",X"00",X"00",X"00",X"02",X"12",X"BC",X"BA",
		X"B8",X"B6",X"B4",X"BD",X"BB",X"B9",X"B7",X"B5",X"C6",X"C4",X"C2",X"C0",X"BE",X"C7",X"C5",X"C3",
		X"C1",X"BF",X"D0",X"CE",X"CC",X"CA",X"C8",X"D1",X"CF",X"CD",X"CB",X"C9",X"7F",X"B2",X"B0",X"AE",
		X"AC",X"7F",X"B3",X"B1",X"AF",X"AD",X"00",X"10",X"88",X"86",X"84",X"89",X"87",X"85",X"8E",X"8C",
		X"8A",X"8F",X"8D",X"8B",X"94",X"92",X"90",X"95",X"93",X"91",X"7F",X"82",X"80",X"7F",X"83",X"81",
		X"01",X"11",X"9E",X"9C",X"9A",X"9F",X"9D",X"9B",X"A4",X"A2",X"A0",X"A5",X"A3",X"A1",X"AA",X"A8",
		X"A6",X"AB",X"A9",X"A7",X"7F",X"98",X"96",X"7F",X"99",X"97",X"09",X"19",X"E6",X"E4",X"E2",X"E0",
		X"DE",X"E7",X"E5",X"E3",X"E1",X"DF",X"E6",X"E4",X"E2",X"E0",X"DE",X"E7",X"E5",X"E3",X"E1",X"DF",
		X"7F",X"DC",X"DA",X"D8",X"D6",X"7F",X"DD",X"DB",X"D9",X"D7",X"7F",X"DC",X"DA",X"D8",X"D6",X"7F",
		X"DD",X"DB",X"D9",X"D7",X"05",X"15",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"50",X"99",
		X"70",X"99",X"90",X"99",X"B0",X"99",X"D0",X"99",X"21",X"8A",X"48",X"C3",X"6D",X"2F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
