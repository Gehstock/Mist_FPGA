library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity snd_rom is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of snd_rom is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"06",X"00",X"21",X"00",X"40",X"C3",X"61",X"01",X"32",X"00",X"C0",X"32",X"01",X"C0",X"C9",X"FF",
		X"32",X"00",X"C0",X"32",X"03",X"C0",X"C9",X"FF",X"32",X"00",X"C0",X"32",X"04",X"C0",X"C9",X"FF",
		X"32",X"00",X"C0",X"32",X"01",X"C0",X"C9",X"FF",X"87",X"85",X"6F",X"7C",X"CE",X"00",X"67",X"7E",
		X"23",X"66",X"6F",X"E9",X"FF",X"FF",X"FF",X"FF",X"D9",X"08",X"CD",X"40",X"00",X"08",X"D9",X"C9",
		X"3A",X"00",X"60",X"47",X"FE",X"20",X"28",X"1A",X"FE",X"A0",X"28",X"16",X"E6",X"60",X"C0",X"78",
		X"FE",X"00",X"28",X"73",X"E6",X"7F",X"FE",X"0D",X"28",X"34",X"FE",X"0E",X"28",X"30",X"FE",X"01",
		X"28",X"2C",X"78",X"B7",X"FA",X"C1",X"00",X"FE",X"1D",X"28",X"05",X"FE",X"1C",X"C8",X"18",X"44",
		X"21",X"00",X"40",X"36",X"1D",X"23",X"36",X"00",X"23",X"36",X"1E",X"23",X"36",X"00",X"C9",X"21",
		X"00",X"40",X"36",X"1C",X"23",X"36",X"00",X"23",X"36",X"1E",X"23",X"36",X"00",X"C9",X"78",X"CB",
		X"7F",X"20",X"17",X"57",X"21",X"09",X"40",X"7E",X"BA",X"C8",X"B7",X"7E",X"C4",X"D9",X"00",X"7A",
		X"32",X"09",X"40",X"3E",X"01",X"32",X"08",X"40",X"78",X"C9",X"AF",X"32",X"08",X"40",X"32",X"09",
		X"40",X"78",X"18",X"0D",X"32",X"0A",X"40",X"3A",X"0A",X"40",X"47",X"B7",X"78",X"50",X"F2",X"F1",
		X"00",X"CB",X"BF",X"CD",X"D9",X"00",X"C9",X"21",X"00",X"40",X"06",X"06",X"AF",X"77",X"23",X"10",
		X"FC",X"AF",X"32",X"08",X"40",X"32",X"09",X"40",X"C9",X"47",X"21",X"00",X"40",X"BE",X"28",X"0B",
		X"23",X"23",X"BE",X"28",X"06",X"23",X"23",X"BE",X"28",X"01",X"C9",X"3E",X"00",X"77",X"23",X"77",
		X"C9",X"CD",X"15",X"01",X"20",X"1B",X"CD",X"15",X"01",X"20",X"15",X"21",X"00",X"40",X"1E",X"03",
		X"7E",X"1D",X"28",X"07",X"2C",X"2C",X"BE",X"38",X"F8",X"18",X"F5",X"BA",X"D0",X"CD",X"15",X"01",
		X"72",X"2C",X"36",X"00",X"C9",X"21",X"00",X"40",X"06",X"03",X"0E",X"04",X"BE",X"28",X"05",X"2C",
		X"2C",X"10",X"F9",X"41",X"79",X"90",X"C9",X"AF",X"4F",X"47",X"C3",X"87",X"01",X"3E",X"91",X"32",
		X"00",X"C0",X"32",X"01",X"C0",X"3D",X"20",X"FD",X"21",X"53",X"00",X"AF",X"37",X"1F",X"E6",X"E0",
		X"47",X"7D",X"E6",X"0F",X"B0",X"32",X"00",X"C0",X"32",X"01",X"C0",X"29",X"29",X"29",X"29",X"7C",
		X"E6",X"3F",X"00",X"00",X"00",X"00",X"32",X"00",X"C0",X"32",X"01",X"C0",X"C3",X"00",X"00",X"16",
		X"8B",X"ED",X"56",X"70",X"7E",X"B8",X"20",X"C5",X"23",X"7C",X"D6",X"44",X"20",X"F3",X"78",X"C6",
		X"55",X"47",X"D2",X"02",X"00",X"06",X"00",X"0E",X"00",X"21",X"00",X"40",X"71",X"7E",X"B8",X"20",
		X"AC",X"0C",X"FE",X"FF",X"28",X"A1",X"04",X"23",X"7C",X"D6",X"44",X"20",X"EF",X"11",X"00",X"00",
		X"21",X"00",X"00",X"06",X"00",X"1A",X"4F",X"09",X"13",X"7A",X"FE",X"20",X"20",X"F7",X"7C",X"FE",
		X"E9",X"20",X"8A",X"7D",X"FE",X"74",X"20",X"85",X"06",X"00",X"21",X"00",X"40",X"70",X"23",X"7C",
		X"D6",X"44",X"20",X"F9",X"F9",X"ED",X"56",X"3E",X"02",X"32",X"11",X"40",X"21",X"FF",X"A1",X"22",
		X"0B",X"40",X"77",X"DD",X"21",X"00",X"00",X"DD",X"21",X"00",X"00",X"FD",X"21",X"00",X"00",X"FD",
		X"21",X"00",X"00",X"3E",X"00",X"32",X"06",X"40",X"CD",X"F5",X"02",X"3E",X"01",X"32",X"06",X"40",
		X"CD",X"F5",X"02",X"3E",X"02",X"32",X"06",X"40",X"CD",X"F5",X"02",X"21",X"80",X"02",X"22",X"E9",
		X"40",X"18",X"00",X"FB",X"3A",X"00",X"80",X"21",X"11",X"40",X"A6",X"20",X"F7",X"3A",X"00",X"80",
		X"21",X"11",X"40",X"A6",X"28",X"F7",X"F3",X"3E",X"00",X"32",X"06",X"40",X"3A",X"01",X"40",X"B7",
		X"3A",X"00",X"40",X"28",X"05",X"CD",X"BE",X"02",X"18",X"03",X"CD",X"A6",X"02",X"FB",X"00",X"00",
		X"F3",X"3E",X"01",X"32",X"06",X"40",X"3A",X"03",X"40",X"B7",X"3A",X"02",X"40",X"28",X"05",X"CD",
		X"BE",X"02",X"18",X"03",X"CD",X"A6",X"02",X"FB",X"00",X"00",X"F3",X"3E",X"02",X"32",X"06",X"40",
		X"3A",X"05",X"40",X"B7",X"3A",X"04",X"40",X"28",X"05",X"CD",X"BE",X"02",X"18",X"06",X"CD",X"A6",
		X"02",X"C3",X"54",X"02",X"CD",X"59",X"02",X"18",X"98",X"3A",X"08",X"40",X"B7",X"C8",X"CD",X"72",
		X"02",X"C8",X"CD",X"82",X"02",X"C0",X"CD",X"92",X"02",X"D0",X"3A",X"09",X"40",X"77",X"23",X"AF",
		X"77",X"C9",X"3A",X"09",X"40",X"21",X"00",X"40",X"BE",X"C8",X"23",X"23",X"BE",X"C8",X"23",X"23",
		X"BE",X"C9",X"21",X"00",X"40",X"7E",X"B7",X"C8",X"23",X"23",X"7E",X"B7",X"C8",X"23",X"23",X"7E",
		X"B7",X"C9",X"3A",X"09",X"40",X"47",X"21",X"00",X"40",X"7E",X"B8",X"D8",X"23",X"23",X"7E",X"B8",
		X"D8",X"23",X"23",X"7E",X"B8",X"C9",X"F5",X"CD",X"F5",X"02",X"F1",X"E6",X"3F",X"21",X"FE",X"05",
		X"EF",X"B7",X"C2",X"C8",X"02",X"21",X"01",X"40",X"CD",X"E2",X"02",X"36",X"01",X"C9",X"B7",X"C8",
		X"E6",X"3F",X"21",X"5E",X"06",X"EF",X"B7",X"C8",X"57",X"3E",X"02",X"32",X"11",X"40",X"3E",X"01",
		X"CD",X"78",X"05",X"21",X"00",X"40",X"CD",X"E2",X"02",X"15",X"06",X"00",X"28",X"01",X"70",X"23",
		X"70",X"C9",X"01",X"00",X"00",X"3A",X"06",X"40",X"4F",X"06",X"00",X"09",X"09",X"C9",X"4B",X"4F",
		X"4E",X"41",X"4D",X"49",X"C9",X"3A",X"06",X"40",X"FE",X"01",X"28",X"21",X"FE",X"02",X"28",X"38",
		X"B7",X"C0",X"3E",X"9F",X"0E",X"20",X"06",X"04",X"CF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DD",X"21",X"00",X"00",X"FD",X"21",X"00",X"00",X"81",X"10",X"ED",X"AF",X"C9",X"3E",X"9F",X"0E",
		X"20",X"06",X"04",X"D7",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DD",X"21",X"00",X"00",X"FD",
		X"21",X"00",X"00",X"81",X"10",X"ED",X"AF",X"C9",X"3E",X"9F",X"0E",X"20",X"06",X"04",X"DF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"DD",X"21",X"00",X"00",X"FD",X"21",X"00",X"00",X"81",X"10",
		X"ED",X"AF",X"C9",X"3A",X"06",X"40",X"FE",X"01",X"28",X"1C",X"FE",X"02",X"28",X"22",X"B7",X"C0",
		X"06",X"03",X"DD",X"21",X"01",X"C0",X"22",X"0D",X"40",X"3E",X"04",X"90",X"CD",X"8A",X"03",X"2A",
		X"0D",X"40",X"29",X"10",X"F1",X"C9",X"06",X"03",X"DD",X"21",X"03",X"C0",X"CD",X"66",X"03",X"C9",
		X"06",X"03",X"DD",X"21",X"04",X"C0",X"CD",X"66",X"03",X"C9",X"3D",X"0F",X"0F",X"37",X"1F",X"E6",
		X"E0",X"4F",X"7D",X"E6",X"0F",X"B1",X"32",X"00",X"C0",X"DD",X"77",X"00",X"FD",X"21",X"00",X"00",
		X"FD",X"21",X"00",X"00",X"FD",X"21",X"00",X"00",X"29",X"29",X"29",X"29",X"7C",X"E6",X"3F",X"32",
		X"00",X"C0",X"DD",X"77",X"00",X"C9",X"47",X"3A",X"06",X"40",X"FE",X"01",X"DD",X"21",X"03",X"C0",
		X"28",X"0E",X"FE",X"02",X"DD",X"21",X"04",X"C0",X"28",X"06",X"B7",X"C0",X"DD",X"21",X"01",X"C0",
		X"78",X"CD",X"8A",X"03",X"C9",X"22",X"0D",X"40",X"EB",X"22",X"0F",X"40",X"3A",X"06",X"40",X"FE",
		X"01",X"DD",X"21",X"03",X"C0",X"28",X"0E",X"FE",X"02",X"DD",X"21",X"04",X"C0",X"28",X"06",X"B7",
		X"C0",X"DD",X"21",X"01",X"C0",X"2A",X"0D",X"40",X"3E",X"01",X"CD",X"8A",X"03",X"2A",X"0D",X"40",
		X"11",X"FF",X"FF",X"19",X"3E",X"02",X"CD",X"8A",X"03",X"2A",X"0D",X"40",X"29",X"3E",X"03",X"CD",
		X"8A",X"03",X"C9",X"22",X"0D",X"40",X"EB",X"22",X"0F",X"40",X"3A",X"06",X"40",X"FE",X"02",X"DD",
		X"21",X"04",X"C0",X"28",X"0E",X"FE",X"01",X"DD",X"21",X"03",X"C0",X"28",X"06",X"B7",X"DD",X"21",
		X"01",X"C0",X"C0",X"2A",X"0D",X"40",X"3E",X"01",X"CD",X"8A",X"03",X"2A",X"0F",X"40",X"EB",X"2A",
		X"0D",X"40",X"19",X"3E",X"02",X"CD",X"8A",X"03",X"2A",X"0F",X"40",X"EB",X"2A",X"0D",X"40",X"19",
		X"19",X"3E",X"03",X"CD",X"8A",X"03",X"C9",X"22",X"0D",X"40",X"EB",X"22",X"0F",X"40",X"3A",X"06",
		X"40",X"FE",X"02",X"DD",X"21",X"04",X"C0",X"28",X"0E",X"FE",X"01",X"DD",X"21",X"03",X"C0",X"28",
		X"06",X"B7",X"C0",X"DD",X"21",X"01",X"C0",X"2A",X"0D",X"40",X"3E",X"01",X"CD",X"8A",X"03",X"2A",
		X"0D",X"40",X"11",X"02",X"00",X"19",X"3E",X"02",X"CD",X"8A",X"03",X"2A",X"0D",X"40",X"29",X"3E",
		X"03",X"CD",X"8A",X"03",X"C9",X"3D",X"47",X"3E",X"0F",X"91",X"4F",X"3A",X"06",X"40",X"FE",X"02",
		X"28",X"10",X"FE",X"01",X"28",X"07",X"B7",X"C0",X"CD",X"B7",X"04",X"CF",X"C9",X"CD",X"B7",X"04",
		X"D7",X"C9",X"CD",X"B7",X"04",X"DF",X"C9",X"FD",X"21",X"00",X"00",X"FD",X"21",X"00",X"00",X"FD",
		X"21",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"58",X"21",X"D6",X"04",X"16",X"00",X"19",X"7E",
		X"47",X"79",X"E6",X"0F",X"B0",X"C9",X"90",X"B0",X"D0",X"F0",X"3E",X"0F",X"91",X"4F",X"3A",X"06",
		X"40",X"FE",X"01",X"DD",X"21",X"03",X"C0",X"28",X"0E",X"FE",X"02",X"DD",X"21",X"04",X"C0",X"28",
		X"06",X"B7",X"C0",X"DD",X"21",X"01",X"C0",X"1E",X"00",X"21",X"D6",X"04",X"16",X"00",X"19",X"46",
		X"79",X"E6",X"0F",X"4F",X"B0",X"32",X"00",X"C0",X"DD",X"77",X"00",X"00",X"00",X"00",X"00",X"FD",
		X"21",X"00",X"00",X"FD",X"21",X"00",X"00",X"FD",X"21",X"00",X"00",X"23",X"46",X"79",X"B0",X"32",
		X"00",X"C0",X"DD",X"77",X"00",X"00",X"00",X"00",X"00",X"FD",X"21",X"00",X"00",X"FD",X"21",X"00",
		X"00",X"FD",X"21",X"00",X"00",X"23",X"46",X"79",X"B0",X"32",X"00",X"C0",X"DD",X"77",X"00",X"FD",
		X"21",X"00",X"00",X"FD",X"21",X"00",X"00",X"FD",X"21",X"00",X"00",X"C9",X"FD",X"21",X"00",X"00",
		X"FD",X"21",X"00",X"00",X"FD",X"21",X"00",X"00",X"FE",X"08",X"D0",X"47",X"3A",X"06",X"40",X"FE",
		X"01",X"28",X"0B",X"FE",X"02",X"28",X"0C",X"B7",X"C0",X"78",X"F6",X"E0",X"CF",X"C9",X"78",X"F6",
		X"E0",X"D7",X"C9",X"78",X"F6",X"E0",X"DF",X"C9",X"E6",X"01",X"5F",X"3A",X"06",X"40",X"FE",X"01",
		X"28",X"24",X"FE",X"02",X"28",X"3C",X"B7",X"C0",X"2A",X"0B",X"40",X"CB",X"43",X"20",X"06",X"CB",
		X"9D",X"CB",X"A5",X"18",X"04",X"3E",X"18",X"B5",X"6F",X"22",X"0B",X"40",X"77",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"C9",X"2A",X"0B",X"40",X"CB",X"43",X"20",X"04",X"CB",X"BD",X"18",
		X"04",X"3E",X"80",X"B5",X"6F",X"22",X"0B",X"40",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C9",X"2A",X"0B",X"40",X"CB",X"43",X"20",X"04",X"CB",X"84",X"18",X"04",X"3E",X"01",X"B4",
		X"67",X"22",X"0B",X"40",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C9",X"21",X"FF",
		X"A1",X"22",X"0B",X"40",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C9",X"21",X"67",
		X"A0",X"22",X"0B",X"40",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C9",X"F5",X"02",
		X"DC",X"06",X"E6",X"08",X"FA",X"09",X"A9",X"0A",X"5B",X"0B",X"91",X"18",X"0B",X"0C",X"79",X"16",
		X"A2",X"0C",X"0D",X"0D",X"E4",X"0D",X"84",X"0E",X"28",X"08",X"81",X"07",X"7F",X"0F",X"50",X"10",
		X"CC",X"10",X"15",X"12",X"C1",X"12",X"23",X"13",X"F8",X"13",X"51",X"15",X"E2",X"15",X"BC",X"17",
		X"55",X"19",X"1B",X"1A",X"EE",X"1A",X"72",X"1B",X"07",X"1C",X"97",X"1C",X"05",X"17",X"EA",X"1C",
		X"97",X"1C",X"EA",X"1C",X"BE",X"06",X"BE",X"06",X"BE",X"06",X"BE",X"06",X"BE",X"06",X"BE",X"06",
		X"BE",X"06",X"BE",X"06",X"BE",X"06",X"BE",X"06",X"BE",X"06",X"BE",X"06",X"BE",X"06",X"00",X"00",
		X"20",X"07",X"14",X"09",X"1F",X"0A",X"ED",X"0A",X"8C",X"0B",X"C9",X"18",X"3D",X"0C",X"AA",X"16",
		X"D2",X"0C",X"3D",X"0D",X"1B",X"0E",X"B8",X"0E",X"69",X"08",X"B4",X"07",X"AA",X"0F",X"7B",X"10",
		X"21",X"11",X"54",X"12",X"07",X"13",X"69",X"13",X"2C",X"14",X"7E",X"15",X"11",X"16",X"08",X"18",
		X"97",X"19",X"84",X"1A",X"27",X"1B",X"9E",X"1B",X"36",X"1C",X"B5",X"1C",X"58",X"17",X"17",X"1D",
		X"B5",X"1C",X"17",X"1D",X"C1",X"06",X"C1",X"06",X"C1",X"06",X"C1",X"06",X"C1",X"06",X"C1",X"06",
		X"C1",X"06",X"C1",X"06",X"C1",X"06",X"C1",X"06",X"C1",X"06",X"C1",X"06",X"C1",X"06",X"3E",X"00",
		X"C9",X"3E",X"FF",X"C9",X"43",X"4F",X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"20",X"62",X"79",
		X"20",X"4B",X"4F",X"4E",X"41",X"4D",X"49",X"20",X"31",X"39",X"38",X"34",X"3E",X"00",X"CD",X"78",
		X"05",X"3E",X"01",X"0E",X"09",X"CD",X"95",X"04",X"3E",X"03",X"0E",X"02",X"CD",X"95",X"04",X"3E",
		X"04",X"0E",X"00",X"CD",X"95",X"04",X"3E",X"03",X"21",X"01",X"00",X"CD",X"B6",X"03",X"21",X"01",
		X"00",X"22",X"17",X"40",X"3E",X"01",X"CD",X"B6",X"03",X"21",X"01",X"00",X"22",X"19",X"40",X"21",
		X"0F",X"00",X"22",X"14",X"40",X"AF",X"32",X"12",X"40",X"32",X"13",X"40",X"32",X"16",X"40",X"C9",
		X"3A",X"12",X"40",X"2F",X"32",X"12",X"40",X"B7",X"20",X"48",X"2A",X"14",X"40",X"22",X"19",X"40",
		X"3E",X"01",X"CD",X"B6",X"03",X"3A",X"13",X"40",X"3D",X"32",X"13",X"40",X"E6",X"03",X"20",X"3C",
		X"3A",X"16",X"40",X"B7",X"20",X"13",X"2A",X"14",X"40",X"01",X"01",X"00",X"09",X"7D",X"FE",X"8F",
		X"38",X"05",X"3E",X"01",X"32",X"16",X"40",X"18",X"11",X"2A",X"14",X"40",X"01",X"FF",X"FF",X"09",
		X"7D",X"FE",X"0F",X"30",X"05",X"3E",X"00",X"32",X"16",X"40",X"22",X"14",X"40",X"3E",X"03",X"CD",
		X"B6",X"03",X"2A",X"17",X"40",X"3E",X"01",X"CD",X"B6",X"03",X"18",X"00",X"AF",X"C9",X"3E",X"FF",
		X"C9",X"3E",X"00",X"CD",X"78",X"05",X"21",X"18",X"00",X"CD",X"53",X"03",X"3E",X"01",X"0E",X"0A",
		X"CD",X"95",X"04",X"3E",X"02",X"0E",X"09",X"CD",X"95",X"04",X"3E",X"03",X"0E",X"08",X"CD",X"95",
		X"04",X"3E",X"18",X"32",X"1E",X"40",X"3E",X"0A",X"32",X"1D",X"40",X"3E",X"00",X"32",X"1B",X"40",
		X"32",X"1C",X"40",X"C9",X"3A",X"1B",X"40",X"2F",X"32",X"1B",X"40",X"B7",X"20",X"64",X"21",X"1C",
		X"40",X"35",X"7E",X"4F",X"06",X"00",X"21",X"00",X"03",X"09",X"3A",X"1E",X"40",X"47",X"7E",X"E6",
		X"01",X"80",X"6F",X"26",X"00",X"CD",X"53",X"03",X"3A",X"1C",X"40",X"4F",X"E6",X"07",X"20",X"42",
		X"06",X"FF",X"CB",X"69",X"20",X"02",X"06",X"01",X"3A",X"1E",X"40",X"80",X"32",X"1E",X"40",X"3A",
		X"1C",X"40",X"4F",X"E6",X"3F",X"20",X"2B",X"CB",X"69",X"3E",X"0B",X"20",X"02",X"3E",X"09",X"32",
		X"1D",X"40",X"4F",X"3E",X"01",X"CD",X"95",X"04",X"3A",X"1D",X"40",X"06",X"01",X"80",X"4F",X"3E",
		X"02",X"CD",X"95",X"04",X"3A",X"1D",X"40",X"06",X"FF",X"80",X"4F",X"3E",X"03",X"CD",X"95",X"04",
		X"18",X"00",X"3E",X"00",X"C9",X"3E",X"FF",X"C9",X"3E",X"00",X"CD",X"78",X"05",X"21",X"18",X"00",
		X"3E",X"01",X"CD",X"B6",X"03",X"0E",X"06",X"3E",X"01",X"CD",X"95",X"04",X"3E",X"0D",X"32",X"22",
		X"40",X"32",X"21",X"40",X"21",X"40",X"00",X"22",X"23",X"40",X"21",X"40",X"00",X"22",X"25",X"40",
		X"21",X"00",X"00",X"22",X"27",X"40",X"3E",X"10",X"32",X"29",X"40",X"3E",X"02",X"32",X"2A",X"40",
		X"3E",X"00",X"32",X"1F",X"40",X"32",X"20",X"40",X"C9",X"3A",X"1F",X"40",X"2F",X"32",X"1F",X"40",
		X"B7",X"20",X"6D",X"3A",X"20",X"40",X"3D",X"32",X"20",X"40",X"E6",X"00",X"20",X"62",X"2A",X"27",
		X"40",X"EB",X"2A",X"23",X"40",X"7D",X"C6",X"20",X"E6",X"FF",X"6F",X"22",X"23",X"40",X"19",X"3E",
		X"01",X"CD",X"B6",X"03",X"3A",X"21",X"40",X"3D",X"FE",X"0B",X"38",X"0B",X"32",X"21",X"40",X"4F",
		X"3E",X"01",X"CD",X"95",X"04",X"18",X"39",X"2A",X"23",X"40",X"EB",X"2A",X"25",X"40",X"22",X"23",
		X"40",X"3A",X"22",X"40",X"32",X"21",X"40",X"21",X"29",X"40",X"35",X"20",X"23",X"36",X"10",X"EB",
		X"22",X"25",X"40",X"11",X"00",X"00",X"2A",X"27",X"40",X"19",X"22",X"27",X"40",X"21",X"2A",X"40",
		X"35",X"20",X"0D",X"36",X"08",X"3A",X"22",X"40",X"4F",X"3E",X"01",X"CD",X"95",X"04",X"18",X"00",
		X"3E",X"00",X"C9",X"3E",X"FF",X"C9",X"3E",X"00",X"CD",X"78",X"05",X"11",X"00",X"00",X"21",X"04",
		X"00",X"CD",X"D5",X"03",X"0E",X"08",X"CD",X"DA",X"04",X"3E",X"08",X"32",X"2E",X"40",X"3E",X"09",
		X"32",X"2D",X"40",X"3E",X"01",X"32",X"2F",X"40",X"3E",X"00",X"32",X"30",X"40",X"32",X"2B",X"40",
		X"32",X"2C",X"40",X"C9",X"3A",X"2B",X"40",X"2F",X"32",X"2B",X"40",X"B7",X"C2",X"3D",X"09",X"3A",
		X"2C",X"40",X"3D",X"32",X"2C",X"40",X"3A",X"2D",X"40",X"06",X"66",X"80",X"E6",X"55",X"06",X"5F",
		X"80",X"32",X"2D",X"40",X"6F",X"26",X"00",X"11",X"00",X"00",X"CD",X"D5",X"03",X"3A",X"2F",X"40",
		X"3D",X"32",X"2F",X"40",X"C2",X"F4",X"09",X"3A",X"30",X"40",X"4F",X"06",X"00",X"21",X"7B",X"09",
		X"09",X"7E",X"FE",X"FF",X"CA",X"F7",X"09",X"5F",X"06",X"01",X"3A",X"2E",X"40",X"CB",X"7B",X"CA",
		X"64",X"09",X"06",X"FF",X"80",X"32",X"2E",X"40",X"4F",X"CB",X"BB",X"21",X"2F",X"40",X"73",X"3A",
		X"30",X"40",X"3C",X"32",X"30",X"40",X"CD",X"DA",X"04",X"18",X"79",X"01",X"01",X"01",X"02",X"02",
		X"03",X"03",X"82",X"82",X"82",X"82",X"82",X"83",X"83",X"83",X"02",X"02",X"02",X"02",X"02",X"03",
		X"03",X"03",X"96",X"96",X"96",X"96",X"16",X"16",X"16",X"16",X"96",X"96",X"96",X"96",X"16",X"16",
		X"16",X"98",X"98",X"98",X"98",X"18",X"18",X"18",X"9A",X"9A",X"9A",X"9A",X"1A",X"1A",X"1A",X"9C",
		X"9C",X"9C",X"9C",X"1C",X"1C",X"1C",X"9E",X"9E",X"9E",X"9E",X"1E",X"1E",X"1E",X"9E",X"9E",X"9E",
		X"9E",X"1E",X"1E",X"1E",X"9E",X"9E",X"9E",X"9E",X"1E",X"1E",X"1E",X"9E",X"9E",X"9E",X"9E",X"1E",
		X"1E",X"1E",X"9E",X"9E",X"9E",X"9E",X"1E",X"1E",X"1E",X"9E",X"9E",X"9E",X"9E",X"1E",X"1E",X"1E",
		X"9E",X"9E",X"9E",X"9E",X"1E",X"1E",X"1E",X"FF",X"B5",X"FF",X"B1",X"FF",X"B2",X"FF",X"BF",X"FF",
		X"B3",X"FF",X"B7",X"FF",X"3E",X"00",X"C9",X"3E",X"FF",X"C9",X"3E",X"00",X"CD",X"78",X"05",X"3E",
		X"01",X"0E",X"09",X"CD",X"95",X"04",X"21",X"05",X"00",X"CD",X"53",X"03",X"3E",X"0A",X"32",X"33",
		X"40",X"3E",X"FF",X"32",X"34",X"40",X"AF",X"32",X"31",X"40",X"32",X"32",X"40",X"18",X"4B",X"3A",
		X"31",X"40",X"2F",X"32",X"31",X"40",X"B7",X"20",X"41",X"3A",X"32",X"40",X"3D",X"32",X"32",X"40",
		X"E6",X"07",X"20",X"15",X"3A",X"34",X"40",X"3C",X"32",X"34",X"40",X"4F",X"06",X"00",X"21",X"6F",
		X"0A",X"09",X"7E",X"6F",X"26",X"00",X"CD",X"53",X"03",X"3A",X"32",X"40",X"E6",X"1F",X"20",X"1A",
		X"3A",X"33",X"40",X"3D",X"32",X"33",X"40",X"28",X"13",X"4F",X"3E",X"01",X"CD",X"95",X"04",X"3A",
		X"33",X"40",X"4F",X"3E",X"02",X"CD",X"95",X"04",X"18",X"00",X"AF",X"C9",X"3E",X"FF",X"C9",X"00",
		X"05",X"09",X"08",X"06",X"04",X"04",X"04",X"05",X"09",X"04",X"04",X"04",X"08",X"09",X"04",X"08",
		X"06",X"05",X"0B",X"0A",X"0B",X"04",X"06",X"05",X"04",X"04",X"0A",X"0A",X"0A",X"06",X"04",X"05",
		X"05",X"09",X"08",X"06",X"04",X"04",X"04",X"05",X"09",X"04",X"04",X"04",X"08",X"09",X"04",X"08",
		X"06",X"05",X"0B",X"0A",X"0B",X"04",X"06",X"05",X"00",X"3E",X"00",X"CD",X"78",X"05",X"3E",X"03",
		X"CD",X"4C",X"05",X"21",X"04",X"00",X"3E",X"03",X"CD",X"B6",X"03",X"21",X"01",X"00",X"3E",X"01",
		X"CD",X"B6",X"03",X"0E",X"0E",X"3E",X"04",X"CD",X"95",X"04",X"3E",X"0C",X"32",X"3C",X"40",X"0E",
		X"0C",X"3E",X"01",X"CD",X"95",X"04",X"21",X"02",X"00",X"22",X"38",X"40",X"21",X"02",X"00",X"22",
		X"3A",X"40",X"21",X"04",X"00",X"22",X"36",X"40",X"AF",X"32",X"35",X"40",X"C9",X"3A",X"35",X"40",
		X"CB",X"47",X"2A",X"38",X"40",X"20",X"03",X"2A",X"3A",X"40",X"3E",X"01",X"CD",X"B6",X"03",X"3A",
		X"35",X"40",X"3D",X"32",X"35",X"40",X"E6",X"0F",X"20",X"0F",X"2A",X"36",X"40",X"11",X"03",X"00",
		X"19",X"22",X"36",X"40",X"3E",X"03",X"CD",X"B6",X"03",X"3A",X"35",X"40",X"E6",X"01",X"20",X"11",
		X"2A",X"38",X"40",X"11",X"02",X"00",X"19",X"22",X"38",X"40",X"11",X"00",X"00",X"19",X"22",X"3A",
		X"40",X"3A",X"35",X"40",X"E6",X"7F",X"20",X"1D",X"3A",X"3C",X"40",X"3D",X"32",X"3C",X"40",X"28",
		X"17",X"4F",X"3E",X"01",X"CD",X"95",X"04",X"3A",X"3C",X"40",X"06",X"02",X"80",X"4F",X"3E",X"04",
		X"CD",X"95",X"04",X"18",X"00",X"3E",X"00",X"C9",X"3E",X"FF",X"C9",X"3E",X"00",X"CD",X"78",X"05",
		X"21",X"20",X"00",X"CD",X"53",X"03",X"0E",X"07",X"CD",X"DA",X"04",X"21",X"02",X"00",X"22",X"42",
		X"40",X"3E",X"0B",X"32",X"41",X"40",X"3E",X"00",X"32",X"44",X"40",X"3E",X"01",X"32",X"40",X"40",
		X"3E",X"00",X"32",X"3D",X"40",X"32",X"3E",X"40",X"32",X"3F",X"40",X"C9",X"3A",X"3D",X"40",X"2F",
		X"32",X"3D",X"40",X"B7",X"20",X"57",X"21",X"3E",X"40",X"35",X"7E",X"E6",X"0F",X"20",X"09",X"3A",
		X"41",X"40",X"3D",X"32",X"41",X"40",X"28",X"48",X"21",X"40",X"40",X"35",X"20",X"3F",X"3A",X"44",
		X"40",X"3E",X"01",X"32",X"44",X"40",X"77",X"3A",X"3F",X"40",X"2F",X"32",X"3F",X"40",X"B7",X"20",
		X"16",X"3A",X"41",X"40",X"06",X"00",X"80",X"4F",X"CD",X"DA",X"04",X"2A",X"42",X"40",X"11",X"04",
		X"00",X"19",X"22",X"42",X"40",X"18",X"11",X"3A",X"41",X"40",X"4F",X"CD",X"DA",X"04",X"2A",X"42",
		X"40",X"11",X"FD",X"FF",X"19",X"22",X"42",X"40",X"CD",X"53",X"03",X"18",X"00",X"3E",X"00",X"C9",
		X"3E",X"FF",X"C9",X"BD",X"B1",X"B0",X"A7",X"AE",X"B7",X"B9",X"B8",X"AC",X"E0",X"9E",X"87",X"E0",
		X"B5",X"B1",X"B2",X"BF",X"B3",X"B7",X"E0",X"CF",X"C7",X"C8",X"CC",X"3E",X"00",X"CD",X"78",X"05",
		X"21",X"20",X"00",X"3E",X"01",X"CD",X"B6",X"03",X"3E",X"01",X"0E",X"0F",X"CD",X"95",X"04",X"3E",
		X"0F",X"32",X"47",X"40",X"21",X"20",X"00",X"22",X"48",X"40",X"3E",X"00",X"32",X"4A",X"40",X"3E",
		X"16",X"32",X"4B",X"40",X"3E",X"00",X"32",X"45",X"40",X"32",X"46",X"40",X"C9",X"3A",X"4A",X"40",
		X"3C",X"FE",X"81",X"20",X"02",X"3E",X"00",X"32",X"4A",X"40",X"3A",X"45",X"40",X"2F",X"32",X"45",
		X"40",X"B7",X"20",X"48",X"3A",X"46",X"40",X"3D",X"32",X"46",X"40",X"47",X"E6",X"01",X"20",X"3C",
		X"CB",X"48",X"2A",X"48",X"40",X"3A",X"4A",X"40",X"5F",X"16",X"00",X"19",X"22",X"48",X"40",X"20",
		X"07",X"2A",X"48",X"40",X"11",X"20",X"00",X"19",X"3E",X"01",X"CD",X"B6",X"03",X"3A",X"4B",X"40",
		X"3D",X"32",X"4B",X"40",X"20",X"16",X"3E",X"0E",X"32",X"4B",X"40",X"3A",X"47",X"40",X"3D",X"32",
		X"47",X"40",X"28",X"0B",X"4F",X"3E",X"01",X"CD",X"95",X"04",X"18",X"00",X"3E",X"00",X"C9",X"3E",
		X"FF",X"C9",X"3E",X"00",X"CD",X"78",X"05",X"3E",X"02",X"32",X"50",X"40",X"3E",X"14",X"32",X"4F",
		X"40",X"3A",X"4F",X"40",X"FE",X"10",X"38",X"02",X"3E",X"0F",X"4F",X"3E",X"01",X"CD",X"95",X"04",
		X"3E",X"00",X"32",X"4E",X"40",X"21",X"40",X"00",X"22",X"4C",X"40",X"3E",X"01",X"CD",X"B6",X"03",
		X"AF",X"C9",X"21",X"50",X"40",X"35",X"20",X"21",X"36",X"02",X"3A",X"4E",X"40",X"06",X"01",X"80",
		X"32",X"4E",X"40",X"3A",X"4E",X"40",X"FE",X"59",X"28",X"11",X"4F",X"06",X"00",X"2A",X"4C",X"40",
		X"09",X"22",X"4C",X"40",X"3E",X"01",X"CD",X"B6",X"03",X"AF",X"C9",X"3A",X"4F",X"40",X"D6",X"02",
		X"38",X"08",X"28",X"06",X"32",X"4F",X"40",X"C3",X"B1",X"0C",X"3E",X"FF",X"C9",X"3E",X"00",X"CD",
		X"78",X"05",X"3E",X"02",X"32",X"55",X"40",X"3E",X"15",X"32",X"54",X"40",X"3A",X"54",X"40",X"FE",
		X"10",X"38",X"02",X"3E",X"0F",X"4F",X"3E",X"01",X"CD",X"95",X"04",X"3E",X"FF",X"32",X"53",X"40",
		X"21",X"31",X"00",X"22",X"51",X"40",X"3E",X"01",X"CD",X"B6",X"03",X"AF",X"C9",X"21",X"55",X"40",
		X"35",X"20",X"21",X"36",X"02",X"3A",X"53",X"40",X"06",X"01",X"80",X"32",X"53",X"40",X"3A",X"53",
		X"40",X"FE",X"5E",X"28",X"11",X"4F",X"06",X"00",X"2A",X"51",X"40",X"09",X"22",X"51",X"40",X"3E",
		X"01",X"CD",X"B6",X"03",X"AF",X"C9",X"3A",X"54",X"40",X"D6",X"02",X"38",X"08",X"28",X"06",X"32",
		X"54",X"40",X"C3",X"1C",X"0D",X"3E",X"FF",X"C9",X"3E",X"00",X"CD",X"78",X"05",X"3E",X"02",X"32",
		X"5A",X"40",X"0E",X"00",X"CD",X"DA",X"04",X"3E",X"0F",X"32",X"59",X"40",X"3E",X"00",X"32",X"58",
		X"40",X"21",X"40",X"00",X"22",X"56",X"40",X"3E",X"03",X"CD",X"B6",X"03",X"3A",X"59",X"40",X"4F",
		X"3E",X"03",X"CD",X"95",X"04",X"AF",X"C9",X"21",X"5A",X"40",X"35",X"20",X"21",X"36",X"02",X"3A",
		X"58",X"40",X"06",X"01",X"80",X"32",X"58",X"40",X"3A",X"58",X"40",X"FE",X"59",X"28",X"11",X"4F",
		X"06",X"00",X"2A",X"56",X"40",X"09",X"22",X"56",X"40",X"3E",X"03",X"CD",X"B6",X"03",X"AF",X"C9",
		X"3A",X"59",X"40",X"D6",X"03",X"DA",X"E1",X"0D",X"CA",X"E1",X"0D",X"32",X"59",X"40",X"C3",X"8C",
		X"0D",X"3E",X"FF",X"C9",X"3E",X"00",X"CD",X"78",X"05",X"21",X"80",X"00",X"3E",X"01",X"CD",X"B6",
		X"03",X"0E",X"0A",X"3E",X"01",X"CD",X"95",X"04",X"3E",X"0A",X"32",X"63",X"40",X"21",X"00",X"00",
		X"22",X"61",X"40",X"21",X"1A",X"00",X"22",X"5D",X"40",X"21",X"00",X"00",X"22",X"5F",X"40",X"3E",
		X"00",X"32",X"5B",X"40",X"32",X"64",X"40",X"32",X"5C",X"40",X"C9",X"3A",X"5B",X"40",X"2F",X"32",
		X"5B",X"40",X"B7",X"20",X"59",X"3A",X"5C",X"40",X"3D",X"32",X"5C",X"40",X"21",X"64",X"40",X"7E",
		X"B7",X"20",X"33",X"3A",X"5C",X"40",X"FE",X"A0",X"30",X"01",X"34",X"47",X"E6",X"03",X"20",X"3E",
		X"CB",X"50",X"20",X"0C",X"11",X"FF",X"FF",X"2A",X"61",X"40",X"19",X"22",X"61",X"40",X"18",X"0A",
		X"11",X"02",X"00",X"2A",X"5F",X"40",X"19",X"22",X"5F",X"40",X"EB",X"2A",X"5D",X"40",X"19",X"3E",
		X"01",X"CD",X"B6",X"03",X"18",X"18",X"3A",X"5C",X"40",X"E6",X"0F",X"20",X"11",X"3A",X"63",X"40",
		X"3D",X"32",X"63",X"40",X"28",X"0B",X"4F",X"3E",X"01",X"CD",X"95",X"04",X"18",X"00",X"3E",X"00",
		X"C9",X"3E",X"FF",X"C9",X"3E",X"00",X"CD",X"78",X"05",X"3E",X"03",X"21",X"01",X"00",X"CD",X"B6",
		X"03",X"3E",X"04",X"0E",X"04",X"CD",X"95",X"04",X"3E",X"07",X"CD",X"4C",X"05",X"3E",X"04",X"32",
		X"6A",X"40",X"21",X"01",X"00",X"22",X"67",X"40",X"3E",X"08",X"32",X"69",X"40",X"AF",X"32",X"6B",
		X"40",X"32",X"65",X"40",X"32",X"66",X"40",X"C9",X"3A",X"65",X"40",X"2F",X"32",X"65",X"40",X"B7",
		X"C2",X"79",X"0F",X"3A",X"6B",X"40",X"B7",X"20",X"7C",X"3A",X"66",X"40",X"3D",X"32",X"66",X"40",
		X"FE",X"C0",X"28",X"59",X"FE",X"E0",X"38",X"12",X"E6",X"03",X"C2",X"79",X"0F",X"3A",X"69",X"40",
		X"3C",X"32",X"69",X"40",X"4F",X"3E",X"04",X"CD",X"95",X"04",X"3A",X"66",X"40",X"FE",X"E8",X"D2",
		X"79",X"0F",X"3A",X"6A",X"40",X"3D",X"32",X"6A",X"40",X"3A",X"66",X"40",X"E6",X"07",X"20",X"0F",
		X"2A",X"67",X"40",X"11",X"08",X"00",X"19",X"22",X"67",X"40",X"3E",X"03",X"CD",X"B6",X"03",X"3A",
		X"6A",X"40",X"B7",X"20",X"64",X"3E",X"10",X"32",X"6A",X"40",X"3A",X"69",X"40",X"3D",X"32",X"69",
		X"40",X"FE",X"02",X"28",X"57",X"4F",X"3E",X"04",X"CD",X"95",X"04",X"18",X"4C",X"3E",X"01",X"32",
		X"6B",X"40",X"21",X"04",X"00",X"22",X"67",X"40",X"3E",X"0B",X"32",X"69",X"40",X"4F",X"3E",X"04",
		X"CD",X"95",X"04",X"18",X"34",X"3A",X"66",X"40",X"3D",X"32",X"66",X"40",X"E6",X"0F",X"20",X"29",
		X"2A",X"67",X"40",X"11",X"02",X"00",X"19",X"22",X"67",X"40",X"3E",X"03",X"CD",X"B6",X"03",X"3A",
		X"66",X"40",X"E6",X"3F",X"20",X"13",X"3A",X"69",X"40",X"3D",X"32",X"69",X"40",X"FE",X"03",X"28",
		X"0B",X"4F",X"3E",X"04",X"CD",X"95",X"04",X"18",X"00",X"3E",X"00",X"C9",X"3E",X"FF",X"C9",X"3E",
		X"00",X"CD",X"78",X"05",X"21",X"10",X"00",X"CD",X"53",X"03",X"0E",X"0E",X"CD",X"DA",X"04",X"3E",
		X"08",X"32",X"70",X"40",X"3E",X"08",X"32",X"6F",X"40",X"3E",X"0F",X"32",X"6E",X"40",X"3E",X"00",
		X"32",X"71",X"40",X"32",X"6C",X"40",X"32",X"6D",X"40",X"C9",X"3A",X"6D",X"40",X"3D",X"32",X"6D",
		X"40",X"3A",X"71",X"40",X"B7",X"20",X"55",X"3A",X"70",X"40",X"4F",X"3A",X"6F",X"40",X"06",X"04",
		X"80",X"E6",X"0F",X"32",X"6F",X"40",X"81",X"6F",X"26",X"00",X"CD",X"53",X"03",X"3A",X"6D",X"40",
		X"E6",X"07",X"20",X"76",X"3A",X"70",X"40",X"06",X"04",X"80",X"32",X"70",X"40",X"E6",X"07",X"20",
		X"69",X"3A",X"6E",X"40",X"3D",X"32",X"6E",X"40",X"FE",X"02",X"28",X"06",X"4F",X"CD",X"DA",X"04",
		X"18",X"58",X"3E",X"01",X"32",X"71",X"40",X"3E",X"09",X"32",X"6E",X"40",X"4F",X"CD",X"DA",X"04",
		X"3E",X"08",X"32",X"70",X"40",X"3E",X"08",X"32",X"6F",X"40",X"18",X"3E",X"3A",X"70",X"40",X"4F",
		X"3A",X"6F",X"40",X"06",X"04",X"80",X"E6",X"0F",X"32",X"6F",X"40",X"81",X"6F",X"26",X"00",X"CD",
		X"53",X"03",X"3A",X"6D",X"40",X"E6",X"1F",X"20",X"21",X"3A",X"70",X"40",X"06",X"01",X"80",X"32",
		X"70",X"40",X"3A",X"6D",X"40",X"E6",X"7F",X"20",X"11",X"3A",X"6E",X"40",X"3D",X"32",X"6E",X"40",
		X"FE",X"02",X"28",X"09",X"4F",X"CD",X"DA",X"04",X"18",X"00",X"3E",X"00",X"C9",X"3E",X"FF",X"C9",
		X"3E",X"00",X"CD",X"78",X"05",X"21",X"72",X"40",X"36",X"00",X"3E",X"03",X"32",X"74",X"40",X"21",
		X"74",X"40",X"35",X"28",X"40",X"0E",X"0F",X"3E",X"01",X"CD",X"95",X"04",X"3E",X"C8",X"32",X"73",
		X"40",X"21",X"C8",X"00",X"3E",X"01",X"CD",X"B6",X"03",X"AF",X"C9",X"21",X"72",X"40",X"35",X"7E",
		X"28",X"DD",X"E6",X"7F",X"0E",X"0B",X"28",X"DF",X"57",X"E6",X"07",X"20",X"13",X"7A",X"0F",X"0F",
		X"0F",X"ED",X"44",X"21",X"73",X"40",X"86",X"77",X"6F",X"26",X"00",X"3E",X"01",X"CD",X"B6",X"03",
		X"AF",X"C9",X"3E",X"00",X"C9",X"3E",X"FF",X"C9",X"3E",X"00",X"C9",X"3E",X"FF",X"C9",X"3E",X"00",
		X"C9",X"3E",X"FF",X"C9",X"BD",X"B1",X"B0",X"A7",X"AE",X"B7",X"B9",X"B8",X"AC",X"E0",X"9E",X"87",
		X"E0",X"B5",X"B1",X"B2",X"BF",X"B3",X"B7",X"E0",X"CF",X"C7",X"C8",X"CC",X"3E",X"00",X"CD",X"78",
		X"05",X"3E",X"03",X"0E",X"00",X"CD",X"95",X"04",X"3E",X"03",X"CD",X"B6",X"03",X"3E",X"04",X"0E",
		X"0F",X"CD",X"95",X"04",X"3E",X"07",X"CD",X"4C",X"05",X"21",X"FF",X"02",X"3E",X"01",X"CD",X"B6",
		X"03",X"21",X"40",X"03",X"3E",X"02",X"CD",X"B6",X"03",X"3E",X"01",X"0E",X"00",X"CD",X"95",X"04",
		X"3E",X"02",X"0E",X"00",X"CD",X"95",X"04",X"3E",X"0F",X"32",X"79",X"40",X"21",X"04",X"00",X"22",
		X"77",X"40",X"3E",X"00",X"32",X"75",X"40",X"32",X"7B",X"40",X"32",X"7A",X"40",X"32",X"76",X"40",
		X"C9",X"3A",X"75",X"40",X"2F",X"32",X"75",X"40",X"B7",X"C2",X"0F",X"12",X"3A",X"76",X"40",X"3D",
		X"32",X"76",X"40",X"3A",X"7A",X"40",X"B7",X"20",X"75",X"3A",X"76",X"40",X"FE",X"D8",X"38",X"24",
		X"E6",X"07",X"C2",X"0F",X"12",X"3A",X"79",X"40",X"3D",X"32",X"79",X"40",X"4F",X"3E",X"04",X"CD",
		X"95",X"04",X"2A",X"77",X"40",X"11",X"05",X"00",X"19",X"22",X"77",X"40",X"3E",X"03",X"CD",X"B6",
		X"03",X"C3",X"0F",X"12",X"E6",X"07",X"C2",X"0F",X"12",X"3A",X"79",X"40",X"3C",X"FE",X"0F",X"20",
		X"11",X"32",X"79",X"40",X"4F",X"3E",X"04",X"CD",X"95",X"04",X"3E",X"01",X"32",X"7A",X"40",X"C3",
		X"0F",X"12",X"32",X"79",X"40",X"4F",X"3E",X"04",X"CD",X"95",X"04",X"3A",X"79",X"40",X"4F",X"3E",
		X"01",X"CD",X"95",X"04",X"3A",X"79",X"40",X"4F",X"3E",X"02",X"CD",X"95",X"04",X"2A",X"77",X"40",
		X"11",X"FD",X"FF",X"19",X"22",X"77",X"40",X"3E",X"03",X"CD",X"B6",X"03",X"18",X"61",X"3A",X"76",
		X"40",X"4F",X"06",X"00",X"21",X"00",X"02",X"09",X"46",X"23",X"7E",X"E6",X"7F",X"32",X"7B",X"40",
		X"26",X"02",X"78",X"E6",X"7F",X"6F",X"3E",X"01",X"CD",X"B6",X"03",X"3A",X"7B",X"40",X"6F",X"26",
		X"02",X"3E",X"02",X"CD",X"B6",X"03",X"3A",X"76",X"40",X"E6",X"1F",X"20",X"32",X"3A",X"79",X"40",
		X"3D",X"32",X"79",X"40",X"28",X"2C",X"4F",X"3E",X"04",X"CD",X"95",X"04",X"3A",X"79",X"40",X"4F",
		X"3E",X"01",X"CD",X"95",X"04",X"3A",X"79",X"40",X"4F",X"3E",X"02",X"CD",X"95",X"04",X"2A",X"77",
		X"40",X"11",X"FF",X"FF",X"19",X"22",X"77",X"40",X"3E",X"03",X"CD",X"B6",X"03",X"18",X"00",X"3E",
		X"00",X"C9",X"3E",X"FF",X"C9",X"3E",X"00",X"CD",X"78",X"05",X"21",X"08",X"00",X"3E",X"01",X"CD",
		X"53",X"03",X"0E",X"0D",X"3E",X"01",X"CD",X"95",X"04",X"0E",X"0D",X"3E",X"02",X"CD",X"95",X"04",
		X"3E",X"0D",X"32",X"80",X"40",X"3E",X"0D",X"32",X"81",X"40",X"3E",X"0D",X"32",X"84",X"40",X"21",
		X"08",X"00",X"22",X"7E",X"40",X"21",X"04",X"00",X"22",X"82",X"40",X"3E",X"00",X"32",X"7C",X"40",
		X"32",X"7D",X"40",X"C9",X"3A",X"7C",X"40",X"2F",X"32",X"7C",X"40",X"B7",X"20",X"5D",X"3A",X"7D",
		X"40",X"3D",X"32",X"7D",X"40",X"E6",X"03",X"20",X"52",X"21",X"84",X"40",X"35",X"21",X"80",X"40",
		X"35",X"20",X"1D",X"3E",X"0D",X"32",X"84",X"40",X"3A",X"81",X"40",X"3D",X"32",X"81",X"40",X"28",
		X"3D",X"32",X"80",X"40",X"21",X"02",X"00",X"22",X"7E",X"40",X"21",X"04",X"00",X"22",X"82",X"40",
		X"3A",X"84",X"40",X"4F",X"3E",X"01",X"CD",X"95",X"04",X"3A",X"84",X"40",X"4F",X"3E",X"02",X"CD",
		X"95",X"04",X"2A",X"82",X"40",X"11",X"02",X"00",X"19",X"22",X"82",X"40",X"EB",X"2A",X"7E",X"40",
		X"19",X"22",X"7E",X"40",X"3E",X"01",X"CD",X"53",X"03",X"18",X"00",X"3E",X"00",X"C9",X"3E",X"FF",
		X"C9",X"3E",X"00",X"CD",X"78",X"05",X"3E",X"04",X"32",X"87",X"40",X"3E",X"0F",X"32",X"88",X"40",
		X"3A",X"87",X"40",X"3D",X"32",X"87",X"40",X"20",X"18",X"3E",X"04",X"32",X"87",X"40",X"3A",X"88",
		X"40",X"FE",X"0D",X"06",X"FF",X"30",X"02",X"06",X"FE",X"80",X"32",X"88",X"40",X"FE",X"04",X"28",
		X"2F",X"3A",X"88",X"40",X"4F",X"3E",X"01",X"CD",X"95",X"04",X"21",X"20",X"00",X"22",X"85",X"40",
		X"3E",X"01",X"CD",X"B6",X"03",X"AF",X"C9",X"2A",X"85",X"40",X"01",X"08",X"00",X"09",X"7C",X"FE",
		X"07",X"28",X"BD",X"22",X"85",X"40",X"3E",X"01",X"CD",X"B6",X"03",X"AF",X"C9",X"3E",X"00",X"C9",
		X"3E",X"FF",X"C9",X"3E",X"00",X"CD",X"78",X"05",X"21",X"18",X"00",X"3E",X"01",X"CD",X"B6",X"03",
		X"0E",X"0D",X"3E",X"01",X"CD",X"95",X"04",X"3E",X"0B",X"32",X"91",X"40",X"3E",X"0D",X"32",X"8C",
		X"40",X"32",X"8B",X"40",X"21",X"10",X"00",X"22",X"8D",X"40",X"21",X"10",X"00",X"22",X"8F",X"40",
		X"21",X"00",X"00",X"22",X"92",X"40",X"3E",X"01",X"32",X"94",X"40",X"3E",X"02",X"32",X"95",X"40",
		X"3E",X"00",X"32",X"89",X"40",X"32",X"8A",X"40",X"C9",X"3A",X"89",X"40",X"2F",X"32",X"89",X"40",
		X"B7",X"20",X"7F",X"3A",X"8A",X"40",X"3D",X"32",X"8A",X"40",X"E6",X"01",X"20",X"74",X"2A",X"92",
		X"40",X"EB",X"2A",X"8D",X"40",X"7D",X"C6",X"21",X"E6",X"3F",X"6F",X"19",X"22",X"8D",X"40",X"19",
		X"22",X"8D",X"40",X"3E",X"01",X"CD",X"B6",X"03",X"3A",X"8B",X"40",X"3D",X"21",X"91",X"40",X"BE",
		X"38",X"0B",X"32",X"8B",X"40",X"4F",X"3E",X"01",X"CD",X"95",X"04",X"18",X"45",X"2A",X"8D",X"40",
		X"EB",X"2A",X"8F",X"40",X"22",X"8D",X"40",X"3A",X"8C",X"40",X"32",X"8B",X"40",X"21",X"94",X"40",
		X"35",X"20",X"2F",X"36",X"02",X"EB",X"22",X"8F",X"40",X"11",X"00",X"00",X"2A",X"92",X"40",X"19",
		X"22",X"92",X"40",X"21",X"95",X"40",X"35",X"20",X"19",X"36",X"12",X"21",X"91",X"40",X"35",X"3A",
		X"8C",X"40",X"3D",X"32",X"8C",X"40",X"FE",X"04",X"28",X"0B",X"4F",X"3E",X"01",X"CD",X"95",X"04",
		X"18",X"00",X"3E",X"00",X"C9",X"3E",X"FF",X"C9",X"3E",X"00",X"32",X"9D",X"40",X"3E",X"5E",X"32",
		X"9C",X"40",X"3E",X"00",X"CD",X"78",X"05",X"21",X"FF",X"02",X"3E",X"01",X"CD",X"B6",X"03",X"0E",
		X"0C",X"3E",X"01",X"CD",X"95",X"04",X"21",X"FF",X"01",X"22",X"9A",X"40",X"21",X"FF",X"01",X"22",
		X"98",X"40",X"3E",X"06",X"32",X"96",X"40",X"AF",X"32",X"97",X"40",X"C9",X"3A",X"9D",X"40",X"FE",
		X"00",X"28",X"0C",X"FE",X"01",X"CA",X"97",X"14",X"FE",X"02",X"CA",X"D0",X"14",X"18",X"4D",X"3A",
		X"96",X"40",X"3D",X"32",X"96",X"40",X"20",X"44",X"3E",X"06",X"32",X"96",X"40",X"3A",X"97",X"40",
		X"B7",X"20",X"16",X"2A",X"9A",X"40",X"11",X"FE",X"FF",X"19",X"22",X"9A",X"40",X"22",X"98",X"40",
		X"3A",X"9C",X"40",X"3D",X"32",X"9C",X"40",X"28",X"26",X"CD",X"6E",X"14",X"18",X"1E",X"3A",X"97",
		X"40",X"3C",X"FE",X"05",X"20",X"02",X"3E",X"FE",X"32",X"97",X"40",X"2A",X"98",X"40",X"CB",X"3C",
		X"AF",X"CB",X"1D",X"22",X"98",X"40",X"3E",X"01",X"CD",X"B6",X"03",X"C9",X"3E",X"00",X"C9",X"3E",
		X"01",X"32",X"9D",X"40",X"3E",X"00",X"C9",X"3E",X"02",X"32",X"A3",X"40",X"3E",X"0F",X"32",X"A2",
		X"40",X"21",X"40",X"00",X"3E",X"01",X"CD",X"B6",X"03",X"0E",X"0F",X"3E",X"01",X"CD",X"95",X"04",
		X"3A",X"A3",X"40",X"3D",X"32",X"A3",X"40",X"3E",X"0F",X"32",X"A2",X"40",X"21",X"40",X"00",X"22",
		X"A0",X"40",X"3E",X"02",X"32",X"9D",X"40",X"3E",X"00",X"32",X"9E",X"40",X"32",X"9F",X"40",X"C9",
		X"3A",X"9E",X"40",X"2F",X"32",X"9E",X"40",X"B7",X"20",X"6B",X"3A",X"9F",X"40",X"3D",X"32",X"9F",
		X"40",X"47",X"E6",X"03",X"20",X"5F",X"CB",X"50",X"28",X"18",X"11",X"04",X"00",X"CB",X"58",X"20",
		X"03",X"11",X"FC",X"FF",X"2A",X"A0",X"40",X"19",X"22",X"A0",X"40",X"3E",X"01",X"CD",X"B6",X"03",
		X"18",X"43",X"2A",X"A0",X"40",X"11",X"20",X"00",X"19",X"3E",X"01",X"CD",X"B6",X"03",X"3A",X"9F",
		X"40",X"E6",X"1F",X"20",X"0A",X"2A",X"A0",X"40",X"11",X"FE",X"FF",X"19",X"22",X"A0",X"40",X"3A",
		X"9F",X"40",X"E6",X"3F",X"20",X"1F",X"3A",X"A2",X"40",X"3D",X"32",X"A2",X"40",X"FE",X"08",X"28",
		X"17",X"4F",X"FE",X"0E",X"C2",X"3E",X"15",X"3A",X"A3",X"40",X"B7",X"C2",X"A1",X"14",X"3E",X"01",
		X"CD",X"95",X"04",X"18",X"00",X"3E",X"00",X"C9",X"3E",X"FF",X"C9",X"3E",X"00",X"C9",X"3E",X"FF",
		X"C9",X"3E",X"00",X"CD",X"78",X"05",X"21",X"C0",X"00",X"11",X"30",X"00",X"CD",X"D5",X"03",X"0E",
		X"0B",X"CD",X"DA",X"04",X"3E",X"03",X"0E",X"0C",X"CD",X"95",X"04",X"3E",X"0B",X"32",X"A7",X"40",
		X"3E",X"78",X"32",X"A6",X"40",X"3E",X"00",X"32",X"A4",X"40",X"32",X"A5",X"40",X"C9",X"3A",X"A4",
		X"40",X"2F",X"32",X"A4",X"40",X"B7",X"20",X"54",X"3A",X"A5",X"40",X"3D",X"32",X"A5",X"40",X"E6",
		X"07",X"20",X"08",X"3A",X"A6",X"40",X"C6",X"F9",X"32",X"A6",X"40",X"3A",X"A5",X"40",X"E6",X"03",
		X"20",X"15",X"3A",X"A6",X"40",X"C6",X"03",X"32",X"A6",X"40",X"FE",X"24",X"38",X"31",X"6F",X"26",
		X"00",X"11",X"30",X"00",X"CD",X"D5",X"03",X"3A",X"A5",X"40",X"47",X"E6",X"01",X"20",X"1D",X"CB",
		X"48",X"0E",X"0A",X"20",X"02",X"0E",X"0C",X"79",X"32",X"A7",X"40",X"CD",X"DA",X"04",X"3A",X"A7",
		X"40",X"06",X"01",X"80",X"4F",X"3E",X"03",X"CD",X"95",X"04",X"18",X"00",X"3E",X"00",X"C9",X"3E",
		X"FF",X"C9",X"3E",X"00",X"CD",X"78",X"05",X"3E",X"20",X"32",X"AF",X"40",X"3E",X"02",X"32",X"A8",
		X"40",X"3E",X"04",X"32",X"AE",X"40",X"3E",X"0E",X"32",X"AD",X"40",X"4F",X"3E",X"01",X"CD",X"95",
		X"04",X"21",X"08",X"00",X"22",X"A9",X"40",X"22",X"AB",X"40",X"3E",X"01",X"CD",X"B6",X"03",X"AF",
		X"C9",X"21",X"A8",X"40",X"35",X"20",X"2A",X"36",X"01",X"2A",X"A9",X"40",X"7D",X"C6",X"80",X"6F",
		X"22",X"A9",X"40",X"3E",X"01",X"CD",X"B6",X"03",X"21",X"AE",X"40",X"35",X"20",X"13",X"36",X"05",
		X"3A",X"AD",X"40",X"3D",X"FE",X"05",X"28",X"0B",X"32",X"AD",X"40",X"4F",X"3E",X"01",X"CD",X"95",
		X"04",X"AF",X"C9",X"3E",X"0E",X"32",X"AD",X"40",X"2A",X"AB",X"40",X"11",X"01",X"00",X"19",X"22",
		X"AB",X"40",X"22",X"A9",X"40",X"21",X"AF",X"40",X"35",X"CA",X"E2",X"15",X"AF",X"C9",X"3E",X"FF",
		X"C9",X"BD",X"B1",X"B0",X"A7",X"AE",X"B7",X"B9",X"B8",X"AC",X"E0",X"9E",X"87",X"E0",X"B5",X"B1",
		X"B2",X"BF",X"B3",X"B7",X"E0",X"CF",X"C7",X"C8",X"CC",X"3E",X"00",X"CD",X"78",X"05",X"11",X"01",
		X"00",X"21",X"48",X"00",X"CD",X"57",X"04",X"0E",X"0E",X"CD",X"DA",X"04",X"21",X"00",X"00",X"22",
		X"B5",X"40",X"3E",X"28",X"32",X"B4",X"40",X"3E",X"0D",X"32",X"B3",X"40",X"3E",X"03",X"32",X"B2",
		X"40",X"3E",X"00",X"32",X"B0",X"40",X"32",X"B1",X"40",X"C9",X"3A",X"B0",X"40",X"2F",X"32",X"B0",
		X"40",X"B7",X"20",X"4B",X"3A",X"B1",X"40",X"3D",X"32",X"B1",X"40",X"3A",X"B2",X"40",X"06",X"40",
		X"80",X"E6",X"3C",X"06",X"48",X"80",X"32",X"B2",X"40",X"6F",X"26",X"00",X"EB",X"2A",X"B5",X"40",
		X"19",X"11",X"02",X"00",X"CD",X"57",X"04",X"3A",X"B1",X"40",X"E6",X"FF",X"20",X"0A",X"2A",X"B5",
		X"40",X"11",X"00",X"00",X"19",X"22",X"B5",X"40",X"21",X"B4",X"40",X"35",X"20",X"11",X"36",X"28",
		X"20",X"0D",X"3A",X"B3",X"40",X"3D",X"32",X"B3",X"40",X"28",X"07",X"4F",X"CD",X"DA",X"04",X"3E",
		X"00",X"C9",X"3E",X"FF",X"C9",X"3E",X"00",X"CD",X"78",X"05",X"21",X"01",X"00",X"11",X"00",X"00",
		X"CD",X"13",X"04",X"0E",X"00",X"3E",X"03",X"CD",X"95",X"04",X"0E",X"0F",X"3E",X"01",X"CD",X"95",
		X"04",X"3E",X"02",X"0E",X"0F",X"CD",X"95",X"04",X"3E",X"10",X"32",X"C0",X"40",X"3A",X"C0",X"40",
		X"3D",X"32",X"C0",X"40",X"32",X"BF",X"40",X"FE",X"08",X"CA",X"B9",X"17",X"21",X"09",X"00",X"22",
		X"B9",X"40",X"22",X"BB",X"40",X"21",X"02",X"00",X"22",X"BD",X"40",X"3E",X"01",X"32",X"B7",X"40",
		X"AF",X"32",X"C1",X"40",X"32",X"B8",X"40",X"C9",X"3A",X"B8",X"40",X"3D",X"32",X"B8",X"40",X"CB",
		X"4F",X"2A",X"B9",X"40",X"20",X"03",X"2A",X"BB",X"40",X"11",X"01",X"00",X"CD",X"13",X"04",X"3A",
		X"B8",X"40",X"E6",X"03",X"20",X"0B",X"2A",X"B9",X"40",X"EB",X"2A",X"BD",X"40",X"19",X"22",X"B9",
		X"40",X"3A",X"B8",X"40",X"E6",X"0F",X"20",X"2E",X"3A",X"BF",X"40",X"3D",X"32",X"BF",X"40",X"FE",
		X"08",X"CA",X"2D",X"17",X"4F",X"3E",X"01",X"CD",X"95",X"04",X"3A",X"BF",X"40",X"4F",X"3E",X"02",
		X"CD",X"95",X"04",X"3A",X"B8",X"40",X"E6",X"1F",X"20",X"0C",X"2A",X"BD",X"40",X"11",X"08",X"00",
		X"19",X"22",X"BD",X"40",X"18",X"00",X"3E",X"00",X"C9",X"3E",X"FF",X"C9",X"3E",X"00",X"32",X"C9",
		X"40",X"21",X"C7",X"40",X"34",X"7E",X"06",X"05",X"80",X"82",X"81",X"E6",X"07",X"77",X"3E",X"00",
		X"CD",X"78",X"05",X"3E",X"05",X"32",X"C7",X"40",X"11",X"01",X"00",X"21",X"10",X"00",X"CD",X"57",
		X"04",X"0E",X"0D",X"CD",X"DA",X"04",X"3E",X"80",X"32",X"CA",X"40",X"3E",X"40",X"32",X"C8",X"40",
		X"3E",X"00",X"32",X"C4",X"40",X"3E",X"09",X"32",X"C6",X"40",X"3E",X"03",X"32",X"C5",X"40",X"3E",
		X"00",X"32",X"C2",X"40",X"32",X"C3",X"40",X"C9",X"3A",X"C2",X"40",X"2F",X"32",X"C2",X"40",X"B7",
		X"20",X"79",X"3A",X"C3",X"40",X"3D",X"32",X"C3",X"40",X"3A",X"C9",X"40",X"B7",X"20",X"3C",X"3A",
		X"C8",X"40",X"3D",X"32",X"C8",X"40",X"20",X"08",X"3E",X"01",X"32",X"C9",X"40",X"C3",X"D3",X"17",
		X"3A",X"C3",X"40",X"E6",X"1F",X"20",X"0B",X"3A",X"C4",X"40",X"3C",X"32",X"C4",X"40",X"4F",X"CD",
		X"DA",X"04",X"3A",X"CA",X"40",X"06",X"11",X"80",X"E6",X"33",X"06",X"68",X"80",X"32",X"CA",X"40",
		X"6F",X"26",X"00",X"11",X"01",X"00",X"CD",X"57",X"04",X"18",X"30",X"3A",X"C5",X"40",X"06",X"11",
		X"80",X"E6",X"33",X"06",X"64",X"80",X"32",X"C5",X"40",X"21",X"C7",X"40",X"46",X"80",X"6F",X"26",
		X"00",X"11",X"01",X"00",X"CD",X"57",X"04",X"3A",X"C3",X"40",X"E6",X"1F",X"20",X"0D",X"3A",X"C6",
		X"40",X"3D",X"32",X"C6",X"40",X"28",X"07",X"4F",X"CD",X"DA",X"04",X"3E",X"00",X"C9",X"3E",X"FF",
		X"C9",X"3E",X"00",X"CD",X"78",X"05",X"21",X"00",X"00",X"3E",X"01",X"CD",X"B6",X"03",X"0E",X"0F",
		X"3E",X"01",X"CD",X"95",X"04",X"3E",X"11",X"32",X"D1",X"40",X"21",X"90",X"00",X"22",X"CC",X"40",
		X"21",X"F0",X"00",X"22",X"CE",X"40",X"3E",X"00",X"32",X"D0",X"40",X"21",X"F0",X"FF",X"22",X"D3",
		X"40",X"AF",X"32",X"D2",X"40",X"32",X"CB",X"40",X"C9",X"3A",X"CB",X"40",X"3D",X"32",X"CB",X"40",
		X"CB",X"4F",X"2A",X"CC",X"40",X"20",X"03",X"2A",X"CE",X"40",X"3E",X"01",X"CD",X"B6",X"03",X"3A",
		X"CB",X"40",X"E6",X"03",X"20",X"0D",X"2A",X"CC",X"40",X"3A",X"D0",X"40",X"4F",X"06",X"00",X"09",
		X"22",X"CC",X"40",X"3A",X"CB",X"40",X"E6",X"3F",X"20",X"1C",X"3A",X"D1",X"40",X"06",X"FF",X"80",
		X"32",X"D1",X"40",X"FE",X"06",X"28",X"4B",X"FE",X"0F",X"38",X"02",X"3E",X"0F",X"4F",X"3E",X"01",
		X"CD",X"95",X"04",X"3A",X"CB",X"40",X"E6",X"07",X"20",X"35",X"3A",X"D0",X"40",X"06",X"04",X"80",
		X"FE",X"38",X"20",X"02",X"3E",X"00",X"32",X"D0",X"40",X"3A",X"CB",X"40",X"E6",X"04",X"20",X"1F",
		X"2A",X"CE",X"40",X"11",X"FC",X"FF",X"3A",X"D2",X"40",X"B7",X"28",X"03",X"11",X"01",X"00",X"19",
		X"22",X"CE",X"40",X"7D",X"FE",X"40",X"30",X"07",X"3E",X"01",X"32",X"D2",X"40",X"18",X"00",X"3E",
		X"00",X"C9",X"3E",X"FF",X"C9",X"3E",X"00",X"CD",X"78",X"05",X"21",X"00",X"00",X"3E",X"01",X"CD",
		X"B6",X"03",X"21",X"00",X"00",X"3E",X"02",X"CD",X"B6",X"03",X"3E",X"01",X"0E",X"0F",X"CD",X"95",
		X"04",X"3E",X"02",X"0E",X"0F",X"CD",X"95",X"04",X"21",X"00",X"00",X"22",X"D7",X"40",X"21",X"0A",
		X"00",X"22",X"D9",X"40",X"3E",X"10",X"32",X"D6",X"40",X"AF",X"32",X"DB",X"40",X"32",X"DC",X"40",
		X"32",X"DD",X"40",X"32",X"D5",X"40",X"C9",X"3E",X"01",X"32",X"11",X"40",X"3A",X"D5",X"40",X"3D",
		X"32",X"D5",X"40",X"CB",X"47",X"28",X"1E",X"3A",X"DB",X"40",X"3C",X"FE",X"66",X"20",X"02",X"3E",
		X"00",X"32",X"DB",X"40",X"4F",X"06",X"00",X"2A",X"D7",X"40",X"09",X"22",X"D7",X"40",X"3E",X"01",
		X"CD",X"B6",X"03",X"18",X"1E",X"3A",X"DC",X"40",X"3C",X"FE",X"11",X"20",X"02",X"3E",X"00",X"32",
		X"DC",X"40",X"4F",X"06",X"00",X"2A",X"D9",X"40",X"09",X"22",X"D9",X"40",X"3E",X"02",X"CD",X"B6",
		X"03",X"18",X"00",X"3A",X"DD",X"40",X"3C",X"32",X"DD",X"40",X"FE",X"FF",X"20",X"27",X"3E",X"00",
		X"32",X"DD",X"40",X"3A",X"D6",X"40",X"3D",X"32",X"D6",X"40",X"FE",X"0F",X"38",X"02",X"3E",X"0F",
		X"FE",X"05",X"28",X"14",X"4F",X"3E",X"01",X"CD",X"95",X"04",X"3A",X"D6",X"40",X"4F",X"3E",X"02",
		X"CD",X"95",X"04",X"18",X"00",X"3E",X"00",X"C9",X"3E",X"FF",X"C9",X"2A",X"E9",X"40",X"7C",X"B5",
		X"28",X"06",X"2B",X"22",X"E9",X"40",X"18",X"59",X"3E",X"00",X"CD",X"78",X"05",X"21",X"80",X"02",
		X"32",X"E9",X"40",X"21",X"01",X"00",X"11",X"00",X"00",X"CD",X"13",X"04",X"0E",X"00",X"3E",X"03",
		X"CD",X"95",X"04",X"0E",X"0F",X"3E",X"01",X"CD",X"95",X"04",X"3E",X"02",X"0E",X"0F",X"CD",X"95",
		X"04",X"3E",X"10",X"32",X"E7",X"40",X"3A",X"E7",X"40",X"3D",X"32",X"E7",X"40",X"32",X"E6",X"40",
		X"FE",X"08",X"CA",X"E5",X"1A",X"21",X"09",X"00",X"22",X"E0",X"40",X"22",X"E2",X"40",X"21",X"02",
		X"00",X"22",X"E4",X"40",X"3E",X"01",X"32",X"DE",X"40",X"AF",X"32",X"E8",X"40",X"32",X"DF",X"40",
		X"C9",X"3E",X"01",X"C9",X"3A",X"DF",X"40",X"3D",X"32",X"DF",X"40",X"CB",X"4F",X"2A",X"E0",X"40",
		X"20",X"03",X"2A",X"E2",X"40",X"11",X"01",X"00",X"CD",X"13",X"04",X"3A",X"DF",X"40",X"E6",X"03",
		X"20",X"0B",X"2A",X"E0",X"40",X"EB",X"2A",X"E4",X"40",X"19",X"22",X"E0",X"40",X"3A",X"DF",X"40",
		X"E6",X"0F",X"20",X"2E",X"3A",X"E6",X"40",X"3D",X"32",X"E6",X"40",X"FE",X"08",X"CA",X"56",X"1A",
		X"4F",X"3E",X"01",X"CD",X"95",X"04",X"3A",X"E6",X"40",X"4F",X"3E",X"02",X"CD",X"95",X"04",X"3A",
		X"DF",X"40",X"E6",X"1F",X"20",X"0C",X"2A",X"E4",X"40",X"11",X"08",X"00",X"19",X"22",X"E4",X"40",
		X"18",X"00",X"3E",X"00",X"C9",X"21",X"80",X"02",X"22",X"E9",X"40",X"3E",X"FF",X"C9",X"3E",X"03",
		X"32",X"F1",X"40",X"3A",X"F1",X"40",X"3D",X"32",X"F1",X"40",X"28",X"73",X"3E",X"00",X"CD",X"78",
		X"05",X"11",X"FE",X"FF",X"21",X"28",X"00",X"CD",X"D5",X"03",X"0E",X"06",X"CD",X"DA",X"04",X"3E",
		X"0E",X"32",X"EE",X"40",X"21",X"28",X"00",X"22",X"EF",X"40",X"3E",X"0E",X"32",X"ED",X"40",X"AF",
		X"32",X"EB",X"40",X"32",X"EC",X"40",X"C9",X"3A",X"EB",X"40",X"2F",X"32",X"EB",X"40",X"B7",X"20",
		X"3C",X"3A",X"EC",X"40",X"3D",X"32",X"EC",X"40",X"47",X"E6",X"3F",X"20",X"0B",X"3A",X"EE",X"40",
		X"3D",X"32",X"EE",X"40",X"FE",X"0A",X"28",X"AB",X"78",X"E6",X"1F",X"20",X"16",X"2A",X"EF",X"40",
		X"01",X"FF",X"FF",X"09",X"22",X"EF",X"40",X"11",X"FE",X"FF",X"CD",X"D5",X"03",X"3A",X"EE",X"40",
		X"32",X"ED",X"40",X"21",X"ED",X"40",X"35",X"4E",X"CD",X"DA",X"04",X"18",X"00",X"AF",X"C9",X"3E",
		X"FF",X"C9",X"3E",X"00",X"CD",X"78",X"05",X"3E",X"01",X"21",X"01",X"01",X"CD",X"B6",X"03",X"0E",
		X"0F",X"3E",X"01",X"CD",X"95",X"04",X"3E",X"08",X"32",X"F3",X"40",X"21",X"80",X"00",X"22",X"F5",
		X"40",X"3E",X"08",X"32",X"F4",X"40",X"AF",X"32",X"FD",X"40",X"32",X"F2",X"40",X"C9",X"3A",X"F3",
		X"40",X"3D",X"32",X"F3",X"40",X"20",X"3D",X"3A",X"F4",X"40",X"32",X"F3",X"40",X"3A",X"F2",X"40",
		X"3D",X"32",X"F2",X"40",X"0E",X"0F",X"CB",X"47",X"20",X"02",X"0E",X"00",X"3E",X"01",X"CD",X"95",
		X"04",X"2A",X"F5",X"40",X"AF",X"11",X"01",X"00",X"ED",X"52",X"22",X"F5",X"40",X"20",X"15",X"21",
		X"00",X"01",X"22",X"F5",X"40",X"3A",X"F4",X"40",X"06",X"FE",X"80",X"FE",X"04",X"28",X"08",X"32",
		X"F4",X"40",X"18",X"00",X"3E",X"00",X"C9",X"3E",X"FF",X"32",X"FD",X"40",X"3E",X"FF",X"C9",X"BD",
		X"B1",X"B0",X"A7",X"AE",X"B7",X"B9",X"B8",X"AC",X"E0",X"9E",X"87",X"E0",X"B5",X"B1",X"B2",X"BF",
		X"B3",X"B7",X"E0",X"CF",X"C7",X"C8",X"CC",X"3E",X"00",X"CD",X"78",X"05",X"3E",X"01",X"21",X"01",
		X"01",X"CD",X"B6",X"03",X"0E",X"0F",X"3E",X"01",X"CD",X"95",X"04",X"3E",X"02",X"32",X"F8",X"40",
		X"21",X"20",X"00",X"22",X"FA",X"40",X"3E",X"08",X"32",X"F9",X"40",X"AF",X"32",X"FD",X"40",X"32",
		X"FC",X"40",X"32",X"F7",X"40",X"C9",X"3A",X"F8",X"40",X"3D",X"32",X"F8",X"40",X"20",X"4F",X"3A",
		X"F9",X"40",X"32",X"F8",X"40",X"3A",X"F7",X"40",X"3D",X"32",X"F7",X"40",X"0E",X"0F",X"CB",X"47",
		X"20",X"02",X"0E",X"00",X"3E",X"01",X"CD",X"95",X"04",X"2A",X"FA",X"40",X"AF",X"11",X"01",X"00",
		X"ED",X"52",X"22",X"FA",X"40",X"20",X"27",X"21",X"70",X"00",X"22",X"FA",X"40",X"3A",X"FC",X"40",
		X"3C",X"32",X"FC",X"40",X"4F",X"06",X"00",X"21",X"85",X"1C",X"09",X"7E",X"FE",X"FF",X"28",X"11",
		X"32",X"F9",X"40",X"18",X"09",X"08",X"06",X"06",X"08",X"06",X"04",X"04",X"04",X"FF",X"3E",X"00",
		X"C9",X"3E",X"FF",X"32",X"FD",X"40",X"C9",X"3E",X"00",X"CD",X"78",X"05",X"3E",X"01",X"21",X"81",
		X"00",X"CD",X"B6",X"03",X"0E",X"0B",X"3E",X"01",X"CD",X"95",X"04",X"3E",X"01",X"32",X"FF",X"40",
		X"AF",X"32",X"FE",X"40",X"C9",X"3A",X"FD",X"40",X"B7",X"20",X"27",X"3A",X"FF",X"40",X"3D",X"32",
		X"FF",X"40",X"20",X"1B",X"3E",X"01",X"32",X"FF",X"40",X"3A",X"FE",X"40",X"3D",X"32",X"FE",X"40",
		X"0E",X"0B",X"CB",X"47",X"20",X"02",X"0E",X"00",X"3E",X"01",X"CD",X"95",X"04",X"18",X"00",X"3E",
		X"00",X"C9",X"3E",X"00",X"32",X"FD",X"40",X"3E",X"FF",X"C9",X"3E",X"00",X"CD",X"78",X"05",X"21",
		X"0E",X"00",X"11",X"01",X"00",X"CD",X"D5",X"03",X"0E",X"0A",X"CD",X"DA",X"04",X"21",X"0D",X"00",
		X"22",X"02",X"41",X"22",X"04",X"41",X"3E",X"0A",X"32",X"06",X"41",X"32",X"07",X"41",X"3E",X"00",
		X"32",X"00",X"41",X"32",X"01",X"41",X"C9",X"3A",X"00",X"41",X"2F",X"32",X"00",X"41",X"B7",X"20",
		X"47",X"3A",X"01",X"41",X"3D",X"32",X"01",X"41",X"E6",X"0F",X"20",X"24",X"2A",X"04",X"41",X"2B",
		X"22",X"04",X"41",X"11",X"01",X"00",X"CD",X"D5",X"03",X"3A",X"07",X"41",X"D6",X"01",X"47",X"3A",
		X"06",X"41",X"3D",X"B8",X"30",X"03",X"3A",X"07",X"41",X"32",X"06",X"41",X"4F",X"CD",X"DA",X"04",
		X"3A",X"01",X"41",X"E6",X"3F",X"20",X"11",X"2A",X"02",X"41",X"7D",X"FE",X"06",X"28",X"0C",X"2B",
		X"22",X"02",X"41",X"22",X"04",X"41",X"18",X"00",X"3E",X"00",X"C9",X"3E",X"FF",X"C9",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
