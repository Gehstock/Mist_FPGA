library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity obj_7s is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of obj_7s is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"78",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"F0",X"E0",X"00",X"00",X"0C",X"0C",X"0C",X"00",X"00",X"00",X"E0",X"F0",X"F8",X"FC",
		X"00",X"00",X"00",X"1C",X"1C",X"1C",X"04",X"00",X"00",X"03",X"03",X"03",X"E0",X"F0",X"F8",X"FC",
		X"00",X"00",X"10",X"38",X"1C",X"14",X"00",X"00",X"04",X"0E",X"0E",X"04",X"E0",X"F0",X"F8",X"FC",
		X"1E",X"1C",X"00",X"00",X"00",X"02",X"07",X"03",X"00",X"00",X"00",X"00",X"E0",X"F0",X"F8",X"FC",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"E0",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"03",X"00",X"F0",X"F8",X"FC",X"FE",X"9C",
		X"3C",X"38",X"00",X"00",X"18",X"18",X"1C",X"10",X"00",X"00",X"00",X"F0",X"F8",X"FC",X"FE",X"BC",
		X"00",X"00",X"0F",X"00",X"00",X"03",X"03",X"00",X"00",X"70",X"FC",X"FE",X"FC",X"00",X"00",X"00",
		X"E0",X"00",X"00",X"20",X"70",X"78",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"06",X"02",X"02",X"00",X"00",X"80",X"C0",X"E0",X"F0",
		X"10",X"38",X"70",X"60",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"07",X"07",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"1C",X"0E",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"0E",X"1E",X"8C",X"C0",X"E0",X"F0",
		X"08",X"1C",X"0E",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"0E",X"1E",X"8C",X"C0",X"E0",X"F0",
		X"08",X"1C",X"0E",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"0E",X"1E",X"8C",X"C0",X"E0",X"F0",
		X"1E",X"00",X"00",X"00",X"00",X"03",X"03",X"00",X"00",X"F0",X"F8",X"FC",X"38",X"20",X"00",X"00",
		X"1E",X"00",X"00",X"03",X"07",X"00",X"00",X"70",X"FC",X"FE",X"3C",X"00",X"00",X"00",X"00",X"00",
		X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"0E",X"07",X"07",X"03",X"00",X"C0",X"E0",X"F0",X"F0",X"F0",X"F0",X"FB",X"DB",X"9A",X"E0",
		X"0C",X"0E",X"07",X"07",X"03",X"01",X"C3",X"E3",X"F0",X"F0",X"F0",X"F0",X"F8",X"D8",X"98",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"10",X"10",X"EE",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"10",X"10",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"10",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"03",X"03",X"03",X"F0",X"88",X"BC",
		X"FE",X"9C",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"06",X"03",X"03",X"01",X"00",X"0E",X"0E",X"06",X"00",X"00",X"E0",X"F0",X"F8",X"FC",
		X"00",X"04",X"06",X"03",X"03",X"01",X"00",X"07",X"03",X"00",X"00",X"F0",X"F8",X"FC",X"FE",X"9C",
		X"00",X"00",X"FC",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"FC",
		X"50",X"90",X"60",X"A0",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EC",X"FE",X"6A",X"40",X"80",X"80",X"44",X"40",X"20",X"20",X"A2",X"40",X"40",X"68",X"68",X"50",
		X"70",X"30",X"20",X"60",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7A",X"FF",X"D2",X"80",X"C9",X"40",X"40",X"90",X"D0",X"D8",X"68",X"28",X"28",X"10",X"10",X"90",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"BE",X"BE",X"3E",X"3E",X"1E",
		X"7E",X"7E",X"7E",X"7E",X"7E",X"FE",X"FE",X"FE",X"FE",X"7E",X"7E",X"FA",X"F2",X"F0",X"F0",X"F0",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"F0",X"FC",X"FE",X"FE",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"FA",X"F2",X"F0",X"F0",X"F0",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"F8",X"FC",X"FE",X"FE",X"7E",X"F0",X"FC",X"FE",X"FE",X"7E",X"7E",X"FA",X"F2",X"F0",X"F0",X"F0",
		X"1E",X"1E",X"1E",X"1E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"52",X"F7",X"F7",X"F7",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FE",X"FE",X"FE",X"FE",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FE",X"FE",X"FE",X"FE",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F7",X"F7",X"F7",X"F7",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F4",X"E2",X"F0",X"48",X"20",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"06",X"03",X"03",X"40",X"80",X"C0",X"D0",X"F0",X"F8",X"F8",X"FC",X"FF",X"77",X"F4",X"F8",
		X"04",X"06",X"03",X"03",X"40",X"81",X"C3",X"D7",X"FE",X"FE",X"FC",X"F8",X"F0",X"70",X"F0",X"F8",
		X"FE",X"FC",X"D0",X"E0",X"F0",X"E8",X"40",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"62",X"77",X"F7",X"EF",X"F0",X"FA",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"FF",X"FF",X"00",
		X"36",X"36",X"36",X"36",X"36",X"36",X"76",X"66",X"EE",X"CC",X"9C",X"38",X"F8",X"E0",X"80",X"00",
		X"36",X"36",X"36",X"36",X"36",X"36",X"36",X"36",X"36",X"36",X"36",X"36",X"36",X"36",X"36",X"36",
		X"00",X"00",X"00",X"00",X"20",X"30",X"38",X"7C",X"DE",X"BE",X"1A",X"50",X"70",X"70",X"50",X"30",
		X"00",X"00",X"00",X"00",X"2C",X"3E",X"3F",X"7F",X"CD",X"A8",X"38",X"A8",X"D8",X"D8",X"C0",X"00",
		X"F0",X"E0",X"C0",X"F0",X"7C",X"70",X"70",X"33",X"3F",X"7F",X"65",X"46",X"46",X"04",X"00",X"00",
		X"E0",X"E0",X"DC",X"F8",X"F0",X"78",X"7C",X"7B",X"37",X"7F",X"65",X"46",X"46",X"04",X"00",X"00",
		X"F0",X"E0",X"C0",X"F0",X"78",X"7C",X"7B",X"37",X"7F",X"65",X"46",X"46",X"04",X"00",X"00",X"00",
		X"C0",X"F8",X"F0",X"C0",X"F0",X"78",X"7C",X"7B",X"37",X"7F",X"65",X"46",X"46",X"04",X"00",X"00",
		X"F8",X"F0",X"C0",X"F0",X"78",X"7C",X"7B",X"37",X"7F",X"65",X"46",X"46",X"04",X"00",X"00",X"00",
		X"00",X"00",X"E0",X"C0",X"00",X"E0",X"E0",X"30",X"00",X"CC",X"9C",X"FC",X"F4",X"0C",X"08",X"80",
		X"C0",X"80",X"00",X"00",X"00",X"E0",X"E0",X"30",X"00",X"CC",X"9C",X"FC",X"F4",X"0C",X"08",X"80",
		X"F0",X"E0",X"00",X"00",X"F0",X"F0",X"18",X"80",X"E6",X"CE",X"FE",X"FA",X"86",X"84",X"40",X"00",
		X"78",X"70",X"E0",X"00",X"00",X"0E",X"7C",X"78",X"80",X"CC",X"9C",X"F4",X"8C",X"8C",X"88",X"C0",
		X"C0",X"80",X"00",X"08",X"0E",X"0E",X"06",X"82",X"00",X"00",X"D8",X"38",X"F8",X"18",X"10",X"00",
		X"2E",X"1E",X"0C",X"08",X"08",X"08",X"0B",X"1F",X"3E",X"FC",X"E0",X"C0",X"80",X"00",X"00",X"00",
		X"20",X"10",X"08",X"08",X"08",X"08",X"08",X"18",X"30",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"20",X"20",X"20",X"60",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"30",X"28",X"28",X"68",X"F8",X"F0",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"20",X"38",X"30",X"70",X"D0",X"9A",X"3E",X"9E",X"0C",X"00",X"00",X"00",
		X"20",X"10",X"08",X"08",X"00",X"00",X"00",X"00",X"1C",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"60",X"10",X"00",X"00",X"00",X"04",X"04",X"08",X"10",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"C0",X"20",X"00",X"04",X"04",X"04",X"08",X"08",X"10",X"20",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"10",X"08",X"08",X"08",X"08",X"08",X"18",X"30",X"E0",
		X"00",X"00",X"00",X"20",X"20",X"10",X"08",X"08",X"08",X"08",X"08",X"18",X"30",X"E0",X"00",X"00",
		X"00",X"20",X"20",X"10",X"08",X"08",X"08",X"08",X"08",X"18",X"30",X"E0",X"00",X"00",X"00",X"00",
		X"FC",X"FE",X"FE",X"FE",X"DE",X"1C",X"3C",X"38",X"38",X"38",X"90",X"D0",X"A0",X"80",X"80",X"00",
		X"7C",X"7E",X"F6",X"E6",X"CE",X"1C",X"2C",X"B8",X"38",X"38",X"10",X"80",X"80",X"80",X"80",X"00",
		X"7C",X"F0",X"E4",X"C8",X"88",X"10",X"28",X"30",X"38",X"08",X"80",X"E0",X"A0",X"80",X"80",X"00",
		X"18",X"14",X"08",X"00",X"00",X"00",X"08",X"04",X"04",X"00",X"00",X"88",X"10",X"00",X"00",X"00",
		X"06",X"03",X"00",X"00",X"00",X"10",X"02",X"01",X"01",X"10",X"20",X"00",X"86",X"80",X"80",X"00",
		X"04",X"0C",X"80",X"02",X"00",X"00",X"60",X"02",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"F0",X"E8",X"DC",X"BE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"0F",X"0F",X"0F",X"0E",X"8C",X"C8",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"F8",X"FE",X"FC",X"F0",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"0E",X"F8",X"E1",X"07",X"1E",X"F8",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"FC",X"00",X"06",X"F6",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"1E",X"F8",X"E1",X"07",X"1E",X"F8",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"0E",X"E1",X"E1",X"10",X"10",X"0E",X"0E",X"E0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"0E",X"0E",X"10",X"10",X"E0",X"E0",X"0E",X"0E",
		X"00",X"00",X"00",X"0E",X"EE",X"E1",X"11",X"10",X"00",X"0E",X"EE",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FE",X"BA",X"BB",X"77",X"FF",X"FF",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"FF",X"FF",X"BB",X"BB",X"B7",X"FF",X"DD",X"EF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"FF",X"FF",X"BB",X"BB",X"B7",X"FF",X"DD",X"EF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E8",X"B0",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"06",X"0C",X"18",X"30",X"EE",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"81",X"C3",X"C3",X"C3",X"FF",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"1D",X"3F",X"3E",X"3C",X"F8",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"83",X"C3",X"CF",X"FC",X"F0",X"C0",X"00",X"00",
		X"00",X"E0",X"70",X"C8",X"80",X"80",X"80",X"44",X"A0",X"B0",X"D0",X"D2",X"A0",X"40",X"80",X"00",
		X"00",X"60",X"90",X"68",X"F4",X"94",X"94",X"94",X"B4",X"6C",X"C8",X"18",X"30",X"E0",X"00",X"00",
		X"00",X"E0",X"10",X"C8",X"68",X"34",X"14",X"D4",X"74",X"94",X"C4",X"48",X"50",X"60",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"40",X"40",X"40",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"70",X"90",X"68",X"A8",X"A8",X"C8",X"30",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"C0",X"20",X"D0",X"50",X"D0",X"50",X"A0",X"60",X"20",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"90",X"50",X"20",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"40",X"A0",X"A0",X"60",X"20",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"20",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"08",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"08",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"E0",X"60",X"B0",X"B0",X"B0",X"B0",X"B0",X"F0",X"E0",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"20",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"3C",X"E0",X"0A",X"E0",X"FE",X"7E",X"FC",X"F8",X"F0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"2A",X"2A",X"12",X"C4",X"FC",X"C0",X"9C",X"C6",X"8E",X"16",X"8C",X"98",X"00",X"00",X"00",X"00",
		X"20",X"29",X"12",X"C2",X"FC",X"C0",X"98",X"C4",X"8E",X"0E",X"8A",X"82",X"04",X"00",X"00",X"00",
		X"94",X"54",X"54",X"14",X"C4",X"F8",X"C0",X"9C",X"CE",X"8B",X"09",X"85",X"80",X"00",X"00",X"00",
		X"29",X"29",X"92",X"86",X"BC",X"E0",X"D8",X"8C",X"C6",X"8F",X"1F",X"3B",X"23",X"87",X"5F",X"3C",
		X"52",X"52",X"84",X"98",X"A0",X"EE",X"D7",X"8F",X"CB",X"8B",X"03",X"07",X"06",X"80",X"40",X"20",
		X"48",X"24",X"84",X"84",X"B8",X"E0",X"DC",X"86",X"CF",X"9F",X"1B",X"17",X"07",X"8E",X"4C",X"20",
		X"0C",X"A6",X"0B",X"0B",X"CF",X"E7",X"DA",X"CC",X"C0",X"9C",X"24",X"12",X"09",X"00",X"00",X"00",
		X"0C",X"A6",X"0B",X"0B",X"CF",X"E7",X"DA",X"CC",X"C0",X"90",X"28",X"28",X"48",X"08",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"C0",X"9C",X"BE",X"60",X"60",X"60",X"70",X"71",X"7F",X"1F",X"1F",X"16",X"1E",X"1C",X"18",
		X"0E",X"FC",X"F8",X"FC",X"F8",X"F8",X"F0",X"F8",X"F8",X"F8",X"78",X"30",X"30",X"20",X"40",X"00",
		X"1E",X"F8",X"FE",X"F0",X"70",X"B0",X"E0",X"C8",X"D0",X"D0",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"3B",X"FE",X"FE",X"E2",X"41",X"C0",X"C0",X"80",X"00",X"04",X"18",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"10",X"10",X"10",X"1F",X"F0",X"1F",X"DF",X"DF",X"DF",X"DF",X"FF",X"FF",X"DF",X"DF",X"FF",
		X"A0",X"A0",X"A0",X"D0",X"E8",X"F7",X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"00",
		X"D0",X"D0",X"D0",X"FF",X"20",X"00",X"20",X"20",X"20",X"20",X"80",X"20",X"20",X"20",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"A0",X"A0",X"A0",X"A0",X"A0",X"20",X"FE",
		X"A0",X"A0",X"A0",X"D0",X"E8",X"F4",X"FB",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"00",
		X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"20",X"FE",X"D0",X"D0",X"D0",X"FF",
		X"FE",X"D3",X"D3",X"D3",X"FF",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",
		X"00",X"7F",X"FF",X"80",X"00",X"7F",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"F3",X"E1",X"E0",X"00",
		X"F0",X"10",X"10",X"10",X"1F",X"F0",X"1F",X"DF",X"DF",X"DF",X"DF",X"FF",X"FF",X"DF",X"DF",X"FF",
		X"70",X"10",X"10",X"10",X"9F",X"70",X"9F",X"DF",X"DF",X"DF",X"DF",X"FF",X"FF",X"DF",X"DF",X"FF",
		X"10",X"10",X"10",X"1F",X"F0",X"1F",X"5F",X"DF",X"DF",X"DF",X"DF",X"DF",X"FF",X"FF",X"DF",X"DF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"10",X"24",X"88",X"98",X"A4",X"EC",X"ED",X"D9",X"FB",X"BB",X"3F",X"9F",X"1F",X"8E",X"4C",X"20",
		X"40",X"20",X"A0",X"E0",X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",
		X"50",X"48",X"08",X"F0",X"F0",X"E0",X"FC",X"E6",X"E3",X"47",X"6D",X"6B",X"6B",X"67",X"6E",X"00",
		X"40",X"20",X"A0",X"E0",X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",
		X"00",X"80",X"D0",X"F0",X"00",X"40",X"40",X"00",X"60",X"E0",X"A0",X"F0",X"58",X"E0",X"F8",X"70",
		X"00",X"80",X"D0",X"F0",X"00",X"40",X"40",X"00",X"70",X"FC",X"BE",X"DE",X"0E",X"04",X"00",X"00",
		X"00",X"A0",X"D0",X"E0",X"00",X"48",X"42",X"06",X"7E",X"FC",X"A0",X"C0",X"00",X"00",X"00",X"00",
		X"C0",X"E8",X"1A",X"26",X"CC",X"88",X"60",X"F0",X"A0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C3",X"AF",X"FE",X"70",X"00",X"40",X"40",X"00",X"F0",X"D0",X"A0",X"00",X"00",X"00",X"00",X"00",
		X"C3",X"AF",X"FE",X"70",X"00",X"40",X"40",X"00",X"F0",X"C8",X"80",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"FE",X"FE",X"FE",X"AE",X"5C",X"FC",X"B8",X"B8",X"B8",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"FE",X"FE",X"AE",X"5E",X"FC",X"00",X"A0",X"A0",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"FE",X"FE",X"00",X"00",X"00",X"00",X"A0",X"A0",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"F8",X"04",X"00",X"00",X"00",X"00",X"A0",X"A0",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"F8",X"04",X"00",X"00",X"00",X"00",X"A0",X"A0",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"FE",X"FE",X"FE",X"AE",X"5C",X"FC",X"B8",X"B8",X"B8",X"B0",X"D0",X"80",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"C0",X"A0",X"80",X"C0",X"E0",X"A0",X"A0",X"C0",X"80",X"00",X"00",
		X"00",X"F8",X"FC",X"06",X"06",X"00",X"FC",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FE",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"FE",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"10",X"18",X"1C",X"1C",X"1E",X"1E",X"1E",X"1E",X"1E",X"1E",X"1C",X"1C",X"18",X"10",X"00",
		X"00",X"30",X"38",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"38",X"30",X"00",
		X"40",X"70",X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"70",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",
		X"00",X"00",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"80",X"80",
		X"00",X"00",X"C0",X"E0",X"60",X"B0",X"B0",X"B0",X"B0",X"B0",X"F0",X"E0",X"C0",X"80",X"80",X"80",
		X"00",X"00",X"00",X"20",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"20",X"00",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",
		X"00",X"00",X"E0",X"10",X"68",X"A8",X"A8",X"A8",X"A8",X"A8",X"E8",X"10",X"E0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"40",X"20",X"00",X"20",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"60",X"10",X"48",X"28",X"00",X"28",X"48",X"10",X"60",X"00",X"00",X"00",X"00",
		X"00",X"00",X"70",X"08",X"64",X"34",X"14",X"00",X"14",X"34",X"64",X"08",X"70",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"60",X"D0",X"70",X"20",X"70",X"D0",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"60",X"20",X"60",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"20",X"C8",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"80",X"A0",X"A0",X"A0",X"20",X"10",X"00",
		X"00",X"00",X"00",X"80",X"00",X"00",X"10",X"10",X"90",X"A0",X"A0",X"C0",X"C0",X"A0",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"20",X"20",X"20",X"20",X"28",X"28",X"20",X"20",X"24",
		X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"20",X"20",X"20",X"20",X"28",X"28",X"20",X"20",X"24",
		X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"20",X"30",X"30",X"20",X"28",X"28",X"20",X"20",X"24",
		X"00",X"00",X"00",X"00",X"2C",X"3E",X"3F",X"7F",X"CF",X"AF",X"3B",X"AB",X"DF",X"DA",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"F0",X"F0",X"78",X"F8",X"F8",X"98",X"F0",
		X"20",X"70",X"70",X"39",X"22",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"84",X"8E",X"CE",X"CC",X"FC",X"0E",X"03",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"A0",X"E0",X"E0",X"C0",X"10",X"F8",X"78",X"24",X"1E",X"0E",X"0C",X"04",X"04",X"00",X"0C",
		X"18",X"3C",X"7A",X"FB",X"7F",X"7F",X"4D",X"5E",X"8C",X"C0",X"E0",X"F0",X"60",X"00",X"00",X"00",
		X"06",X"56",X"03",X"0F",X"C7",X"E3",X"EA",X"E6",X"F0",X"EE",X"12",X"09",X"04",X"00",X"00",X"00",
		X"00",X"40",X"20",X"20",X"08",X"84",X"C4",X"E0",X"E2",X"F3",X"E1",X"E5",X"57",X"5F",X"8E",X"00",
		X"04",X"8E",X"5F",X"57",X"15",X"C5",X"E3",X"E2",X"E0",X"E4",X"E4",X"88",X"00",X"20",X"40",X"00",
		X"00",X"00",X"00",X"10",X"92",X"A4",X"18",X"C0",X"CE",X"F3",X"E7",X"CF",X"0B",X"0B",X"A6",X"0C",
		X"80",X"00",X"00",X"C0",X"00",X"10",X"94",X"C4",X"D8",X"C0",X"F8",X"CC",X"1C",X"2C",X"1C",X"78",
		X"38",X"3C",X"66",X"1E",X"04",X"98",X"C0",X"D8",X"E4",X"D4",X"90",X"00",X"C0",X"00",X"00",X"80",
		X"C0",X"A0",X"E0",X"70",X"06",X"4F",X"4F",X"06",X"F0",X"D0",X"A0",X"00",X"00",X"00",X"00",X"00",
		X"18",X"BC",X"2C",X"18",X"46",X"8F",X"2B",X"46",X"10",X"A4",X"CC",X"D4",X"F4",X"AC",X"18",X"00",
		X"00",X"0C",X"9E",X"58",X"D2",X"CC",X"A4",X"10",X"46",X"2B",X"8F",X"46",X"18",X"2C",X"3C",X"18",
		X"00",X"00",X"00",X"00",X"00",X"D0",X"E8",X"F8",X"01",X"A5",X"A3",X"8E",X"3C",X"70",X"50",X"60",
		X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"E0",X"68",X"18",X"00",X"70",X"B8",X"98",X"50",
		X"30",X"F8",X"98",X"68",X"00",X"10",X"68",X"E0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0E",X"D3",X"D3",X"D3",X"D3",X"CE",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"1B",X"9B",X"9B",X"9F",X"8F",X"87",X"8F",X"9B",X"13",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FE",X"FE",X"00",X"83",X"C3",X"CF",X"D3",X"D3",X"D3",X"D3",X"8F",X"00",X"FE",X"FE",X"00",
		X"00",X"00",X"00",X"00",X"FE",X"FE",X"00",X"83",X"CF",X"D3",X"D3",X"8F",X"00",X"FE",X"FE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FE",X"CF",X"D3",X"DF",X"FE",X"FE",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
