library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity prog is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of prog is
	type rom is array(0 to  32767) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"F3",X"31",X"00",X"E8",X"01",X"00",X"00",X"FD",X"21",X"00",X"00",X"10",X"FA",X"0D",X"20",X"F7",
		X"ED",X"56",X"21",X"B3",X"E6",X"36",X"01",X"DB",X"04",X"CB",X"7F",X"CA",X"41",X"6F",X"35",X"CD",
		X"7A",X"00",X"00",X"00",X"00",X"FB",X"C3",X"CF",X"25",X"CD",X"00",X"1D",X"CD",X"4C",X"04",X"CD",
		X"2C",X"07",X"18",X"F5",X"C7",X"C7",X"C7",X"C7",X"08",X"D9",X"DD",X"E5",X"FD",X"E5",X"CD",X"28",
		X"01",X"CD",X"A2",X"00",X"CD",X"68",X"31",X"3A",X"6A",X"E5",X"B7",X"C4",X"4B",X"2A",X"3A",X"9D",
		X"E5",X"FE",X"02",X"CC",X"41",X"01",X"CD",X"90",X"01",X"FD",X"E1",X"DD",X"E1",X"D9",X"08",X"FB",
		X"C9",X"C7",X"C7",X"C7",X"C7",X"C7",X"FB",X"ED",X"45",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"93",X"24",X"6C",X"DB",X"7A",X"FB",X"85",X"91",X"A3",X"80",X"AF",X"32",X"9D",X"E5",X"D3",X"01",
		X"21",X"00",X"D0",X"36",X"00",X"54",X"5D",X"13",X"01",X"F0",X"17",X"ED",X"B0",X"CD",X"28",X"01",
		X"CD",X"F4",X"08",X"CD",X"D6",X"08",X"CD",X"A6",X"6D",X"3E",X"00",X"D3",X"00",X"F6",X"80",X"D3",
		X"00",X"C9",X"21",X"B5",X"E5",X"35",X"23",X"35",X"21",X"B5",X"E6",X"35",X"3A",X"B9",X"E5",X"B7",
		X"20",X"04",X"DB",X"01",X"18",X"02",X"DB",X"02",X"2F",X"32",X"4D",X"E4",X"21",X"CF",X"E5",X"07",
		X"CB",X"16",X"07",X"07",X"CB",X"16",X"3A",X"4D",X"E4",X"21",X"D0",X"E5",X"0F",X"CB",X"16",X"0F",
		X"CB",X"16",X"DB",X"00",X"2F",X"21",X"AA",X"E5",X"1F",X"CB",X"16",X"1F",X"CB",X"16",X"DB",X"04",
		X"CB",X"67",X"20",X"29",X"21",X"B4",X"E5",X"7E",X"B7",X"20",X"11",X"3A",X"AA",X"E5",X"E6",X"05",
		X"FE",X"05",X"20",X"06",X"36",X"01",X"F1",X"C3",X"59",X"00",X"18",X"11",X"3A",X"AA",X"E5",X"E6",
		X"0A",X"FE",X"0A",X"20",X"04",X"36",X"00",X"18",X"04",X"F1",X"C3",X"59",X"00",X"CD",X"23",X"09",
		X"3A",X"AF",X"E5",X"B7",X"20",X"05",X"3E",X"02",X"32",X"B2",X"E5",X"3A",X"A7",X"E5",X"B7",X"C8",
		X"3A",X"B2",X"E5",X"B7",X"C8",X"C3",X"A0",X"68",X"3A",X"B3",X"E6",X"B7",X"28",X"07",X"CD",X"39",
		X"7C",X"F1",X"C3",X"59",X"00",X"01",X"00",X"01",X"11",X"00",X"C0",X"21",X"00",X"E3",X"ED",X"B0",
		X"C9",X"CD",X"E6",X"03",X"CD",X"00",X"0B",X"CD",X"00",X"13",X"CD",X"00",X"24",X"C9",X"FD",X"E5",
		X"3A",X"E9",X"E4",X"32",X"88",X"E5",X"FD",X"21",X"58",X"E4",X"11",X"18",X"00",X"DD",X"7E",X"06",
		X"FD",X"BE",X"06",X"20",X"20",X"DD",X"7E",X"07",X"FD",X"96",X"07",X"30",X"02",X"ED",X"44",X"FE",
		X"04",X"30",X"12",X"FD",X"7E",X"0D",X"B7",X"28",X"0C",X"FD",X"7E",X"08",X"FE",X"09",X"30",X"02",
		X"0E",X"FF",X"FD",X"E1",X"C9",X"FD",X"19",X"21",X"88",X"E5",X"35",X"20",X"D0",X"FD",X"E1",X"C9",
		X"3A",X"9D",X"E5",X"B7",X"C8",X"3A",X"6A",X"E5",X"B7",X"CC",X"03",X"32",X"DD",X"21",X"40",X"E4",
		X"FD",X"21",X"B0",X"E3",X"3A",X"6A",X"E5",X"FE",X"02",X"20",X"04",X"FD",X"21",X"F0",X"E3",X"AF",
		X"32",X"E8",X"E4",X"DD",X"4E",X"0A",X"3A",X"E8",X"E4",X"B7",X"28",X"17",X"DD",X"7E",X"0D",X"B7",
		X"28",X"0E",X"DD",X"34",X"08",X"DD",X"7E",X"08",X"FE",X"18",X"38",X"04",X"DD",X"36",X"08",X"00",
		X"CD",X"4E",X"01",X"79",X"FE",X"FF",X"20",X"0B",X"FD",X"36",X"04",X"00",X"FD",X"36",X"0C",X"00",
		X"C3",X"11",X"03",X"06",X"00",X"2A",X"F6",X"E4",X"3A",X"E8",X"E4",X"B7",X"20",X"05",X"21",X"00",
		X"00",X"18",X"19",X"57",X"3A",X"02",X"E5",X"B7",X"28",X"12",X"3A",X"E9",X"E4",X"BA",X"20",X"0C",
		X"11",X"30",X"00",X"19",X"3A",X"CD",X"E5",X"FE",X"08",X"20",X"01",X"EB",X"09",X"22",X"F9",X"E4",
		X"01",X"60",X"45",X"09",X"46",X"DD",X"6E",X"00",X"DD",X"7E",X"01",X"C6",X"04",X"67",X"29",X"29",
		X"29",X"0E",X"00",X"CB",X"28",X"CB",X"19",X"DD",X"7E",X"0B",X"B7",X"20",X"04",X"ED",X"42",X"18",
		X"01",X"09",X"29",X"FD",X"74",X"06",X"3E",X"00",X"17",X"FD",X"77",X"07",X"3A",X"F8",X"E4",X"4F",
		X"DD",X"CB",X"17",X"66",X"28",X"01",X"0C",X"3A",X"E8",X"E4",X"B7",X"20",X"04",X"0E",X"03",X"18",
		X"11",X"47",X"3A",X"02",X"E5",X"B7",X"28",X"0A",X"3A",X"E9",X"E4",X"B8",X"20",X"04",X"3A",X"6E",
		X"E5",X"4F",X"CB",X"E1",X"FD",X"71",X"00",X"11",X"B0",X"43",X"2A",X"F9",X"E4",X"19",X"56",X"DD",
		X"7E",X"0B",X"B7",X"20",X"04",X"3E",X"40",X"AA",X"57",X"7A",X"E6",X"C0",X"FD",X"77",X"05",X"2A",
		X"F9",X"E4",X"7A",X"11",X"00",X"42",X"19",X"57",X"5E",X"D5",X"FD",X"73",X"04",X"11",X"C0",X"48",
		X"2A",X"F9",X"E4",X"19",X"AF",X"57",X"5E",X"CB",X"7B",X"28",X"01",X"15",X"DD",X"6E",X"02",X"DD",
		X"66",X"03",X"29",X"29",X"29",X"17",X"6C",X"67",X"19",X"EB",X"21",X"E9",X"00",X"B7",X"ED",X"52",
		X"ED",X"5B",X"E3",X"E5",X"19",X"FD",X"75",X"02",X"FD",X"74",X"03",X"D1",X"CB",X"42",X"28",X"4D",
		X"1C",X"FD",X"73",X"0C",X"FD",X"71",X"08",X"E5",X"01",X"70",X"4A",X"2A",X"F9",X"E4",X"09",X"7E",
		X"06",X"00",X"ED",X"44",X"4F",X"CB",X"79",X"28",X"01",X"05",X"E1",X"09",X"FD",X"75",X"0A",X"FD",
		X"74",X"0B",X"7A",X"E6",X"C0",X"FD",X"77",X"0D",X"01",X"10",X"47",X"2A",X"F9",X"E4",X"09",X"7E",
		X"CB",X"72",X"28",X"02",X"ED",X"44",X"4F",X"06",X"00",X"CB",X"79",X"28",X"01",X"05",X"FD",X"66",
		X"07",X"FD",X"6E",X"06",X"09",X"FD",X"75",X"0E",X"FD",X"74",X"0F",X"18",X"04",X"FD",X"36",X"0C",
		X"00",X"11",X"F0",X"FF",X"FD",X"19",X"01",X"18",X"00",X"DD",X"09",X"21",X"E8",X"E4",X"34",X"3A",
		X"E9",X"E4",X"BE",X"D2",X"B3",X"01",X"3A",X"6A",X"E5",X"FE",X"02",X"C8",X"FD",X"21",X"00",X"E3",
		X"3A",X"17",X"E5",X"87",X"87",X"87",X"21",X"12",X"E5",X"86",X"ED",X"44",X"3C",X"4F",X"06",X"00",
		X"2A",X"E3",X"E5",X"09",X"FD",X"75",X"02",X"FD",X"74",X"03",X"FD",X"36",X"00",X"12",X"3A",X"16",
		X"E5",X"C6",X"04",X"87",X"87",X"87",X"6F",X"26",X"00",X"29",X"FD",X"75",X"06",X"FD",X"74",X"07",
		X"3A",X"10",X"E5",X"FD",X"77",X"04",X"FD",X"21",X"08",X"E3",X"FD",X"36",X"04",X"00",X"FD",X"36",
		X"0C",X"00",X"16",X"14",X"1E",X"02",X"DD",X"21",X"18",X"E5",X"DD",X"7E",X"01",X"FE",X"00",X"28",
		X"3A",X"DD",X"7E",X"03",X"87",X"87",X"87",X"47",X"3E",X"F1",X"90",X"4F",X"06",X"00",X"2A",X"E3",
		X"E5",X"09",X"FD",X"75",X"02",X"FD",X"74",X"03",X"DD",X"7E",X"02",X"C6",X"04",X"87",X"87",X"87",
		X"6F",X"26",X"00",X"29",X"FD",X"75",X"06",X"FD",X"74",X"07",X"FD",X"36",X"00",X"12",X"DD",X"7E",
		X"01",X"FD",X"77",X"04",X"01",X"08",X"00",X"FD",X"09",X"1D",X"C8",X"01",X"04",X"00",X"DD",X"09",
		X"15",X"20",X"B7",X"21",X"9E",X"E5",X"06",X"00",X"7E",X"B7",X"28",X"12",X"35",X"20",X"0F",X"E5",
		X"78",X"87",X"87",X"87",X"5F",X"16",X"00",X"21",X"C4",X"E3",X"19",X"36",X"00",X"E1",X"23",X"04",
		X"78",X"FE",X"08",X"38",X"E3",X"C9",X"21",X"8A",X"E5",X"7E",X"23",X"B6",X"23",X"47",X"7E",X"E6",
		X"F0",X"B0",X"20",X"0B",X"AF",X"77",X"3E",X"01",X"32",X"CE",X"E5",X"CD",X"03",X"32",X"C9",X"0E",
		X"00",X"21",X"B1",X"E6",X"3A",X"8B",X"E5",X"BE",X"20",X"01",X"0C",X"ED",X"5B",X"E1",X"E5",X"21",
		X"8D",X"E5",X"7E",X"93",X"27",X"77",X"2B",X"7E",X"9A",X"27",X"77",X"06",X"02",X"2B",X"7E",X"DE",
		X"00",X"27",X"77",X"10",X"F8",X"CB",X"41",X"C8",X"3A",X"8B",X"E5",X"21",X"B1",X"E6",X"BE",X"C8",
		X"7E",X"FE",X"15",X"20",X"04",X"3E",X"1C",X"18",X"0A",X"FE",X"10",X"20",X"04",X"3E",X"1D",X"18",
		X"02",X"3E",X"1E",X"CD",X"42",X"31",X"7E",X"D6",X"05",X"27",X"77",X"C9",X"3A",X"FC",X"E4",X"B7",
		X"C0",X"21",X"B6",X"E5",X"3A",X"04",X"E5",X"B7",X"20",X"02",X"36",X"FF",X"7E",X"FE",X"80",X"38",
		X"02",X"36",X"18",X"7E",X"21",X"04",X"E5",X"FE",X"09",X"30",X"0D",X"7E",X"FE",X"01",X"28",X"06",
		X"3E",X"01",X"77",X"CD",X"89",X"63",X"18",X"0B",X"7E",X"FE",X"02",X"28",X"06",X"3E",X"02",X"77",
		X"CD",X"89",X"63",X"3A",X"41",X"E4",X"21",X"7B",X"E5",X"BE",X"20",X"0C",X"3A",X"43",X"E4",X"23",
		X"BE",X"20",X"05",X"3E",X"01",X"32",X"AF",X"E6",X"3A",X"AF",X"E6",X"B7",X"C8",X"3A",X"46",X"E4",
		X"FE",X"08",X"C0",X"AF",X"CD",X"89",X"63",X"F1",X"3E",X"00",X"32",X"9D",X"E5",X"3E",X"00",X"CD",
		X"42",X"31",X"3E",X"23",X"CD",X"42",X"31",X"3E",X"54",X"CD",X"3E",X"30",X"CD",X"8D",X"32",X"3A",
		X"00",X"E5",X"B7",X"20",X"47",X"21",X"21",X"D7",X"36",X"05",X"2B",X"36",X"00",X"11",X"22",X"D7",
		X"01",X"3E",X"00",X"ED",X"B0",X"21",X"A1",X"D7",X"36",X"05",X"2B",X"36",X"00",X"11",X"A2",X"D7",
		X"01",X"3E",X"00",X"ED",X"B0",X"21",X"21",X"D8",X"36",X"05",X"2B",X"36",X"00",X"11",X"22",X"D8",
		X"01",X"3E",X"00",X"ED",X"B0",X"0E",X"47",X"21",X"A2",X"D7",X"11",X"F8",X"06",X"CD",X"2D",X"30",
		X"3E",X"1F",X"CD",X"42",X"31",X"0E",X"02",X"CD",X"CF",X"2F",X"18",X"4C",X"3A",X"FF",X"E4",X"B7",
		X"C2",X"64",X"05",X"21",X"25",X"D7",X"36",X"05",X"2B",X"36",X"00",X"11",X"26",X"D7",X"01",X"38",
		X"00",X"ED",X"B0",X"21",X"A5",X"D7",X"36",X"05",X"2B",X"36",X"00",X"11",X"A6",X"D7",X"01",X"38",
		X"00",X"ED",X"B0",X"21",X"25",X"D8",X"36",X"05",X"2B",X"36",X"00",X"11",X"26",X"D8",X"01",X"38",
		X"00",X"ED",X"B0",X"0E",X"47",X"21",X"A6",X"D7",X"11",X"DC",X"06",X"CD",X"2D",X"30",X"3E",X"1F",
		X"CD",X"42",X"31",X"0E",X"01",X"CD",X"CF",X"2F",X"CD",X"03",X"32",X"3A",X"00",X"E5",X"32",X"89",
		X"E5",X"CD",X"89",X"06",X"21",X"6C",X"E5",X"3A",X"8B",X"E5",X"BE",X"38",X"57",X"CD",X"B9",X"32",
		X"21",X"A3",X"D1",X"36",X"05",X"2B",X"36",X"00",X"11",X"A4",X"D1",X"01",X"34",X"00",X"ED",X"B0",
		X"21",X"23",X"D2",X"36",X"05",X"2B",X"36",X"00",X"11",X"24",X"D2",X"01",X"34",X"00",X"ED",X"B0",
		X"21",X"A3",X"D2",X"36",X"05",X"2B",X"36",X"00",X"11",X"A4",X"D2",X"01",X"34",X"00",X"ED",X"B0",
		X"0E",X"47",X"21",X"24",X"D2",X"11",X"6F",X"06",X"CD",X"2D",X"30",X"2A",X"8B",X"E5",X"22",X"B6",
		X"E6",X"3E",X"FF",X"32",X"B5",X"E6",X"3E",X"01",X"32",X"05",X"E5",X"CD",X"E4",X"05",X"2A",X"B6",
		X"E6",X"22",X"8B",X"E5",X"CD",X"E4",X"05",X"21",X"8E",X"E5",X"4E",X"34",X"7E",X"FE",X"61",X"20",
		X"02",X"36",X"49",X"79",X"CD",X"EC",X"31",X"B7",X"C2",X"00",X"5D",X"79",X"E6",X"07",X"CA",X"34",
		X"28",X"C3",X"ED",X"26",X"3A",X"8F",X"E5",X"32",X"89",X"E5",X"3E",X"14",X"32",X"88",X"E5",X"2A",
		X"8B",X"E5",X"7C",X"E6",X"F0",X"B5",X"28",X"32",X"21",X"8C",X"E5",X"7E",X"D6",X"10",X"27",X"77",
		X"2B",X"7E",X"DE",X"00",X"27",X"77",X"01",X"10",X"00",X"CD",X"DB",X"2F",X"CD",X"03",X"32",X"21",
		X"88",X"E5",X"35",X"20",X"DA",X"21",X"8F",X"E5",X"3A",X"89",X"E5",X"BE",X"20",X"05",X"3E",X"11",
		X"CD",X"42",X"31",X"3E",X"04",X"CD",X"30",X"06",X"18",X"C0",X"3E",X"1C",X"CD",X"30",X"06",X"C9",
		X"32",X"B5",X"E5",X"3A",X"05",X"E5",X"B7",X"28",X"2A",X"21",X"B5",X"E6",X"7E",X"FE",X"80",X"38",
		X"02",X"36",X"28",X"7E",X"FE",X"14",X"30",X"12",X"21",X"2B",X"D1",X"36",X"05",X"2B",X"36",X"00",
		X"11",X"2C",X"D1",X"01",X"02",X"00",X"ED",X"B0",X"18",X"09",X"21",X"2A",X"D1",X"11",X"6B",X"06",
		X"CD",X"2D",X"30",X"3A",X"B5",X"E5",X"FE",X"00",X"20",X"C9",X"C9",X"06",X"58",X"32",X"00",X"42",
		X"45",X"4C",X"4F",X"57",X"20",X"48",X"41",X"4C",X"46",X"20",X"54",X"49",X"4D",X"45",X"20",X"43",
		X"4C",X"45",X"41",X"52",X"41",X"4E",X"43",X"45",X"00",X"3E",X"09",X"32",X"88",X"E5",X"21",X"B9",
		X"D8",X"36",X"05",X"2B",X"36",X"00",X"11",X"BA",X"D8",X"01",X"0C",X"00",X"ED",X"B0",X"21",X"39",
		X"D9",X"36",X"05",X"2B",X"36",X"00",X"11",X"3A",X"D9",X"01",X"0C",X"00",X"ED",X"B0",X"0E",X"47",
		X"11",X"26",X"07",X"3A",X"88",X"E5",X"1F",X"30",X"0C",X"11",X"18",X"07",X"3A",X"89",X"E5",X"B7",
		X"20",X"03",X"11",X"1F",X"07",X"21",X"BA",X"D8",X"CD",X"2D",X"30",X"3E",X"0E",X"CD",X"3E",X"30",
		X"21",X"88",X"E5",X"35",X"20",X"D8",X"3E",X"70",X"CD",X"3E",X"30",X"C9",X"59",X"4F",X"55",X"20",
		X"48",X"41",X"56",X"45",X"20",X"4B",X"49",X"4C",X"4C",X"45",X"44",X"20",X"4E",X"4F",X"20",X"45",
		X"4E",X"45",X"4D",X"49",X"45",X"53",X"2E",X"00",X"59",X"4F",X"55",X"20",X"4D",X"41",X"44",X"45",
		X"20",X"49",X"54",X"20",X"57",X"49",X"54",X"48",X"4F",X"55",X"54",X"20",X"45",X"4E",X"54",X"52",
		X"41",X"50",X"50",X"49",X"4E",X"47",X"2E",X"00",X"04",X"31",X"30",X"30",X"30",X"30",X"00",X"04",
		X"32",X"30",X"30",X"30",X"30",X"00",X"20",X"20",X"20",X"20",X"20",X"00",X"CD",X"CE",X"07",X"CD",
		X"1D",X"08",X"CD",X"AA",X"09",X"3A",X"50",X"E4",X"B7",X"C0",X"3A",X"A7",X"E5",X"B7",X"28",X"0E",
		X"3E",X"00",X"32",X"9D",X"E5",X"3E",X"38",X"CD",X"3E",X"30",X"F1",X"C3",X"85",X"68",X"DB",X"04",
		X"CB",X"77",X"C8",X"3E",X"0C",X"32",X"4A",X"E4",X"3E",X"01",X"32",X"9D",X"E5",X"3E",X"00",X"CD",
		X"42",X"31",X"3E",X"06",X"CD",X"42",X"31",X"3E",X"38",X"CD",X"3E",X"30",X"3E",X"00",X"32",X"9D",
		X"E5",X"F1",X"21",X"8F",X"E5",X"35",X"7E",X"FE",X"FF",X"20",X"2A",X"21",X"34",X"D7",X"11",X"A8",
		X"07",X"CD",X"2D",X"30",X"21",X"B4",X"D7",X"11",X"B5",X"07",X"CD",X"2D",X"30",X"21",X"34",X"D8",
		X"11",X"A8",X"07",X"CD",X"2D",X"30",X"3E",X"21",X"CD",X"42",X"31",X"3E",X"8C",X"CD",X"3E",X"30",
		X"3E",X"02",X"32",X"90",X"E5",X"C3",X"E3",X"6A",X"06",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"00",X"06",X"20",X"47",X"41",X"4D",X"45",X"20",X"4F",X"56",X"45",X"52",
		X"20",X"00",X"20",X"54",X"49",X"4D",X"45",X"20",X"4F",X"56",X"45",X"52",X"20",X"00",X"3A",X"CE",
		X"E5",X"B7",X"C8",X"DB",X"04",X"CB",X"77",X"C8",X"F1",X"AF",X"32",X"CE",X"E5",X"32",X"9D",X"E5",
		X"3E",X"00",X"CD",X"42",X"31",X"3E",X"25",X"CD",X"42",X"31",X"21",X"35",X"D7",X"36",X"05",X"2B",
		X"36",X"00",X"11",X"36",X"D7",X"01",X"14",X"00",X"ED",X"B0",X"0E",X"47",X"21",X"B4",X"D7",X"11",
		X"C2",X"07",X"CD",X"2D",X"30",X"21",X"35",X"D8",X"36",X"05",X"2B",X"36",X"00",X"11",X"36",X"D8",
		X"01",X"14",X"00",X"ED",X"B0",X"3E",X"8C",X"CD",X"3E",X"30",X"C3",X"67",X"07",X"2A",X"55",X"E4",
		X"01",X"C0",X"FE",X"09",X"D0",X"AF",X"32",X"50",X"E4",X"32",X"9D",X"E5",X"CD",X"8D",X"32",X"21",
		X"29",X"D7",X"36",X"05",X"2B",X"36",X"00",X"11",X"2A",X"D7",X"01",X"2A",X"00",X"ED",X"B0",X"21",
		X"A9",X"D7",X"36",X"05",X"2B",X"36",X"00",X"11",X"AA",X"D7",X"01",X"2A",X"00",X"ED",X"B0",X"21",
		X"29",X"D8",X"36",X"05",X"2B",X"36",X"00",X"11",X"2A",X"D8",X"01",X"2A",X"00",X"ED",X"B0",X"3E",
		X"02",X"32",X"89",X"E5",X"3E",X"10",X"CD",X"42",X"31",X"3E",X"04",X"32",X"88",X"E5",X"3A",X"88",
		X"E5",X"1F",X"30",X"12",X"21",X"AB",X"D7",X"36",X"05",X"2B",X"36",X"00",X"11",X"AC",X"D7",X"01",
		X"28",X"00",X"ED",X"B0",X"18",X"0B",X"0E",X"47",X"21",X"AA",X"D7",X"11",X"C0",X"08",X"CD",X"2D",
		X"30",X"3E",X"15",X"CD",X"3E",X"30",X"21",X"88",X"E5",X"35",X"20",X"D2",X"21",X"89",X"E5",X"35",
		X"20",X"C2",X"3E",X"10",X"CD",X"42",X"31",X"0E",X"47",X"21",X"AA",X"D7",X"11",X"C0",X"08",X"CD",
		X"2D",X"30",X"3E",X"54",X"CD",X"3E",X"30",X"3A",X"8F",X"E5",X"B7",X"C0",X"CD",X"B9",X"32",X"C9",
		X"59",X"4F",X"55",X"20",X"41",X"52",X"45",X"20",X"42",X"4F",X"55",X"4E",X"44",X"20",X"54",X"4F",
		X"20",X"44",X"49",X"45",X"2E",X"00",X"DB",X"03",X"2F",X"47",X"E6",X"03",X"32",X"DF",X"E5",X"78",
		X"1F",X"1F",X"E6",X"03",X"4F",X"06",X"00",X"21",X"F0",X"08",X"09",X"7E",X"32",X"E0",X"E5",X"C9",
		X"02",X"01",X"03",X"04",X"DB",X"03",X"2F",X"1F",X"1F",X"1F",X"1F",X"47",X"21",X"AF",X"E5",X"DB",
		X"04",X"CB",X"57",X"20",X"11",X"78",X"3C",X"E6",X"03",X"77",X"23",X"78",X"1F",X"1F",X"E6",X"03",
		X"FE",X"02",X"DE",X"F5",X"77",X"C9",X"78",X"3C",X"E6",X"0F",X"CB",X"5F",X"28",X"01",X"3C",X"77",
		X"23",X"77",X"C9",X"21",X"AD",X"E5",X"11",X"AF",X"E5",X"DB",X"00",X"CD",X"58",X"09",X"21",X"AE",
		X"E5",X"13",X"DB",X"02",X"1F",X"F6",X"04",X"CD",X"58",X"09",X"3A",X"B9",X"E5",X"47",X"21",X"AB",
		X"E5",X"7E",X"B7",X"28",X"05",X"35",X"3E",X"02",X"B0",X"47",X"23",X"7E",X"B7",X"28",X"05",X"35",
		X"3E",X"04",X"B0",X"47",X"78",X"D3",X"01",X"C9",X"1F",X"1F",X"1F",X"CB",X"16",X"1F",X"CB",X"16",
		X"7E",X"E6",X"55",X"FE",X"50",X"20",X"2B",X"2B",X"2B",X"36",X"0C",X"3A",X"B2",X"E6",X"B7",X"20",
		X"08",X"3E",X"12",X"D3",X"00",X"F6",X"80",X"D3",X"00",X"1A",X"FE",X"01",X"28",X"12",X"FE",X"08",
		X"30",X"0C",X"21",X"B1",X"E5",X"34",X"BE",X"C0",X"AF",X"77",X"3E",X"01",X"18",X"02",X"D6",X"08",
		X"18",X"0D",X"7E",X"E6",X"AA",X"C0",X"21",X"B3",X"E5",X"34",X"7E",X"E6",X"0F",X"C0",X"3C",X"21",
		X"B2",X"E5",X"86",X"27",X"30",X"02",X"3E",X"99",X"77",X"C9",X"DB",X"04",X"CB",X"6F",X"C0",X"CB",
		X"67",X"C8",X"DB",X"00",X"CB",X"47",X"C0",X"F1",X"F1",X"AF",X"32",X"9D",X"E5",X"3E",X"00",X"CD",
		X"42",X"31",X"21",X"10",X"D0",X"36",X"00",X"54",X"5D",X"13",X"01",X"EF",X"13",X"ED",X"B0",X"21",
		X"22",X"D7",X"11",X"29",X"0A",X"CD",X"2D",X"30",X"21",X"1A",X"D9",X"11",X"48",X"0A",X"CD",X"2D",
		X"30",X"11",X"00",X"00",X"0E",X"04",X"3A",X"8E",X"E5",X"21",X"60",X"D9",X"CD",X"48",X"30",X"21",
		X"8E",X"E5",X"DB",X"01",X"CB",X"7F",X"28",X"0E",X"CB",X"42",X"28",X"08",X"16",X"00",X"7E",X"FE",
		X"02",X"38",X"01",X"35",X"18",X"02",X"16",X"01",X"DB",X"01",X"CB",X"6F",X"28",X"09",X"CB",X"43",
		X"28",X"03",X"1E",X"00",X"34",X"18",X"02",X"1E",X"01",X"3E",X"01",X"CD",X"3E",X"30",X"DB",X"00",
		X"CB",X"4F",X"20",X"C0",X"7E",X"3D",X"C3",X"D4",X"05",X"02",X"53",X"45",X"4C",X"45",X"43",X"54",
		X"20",X"42",X"55",X"54",X"54",X"4F",X"4E",X"20",X"54",X"4F",X"20",X"43",X"48",X"41",X"4E",X"47",
		X"45",X"20",X"52",X"4F",X"55",X"4E",X"44",X"00",X"02",X"44",X"49",X"47",X"4C",X"45",X"46",X"54",
		X"2D",X"2D",X"44",X"4F",X"57",X"4E",X"20",X"20",X"44",X"49",X"47",X"52",X"49",X"47",X"48",X"54",
		X"2D",X"2D",X"55",X"50",X"20",X"20",X"4C",X"45",X"56",X"45",X"4C",X"2D",X"30",X"30",X"00",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"3A",X"A7",X"E5",X"B7",X"28",X"0E",X"CD",X"12",X"5C",X"32",X"4D",X"E4",X"FE",X"FF",X"20",X"04",
		X"AF",X"32",X"50",X"E4",X"2A",X"44",X"E4",X"7D",X"6C",X"2C",X"2C",X"CD",X"D5",X"62",X"7E",X"2A",
		X"55",X"E4",X"FE",X"0E",X"38",X"03",X"23",X"18",X"03",X"21",X"00",X"00",X"22",X"55",X"E4",X"DD",
		X"21",X"40",X"E4",X"21",X"08",X"E5",X"7E",X"B7",X"28",X"01",X"35",X"21",X"06",X"E5",X"7E",X"B7",
		X"28",X"18",X"35",X"3A",X"0A",X"E5",X"DD",X"BE",X"0B",X"20",X"0F",X"21",X"0B",X"E5",X"3A",X"44",
		X"E4",X"BE",X"28",X"06",X"77",X"3E",X"0C",X"CD",X"73",X"30",X"3A",X"4E",X"E4",X"B7",X"FA",X"B4",
		X"0F",X"C2",X"43",X"10",X"21",X"4C",X"E4",X"7E",X"B7",X"28",X"11",X"35",X"C0",X"36",X"08",X"21",
		X"4A",X"E4",X"34",X"7E",X"E6",X"FC",X"FE",X"14",X"C8",X"36",X"14",X"C9",X"3A",X"54",X"E4",X"FE",
		X"02",X"20",X"0D",X"06",X"1C",X"CD",X"9F",X"10",X"D0",X"AF",X"32",X"54",X"E4",X"CD",X"37",X"12",
		X"3A",X"54",X"E4",X"FE",X"01",X"20",X"0E",X"CD",X"0E",X"12",X"06",X"20",X"CD",X"9F",X"10",X"D0",
		X"3E",X"03",X"32",X"54",X"E4",X"AF",X"32",X"51",X"E4",X"3A",X"44",X"E4",X"2A",X"45",X"E4",X"CD",
		X"00",X"2D",X"06",X"F8",X"0E",X"10",X"CD",X"8D",X"2E",X"CA",X"9F",X"0C",X"AF",X"32",X"87",X"E5",
		X"32",X"54",X"E4",X"7E",X"E6",X"FC",X"FE",X"18",X"20",X"13",X"3E",X"01",X"32",X"87",X"E5",X"3A",
		X"42",X"E4",X"B7",X"20",X"08",X"3E",X"01",X"32",X"51",X"E4",X"CA",X"9F",X"0C",X"3A",X"45",X"E4",
		X"FE",X"1D",X"30",X"0E",X"1A",X"E6",X"F8",X"FE",X"10",X"28",X"07",X"1A",X"E6",X"F8",X"FE",X"08",
		X"20",X"0D",X"3E",X"01",X"32",X"87",X"E5",X"3A",X"42",X"E4",X"FE",X"80",X"DA",X"9F",X"0C",X"2A",
		X"47",X"E4",X"3A",X"46",X"E4",X"CD",X"15",X"2D",X"DA",X"B1",X"0C",X"21",X"4F",X"E4",X"7E",X"B7",
		X"20",X"06",X"34",X"3E",X"15",X"CD",X"42",X"31",X"3E",X"0C",X"32",X"4A",X"E4",X"21",X"09",X"E5",
		X"7E",X"B7",X"28",X"04",X"35",X"C3",X"B1",X"0C",X"CD",X"0E",X"12",X"2A",X"42",X"E4",X"7C",X"11",
		X"1E",X"00",X"19",X"22",X"42",X"E4",X"BC",X"28",X"0A",X"3A",X"87",X"E5",X"B7",X"28",X"04",X"AF",
		X"32",X"42",X"E4",X"2A",X"42",X"E4",X"29",X"7C",X"3C",X"1F",X"32",X"45",X"E4",X"29",X"29",X"7C",
		X"32",X"46",X"E4",X"CD",X"88",X"11",X"3A",X"42",X"E4",X"B7",X"C0",X"3A",X"44",X"E4",X"2A",X"45",
		X"E4",X"CD",X"00",X"2D",X"3A",X"45",X"E4",X"FE",X"1D",X"30",X"06",X"1A",X"E6",X"F8",X"FE",X"08",
		X"C0",X"15",X"0E",X"04",X"CD",X"A9",X"2E",X"C0",X"1D",X"1D",X"1D",X"1D",X"3A",X"44",X"E4",X"B7",
		X"28",X"06",X"1A",X"E6",X"F8",X"FE",X"08",X"C0",X"3A",X"44",X"E4",X"FE",X"17",X"30",X"0A",X"7B",
		X"C6",X"08",X"5F",X"1A",X"E6",X"F8",X"FE",X"08",X"C0",X"3E",X"08",X"32",X"4C",X"E4",X"C9",X"21",
		X"4F",X"E4",X"7E",X"B7",X"28",X"07",X"36",X"00",X"3E",X"16",X"CD",X"42",X"31",X"AF",X"32",X"52",
		X"E4",X"3A",X"4D",X"E4",X"CB",X"7F",X"C2",X"42",X"0F",X"CB",X"6F",X"C2",X"CF",X"0F",X"CB",X"5F",
		X"28",X"06",X"CD",X"4C",X"0E",X"D8",X"18",X"08",X"CB",X"57",X"28",X"04",X"CD",X"B7",X"0E",X"D8",
		X"3A",X"4D",X"E4",X"CB",X"47",X"C2",X"5E",X"0D",X"CB",X"4F",X"C2",X"21",X"0D",X"3A",X"44",X"E4",
		X"2A",X"45",X"E4",X"CD",X"00",X"2D",X"1A",X"E6",X"F8",X"FE",X"08",X"20",X"0B",X"3E",X"12",X"32",
		X"4A",X"E4",X"3E",X"01",X"32",X"49",X"E4",X"C9",X"06",X"F8",X"0E",X"10",X"CD",X"8D",X"2E",X"20",
		X"0D",X"15",X"1A",X"E6",X"F8",X"FE",X"10",X"C0",X"3E",X"08",X"32",X"4A",X"E4",X"C9",X"7E",X"E6",
		X"FC",X"FE",X"18",X"20",X"06",X"3E",X"07",X"32",X"4A",X"E4",X"C9",X"3E",X"12",X"32",X"4A",X"E4",
		X"C9",X"AF",X"32",X"87",X"E5",X"3A",X"44",X"E4",X"2A",X"45",X"E4",X"CD",X"00",X"2D",X"3A",X"44",
		X"E4",X"B7",X"28",X"0E",X"15",X"1B",X"1B",X"1B",X"1B",X"06",X"F8",X"0E",X"08",X"CD",X"71",X"2E",
		X"20",X"0C",X"3E",X"01",X"32",X"87",X"E5",X"3A",X"40",X"E4",X"3D",X"FE",X"7F",X"D0",X"3E",X"01",
		X"32",X"4B",X"E4",X"CD",X"37",X"12",X"CD",X"D4",X"0D",X"11",X"EC",X"FF",X"18",X"3D",X"AF",X"32",
		X"87",X"E5",X"3A",X"44",X"E4",X"2A",X"45",X"E4",X"CD",X"00",X"2D",X"3A",X"44",X"E4",X"FE",X"17",
		X"30",X"0E",X"15",X"13",X"13",X"13",X"13",X"06",X"F8",X"0E",X"08",X"CD",X"71",X"2E",X"20",X"0E",
		X"3E",X"01",X"32",X"87",X"E5",X"3A",X"40",X"E4",X"FE",X"80",X"30",X"02",X"B7",X"C9",X"AF",X"32",
		X"4B",X"E4",X"CD",X"37",X"12",X"CD",X"D4",X"0D",X"11",X"14",X"00",X"2A",X"40",X"E4",X"7C",X"19",
		X"22",X"40",X"E4",X"BC",X"28",X"14",X"3A",X"87",X"E5",X"B7",X"28",X"0E",X"2A",X"40",X"E4",X"7D",
		X"FE",X"80",X"38",X"01",X"24",X"2E",X"00",X"22",X"40",X"E4",X"2A",X"40",X"E4",X"29",X"7C",X"3C",
		X"1F",X"32",X"44",X"E4",X"29",X"29",X"7C",X"32",X"47",X"E4",X"CD",X"88",X"11",X"06",X"00",X"CD",
		X"F1",X"10",X"37",X"C9",X"3A",X"51",X"E4",X"B7",X"C8",X"F1",X"3A",X"4A",X"E4",X"E6",X"FC",X"21",
		X"49",X"E4",X"FE",X"2C",X"28",X"02",X"36",X"01",X"35",X"C0",X"21",X"4A",X"E4",X"34",X"7E",X"E6",
		X"FC",X"FE",X"2C",X"28",X"02",X"36",X"2C",X"7E",X"D6",X"18",X"4F",X"06",X"00",X"21",X"20",X"4C",
		X"09",X"7E",X"32",X"49",X"E4",X"21",X"D0",X"4D",X"09",X"7E",X"87",X"87",X"87",X"87",X"5F",X"3A",
		X"87",X"E5",X"57",X"2A",X"40",X"E4",X"3A",X"4B",X"E4",X"B7",X"7D",X"28",X"0D",X"93",X"30",X"08",
		X"CB",X"42",X"28",X"03",X"AF",X"18",X"01",X"25",X"18",X"09",X"83",X"30",X"06",X"24",X"CB",X"42",
		X"28",X"01",X"AF",X"6F",X"22",X"40",X"E4",X"2A",X"40",X"E4",X"29",X"7C",X"3C",X"1F",X"32",X"44",
		X"E4",X"29",X"29",X"7C",X"32",X"47",X"E4",X"CD",X"88",X"11",X"37",X"C9",X"AF",X"32",X"87",X"E5",
		X"3A",X"44",X"E4",X"2A",X"45",X"E4",X"CD",X"00",X"2D",X"06",X"F8",X"0E",X"10",X"CD",X"8D",X"2E",
		X"20",X"14",X"3A",X"45",X"E4",X"FE",X"01",X"28",X"16",X"15",X"15",X"1A",X"E6",X"F8",X"FE",X"08",
		X"28",X"0D",X"18",X"17",X"18",X"09",X"1A",X"E6",X"F8",X"FE",X"10",X"28",X"02",X"B7",X"C9",X"3A",
		X"42",X"E4",X"3D",X"FE",X"7F",X"D0",X"3E",X"01",X"32",X"87",X"E5",X"CD",X"0E",X"12",X"3A",X"44",
		X"E4",X"2A",X"45",X"E4",X"CD",X"00",X"2D",X"15",X"1A",X"E6",X"F8",X"11",X"E2",X"FF",X"FE",X"10",
		X"CA",X"07",X"0F",X"21",X"54",X"E4",X"7E",X"FE",X"03",X"C2",X"07",X"0F",X"35",X"3E",X"1C",X"32",
		X"4A",X"E4",X"CD",X"AB",X"10",X"37",X"C9",X"AF",X"32",X"87",X"E5",X"3A",X"45",X"E4",X"FE",X"1D",
		X"30",X"07",X"1A",X"E6",X"F8",X"FE",X"08",X"20",X"0E",X"3A",X"42",X"E4",X"FE",X"80",X"30",X"02",
		X"B7",X"C9",X"3E",X"01",X"32",X"87",X"E5",X"CD",X"0E",X"12",X"3A",X"44",X"E4",X"2A",X"43",X"E4",
		X"CD",X"00",X"2D",X"1A",X"15",X"E6",X"F8",X"FE",X"10",X"1A",X"11",X"1E",X"00",X"20",X"18",X"E6",
		X"F8",X"FE",X"10",X"28",X"12",X"21",X"54",X"E4",X"7E",X"B7",X"20",X"0B",X"34",X"3E",X"20",X"32",
		X"4A",X"E4",X"CD",X"AB",X"10",X"37",X"C9",X"2A",X"42",X"E4",X"7C",X"19",X"22",X"42",X"E4",X"BC",
		X"28",X"11",X"3A",X"87",X"E5",X"B7",X"28",X"0B",X"7D",X"FE",X"80",X"38",X"01",X"24",X"2E",X"00",
		X"22",X"42",X"E4",X"2A",X"42",X"E4",X"29",X"7C",X"3C",X"1F",X"32",X"45",X"E4",X"29",X"29",X"7C",
		X"32",X"46",X"E4",X"CD",X"88",X"11",X"06",X"08",X"CD",X"F1",X"10",X"3E",X"03",X"32",X"54",X"E4",
		X"37",X"C9",X"AF",X"32",X"0F",X"E5",X"3A",X"45",X"E4",X"FE",X"1C",X"D0",X"3A",X"44",X"E4",X"B7",
		X"C8",X"3A",X"45",X"E4",X"6F",X"C6",X"03",X"32",X"17",X"E5",X"3A",X"44",X"E4",X"3D",X"32",X"16",
		X"E5",X"CD",X"00",X"2D",X"06",X"FC",X"0E",X"08",X"CD",X"7F",X"2E",X"C0",X"ED",X"53",X"13",X"E5",
		X"15",X"06",X"F8",X"0E",X"00",X"CD",X"7F",X"2E",X"C0",X"3E",X"10",X"32",X"4A",X"E4",X"14",X"1C",
		X"1C",X"1C",X"1C",X"1A",X"E6",X"F8",X"FE",X"08",X"28",X"17",X"2C",X"2C",X"2C",X"2C",X"7E",X"E6",
		X"FC",X"FE",X"18",X"28",X"07",X"7E",X"E6",X"F8",X"FE",X"10",X"20",X"05",X"3E",X"11",X"32",X"4A",
		X"E4",X"3E",X"FF",X"32",X"4E",X"E4",X"21",X"40",X"01",X"22",X"11",X"E5",X"3E",X"01",X"32",X"4B",
		X"E4",X"32",X"07",X"E5",X"3A",X"0F",X"E5",X"FE",X"0E",X"D2",X"59",X"10",X"2A",X"46",X"E4",X"7D",
		X"C6",X"08",X"6F",X"7C",X"D6",X"06",X"CD",X"EF",X"2D",X"DA",X"92",X"10",X"C3",X"59",X"10",X"AF",
		X"32",X"0F",X"E5",X"3A",X"45",X"E4",X"FE",X"1C",X"D0",X"3A",X"44",X"E4",X"FE",X"17",X"D0",X"3A",
		X"45",X"E4",X"6F",X"C6",X"03",X"32",X"17",X"E5",X"3A",X"44",X"E4",X"3C",X"32",X"16",X"E5",X"CD",
		X"00",X"2D",X"06",X"FC",X"0E",X"08",X"CD",X"7F",X"2E",X"C0",X"ED",X"53",X"13",X"E5",X"15",X"06",
		X"F8",X"0E",X"00",X"CD",X"7F",X"2E",X"C0",X"3E",X"10",X"32",X"4A",X"E4",X"14",X"1D",X"1D",X"1D",
		X"1D",X"1A",X"E6",X"F8",X"FE",X"08",X"28",X"17",X"2D",X"2D",X"2D",X"2D",X"7E",X"E6",X"FC",X"FE",
		X"18",X"28",X"07",X"7E",X"E6",X"F8",X"FE",X"10",X"20",X"05",X"3E",X"11",X"32",X"4A",X"E4",X"3E",
		X"01",X"32",X"4E",X"E4",X"21",X"40",X"01",X"22",X"11",X"E5",X"AF",X"32",X"4B",X"E4",X"3E",X"01",
		X"32",X"07",X"E5",X"3A",X"0F",X"E5",X"FE",X"0E",X"30",X"0F",X"2A",X"46",X"E4",X"7D",X"C6",X"08",
		X"6F",X"7C",X"C6",X"06",X"CD",X"31",X"2E",X"38",X"39",X"21",X"07",X"E5",X"7E",X"B7",X"28",X"07",
		X"36",X"00",X"3E",X"01",X"CD",X"42",X"31",X"CD",X"0E",X"12",X"CD",X"37",X"12",X"3A",X"0F",X"E5",
		X"FE",X"14",X"D2",X"03",X"11",X"21",X"10",X"E5",X"36",X"F3",X"3A",X"0F",X"E5",X"1F",X"1F",X"30",
		X"02",X"36",X"F2",X"2A",X"11",X"E5",X"11",X"C0",X"00",X"19",X"22",X"11",X"E5",X"21",X"0F",X"E5",
		X"34",X"C9",X"3E",X"00",X"32",X"10",X"E5",X"AF",X"32",X"4E",X"E4",X"32",X"07",X"E5",X"C9",X"21",
		X"49",X"E4",X"35",X"28",X"02",X"B7",X"C9",X"21",X"4A",X"E4",X"34",X"3A",X"4A",X"E4",X"D6",X"18",
		X"4F",X"06",X"00",X"21",X"20",X"4C",X"09",X"7E",X"32",X"49",X"E4",X"B7",X"20",X"07",X"3E",X"01",
		X"32",X"49",X"E4",X"37",X"C9",X"21",X"A8",X"4E",X"09",X"56",X"1E",X"00",X"CB",X"2A",X"CB",X"1B",
		X"CB",X"2A",X"CB",X"1B",X"CB",X"2A",X"CB",X"1B",X"2A",X"42",X"E4",X"19",X"22",X"42",X"E4",X"2A",
		X"42",X"E4",X"29",X"7C",X"3C",X"1F",X"32",X"45",X"E4",X"29",X"29",X"7C",X"32",X"46",X"E4",X"B7",
		X"C9",X"21",X"49",X"E4",X"35",X"C0",X"36",X"06",X"21",X"4A",X"E4",X"34",X"7E",X"E6",X"FC",X"B8",
		X"C8",X"70",X"C9",X"AF",X"32",X"4E",X"E4",X"32",X"0C",X"E5",X"3D",X"32",X"0B",X"E5",X"CD",X"DD",
		X"0C",X"ED",X"5B",X"13",X"E5",X"3E",X"04",X"CD",X"BE",X"2F",X"3E",X"00",X"32",X"10",X"E5",X"21",
		X"18",X"E5",X"06",X"14",X"7E",X"B7",X"28",X"07",X"23",X"23",X"23",X"23",X"10",X"F6",X"C9",X"36",
		X"A0",X"23",X"23",X"3A",X"16",X"E5",X"77",X"5F",X"23",X"3A",X"17",X"E5",X"77",X"57",X"2A",X"71",
		X"E5",X"B7",X"ED",X"52",X"C0",X"22",X"71",X"E5",X"3E",X"01",X"32",X"02",X"E5",X"21",X"E9",X"E4",
		X"7E",X"FD",X"21",X"58",X"E4",X"01",X"18",X"00",X"FD",X"09",X"3D",X"20",X"FB",X"34",X"FD",X"77",
		X"00",X"FD",X"77",X"02",X"FD",X"73",X"01",X"FD",X"73",X"04",X"15",X"FD",X"72",X"03",X"FD",X"72",
		X"05",X"7B",X"87",X"87",X"87",X"FD",X"77",X"07",X"7A",X"87",X"87",X"87",X"FD",X"77",X"06",X"FD",
		X"36",X"09",X"01",X"FD",X"36",X"0C",X"B0",X"C9",X"3A",X"51",X"E4",X"B7",X"20",X"18",X"3A",X"40",
		X"E4",X"FE",X"80",X"38",X"02",X"ED",X"44",X"FE",X"14",X"D0",X"3A",X"42",X"E4",X"FE",X"80",X"38",
		X"02",X"ED",X"44",X"FE",X"1E",X"D0",X"3A",X"44",X"E4",X"2A",X"45",X"E4",X"CD",X"00",X"2D",X"15",
		X"1A",X"E6",X"FC",X"FE",X"60",X"20",X"20",X"CD",X"83",X"2F",X"ED",X"5F",X"FE",X"33",X"38",X"04",
		X"3E",X"08",X"18",X"0A",X"FE",X"0D",X"38",X"04",X"3E",X"09",X"18",X"02",X"3E",X"0A",X"CD",X"73",
		X"30",X"3E",X"02",X"CD",X"42",X"31",X"C9",X"FE",X"70",X"C0",X"21",X"FC",X"E4",X"35",X"CD",X"5C",
		X"2F",X"0E",X"00",X"14",X"1A",X"FE",X"04",X"20",X"02",X"0E",X"04",X"21",X"0D",X"E5",X"3A",X"08",
		X"E5",X"B7",X"20",X"04",X"36",X"00",X"18",X"06",X"7E",X"FE",X"03",X"30",X"01",X"34",X"7E",X"81",
		X"CD",X"73",X"30",X"3E",X"13",X"32",X"08",X"E5",X"3E",X"02",X"CD",X"42",X"31",X"C9",X"2A",X"40",
		X"E4",X"7D",X"FE",X"80",X"30",X"07",X"D6",X"14",X"30",X"01",X"AF",X"18",X"06",X"C6",X"14",X"30",
		X"02",X"24",X"AF",X"6F",X"22",X"40",X"E4",X"29",X"7C",X"3C",X"1F",X"32",X"44",X"E4",X"29",X"29",
		X"7C",X"32",X"47",X"E4",X"C3",X"88",X"11",X"3A",X"52",X"E4",X"B7",X"C0",X"2A",X"42",X"E4",X"7D",
		X"FE",X"80",X"30",X"07",X"D6",X"1E",X"30",X"01",X"AF",X"18",X"06",X"C6",X"1E",X"30",X"02",X"24",
		X"AF",X"6F",X"22",X"42",X"E4",X"29",X"7C",X"3C",X"1F",X"32",X"45",X"E4",X"29",X"29",X"7C",X"32",
		X"46",X"E4",X"C3",X"88",X"11",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"3A",X"E9",X"E4",X"32",X"E8",X"E4",X"DD",X"21",X"58",X"E4",X"CD",X"19",X"13",X"11",X"18",X"00",
		X"DD",X"19",X"21",X"E8",X"E4",X"35",X"20",X"F2",X"C9",X"21",X"6D",X"E5",X"36",X"00",X"3A",X"02",
		X"E5",X"B7",X"28",X"19",X"3A",X"E8",X"E4",X"FE",X"01",X"20",X"12",X"34",X"3A",X"03",X"E5",X"B7",
		X"28",X"0B",X"DD",X"7E",X"0C",X"FE",X"20",X"20",X"04",X"DD",X"36",X"0C",X"40",X"DD",X"7E",X"0E",
		X"B7",X"C0",X"3A",X"F5",X"E4",X"B7",X"28",X"03",X"DD",X"34",X"17",X"DD",X"7E",X"0C",X"B7",X"28",
		X"32",X"DD",X"35",X"0C",X"DD",X"7E",X"0C",X"FE",X"20",X"DA",X"23",X"15",X"DD",X"6E",X"07",X"DD",
		X"7E",X"06",X"CD",X"F2",X"2E",X"DD",X"7E",X"0C",X"FE",X"B0",X"D0",X"DD",X"35",X"09",X"C0",X"DD",
		X"36",X"09",X"08",X"DD",X"34",X"0A",X"DD",X"7E",X"0A",X"E6",X"FC",X"FE",X"14",X"C8",X"DD",X"36",
		X"0A",X"14",X"C9",X"DD",X"7E",X"14",X"FE",X"14",X"20",X"0F",X"CD",X"F7",X"18",X"D8",X"06",X"1C",
		X"CD",X"66",X"1A",X"D0",X"DD",X"36",X"14",X"00",X"C9",X"DD",X"7E",X"14",X"FE",X"01",X"20",X"12",
		X"CD",X"C1",X"1B",X"CD",X"F7",X"18",X"D8",X"06",X"20",X"CD",X"66",X"1A",X"D0",X"DD",X"36",X"14",
		X"15",X"C9",X"DD",X"7E",X"15",X"FE",X"02",X"20",X"19",X"CD",X"C1",X"1B",X"CD",X"F7",X"18",X"D8",
		X"06",X"28",X"CD",X"66",X"1A",X"D0",X"DD",X"36",X"15",X"00",X"DD",X"34",X"09",X"DD",X"36",X"0F",
		X"02",X"C9",X"DD",X"7E",X"15",X"FE",X"01",X"20",X"0F",X"CD",X"F7",X"18",X"D8",X"06",X"24",X"CD",
		X"66",X"1A",X"D0",X"DD",X"36",X"15",X"03",X"C9",X"DD",X"7E",X"06",X"DD",X"6E",X"07",X"CD",X"9E",
		X"2D",X"DA",X"75",X"15",X"DD",X"7E",X"04",X"DD",X"6E",X"05",X"CD",X"00",X"2D",X"06",X"F8",X"0E",
		X"10",X"CD",X"8D",X"2E",X"CA",X"75",X"15",X"AF",X"32",X"87",X"E5",X"DD",X"77",X"14",X"7E",X"E6",
		X"FC",X"FE",X"18",X"20",X"0C",X"3E",X"01",X"32",X"87",X"E5",X"DD",X"7E",X"02",X"B7",X"CA",X"75",
		X"15",X"DD",X"7E",X"05",X"FE",X"1D",X"30",X"29",X"1A",X"E6",X"F8",X"FE",X"10",X"28",X"22",X"1A",
		X"E6",X"F8",X"FE",X"08",X"28",X"1B",X"DD",X"7E",X"16",X"B7",X"28",X"08",X"3C",X"DD",X"BE",X"05",
		X"30",X"1C",X"18",X"0D",X"1A",X"FE",X"04",X"20",X"15",X"DD",X"7E",X"05",X"DD",X"77",X"16",X"18",
		X"0D",X"3E",X"01",X"32",X"87",X"E5",X"DD",X"7E",X"02",X"FE",X"80",X"DA",X"75",X"15",X"DD",X"36",
		X"10",X"00",X"CD",X"C1",X"1B",X"DD",X"7E",X"02",X"C6",X"15",X"DD",X"77",X"02",X"30",X"0D",X"DD",
		X"34",X"03",X"3A",X"87",X"E5",X"B7",X"28",X"04",X"AF",X"DD",X"77",X"02",X"DD",X"6E",X"02",X"DD",
		X"66",X"03",X"29",X"7C",X"3C",X"1F",X"DD",X"77",X"05",X"29",X"29",X"7C",X"DD",X"77",X"06",X"DD",
		X"7E",X"06",X"DD",X"6E",X"07",X"CD",X"D3",X"2E",X"CD",X"39",X"1B",X"06",X"0C",X"CD",X"2E",X"1A",
		X"DD",X"7E",X"04",X"DD",X"6E",X"05",X"CD",X"00",X"2D",X"24",X"7E",X"25",X"FE",X"04",X"20",X"3E",
		X"DD",X"7E",X"0D",X"B7",X"28",X"19",X"DD",X"36",X"0D",X"00",X"EB",X"06",X"FC",X"0E",X"00",X"CD",
		X"7F",X"2E",X"20",X"04",X"CD",X"0E",X"2F",X"C9",X"21",X"FC",X"E4",X"35",X"C9",X"18",X"1F",X"3A",
		X"6D",X"E5",X"B7",X"28",X"19",X"3A",X"03",X"E5",X"B7",X"20",X"13",X"3E",X"01",X"32",X"03",X"E5",
		X"EB",X"06",X"FC",X"0E",X"00",X"CD",X"7F",X"2E",X"20",X"03",X"CD",X"35",X"2F",X"C9",X"DD",X"7E",
		X"02",X"B7",X"C0",X"15",X"1A",X"FE",X"04",X"C0",X"3A",X"87",X"E5",X"B7",X"C8",X"DD",X"36",X"16",
		X"00",X"DD",X"36",X"0C",X"C0",X"DD",X"36",X"10",X"00",X"DD",X"36",X"0A",X"10",X"3E",X"05",X"CD",
		X"42",X"31",X"3A",X"6D",X"E5",X"B7",X"C0",X"01",X"00",X"01",X"CD",X"DB",X"2F",X"3E",X"01",X"32",
		X"00",X"E5",X"C9",X"B7",X"28",X"3C",X"FE",X"1F",X"20",X"0F",X"DD",X"36",X"10",X"01",X"DD",X"36",
		X"0F",X"FE",X"DD",X"35",X"05",X"DD",X"35",X"05",X"C9",X"FE",X"18",X"38",X"06",X"DD",X"7E",X"0F",
		X"FE",X"FE",X"C8",X"DD",X"36",X"10",X"00",X"DD",X"34",X"05",X"DD",X"34",X"05",X"DD",X"7E",X"0F",
		X"DD",X"77",X"0B",X"FE",X"FE",X"38",X"04",X"DD",X"77",X"0C",X"C9",X"DD",X"36",X"0A",X"18",X"CD",
		X"76",X"1A",X"DD",X"36",X"0C",X"01",X"CD",X"F7",X"18",X"D8",X"06",X"18",X"CD",X"66",X"1A",X"D0",
		X"DD",X"36",X"0C",X"00",X"C9",X"DD",X"36",X"16",X"00",X"DD",X"36",X"10",X"01",X"DD",X"7E",X"0F",
		X"B7",X"CA",X"85",X"17",X"3D",X"CA",X"29",X"17",X"3D",X"CA",X"5D",X"16",X"3D",X"CA",X"9A",X"15",
		X"DD",X"6E",X"07",X"DD",X"7E",X"06",X"CD",X"F2",X"2E",X"C9",X"AF",X"32",X"87",X"E5",X"DD",X"7E",
		X"05",X"FE",X"01",X"28",X"23",X"DD",X"7E",X"04",X"DD",X"6E",X"05",X"CD",X"00",X"2D",X"06",X"F8",
		X"0E",X"10",X"CD",X"8D",X"2E",X"20",X"0B",X"15",X"15",X"1A",X"E6",X"F8",X"FE",X"08",X"20",X"14",
		X"18",X"06",X"1A",X"E6",X"F8",X"FE",X"10",X"C0",X"DD",X"7E",X"02",X"3D",X"FE",X"7F",X"D0",X"3E",
		X"01",X"32",X"87",X"E5",X"CD",X"C1",X"1B",X"DD",X"7E",X"04",X"DD",X"6E",X"03",X"CD",X"00",X"2D",
		X"24",X"24",X"7E",X"E6",X"F8",X"FE",X"10",X"20",X"30",X"1A",X"E6",X"F8",X"FE",X"10",X"20",X"29",
		X"15",X"1A",X"E6",X"F8",X"FE",X"10",X"28",X"21",X"DD",X"7E",X"14",X"FE",X"15",X"20",X"1A",X"DD",
		X"35",X"14",X"DD",X"46",X"0A",X"DD",X"4E",X"09",X"C5",X"DD",X"36",X"0A",X"1C",X"CD",X"76",X"1A",
		X"C1",X"30",X"41",X"DD",X"70",X"0A",X"DD",X"71",X"09",X"DD",X"7E",X"02",X"D6",X"15",X"DD",X"77",
		X"02",X"30",X"0F",X"3A",X"87",X"E5",X"B7",X"28",X"06",X"AF",X"DD",X"77",X"02",X"18",X"03",X"DD",
		X"35",X"03",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"29",X"7C",X"3C",X"1F",X"DD",X"77",X"05",X"29",
		X"29",X"7C",X"DD",X"77",X"06",X"CD",X"39",X"1B",X"CD",X"7A",X"1B",X"06",X"08",X"CD",X"2E",X"1A",
		X"DD",X"36",X"14",X"15",X"DD",X"7E",X"06",X"DD",X"6E",X"07",X"C3",X"D3",X"2E",X"DD",X"7E",X"06",
		X"DD",X"6E",X"07",X"CD",X"9E",X"2D",X"D8",X"AF",X"32",X"87",X"E5",X"DD",X"7E",X"05",X"FE",X"1D",
		X"30",X"10",X"DD",X"7E",X"04",X"DD",X"6E",X"05",X"CD",X"00",X"2D",X"1A",X"E6",X"F8",X"FE",X"08",
		X"20",X"0B",X"DD",X"7E",X"02",X"FE",X"80",X"D8",X"3E",X"01",X"32",X"87",X"E5",X"7E",X"E6",X"FC",
		X"FE",X"18",X"20",X"17",X"DD",X"7E",X"15",X"FE",X"03",X"20",X"10",X"DD",X"35",X"15",X"DD",X"36",
		X"0A",X"28",X"CD",X"76",X"1A",X"D0",X"DD",X"36",X"0A",X"0C",X"C9",X"CD",X"C1",X"1B",X"DD",X"7E",
		X"04",X"DD",X"6E",X"03",X"CD",X"00",X"2D",X"1A",X"E6",X"F8",X"FE",X"10",X"20",X"29",X"15",X"1A",
		X"E6",X"F8",X"FE",X"10",X"28",X"21",X"DD",X"7E",X"14",X"FE",X"15",X"28",X"1A",X"DD",X"34",X"14",
		X"DD",X"46",X"0A",X"DD",X"4E",X"09",X"C5",X"DD",X"36",X"0A",X"20",X"CD",X"76",X"1A",X"C1",X"30",
		X"3F",X"DD",X"70",X"0A",X"DD",X"71",X"09",X"DD",X"7E",X"02",X"C6",X"15",X"DD",X"77",X"02",X"30",
		X"0D",X"DD",X"34",X"03",X"3A",X"87",X"E5",X"B7",X"28",X"04",X"AF",X"DD",X"77",X"02",X"DD",X"6E",
		X"02",X"DD",X"66",X"03",X"29",X"7C",X"3C",X"1F",X"DD",X"77",X"05",X"29",X"29",X"7C",X"DD",X"77",
		X"06",X"CD",X"39",X"1B",X"CD",X"7A",X"1B",X"06",X"08",X"CD",X"2E",X"1A",X"DD",X"36",X"14",X"15",
		X"DD",X"7E",X"06",X"DD",X"6E",X"07",X"C3",X"D3",X"2E",X"DD",X"6E",X"06",X"DD",X"7E",X"07",X"CD",
		X"EF",X"2D",X"D8",X"AF",X"32",X"87",X"E5",X"DD",X"7E",X"04",X"B7",X"28",X"16",X"DD",X"7E",X"04",
		X"DD",X"6E",X"05",X"CD",X"00",X"2D",X"2B",X"2B",X"2B",X"2B",X"06",X"F8",X"0E",X"08",X"CD",X"8D",
		X"2E",X"20",X"0C",X"DD",X"7E",X"00",X"3D",X"FE",X"7F",X"D0",X"3E",X"01",X"32",X"87",X"E5",X"3E",
		X"01",X"DD",X"77",X"0B",X"CD",X"EE",X"1B",X"CD",X"4C",X"18",X"DD",X"7E",X"00",X"D6",X"0E",X"DD",
		X"77",X"00",X"30",X"0F",X"3A",X"87",X"E5",X"B7",X"28",X"06",X"AF",X"DD",X"77",X"00",X"18",X"03",
		X"DD",X"35",X"01",X"18",X"57",X"DD",X"6E",X"06",X"DD",X"7E",X"07",X"CD",X"31",X"2E",X"D8",X"AF",
		X"32",X"87",X"E5",X"DD",X"7E",X"04",X"FE",X"17",X"30",X"16",X"DD",X"7E",X"04",X"DD",X"6E",X"05",
		X"CD",X"00",X"2D",X"23",X"23",X"23",X"23",X"06",X"F8",X"0E",X"08",X"CD",X"8D",X"2E",X"20",X"0B",
		X"DD",X"7E",X"00",X"FE",X"80",X"D8",X"3E",X"01",X"32",X"87",X"E5",X"AF",X"DD",X"77",X"0B",X"CD",
		X"EE",X"1B",X"CD",X"4C",X"18",X"DD",X"7E",X"00",X"C6",X"0E",X"DD",X"77",X"00",X"30",X"0D",X"DD",
		X"34",X"01",X"3A",X"87",X"E5",X"B7",X"28",X"AB",X"AF",X"DD",X"77",X"00",X"DD",X"6E",X"00",X"DD",
		X"66",X"01",X"29",X"7C",X"3C",X"1F",X"DD",X"77",X"04",X"29",X"29",X"7C",X"DD",X"77",X"07",X"CD",
		X"39",X"1B",X"CD",X"7A",X"1B",X"DD",X"6E",X"06",X"DD",X"7E",X"0B",X"B7",X"DD",X"7E",X"07",X"28",
		X"05",X"CD",X"B9",X"2E",X"18",X"03",X"CD",X"B5",X"2E",X"DD",X"7E",X"04",X"DD",X"6E",X"05",X"CD",
		X"00",X"2D",X"E6",X"FC",X"FE",X"18",X"20",X"19",X"DD",X"7E",X"15",X"B7",X"20",X"0B",X"DD",X"34",
		X"15",X"DD",X"36",X"0A",X"24",X"CD",X"76",X"1A",X"D0",X"DD",X"36",X"15",X"03",X"06",X"04",X"18",
		X"18",X"DD",X"7E",X"15",X"FE",X"03",X"20",X"0B",X"DD",X"35",X"15",X"DD",X"36",X"0A",X"28",X"CD",
		X"76",X"1A",X"D0",X"DD",X"36",X"15",X"00",X"06",X"00",X"C3",X"2E",X"1A",X"3A",X"6D",X"E5",X"B7",
		X"20",X"07",X"3A",X"FB",X"E4",X"B7",X"C8",X"18",X"05",X"3A",X"6F",X"E5",X"B7",X"C8",X"DD",X"7E",
		X"04",X"DD",X"6E",X"05",X"CD",X"00",X"2D",X"E6",X"FC",X"FE",X"18",X"C0",X"F1",X"DD",X"6E",X"06",
		X"DD",X"7E",X"0B",X"B7",X"DD",X"7E",X"07",X"28",X"05",X"CD",X"B9",X"2E",X"18",X"03",X"CD",X"B5",
		X"2E",X"DD",X"7E",X"0A",X"E6",X"FC",X"FE",X"2C",X"28",X"04",X"DD",X"36",X"09",X"01",X"DD",X"35",
		X"09",X"C0",X"DD",X"34",X"0A",X"DD",X"7E",X"0A",X"E6",X"FC",X"FE",X"2C",X"28",X"04",X"DD",X"36",
		X"0A",X"2C",X"CD",X"19",X"1B",X"21",X"20",X"4C",X"09",X"7E",X"DD",X"77",X"09",X"21",X"D0",X"4D",
		X"09",X"7E",X"B7",X"C8",X"87",X"87",X"87",X"87",X"5F",X"3A",X"87",X"E5",X"57",X"DD",X"7E",X"00",
		X"DD",X"CB",X"0B",X"46",X"28",X"0F",X"93",X"30",X"0A",X"CB",X"42",X"28",X"03",X"AF",X"18",X"03",
		X"DD",X"35",X"01",X"18",X"0B",X"83",X"30",X"08",X"DD",X"34",X"01",X"CB",X"42",X"28",X"01",X"AF",
		X"DD",X"77",X"00",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"29",X"7C",X"3C",X"1F",X"DD",X"77",X"04",
		X"29",X"29",X"7C",X"DD",X"77",X"07",X"C9",X"DD",X"7E",X"0F",X"FE",X"FF",X"C8",X"E6",X"03",X"CA",
		X"A6",X"19",X"3D",X"CA",X"EA",X"19",X"3D",X"28",X"59",X"DD",X"7E",X"0C",X"B7",X"28",X"0F",X"DD",
		X"7E",X"04",X"DD",X"6E",X"05",X"CD",X"00",X"2D",X"E6",X"F8",X"FE",X"08",X"37",X"C8",X"DD",X"CB",
		X"0F",X"6E",X"20",X"0A",X"DD",X"7E",X"06",X"DD",X"6E",X"07",X"CD",X"A2",X"2D",X"D8",X"DD",X"46",
		X"0F",X"CB",X"78",X"20",X"20",X"DD",X"7E",X"02",X"D6",X"20",X"DD",X"77",X"02",X"30",X"03",X"DD",
		X"35",X"03",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"29",X"7C",X"3C",X"1F",X"DD",X"77",X"05",X"29",
		X"29",X"7C",X"DD",X"77",X"06",X"DD",X"7E",X"06",X"DD",X"6E",X"07",X"CB",X"70",X"CC",X"D3",X"2E",
		X"B7",X"C9",X"DD",X"CB",X"0F",X"6E",X"20",X"0A",X"DD",X"7E",X"06",X"DD",X"6E",X"07",X"CD",X"9E",
		X"2D",X"D8",X"DD",X"46",X"0F",X"CB",X"78",X"20",X"20",X"DD",X"7E",X"02",X"C6",X"20",X"DD",X"77",
		X"02",X"30",X"03",X"DD",X"34",X"03",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"29",X"7C",X"3C",X"1F",
		X"DD",X"77",X"05",X"29",X"29",X"7C",X"DD",X"77",X"06",X"DD",X"7E",X"06",X"DD",X"6E",X"07",X"CB",
		X"70",X"CC",X"D3",X"2E",X"B7",X"C9",X"DD",X"CB",X"0F",X"6E",X"20",X"0A",X"DD",X"6E",X"06",X"DD",
		X"7E",X"07",X"CD",X"31",X"2E",X"D8",X"DD",X"46",X"0F",X"CB",X"78",X"20",X"20",X"DD",X"7E",X"00",
		X"C6",X"10",X"DD",X"77",X"00",X"30",X"03",X"DD",X"34",X"01",X"DD",X"6E",X"00",X"DD",X"66",X"01",
		X"29",X"7C",X"3C",X"1F",X"DD",X"77",X"04",X"29",X"29",X"7C",X"DD",X"77",X"07",X"DD",X"6E",X"06",
		X"DD",X"7E",X"07",X"CB",X"70",X"CC",X"B5",X"2E",X"B7",X"C9",X"DD",X"CB",X"0F",X"6E",X"20",X"0A",
		X"DD",X"6E",X"06",X"DD",X"7E",X"07",X"CD",X"EF",X"2D",X"D8",X"DD",X"46",X"0F",X"CB",X"78",X"20",
		X"20",X"DD",X"7E",X"00",X"D6",X"10",X"DD",X"77",X"00",X"30",X"03",X"DD",X"35",X"01",X"DD",X"6E",
		X"00",X"DD",X"66",X"01",X"29",X"7C",X"3C",X"1F",X"DD",X"77",X"04",X"29",X"29",X"7C",X"DD",X"77",
		X"07",X"DD",X"6E",X"06",X"DD",X"7E",X"07",X"CB",X"70",X"CC",X"B9",X"2E",X"B7",X"C9",X"DD",X"35",
		X"09",X"C0",X"DD",X"36",X"09",X"06",X"DD",X"34",X"0A",X"DD",X"7E",X"0A",X"FE",X"03",X"20",X"12",
		X"3A",X"CD",X"E5",X"5F",X"16",X"00",X"21",X"5D",X"1A",X"19",X"7E",X"B7",X"28",X"04",X"DD",X"70",
		X"0A",X"C9",X"DD",X"7E",X"0A",X"E6",X"FC",X"B8",X"C8",X"DD",X"70",X"0A",X"C9",X"00",X"00",X"01",
		X"01",X"00",X"00",X"01",X"00",X"00",X"DD",X"35",X"09",X"C0",X"DD",X"34",X"0A",X"DD",X"7E",X"0A",
		X"E6",X"FC",X"B8",X"C2",X"0D",X"1B",X"DD",X"36",X"10",X"00",X"CD",X"19",X"1B",X"21",X"20",X"4C",
		X"09",X"7E",X"DD",X"77",X"09",X"B7",X"CA",X"0D",X"1B",X"21",X"F8",X"4C",X"09",X"7E",X"57",X"E6",
		X"03",X"20",X"07",X"DD",X"CB",X"0B",X"46",X"28",X"01",X"14",X"DD",X"72",X"0F",X"21",X"D0",X"4D",
		X"09",X"7E",X"B7",X"28",X"30",X"87",X"87",X"87",X"87",X"16",X"00",X"DD",X"CB",X"0B",X"46",X"28",
		X"03",X"ED",X"44",X"15",X"5F",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"19",X"DD",X"75",X"00",X"DD",
		X"74",X"01",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"29",X"7C",X"3C",X"1F",X"DD",X"77",X"04",X"29",
		X"29",X"7C",X"DD",X"77",X"07",X"21",X"A8",X"4E",X"09",X"7E",X"B7",X"28",X"2F",X"56",X"1E",X"00",
		X"CB",X"2A",X"CB",X"1B",X"CB",X"2A",X"CB",X"1B",X"CB",X"2A",X"CB",X"1B",X"DD",X"6E",X"02",X"DD",
		X"66",X"03",X"19",X"DD",X"75",X"02",X"DD",X"74",X"03",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"29",
		X"7C",X"3C",X"1F",X"DD",X"77",X"05",X"29",X"29",X"7C",X"DD",X"77",X"06",X"C9",X"DD",X"35",X"0A",
		X"DD",X"34",X"09",X"DD",X"36",X"0F",X"FF",X"37",X"C9",X"3A",X"6D",X"E5",X"B7",X"28",X"08",X"3A",
		X"CD",X"E5",X"E6",X"07",X"3C",X"18",X"03",X"3A",X"CD",X"E5",X"47",X"87",X"80",X"87",X"87",X"87",
		X"DD",X"86",X"0A",X"D6",X"18",X"4F",X"06",X"00",X"C9",X"3A",X"6D",X"E5",X"B7",X"C0",X"DD",X"7E",
		X"00",X"FE",X"80",X"38",X"02",X"ED",X"44",X"FE",X"0E",X"D0",X"DD",X"7E",X"02",X"FE",X"80",X"38",
		X"02",X"ED",X"44",X"FE",X"15",X"D0",X"DD",X"7E",X"04",X"DD",X"6E",X"05",X"CD",X"00",X"2D",X"15",
		X"1A",X"E6",X"FC",X"FE",X"70",X"C0",X"DD",X"7E",X"0D",X"B7",X"C0",X"3A",X"68",X"E5",X"C6",X"04",
		X"87",X"87",X"87",X"DD",X"77",X"0D",X"CD",X"5C",X"2F",X"C9",X"DD",X"7E",X"0D",X"B7",X"C8",X"DD",
		X"7E",X"0F",X"FE",X"02",X"D0",X"DD",X"7E",X"0A",X"FE",X"04",X"38",X"03",X"FE",X"08",X"D8",X"DD",
		X"7E",X"04",X"DD",X"6E",X"05",X"CD",X"00",X"2D",X"15",X"06",X"FC",X"0E",X"00",X"CD",X"7F",X"2E",
		X"C0",X"DD",X"35",X"0D",X"C0",X"DD",X"7E",X"0F",X"FE",X"00",X"DD",X"7E",X"00",X"20",X"06",X"FE",
		X"80",X"30",X"0A",X"18",X"04",X"FE",X"80",X"38",X"04",X"CD",X"0E",X"2F",X"C9",X"DD",X"34",X"0D",
		X"C9",X"DD",X"7E",X"00",X"FE",X"80",X"30",X"07",X"D6",X"0E",X"30",X"01",X"AF",X"18",X"08",X"C6",
		X"0E",X"30",X"04",X"DD",X"34",X"01",X"AF",X"DD",X"77",X"00",X"6F",X"DD",X"66",X"01",X"29",X"7C",
		X"3C",X"1F",X"DD",X"77",X"04",X"29",X"29",X"7C",X"DD",X"77",X"07",X"C3",X"39",X"1B",X"DD",X"7E",
		X"02",X"FE",X"80",X"30",X"07",X"D6",X"15",X"30",X"01",X"AF",X"18",X"08",X"C6",X"15",X"30",X"04",
		X"DD",X"34",X"03",X"AF",X"DD",X"77",X"02",X"6F",X"DD",X"66",X"03",X"29",X"7C",X"3C",X"1F",X"DD",
		X"77",X"05",X"29",X"29",X"7C",X"DD",X"77",X"06",X"C3",X"39",X"1B",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"3A",X"E9",X"E4",X"32",X"EA",X"E4",X"DD",X"21",X"58",X"E4",X"FD",X"21",X"EB",X"E4",X"DD",X"7E",
		X"10",X"B7",X"28",X"1C",X"DD",X"6E",X"04",X"DD",X"66",X"05",X"22",X"EF",X"E4",X"DD",X"7E",X"07",
		X"32",X"F2",X"E4",X"CD",X"FD",X"1D",X"47",X"DD",X"7E",X"10",X"B7",X"28",X"03",X"DD",X"70",X"0F",
		X"11",X"18",X"00",X"DD",X"19",X"21",X"EA",X"E4",X"35",X"20",X"D3",X"3A",X"E9",X"E4",X"32",X"EA",
		X"E4",X"DD",X"21",X"58",X"E4",X"DD",X"7E",X"04",X"DD",X"6E",X"05",X"2C",X"2C",X"CD",X"D5",X"62",
		X"7E",X"E6",X"0D",X"FE",X"0D",X"28",X"0A",X"21",X"01",X"E5",X"7E",X"FE",X"39",X"D0",X"36",X"00",
		X"C9",X"11",X"18",X"00",X"DD",X"19",X"21",X"EA",X"E4",X"35",X"20",X"D9",X"21",X"01",X"E5",X"7E",
		X"FE",X"38",X"30",X"02",X"34",X"C9",X"C0",X"34",X"3E",X"00",X"32",X"9D",X"E5",X"21",X"B5",X"E5",
		X"7E",X"BE",X"28",X"FD",X"CD",X"8D",X"32",X"21",X"29",X"D7",X"36",X"05",X"2B",X"36",X"00",X"11",
		X"2A",X"D7",X"01",X"2E",X"00",X"ED",X"B0",X"21",X"A9",X"D7",X"36",X"05",X"2B",X"36",X"00",X"11",
		X"AA",X"D7",X"01",X"2E",X"00",X"ED",X"B0",X"21",X"29",X"D8",X"36",X"05",X"2B",X"36",X"00",X"11",
		X"2A",X"D8",X"01",X"2E",X"00",X"ED",X"B0",X"0E",X"47",X"21",X"AA",X"D7",X"11",X"E5",X"1D",X"CD",
		X"2D",X"30",X"3E",X"1F",X"CD",X"42",X"31",X"0E",X"01",X"CD",X"CF",X"2F",X"CD",X"03",X"32",X"3E",
		X"01",X"32",X"89",X"E5",X"CD",X"89",X"06",X"CD",X"B9",X"32",X"3E",X"26",X"CD",X"42",X"31",X"3E",
		X"02",X"32",X"9D",X"E5",X"C9",X"41",X"4C",X"4C",X"20",X"45",X"4E",X"45",X"4D",X"49",X"45",X"53",
		X"20",X"41",X"52",X"45",X"20",X"53",X"45",X"41",X"4C",X"45",X"44",X"2E",X"00",X"3A",X"45",X"E4",
		X"FD",X"BE",X"05",X"C2",X"B9",X"1E",X"FD",X"46",X"04",X"FD",X"7E",X"07",X"21",X"47",X"E4",X"BE",
		X"38",X"05",X"20",X"54",X"3E",X"FF",X"C9",X"3A",X"44",X"E4",X"B8",X"20",X"03",X"3E",X"00",X"C9",
		X"04",X"78",X"FD",X"6E",X"05",X"CD",X"00",X"2D",X"E6",X"FC",X"FE",X"18",X"28",X"E9",X"7E",X"E6",
		X"F8",X"FE",X"10",X"28",X"E2",X"24",X"7E",X"25",X"E6",X"F8",X"FE",X"10",X"28",X"D9",X"FD",X"7E",
		X"05",X"FE",X"1D",X"30",X"D2",X"7E",X"E6",X"F8",X"FE",X"08",X"28",X"6D",X"24",X"7E",X"E6",X"F8",
		X"FE",X"08",X"28",X"65",X"1A",X"E6",X"F8",X"FE",X"10",X"28",X"BC",X"1A",X"FE",X"04",X"28",X"B7",
		X"E6",X"F8",X"FE",X"08",X"28",X"B1",X"18",X"51",X"3A",X"44",X"E4",X"B8",X"20",X"03",X"3E",X"01",
		X"C9",X"05",X"78",X"FD",X"6E",X"05",X"CD",X"00",X"2D",X"E6",X"FC",X"FE",X"18",X"28",X"E9",X"7E",
		X"E6",X"F8",X"FE",X"10",X"28",X"E2",X"24",X"7E",X"25",X"E6",X"F8",X"FE",X"10",X"28",X"D9",X"FD",
		X"7E",X"05",X"FE",X"1D",X"30",X"D2",X"7E",X"E6",X"F8",X"FE",X"08",X"28",X"1C",X"24",X"7E",X"E6",
		X"F8",X"FE",X"08",X"28",X"14",X"1A",X"E6",X"F8",X"FE",X"10",X"28",X"BC",X"1A",X"FE",X"04",X"28",
		X"B7",X"E6",X"F8",X"FE",X"08",X"28",X"B1",X"18",X"00",X"3E",X"FF",X"32",X"ED",X"E4",X"32",X"EE",
		X"E4",X"FD",X"7E",X"04",X"32",X"EB",X"E4",X"32",X"EC",X"E4",X"CD",X"E0",X"1E",X"CD",X"2B",X"1F",
		X"CD",X"77",X"1F",X"CD",X"96",X"1F",X"CD",X"B9",X"1F",X"CD",X"F1",X"1F",X"3A",X"ED",X"E4",X"C9",
		X"3A",X"EB",X"E4",X"B7",X"28",X"44",X"3D",X"FD",X"6E",X"05",X"CD",X"00",X"2D",X"06",X"F8",X"0E",
		X"08",X"CD",X"8D",X"2E",X"C8",X"06",X"F8",X"0E",X"10",X"CD",X"8D",X"2E",X"28",X"25",X"7E",X"E6",
		X"FC",X"FE",X"18",X"28",X"1E",X"FD",X"7E",X"05",X"FE",X"1D",X"30",X"17",X"1A",X"E6",X"F8",X"FE",
		X"10",X"28",X"10",X"1A",X"FE",X"04",X"28",X"0B",X"E6",X"F8",X"FE",X"08",X"28",X"05",X"21",X"EB",
		X"E4",X"35",X"C9",X"21",X"EB",X"E4",X"35",X"7E",X"18",X"B9",X"C9",X"3A",X"EC",X"E4",X"FE",X"17",
		X"30",X"44",X"3C",X"FD",X"6E",X"05",X"CD",X"00",X"2D",X"06",X"F8",X"0E",X"08",X"CD",X"8D",X"2E",
		X"C8",X"06",X"F8",X"0E",X"10",X"CD",X"8D",X"2E",X"28",X"25",X"7E",X"E6",X"FC",X"FE",X"18",X"28",
		X"1E",X"FD",X"7E",X"05",X"FE",X"1D",X"30",X"17",X"1A",X"E6",X"F8",X"FE",X"10",X"28",X"10",X"1A",
		X"FE",X"04",X"28",X"0B",X"E6",X"F8",X"FE",X"08",X"28",X"05",X"21",X"EC",X"E4",X"34",X"C9",X"21",
		X"EC",X"E4",X"34",X"7E",X"18",X"B8",X"C9",X"FD",X"7E",X"04",X"CD",X"2A",X"20",X"FD",X"BE",X"05",
		X"C8",X"32",X"F3",X"E4",X"FD",X"4E",X"04",X"CD",X"3D",X"21",X"21",X"EE",X"E4",X"BE",X"D0",X"77",
		X"3E",X"02",X"32",X"ED",X"E4",X"C9",X"FD",X"7E",X"04",X"CD",X"B6",X"20",X"FD",X"BE",X"05",X"C8",
		X"FD",X"4E",X"04",X"32",X"F4",X"E4",X"CD",X"3D",X"21",X"21",X"EE",X"E4",X"47",X"78",X"18",X"00",
		X"BE",X"D0",X"77",X"3E",X"03",X"32",X"ED",X"E4",X"C9",X"21",X"EB",X"E4",X"7E",X"FD",X"BE",X"04",
		X"30",X"15",X"CD",X"2A",X"20",X"CD",X"D8",X"1F",X"3A",X"EB",X"E4",X"CD",X"B6",X"20",X"CD",X"D8",
		X"1F",X"21",X"EB",X"E4",X"34",X"18",X"E5",X"C9",X"FD",X"BE",X"05",X"C8",X"21",X"EB",X"E4",X"4E",
		X"CD",X"3D",X"21",X"21",X"EE",X"E4",X"BE",X"D0",X"32",X"EE",X"E4",X"3E",X"01",X"32",X"ED",X"E4",
		X"C9",X"21",X"EC",X"E4",X"FD",X"7E",X"04",X"BE",X"30",X"16",X"7E",X"CD",X"2A",X"20",X"CD",X"11",
		X"20",X"3A",X"EC",X"E4",X"CD",X"B6",X"20",X"CD",X"11",X"20",X"21",X"EC",X"E4",X"35",X"18",X"E4",
		X"C9",X"FD",X"BE",X"05",X"C8",X"21",X"EC",X"E4",X"4E",X"CD",X"3D",X"21",X"21",X"EE",X"E4",X"BE",
		X"D0",X"32",X"EE",X"E4",X"3E",X"00",X"32",X"ED",X"E4",X"C9",X"47",X"FD",X"4E",X"05",X"79",X"FE",
		X"1D",X"30",X"52",X"61",X"78",X"07",X"07",X"07",X"CB",X"3C",X"1F",X"6F",X"11",X"10",X"D0",X"19",
		X"E5",X"11",X"80",X"01",X"19",X"D1",X"EB",X"1A",X"FE",X"04",X"28",X"3A",X"E6",X"F8",X"FE",X"08",
		X"28",X"34",X"0C",X"1A",X"24",X"24",X"15",X"EB",X"E6",X"FC",X"FE",X"00",X"28",X"25",X"3A",X"44",
		X"E4",X"B8",X"30",X"0D",X"2D",X"2D",X"2D",X"2D",X"1D",X"1D",X"1D",X"1D",X"CD",X"88",X"20",X"18",
		X"12",X"20",X"05",X"CD",X"AD",X"20",X"18",X"0B",X"2C",X"2C",X"2C",X"2C",X"1C",X"1C",X"1C",X"1C",
		X"CD",X"88",X"20",X"18",X"A9",X"C9",X"79",X"C9",X"7E",X"E6",X"FC",X"FE",X"18",X"28",X"1E",X"7E",
		X"E6",X"F8",X"FE",X"08",X"C8",X"24",X"7E",X"E6",X"F8",X"FE",X"08",X"C8",X"1A",X"E6",X"F8",X"FE",
		X"10",X"28",X"0A",X"1A",X"FE",X"04",X"28",X"05",X"E6",X"F8",X"FE",X"08",X"C0",X"21",X"45",X"E4",
		X"79",X"BE",X"D8",X"F1",X"79",X"C9",X"47",X"FD",X"4E",X"05",X"79",X"FE",X"01",X"28",X"50",X"61",
		X"78",X"07",X"07",X"07",X"CB",X"3C",X"1F",X"6F",X"11",X"10",X"D0",X"19",X"E5",X"11",X"80",X"01",
		X"19",X"D1",X"EB",X"7E",X"E6",X"F8",X"FE",X"10",X"28",X"09",X"24",X"7E",X"25",X"E6",X"F8",X"FE",
		X"10",X"79",X"C0",X"0D",X"15",X"15",X"24",X"EB",X"3A",X"44",X"E4",X"B8",X"30",X"0D",X"2D",X"2D",
		X"2D",X"2D",X"1D",X"1D",X"1D",X"1D",X"CD",X"10",X"21",X"18",X"12",X"20",X"05",X"CD",X"35",X"21",
		X"18",X"0B",X"2C",X"2C",X"2C",X"2C",X"1C",X"1C",X"1C",X"1C",X"CD",X"10",X"21",X"18",X"AB",X"C9",
		X"7E",X"E6",X"FC",X"FE",X"18",X"28",X"1E",X"7E",X"E6",X"F8",X"FE",X"08",X"C8",X"24",X"7E",X"E6",
		X"F8",X"FE",X"08",X"C8",X"1A",X"E6",X"F8",X"FE",X"10",X"28",X"0A",X"1A",X"FE",X"04",X"28",X"05",
		X"E6",X"F8",X"FE",X"08",X"C0",X"3A",X"45",X"E4",X"B9",X"D8",X"F1",X"79",X"C9",X"47",X"78",X"18",
		X"14",X"2A",X"44",X"E4",X"94",X"30",X"02",X"ED",X"44",X"87",X"87",X"87",X"47",X"79",X"95",X"30",
		X"02",X"ED",X"44",X"80",X"C9",X"21",X"45",X"E4",X"BE",X"20",X"08",X"79",X"FD",X"96",X"04",X"D0",
		X"ED",X"44",X"C9",X"78",X"96",X"30",X"05",X"ED",X"44",X"C6",X"64",X"C9",X"C6",X"C8",X"C9",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"21",X"0E",X"E5",X"7E",X"B7",X"28",X"02",X"35",X"C9",X"34",X"CD",X"BE",X"24",X"21",X"68",X"E5",
		X"35",X"20",X"02",X"36",X"17",X"DD",X"21",X"18",X"E5",X"3E",X"14",X"32",X"88",X"E5",X"DD",X"7E",
		X"00",X"B7",X"28",X"39",X"DD",X"35",X"00",X"20",X"06",X"DD",X"36",X"01",X"00",X"18",X"2E",X"DD",
		X"7E",X"00",X"FE",X"10",X"20",X"04",X"DD",X"36",X"01",X"F4",X"30",X"21",X"FE",X"0F",X"20",X"12",
		X"DD",X"7E",X"02",X"DD",X"6E",X"03",X"CD",X"00",X"2D",X"EB",X"CD",X"19",X"30",X"CD",X"69",X"24",
		X"18",X"0B",X"CB",X"3F",X"CB",X"3F",X"47",X"3E",X"F7",X"90",X"DD",X"77",X"01",X"01",X"04",X"00",
		X"DD",X"09",X"21",X"88",X"E5",X"35",X"20",X"B6",X"C9",X"3A",X"44",X"E4",X"DD",X"BE",X"02",X"20",
		X"17",X"DD",X"7E",X"03",X"21",X"45",X"E4",X"96",X"38",X"0E",X"FE",X"03",X"30",X"0A",X"3E",X"00",
		X"32",X"48",X"E4",X"AF",X"32",X"50",X"E4",X"C9",X"FD",X"21",X"58",X"E4",X"3A",X"E9",X"E4",X"32",
		X"89",X"E5",X"FD",X"7E",X"04",X"DD",X"BE",X"02",X"20",X"18",X"DD",X"7E",X"03",X"FD",X"96",X"05",
		X"38",X"10",X"FE",X"03",X"30",X"0C",X"FD",X"36",X"0C",X"FF",X"FD",X"36",X"09",X"2A",X"FD",X"36",
		X"0E",X"3C",X"11",X"18",X"00",X"FD",X"19",X"21",X"89",X"E5",X"35",X"20",X"D5",X"C9",X"3A",X"E9",
		X"E4",X"32",X"E8",X"E4",X"DD",X"21",X"58",X"E4",X"21",X"6D",X"E5",X"36",X"00",X"3A",X"02",X"E5",
		X"B7",X"28",X"08",X"3A",X"E8",X"E4",X"FE",X"01",X"20",X"01",X"34",X"DD",X"7E",X"0E",X"B7",X"28",
		X"5B",X"DD",X"35",X"09",X"20",X"25",X"3A",X"6D",X"E5",X"B7",X"28",X"0A",X"AF",X"32",X"02",X"E5",
		X"21",X"E9",X"E4",X"35",X"18",X"15",X"DD",X"36",X"09",X"03",X"DD",X"7E",X"0A",X"FE",X"FF",X"20",
		X"06",X"DD",X"36",X"0A",X"0C",X"18",X"04",X"DD",X"36",X"0A",X"FF",X"DD",X"35",X"0E",X"20",X"24",
		X"FD",X"21",X"40",X"E4",X"FD",X"7E",X"04",X"DD",X"BE",X"04",X"20",X"10",X"FD",X"7E",X"05",X"FE",
		X"01",X"38",X"09",X"FE",X"04",X"30",X"05",X"DD",X"34",X"0E",X"18",X"10",X"DD",X"36",X"0C",X"00",
		X"DD",X"36",X"0A",X"0C",X"DD",X"7E",X"0E",X"FE",X"30",X"CC",X"48",X"25",X"11",X"18",X"00",X"DD",
		X"19",X"21",X"E8",X"E4",X"35",X"20",X"81",X"C9",X"3A",X"6D",X"E5",X"B7",X"20",X"0D",X"3E",X"01",
		X"32",X"FF",X"E4",X"01",X"00",X"01",X"CD",X"DB",X"2F",X"18",X"13",X"DD",X"7E",X"04",X"DD",X"6E",
		X"05",X"CD",X"00",X"2D",X"15",X"15",X"1A",X"E6",X"FC",X"FE",X"60",X"CC",X"83",X"2F",X"3E",X"04",
		X"CD",X"42",X"31",X"DD",X"7E",X"0D",X"B7",X"28",X"04",X"21",X"FC",X"E4",X"35",X"DD",X"36",X"0A",
		X"FF",X"11",X"10",X"D1",X"3A",X"68",X"E5",X"87",X"87",X"6F",X"26",X"00",X"19",X"EB",X"06",X"F8",
		X"0E",X"08",X"CD",X"71",X"2E",X"EB",X"20",X"0A",X"21",X"68",X"E5",X"35",X"20",X"02",X"36",X"17",
		X"18",X"E2",X"3A",X"68",X"E5",X"DD",X"77",X"01",X"DD",X"77",X"04",X"87",X"87",X"87",X"DD",X"77",
		X"07",X"AF",X"DD",X"77",X"00",X"DD",X"77",X"02",X"DD",X"77",X"0D",X"3C",X"DD",X"77",X"03",X"DD",
		X"77",X"05",X"DD",X"36",X"06",X"08",X"21",X"68",X"E5",X"35",X"20",X"02",X"36",X"17",X"C9",X"3E",
		X"01",X"32",X"A7",X"E5",X"21",X"22",X"D2",X"CD",X"A1",X"29",X"3E",X"0E",X"CD",X"3E",X"30",X"21",
		X"DE",X"D3",X"11",X"E9",X"26",X"CD",X"2D",X"30",X"21",X"23",X"D2",X"16",X"CB",X"CD",X"DF",X"29",
		X"3E",X"1C",X"CD",X"3E",X"30",X"21",X"23",X"D2",X"16",X"CC",X"CD",X"DF",X"29",X"3E",X"1C",X"CD",
		X"3E",X"30",X"21",X"23",X"D2",X"16",X"CD",X"CD",X"DF",X"29",X"3E",X"1C",X"CD",X"3E",X"30",X"7A",
		X"32",X"6B",X"E5",X"21",X"40",X"E4",X"11",X"41",X"E4",X"01",X"28",X"01",X"36",X"00",X"ED",X"B0",
		X"3E",X"01",X"32",X"CD",X"E5",X"32",X"4B",X"E4",X"32",X"49",X"E4",X"3E",X"16",X"32",X"41",X"E4",
		X"3E",X"0C",X"32",X"43",X"E4",X"3E",X"00",X"32",X"4A",X"E4",X"32",X"46",X"E4",X"3E",X"1E",X"32",
		X"53",X"E4",X"16",X"18",X"1E",X"0C",X"3E",X"01",X"DD",X"21",X"58",X"E4",X"06",X"05",X"DD",X"77",
		X"0B",X"DD",X"77",X"09",X"DD",X"72",X"01",X"DD",X"73",X"03",X"DD",X"36",X"0A",X"00",X"DD",X"36",
		X"06",X"00",X"C5",X"01",X"18",X"00",X"DD",X"09",X"C1",X"14",X"10",X"E2",X"21",X"80",X"00",X"DB",
		X"04",X"CB",X"47",X"20",X"02",X"2D",X"2D",X"22",X"E3",X"E5",X"CD",X"D7",X"63",X"3E",X"05",X"32",
		X"E9",X"E4",X"3E",X"03",X"32",X"6A",X"E5",X"3E",X"01",X"32",X"9D",X"E5",X"3E",X"30",X"32",X"89",
		X"E5",X"21",X"6B",X"E5",X"34",X"7E",X"FE",X"D0",X"38",X"02",X"36",X"CD",X"56",X"21",X"23",X"D2",
		X"CD",X"DF",X"29",X"3E",X"08",X"CD",X"3E",X"30",X"21",X"89",X"E5",X"35",X"20",X"E3",X"3E",X"00",
		X"32",X"9D",X"E5",X"3E",X"00",X"32",X"6A",X"E5",X"CD",X"00",X"65",X"3A",X"DE",X"E5",X"CD",X"00",
		X"5C",X"06",X"03",X"21",X"DE",X"E5",X"7E",X"B7",X"28",X"05",X"36",X"00",X"04",X"18",X"01",X"34",
		X"78",X"32",X"8E",X"E5",X"AF",X"32",X"B8",X"E5",X"32",X"8F",X"E5",X"67",X"6F",X"22",X"91",X"E5",
		X"22",X"92",X"E5",X"CD",X"5E",X"5F",X"C3",X"97",X"5D",X"06",X"54",X"4D",X"00",X"3E",X"13",X"CD",
		X"42",X"31",X"3E",X"01",X"32",X"A9",X"E5",X"CD",X"5E",X"5F",X"21",X"00",X"52",X"CD",X"51",X"64",
		X"21",X"C0",X"D0",X"DD",X"21",X"BE",X"D0",X"0E",X"1F",X"06",X"18",X"7E",X"DD",X"77",X"00",X"2C",
		X"7E",X"EE",X"20",X"DD",X"77",X"01",X"2C",X"DD",X"2B",X"DD",X"2B",X"10",X"EE",X"11",X"50",X"00",
		X"19",X"11",X"B0",X"00",X"DD",X"19",X"0D",X"20",X"E0",X"21",X"24",X"E0",X"11",X"23",X"E0",X"0E",
		X"1F",X"06",X"0C",X"7E",X"07",X"07",X"07",X"07",X"12",X"23",X"1B",X"10",X"F6",X"C5",X"01",X"0C",
		X"00",X"09",X"EB",X"01",X"24",X"00",X"09",X"EB",X"C1",X"0D",X"20",X"E5",X"FD",X"21",X"39",X"54",
		X"CD",X"F0",X"29",X"3E",X"14",X"CD",X"42",X"31",X"3E",X"01",X"32",X"A6",X"E5",X"CD",X"43",X"5F",
		X"3E",X"24",X"CD",X"42",X"31",X"21",X"40",X"E4",X"11",X"41",X"E4",X"01",X"28",X"01",X"36",X"00",
		X"ED",X"B0",X"21",X"CD",X"E5",X"34",X"3E",X"01",X"32",X"4B",X"E4",X"32",X"49",X"E4",X"3E",X"06",
		X"32",X"44",X"E4",X"3E",X"10",X"32",X"41",X"E4",X"3E",X"1D",X"32",X"43",X"E4",X"3E",X"00",X"32",
		X"4A",X"E4",X"32",X"46",X"E4",X"16",X"12",X"1E",X"1F",X"3E",X"01",X"0E",X"05",X"DD",X"21",X"58",
		X"E4",X"06",X"04",X"DD",X"77",X"0B",X"DD",X"77",X"09",X"DD",X"71",X"04",X"DD",X"72",X"01",X"DD",
		X"73",X"03",X"DD",X"36",X"0A",X"00",X"DD",X"36",X"06",X"00",X"C5",X"01",X"18",X"00",X"DD",X"09",
		X"C1",X"14",X"1C",X"10",X"DE",X"CD",X"D7",X"63",X"3E",X"04",X"32",X"E9",X"E4",X"3E",X"02",X"32",
		X"6A",X"E5",X"3E",X"01",X"32",X"9D",X"E5",X"3E",X"A8",X"CD",X"3E",X"30",X"3E",X"03",X"CD",X"42",
		X"31",X"0E",X"30",X"DD",X"21",X"00",X"E3",X"06",X"0B",X"DD",X"34",X"06",X"DD",X"35",X"0E",X"11",
		X"10",X"00",X"DD",X"19",X"10",X"F3",X"3E",X"01",X"CD",X"3E",X"30",X"0D",X"20",X"E5",X"21",X"B6",
		X"D5",X"CD",X"9A",X"31",X"21",X"B8",X"D6",X"CD",X"85",X"31",X"21",X"3C",X"D8",X"11",X"2D",X"28",
		X"CD",X"2D",X"30",X"3E",X"70",X"CD",X"3E",X"30",X"3E",X"00",X"32",X"9D",X"E5",X"3E",X"00",X"32",
		X"6A",X"E5",X"3E",X"13",X"CD",X"42",X"31",X"CD",X"5E",X"5F",X"C3",X"97",X"5D",X"06",X"52",X"45",
		X"41",X"44",X"59",X"00",X"3E",X"13",X"CD",X"42",X"31",X"3E",X"01",X"32",X"A9",X"E5",X"CD",X"5E",
		X"5F",X"21",X"00",X"E3",X"11",X"01",X"E3",X"01",X"68",X"02",X"36",X"00",X"ED",X"B0",X"21",X"00",
		X"E0",X"11",X"01",X"E0",X"01",X"9F",X"02",X"36",X"00",X"ED",X"B0",X"23",X"13",X"01",X"5F",X"00",
		X"36",X"01",X"ED",X"B0",X"3E",X"0A",X"32",X"D8",X"E5",X"3E",X"00",X"32",X"A6",X"E5",X"3E",X"14",
		X"CD",X"42",X"31",X"CD",X"43",X"5F",X"3E",X"27",X"CD",X"42",X"31",X"06",X"00",X"0E",X"47",X"11",
		X"EF",X"28",X"3E",X"01",X"CD",X"3E",X"30",X"3E",X"2E",X"80",X"47",X"30",X"F5",X"1A",X"FE",X"01",
		X"20",X"07",X"13",X"1A",X"6F",X"13",X"1A",X"67",X"13",X"1A",X"77",X"FE",X"20",X"28",X"2E",X"3E",
		X"17",X"CD",X"42",X"31",X"1A",X"FE",X"32",X"20",X"24",X"AF",X"32",X"CD",X"E5",X"32",X"57",X"E4",
		X"3E",X"0B",X"32",X"41",X"E4",X"3E",X"0C",X"32",X"53",X"E4",X"32",X"4A",X"E4",X"3E",X"01",X"32",
		X"4B",X"E4",X"32",X"49",X"E4",X"32",X"6A",X"E5",X"3E",X"01",X"32",X"9D",X"E5",X"13",X"23",X"71",
		X"23",X"1A",X"B7",X"20",X"AD",X"3E",X"FF",X"CD",X"3E",X"30",X"3E",X"00",X"32",X"9D",X"E5",X"3E",
		X"00",X"32",X"6A",X"E5",X"3E",X"13",X"CD",X"42",X"31",X"CD",X"5E",X"5F",X"C3",X"FA",X"26",X"01",
		X"30",X"D3",X"43",X"4F",X"4E",X"47",X"52",X"41",X"54",X"55",X"4C",X"41",X"54",X"49",X"4F",X"4E",
		X"53",X"21",X"20",X"20",X"20",X"20",X"01",X"1E",X"D5",X"59",X"4F",X"55",X"20",X"20",X"48",X"41",
		X"56",X"45",X"20",X"20",X"44",X"4F",X"4E",X"45",X"20",X"20",X"49",X"54",X"20",X"20",X"56",X"45",
		X"52",X"59",X"20",X"20",X"57",X"45",X"4C",X"4C",X"2C",X"20",X"20",X"01",X"A8",X"D6",X"48",X"41",
		X"56",X"49",X"4E",X"47",X"20",X"20",X"50",X"41",X"53",X"53",X"45",X"44",X"20",X"20",X"54",X"48",
		X"52",X"4F",X"55",X"47",X"48",X"20",X"20",X"01",X"2A",X"D8",X"32",X"34",X"20",X"20",X"44",X"41",
		X"4E",X"47",X"45",X"52",X"4F",X"55",X"53",X"20",X"20",X"50",X"4C",X"41",X"43",X"45",X"53",X"2E",
		X"20",X"20",X"20",X"20",X"01",X"A0",X"D9",X"42",X"55",X"54",X"20",X"20",X"54",X"48",X"45",X"52",
		X"45",X"20",X"20",X"41",X"52",X"45",X"20",X"20",X"53",X"54",X"49",X"4C",X"4C",X"20",X"20",X"4F",
		X"54",X"48",X"45",X"52",X"20",X"20",X"01",X"28",X"DB",X"45",X"4E",X"45",X"4D",X"49",X"45",X"53",
		X"20",X"20",X"4F",X"4E",X"20",X"20",X"59",X"4F",X"55",X"52",X"20",X"20",X"57",X"41",X"59",X"2E",
		X"00",X"16",X"88",X"1E",X"04",X"06",X"1E",X"72",X"2C",X"2C",X"14",X"14",X"14",X"14",X"10",X"F7",
		X"7A",X"C6",X"89",X"57",X"01",X"44",X"00",X"09",X"1D",X"20",X"EA",X"C9",X"1E",X"04",X"7E",X"E6",
		X"F0",X"47",X"7A",X"E6",X"0F",X"B0",X"77",X"23",X"06",X"0E",X"72",X"23",X"10",X"FC",X"7E",X"E6",
		X"0F",X"47",X"7A",X"E6",X"F0",X"B0",X"77",X"01",X"09",X"00",X"09",X"1D",X"20",X"E0",X"C9",X"1E",
		X"04",X"06",X"1E",X"72",X"2C",X"2C",X"10",X"FB",X"01",X"44",X"00",X"09",X"1D",X"20",X"F2",X"C9",
		X"DD",X"21",X"00",X"E3",X"FD",X"7E",X"00",X"B7",X"C8",X"DD",X"77",X"04",X"DD",X"77",X"0C",X"FD",
		X"7E",X"01",X"47",X"E6",X"1F",X"DD",X"77",X"00",X"DD",X"77",X"08",X"78",X"E6",X"C0",X"DD",X"77",
		X"05",X"EE",X"40",X"DD",X"77",X"0D",X"FD",X"5E",X"02",X"16",X"00",X"2A",X"E3",X"E5",X"19",X"DD",
		X"75",X"02",X"DD",X"75",X"0A",X"DD",X"74",X"03",X"DD",X"74",X"0B",X"FD",X"5E",X"03",X"DD",X"73",
		X"06",X"DD",X"36",X"07",X"01",X"3E",X"F0",X"93",X"DD",X"77",X"0E",X"DD",X"36",X"0F",X"00",X"11",
		X"04",X"00",X"FD",X"19",X"11",X"10",X"00",X"DD",X"19",X"18",X"A9",X"3A",X"6A",X"E5",X"FE",X"01",
		X"20",X"05",X"CD",X"5B",X"2A",X"18",X"03",X"CD",X"D4",X"2A",X"C9",X"3A",X"53",X"E4",X"FE",X"0C",
		X"20",X"2E",X"11",X"15",X"00",X"2A",X"42",X"E4",X"19",X"22",X"42",X"E4",X"7C",X"2A",X"57",X"E4",
		X"26",X"00",X"01",X"9B",X"2B",X"09",X"BE",X"20",X"15",X"23",X"7E",X"32",X"4B",X"E4",X"3E",X"00",
		X"32",X"53",X"E4",X"32",X"4A",X"E4",X"3A",X"57",X"E4",X"C6",X"02",X"32",X"57",X"E4",X"18",X"43",
		X"3A",X"4B",X"E4",X"FE",X"01",X"20",X"05",X"11",X"F2",X"FF",X"18",X"03",X"11",X"0E",X"00",X"2A",
		X"40",X"E4",X"19",X"22",X"40",X"E4",X"7C",X"2A",X"57",X"E4",X"26",X"00",X"01",X"9B",X"2B",X"09",
		X"BE",X"20",X"15",X"23",X"7E",X"32",X"4B",X"E4",X"3E",X"0C",X"32",X"53",X"E4",X"32",X"4A",X"E4",
		X"3A",X"57",X"E4",X"C6",X"02",X"32",X"57",X"E4",X"3A",X"53",X"E4",X"FE",X"0C",X"28",X"04",X"47",
		X"CD",X"F1",X"10",X"C9",X"3A",X"6A",X"E5",X"FE",X"02",X"20",X"65",X"DD",X"21",X"40",X"E4",X"0E",
		X"05",X"DD",X"7E",X"0B",X"FE",X"01",X"20",X"1C",X"11",X"F4",X"FF",X"DD",X"6E",X"00",X"DD",X"66",
		X"01",X"19",X"DD",X"75",X"00",X"DD",X"74",X"01",X"7C",X"DD",X"BE",X"04",X"20",X"04",X"DD",X"36",
		X"0B",X"00",X"18",X"10",X"11",X"0C",X"00",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"19",X"DD",X"75",
		X"00",X"DD",X"74",X"01",X"11",X"F9",X"FF",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"19",X"DD",X"75",
		X"02",X"DD",X"74",X"03",X"C5",X"DD",X"46",X"06",X"79",X"FE",X"05",X"20",X"05",X"CD",X"F1",X"10",
		X"18",X"03",X"CD",X"2E",X"1A",X"C1",X"11",X"18",X"00",X"DD",X"19",X"0D",X"20",X"A3",X"18",X"5A",
		X"3A",X"6A",X"E5",X"FE",X"03",X"20",X"53",X"DD",X"21",X"40",X"E4",X"0E",X"06",X"11",X"EC",X"FF",
		X"DD",X"6E",X"00",X"DD",X"66",X"01",X"19",X"DD",X"75",X"00",X"DD",X"74",X"01",X"7C",X"FE",X"FE",
		X"20",X"04",X"DD",X"36",X"0A",X"FF",X"C5",X"DD",X"46",X"06",X"79",X"FE",X"06",X"20",X"05",X"CD",
		X"F1",X"10",X"18",X"03",X"CD",X"2E",X"1A",X"C1",X"11",X"18",X"00",X"DD",X"19",X"0D",X"20",X"CD",
		X"3A",X"53",X"E4",X"3C",X"32",X"53",X"E4",X"FE",X"24",X"20",X"0F",X"3E",X"00",X"32",X"53",X"E4",
		X"3A",X"57",X"E4",X"3C",X"32",X"57",X"E4",X"CD",X"9D",X"65",X"C9",X"03",X"01",X"06",X"00",X"07",
		X"00",X"08",X"00",X"0A",X"00",X"09",X"00",X"0D",X"00",X"0D",X"00",X"10",X"00",X"0F",X"00",X"13",
		X"00",X"11",X"00",X"19",X"00",X"32",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"65",X"07",X"07",X"07",X"CB",X"3C",X"1F",X"6F",X"11",X"10",X"D0",X"19",X"E5",X"11",X"80",X"01",
		X"19",X"D1",X"EB",X"7E",X"C9",X"67",X"FD",X"21",X"58",X"E4",X"11",X"18",X"00",X"3A",X"E9",X"E4",
		X"47",X"FD",X"7E",X"06",X"94",X"FE",X"12",X"30",X"6D",X"FE",X"08",X"38",X"69",X"FD",X"7E",X"07",
		X"95",X"30",X"02",X"ED",X"44",X"FE",X"06",X"30",X"5D",X"FD",X"7E",X"0C",X"B7",X"20",X"28",X"FD",
		X"7E",X"16",X"B7",X"20",X"22",X"3A",X"4F",X"E4",X"B7",X"28",X"15",X"FD",X"7E",X"0F",X"FE",X"FF",
		X"28",X"0E",X"21",X"52",X"E4",X"7E",X"B7",X"20",X"07",X"36",X"01",X"3E",X"0B",X"CD",X"73",X"30",
		X"3E",X"06",X"32",X"09",X"E5",X"18",X"2D",X"21",X"0B",X"E5",X"3A",X"44",X"E4",X"BE",X"28",X"24",
		X"7F",X"77",X"21",X"0A",X"E5",X"3A",X"4B",X"E4",X"BE",X"20",X"10",X"21",X"0C",X"E5",X"34",X"7E",
		X"FE",X"03",X"38",X"05",X"3E",X"13",X"32",X"06",X"E5",X"18",X"09",X"3A",X"4B",X"E4",X"77",X"3E",
		X"01",X"32",X"0C",X"E5",X"37",X"C9",X"11",X"18",X"00",X"FD",X"19",X"10",X"84",X"C9",X"C6",X"13",
		X"18",X"00",X"67",X"DD",X"E5",X"C1",X"FD",X"21",X"58",X"E4",X"3A",X"E9",X"E4",X"47",X"FD",X"E5",
		X"D1",X"7B",X"B9",X"28",X"32",X"FD",X"7E",X"0E",X"B7",X"20",X"2C",X"FD",X"7E",X"06",X"BC",X"30",
		X"26",X"C6",X"12",X"BC",X"38",X"21",X"FD",X"7E",X"07",X"95",X"30",X"02",X"ED",X"44",X"FE",X"06",
		X"30",X"15",X"DD",X"7E",X"0F",X"FD",X"BE",X"0F",X"20",X"04",X"37",X"C9",X"18",X"09",X"AF",X"FD",
		X"96",X"0C",X"D8",X"DD",X"96",X"0C",X"D8",X"11",X"18",X"00",X"FD",X"19",X"10",X"C0",X"C9",X"67",
		X"DD",X"E5",X"C1",X"FD",X"21",X"58",X"E4",X"3A",X"E9",X"E4",X"47",X"FD",X"E5",X"D1",X"7B",X"91",
		X"5F",X"28",X"26",X"FD",X"7E",X"0E",X"B7",X"20",X"20",X"FD",X"7E",X"07",X"C6",X"07",X"BC",X"38",
		X"18",X"D6",X"08",X"BC",X"30",X"13",X"3C",X"BC",X"20",X"04",X"CB",X"7B",X"20",X"0B",X"FD",X"7E",
		X"06",X"95",X"30",X"02",X"ED",X"44",X"FE",X"0F",X"D8",X"11",X"18",X"00",X"FD",X"19",X"10",X"CB",
		X"C9",X"C6",X"08",X"67",X"DD",X"E5",X"C1",X"FD",X"21",X"58",X"E4",X"3A",X"E9",X"E4",X"47",X"FD",
		X"E5",X"D1",X"7B",X"91",X"5F",X"28",X"22",X"FD",X"7E",X"0E",X"B7",X"20",X"1C",X"FD",X"7E",X"07",
		X"BC",X"30",X"16",X"C6",X"08",X"BC",X"38",X"11",X"20",X"04",X"CB",X"7B",X"20",X"0B",X"FD",X"7E",
		X"06",X"95",X"30",X"02",X"ED",X"44",X"FE",X"0F",X"D8",X"11",X"18",X"00",X"FD",X"19",X"10",X"CF",
		X"C9",X"1A",X"A0",X"B9",X"C8",X"E5",X"21",X"80",X"00",X"19",X"7E",X"E1",X"A0",X"B9",X"C9",X"1A",
		X"A0",X"B9",X"C0",X"E5",X"21",X"80",X"00",X"19",X"7E",X"E1",X"A0",X"B9",X"C9",X"7E",X"A0",X"B9",
		X"C8",X"24",X"7E",X"25",X"A0",X"B9",X"C9",X"7E",X"A0",X"B9",X"C0",X"24",X"7E",X"25",X"A0",X"B9",
		X"C9",X"7E",X"B9",X"C8",X"24",X"7E",X"25",X"B9",X"C9",X"1A",X"B9",X"C0",X"E5",X"21",X"80",X"00",
		X"19",X"7E",X"E1",X"B9",X"C9",X"C6",X"05",X"18",X"00",X"4F",X"3A",X"47",X"E4",X"B9",X"D0",X"C6",
		X"04",X"B9",X"D8",X"3A",X"46",X"E4",X"95",X"30",X"02",X"ED",X"44",X"FE",X"0A",X"D0",X"AF",X"32",
		X"50",X"E4",X"C9",X"4F",X"3A",X"46",X"E4",X"C6",X"0E",X"B9",X"D8",X"D6",X"1D",X"30",X"01",X"AF",
		X"B9",X"D0",X"3A",X"47",X"E4",X"95",X"30",X"02",X"ED",X"44",X"FE",X"03",X"D0",X"AF",X"32",X"50",
		X"E4",X"C9",X"4F",X"3A",X"46",X"E4",X"91",X"30",X"02",X"ED",X"44",X"FE",X"0E",X"D0",X"3A",X"47",
		X"E4",X"95",X"30",X"02",X"ED",X"44",X"FE",X"03",X"D0",X"AF",X"32",X"50",X"E4",X"C9",X"EB",X"7E",
		X"C6",X"70",X"77",X"2C",X"36",X"0A",X"2C",X"7E",X"C6",X"74",X"77",X"2C",X"36",X"0A",X"01",X"80",
		X"00",X"09",X"36",X"0A",X"2D",X"7E",X"C6",X"7C",X"77",X"2D",X"36",X"0A",X"2D",X"7E",X"C6",X"78",
		X"77",X"ED",X"42",X"EB",X"C9",X"EB",X"7E",X"C6",X"60",X"77",X"2C",X"36",X"0A",X"2C",X"7E",X"C6",
		X"64",X"77",X"2C",X"36",X"0A",X"01",X"80",X"00",X"09",X"36",X"0A",X"2D",X"7E",X"C6",X"6C",X"77",
		X"2D",X"36",X"0A",X"2D",X"7E",X"C6",X"68",X"77",X"ED",X"42",X"EB",X"C9",X"EB",X"7E",X"D6",X"70",
		X"77",X"2C",X"36",X"05",X"2C",X"7E",X"D6",X"74",X"77",X"2C",X"36",X"05",X"01",X"80",X"00",X"09",
		X"36",X"05",X"2D",X"7E",X"D6",X"7C",X"77",X"2D",X"36",X"05",X"2D",X"7E",X"D6",X"78",X"77",X"ED",
		X"42",X"EB",X"C9",X"EB",X"7E",X"D6",X"60",X"77",X"2C",X"36",X"05",X"2C",X"7E",X"D6",X"64",X"77",
		X"2C",X"36",X"05",X"01",X"80",X"00",X"09",X"36",X"05",X"2D",X"7E",X"D6",X"6C",X"77",X"2D",X"36",
		X"05",X"2D",X"7E",X"D6",X"68",X"77",X"ED",X"42",X"EB",X"C9",X"D5",X"07",X"07",X"07",X"CB",X"3C",
		X"1F",X"6F",X"11",X"10",X"D0",X"19",X"EB",X"C5",X"CD",X"0E",X"2F",X"C1",X"D1",X"C9",X"EB",X"77",
		X"23",X"23",X"77",X"01",X"80",X"00",X"09",X"77",X"2B",X"2B",X"77",X"ED",X"42",X"EB",X"C9",X"21",
		X"91",X"E5",X"7E",X"47",X"81",X"27",X"77",X"38",X"36",X"18",X"17",X"21",X"93",X"E5",X"7E",X"81",
		X"27",X"77",X"2B",X"7E",X"88",X"27",X"77",X"2B",X"7E",X"47",X"CE",X"00",X"27",X"77",X"38",X"1F",
		X"B8",X"C8",X"4F",X"78",X"C6",X"01",X"27",X"47",X"C5",X"FE",X"05",X"20",X"0C",X"21",X"8F",X"E5",
		X"34",X"3E",X"12",X"CD",X"42",X"31",X"CD",X"F7",X"31",X"C1",X"78",X"B9",X"38",X"E5",X"C9",X"21",
		X"99",X"99",X"22",X"91",X"E5",X"22",X"92",X"E5",X"C9",X"D5",X"EB",X"3A",X"D8",X"E5",X"77",X"2C",
		X"2C",X"77",X"01",X"80",X"00",X"09",X"77",X"2D",X"2D",X"77",X"EB",X"D1",X"C9",X"1A",X"B7",X"C8",
		X"FE",X"20",X"30",X"03",X"4F",X"18",X"04",X"77",X"2C",X"71",X"2C",X"13",X"18",X"EF",X"32",X"B5",
		X"E5",X"3A",X"B5",X"E5",X"A7",X"20",X"FA",X"C9",X"06",X"00",X"D6",X"0A",X"04",X"30",X"FB",X"C6",
		X"0A",X"05",X"F5",X"78",X"CD",X"58",X"30",X"F1",X"C6",X"30",X"77",X"23",X"71",X"23",X"C9",X"1A",
		X"F5",X"0F",X"0F",X"0F",X"0F",X"CD",X"6A",X"30",X"F1",X"13",X"E6",X"0F",X"C6",X"30",X"77",X"23",
		X"71",X"23",X"C9",X"4F",X"06",X"00",X"21",X"28",X"31",X"09",X"56",X"21",X"FE",X"E4",X"5E",X"34",
		X"7A",X"32",X"88",X"E5",X"B7",X"28",X"09",X"34",X"7B",X"FE",X"07",X"20",X"03",X"1E",X"00",X"34",
		X"CB",X"9E",X"7B",X"32",X"89",X"E5",X"87",X"87",X"87",X"FD",X"21",X"C0",X"E3",X"5F",X"16",X"00",
		X"FD",X"19",X"FD",X"36",X"00",X"11",X"FD",X"36",X"08",X"11",X"16",X"15",X"79",X"FE",X"0B",X"38",
		X"02",X"16",X"03",X"3A",X"46",X"E4",X"82",X"ED",X"44",X"5F",X"16",X"00",X"2A",X"E3",X"E5",X"19",
		X"FD",X"75",X"02",X"FD",X"74",X"03",X"1E",X"00",X"3A",X"88",X"E5",X"B7",X"28",X"0A",X"1C",X"FD",
		X"77",X"0C",X"FD",X"75",X"0A",X"FD",X"74",X"0B",X"21",X"1B",X"31",X"09",X"7E",X"FD",X"77",X"04",
		X"21",X"35",X"31",X"09",X"46",X"0E",X"00",X"CD",X"DB",X"2F",X"3A",X"47",X"E4",X"C6",X"20",X"6F",
		X"26",X"00",X"29",X"FD",X"75",X"06",X"FD",X"74",X"07",X"CB",X"43",X"28",X"0A",X"01",X"F0",X"FF",
		X"09",X"FD",X"75",X"0E",X"FD",X"74",X"0F",X"3A",X"89",X"E5",X"4F",X"06",X"00",X"21",X"9E",X"E5",
		X"09",X"36",X"70",X"CB",X"43",X"28",X"03",X"23",X"36",X"70",X"C9",X"F8",X"F9",X"FB",X"FC",X"FA",
		X"FD",X"FA",X"FD",X"E1",X"E1",X"E1",X"E1",X"E1",X"00",X"00",X"00",X"00",X"00",X"FE",X"FE",X"FF",
		X"F0",X"AA",X"AB",X"F1",X"F0",X"02",X"04",X"06",X"08",X"05",X"10",X"15",X"20",X"30",X"50",X"80",
		X"10",X"30",X"D5",X"57",X"FE",X"12",X"28",X"08",X"3A",X"A7",X"E5",X"B7",X"28",X"02",X"D1",X"C9",
		X"7A",X"E5",X"21",X"BB",X"E5",X"5E",X"16",X"00",X"21",X"BC",X"E5",X"19",X"57",X"1C",X"7B",X"E6",
		X"0F",X"32",X"BB",X"E5",X"72",X"E1",X"D1",X"C9",X"3A",X"BA",X"E5",X"21",X"BB",X"E5",X"BE",X"C8",
		X"5F",X"16",X"00",X"21",X"BC",X"E5",X"19",X"3C",X"E6",X"0F",X"32",X"BA",X"E5",X"7E",X"D3",X"00",
		X"F6",X"80",X"D3",X"00",X"C9",X"11",X"92",X"31",X"CD",X"2D",X"30",X"3A",X"8E",X"E5",X"CD",X"48",
		X"30",X"C9",X"06",X"52",X"4F",X"55",X"4E",X"44",X"2D",X"00",X"3A",X"8E",X"E5",X"3D",X"CD",X"EC",
		X"31",X"79",X"3C",X"32",X"CC",X"E5",X"0E",X"06",X"FE",X"0A",X"38",X"05",X"CD",X"48",X"30",X"18",
		X"05",X"2C",X"2C",X"CD",X"6A",X"30",X"3A",X"CC",X"E5",X"FE",X"04",X"38",X"01",X"AF",X"87",X"87",
		X"5F",X"16",X"00",X"E5",X"21",X"D4",X"31",X"19",X"EB",X"E1",X"CD",X"2D",X"30",X"11",X"E4",X"31",
		X"CD",X"2D",X"30",X"C9",X"06",X"54",X"48",X"00",X"06",X"53",X"54",X"00",X"06",X"4E",X"44",X"00",
		X"06",X"52",X"44",X"00",X"06",X"20",X"42",X"4C",X"4F",X"43",X"4B",X"00",X"0E",X"00",X"0C",X"D6",
		X"03",X"30",X"FB",X"0D",X"C6",X"03",X"C9",X"0E",X"1E",X"21",X"56",X"D0",X"3A",X"8F",X"E5",X"CD",
		X"6A",X"30",X"C9",X"21",X"26",X"D0",X"11",X"8A",X"E5",X"0E",X"1E",X"1A",X"E6",X"0F",X"CD",X"6A",
		X"30",X"13",X"CD",X"5F",X"30",X"1A",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"CD",X"6A",X"30",X"0E",
		X"04",X"21",X"18",X"D0",X"3A",X"B8",X"E5",X"B7",X"28",X"03",X"21",X"60",X"D0",X"3A",X"AD",X"E6",
		X"B7",X"28",X"26",X"E5",X"21",X"B6",X"E5",X"7E",X"B7",X"20",X"06",X"36",X"16",X"21",X"AD",X"E6",
		X"35",X"3A",X"AD",X"E6",X"E1",X"1F",X"30",X"0C",X"36",X"00",X"54",X"5D",X"13",X"01",X"0B",X"00",
		X"ED",X"B0",X"18",X"03",X"CD",X"82",X"32",X"18",X"03",X"CD",X"82",X"32",X"11",X"9A",X"E5",X"21",
		X"91",X"E5",X"06",X"03",X"1A",X"BE",X"13",X"23",X"20",X"02",X"10",X"F8",X"D0",X"3A",X"A7",X"E5",
		X"B7",X"C0",X"01",X"03",X"00",X"11",X"9A",X"E5",X"21",X"91",X"E5",X"ED",X"B0",X"0E",X"06",X"21",
		X"38",X"D0",X"11",X"91",X"E5",X"06",X"03",X"CD",X"5F",X"30",X"10",X"FB",X"C9",X"11",X"B8",X"E6",
		X"21",X"20",X"D7",X"01",X"40",X"00",X"ED",X"B0",X"21",X"A0",X"D7",X"01",X"40",X"00",X"ED",X"B0",
		X"21",X"20",X"D8",X"01",X"40",X"00",X"ED",X"B0",X"21",X"B8",X"D8",X"01",X"0E",X"00",X"ED",X"B0",
		X"21",X"38",X"D9",X"01",X"0E",X"00",X"ED",X"B0",X"C9",X"21",X"B8",X"E6",X"11",X"20",X"D7",X"01",
		X"40",X"00",X"ED",X"B0",X"11",X"A0",X"D7",X"01",X"40",X"00",X"ED",X"B0",X"11",X"20",X"D8",X"01",
		X"40",X"00",X"ED",X"B0",X"11",X"B8",X"D8",X"01",X"0E",X"00",X"ED",X"B0",X"11",X"38",X"D9",X"01",
		X"0E",X"00",X"ED",X"B0",X"C9",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"00",X"00",X"32",X"34",X"01",X"35",X"72",X"35",X"4B",X"3C",X"62",X"36",X"CE",X"36",X"45",X"37",
		X"89",X"34",X"CA",X"3C",X"A8",X"3B",X"04",X"3E",X"E2",X"35",X"59",X"3D",X"8C",X"3F",X"9B",X"39",
		X"A9",X"3E",X"F9",X"38",X"CC",X"3A",X"1E",X"3F",X"2F",X"3A",X"C5",X"37",X"71",X"38",X"7D",X"40",
		X"F7",X"3F",X"00",X"01",X"AE",X"E5",X"A4",X"EB",X"A9",X"CF",X"F7",X"A9",X"8D",X"CA",X"AE",X"CA",
		X"F7",X"B3",X"F1",X"B9",X"C5",X"E8",X"D2",X"F7",X"BE",X"F7",X"03",X"84",X"8D",X"C5",X"8E",X"92",
		X"C2",X"89",X"8D",X"D5",X"CB",X"8E",X"98",X"D2",X"99",X"9D",X"C4",X"D7",X"93",X"98",X"C7",X"04",
		X"A6",X"C6",X"EE",X"04",X"B6",X"C8",X"F1",X"04",X"06",X"81",X"88",X"CF",X"07",X"A2",X"C3",X"A7",
		X"D3",X"AC",X"D1",X"B7",X"C6",X"D5",X"BC",X"CF",X"0A",X"A4",X"CB",X"A9",X"CA",X"BE",X"C0",X"09",
		X"BB",X"CC",X"08",X"AB",X"C3",X"D3",X"B0",X"CC",X"1F",X"00",X"01",X"A4",X"C2",X"A9",X"C1",X"E3",
		X"A5",X"CA",X"F1",X"A7",X"D3",X"F6",X"AC",X"CF",X"F6",X"B0",X"95",X"C1",X"E3",X"B4",X"D3",X"F7",
		X"B0",X"C6",X"E7",X"CA",X"ED",X"B9",X"EC",X"D4",X"F7",X"BE",X"F7",X"02",X"A4",X"C1",X"C3",X"90",
		X"98",X"C0",X"C4",X"B0",X"C5",X"C8",X"04",X"A9",X"C5",X"ED",X"B6",X"CD",X"F1",X"03",X"84",X"8F",
		X"C0",X"C4",X"85",X"8B",X"D2",X"8C",X"91",X"CE",X"87",X"93",X"D7",X"85",X"98",X"C9",X"94",X"98",
		X"D5",X"94",X"9D",X"D2",X"99",X"9D",X"C7",X"06",X"A1",X"86",X"D7",X"07",X"A2",X"C2",X"A3",X"CF",
		X"A5",X"D4",X"A7",X"C1",X"AB",X"C2",X"AE",X"C6",X"CB",X"B7",X"C1",X"C5",X"D7",X"BC",X"C0",X"D7",
		X"09",X"BB",X"CA",X"08",X"A6",X"C3",X"A9",X"D1",X"AD",X"C3",X"0A",X"B9",X"D4",X"BE",X"C0",X"D7",
		X"1F",X"00",X"01",X"A5",X"CA",X"F2",X"A6",X"E3",X"A8",X"D4",X"F7",X"AB",X"C5",X"F3",X"AF",X"E4",
		X"B0",X"CA",X"F1",X"B3",X"D7",X"B5",X"CC",X"F3",X"B7",X"CC",X"D3",X"B9",X"EC",X"D3",X"F7",X"BA",
		X"9D",X"CF",X"F0",X"BE",X"F7",X"04",X"AE",X"D4",X"AF",X"D5",X"B0",X"D6",X"B2",X"C4",X"E8",X"03",
		X"99",X"9D",X"C2",X"D6",X"9A",X"9D",X"CE",X"D1",X"95",X"98",X"CB",X"D4",X"90",X"94",X"C9",X"CF",
		X"8F",X"98",X"C3",X"8B",X"8F",X"CC",X"D1",X"86",X"8E",X"C4",X"85",X"8A",X"C9",X"D3",X"06",X"A1",
		X"87",X"D7",X"07",X"A3",X"CE",X"A4",X"C2",X"A9",X"CF",X"AD",X"C1",X"B1",X"D7",X"B8",X"D0",X"BC",
		X"D4",X"08",X"A8",X"C6",X"AD",X"CE",X"B2",X"D2",X"09",X"B6",X"C9",X"0A",X"B3",X"D7",X"BE",X"C0",
		X"D7",X"1F",X"00",X"01",X"A4",X"C0",X"D0",X"F7",X"A6",X"E1",X"CF",X"F0",X"A8",X"C1",X"C2",X"CE",
		X"CF",X"A9",X"D2",X"F6",X"AA",X"C2",X"C3",X"CD",X"CE",X"AC",X"C3",X"C4",X"CC",X"CD",X"AE",X"C3",
		X"E5",X"CB",X"ED",X"AF",X"E5",X"CB",X"F7",X"B0",X"C6",X"CA",X"B2",X"C6",X"EA",X"B4",X"C1",X"E3",
		X"CD",X"F3",X"B9",X"C5",X"F7",X"BE",X"F7",X"03",X"A4",X"8E",X"D3",X"AF",X"93",X"C2",X"AF",X"95",
		X"CE",X"B2",X"95",X"C8",X"B4",X"9A",X"C4",X"D1",X"B4",X"9D",X"C0",X"B9",X"9D",X"CB",X"D5",X"06",
		X"A1",X"91",X"C8",X"07",X"A2",X"D1",X"A7",X"D6",X"AC",X"CB",X"AD",X"C0",X"B2",X"C3",X"D3",X"B7",
		X"C8",X"08",X"AC",X"C1",X"B1",X"C4",X"B6",X"CE",X"09",X"BB",X"CE",X"0A",X"A9",X"D2",X"D6",X"BE",
		X"D7",X"1F",X"01",X"01",X"A6",X"98",X"C9",X"CE",X"A8",X"9A",X"C1",X"C4",X"D3",X"D6",X"A8",X"C2",
		X"C3",X"D4",X"D5",X"AF",X"C2",X"C3",X"D4",X"D5",X"B2",X"CB",X"CC",X"B9",X"C1",X"E5",X"C9",X"CA",
		X"CD",X"CE",X"D2",X"F6",X"BB",X"9D",X"C6",X"D1",X"BE",X"F7",X"02",X"B9",X"CB",X"CC",X"04",X"A8",
		X"C6",X"C7",X"D0",X"D1",X"B3",X"C6",X"E8",X"CF",X"F1",X"03",X"A6",X"8A",X"C8",X"CF",X"A8",X"94",
		X"C5",X"D2",X"B2",X"98",X"CA",X"CD",X"B6",X"9D",X"C8",X"CF",X"A8",X"9D",X"C0",X"D7",X"06",X"A1",
		X"91",X"CA",X"CD",X"07",X"A6",X"C2",X"D5",X"AD",X"C3",X"D4",X"B7",X"C2",X"CB",X"D5",X"08",X"A5",
		X"C4",X"D3",X"B6",X"CC",X"BB",X"C7",X"09",X"BB",X"CC",X"0A",X"A6",X"CE",X"BE",X"C5",X"BE",X"D2",
		X"0D",X"8E",X"C2",X"C3",X"D4",X"D5",X"98",X"C2",X"C3",X"D4",X"D5",X"98",X"CB",X"CC",X"91",X"CA",
		X"ED",X"1F",X"00",X"01",X"A4",X"C0",X"C2",X"C4",X"C6",X"C8",X"CA",X"CC",X"CE",X"D0",X"D2",X"D4",
		X"A9",X"8B",X"C0",X"C2",X"C4",X"C6",X"C8",X"CA",X"CC",X"CE",X"D0",X"D2",X"D4",X"AF",X"C0",X"C2",
		X"C4",X"C6",X"C8",X"CA",X"CC",X"CE",X"D0",X"D2",X"D4",X"A4",X"93",X"D6",X"B4",X"C1",X"F6",X"BE",
		X"F7",X"02",X"B9",X"C1",X"F6",X"03",X"A4",X"93",X"C1",X"C3",X"C5",X"C7",X"C9",X"CB",X"CD",X"CF",
		X"D1",X"D3",X"D5",X"B4",X"9D",X"C0",X"06",X"A1",X"9D",X"D7",X"07",X"A7",X"C0",X"C8",X"D0",X"AD",
		X"C4",X"CC",X"D4",X"B2",X"C0",X"B7",X"C6",X"CA",X"CE",X"BC",X"C1",X"D6",X"08",X"A1",X"CA",X"D3",
		X"B6",X"C8",X"D0",X"09",X"BB",X"C8",X"0A",X"A4",X"C0",X"A9",X"C0",X"AF",X"C0",X"1F",X"00",X"01",
		X"A5",X"C0",X"E2",X"C6",X"EB",X"CE",X"F0",X"AD",X"91",X"D3",X"D6",X"AD",X"D7",X"AF",X"C1",X"EA",
		X"B0",X"D4",X"B0",X"94",X"D5",X"B4",X"C0",X"E3",X"CA",X"EC",X"B5",X"D3",X"F6",X"B9",X"C0",X"E6",
		X"BE",X"F7",X"04",X"A2",X"C4",X"C5",X"A5",X"D2",X"F7",X"A9",X"C4",X"E8",X"B6",X"CE",X"F0",X"03",
		X"A5",X"8A",X"C3",X"A5",X"9D",X"D1",X"A7",X"95",X"C9",X"AF",X"93",X"C0",X"B2",X"9D",X"D7",X"B4",
		X"98",X"C4",X"CD",X"B9",X"9D",X"C7",X"06",X"A1",X"86",X"CC",X"07",X"A3",X"C0",X"C6",X"D0",X"AD",
		X"C6",X"CA",X"AE",X"D4",X"B1",X"CF",X"B3",X"D3",X"D6",X"B7",X"C1",X"BC",X"C1",X"CD",X"D6",X"08",
		X"A2",X"C1",X"C9",X"CF",X"AC",X"C3",X"09",X"BB",X"CB",X"0A",X"A5",X"CA",X"B5",X"D4",X"BE",X"C0",
		X"0D",X"8F",X"D4",X"D5",X"1F",X"00",X"01",X"A4",X"C1",X"E8",X"A6",X"CA",X"EE",X"D2",X"F7",X"A8",
		X"8A",X"CE",X"A9",X"C2",X"E7",X"AB",X"CE",X"F7",X"AD",X"92",X"D6",X"B1",X"D2",X"F4",X"B0",X"95",
		X"C2",X"E4",X"C7",X"B2",X"C6",X"B4",X"C5",X"C6",X"B7",X"CE",X"F2",X"B6",X"D6",X"D7",X"B9",X"C5",
		X"BE",X"F7",X"02",X"AB",X"9A",X"CB",X"AB",X"CC",X"B1",X"9A",X"CC",X"B9",X"C1",X"E4",X"C6",X"EA",
		X"04",X"AE",X"CC",X"F1",X"03",X"A4",X"9D",X"C0",X"A4",X"98",X"C9",X"A6",X"8A",X"CF",X"D4",X"B0",
		X"95",X"D7",X"B1",X"9D",X"D5",X"06",X"A1",X"85",X"D2",X"07",X"A4",X"CF",X"D3",X"D7",X"A6",X"D1",
		X"A7",X"C2",X"C7",X"A9",X"CB",X"CC",X"D7",X"AE",X"D7",X"AF",X"CC",X"D3",X"B2",X"C5",X"B5",X"D0",
		X"08",X"A1",X"C4",X"A3",X"CC",X"A8",X"D2",X"09",X"BB",X"CC",X"0A",X"A9",X"C6",X"B1",X"D3",X"BE",
		X"D7",X"0E",X"93",X"C5",X"1F",X"01",X"01",X"A5",X"C0",X"E2",X"C4",X"A8",X"D3",X"F6",X"AA",X"C6",
		X"F1",X"AA",X"8C",X"D5",X"AB",X"C1",X"E3",X"AA",X"9D",X"C6",X"AA",X"9A",X"D1",X"AD",X"D3",X"F7",
		X"AF",X"C7",X"E9",X"CD",X"EF",X"AF",X"94",X"D3",X"B0",X"92",X"C3",X"B2",X"C0",X"E2",X"B3",X"D3",
		X"F7",X"B4",X"96",X"C5",X"C9",X"CD",X"B6",X"98",X"C4",X"B7",X"C7",X"F0",X"B8",X"9A",X"C3",X"B9",
		X"D2",X"B8",X"D5",X"F7",X"BC",X"C2",X"D3",X"BE",X"C0",X"F7",X"04",X"A7",X"C4",X"C5",X"A5",X"D1",
		X"F3",X"AC",X"C8",X"EF",X"B1",X"C7",X"EF",X"AA",X"D2",X"03",X"A1",X"84",X"C0",X"A8",X"8C",X"D7",
		X"A9",X"C3",X"AA",X"8D",X"CB",X"AB",X"91",X"C0",X"AC",X"96",X"D0",X"AD",X"92",X"D6",X"B1",X"96",
		X"CB",X"B2",X"9D",X"C1",X"B3",X"97",X"D5",X"B4",X"96",X"C7",X"CE",X"B8",X"9D",X"D4",X"06",X"A5",
		X"89",X"C3",X"07",X"AB",X"D4",X"AD",X"C7",X"CF",X"B1",X"D4",X"B5",X"C8",X"CA",X"CC",X"CF",X"B6",
		X"C3",X"D7",X"B7",X"D2",X"BC",X"C0",X"C4",X"CA",X"CC",X"D7",X"08",X"A5",X"D4",X"A7",X"C8",X"BB",
		X"C5",X"09",X"A8",X"C2",X"0A",X"A5",X"C2",X"BE",X"C0",X"D7",X"0F",X"9D",X"C3",X"E5",X"C7",X"F2",
		X"1F",X"00",X"01",X"A4",X"C1",X"C2",X"A9",X"C1",X"E6",X"CA",X"F6",X"A9",X"9B",X"CA",X"AE",X"C0",
		X"E7",X"CD",X"F5",X"B0",X"92",X"CD",X"D5",X"B3",X"C4",X"E6",X"CB",X"ED",X"D0",X"F5",X"B5",X"97",
		X"C6",X"D5",X"B8",X"C2",X"E6",X"CB",X"F5",X"BA",X"C0",X"E2",X"BD",X"C4",X"C8",X"C9",X"CF",X"F7",
		X"02",X"9F",X"C0",X"F7",X"04",X"A3",X"C7",X"F6",X"BA",X"C4",X"E7",X"03",X"A4",X"8D",X"C0",X"A6",
		X"88",X"C6",X"A9",X"97",X"C3",X"A9",X"9C",X"D7",X"AE",X"9C",X"C8",X"B3",X"97",X"CF",X"D4",X"BA",
		X"9E",X"C3",X"BD",X"CE",X"06",X"A1",X"85",X"C3",X"07",X"A2",X"C1",X"A7",X"D3",X"AC",X"C1",X"C4",
		X"CE",X"B1",X"C6",X"CB",X"D1",X"B6",X"C5",X"D0",X"D3",X"B8",X"C0",X"C1",X"BD",X"C0",X"C5",X"CA",
		X"08",X"A6",X"CD",X"B0",X"C4",X"BC",X"C6",X"09",X"A1",X"C2",X"0A",X"B3",X"D1",X"AE",X"CD",X"D5",
		X"0D",X"99",X"C0",X"C1",X"0F",X"9E",X"C5",X"E7",X"1F",X"00",X"01",X"AA",X"C2",X"CE",X"AC",X"C0",
		X"E2",X"AE",X"90",X"C2",X"B1",X"C0",X"E3",X"D3",X"F6",X"B3",X"9D",X"C0",X"B6",X"C1",X"E4",X"CD",
		X"B7",X"D0",X"F6",X"B8",X"C7",X"ED",X"B9",X"CD",X"D0",X"D4",X"9B",X"C5",X"D4",X"BC",X"C4",X"C5",
		X"D1",X"F7",X"BE",X"C0",X"F7",X"02",X"A5",X"C0",X"E2",X"C4",X"ED",X"AA",X"95",X"CD",X"AC",X"90",
		X"CE",X"AF",X"CF",X"D0",X"04",X"A4",X"CE",X"F4",X"A7",X"CA",X"EC",X"AB",X"D0",X"F5",X"AE",X"C4",
		X"EC",X"B1",X"CE",X"F1",X"B8",X"C2",X"E4",X"03",X"A1",X"84",X"D5",X"A7",X"90",X"C3",X"A7",X"C9",
		X"AA",X"8E",X"CF",X"AB",X"90",X"D6",X"AC",X"97",X"C9",X"B1",X"97",X"CC",X"B4",X"9D",X"CE",X"AE",
		X"9B",X"D7",X"B8",X"9D",X"C1",X"C6",X"BA",X"9D",X"CC",X"06",X"A5",X"C3",X"07",X"AA",X"C1",X"CC",
		X"AD",X"D0",X"AF",X"C5",X"C8",X"CB",X"C0",X"B4",X"C1",X"B5",X"D2",X"BA",X"D1",X"D3",X"D6",X"BC",
		X"C3",X"C7",X"CB",X"08",X"A7",X"CE",X"B3",X"C3",X"B4",X"D1",X"BB",X"C9",X"09",X"B5",X"C7",X"0A",
		X"AA",X"CE",X"BC",X"D3",X"BC",X"D5",X"0D",X"8B",X"C0",X"C1",X"1F",X"00",X"01",X"A4",X"CC",X"F7",
		X"A5",X"C7",X"E9",X"A9",X"CD",X"F6",X"AA",X"C1",X"E4",X"AF",X"C5",X"C7",X"E9",X"B4",X"C4",X"B9",
		X"C2",X"C3",X"C7",X"E9",X"CD",X"F7",X"BE",X"C0",X"F7",X"02",X"AA",X"C8",X"EA",X"8B",X"CD",X"F6",
		X"AC",X"98",X"CD",X"AC",X"95",X"D6",X"AF",X"CF",X"F4",X"B1",X"93",X"CF",X"B4",X"C8",X"EA",X"CF",
		X"F6",X"04",X"A2",X"C1",X"E5",X"03",X"A4",X"88",X"D1",X"A5",X"89",X"CA",X"A5",X"9D",X"C0",X"A9",
		X"9D",X"CC",X"A9",X"98",X"D7",X"AA",X"8E",X"C5",X"C7",X"AF",X"93",X"C4",X"CA",X"D5",X"AF",X"98",
		X"CE",X"B4",X"98",X"C3",X"C7",X"B9",X"9D",X"C1",X"B9",X"CA",X"06",X"A1",X"86",X"C6",X"BB",X"9D",
		X"CA",X"07",X"A2",X"CC",X"D6",X"A3",X"C9",X"A8",X"C2",X"C4",X"C9",X"AD",X"C9",X"D0",X"D3",X"B2",
		X"C9",X"D1",X"D3",X"B7",X"C4",X"C9",X"D1",X"BC",X"C2",X"CE",X"D6",X"08",X"A1",X"D4",X"A7",X"C3",
		X"A6",X"D4",X"AC",X"CB",X"09",X"A6",X"CB",X"0A",X"A5",X"C9",X"AF",X"C9",X"BE",X"D7",X"1F",X"00",
		X"01",X"A7",X"C1",X"C5",X"EA",X"CD",X"F3",X"D5",X"F7",X"A9",X"D6",X"AF",X"C5",X"E8",X"D2",X"F7",
		X"B6",X"C0",X"E6",X"B8",X"C6",X"EA",X"CF",X"F1",X"D3",X"D5",X"F7",X"BA",X"D3",X"F7",X"BC",X"D4",
		X"F7",X"BD",X"C0",X"EA",X"CF",X"F7",X"02",X"A5",X"D5",X"AF",X"CA",X"F1",X"B8",X"CC",X"ED",X"9F",
		X"C0",X"F7",X"04",X"A2",X"C3",X"CB",X"CC",X"D4",X"F7",X"A9",X"C6",X"F3",X"AB",X"D6",X"B0",X"C1",
		X"C2",X"B1",X"D2",X"F4",X"B5",X"D2",X"03",X"A1",X"92",X"C0",X"A2",X"86",X"D3",X"A5",X"89",X"C4",
		X"A5",X"CA",X"A7",X"8A",X"D4",X"A9",X"8B",X"D5",X"A9",X"8E",X"C5",X"D7",X"AF",X"97",X"C9",X"B4",
		X"97",X"D1",X"B6",X"C7",X"B8",X"9E",X"CB",X"CE",X"06",X"A1",X"84",X"CA",X"07",X"A5",X"C1",X"C5",
		X"C9",X"CE",X"D1",X"D7",X"AA",X"C7",X"CB",X"D0",X"B4",X"C0",X"C3",X"B6",X"D7",X"B8",X"D4",X"BB",
		X"C0",X"C2",X"BD",X"CC",X"08",X"A4",X"C7",X"D0",X"AC",X"D4",X"09",X"B5",X"CC",X"0A",X"A7",X"C1",
		X"B8",X"D7",X"BD",X"C0",X"0D",X"86",X"D6",X"D7",X"0E",X"99",X"D4",X"1F",X"01",X"01",X"A2",X"C8",
		X"CF",X"D5",X"A3",X"C8",X"D0",X"D4",X"A4",X"C7",X"D4",X"A5",X"C1",X"E6",X"CD",X"D1",X"F3",X"85",
		X"CD",X"F0",X"A7",X"C6",X"CD",X"D1",X"A9",X"C6",X"F6",X"AA",X"C0",X"E4",X"AE",X"C6",X"F7",X"AF",
		X"C1",X"E4",X"B0",X"93",X"C4",X"C6",X"D1",X"D3",X"B3",X"D4",X"B3",X"95",X"C7",X"D5",X"94",X"C4",
		X"B4",X"96",X"C3",X"D1",X"B5",X"97",X"C8",X"B6",X"98",X"C2",X"B6",X"D0",X"D1",X"D5",X"F7",X"B7",
		X"9A",X"C9",X"B8",X"9A",X"C1",X"B8",X"CE",X"F1",X"B9",X"C6",X"BA",X"C4",X"CA",X"EE",X"BC",X"C3",
		X"C4",X"C7",X"BB",X"9D",X"D5",X"D7",X"BD",X"CF",X"F1",X"BE",X"C0",X"E8",X"CF",X"F7",X"02",X"A5",
		X"C0",X"C2",X"C3",X"9F",X"C9",X"EE",X"04",X"A6",X"C7",X"F0",X"B0",X"C7",X"F0",X"B1",X"C1",X"E3",
		X"03",X"A5",X"9D",X"C5",X"D2",X"A9",X"8D",X"D7",X"AA",X"8E",X"C3",X"AF",X"9D",X"C0",X"B8",X"CD",
		X"BA",X"9E",X"CC",X"BB",X"9D",X"C8",X"BB",X"9E",X"C9",X"06",X"A1",X"88",X"CB",X"BB",X"9D",X"D6",
		X"07",X"A3",X"C0",X"C6",X"D3",X"A7",X"C8",X"CE",X"D0",X"D4",X"A8",X"C0",X"B1",X"C8",X"B3",X"CA",
		X"CE",X"B2",X"C3",X"B4",X"D6",X"B9",X"D7",X"BA",X"C3",X"BB",X"D1",X"BC",X"C1",X"C6",X"D3",X"BD",
		X"CA",X"CE",X"08",X"A2",X"C3",X"BB",X"C2",X"D4",X"09",X"AB",X"CA",X"0A",X"B3",X"D4",X"B8",X"CE",
		X"BC",X"C3",X"0D",X"88",X"C7",X"EC",X"CE",X"F0",X"92",X"D4",X"D5",X"95",X"D6",X"D7",X"97",X"CD",
		X"EF",X"99",X"CA",X"EC",X"0E",X"9D",X"D6",X"1F",X"00",X"01",X"A4",X"C9",X"F6",X"A6",X"C7",X"E9",
		X"A6",X"9B",X"D6",X"A6",X"99",X"C7",X"A9",X"CB",X"F4",X"A9",X"9B",X"D4",X"AB",X"C9",X"EB",X"D4",
		X"AD",X"9B",X"C9",X"AC",X"C2",X"C3",X"AE",X"C3",X"E5",X"AE",X"CD",X"F2",X"B0",X"CB",X"ED",X"B0",
		X"9B",X"CB",X"D2",X"B1",X"C2",X"C3",X"B3",X"C5",X"CF",X"D0",X"B5",X"CD",X"F0",X"B7",X"99",X"CD",
		X"D0",X"B8",X"C2",X"C4",X"C5",X"BA",X"CD",X"F0",X"BD",X"C0",X"E7",X"02",X"9F",X"C0",X"F7",X"04",
		X"A1",X"C7",X"E9",X"A4",X"C4",X"C5",X"A7",X"C1",X"C2",X"03",X"A1",X"85",X"C6",X"A4",X"88",X"C3",
		X"A7",X"9C",X"C0",X"A4",X"9E",X"D7",X"A9",X"9E",X"D5",X"AE",X"9E",X"D3",X"B3",X"9E",X"D1",X"06",
		X"A1",X"86",X"C0",X"07",X"A2",X"CC",X"D2",X"A7",X"CC",X"D1",X"A9",X"C9",X"AA",X"C2",X"AC",X"C5",
		X"AC",X"D0",X"AE",X"CC",X"AF",X"C2",X"B1",X"C5",X"CF",X"B3",X"CD",X"B6",X"C2",X"C5",X"B8",X"CE",
		X"BB",X"C2",X"C5",X"08",X"A3",X"C8",X"A8",X"CA",X"AD",X"CB",X"B2",X"CE",X"09",X"BA",X"C3",X"0A",
		X"A6",X"C7",X"AB",X"C9",X"B0",X"CB",X"0D",X"99",X"CE",X"CF",X"1F",X"00",X"01",X"A5",X"CB",X"ED",
		X"D4",X"D5",X"A7",X"C0",X"C1",X"C6",X"E8",X"D5",X"AA",X"D1",X"F5",X"AC",X"C8",X"EE",X"AE",X"90",
		X"C8",X"AF",X"CE",X"B1",X"C3",X"EE",X"B9",X"C3",X"E6",X"BE",X"C0",X"F7",X"02",X"A5",X"D1",X"F3",
		X"A7",X"89",X"D1",X"B3",X"98",X"C3",X"C6",X"BE",X"C2",X"E5",X"C9",X"ED",X"D0",X"F3",X"D6",X"D7",
		X"04",X"A2",X"C0",X"E4",X"C9",X"F1",X"A9",X"CF",X"D0",X"AC",X"CF",X"D0",X"03",X"A5",X"C0",X"A5",
		X"9D",X"D6",X"A7",X"92",X"C2",X"B1",X"9D",X"C7",X"06",X"A1",X"84",X"D6",X"07",X"A3",X"D4",X"A5",
		X"C1",X"C6",X"C8",X"A8",X"D2",X"D4",X"AF",X"C9",X"CB",X"CD",X"B7",X"C4",X"C5",X"BC",X"C0",X"C5",
		X"CE",X"D4",X"08",X"A2",X"CC",X"D2",X"A9",X"CB",X"09",X"BB",X"CB",X"0A",X"A5",X"CB",X"AC",X"C8",
		X"BE",X"C0",X"0D",X"89",X"D2",X"F4",X"98",X"C4",X"C5",X"1F",X"00",X"01",X"A5",X"C3",X"F0",X"A7",
		X"C9",X"CD",X"AA",X"C0",X"F7",X"AC",X"C9",X"CF",X"AF",X"C6",X"F7",X"B1",X"C9",X"CD",X"C6",X"B2",
		X"C0",X"E5",X"B4",X"CA",X"F6",X"B6",X"CD",X"B7",X"C1",X"E6",X"B9",X"C6",X"F7",X"BB",X"CD",X"BE",
		X"C0",X"F7",X"02",X"89",X"C9",X"CD",X"8E",X"C9",X"CF",X"93",X"CD",X"B3",X"96",X"C6",X"B3",X"95",
		X"C9",X"B8",X"CD",X"BD",X"CD",X"04",X"A2",X"C1",X"C2",X"D2",X"F7",X"03",X"A2",X"89",X"C0",X"A5",
		X"89",X"D1",X"AA",X"91",X"C1",X"AA",X"8E",X"D4",X"AF",X"93",X"D1",X"B2",X"96",X"C3",X"B4",X"98",
		X"D7",X"B7",X"9D",X"C0",X"B9",X"9D",X"D2",X"06",X"A1",X"84",X"C3",X"07",X"A3",X"C5",X"C9",X"A8",
		X"C4",X"CB",X"CF",X"D7",X"AD",X"CB",X"D2",X"D7",X"B0",X"C2",X"B2",X"CB",X"CF",X"B5",X"C1",X"B7",
		X"C8",X"CB",X"D5",X"BC",X"C2",X"CB",X"CF",X"08",X"A2",X"CB",X"A7",X"D2",X"B1",X"D3",X"BB",X"C7",
		X"09",X"BB",X"C3",X"0A",X"BE",X"CC",X"CE",X"D7",X"1F",X"00",X"01",X"A4",X"C5",X"F2",X"A6",X"88",
		X"C5",X"CB",X"D2",X"D3",X"A9",X"C3",X"E7",X"CB",X"CF",X"F3",X"A6",X"D4",X"F6",X"AB",X"8F",X"C3",
		X"C7",X"CF",X"A6",X"94",X"D7",X"AB",X"C7",X"EF",X"D3",X"F7",X"AE",X"C1",X"E7",X"B0",X"97",X"C1",
		X"C7",X"B0",X"CD",X"F4",X"B2",X"94",X"CD",X"B3",X"9A",X"C4",X"B3",X"C5",X"C6",X"B5",X"CA",X"EE",
		X"D1",X"D5",X"F7",X"B6",X"C2",X"C3",X"B7",X"C7",X"EA",X"CE",X"D1",X"F5",X"B9",X"C4",X"E7",X"CA",
		X"CE",X"F1",X"BE",X"C0",X"F7",X"02",X"BE",X"C1",X"C3",X"C5",X"C7",X"C9",X"CB",X"CD",X"CF",X"D1",
		X"D3",X"D5",X"D7",X"04",X"AD",X"D5",X"03",X"A4",X"88",X"D1",X"A9",X"8F",X"D0",X"B0",X"94",X"CC",
		X"D6",X"B5",X"9D",X"CB",X"B5",X"98",X"D0",X"B5",X"D2",X"D4",X"06",X"A1",X"9D",X"C0",X"07",X"A7",
		X"C7",X"A9",X"C9",X"CD",X"D5",X"AC",X"C5",X"AE",X"CD",X"D4",X"B3",X"CE",X"B4",X"C2",X"B5",X"C8",
		X"D3",X"B7",X"C5",X"CF",X"BC",X"C2",X"D3",X"D7",X"08",X"A1",X"CA",X"A3",X"D4",X"AD",X"D2",X"09",
		X"BB",X"C9",X"0A",X"A4",X"C5",X"A4",X"CB",X"AE",X"C1",X"0D",X"85",X"D3",X"F7",X"8A",X"CC",X"EE",
		X"96",X"C8",X"C9",X"1F",X"00",X"01",X"A7",X"99",X"D6",X"A7",X"8E",X"D4",X"A7",X"D0",X"F3",X"A9",
		X"91",X"D0",X"AA",X"CC",X"EF",X"AC",X"94",X"CC",X"AD",X"C8",X"EB",X"D1",X"F3",X"AF",X"97",X"C8",
		X"B0",X"C4",X"E7",X"CD",X"EF",X"B2",X"9B",X"C4",X"B3",X"C0",X"E3",X"C9",X"EB",X"B5",X"9B",X"C0",
		X"B6",X"C5",X"E7",X"BA",X"C1",X"E3",X"B2",X"99",X"D3",X"B2",X"D4",X"D5",X"B8",X"D4",X"D5",X"B5",
		X"CF",X"F2",X"B7",X"CF",X"B9",X"CC",X"EF",X"BB",X"CC",X"F2",X"BD",X"C7",X"F7",X"02",X"9F",X"C0",
		X"F7",X"03",X"A7",X"9C",X"D7",X"A7",X"91",X"D5",X"A7",X"89",X"CF",X"AA",X"8C",X"CB",X"AD",X"8F",
		X"C7",X"B0",X"92",X"C3",X"B2",X"94",X"D2",X"B5",X"98",X"CE",X"B9",X"9C",X"CB",X"06",X"A1",X"86",
		X"D7",X"BD",X"C6",X"07",X"AB",X"D1",X"D3",X"AE",X"CD",X"CF",X"B1",X"C9",X"CB",X"B0",X"D4",X"B3",
		X"D0",X"B4",X"C5",X"C7",X"B7",X"CC",X"B8",X"C1",X"C3",X"B9",X"D0",X"D2",X"BB",X"D3",X"D5",X"C8",
		X"CA",X"08",X"A4",X"D2",X"A7",X"CD",X"AA",X"C9",X"BC",X"C0",X"09",X"B5",X"D4",X"0A",X"B3",X"C0",
		X"BD",X"D3",X"BA",X"C1",X"0D",X"8C",X"D1",X"F3",X"1F",X"00",X"02",X"9F",X"C0",X"F7",X"04",X"A4",
		X"C4",X"CA",X"D2",X"D6",X"A7",X"C1",X"C2",X"C5",X"C8",X"CB",X"D0",X"D3",X"D5",X"AA",X"C6",X"CC",
		X"D4",X"AD",X"C2",X"C7",X"CD",X"D0",X"D5",X"B0",X"C1",X"C6",X"C8",X"CB",X"CE",X"D4",X"D6",X"B3",
		X"C5",X"C8",X"CA",X"CD",X"CF",X"D3",X"D5",X"B6",X"C1",X"C4",X"C9",X"CC",X"D0",X"D2",X"B9",X"C2",
		X"C5",X"CB",X"D4",X"D6",X"03",X"A4",X"87",X"C3",X"D1",X"A4",X"90",X"C9",X"D7",X"A7",X"90",X"C0",
		X"A7",X"8D",X"CF",X"AD",X"99",X"C3",X"AD",X"9E",X"D1",X"B6",X"9E",X"C0",X"06",X"A1",X"86",X"C0",
		X"07",X"A5",X"CA",X"CF",X"A9",X"C2",X"D2",X"D6",X"AD",X"C6",X"B1",X"D4",X"B4",X"CF",X"BA",X"C5",
		X"D4",X"AC",X"CB",X"08",X"AA",X"CC",X"B6",X"C9",X"CC",X"D2",X"09",X"BC",X"CB",X"1F",X"00",X"01",
		X"A5",X"87",X"C2",X"C6",X"D1",X"A8",X"98",X"C2",X"F7",X"00",X"A8",X"8D",X"C8",X"AB",X"8D",X"C6",
		X"C7",X"AB",X"98",X"C5",X"AE",X"90",X"CB",X"F0",X"AE",X"D3",X"AC",X"D6",X"B5",X"97",X"CD",X"EF",
		X"B7",X"CC",X"01",X"AE",X"CD",X"EE",X"B9",X"CD",X"EE",X"BA",X"CC",X"ED",X"BC",X"9E",X"CB",X"ED",
		X"02",X"9F",X"C0",X"F7",X"04",X"A2",X"C1",X"F7",X"B9",X"D0",X"F5",X"03",X"A5",X"9E",X"C0",X"AE",
		X"9A",X"D6",X"B8",X"9A",X"CF",X"06",X"A1",X"84",X"C0",X"07",X"AF",X"CB",X"D0",X"AE",X"D3",X"08",
		X"A5",X"C9",X"CC",X"AB",X"C7",X"BC",X"D2",X"09",X"B5",X"CE",X"0A",X"A8",X"D0",X"AE",X"C6",X"BC",
		X"CB",X"0E",X"90",X"CB",X"CC",X"CF",X"D0",X"8F",X"D3",X"99",X"CC",X"1F",X"00",X"01",X"A8",X"95",
		X"C0",X"EA",X"A8",X"CC",X"EF",X"AD",X"CB",X"F6",X"B4",X"D1",X"F6",X"B9",X"C0",X"ED",X"BB",X"C5",
		X"BC",X"CE",X"BE",X"C0",X"F7",X"00",X"B0",X"93",X"C2",X"E4",X"B3",X"95",X"C9",X"AF",X"95",X"CA",
		X"04",X"A3",X"C1",X"EE",X"A5",X"D0",X"F6",X"B1",X"CA",X"F0",X"03",X"A2",X"87",X"C0",X"CF",X"A8",
		X"8A",X"CB",X"AA",X"8E",X"CA",X"AE",X"92",X"C9",X"B2",X"95",X"C8",X"B9",X"9D",X"C6",X"CC",X"A5",
		X"9D",X"D7",X"06",X"A1",X"84",X"D7",X"07",X"A8",X"D0",X"D2",X"D4",X"B2",X"C2",X"C4",X"B7",X"C2",
		X"08",X"AA",X"CE",X"D3",X"B1",X"D3",X"BB",X"D3",X"09",X"BB",X"C9",X"0A",X"B9",X"C0",X"BE",X"C4",
		X"BE",X"CD",X"0F",X"9D",X"C0",X"E4",X"1F",X"00",X"01",X"A8",X"C9",X"EC",X"D1",X"F4",X"AC",X"C1",
		X"E7",X"AD",X"CE",X"F6",X"B6",X"C1",X"E7",X"B9",X"C9",X"F4",X"A5",X"8A",X"C1",X"AE",X"92",X"C1",
		X"B8",X"9D",X"C1",X"B8",X"C7",X"A5",X"87",X"C9",X"CC",X"B1",X"98",X"C9",X"AF",X"9C",X"D6",X"02",
		X"B1",X"C2",X"E8",X"BE",X"C0",X"F7",X"BA",X"9D",X"C7",X"04",X"A2",X"C1",X"E8",X"CF",X"F6",X"A5",
		X"C2",X"E8",X"AA",X"C9",X"ED",X"B2",X"CB",X"F5",X"03",X"A5",X"9D",X"C0",X"AC",X"90",X"C2",X"A9",
		X"8D",X"C8",X"B1",X"98",X"CA",X"B9",X"9D",X"D5",X"A5",X"9A",X"D7",X"06",X"A1",X"84",X"D7",X"07",
		X"A4",X"D0",X"D5",X"A6",X"CA",X"D2",X"A8",X"C3",X"C5",X"B5",X"CD",X"D2",X"B8",X"C6",X"BC",X"CD",
		X"08",X"A5",X"D4",X"AA",X"D3",X"AE",X"C5",X"BB",X"D0",X"09",X"B3",X"C5",X"0A",X"A8",X"D1",X"B6",
		X"C4",X"B6",X"C7",X"0D",X"87",X"CA",X"CB",X"0F",X"9D",X"C2",X"E6",X"D7",X"1F",X"01",X"01",X"A8",
		X"95",X"C0",X"E5",X"D1",X"F7",X"AA",X"95",X"C8",X"EE",X"A5",X"C8",X"EE",X"B9",X"C1",X"E5",X"C8",
		X"EE",X"D1",X"F6",X"BE",X"C0",X"F7",X"A2",X"84",X"CB",X"00",X"AE",X"91",X"C1",X"C2",X"D6",X"D7",
		X"B4",X"C4",X"D2",X"D3",X"CB",X"04",X"A2",X"C0",X"E5",X"D1",X"F7",X"A7",X"C8",X"EE",X"03",X"A5",
		X"9A",X"C6",X"D0",X"B9",X"9D",X"C0",X"D7",X"06",X"A1",X"84",X"C6",X"D0",X"07",X"A3",X"C0",X"D7",
		X"B0",X"C2",X"D6",X"B4",X"C4",X"CB",X"D2",X"D3",X"BC",X"C4",X"D3",X"08",X"A7",X"CB",X"B6",X"CA",
		X"CC",X"09",X"BB",X"CB",X"0A",X"B9",X"C9",X"CB",X"CD",X"0E",X"91",X"C1",X"C2",X"D6",X"D7",X"1F",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"02",X"C0",X"02",X"C1",X"C4",X"06",X"C2",X"04",X"08",X"08",X"08",X"08",X"0C",X"00",X"00",X"00",
		X"C8",X"C6",X"10",X"00",X"0C",X"0E",X"0C",X"0E",X"00",X"00",X"00",X"00",X"0A",X"CA",X"CA",X"02",
		X"CA",X"0A",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C4",X"06",X"C2",X"04",
		X"20",X"AC",X"20",X"AE",X"00",X"00",X"00",X"00",X"16",X"16",X"16",X"16",X"1C",X"1E",X"1C",X"1E",
		X"B4",X"00",X"00",X"00",X"B4",X"B5",X"B4",X"B5",X"16",X"18",X"1A",X"20",X"18",X"1A",X"20",X"20",
		X"1A",X"18",X"16",X"16",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"14",X"12",X"B0",X"B2",
		X"A0",X"9C",X"9E",X"A0",X"00",X"00",X"00",X"00",X"A6",X"A6",X"A6",X"A6",X"A1",X"A0",X"A1",X"A0",
		X"A0",X"00",X"00",X"00",X"A0",X"A1",X"A0",X"A1",X"A6",X"A6",X"A0",X"A0",X"A6",X"A6",X"A6",X"A0",
		X"A6",X"A6",X"A6",X"A6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A2",X"38",X"A4",X"36",
		X"92",X"90",X"8E",X"00",X"00",X"00",X"00",X"00",X"3A",X"3A",X"3A",X"3A",X"98",X"99",X"98",X"99",
		X"99",X"00",X"00",X"00",X"98",X"99",X"98",X"99",X"98",X"99",X"92",X"92",X"3C",X"3C",X"3C",X"3C",
		X"3C",X"3C",X"3C",X"3A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"94",X"96",X"94",X"96",
		X"B6",X"BA",X"B6",X"BA",X"E6",X"E8",X"EA",X"EC",X"22",X"22",X"22",X"22",X"24",X"24",X"24",X"24",
		X"EE",X"00",X"00",X"00",X"EE",X"EF",X"EE",X"EF",X"E4",X"E2",X"B6",X"B6",X"E2",X"E4",X"B6",X"B6",
		X"E4",X"E2",X"22",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DD",X"DE",X"DF",X"DE",X"00",X"00",X"00",X"00",X"DE",X"A7",X"DE",X"A7",X"40",X"40",X"40",X"40",
		X"BF",X"00",X"00",X"00",X"DD",X"BF",X"DD",X"BF",X"DD",X"3E",X"BC",X"DF",X"A7",X"DE",X"A7",X"DE",
		X"DE",X"A7",X"DE",X"A7",X"DD",X"34",X"DD",X"00",X"DD",X"34",X"DD",X"DD",X"DE",X"DF",X"DE",X"DD",
		X"80",X"84",X"82",X"00",X"00",X"00",X"00",X"00",X"8A",X"8A",X"8A",X"8A",X"2A",X"2A",X"2A",X"2A",
		X"8C",X"00",X"00",X"00",X"8C",X"8D",X"8C",X"8D",X"8C",X"84",X"82",X"80",X"8A",X"8A",X"8A",X"8A",
		X"8A",X"8A",X"8A",X"8A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"86",X"28",X"88",X"26",
		X"CE",X"CC",X"CE",X"CC",X"30",X"32",X"30",X"32",X"CE",X"CF",X"CE",X"CF",X"CE",X"CF",X"CE",X"CF",
		X"CF",X"00",X"00",X"00",X"CE",X"CF",X"CE",X"CF",X"CE",X"CF",X"CE",X"CF",X"CE",X"CF",X"CE",X"CF",
		X"CE",X"CF",X"CE",X"CF",X"2C",X"2E",X"30",X"00",X"2E",X"2C",X"CE",X"00",X"00",X"00",X"00",X"00",
		X"D0",X"D1",X"D0",X"D1",X"00",X"00",X"00",X"00",X"D4",X"D4",X"D4",X"D4",X"D4",X"D4",X"D4",X"D4",
		X"D8",X"00",X"00",X"00",X"D4",X"D4",X"D4",X"D4",X"D8",X"D0",X"D1",X"00",X"D4",X"D4",X"D4",X"D4",
		X"D4",X"D4",X"D4",X"D4",X"D1",X"DB",X"D9",X"D5",X"D5",X"D9",X"DB",X"D1",X"D5",X"D7",X"D5",X"D7",
		X"00",X"00",X"00",X"00",X"41",X"40",X"41",X"40",X"00",X"40",X"00",X"40",X"00",X"00",X"00",X"00",
		X"01",X"01",X"00",X"00",X"00",X"00",X"40",X"40",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"41",X"40",X"41",X"40",
		X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"40",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"41",X"41",
		X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"40",X"00",X"00",X"40",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"40",X"40",X"00",X"00",X"00",X"40",X"00",X"00",
		X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"41",X"40",X"41",X"40",
		X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"40",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"40",X"00",X"00",
		X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"41",X"41",X"41",X"41",
		X"01",X"01",X"01",X"01",X"41",X"41",X"41",X"41",X"00",X"40",X"00",X"40",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"00",X"00",X"40",X"00",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"01",X"01",X"00",X"00",X"40",X"40",
		X"00",X"00",X"40",X"40",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"81",X"80",X"80",
		X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"41",X"01",X"41",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"41",X"01",X"01",
		X"01",X"41",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"41",X"40",X"41",X"40",
		X"40",X"41",X"40",X"41",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"40",X"00",X"00",X"40",X"40",
		X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"40",X"00",X"00",X"01",X"00",X"00",X"40",X"00",X"40",
		X"00",X"40",X"00",X"40",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"01",X"00",
		X"FE",X"00",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FE",X"00",
		X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"F5",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FA",X"FC",X"F5",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"F8",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"FC",X"FC",X"FC",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"01",X"FF",X"FF",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"00",X"FE",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FD",X"FD",X"FD",X"00",X"00",X"00",X"00",X"00",X"F8",X"08",X"F8",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FD",X"FD",X"FD",X"F8",X"08",X"F8",X"F8",
		X"F8",X"08",X"F8",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FC",X"00",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FC",X"F8",X"F8",X"FC",X"FC",X"F8",X"F8",X"FC",X"FC",X"00",X"FC",X"00",
		X"00",X"00",X"00",X"00",X"FD",X"00",X"FD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"00",
		X"10",X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"FD",X"00",X"FD",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FE",
		X"00",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"00",X"01",X"00",
		X"10",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"04",X"04",X"04",
		X"02",X"02",X"02",X"02",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"00",
		X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"10",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",
		X"10",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"04",X"00",
		X"10",X"10",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"10",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"00",X"FF",X"00",X"FF",X"F8",X"00",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",
		X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"00",X"F8",X"00",
		X"00",X"FC",X"00",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"00",X"08",X"09",X"00",X"00",
		X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"00",X"F8",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"04",X"04",X"07",X"07",
		X"04",X"04",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"F8",X"F8",X"F8",
		X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F9",X"FD",X"FC",X"FC",X"FD",X"FD",X"FC",X"00",
		X"FD",X"FD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"00",X"F8",X"00",X"00",X"00",X"F9",X"F9",X"F9",X"F9",
		X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"FF",X"00",X"00",X"00",X"03",X"03",
		X"00",X"00",X"FD",X"FD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"08",X"F8",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"F8",X"F8",X"FC",X"00",X"00",X"F8",X"F9",X"F8",X"F9",
		X"00",X"00",X"00",X"00",X"08",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"08",X"00",
		X"00",X"04",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"08",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"05",X"05",X"05",
		X"04",X"04",X"04",X"04",X"FC",X"FC",X"FC",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"07",X"04",X"04",X"07",X"07",X"04",X"00",
		X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"0C",X"07",X"01",X"08",X"07",X"01",X"00",X"08",X"07",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"06",X"06",X"06",X"06",X"08",X"08",X"08",X"01",X"0A",X"06",X"00",X"00",
		X"0A",X"06",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"08",X"09",X"07",
		X"08",X"08",X"01",X"00",X"06",X"06",X"06",X"01",X"06",X"06",X"06",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"05",X"04",X"03",X"03",X"08",X"08",X"01",X"00",X"06",X"06",X"06",X"00",
		X"06",X"06",X"06",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"04",X"03",X"04",
		X"08",X"08",X"01",X"00",X"0A",X"06",X"00",X"00",X"0A",X"06",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"06",X"06",X"04",X"05",X"05",X"05",X"05",
		X"05",X"05",X"05",X"05",X"06",X"08",X"04",X"00",X"06",X"08",X"04",X"00",X"04",X"03",X"04",X"04",
		X"08",X"08",X"04",X"00",X"06",X"06",X"06",X"00",X"06",X"06",X"06",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"05",X"05",X"05",X"05",X"08",X"08",X"08",X"02",X"05",X"05",X"05",X"00",
		X"05",X"05",X"05",X"00",X"04",X"04",X"04",X"00",X"04",X"04",X"04",X"00",X"00",X"00",X"00",X"00",
		X"08",X"0C",X"08",X"00",X"05",X"05",X"05",X"00",X"05",X"05",X"05",X"00",X"04",X"04",X"04",X"04",
		X"04",X"04",X"04",X"04",X"05",X"05",X"05",X"05",X"43",X"03",X"20",X"FF",X"A3",X"FF",X"A3",X"FF",
		X"A2",X"FF",X"A2",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"83",X"83",X"A3",X"FF",X"A3",X"A3",X"FF",X"FF",X"A2",X"A2",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"43",X"A0",X"FF",X"FF",X"A3",X"A3",X"A3",X"FF",
		X"A2",X"A2",X"A2",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"43",X"A0",X"FF",X"FF",X"A3",X"A3",X"A3",X"FF",X"A2",X"A2",X"A2",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"43",X"A0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"A2",X"A2",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"83",X"20",X"20",X"A3",X"A3",X"A3",X"A3",X"A2",X"A2",X"A2",X"A2",X"FF",X"FF",X"FF",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"43",X"A0",X"A0",X"FF",X"A3",X"A3",X"A3",X"FF",
		X"A2",X"A2",X"A2",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"23",X"20",X"20",X"23",X"23",X"23",X"FF",X"22",X"22",X"22",X"FF",X"FF",X"FF",X"FF",X"00",
		X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"03",X"20",X"FF",X"23",X"23",X"23",X"FF",
		X"22",X"22",X"22",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"06",X"07",X"06",X"00",X"04",X"04",X"02",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"06",X"07",X"08",
		X"00",X"05",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"05",X"04",X"02",X"00",X"05",X"05",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"03",X"03",
		X"00",X"08",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"02",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"04",X"00",X"00",X"04",X"04",X"00",X"04",
		X"00",X"05",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"04",X"04",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"00",X"00",X"03",X"03",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"04",
		X"00",X"04",X"00",X"04",X"04",X"04",X"04",X"04",X"00",X"00",X"00",X"00",X"FC",X"FA",X"00",X"00",
		X"02",X"06",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"F8",X"F8",X"00",X"FA",X"F7",X"00",X"00",X"01",X"07",X"07",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"00",X"00",X"FC",X"FC",X"FC",X"FC",
		X"04",X"04",X"04",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"F8",X"00",X"00",X"FC",X"FC",X"F9",X"00",X"04",X"04",X"04",X"04",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"00",X"00",X"F8",X"F9",X"00",X"00",
		X"00",X"08",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"F8",X"F8",X"FC",X"FC",X"FC",X"FC",X"04",X"04",X"04",X"04",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"00",X"00",X"FC",X"FC",X"F9",X"00",
		X"04",X"04",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"02",X"51",X"01",X"01",X"00",X"03",X"92",X"D4",X"01",X"01",X"18",X"03",X"0F",X"D0",X"D5",X"CF",
		X"D2",X"01",X"02",X"18",X"03",X"0E",X"D0",X"D1",X"D5",X"D3",X"01",X"03",X"18",X"03",X"0C",X"D0",
		X"D1",X"D2",X"D4",X"D5",X"D3",X"01",X"04",X"18",X"03",X"0A",X"D0",X"D1",X"D2",X"D4",X"D4",X"D4",
		X"D5",X"D3",X"01",X"05",X"27",X"D5",X"D3",X"01",X"06",X"27",X"D5",X"D3",X"01",X"07",X"28",X"D3",
		X"01",X"08",X"28",X"D3",X"01",X"09",X"27",X"D5",X"D3",X"01",X"0A",X"27",X"D5",X"D3",X"01",X"0B",
		X"27",X"D5",X"D3",X"01",X"0C",X"27",X"D5",X"D3",X"01",X"0D",X"27",X"D5",X"D3",X"01",X"0E",X"27",
		X"D5",X"D3",X"01",X"0F",X"27",X"D5",X"D3",X"01",X"10",X"27",X"D5",X"D3",X"01",X"11",X"27",X"D5",
		X"D3",X"01",X"12",X"27",X"D5",X"D3",X"02",X"53",X"01",X"07",X"26",X"CA",X"01",X"08",X"25",X"CB",
		X"CC",X"02",X"54",X"01",X"07",X"27",X"CD",X"01",X"08",X"27",X"CE",X"02",X"52",X"01",X"05",X"18",
		X"03",X"0A",X"EB",X"01",X"06",X"18",X"03",X"0A",X"EB",X"01",X"07",X"18",X"03",X"08",X"EC",X"ED",
		X"EB",X"01",X"08",X"18",X"03",X"08",X"5C",X"EE",X"EB",X"01",X"09",X"1E",X"5C",X"5C",X"EE",X"EB",
		X"01",X"0A",X"1E",X"5C",X"5C",X"EE",X"EB",X"01",X"0B",X"1E",X"5C",X"5C",X"EE",X"EB",X"01",X"0C",
		X"1E",X"5C",X"5C",X"EE",X"EB",X"01",X"0D",X"1E",X"5C",X"5C",X"EE",X"EB",X"01",X"0E",X"1E",X"5C",
		X"5C",X"EE",X"EB",X"01",X"0F",X"1E",X"5C",X"5C",X"EE",X"EB",X"01",X"10",X"1E",X"5C",X"5C",X"EE",
		X"EB",X"01",X"11",X"1E",X"5C",X"5C",X"EE",X"EB",X"01",X"12",X"1E",X"5C",X"5C",X"EE",X"EB",X"01",
		X"13",X"1C",X"FD",X"EF",X"F0",X"F1",X"F2",X"F3",X"01",X"14",X"18",X"03",X"04",X"F8",X"F7",X"F6",
		X"F4",X"F5",X"01",X"15",X"18",X"03",X"05",X"F8",X"F7",X"F6",X"F6",X"EF",X"FC",X"01",X"16",X"18",
		X"03",X"06",X"F8",X"F7",X"F6",X"F6",X"F4",X"F5",X"01",X"17",X"18",X"03",X"07",X"F8",X"F7",X"F6",
		X"F6",X"F6",X"EF",X"FC",X"01",X"18",X"18",X"03",X"08",X"F8",X"F7",X"F6",X"F6",X"F6",X"F4",X"F5",
		X"01",X"19",X"18",X"03",X"09",X"F8",X"F7",X"03",X"04",X"F6",X"EF",X"F9",X"01",X"1A",X"18",X"03",
		X"0A",X"F8",X"F7",X"03",X"04",X"F6",X"F4",X"F5",X"01",X"1B",X"18",X"03",X"0B",X"F8",X"F7",X"03",
		X"05",X"F6",X"EF",X"FC",X"01",X"1C",X"18",X"03",X"0C",X"F8",X"F7",X"03",X"05",X"F6",X"F4",X"F5",
		X"01",X"1D",X"18",X"03",X"0D",X"F8",X"F7",X"03",X"06",X"F6",X"EF",X"FC",X"01",X"1E",X"18",X"03",
		X"0E",X"F8",X"F7",X"03",X"06",X"F6",X"F4",X"F5",X"01",X"1F",X"18",X"03",X"0F",X"F8",X"F7",X"03",
		X"07",X"F6",X"EF",X"02",X"10",X"01",X"09",X"18",X"03",X"06",X"04",X"01",X"0A",X"18",X"03",X"06",
		X"04",X"01",X"0B",X"18",X"03",X"06",X"04",X"01",X"0C",X"18",X"03",X"06",X"04",X"01",X"0D",X"18",
		X"03",X"06",X"04",X"01",X"0E",X"18",X"03",X"06",X"04",X"01",X"0F",X"18",X"03",X"06",X"04",X"01",
		X"10",X"18",X"03",X"06",X"04",X"01",X"11",X"18",X"03",X"06",X"04",X"01",X"12",X"18",X"03",X"06",
		X"04",X"01",X"13",X"18",X"03",X"04",X"04",X"02",X"55",X"01",X"13",X"22",X"03",X"05",X"94",X"D5",
		X"FA",X"03",X"07",X"94",X"01",X"14",X"20",X"03",X"07",X"94",X"D5",X"FA",X"03",X"07",X"94",X"01",
		X"15",X"22",X"03",X"05",X"94",X"D5",X"FA",X"03",X"07",X"94",X"01",X"16",X"23",X"03",X"04",X"94",
		X"D5",X"FA",X"03",X"07",X"94",X"01",X"17",X"25",X"94",X"D6",X"D7",X"D8",X"D9",X"03",X"06",X"94",
		X"01",X"18",X"26",X"DA",X"DB",X"DC",X"DD",X"DE",X"03",X"05",X"94",X"01",X"19",X"28",X"E0",X"E1",
		X"E2",X"E3",X"E4",X"94",X"94",X"94",X"01",X"1A",X"29",X"94",X"94",X"E5",X"E6",X"E3",X"E4",X"94",
		X"01",X"1B",X"2B",X"94",X"94",X"E5",X"E6",X"E3",X"01",X"1C",X"2C",X"94",X"94",X"94",X"E5",X"01",
		X"1D",X"2E",X"94",X"94",X"01",X"1E",X"2F",X"94",X"00",X"4C",X"0C",X"99",X"00",X"4E",X"0C",X"99",
		X"10",X"50",X"0C",X"99",X"20",X"52",X"0C",X"79",X"00",X"54",X"0C",X"79",X"10",X"A8",X"0C",X"79",
		X"20",X"A8",X"0C",X"89",X"20",X"70",X"0C",X"59",X"00",X"72",X"0C",X"59",X"10",X"74",X"0C",X"59",
		X"20",X"76",X"4C",X"7D",X"00",X"00",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"21",X"2A",X"5C",X"A7",X"28",X"03",X"21",X"5C",X"5C",X"7E",X"32",X"DB",X"E5",X"23",X"22",X"DC",
		X"E5",X"C9",X"21",X"DB",X"E5",X"35",X"2A",X"DC",X"E5",X"20",X"0D",X"7E",X"3C",X"28",X"09",X"23",
		X"7E",X"32",X"DB",X"E5",X"23",X"22",X"DC",X"E5",X"7E",X"C9",X"0C",X"02",X"78",X"80",X"14",X"02",
		X"32",X"80",X"24",X"08",X"32",X"02",X"23",X"20",X"32",X"01",X"5A",X"02",X"1E",X"20",X"0C",X"02",
		X"1E",X"20",X"0C",X"02",X"5A",X"20",X"73",X"01",X"24",X"08",X"5A",X"01",X"24",X"08",X"64",X"01",
		X"32",X"04",X"5F",X"02",X"23",X"20",X"14",X"80",X"1E",X"08",X"FF",X"FF",X"8C",X"01",X"DC",X"08",
		X"19",X"02",X"19",X"01",X"14",X"80",X"14",X"04",X"14",X"80",X"4A",X"02",X"C8",X"01",X"EB",X"02",
		X"6E",X"80",X"37",X"02",X"50",X"01",X"14",X"80",X"0A",X"01",X"0A",X"02",X"0F",X"01",X"0A",X"02",
		X"05",X"01",X"0A",X"02",X"28",X"08",X"FF",X"FF",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"3E",X"13",X"CD",X"42",X"31",X"CD",X"5E",X"5F",X"3E",X"01",X"32",X"AE",X"E6",X"18",X"04",X"AF",
		X"32",X"AE",X"E6",X"3A",X"90",X"E5",X"FE",X"00",X"20",X"05",X"3E",X"20",X"CD",X"42",X"31",X"CD",
		X"C9",X"5E",X"3A",X"B7",X"E5",X"B7",X"28",X"35",X"3A",X"AE",X"E6",X"B7",X"20",X"2F",X"CD",X"D6",
		X"5E",X"3E",X"02",X"32",X"88",X"E5",X"3E",X"0E",X"CD",X"3E",X"30",X"21",X"2E",X"D6",X"36",X"00",
		X"54",X"5D",X"13",X"01",X"27",X"00",X"ED",X"B0",X"3E",X"0E",X"CD",X"3E",X"30",X"CD",X"D6",X"5E",
		X"21",X"88",X"E5",X"35",X"20",X"E0",X"3E",X"70",X"CD",X"3E",X"30",X"18",X"35",X"3A",X"90",X"E5",
		X"FE",X"00",X"21",X"36",X"D6",X"CC",X"9A",X"31",X"3E",X"02",X"32",X"88",X"E5",X"3E",X"0E",X"CD",
		X"3E",X"30",X"21",X"32",X"D7",X"36",X"00",X"54",X"5D",X"13",X"01",X"1B",X"00",X"ED",X"B0",X"3E",
		X"0E",X"CD",X"3E",X"30",X"CD",X"C9",X"5E",X"21",X"88",X"E5",X"35",X"20",X"E0",X"3E",X"38",X"CD",
		X"3E",X"30",X"3E",X"01",X"32",X"90",X"E5",X"3A",X"8E",X"E5",X"3D",X"CD",X"EC",X"31",X"79",X"3C",
		X"32",X"CC",X"E5",X"79",X"E6",X"07",X"3C",X"32",X"CD",X"E5",X"21",X"00",X"00",X"22",X"8A",X"E5",
		X"22",X"8B",X"E5",X"21",X"6C",X"E5",X"FE",X"01",X"20",X"09",X"36",X"30",X"3E",X"60",X"32",X"8B",
		X"E5",X"18",X"14",X"FE",X"02",X"20",X"09",X"36",X"40",X"3E",X"80",X"32",X"8B",X"E5",X"18",X"07",
		X"36",X"50",X"3E",X"01",X"32",X"8A",X"E5",X"79",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"21",X"DF",
		X"E5",X"86",X"87",X"5F",X"16",X"00",X"21",X"35",X"5F",X"19",X"5E",X"23",X"56",X"ED",X"53",X"E1",
		X"E5",X"3E",X"14",X"CD",X"42",X"31",X"CD",X"80",X"61",X"CD",X"D7",X"63",X"AF",X"32",X"A6",X"E5",
		X"CD",X"43",X"5F",X"CD",X"E7",X"62",X"21",X"10",X"D0",X"11",X"ED",X"5E",X"CD",X"2D",X"30",X"CD",
		X"03",X"32",X"0E",X"1E",X"21",X"4A",X"D0",X"3A",X"8E",X"E5",X"CD",X"48",X"30",X"CD",X"F7",X"31",
		X"0E",X"04",X"11",X"97",X"E5",X"21",X"60",X"D0",X"3A",X"B8",X"E5",X"B7",X"28",X"03",X"21",X"18",
		X"D0",X"06",X"03",X"CD",X"5F",X"30",X"10",X"FB",X"0E",X"06",X"11",X"9A",X"E5",X"21",X"38",X"D0",
		X"06",X"03",X"CD",X"5F",X"30",X"10",X"FB",X"3A",X"B4",X"E6",X"FE",X"0C",X"20",X"14",X"21",X"BA",
		X"E1",X"06",X"07",X"36",X"0D",X"23",X"23",X"23",X"36",X"0D",X"11",X"15",X"00",X"19",X"10",X"F3",
		X"18",X"0C",X"FE",X"10",X"20",X"08",X"3E",X"01",X"32",X"FF",X"E4",X"32",X"00",X"E5",X"3A",X"A7",
		X"E5",X"B7",X"20",X"43",X"3A",X"AE",X"E6",X"B7",X"20",X"10",X"3A",X"B7",X"E5",X"B7",X"28",X"0A",
		X"3E",X"16",X"32",X"B6",X"E5",X"3E",X"18",X"32",X"AD",X"E6",X"3E",X"01",X"32",X"9D",X"E5",X"21",
		X"4A",X"E4",X"06",X"0A",X"78",X"C6",X"02",X"E6",X"03",X"20",X"05",X"3E",X"17",X"CD",X"42",X"31",
		X"7E",X"FE",X"FF",X"20",X"04",X"36",X"12",X"18",X"02",X"36",X"FF",X"3E",X"09",X"CD",X"3E",X"30",
		X"10",X"E2",X"3E",X"26",X"CD",X"42",X"31",X"3E",X"02",X"32",X"9D",X"E5",X"3E",X"15",X"32",X"B1",
		X"E6",X"3E",X"01",X"32",X"68",X"E5",X"C3",X"29",X"00",X"21",X"32",X"D7",X"CD",X"85",X"31",X"11",
		X"23",X"5F",X"CD",X"2D",X"30",X"C9",X"0E",X"06",X"3A",X"B8",X"E5",X"C6",X"31",X"21",X"2E",X"D6",
		X"CD",X"6A",X"30",X"11",X"2B",X"5F",X"CD",X"2D",X"30",X"CD",X"9A",X"31",X"C9",X"06",X"20",X"31",
		X"50",X"2D",X"20",X"20",X"20",X"20",X"20",X"20",X"1E",X"3C",X"31",X"30",X"30",X"30",X"30",X"3E",
		X"06",X"48",X"49",X"2D",X"20",X"20",X"20",X"20",X"20",X"20",X"1E",X"3C",X"52",X"2D",X"20",X"20",
		X"20",X"5E",X"5F",X"2D",X"20",X"3E",X"06",X"32",X"50",X"2D",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"00",X"06",X"20",X"52",X"45",X"41",X"44",X"59",X"00",X"06",X"2D",X"50",X"4C",X"41",
		X"59",X"45",X"52",X"20",X"00",X"98",X"00",X"04",X"01",X"10",X"01",X"14",X"01",X"17",X"01",X"21",
		X"01",X"26",X"01",X"3E",X"01",X"32",X"74",X"E5",X"AF",X"32",X"73",X"E5",X"CD",X"91",X"5F",X"3E",
		X"02",X"CD",X"3E",X"30",X"21",X"73",X"E5",X"34",X"7E",X"FE",X"1E",X"38",X"EF",X"C9",X"DD",X"21",
		X"00",X"E3",X"06",X"10",X"DD",X"36",X"04",X"00",X"DD",X"36",X"0C",X"00",X"11",X"10",X"00",X"DD",
		X"19",X"10",X"F1",X"AF",X"32",X"74",X"E5",X"32",X"A6",X"E5",X"3E",X"1C",X"32",X"73",X"E5",X"CD",
		X"91",X"5F",X"3E",X"02",X"CD",X"3E",X"30",X"21",X"73",X"E5",X"35",X"7E",X"FE",X"FF",X"20",X"EF",
		X"C9",X"87",X"4F",X"AF",X"47",X"91",X"57",X"CB",X"21",X"78",X"E6",X"03",X"CC",X"AD",X"5F",X"7A",
		X"CB",X"7F",X"20",X"02",X"0D",X"91",X"04",X"80",X"57",X"79",X"B8",X"30",X"EC",X"C5",X"D5",X"CB",
		X"38",X"CB",X"38",X"30",X"01",X"04",X"CB",X"39",X"CB",X"39",X"30",X"01",X"0C",X"2E",X"10",X"CD",
		X"D2",X"5F",X"3A",X"74",X"E5",X"B7",X"28",X"03",X"0D",X"18",X"01",X"0C",X"CD",X"D2",X"5F",X"D1",
		X"C1",X"C9",X"51",X"3E",X"18",X"80",X"FE",X"30",X"DC",X"F1",X"5F",X"3E",X"18",X"90",X"D4",X"F1",
		X"5F",X"50",X"3E",X"18",X"81",X"FE",X"30",X"DC",X"F1",X"5F",X"3E",X"18",X"91",X"D4",X"F1",X"5F",
		X"C9",X"67",X"7D",X"82",X"FE",X"20",X"DC",X"00",X"60",X"7D",X"92",X"D8",X"CD",X"00",X"60",X"C9",
		X"C5",X"D5",X"E5",X"6F",X"3A",X"A6",X"E5",X"B7",X"C2",X"3C",X"61",X"7C",X"CB",X"3F",X"CB",X"12",
		X"67",X"22",X"D6",X"E5",X"CD",X"D5",X"62",X"7E",X"FE",X"01",X"20",X"08",X"3A",X"D8",X"E5",X"47",
		X"0E",X"1F",X"18",X"11",X"FE",X"02",X"20",X"08",X"3A",X"D9",X"E5",X"47",X"0E",X"1D",X"18",X"05",
		X"CD",X"55",X"60",X"0E",X"05",X"2A",X"D6",X"E5",X"7C",X"D5",X"CD",X"00",X"2D",X"D1",X"CB",X"42",
		X"28",X"02",X"2C",X"2C",X"3A",X"74",X"E5",X"B7",X"20",X"04",X"06",X"04",X"0E",X"00",X"70",X"2C",
		X"71",X"E1",X"D1",X"C1",X"C9",X"FE",X"07",X"38",X"01",X"AF",X"FE",X"03",X"38",X"02",X"3D",X"3D",
		X"47",X"3A",X"D6",X"E5",X"B7",X"C8",X"3A",X"D7",X"E5",X"B7",X"28",X"0C",X"2B",X"7E",X"FE",X"07",
		X"38",X"01",X"AF",X"FE",X"02",X"38",X"01",X"3D",X"4F",X"2A",X"D6",X"E5",X"2D",X"7C",X"C5",X"CD",
		X"D5",X"62",X"C1",X"7E",X"FE",X"04",X"38",X"01",X"AF",X"FE",X"02",X"38",X"01",X"3D",X"5F",X"3A",
		X"D7",X"E5",X"B7",X"28",X"0C",X"2B",X"7E",X"FE",X"04",X"38",X"01",X"AF",X"FE",X"02",X"38",X"01",
		X"3D",X"6F",X"CB",X"42",X"28",X"0D",X"78",X"87",X"80",X"83",X"4F",X"06",X"00",X"21",X"C7",X"60",
		X"09",X"46",X"C9",X"78",X"87",X"80",X"83",X"5F",X"87",X"83",X"85",X"87",X"87",X"81",X"4F",X"06",
		X"00",X"21",X"D0",X"60",X"09",X"46",X"C9",X"00",X"03",X"00",X"14",X"15",X"14",X"18",X"1B",X"18",
		X"00",X"02",X"00",X"00",X"03",X"03",X"03",X"03",X"00",X"02",X"00",X"00",X"01",X"03",X"01",X"01",
		X"03",X"03",X"03",X"03",X"01",X"03",X"01",X"01",X"00",X"02",X"00",X"00",X"03",X"03",X"03",X"03",
		X"00",X"02",X"00",X"00",X"10",X"12",X"10",X"10",X"13",X"13",X"13",X"13",X"10",X"12",X"10",X"10",
		X"11",X"13",X"11",X"11",X"13",X"13",X"13",X"13",X"11",X"13",X"11",X"11",X"10",X"12",X"10",X"10",
		X"13",X"13",X"13",X"13",X"10",X"12",X"10",X"10",X"18",X"1A",X"18",X"18",X"1B",X"1B",X"1B",X"1B",
		X"18",X"1A",X"18",X"18",X"19",X"1B",X"19",X"19",X"1B",X"1B",X"1B",X"1B",X"19",X"1B",X"19",X"19",
		X"18",X"1A",X"18",X"18",X"1B",X"1B",X"1B",X"1B",X"18",X"1A",X"18",X"18",X"7C",X"CB",X"3F",X"CB",
		X"12",X"67",X"E5",X"CD",X"D5",X"62",X"7E",X"E1",X"CB",X"42",X"20",X"04",X"0F",X"0F",X"0F",X"0F",
		X"E6",X"0F",X"4F",X"42",X"7C",X"CD",X"00",X"2D",X"2C",X"CB",X"40",X"28",X"02",X"2C",X"2C",X"7E",
		X"B1",X"77",X"E6",X"C0",X"20",X"0A",X"2D",X"7E",X"FE",X"04",X"20",X"02",X"36",X"00",X"18",X"0C",
		X"FE",X"40",X"20",X"08",X"2D",X"7E",X"FE",X"FD",X"20",X"02",X"36",X"FB",X"E1",X"D1",X"C1",X"C9",
		X"21",X"00",X"E0",X"54",X"5D",X"13",X"36",X"00",X"01",X"68",X"05",X"ED",X"B0",X"ED",X"5F",X"CD",
		X"EC",X"31",X"32",X"70",X"E5",X"FD",X"21",X"58",X"E4",X"3A",X"8E",X"E5",X"FE",X"19",X"38",X"04",
		X"D6",X"18",X"18",X"F8",X"32",X"B4",X"E6",X"6F",X"26",X"00",X"29",X"EB",X"21",X"00",X"34",X"19",
		X"5E",X"23",X"56",X"1A",X"32",X"AF",X"E6",X"13",X"AF",X"32",X"7A",X"E5",X"1A",X"CB",X"7F",X"20",
		X"07",X"FE",X"1F",X"C8",X"32",X"7A",X"E5",X"13",X"1A",X"CB",X"7F",X"28",X"EF",X"CB",X"77",X"28",
		X"03",X"13",X"18",X"F4",X"3E",X"01",X"32",X"79",X"E5",X"1A",X"E6",X"1F",X"32",X"78",X"E5",X"32",
		X"77",X"E5",X"1A",X"CB",X"6F",X"28",X"09",X"3E",X"02",X"32",X"79",X"E5",X"21",X"77",X"E5",X"34",
		X"AF",X"32",X"75",X"E5",X"13",X"1A",X"E6",X"C0",X"FE",X"80",X"20",X"10",X"1A",X"E6",X"1F",X"32",
		X"77",X"E5",X"21",X"78",X"E5",X"96",X"3C",X"32",X"79",X"E5",X"18",X"E8",X"1A",X"E6",X"C0",X"FE",
		X"C0",X"20",X"B5",X"1A",X"CB",X"6F",X"20",X"06",X"E6",X"1F",X"32",X"75",X"E5",X"13",X"1A",X"E6",
		X"E0",X"FE",X"E0",X"20",X"15",X"1A",X"E6",X"1F",X"32",X"76",X"E5",X"13",X"3A",X"76",X"E5",X"21",
		X"75",X"E5",X"BE",X"38",X"D7",X"CD",X"3F",X"62",X"18",X"F2",X"CD",X"3F",X"62",X"18",X"CD",X"3A",
		X"7A",X"E5",X"FE",X"04",X"28",X"7F",X"FE",X"0B",X"30",X"04",X"FE",X"07",X"30",X"42",X"FE",X"06",
		X"28",X"1D",X"3A",X"79",X"E5",X"B7",X"28",X"78",X"21",X"77",X"E5",X"4E",X"47",X"C5",X"3A",X"75",
		X"E5",X"69",X"CD",X"D5",X"62",X"C1",X"3A",X"7A",X"E5",X"77",X"0D",X"10",X"F0",X"18",X"61",X"21",
		X"FD",X"E4",X"7E",X"FE",X"04",X"30",X"59",X"34",X"47",X"87",X"80",X"4F",X"06",X"00",X"21",X"7B",
		X"E5",X"09",X"3A",X"75",X"E5",X"77",X"23",X"ED",X"4B",X"77",X"E5",X"70",X"23",X"71",X"18",X"40",
		X"FE",X"08",X"20",X"0E",X"CD",X"0B",X"63",X"01",X"18",X"00",X"FD",X"09",X"21",X"E9",X"E4",X"34",
		X"18",X"21",X"FE",X"09",X"20",X"0D",X"FD",X"E5",X"FD",X"21",X"40",X"E4",X"CD",X"0B",X"63",X"FD",
		X"E1",X"18",X"10",X"FE",X"07",X"20",X"05",X"CD",X"5A",X"63",X"18",X"07",X"FE",X"0A",X"20",X"03",
		X"CD",X"74",X"63",X"18",X"0B",X"3A",X"75",X"E5",X"2A",X"78",X"E5",X"CD",X"D5",X"62",X"36",X"04",
		X"21",X"75",X"E5",X"34",X"C9",X"26",X"00",X"29",X"29",X"29",X"44",X"4D",X"29",X"09",X"4F",X"06",
		X"00",X"09",X"01",X"00",X"E0",X"09",X"C9",X"11",X"00",X"E4",X"3A",X"FC",X"E4",X"B7",X"28",X"0D",
		X"47",X"1A",X"6F",X"13",X"1A",X"67",X"13",X"7D",X"CD",X"AA",X"2F",X"10",X"F4",X"C9",X"00",X"08",
		X"0D",X"10",X"18",X"00",X"08",X"08",X"09",X"0B",X"0B",X"0A",X"08",X"FD",X"36",X"0A",X"00",X"FE",
		X"09",X"20",X"08",X"AF",X"32",X"0C",X"E5",X"3D",X"32",X"0B",X"E5",X"3E",X"01",X"FD",X"77",X"0F",
		X"FD",X"77",X"10",X"3A",X"75",X"E5",X"FD",X"77",X"01",X"FD",X"77",X"04",X"87",X"87",X"87",X"FD",
		X"77",X"07",X"3A",X"78",X"E5",X"FD",X"77",X"03",X"FD",X"77",X"05",X"87",X"87",X"87",X"FD",X"77",
		X"06",X"3E",X"06",X"FD",X"77",X"09",X"AF",X"FD",X"77",X"00",X"FD",X"77",X"02",X"FD",X"77",X"0A",
		X"FD",X"77",X"0C",X"FD",X"77",X"0D",X"FD",X"77",X"0E",X"C9",X"21",X"FC",X"E4",X"7E",X"FE",X"20",
		X"D0",X"34",X"87",X"4F",X"06",X"00",X"21",X"00",X"E4",X"09",X"3A",X"75",X"E5",X"77",X"23",X"3A",
		X"78",X"E5",X"77",X"C9",X"21",X"70",X"E5",X"7E",X"B7",X"20",X"0C",X"3A",X"78",X"E5",X"32",X"72",
		X"E5",X"3A",X"75",X"E5",X"32",X"71",X"E5",X"35",X"C9",X"1F",X"CB",X"11",X"3A",X"FD",X"E4",X"32",
		X"69",X"E5",X"DD",X"21",X"7B",X"E5",X"21",X"69",X"E5",X"7E",X"B7",X"C8",X"35",X"DD",X"7E",X"00",
		X"DD",X"66",X"01",X"87",X"87",X"87",X"CB",X"3C",X"1F",X"6F",X"11",X"10",X"D0",X"19",X"DD",X"7E",
		X"02",X"DD",X"96",X"01",X"3C",X"47",X"CB",X"41",X"28",X"08",X"36",X"17",X"2C",X"2C",X"36",X"17",
		X"18",X"06",X"36",X"10",X"2C",X"2C",X"36",X"14",X"2D",X"2D",X"11",X"80",X"00",X"19",X"10",X"E6",
		X"11",X"03",X"00",X"DD",X"19",X"18",X"BF",X"3A",X"CD",X"E5",X"4F",X"87",X"81",X"6F",X"26",X"00",
		X"29",X"29",X"29",X"29",X"22",X"F6",X"E4",X"21",X"30",X"64",X"06",X"00",X"09",X"7E",X"32",X"F8",
		X"E4",X"21",X"39",X"64",X"09",X"7E",X"32",X"F5",X"E4",X"21",X"42",X"64",X"09",X"7E",X"32",X"FB",
		X"E4",X"79",X"E6",X"07",X"3C",X"4F",X"21",X"30",X"64",X"09",X"7E",X"32",X"6E",X"E5",X"21",X"42",
		X"64",X"09",X"7E",X"32",X"6F",X"E5",X"3A",X"8E",X"E5",X"CD",X"EC",X"31",X"4F",X"06",X"00",X"21",
		X"4B",X"64",X"09",X"7E",X"32",X"D8",X"E5",X"21",X"4E",X"64",X"09",X"7E",X"32",X"D9",X"E5",X"C9",
		X"00",X"04",X"08",X"0E",X"0A",X"07",X"0F",X"05",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",
		X"01",X"00",X"00",X"01",X"01",X"01",X"00",X"01",X"01",X"00",X"01",X"09",X"0A",X"08",X"0D",X"0E",
		X"0C",X"AF",X"32",X"89",X"E5",X"7E",X"B7",X"C8",X"3D",X"20",X"24",X"23",X"EB",X"1A",X"6F",X"13",
		X"1A",X"13",X"D5",X"CB",X"3F",X"CB",X"10",X"5D",X"57",X"D5",X"CD",X"00",X"2D",X"D1",X"CB",X"40",
		X"28",X"02",X"2C",X"2C",X"EB",X"7C",X"CD",X"D5",X"62",X"E5",X"DD",X"E1",X"E1",X"18",X"D6",X"3D",
		X"20",X"08",X"23",X"7E",X"32",X"88",X"E5",X"23",X"18",X"CB",X"06",X"01",X"3D",X"20",X"14",X"23",
		X"46",X"23",X"CB",X"78",X"28",X"0D",X"78",X"06",X"30",X"E6",X"7F",X"FE",X"02",X"38",X"04",X"3D",
		X"32",X"89",X"E5",X"3A",X"88",X"E5",X"E6",X"0F",X"CB",X"4B",X"28",X"0E",X"4F",X"DD",X"7E",X"00",
		X"E6",X"F0",X"B1",X"DD",X"77",X"00",X"DD",X"23",X"18",X"0E",X"0F",X"0F",X"0F",X"0F",X"4F",X"DD",
		X"7E",X"00",X"E6",X"0F",X"B1",X"DD",X"77",X"00",X"7E",X"12",X"13",X"3A",X"88",X"E5",X"E6",X"F0",
		X"12",X"13",X"7B",X"FE",X"70",X"20",X"02",X"1E",X"90",X"FE",X"F0",X"20",X"03",X"1E",X"10",X"14",
		X"10",X"C1",X"3A",X"89",X"E5",X"B7",X"28",X"08",X"3D",X"32",X"89",X"E5",X"06",X"30",X"18",X"B3",
		X"23",X"C3",X"55",X"64",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"21",X"36",X"D5",X"11",X"1F",X"68",X"CD",X"2D",X"30",X"3E",X"24",X"CD",X"3E",X"30",X"DB",X"04",
		X"CB",X"57",X"28",X"2D",X"DB",X"03",X"0F",X"0F",X"E6",X"3C",X"C6",X"10",X"21",X"FA",X"65",X"5F",
		X"16",X"00",X"19",X"5E",X"23",X"56",X"23",X"D5",X"7E",X"23",X"66",X"6F",X"11",X"B0",X"D6",X"EB",
		X"CD",X"2D",X"30",X"3E",X"24",X"CD",X"3E",X"30",X"D1",X"21",X"B0",X"D7",X"CD",X"2D",X"30",X"18",
		X"39",X"DB",X"03",X"07",X"07",X"07",X"F5",X"E6",X"06",X"5F",X"16",X"00",X"21",X"FA",X"65",X"19",
		X"5E",X"23",X"56",X"23",X"F1",X"D5",X"07",X"07",X"E6",X"06",X"C6",X"08",X"5F",X"16",X"00",X"21",
		X"FA",X"65",X"19",X"7E",X"23",X"66",X"6F",X"11",X"AC",X"D6",X"EB",X"CD",X"2D",X"30",X"3E",X"24",
		X"CD",X"3E",X"30",X"D1",X"21",X"AC",X"D7",X"CD",X"2D",X"30",X"06",X"06",X"C5",X"21",X"36",X"D5",
		X"11",X"2D",X"68",X"CD",X"2D",X"30",X"3E",X"0C",X"CD",X"3E",X"30",X"21",X"36",X"D5",X"11",X"1F",
		X"68",X"CD",X"2D",X"30",X"3E",X"18",X"CD",X"3E",X"30",X"C1",X"10",X"E0",X"C9",X"3A",X"57",X"E4",
		X"FE",X"01",X"20",X"0B",X"21",X"28",X"DA",X"11",X"3B",X"68",X"CD",X"2D",X"30",X"18",X"4A",X"3A",
		X"57",X"E4",X"FE",X"02",X"20",X"16",X"0E",X"C6",X"21",X"3C",X"DB",X"11",X"55",X"68",X"CD",X"2D",
		X"30",X"21",X"BC",X"DB",X"11",X"5A",X"68",X"CD",X"2D",X"30",X"18",X"2D",X"3A",X"57",X"E4",X"FE",
		X"03",X"20",X"0B",X"21",X"B2",X"DC",X"11",X"5F",X"68",X"CD",X"2D",X"30",X"18",X"1B",X"3A",X"57",
		X"E4",X"FE",X"04",X"20",X"14",X"0E",X"C6",X"21",X"B6",X"DD",X"11",X"6F",X"68",X"CD",X"2D",X"30",
		X"21",X"36",X"DE",X"11",X"7A",X"68",X"CD",X"2D",X"30",X"C9",X"C6",X"67",X"DC",X"67",X"F2",X"67",
		X"08",X"68",X"1E",X"68",X"87",X"67",X"9C",X"67",X"B1",X"67",X"1E",X"68",X"1E",X"68",X"1E",X"68",
		X"1E",X"68",X"1E",X"68",X"1E",X"68",X"1E",X"68",X"28",X"67",X"1E",X"68",X"3B",X"67",X"1E",X"68",
		X"4E",X"67",X"1E",X"68",X"61",X"67",X"1E",X"68",X"74",X"67",X"1E",X"68",X"1E",X"68",X"1E",X"68",
		X"1E",X"68",X"5C",X"66",X"4A",X"66",X"81",X"66",X"6F",X"66",X"A6",X"66",X"94",X"66",X"CB",X"66",
		X"B9",X"66",X"F0",X"66",X"DE",X"66",X"15",X"67",X"03",X"67",X"20",X"36",X"20",X"43",X"4F",X"49",
		X"4E",X"53",X"20",X"31",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"00",X"31",X"32",X"20",X"43",
		X"4F",X"49",X"4E",X"53",X"20",X"32",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"53",X"00",X"20",
		X"35",X"20",X"43",X"4F",X"49",X"4E",X"53",X"20",X"31",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",
		X"00",X"31",X"30",X"20",X"43",X"4F",X"49",X"4E",X"53",X"20",X"32",X"20",X"50",X"4C",X"41",X"59",
		X"45",X"52",X"53",X"00",X"20",X"34",X"20",X"43",X"4F",X"49",X"4E",X"53",X"20",X"31",X"20",X"50",
		X"4C",X"41",X"59",X"45",X"52",X"00",X"20",X"38",X"20",X"43",X"4F",X"49",X"4E",X"53",X"20",X"32",
		X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"53",X"00",X"20",X"33",X"20",X"43",X"4F",X"49",X"4E",
		X"53",X"20",X"31",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"00",X"20",X"36",X"20",X"43",X"4F",
		X"49",X"4E",X"53",X"20",X"32",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"53",X"00",X"20",X"32",
		X"20",X"43",X"4F",X"49",X"4E",X"53",X"20",X"31",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"00",
		X"20",X"34",X"20",X"43",X"4F",X"49",X"4E",X"53",X"20",X"32",X"20",X"50",X"4C",X"41",X"59",X"45",
		X"52",X"53",X"00",X"20",X"31",X"20",X"43",X"4F",X"49",X"4E",X"20",X"20",X"31",X"20",X"50",X"4C",
		X"41",X"59",X"45",X"52",X"00",X"20",X"32",X"20",X"43",X"4F",X"49",X"4E",X"53",X"20",X"32",X"20",
		X"50",X"4C",X"41",X"59",X"45",X"52",X"53",X"00",X"20",X"31",X"20",X"43",X"4F",X"49",X"4E",X"20",
		X"20",X"36",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"53",X"00",X"20",X"31",X"20",X"43",X"4F",
		X"49",X"4E",X"20",X"20",X"35",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"53",X"00",X"20",X"31",
		X"20",X"43",X"4F",X"49",X"4E",X"20",X"20",X"34",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"53",
		X"00",X"20",X"31",X"20",X"43",X"4F",X"49",X"4E",X"20",X"20",X"33",X"20",X"50",X"4C",X"41",X"59",
		X"45",X"52",X"53",X"00",X"20",X"31",X"20",X"43",X"4F",X"49",X"4E",X"20",X"20",X"32",X"20",X"50",
		X"4C",X"41",X"59",X"45",X"52",X"53",X"00",X"41",X"20",X"2D",X"20",X"33",X"20",X"43",X"4F",X"49",
		X"4E",X"53",X"20",X"31",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"00",X"41",X"20",X"2D",X"20",
		X"32",X"20",X"43",X"4F",X"49",X"4E",X"53",X"20",X"31",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",
		X"00",X"41",X"20",X"2D",X"20",X"31",X"20",X"43",X"4F",X"49",X"4E",X"20",X"20",X"31",X"20",X"50",
		X"4C",X"41",X"59",X"45",X"52",X"00",X"42",X"20",X"2D",X"20",X"31",X"20",X"43",X"4F",X"49",X"4E",
		X"20",X"20",X"36",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"53",X"00",X"42",X"20",X"2D",X"20",
		X"31",X"20",X"43",X"4F",X"49",X"4E",X"20",X"20",X"35",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",
		X"53",X"00",X"42",X"20",X"2D",X"20",X"31",X"20",X"43",X"4F",X"49",X"4E",X"20",X"20",X"33",X"20",
		X"50",X"4C",X"41",X"59",X"45",X"52",X"53",X"00",X"42",X"20",X"2D",X"20",X"31",X"20",X"43",X"4F",
		X"49",X"4E",X"20",X"20",X"32",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"53",X"00",X"00",X"02",
		X"49",X"4E",X"53",X"45",X"52",X"54",X"20",X"20",X"43",X"4F",X"49",X"4E",X"00",X"02",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"00",X"06",X"40",X"31",X"39",X"38",
		X"34",X"20",X"20",X"20",X"49",X"52",X"45",X"4D",X"20",X"43",X"4F",X"52",X"50",X"4F",X"52",X"41",
		X"54",X"49",X"4F",X"4E",X"00",X"80",X"82",X"84",X"86",X"00",X"81",X"83",X"85",X"87",X"00",X"02",
		X"4C",X"49",X"43",X"45",X"4E",X"53",X"45",X"44",X"20",X"20",X"46",X"52",X"4F",X"4D",X"00",X"68",
		X"6A",X"6C",X"6E",X"70",X"72",X"74",X"76",X"78",X"7A",X"00",X"69",X"6B",X"6D",X"6F",X"71",X"73",
		X"75",X"77",X"79",X"7B",X"00",X"CD",X"5E",X"5F",X"3E",X"FF",X"32",X"D1",X"E5",X"CD",X"28",X"6D",
		X"3E",X"A8",X"CD",X"3E",X"30",X"3E",X"01",X"32",X"A9",X"E5",X"CD",X"5E",X"5F",X"C3",X"CF",X"25",
		X"31",X"00",X"E8",X"21",X"10",X"D0",X"36",X"00",X"54",X"5D",X"13",X"01",X"57",X"15",X"ED",X"B0",
		X"AF",X"32",X"A7",X"E5",X"32",X"9D",X"E5",X"32",X"6A",X"E5",X"FB",X"3E",X"50",X"32",X"B5",X"E5",
		X"21",X"B5",X"E5",X"7E",X"FE",X"14",X"38",X"0B",X"21",X"36",X"D5",X"11",X"91",X"69",X"CD",X"2D",
		X"30",X"18",X"12",X"B7",X"20",X"02",X"36",X"28",X"21",X"26",X"D5",X"36",X"00",X"54",X"5D",X"13",
		X"01",X"35",X"00",X"ED",X"B0",X"11",X"A0",X"69",X"3A",X"B2",X"E5",X"FE",X"02",X"38",X"03",X"11",
		X"B2",X"69",X"21",X"34",X"D7",X"CD",X"2D",X"30",X"CD",X"7F",X"69",X"21",X"AA",X"E5",X"7E",X"E6",
		X"0A",X"FE",X"0A",X"20",X"0E",X"3A",X"B2",X"E5",X"3D",X"27",X"32",X"B2",X"E5",X"AF",X"32",X"B7",
		X"E5",X"18",X"1B",X"7E",X"E6",X"05",X"FE",X"05",X"C2",X"C0",X"68",X"3A",X"B2",X"E5",X"FE",X"02",
		X"DA",X"C0",X"68",X"D6",X"02",X"27",X"32",X"B2",X"E5",X"3E",X"01",X"32",X"B7",X"E5",X"AF",X"32",
		X"B9",X"E5",X"32",X"B8",X"E5",X"32",X"90",X"E5",X"32",X"96",X"E5",X"3C",X"32",X"B2",X"E6",X"CB",
		X"41",X"20",X"06",X"32",X"8E",X"E5",X"32",X"94",X"E5",X"3A",X"E0",X"E5",X"32",X"8F",X"E5",X"32",
		X"95",X"E5",X"21",X"00",X"00",X"22",X"91",X"E5",X"22",X"92",X"E5",X"22",X"97",X"E5",X"22",X"98",
		X"E5",X"21",X"80",X"00",X"DB",X"04",X"CB",X"47",X"20",X"02",X"2D",X"2D",X"22",X"E3",X"E5",X"21",
		X"10",X"D3",X"36",X"00",X"54",X"5D",X"13",X"01",X"7F",X"09",X"ED",X"B0",X"C3",X"0F",X"5D",X"21",
		X"42",X"DC",X"11",X"C6",X"69",X"CD",X"2D",X"30",X"0E",X"02",X"11",X"B2",X"E5",X"CD",X"5F",X"30",
		X"C9",X"04",X"50",X"55",X"53",X"48",X"20",X"20",X"20",X"42",X"55",X"54",X"54",X"4F",X"4E",X"00",
		X"04",X"4F",X"4E",X"4C",X"59",X"20",X"20",X"02",X"31",X"20",X"04",X"50",X"4C",X"41",X"59",X"45",
		X"52",X"00",X"02",X"31",X"20",X"04",X"4F",X"52",X"20",X"02",X"32",X"20",X"20",X"04",X"50",X"4C",
		X"41",X"59",X"45",X"52",X"53",X"00",X"04",X"43",X"52",X"45",X"44",X"49",X"54",X"20",X"00",X"06",
		X"31",X"53",X"54",X"20",X"20",X"42",X"4C",X"4F",X"43",X"4B",X"00",X"21",X"30",X"D3",X"11",X"8F",
		X"6A",X"CD",X"2D",X"30",X"3E",X"22",X"CD",X"42",X"31",X"3E",X"0A",X"32",X"88",X"E5",X"3E",X"38",
		X"32",X"B6",X"E5",X"3E",X"50",X"32",X"B5",X"E5",X"21",X"B6",X"E5",X"7E",X"B7",X"20",X"09",X"36",
		X"38",X"21",X"88",X"E5",X"35",X"CA",X"89",X"6A",X"21",X"B5",X"E5",X"7E",X"FE",X"14",X"38",X"1C",
		X"3A",X"B2",X"E5",X"B7",X"20",X"0B",X"21",X"24",X"D5",X"11",X"A1",X"6A",X"CD",X"2D",X"30",X"18",
		X"09",X"21",X"24",X"D5",X"11",X"C6",X"6A",X"CD",X"2D",X"30",X"18",X"12",X"B7",X"20",X"02",X"36",
		X"27",X"21",X"24",X"D5",X"36",X"00",X"54",X"5D",X"13",X"01",X"35",X"00",X"ED",X"B0",X"CD",X"7F",
		X"69",X"21",X"3A",X"D9",X"11",X"BE",X"6A",X"CD",X"2D",X"30",X"0E",X"06",X"3A",X"88",X"E5",X"3D",
		X"CD",X"6A",X"30",X"21",X"AA",X"E5",X"7E",X"E6",X"0A",X"FE",X"0A",X"28",X"07",X"7E",X"E6",X"05",
		X"FE",X"05",X"20",X"22",X"3A",X"B2",X"E5",X"B7",X"CA",X"F8",X"69",X"D6",X"01",X"27",X"32",X"B2",
		X"E5",X"AF",X"32",X"90",X"E5",X"3A",X"E0",X"E5",X"32",X"8F",X"E5",X"21",X"00",X"00",X"22",X"91",
		X"E5",X"22",X"92",X"E5",X"18",X"03",X"C3",X"F8",X"69",X"3E",X"00",X"CD",X"42",X"31",X"C9",X"03",
		X"54",X"4F",X"20",X"43",X"4F",X"4E",X"54",X"49",X"4E",X"55",X"45",X"20",X"47",X"41",X"4D",X"45",
		X"00",X"04",X"49",X"4E",X"53",X"45",X"52",X"54",X"20",X"43",X"4F",X"49",X"4E",X"20",X"41",X"4E",
		X"44",X"20",X"50",X"55",X"53",X"48",X"20",X"42",X"55",X"54",X"54",X"4F",X"4E",X"00",X"03",X"54",
		X"49",X"4D",X"45",X"20",X"20",X"00",X"04",X"20",X"20",X"20",X"20",X"20",X"50",X"55",X"53",X"48",
		X"20",X"53",X"54",X"41",X"52",X"54",X"20",X"42",X"55",X"54",X"54",X"4F",X"4E",X"20",X"20",X"20",
		X"20",X"20",X"00",X"3E",X"13",X"CD",X"42",X"31",X"CD",X"5E",X"5F",X"3A",X"90",X"E5",X"FE",X"02",
		X"20",X"26",X"AF",X"32",X"B2",X"E6",X"CD",X"A8",X"6B",X"CD",X"DB",X"69",X"3E",X"01",X"32",X"B2",
		X"E6",X"3A",X"90",X"E5",X"FE",X"00",X"20",X"10",X"21",X"10",X"D3",X"36",X"00",X"54",X"5D",X"13",
		X"01",X"7F",X"09",X"ED",X"B0",X"C3",X"0F",X"5D",X"3A",X"B7",X"E5",X"FE",X"00",X"28",X"07",X"3A",
		X"96",X"E5",X"FE",X"02",X"20",X"2E",X"3A",X"90",X"E5",X"FE",X"02",X"28",X"10",X"21",X"10",X"D3",
		X"36",X"00",X"54",X"5D",X"13",X"01",X"7F",X"09",X"ED",X"B0",X"C3",X"0F",X"5D",X"CD",X"5E",X"5F",
		X"AF",X"32",X"B2",X"E6",X"32",X"B9",X"E5",X"3E",X"01",X"CD",X"3E",X"30",X"3E",X"01",X"32",X"A7",
		X"E5",X"C3",X"CF",X"25",X"21",X"10",X"D3",X"36",X"00",X"54",X"5D",X"13",X"01",X"7F",X"09",X"ED",
		X"B0",X"21",X"B8",X"E5",X"7E",X"B7",X"20",X"03",X"34",X"18",X"02",X"36",X"00",X"CD",X"96",X"6B",
		X"DB",X"04",X"CB",X"4F",X"28",X"1D",X"21",X"B9",X"E5",X"CB",X"46",X"20",X"03",X"34",X"18",X"01",
		X"35",X"E6",X"01",X"AE",X"21",X"80",X"00",X"20",X"02",X"2D",X"2D",X"22",X"E3",X"E5",X"3E",X"01",
		X"CD",X"3E",X"30",X"C3",X"0F",X"5D",X"21",X"8E",X"E5",X"11",X"94",X"E5",X"06",X"06",X"1A",X"4E",
		X"77",X"79",X"12",X"23",X"13",X"10",X"F7",X"C9",X"0E",X"00",X"16",X"15",X"21",X"E5",X"E5",X"06",
		X"00",X"09",X"DD",X"21",X"91",X"E5",X"06",X"03",X"DD",X"7E",X"00",X"BE",X"38",X"12",X"28",X"0B",
		X"15",X"3E",X"0A",X"81",X"4F",X"FE",X"C8",X"28",X"07",X"18",X"E1",X"DD",X"23",X"23",X"10",X"E8",
		X"7A",X"32",X"D1",X"E5",X"79",X"B7",X"C8",X"D6",X"0A",X"11",X"E5",X"E5",X"28",X"08",X"4F",X"06",
		X"00",X"21",X"EF",X"E5",X"ED",X"B0",X"21",X"91",X"E5",X"01",X"03",X"00",X"ED",X"B0",X"62",X"6B",
		X"36",X"00",X"13",X"01",X"05",X"00",X"ED",X"B0",X"3A",X"8E",X"E5",X"12",X"CD",X"28",X"6D",X"21",
		X"B8",X"D2",X"11",X"22",X"6D",X"CD",X"2D",X"30",X"DD",X"2A",X"D2",X"E5",X"11",X"16",X"00",X"DD",
		X"19",X"FD",X"2A",X"D4",X"E5",X"FD",X"23",X"FD",X"23",X"FD",X"23",X"0E",X"41",X"1E",X"03",X"3E",
		X"14",X"32",X"88",X"E5",X"21",X"C2",X"D2",X"C5",X"0E",X"06",X"3A",X"88",X"E5",X"CD",X"48",X"30",
		X"C1",X"06",X"04",X"3E",X"0E",X"32",X"B6",X"E5",X"AF",X"32",X"89",X"E5",X"3A",X"D0",X"E5",X"B7",
		X"20",X"03",X"57",X"18",X"44",X"7A",X"B7",X"20",X"13",X"3A",X"D0",X"E5",X"FE",X"0A",X"20",X"04",
		X"14",X"0C",X"18",X"06",X"FE",X"05",X"20",X"02",X"15",X"0D",X"18",X"1F",X"3A",X"D0",X"E5",X"FE",
		X"AA",X"20",X"0B",X"14",X"7A",X"FE",X"18",X"20",X"03",X"0C",X"16",X"0C",X"18",X"0D",X"FE",X"55",
		X"20",X"09",X"15",X"7A",X"FE",X"E8",X"20",X"03",X"0D",X"16",X"F4",X"79",X"FE",X"5D",X"38",X"02",
		X"0E",X"41",X"79",X"FE",X"41",X"30",X"02",X"0E",X"5C",X"3A",X"CF",X"E5",X"FE",X"05",X"28",X"04",
		X"FE",X"0A",X"20",X"21",X"21",X"89",X"E5",X"3A",X"B6",X"E5",X"BE",X"38",X"18",X"3C",X"77",X"79",
		X"FE",X"5C",X"28",X"3D",X"FD",X"71",X"00",X"FD",X"23",X"DD",X"71",X"00",X"0E",X"41",X"DD",X"23",
		X"DD",X"23",X"1D",X"28",X"2C",X"CB",X"40",X"28",X"05",X"DD",X"71",X"00",X"18",X"03",X"DD",X"71",
		X"00",X"3A",X"AA",X"E5",X"B7",X"20",X"1A",X"3E",X"01",X"CD",X"3E",X"30",X"3A",X"B6",X"E5",X"B7",
		X"C2",X"3C",X"6C",X"05",X"C2",X"33",X"6C",X"21",X"88",X"E5",X"35",X"7E",X"FE",X"FF",X"C2",X"24",
		X"6C",X"DD",X"36",X"00",X"00",X"3E",X"38",X"CD",X"3E",X"30",X"3E",X"13",X"CD",X"42",X"31",X"CD",
		X"5E",X"5F",X"C9",X"03",X"42",X"45",X"53",X"54",X"20",X"20",X"06",X"32",X"30",X"20",X"20",X"03",
		X"50",X"4C",X"41",X"59",X"45",X"52",X"53",X"00",X"02",X"20",X"4E",X"4F",X"2E",X"53",X"43",X"4F",
		X"52",X"45",X"53",X"20",X"20",X"4E",X"41",X"4D",X"45",X"20",X"52",X"4F",X"55",X"4E",X"44",X"20",
		X"20",X"00",X"02",X"54",X"49",X"4D",X"45",X"00",X"21",X"B0",X"D1",X"11",X"F3",X"6C",X"CD",X"2D",
		X"30",X"21",X"90",X"D3",X"11",X"08",X"6D",X"CD",X"2D",X"30",X"11",X"08",X"6D",X"CD",X"2D",X"30",
		X"11",X"E5",X"E5",X"21",X"C2",X"DD",X"3A",X"D1",X"E5",X"4F",X"06",X"14",X"78",X"FE",X"0A",X"20",
		X"03",X"21",X"92",X"DD",X"B9",X"20",X"07",X"22",X"D2",X"E5",X"ED",X"53",X"D4",X"E5",X"C5",X"E5",
		X"41",X"0E",X"02",X"B8",X"20",X"02",X"0E",X"06",X"FE",X"0A",X"30",X"07",X"2C",X"2C",X"CD",X"6A",
		X"30",X"18",X"03",X"CD",X"48",X"30",X"2C",X"2C",X"79",X"FE",X"02",X"20",X"02",X"0E",X"04",X"06",
		X"03",X"CD",X"5F",X"30",X"10",X"FB",X"2C",X"2C",X"2C",X"2C",X"06",X"03",X"1A",X"77",X"2C",X"71",
		X"2C",X"13",X"10",X"F8",X"7D",X"C6",X"06",X"6F",X"13",X"13",X"13",X"1A",X"CD",X"48",X"30",X"13",
		X"E1",X"C1",X"25",X"10",X"A7",X"C9",X"01",X"03",X"00",X"11",X"9A",X"E5",X"21",X"7B",X"6E",X"ED",
		X"B0",X"01",X"C8",X"00",X"11",X"E5",X"E5",X"21",X"BD",X"6D",X"ED",X"B0",X"C9",X"01",X"01",X"00",
		X"53",X"54",X"45",X"20",X"20",X"20",X"01",X"01",X"03",X"50",X"4F",X"49",X"4E",X"20",X"20",X"20",
		X"01",X"01",X"08",X"80",X"45",X"48",X"45",X"20",X"20",X"20",X"02",X"01",X"10",X"30",X"4D",X"49",
		X"54",X"20",X"20",X"20",X"01",X"01",X"21",X"50",X"41",X"41",X"54",X"20",X"20",X"20",X"01",X"01",
		X"23",X"50",X"47",X"4E",X"41",X"20",X"20",X"20",X"02",X"01",X"28",X"00",X"4F",X"41",X"59",X"20",
		X"20",X"20",X"02",X"01",X"38",X"70",X"4E",X"52",X"41",X"20",X"20",X"20",X"02",X"01",X"60",X"10",
		X"4F",X"49",X"57",X"20",X"20",X"20",X"02",X"01",X"89",X"90",X"4B",X"48",X"4F",X"20",X"20",X"20",
		X"02",X"02",X"66",X"00",X"48",X"4E",X"49",X"20",X"20",X"20",X"02",X"02",X"77",X"50",X"53",X"41",
		X"4F",X"20",X"20",X"20",X"02",X"03",X"12",X"50",X"55",X"48",X"59",X"20",X"20",X"20",X"02",X"03",
		X"33",X"00",X"42",X"53",X"41",X"20",X"20",X"20",X"03",X"03",X"65",X"00",X"41",X"49",X"57",X"20",
		X"20",X"20",X"03",X"03",X"70",X"50",X"4B",X"41",X"45",X"20",X"20",X"20",X"04",X"03",X"88",X"00",
		X"4D",X"4B",X"4D",X"20",X"20",X"20",X"03",X"04",X"01",X"50",X"45",X"49",X"41",X"20",X"20",X"20",
		X"03",X"04",X"32",X"00",X"52",X"4B",X"47",X"20",X"20",X"20",X"03",X"04",X"85",X"40",X"49",X"49",
		X"4F",X"20",X"20",X"20",X"04",X"F9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"31",X"00",X"E8",X"11",X"00",X"20",X"CD",X"2D",X"6F",X"22",X"74",X"00",X"CD",X"2D",X"6F",X"22",
		X"76",X"00",X"CD",X"2D",X"6F",X"22",X"78",X"00",X"11",X"00",X"00",X"CD",X"2D",X"6F",X"22",X"72",
		X"00",X"11",X"FF",X"FF",X"EB",X"A7",X"ED",X"52",X"22",X"70",X"00",X"18",X"FE",X"01",X"00",X"20",
		X"21",X"00",X"00",X"1A",X"85",X"6F",X"3E",X"00",X"8C",X"67",X"13",X"0B",X"78",X"B1",X"20",X"F3",
		X"C9",X"F3",X"ED",X"46",X"31",X"00",X"E8",X"DD",X"21",X"4E",X"6F",X"C3",X"90",X"72",X"0E",X"05",
		X"3E",X"FF",X"ED",X"79",X"0C",X"ED",X"79",X"0C",X"ED",X"79",X"21",X"00",X"E1",X"36",X"00",X"54",
		X"5D",X"13",X"01",X"FF",X"01",X"ED",X"B0",X"FB",X"01",X"00",X"80",X"0B",X"79",X"B0",X"20",X"FB",
		X"F3",X"AF",X"5F",X"16",X"20",X"21",X"00",X"E0",X"0E",X"10",X"06",X"00",X"77",X"23",X"3C",X"15",
		X"28",X"07",X"10",X"F8",X"0D",X"20",X"F3",X"18",X"05",X"16",X"20",X"3C",X"18",X"F4",X"7B",X"16",
		X"20",X"21",X"00",X"E0",X"0E",X"10",X"06",X"00",X"BE",X"C2",X"95",X"71",X"23",X"3C",X"15",X"28",
		X"07",X"10",X"F5",X"0D",X"20",X"F0",X"18",X"05",X"3C",X"16",X"20",X"18",X"F4",X"7B",X"3C",X"FE",
		X"0F",X"20",X"BF",X"31",X"00",X"E8",X"CD",X"F2",X"77",X"AF",X"32",X"01",X"E0",X"16",X"20",X"0E",
		X"10",X"21",X"00",X"D0",X"06",X"00",X"77",X"23",X"3C",X"15",X"28",X"07",X"10",X"F8",X"0D",X"20",
		X"F3",X"18",X"05",X"3C",X"16",X"20",X"18",X"F4",X"3A",X"01",X"E0",X"16",X"20",X"21",X"00",X"D0",
		X"0E",X"10",X"06",X"00",X"CD",X"35",X"72",X"23",X"3C",X"15",X"28",X"07",X"10",X"F6",X"0D",X"20",
		X"F1",X"18",X"05",X"3C",X"16",X"20",X"18",X"F4",X"3A",X"01",X"E0",X"3C",X"FE",X"0F",X"20",X"BA",
		X"DD",X"21",X"BF",X"70",X"CD",X"90",X"72",X"21",X"0F",X"7A",X"DD",X"21",X"BF",X"70",X"CD",X"28",
		X"71",X"CD",X"AF",X"70",X"CD",X"F2",X"77",X"3E",X"03",X"32",X"01",X"E7",X"CD",X"9E",X"79",X"3E",
		X"01",X"32",X"00",X"E3",X"32",X"02",X"E3",X"DB",X"00",X"2F",X"0F",X"0F",X"30",X"F9",X"3E",X"03",
		X"32",X"01",X"E7",X"CD",X"B6",X"77",X"21",X"AA",X"7B",X"CD",X"D5",X"77",X"3A",X"01",X"E7",X"06",
		X"06",X"CD",X"4A",X"7D",X"CD",X"95",X"79",X"CD",X"95",X"79",X"DB",X"00",X"2F",X"0F",X"30",X"14",
		X"3A",X"01",X"E7",X"07",X"4F",X"06",X"00",X"DD",X"21",X"98",X"7B",X"DD",X"09",X"DD",X"66",X"01",
		X"DD",X"6E",X"00",X"E9",X"CD",X"9E",X"79",X"CD",X"9E",X"79",X"CD",X"95",X"79",X"CD",X"95",X"79",
		X"DB",X"01",X"2F",X"0F",X"38",X"05",X"0F",X"38",X"1C",X"18",X"C9",X"3A",X"01",X"E7",X"FE",X"08",
		X"CA",X"44",X"70",X"06",X"04",X"CD",X"4A",X"7D",X"C6",X"01",X"32",X"01",X"E7",X"06",X"06",X"CD",
		X"4A",X"7D",X"C3",X"44",X"70",X"3A",X"01",X"E7",X"FE",X"03",X"CA",X"44",X"70",X"06",X"04",X"CD",
		X"4A",X"7D",X"C6",X"FF",X"32",X"01",X"E7",X"06",X"06",X"CD",X"4A",X"7D",X"C3",X"44",X"70",X"11",
		X"00",X"00",X"AF",X"32",X"00",X"E7",X"06",X"04",X"C5",X"CD",X"C0",X"70",X"C1",X"10",X"F9",X"C9",
		X"21",X"00",X"00",X"06",X"20",X"1A",X"85",X"30",X"01",X"24",X"6F",X"1C",X"20",X"F7",X"14",X"10",
		X"F4",X"D5",X"E5",X"3A",X"00",X"E7",X"21",X"72",X"00",X"87",X"85",X"6F",X"5E",X"23",X"56",X"E1",
		X"7A",X"BC",X"20",X"09",X"7B",X"BD",X"20",X"05",X"21",X"2F",X"7A",X"18",X"03",X"21",X"38",X"7A",
		X"11",X"83",X"E7",X"01",X"09",X"00",X"ED",X"B0",X"11",X"00",X"01",X"21",X"A0",X"D1",X"3A",X"00",
		X"E7",X"A7",X"28",X"04",X"47",X"19",X"10",X"FD",X"22",X"81",X"E7",X"3E",X"08",X"32",X"80",X"E7",
		X"3A",X"00",X"E7",X"C6",X"30",X"32",X"86",X"E7",X"21",X"00",X"E7",X"34",X"21",X"80",X"E7",X"DD",
		X"21",X"BF",X"70",X"CD",X"28",X"71",X"D1",X"C9",X"7E",X"23",X"FE",X"00",X"28",X"12",X"5E",X"23",
		X"56",X"23",X"4F",X"7E",X"12",X"13",X"3E",X"04",X"12",X"23",X"13",X"0D",X"20",X"F5",X"18",X"E8",
		X"DD",X"E9",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"C6",X"30",X"FE",X"3A",X"38",X"02",X"C6",X"07",
		X"FD",X"77",X"00",X"FD",X"36",X"01",X"04",X"DD",X"E9",X"E6",X"0F",X"C6",X"30",X"FE",X"3A",X"38",
		X"02",X"C6",X"07",X"FD",X"77",X"00",X"FD",X"36",X"01",X"04",X"DD",X"E9",X"F5",X"0F",X"0F",X"0F",
		X"0F",X"E6",X"0F",X"C6",X"30",X"FE",X"3A",X"38",X"02",X"C6",X"07",X"FD",X"77",X"00",X"FD",X"36",
		X"01",X"04",X"F1",X"E6",X"0F",X"C6",X"30",X"FE",X"3A",X"38",X"02",X"C6",X"07",X"FD",X"77",X"02",
		X"FD",X"36",X"03",X"04",X"C9",X"08",X"D9",X"DD",X"21",X"9E",X"71",X"C3",X"15",X"72",X"21",X"1B",
		X"7A",X"DD",X"21",X"A8",X"71",X"C3",X"28",X"71",X"D9",X"FD",X"21",X"B8",X"D0",X"DD",X"21",X"B5",
		X"71",X"7C",X"C3",X"42",X"71",X"FD",X"23",X"FD",X"23",X"DD",X"21",X"C1",X"71",X"7C",X"C3",X"59",
		X"71",X"DD",X"21",X"CD",X"71",X"7D",X"FD",X"23",X"FD",X"23",X"C3",X"42",X"71",X"DD",X"21",X"D9",
		X"71",X"7D",X"FD",X"23",X"FD",X"23",X"C3",X"59",X"71",X"08",X"D9",X"FD",X"23",X"FD",X"23",X"FD",
		X"23",X"FD",X"23",X"DD",X"21",X"EB",X"71",X"5F",X"C3",X"42",X"71",X"FD",X"23",X"FD",X"23",X"DD",
		X"21",X"F7",X"71",X"7B",X"C3",X"59",X"71",X"08",X"D9",X"FD",X"23",X"FD",X"23",X"FD",X"23",X"FD",
		X"23",X"DD",X"21",X"09",X"72",X"7E",X"C3",X"42",X"71",X"FD",X"23",X"FD",X"23",X"7E",X"DD",X"21",
		X"23",X"72",X"C3",X"59",X"71",X"21",X"01",X"D0",X"01",X"FF",X"0F",X"36",X"00",X"54",X"5D",X"ED",
		X"B0",X"DD",X"E9",X"CD",X"9E",X"79",X"DB",X"00",X"0F",X"38",X"06",X"0F",X"DA",X"B3",X"6F",X"18",
		X"F2",X"08",X"C3",X"9C",X"6F",X"BE",X"C8",X"F5",X"E5",X"DD",X"21",X"40",X"72",X"C3",X"90",X"72",
		X"21",X"1B",X"7A",X"DD",X"21",X"4A",X"72",X"C3",X"28",X"71",X"E1",X"FD",X"21",X"B8",X"D0",X"7C",
		X"CD",X"6C",X"71",X"FD",X"23",X"FD",X"23",X"FD",X"23",X"FD",X"23",X"7D",X"CD",X"6C",X"71",X"F1",
		X"F5",X"FD",X"23",X"FD",X"23",X"FD",X"23",X"FD",X"23",X"CD",X"6C",X"71",X"FD",X"23",X"FD",X"23",
		X"FD",X"23",X"FD",X"23",X"7E",X"CD",X"6C",X"71",X"CD",X"9E",X"79",X"CD",X"9E",X"79",X"DB",X"00",
		X"0F",X"DA",X"89",X"72",X"0F",X"38",X"04",X"18",X"EF",X"F1",X"C9",X"F1",X"C1",X"C3",X"00",X"70",
		X"21",X"01",X"D0",X"01",X"FF",X"07",X"36",X"00",X"54",X"5D",X"13",X"13",X"CD",X"A7",X"79",X"21",
		X"00",X"D0",X"01",X"FF",X"07",X"36",X"00",X"54",X"5D",X"13",X"13",X"CD",X"A7",X"79",X"DD",X"E9",
		X"3E",X"FF",X"D3",X"05",X"CD",X"B6",X"77",X"21",X"41",X"7A",X"CD",X"D5",X"77",X"DB",X"03",X"21",
		X"AE",X"D1",X"CD",X"33",X"76",X"DB",X"04",X"21",X"AE",X"D2",X"CD",X"33",X"76",X"CD",X"E4",X"72",
		X"CD",X"72",X"73",X"CD",X"95",X"79",X"CD",X"95",X"79",X"DB",X"00",X"EE",X"FF",X"0F",X"0F",X"DA",
		X"33",X"70",X"18",X"D9",X"21",X"87",X"74",X"CD",X"D5",X"77",X"CD",X"B0",X"73",X"DB",X"04",X"EE",
		X"FF",X"CB",X"57",X"28",X"4B",X"21",X"FC",X"73",X"CD",X"D5",X"77",X"DB",X"03",X"EE",X"FF",X"0F",
		X"0F",X"0F",X"0F",X"11",X"00",X"00",X"21",X"90",X"73",X"01",X"00",X"05",X"E6",X"0F",X"20",X"0A",
		X"19",X"5E",X"23",X"66",X"6B",X"CD",X"D5",X"77",X"18",X"25",X"0C",X"1C",X"1C",X"B9",X"20",X"02",
		X"18",X"EE",X"10",X"F6",X"01",X"08",X"05",X"1C",X"1C",X"B9",X"20",X"02",X"18",X"09",X"0C",X"10",
		X"F6",X"FE",X"0F",X"20",X"0A",X"1C",X"1C",X"19",X"5E",X"23",X"66",X"6B",X"CD",X"D5",X"77",X"C9",
		X"21",X"2A",X"74",X"CD",X"D5",X"77",X"DB",X"03",X"EE",X"FF",X"21",X"A8",X"73",X"11",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"28",X"11",X"1C",X"1C",X"FE",X"08",X"28",X"0B",X"1C",X"1C",
		X"FE",X"0A",X"28",X"05",X"1C",X"1C",X"FE",X"0F",X"C0",X"19",X"5E",X"23",X"66",X"6B",X"CD",X"D5",
		X"77",X"C9",X"DB",X"04",X"2F",X"0F",X"0F",X"38",X"13",X"AF",X"87",X"21",X"AE",X"74",X"85",X"6F",
		X"3E",X"00",X"8C",X"67",X"5E",X"23",X"66",X"6B",X"CD",X"D5",X"77",X"C9",X"3E",X"01",X"18",X"EA",
		X"D2",X"74",X"E3",X"74",X"F5",X"74",X"07",X"75",X"19",X"75",X"2B",X"75",X"3D",X"75",X"4F",X"75",
		X"61",X"75",X"73",X"75",X"85",X"75",X"97",X"75",X"A8",X"75",X"CB",X"75",X"EE",X"75",X"11",X"76",
		X"DB",X"03",X"EE",X"FF",X"47",X"E6",X"03",X"28",X"25",X"FE",X"01",X"28",X"26",X"FE",X"02",X"28",
		X"27",X"21",X"47",X"74",X"CD",X"D5",X"77",X"78",X"0F",X"0F",X"47",X"E6",X"03",X"28",X"1E",X"FE",
		X"01",X"28",X"1F",X"FE",X"02",X"28",X"20",X"21",X"52",X"74",X"CD",X"D5",X"77",X"C9",X"21",X"57",
		X"74",X"18",X"E1",X"21",X"67",X"74",X"18",X"DC",X"21",X"77",X"74",X"18",X"D7",X"21",X"62",X"74",
		X"18",X"E8",X"21",X"72",X"74",X"18",X"E3",X"21",X"82",X"74",X"18",X"DE",X"0B",X"92",X"D3",X"43",
		X"4F",X"49",X"4E",X"20",X"4D",X"4F",X"44",X"45",X"20",X"20",X"0B",X"12",X"D4",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"0E",X"30",X"D4",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"00",X"0B",X"92",X"D3",X"43",X"4F",X"49",
		X"4E",X"20",X"4D",X"4F",X"44",X"45",X"20",X"41",X"0B",X"12",X"D4",X"43",X"4F",X"49",X"4E",X"20",
		X"4D",X"4F",X"44",X"45",X"20",X"42",X"00",X"07",X"30",X"D6",X"31",X"35",X"35",X"20",X"53",X"45",
		X"43",X"00",X"01",X"B0",X"D6",X"35",X"00",X"07",X"30",X"D6",X"31",X"38",X"30",X"20",X"53",X"45",
		X"43",X"00",X"01",X"B0",X"D6",X"33",X"00",X"07",X"30",X"D6",X"31",X"37",X"30",X"20",X"53",X"45",
		X"43",X"00",X"01",X"B0",X"D6",X"32",X"00",X"07",X"30",X"D6",X"31",X"36",X"30",X"20",X"53",X"45",
		X"43",X"00",X"01",X"B0",X"D6",X"34",X"00",X"09",X"12",X"D5",X"42",X"4F",X"44",X"59",X"20",X"54",
		X"59",X"50",X"45",X"09",X"12",X"D6",X"50",X"4C",X"41",X"59",X"20",X"54",X"49",X"4D",X"45",X"0B",
		X"92",X"D6",X"43",X"4F",X"4D",X"4D",X"41",X"4E",X"44",X"4F",X"4D",X"45",X"4E",X"00",X"B2",X"74",
		X"C2",X"74",X"0C",X"30",X"D5",X"54",X"41",X"42",X"4C",X"45",X"20",X"54",X"59",X"50",X"45",X"20",
		X"20",X"00",X"0C",X"30",X"D5",X"55",X"50",X"52",X"49",X"47",X"48",X"54",X"20",X"54",X"59",X"50",
		X"45",X"00",X"0D",X"B0",X"D3",X"31",X"20",X"43",X"4F",X"49",X"4E",X"20",X"31",X"20",X"50",X"4C",
		X"41",X"59",X"00",X"0E",X"B0",X"D3",X"32",X"20",X"43",X"4F",X"49",X"4E",X"53",X"20",X"31",X"20",
		X"50",X"4C",X"41",X"59",X"00",X"0E",X"B0",X"D3",X"33",X"20",X"43",X"4F",X"49",X"4E",X"53",X"20",
		X"31",X"20",X"50",X"4C",X"41",X"59",X"00",X"0E",X"B0",X"D3",X"34",X"20",X"43",X"4F",X"49",X"4E",
		X"53",X"20",X"31",X"20",X"50",X"4C",X"41",X"59",X"00",X"0E",X"B0",X"D3",X"35",X"20",X"43",X"4F",
		X"49",X"4E",X"53",X"20",X"31",X"20",X"50",X"4C",X"41",X"59",X"00",X"0E",X"B0",X"D3",X"36",X"20",
		X"43",X"4F",X"49",X"4E",X"53",X"20",X"31",X"20",X"50",X"4C",X"41",X"59",X"00",X"0E",X"B0",X"D3",
		X"31",X"20",X"43",X"4F",X"49",X"4E",X"20",X"32",X"20",X"50",X"4C",X"41",X"59",X"53",X"00",X"0E",
		X"B0",X"D3",X"31",X"20",X"43",X"4F",X"49",X"4E",X"20",X"33",X"20",X"50",X"4C",X"41",X"59",X"53",
		X"00",X"0E",X"B0",X"D3",X"31",X"20",X"43",X"4F",X"49",X"4E",X"20",X"34",X"20",X"50",X"4C",X"41",
		X"59",X"53",X"00",X"0E",X"B0",X"D3",X"31",X"20",X"43",X"4F",X"49",X"4E",X"20",X"35",X"20",X"50",
		X"4C",X"41",X"59",X"53",X"00",X"0E",X"B0",X"D3",X"31",X"20",X"43",X"4F",X"49",X"4E",X"20",X"36",
		X"20",X"50",X"4C",X"41",X"59",X"53",X"00",X"0E",X"B0",X"D3",X"20",X"20",X"20",X"20",X"46",X"52",
		X"45",X"45",X"20",X"20",X"20",X"20",X"20",X"00",X"0E",X"B0",X"D3",X"31",X"20",X"43",X"4F",X"49",
		X"4E",X"20",X"31",X"20",X"50",X"4C",X"41",X"59",X"20",X"0E",X"30",X"D4",X"31",X"20",X"43",X"4F",
		X"49",X"4E",X"20",X"32",X"20",X"50",X"4C",X"41",X"59",X"53",X"00",X"0E",X"B0",X"D3",X"32",X"20",
		X"43",X"4F",X"49",X"4E",X"53",X"20",X"31",X"20",X"50",X"4C",X"41",X"59",X"0E",X"30",X"D4",X"31",
		X"20",X"43",X"4F",X"49",X"4E",X"20",X"33",X"20",X"50",X"4C",X"41",X"59",X"53",X"00",X"0E",X"B0",
		X"D3",X"33",X"20",X"43",X"4F",X"49",X"4E",X"53",X"20",X"31",X"20",X"50",X"4C",X"41",X"59",X"0E",
		X"30",X"D4",X"31",X"20",X"43",X"4F",X"49",X"4E",X"20",X"35",X"20",X"50",X"4C",X"41",X"59",X"53",
		X"00",X"0E",X"B0",X"D3",X"20",X"20",X"20",X"20",X"46",X"52",X"45",X"45",X"20",X"20",X"20",X"20",
		X"20",X"0E",X"30",X"D4",X"31",X"20",X"43",X"4F",X"49",X"4E",X"20",X"36",X"20",X"50",X"4C",X"41",
		X"59",X"53",X"00",X"EE",X"FF",X"06",X"08",X"23",X"36",X"04",X"2B",X"0F",X"38",X"04",X"36",X"30",
		X"18",X"02",X"36",X"31",X"23",X"23",X"23",X"23",X"10",X"ED",X"C9",X"CD",X"B6",X"77",X"21",X"00",
		X"D0",X"11",X"05",X"08",X"01",X"00",X"08",X"72",X"23",X"73",X"23",X"0B",X"78",X"B1",X"20",X"F7",
		X"21",X"00",X"E1",X"11",X"01",X"E1",X"36",X"00",X"01",X"00",X"01",X"ED",X"B0",X"FB",X"21",X"A3",
		X"76",X"11",X"00",X"E1",X"01",X"20",X"00",X"ED",X"B0",X"CD",X"95",X"79",X"CD",X"95",X"79",X"CD",
		X"95",X"79",X"DB",X"00",X"2F",X"0F",X"0F",X"30",X"F0",X"21",X"00",X"E1",X"11",X"01",X"E1",X"36",
		X"00",X"01",X"00",X"01",X"ED",X"B0",X"CD",X"95",X"79",X"CD",X"95",X"79",X"CD",X"95",X"79",X"F3",
		X"C3",X"33",X"70",X"13",X"00",X"C0",X"00",X"10",X"80",X"A0",X"00",X"13",X"00",X"40",X"01",X"10",
		X"00",X"A0",X"00",X"13",X"00",X"C0",X"00",X"10",X"C0",X"60",X"01",X"13",X"00",X"40",X"01",X"10",
		X"40",X"60",X"01",X"00",X"03",X"00",X"80",X"00",X"10",X"00",X"80",X"00",X"03",X"00",X"80",X"00",
		X"10",X"01",X"80",X"00",X"03",X"01",X"80",X"00",X"10",X"00",X"80",X"00",X"03",X"01",X"80",X"00",
		X"10",X"01",X"80",X"11",X"00",X"C0",X"01",X"00",X"01",X"ED",X"B0",X"C9",X"21",X"00",X"E1",X"11",
		X"01",X"E1",X"36",X"00",X"01",X"00",X"01",X"ED",X"B0",X"AF",X"32",X"06",X"E3",X"67",X"6F",X"22",
		X"0D",X"E7",X"CD",X"B6",X"77",X"21",X"DF",X"7A",X"CD",X"D5",X"77",X"FB",X"06",X"08",X"DB",X"00",
		X"2F",X"21",X"C0",X"D2",X"CD",X"38",X"77",X"06",X"08",X"DB",X"01",X"2F",X"21",X"C0",X"D4",X"CD",
		X"38",X"77",X"06",X"08",X"DB",X"02",X"2F",X"21",X"C0",X"D6",X"CD",X"38",X"77",X"06",X"08",X"21",
		X"40",X"D1",X"7B",X"CD",X"38",X"77",X"18",X"14",X"23",X"36",X"04",X"2B",X"0F",X"38",X"04",X"36",
		X"30",X"18",X"02",X"36",X"31",X"23",X"23",X"23",X"23",X"10",X"ED",X"C9",X"CD",X"95",X"77",X"3A",
		X"0D",X"E7",X"21",X"C0",X"D7",X"CD",X"78",X"77",X"3A",X"0E",X"E7",X"CD",X"78",X"77",X"CD",X"9E",
		X"79",X"CD",X"9E",X"79",X"DB",X"01",X"2F",X"0F",X"0F",X"38",X"02",X"18",X"9E",X"DB",X"00",X"2F",
		X"0F",X"0F",X"30",X"97",X"F3",X"C3",X"33",X"70",X"23",X"36",X"04",X"2B",X"F5",X"0F",X"0F",X"0F",
		X"0F",X"E6",X"0F",X"C6",X"30",X"77",X"23",X"23",X"23",X"36",X"04",X"2B",X"F1",X"E6",X"0F",X"C6",
		X"30",X"77",X"23",X"23",X"C9",X"21",X"0F",X"E7",X"3A",X"09",X"E0",X"E6",X"C0",X"BE",X"C8",X"32",
		X"0F",X"E7",X"3A",X"0E",X"E7",X"C6",X"01",X"27",X"32",X"0E",X"E7",X"D0",X"3A",X"0D",X"E7",X"C6",
		X"01",X"27",X"32",X"0D",X"E7",X"C9",X"21",X"00",X"D0",X"01",X"FF",X"07",X"36",X"00",X"54",X"5D",
		X"13",X"13",X"CD",X"A7",X"79",X"21",X"01",X"D0",X"01",X"FF",X"07",X"36",X"00",X"54",X"5D",X"13",
		X"13",X"CD",X"A7",X"79",X"C9",X"7E",X"FE",X"00",X"C8",X"CD",X"DE",X"77",X"18",X"F7",X"4E",X"06",
		X"00",X"23",X"5E",X"23",X"56",X"23",X"7E",X"12",X"3E",X"04",X"13",X"12",X"13",X"23",X"0D",X"20",
		X"F5",X"C9",X"21",X"00",X"E0",X"0E",X"06",X"AF",X"06",X"00",X"77",X"10",X"FD",X"0D",X"20",X"F8",
		X"C9",X"0E",X"00",X"06",X"00",X"10",X"FE",X"0D",X"20",X"F9",X"3D",X"20",X"F4",X"C9",X"C5",X"E5",
		X"77",X"23",X"10",X"FC",X"E1",X"0E",X"20",X"09",X"C1",X"0D",X"20",X"F2",X"C9",X"CD",X"B6",X"77",
		X"CD",X"36",X"78",X"CD",X"95",X"79",X"CD",X"95",X"79",X"CD",X"95",X"79",X"DB",X"00",X"2F",X"0F",
		X"0F",X"DA",X"33",X"70",X"18",X"ED",X"21",X"00",X"D0",X"01",X"FF",X"0F",X"3E",X"86",X"77",X"23",
		X"0B",X"78",X"B1",X"20",X"F7",X"21",X"0C",X"D0",X"06",X"10",X"E5",X"C5",X"CD",X"71",X"78",X"C1",
		X"E1",X"11",X"00",X"01",X"19",X"10",X"F3",X"06",X"40",X"21",X"BF",X"D7",X"7E",X"B0",X"77",X"23",
		X"23",X"7E",X"B0",X"77",X"11",X"80",X"00",X"19",X"7E",X"B0",X"77",X"2B",X"2B",X"7E",X"B0",X"77",
		X"C9",X"06",X"19",X"CD",X"7D",X"78",X"23",X"23",X"23",X"23",X"10",X"F7",X"C9",X"E5",X"3E",X"03",
		X"77",X"23",X"23",X"3E",X"02",X"77",X"E1",X"E5",X"11",X"80",X"00",X"19",X"3E",X"01",X"77",X"23",
		X"23",X"3E",X"00",X"77",X"E1",X"C9",X"F3",X"CD",X"B6",X"77",X"21",X"B3",X"79",X"CD",X"D5",X"77",
		X"CD",X"95",X"79",X"CD",X"95",X"79",X"CD",X"95",X"79",X"DB",X"00",X"2F",X"0F",X"38",X"02",X"18",
		X"EC",X"11",X"01",X"46",X"CD",X"85",X"79",X"CD",X"95",X"79",X"CD",X"95",X"79",X"CD",X"95",X"79",
		X"DB",X"00",X"2F",X"0F",X"38",X"02",X"18",X"E9",X"13",X"CD",X"85",X"79",X"CD",X"95",X"79",X"CD",
		X"95",X"79",X"CD",X"95",X"79",X"DB",X"00",X"2F",X"0F",X"38",X"02",X"18",X"EF",X"13",X"CD",X"85",
		X"79",X"CD",X"95",X"79",X"CD",X"95",X"79",X"CD",X"95",X"79",X"DB",X"00",X"2F",X"0F",X"38",X"02",
		X"18",X"EC",X"3E",X"10",X"21",X"10",X"D0",X"0E",X"03",X"11",X"01",X"46",X"06",X"10",X"73",X"23",
		X"72",X"23",X"10",X"FA",X"13",X"0D",X"20",X"F4",X"11",X"20",X"00",X"19",X"3D",X"20",X"E8",X"3E",
		X"03",X"11",X"01",X"52",X"0E",X"04",X"06",X"30",X"73",X"23",X"72",X"23",X"10",X"FA",X"D5",X"11",
		X"20",X"00",X"19",X"D1",X"0D",X"20",X"EF",X"13",X"3D",X"20",X"E9",X"11",X"01",X"49",X"0E",X"04",
		X"06",X"30",X"73",X"23",X"72",X"23",X"10",X"FA",X"D5",X"11",X"20",X"00",X"19",X"D1",X"0D",X"20",
		X"EF",X"CD",X"95",X"79",X"CD",X"95",X"79",X"CD",X"95",X"79",X"DB",X"00",X"2F",X"0F",X"38",X"02",
		X"18",X"A0",X"CD",X"95",X"79",X"CD",X"95",X"79",X"CD",X"95",X"79",X"3E",X"01",X"D3",X"01",X"CD",
		X"95",X"79",X"CD",X"95",X"79",X"CD",X"95",X"79",X"DB",X"00",X"2F",X"0F",X"30",X"F1",X"AF",X"D3",
		X"01",X"CD",X"95",X"79",X"CD",X"95",X"79",X"CD",X"95",X"79",X"DB",X"00",X"2F",X"0F",X"0F",X"DA",
		X"33",X"70",X"C3",X"71",X"79",X"21",X"00",X"D0",X"01",X"00",X"08",X"73",X"23",X"72",X"23",X"0B",
		X"78",X"B1",X"20",X"F7",X"C9",X"01",X"00",X"40",X"0B",X"78",X"B1",X"20",X"FB",X"C9",X"01",X"00",
		X"90",X"0B",X"78",X"B1",X"20",X"FB",X"C9",X"7E",X"12",X"23",X"23",X"13",X"13",X"0B",X"78",X"B1",
		X"20",X"F5",X"C9",X"0E",X"A0",X"D1",X"41",X"20",X"42",X"20",X"43",X"20",X"44",X"20",X"45",X"20",
		X"46",X"20",X"47",X"20",X"0E",X"20",X"D2",X"48",X"20",X"49",X"20",X"4A",X"20",X"4B",X"20",X"4C",
		X"20",X"4D",X"20",X"4E",X"20",X"0E",X"A0",X"D2",X"4F",X"20",X"50",X"20",X"51",X"20",X"52",X"20",
		X"53",X"20",X"54",X"20",X"55",X"20",X"0E",X"20",X"D3",X"56",X"20",X"57",X"20",X"58",X"20",X"59",
		X"20",X"5A",X"20",X"20",X"20",X"20",X"20",X"14",X"A0",X"D3",X"31",X"20",X"32",X"20",X"33",X"20",
		X"34",X"20",X"35",X"20",X"36",X"20",X"37",X"20",X"38",X"20",X"39",X"20",X"30",X"20",X"00",X"08",
		X"A0",X"D0",X"52",X"41",X"4D",X"20",X"20",X"20",X"4F",X"4B",X"00",X"10",X"A0",X"D0",X"52",X"41",
		X"4D",X"20",X"20",X"20",X"4E",X"47",X"20",X"20",X"28",X"20",X"20",X"20",X"20",X"29",X"00",X"52",
		X"4F",X"4D",X"20",X"20",X"20",X"4F",X"4B",X"00",X"52",X"4F",X"4D",X"20",X"20",X"20",X"4E",X"47",
		X"00",X"16",X"A0",X"D0",X"44",X"49",X"50",X"20",X"53",X"57",X"20",X"31",X"20",X"32",X"20",X"33",
		X"20",X"34",X"20",X"35",X"20",X"36",X"20",X"37",X"20",X"38",X"03",X"A0",X"D1",X"53",X"57",X"31",
		X"03",X"A0",X"D2",X"53",X"57",X"32",X"00",X"01",X"98",X"D2",X"20",X"1B",X"C4",X"D2",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"00",X"0C",X"A0",X"D0",X"49",X"4E",X"54",
		X"45",X"52",X"46",X"41",X"43",X"45",X"20",X"4F",X"4B",X"00",X"A0",X"7A",X"B5",X"7A",X"CA",X"7A",
		X"11",X"A0",X"D0",X"43",X"48",X"45",X"43",X"4B",X"20",X"49",X"4E",X"54",X"45",X"52",X"46",X"41",
		X"43",X"45",X"20",X"31",X"00",X"11",X"A0",X"D0",X"43",X"48",X"45",X"43",X"4B",X"20",X"49",X"4E",
		X"54",X"45",X"52",X"46",X"41",X"43",X"45",X"20",X"32",X"00",X"11",X"A0",X"D0",X"43",X"48",X"45",
		X"43",X"4B",X"20",X"49",X"4E",X"54",X"45",X"52",X"46",X"41",X"43",X"45",X"20",X"33",X"00",X"0A",
		X"20",X"D1",X"57",X"52",X"49",X"54",X"45",X"20",X"44",X"41",X"54",X"41",X"0C",X"20",X"D2",X"49",
		X"4E",X"54",X"45",X"52",X"46",X"41",X"43",X"45",X"20",X"31",X"20",X"0C",X"A0",X"D2",X"20",X"20",
		X"20",X"52",X"45",X"41",X"44",X"20",X"44",X"41",X"54",X"41",X"0C",X"20",X"D4",X"49",X"4E",X"54",
		X"45",X"52",X"46",X"41",X"43",X"45",X"20",X"32",X"20",X"0C",X"A0",X"D4",X"20",X"20",X"20",X"52",
		X"45",X"41",X"44",X"20",X"44",X"41",X"54",X"41",X"0C",X"20",X"D6",X"49",X"4E",X"54",X"45",X"52",
		X"46",X"41",X"43",X"45",X"20",X"33",X"20",X"0C",X"A0",X"D6",X"20",X"20",X"20",X"52",X"45",X"41",
		X"44",X"20",X"44",X"41",X"54",X"41",X"0F",X"40",X"D2",X"30",X"20",X"31",X"20",X"32",X"20",X"33",
		X"20",X"34",X"20",X"35",X"20",X"36",X"20",X"37",X"0F",X"40",X"D4",X"30",X"20",X"31",X"20",X"32",
		X"20",X"33",X"20",X"34",X"20",X"35",X"20",X"36",X"20",X"37",X"0F",X"40",X"D6",X"30",X"20",X"31",
		X"20",X"32",X"20",X"33",X"20",X"34",X"20",X"35",X"20",X"36",X"20",X"37",X"0F",X"40",X"D1",X"30",
		X"20",X"31",X"20",X"32",X"20",X"33",X"20",X"34",X"20",X"35",X"20",X"36",X"20",X"37",X"06",X"A0",
		X"D7",X"54",X"49",X"4D",X"49",X"4E",X"47",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"72",
		X"EC",X"76",X"5E",X"7C",X"4B",X"76",X"96",X"78",X"1D",X"78",X"0D",X"20",X"D1",X"30",X"31",X"20",
		X"44",X"49",X"50",X"20",X"53",X"57",X"49",X"54",X"43",X"48",X"0B",X"A0",X"D1",X"30",X"32",X"20",
		X"49",X"2F",X"4F",X"20",X"50",X"4F",X"52",X"54",X"08",X"20",X"D2",X"30",X"33",X"20",X"53",X"4F",
		X"55",X"4E",X"44",X"0C",X"A0",X"D2",X"30",X"34",X"20",X"43",X"48",X"41",X"52",X"41",X"43",X"54",
		X"45",X"52",X"08",X"20",X"D3",X"30",X"35",X"20",X"43",X"4F",X"4C",X"4F",X"52",X"16",X"A0",X"D3",
		X"30",X"36",X"20",X"43",X"52",X"4F",X"53",X"53",X"20",X"48",X"41",X"54",X"43",X"48",X"20",X"50",
		X"41",X"54",X"54",X"45",X"52",X"4E",X"00",X"7C",X"B8",X"C0",X"7D",X"B9",X"C9",X"21",X"00",X"80",
		X"01",X"00",X"08",X"AF",X"77",X"23",X"0B",X"78",X"B1",X"20",X"F8",X"C9",X"72",X"23",X"0B",X"78",
		X"B1",X"20",X"F9",X"C9",X"72",X"23",X"23",X"0B",X"78",X"B1",X"20",X"F8",X"C9",X"08",X"D9",X"C3",
		X"39",X"7C",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"21",X"09",X"E0",X"34",X"CD",X"52",X"7C",
		X"3A",X"02",X"E3",X"0F",X"38",X"07",X"21",X"06",X"E3",X"3E",X"80",X"86",X"77",X"C9",X"D9",X"08",
		X"FB",X"C9",X"21",X"00",X"E1",X"11",X"00",X"C0",X"01",X"00",X"01",X"ED",X"B0",X"C9",X"CD",X"B6",
		X"77",X"21",X"B9",X"7D",X"CD",X"D5",X"77",X"2A",X"9C",X"7D",X"22",X"06",X"E7",X"DD",X"21",X"08",
		X"E7",X"FD",X"21",X"A0",X"7D",X"CD",X"95",X"79",X"CD",X"95",X"79",X"CD",X"95",X"79",X"CD",X"8B",
		X"7C",X"DB",X"00",X"2F",X"0F",X"0F",X"DA",X"33",X"70",X"18",X"D3",X"FD",X"22",X"0B",X"E7",X"3E",
		X"01",X"32",X"05",X"E7",X"06",X"06",X"CD",X"50",X"7D",X"CD",X"E5",X"7C",X"CD",X"CF",X"7C",X"01",
		X"00",X"00",X"ED",X"43",X"13",X"E3",X"DB",X"00",X"2F",X"0F",X"0F",X"30",X"04",X"C1",X"C3",X"33",
		X"70",X"DB",X"00",X"2F",X"0F",X"DC",X"CF",X"7C",X"DB",X"01",X"2F",X"0F",X"38",X"34",X"0F",X"38",
		X"5D",X"ED",X"4B",X"13",X"E3",X"0B",X"78",X"B1",X"20",X"D8",X"CD",X"E5",X"7C",X"18",X"4F",X"3A",
		X"05",X"E7",X"4F",X"06",X"00",X"FD",X"2A",X"0B",X"E7",X"FD",X"09",X"FD",X"7E",X"00",X"D3",X"00",
		X"F6",X"80",X"D3",X"00",X"C9",X"3E",X"00",X"D3",X"00",X"3E",X"80",X"D3",X"00",X"06",X"00",X"10",
		X"FE",X"C9",X"CD",X"E5",X"7C",X"CD",X"95",X"79",X"CD",X"95",X"79",X"CD",X"95",X"79",X"3A",X"07",
		X"E7",X"5F",X"3A",X"05",X"E7",X"BB",X"C8",X"06",X"04",X"CD",X"50",X"7D",X"3D",X"32",X"05",X"E7",
		X"06",X"06",X"CD",X"50",X"7D",X"CD",X"CF",X"7C",X"01",X"00",X"00",X"C3",X"A2",X"7C",X"CD",X"E5",
		X"7C",X"CD",X"95",X"79",X"CD",X"95",X"79",X"CD",X"95",X"79",X"3A",X"06",X"E7",X"5F",X"3A",X"05",
		X"E7",X"BB",X"C8",X"06",X"04",X"CD",X"50",X"7D",X"3C",X"32",X"05",X"E7",X"06",X"06",X"CD",X"50",
		X"7D",X"CD",X"CF",X"7C",X"01",X"00",X"00",X"C3",X"A2",X"7C",X"4F",X"D6",X"03",X"3C",X"18",X"17",
		X"4F",X"C5",X"21",X"20",X"D1",X"11",X"80",X"00",X"47",X"05",X"28",X"03",X"19",X"18",X"FA",X"C1",
		X"23",X"70",X"23",X"23",X"70",X"79",X"C9",X"C5",X"21",X"20",X"D1",X"11",X"80",X"00",X"47",X"FE",
		X"01",X"28",X"04",X"05",X"19",X"10",X"FD",X"C1",X"23",X"70",X"23",X"23",X"70",X"79",X"C9",X"C5",
		X"0E",X"00",X"06",X"00",X"10",X"FE",X"F5",X"3A",X"00",X"D0",X"CB",X"4F",X"28",X"09",X"F1",X"0D",
		X"20",X"F0",X"3D",X"20",X"EB",X"C1",X"C9",X"F1",X"C1",X"06",X"01",X"C9",X"15",X"01",X"00",X"00",
		X"00",X"01",X"02",X"03",X"04",X"05",X"06",X"1C",X"11",X"12",X"13",X"14",X"15",X"20",X"21",X"22",
		X"23",X"24",X"25",X"26",X"27",X"00",X"00",X"00",X"00",X"0B",X"A0",X"D0",X"53",X"20",X"4F",X"20",
		X"55",X"20",X"4E",X"20",X"44",X"20",X"53",X"0F",X"20",X"D1",X"30",X"31",X"20",X"48",X"4F",X"4C",
		X"45",X"20",X"44",X"49",X"47",X"47",X"49",X"4E",X"47",X"15",X"A0",X"D1",X"30",X"32",X"20",X"50",
		X"49",X"43",X"4B",X"49",X"4E",X"47",X"20",X"55",X"50",X"20",X"46",X"4F",X"52",X"54",X"49",X"4E",
		X"45",X"0F",X"20",X"D2",X"30",X"33",X"20",X"44",X"4F",X"4F",X"52",X"20",X"4F",X"50",X"45",X"4E",
		X"49",X"4E",X"47",X"13",X"A0",X"D2",X"30",X"34",X"20",X"42",X"55",X"52",X"49",X"45",X"44",X"20",
		X"49",X"4E",X"54",X"4F",X"20",X"48",X"4F",X"4C",X"45",X"14",X"20",X"D3",X"30",X"35",X"20",X"46",
		X"41",X"4C",X"4C",X"49",X"4E",X"47",X"20",X"49",X"4E",X"54",X"4F",X"20",X"48",X"4F",X"4C",X"45",
		X"10",X"A0",X"D3",X"30",X"36",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"20",X"4B",X"49",X"4C",
		X"4C",X"45",X"44",X"12",X"20",X"D4",X"30",X"37",X"20",X"54",X"49",X"4D",X"45",X"20",X"55",X"50",
		X"20",X"57",X"41",X"52",X"4E",X"49",X"4E",X"47",X"16",X"A0",X"D4",X"30",X"38",X"20",X"54",X"49",
		X"4D",X"45",X"20",X"53",X"43",X"4F",X"52",X"45",X"20",X"43",X"4F",X"55",X"4E",X"54",X"49",X"4E",
		X"47",X"11",X"20",X"D5",X"30",X"39",X"20",X"43",X"4F",X"49",X"4E",X"20",X"49",X"4E",X"53",X"45",
		X"52",X"54",X"49",X"4E",X"47",X"0F",X"A0",X"D5",X"31",X"30",X"20",X"5A",X"4F",X"4F",X"4D",X"20",
		X"49",X"4E",X"20",X"20",X"20",X"20",X"20",X"0F",X"20",X"D6",X"31",X"31",X"20",X"5A",X"4F",X"4F",
		X"4D",X"20",X"4F",X"55",X"54",X"20",X"20",X"20",X"20",X"16",X"A0",X"D6",X"31",X"32",X"20",X"50",
		X"4C",X"41",X"59",X"45",X"52",X"20",X"46",X"41",X"4C",X"4C",X"49",X"4E",X"47",X"20",X"20",X"20",
		X"20",X"20",X"0D",X"20",X"D7",X"31",X"33",X"20",X"47",X"41",X"4D",X"45",X"20",X"53",X"54",X"41",
		X"52",X"54",X"0C",X"A0",X"D7",X"31",X"34",X"20",X"47",X"41",X"4D",X"45",X"20",X"4F",X"56",X"45",
		X"52",X"1B",X"20",X"D8",X"31",X"35",X"20",X"42",X"47",X"4D",X"20",X"28",X"43",X"4F",X"4E",X"54",
		X"49",X"4E",X"55",X"49",X"54",X"59",X"20",X"44",X"49",X"53",X"50",X"4C",X"41",X"59",X"29",X"0E",
		X"A0",X"D8",X"31",X"36",X"20",X"52",X"4F",X"55",X"4E",X"44",X"20",X"43",X"4C",X"45",X"41",X"52",
		X"0E",X"20",X"D9",X"31",X"37",X"20",X"42",X"4C",X"4F",X"43",X"4B",X"20",X"43",X"4C",X"45",X"41",
		X"52",X"0D",X"A0",X"D9",X"31",X"38",X"20",X"54",X"49",X"4D",X"45",X"20",X"55",X"50",X"20",X"20",
		X"20",X"12",X"20",X"DA",X"31",X"39",X"20",X"42",X"47",X"4D",X"20",X"28",X"47",X"41",X"4D",X"45",
		X"20",X"50",X"4C",X"41",X"59",X"29",X"12",X"A0",X"DA",X"32",X"30",X"20",X"47",X"41",X"4D",X"45",
		X"20",X"43",X"4F",X"4D",X"50",X"4C",X"45",X"54",X"49",X"4E",X"47",X"0C",X"20",X"DB",X"20",X"20",
		X"4D",X"55",X"53",X"49",X"43",X"20",X"45",X"4E",X"44",X"20",X"00",X"00",X"00",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
