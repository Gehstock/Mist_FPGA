`define BUILD_DATE "210618"
`define BUILD_TIME "214731"
