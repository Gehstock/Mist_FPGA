library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_7L is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_7L is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"1E",X"0F",X"13",X"13",X"6E",X"00",X"00",X"30",X"1B",X"89",X"C1",X"B1",X"8F",
		X"7E",X"62",X"62",X"32",X"1C",X"00",X"00",X"00",X"87",X"31",X"3D",X"CB",X"4B",X"30",X"00",X"00",
		X"00",X"00",X"00",X"3C",X"1E",X"26",X"26",X"DC",X"00",X"0C",X"36",X"4B",X"8F",X"CC",X"B0",X"84",
		X"FC",X"C4",X"C4",X"64",X"38",X"00",X"00",X"00",X"84",X"16",X"2B",X"CD",X"4C",X"2C",X"08",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"1E",X"02",X"00",X"00",X"00",X"00",X"08",X"28",X"29",X"D9",
		X"12",X"72",X"6C",X"78",X"7C",X"3E",X"1C",X"00",X"AF",X"AB",X"EB",X"6F",X"7F",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"1E",X"02",X"00",X"00",X"00",X"00",X"0A",X"2A",X"29",X"D9",
		X"12",X"72",X"6C",X"78",X"7C",X"3E",X"1C",X"00",X"A9",X"AC",X"AB",X"69",X"79",X"39",X"07",X"00",
		X"00",X"00",X"00",X"00",X"00",X"12",X"1E",X"02",X"00",X"00",X"00",X"03",X"0F",X"2B",X"29",X"DD",
		X"12",X"72",X"6C",X"78",X"7C",X"3E",X"1C",X"00",X"AF",X"AC",X"EF",X"69",X"79",X"09",X"0D",X"0E",
		X"00",X"1C",X"3E",X"7C",X"78",X"6C",X"72",X"12",X"00",X"00",X"00",X"7F",X"6F",X"EB",X"AB",X"AF",
		X"1E",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"D9",X"29",X"28",X"08",X"00",X"00",X"00",X"00",
		X"00",X"1C",X"3E",X"7C",X"78",X"6C",X"72",X"12",X"00",X"07",X"39",X"79",X"69",X"AB",X"AC",X"A9",
		X"1E",X"02",X"12",X"00",X"00",X"00",X"00",X"00",X"D9",X"29",X"2A",X"0A",X"00",X"00",X"00",X"00",
		X"00",X"1C",X"3E",X"7C",X"78",X"6C",X"72",X"12",X"0E",X"0D",X"09",X"79",X"69",X"EF",X"AC",X"AF",
		X"1E",X"02",X"12",X"00",X"00",X"00",X"00",X"00",X"DD",X"29",X"29",X"0D",X"03",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"07",X"04",X"04",X"00",X"00",X"00",X"00",X"60",X"F0",X"90",X"90",
		X"04",X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"90",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"07",X"0F",X"18",X"30",X"24",X"04",X"00",X"00",X"F0",X"F0",X"00",X"00",X"90",X"90",
		X"04",X"07",X"07",X"07",X"00",X"00",X"00",X"00",X"90",X"F8",X"F8",X"F0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"F0",X"0E",X"0E",
		X"00",X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"0E",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"07",X"0F",X"1B",X"3F",X"3C",X"34",X"00",X"00",X"F0",X"F8",X"6C",X"FE",X"9E",X"96",
		X"34",X"3F",X"3F",X"1F",X"08",X"00",X"00",X"00",X"96",X"FE",X"FE",X"FC",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"04",X"04",X"04",X"00",X"00",X"00",X"00",X"10",X"90",X"90",X"90",
		X"04",X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"90",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"07",X"0F",X"18",X"30",X"24",X"04",X"00",X"00",X"F0",X"F0",X"00",X"00",X"90",X"90",
		X"04",X"07",X"07",X"07",X"00",X"00",X"00",X"00",X"90",X"F8",X"F8",X"F0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"90",X"0E",X"0E",
		X"00",X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"0E",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"07",X"0F",X"1C",X"3C",X"3C",X"34",X"00",X"00",X"F0",X"F8",X"1C",X"9E",X"9E",X"96",
		X"34",X"3F",X"3F",X"1F",X"08",X"00",X"00",X"00",X"96",X"FE",X"FE",X"FC",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"06",X"04",X"04",X"00",X"00",X"00",X"00",X"60",X"F0",X"90",X"90",
		X"04",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"90",X"B0",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"07",X"0F",X"18",X"30",X"24",X"04",X"00",X"00",X"F0",X"F0",X"00",X"00",X"90",X"90",
		X"04",X"07",X"07",X"07",X"00",X"00",X"00",X"00",X"90",X"B8",X"F8",X"F0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"F0",X"0E",X"0E",
		X"00",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"0E",X"B0",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"07",X"0F",X"1A",X"3E",X"3C",X"34",X"00",X"00",X"F0",X"F8",X"6C",X"FE",X"9E",X"96",
		X"34",X"3F",X"3F",X"1F",X"08",X"00",X"00",X"00",X"96",X"BE",X"FE",X"FC",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"E0",X"70",X"7A",X"C7",X"C7",X"00",X"00",X"1C",X"1C",X"3C",X"24",X"20",X"20",
		X"FF",X"C7",X"C7",X"7A",X"70",X"E0",X"00",X"00",X"24",X"20",X"20",X"24",X"3C",X"1C",X"18",X"00",
		X"00",X"00",X"00",X"E1",X"70",X"7E",X"C7",X"C7",X"00",X"18",X"FC",X"FC",X"F8",X"24",X"20",X"20",
		X"FF",X"C7",X"C7",X"7E",X"70",X"E0",X"00",X"00",X"24",X"20",X"20",X"24",X"FC",X"F8",X"38",X"08",
		X"00",X"00",X"00",X"1C",X"0E",X"0F",X"18",X"38",X"00",X"00",X"00",X"06",X"02",X"D0",X"D0",X"D4",
		X"3E",X"38",X"18",X"0F",X"0E",X"1C",X"00",X"00",X"D6",X"D4",X"D0",X"D0",X"02",X"06",X"00",X"00",
		X"00",X"00",X"00",X"24",X"46",X"E7",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"20",X"24",X"2C",
		X"FF",X"7D",X"78",X"E0",X"00",X"00",X"00",X"00",X"24",X"20",X"20",X"30",X"38",X"1C",X"0C",X"00",
		X"00",X"00",X"00",X"24",X"46",X"E7",X"FF",X"FF",X"00",X"00",X"00",X"00",X"20",X"20",X"A0",X"20",
		X"FF",X"7D",X"78",X"E0",X"00",X"00",X"00",X"00",X"20",X"00",X"04",X"84",X"7C",X"3C",X"18",X"00",
		X"00",X"00",X"00",X"24",X"46",X"E7",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"20",X"A0",X"20",
		X"FF",X"7D",X"79",X"E0",X"00",X"00",X"00",X"00",X"20",X"A0",X"E0",X"F8",X"3C",X"08",X"00",X"00",
		X"00",X"00",X"00",X"24",X"46",X"E7",X"FF",X"FF",X"00",X"00",X"00",X"00",X"20",X"20",X"20",X"20",
		X"FF",X"7D",X"79",X"F0",X"00",X"00",X"00",X"00",X"00",X"04",X"9C",X"FC",X"7C",X"18",X"00",X"00",
		X"00",X"00",X"00",X"00",X"F0",X"78",X"7D",X"FF",X"00",X"0C",X"1C",X"38",X"30",X"20",X"20",X"24",
		X"FF",X"FF",X"E7",X"46",X"24",X"00",X"00",X"00",X"2C",X"24",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"F0",X"78",X"7D",X"FF",X"00",X"18",X"3C",X"7C",X"84",X"04",X"00",X"20",
		X"FF",X"FF",X"E7",X"46",X"24",X"00",X"00",X"00",X"20",X"20",X"20",X"20",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"F0",X"79",X"7D",X"FF",X"00",X"00",X"08",X"3C",X"F8",X"E0",X"A0",X"20",
		X"FF",X"FF",X"E7",X"46",X"24",X"00",X"00",X"00",X"20",X"20",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"F0",X"79",X"7D",X"FF",X"00",X"00",X"18",X"7C",X"9C",X"9C",X"04",X"00",
		X"FF",X"FF",X"E7",X"46",X"24",X"00",X"00",X"00",X"20",X"20",X"20",X"20",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"70",X"38",X"3F",X"63",X"E3",X"00",X"06",X"1E",X"3C",X"7E",X"12",X"90",X"90",
		X"FF",X"E3",X"63",X"3F",X"38",X"70",X"00",X"00",X"92",X"90",X"90",X"12",X"7C",X"3E",X"0E",X"00",
		X"00",X"60",X"78",X"FC",X"FE",X"7F",X"F1",X"F1",X"00",X"00",X"00",X"00",X"00",X"88",X"C8",X"C8",
		X"FF",X"F1",X"F1",X"7F",X"FE",X"FC",X"78",X"00",X"C8",X"C8",X"C8",X"88",X"00",X"00",X"00",X"00",
		X"00",X"00",X"3D",X"47",X"C7",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"90",X"10",X"B0",X"A0",
		X"7F",X"3F",X"3A",X"70",X"01",X"00",X"00",X"00",X"A2",X"22",X"62",X"32",X"38",X"1C",X"3E",X"1C",
		X"00",X"00",X"00",X"00",X"E0",X"78",X"46",X"C6",X"00",X"00",X"00",X"00",X"00",X"40",X"64",X"22",
		X"FF",X"E3",X"E3",X"FF",X"7E",X"3D",X"38",X"70",X"20",X"20",X"20",X"26",X"26",X"06",X"86",X"3C",
		X"00",X"00",X"00",X"01",X"00",X"72",X"3F",X"3F",X"1C",X"3E",X"1C",X"38",X"32",X"62",X"22",X"A2",
		X"7F",X"FF",X"FF",X"C7",X"47",X"3D",X"00",X"00",X"A0",X"B0",X"10",X"90",X"00",X"00",X"00",X"00",
		X"70",X"38",X"3D",X"7E",X"FF",X"E3",X"E3",X"FE",X"3C",X"86",X"06",X"2E",X"26",X"20",X"20",X"20",
		X"C7",X"46",X"78",X"E0",X"00",X"00",X"00",X"00",X"22",X"64",X"40",X"00",X"00",X"00",X"00",X"00",
		X"40",X"46",X"47",X"67",X"67",X"66",X"76",X"74",X"F3",X"0C",X"30",X"C0",X"C0",X"40",X"40",X"40",
		X"78",X"7C",X"7C",X"7C",X"19",X"07",X"04",X"04",X"40",X"00",X"00",X"00",X"00",X"80",X"A0",X"30",
		X"03",X"22",X"25",X"36",X"36",X"38",X"3C",X"3C",X"E0",X"18",X"8E",X"70",X"40",X"40",X"40",X"40",
		X"3C",X"3C",X"3C",X"1E",X"01",X"07",X"04",X"04",X"40",X"00",X"00",X"00",X"00",X"80",X"A0",X"30",
		X"03",X"16",X"1F",X"1B",X"1C",X"1E",X"1E",X"1F",X"80",X"40",X"A0",X"E8",X"9C",X"C0",X"40",X"40",
		X"1F",X"1F",X"1C",X"1C",X"01",X"07",X"04",X"04",X"40",X"00",X"00",X"00",X"00",X"80",X"E0",X"30",
		X"10",X"30",X"20",X"60",X"7F",X"1F",X"04",X"04",X"00",X"00",X"00",X"00",X"80",X"C0",X"FC",X"10",
		X"0C",X"17",X"30",X"60",X"20",X"30",X"10",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"0C",X"18",X"18",X"1F",X"0F",X"04",X"04",X"00",X"00",X"00",X"00",X"80",X"C0",X"F8",X"10",
		X"0C",X"0F",X"18",X"18",X"18",X"0C",X"06",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"16",X"18",X"18",X"1F",X"0F",X"04",X"04",X"00",X"00",X"00",X"00",X"80",X"C0",X"F0",X"10",
		X"0C",X"0F",X"18",X"18",X"18",X"1E",X"07",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"80",X"00",
		X"40",X"47",X"67",X"64",X"74",X"7C",X"7E",X"7E",X"00",X"00",X"88",X"E0",X"40",X"40",X"40",X"40",
		X"1E",X"07",X"05",X"16",X"24",X"04",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"20",X"00",X"00",
		X"00",X"00",X"04",X"24",X"16",X"05",X"07",X"1E",X"00",X"00",X"20",X"40",X"80",X"00",X"00",X"00",
		X"7E",X"7E",X"7C",X"74",X"64",X"67",X"47",X"40",X"40",X"40",X"40",X"40",X"E0",X"88",X"00",X"00",
		X"00",X"00",X"00",X"E0",X"70",X"7E",X"C7",X"C7",X"00",X"00",X"0C",X"1C",X"1C",X"04",X"20",X"20",
		X"FF",X"C7",X"C7",X"7E",X"70",X"E0",X"00",X"00",X"24",X"20",X"20",X"04",X"1C",X"1C",X"08",X"00",
		X"00",X"00",X"00",X"70",X"38",X"3C",X"7E",X"FF",X"00",X"1C",X"3C",X"70",X"70",X"20",X"20",X"24",
		X"C7",X"C7",X"FF",X"44",X"78",X"F0",X"00",X"00",X"24",X"24",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"E1",X"70",X"7E",X"C3",X"C3",X"00",X"18",X"FC",X"FC",X"F8",X"24",X"20",X"20",
		X"FB",X"C3",X"C3",X"7E",X"70",X"E0",X"00",X"00",X"24",X"20",X"20",X"24",X"FC",X"F8",X"38",X"08",
		X"00",X"03",X"01",X"01",X"01",X"03",X"02",X"3C",X"00",X"E0",X"F0",X"F8",X"BC",X"24",X"20",X"F0",
		X"7C",X"7E",X"7E",X"3F",X"1F",X"0F",X"02",X"00",X"F0",X"60",X"64",X"3C",X"08",X"60",X"00",X"00",
		X"00",X"03",X"01",X"01",X"01",X"03",X"02",X"3C",X"00",X"E0",X"F1",X"FF",X"BC",X"24",X"21",X"F0",
		X"7C",X"7E",X"7E",X"3F",X"1F",X"0F",X"02",X"00",X"F0",X"60",X"64",X"3C",X"08",X"61",X"00",X"00",
		X"00",X"03",X"01",X"00",X"00",X"00",X"00",X"38",X"00",X"E0",X"F0",X"78",X"3C",X"24",X"00",X"10",
		X"7C",X"7E",X"7E",X"3F",X"1F",X"0F",X"02",X"00",X"10",X"00",X"04",X"0C",X"08",X"00",X"00",X"00",
		X"00",X"07",X"03",X"1B",X"27",X"76",X"64",X"79",X"00",X"CA",X"E4",X"F8",X"78",X"48",X"40",X"E0",
		X"F9",X"FC",X"FC",X"7E",X"3E",X"1E",X"04",X"00",X"E0",X"C0",X"C8",X"78",X"1C",X"C4",X"0A",X"00",
		X"00",X"90",X"08",X"27",X"30",X"20",X"08",X"1C",X"00",X"02",X"04",X"0A",X"44",X"62",X"00",X"39",
		X"0C",X"0B",X"03",X"06",X"00",X"00",X"00",X"00",X"79",X"89",X"09",X"02",X"02",X"C0",X"D0",X"00",
		X"00",X"B0",X"44",X"67",X"10",X"10",X"18",X"18",X"00",X"00",X"02",X"04",X"C2",X"54",X"00",X"39",
		X"04",X"07",X"07",X"06",X"01",X"01",X"00",X"00",X"79",X"89",X"09",X"02",X"82",X"80",X"10",X"00",
		X"00",X"B0",X"4C",X"46",X"11",X"30",X"18",X"14",X"00",X"00",X"00",X"02",X"C4",X"32",X"00",X"39",
		X"04",X"0C",X"05",X"06",X"00",X"00",X"00",X"00",X"49",X"89",X"09",X"C2",X"C2",X"00",X"30",X"00",
		X"00",X"A0",X"4C",X"41",X"31",X"30",X"14",X"0C",X"00",X"00",X"00",X"00",X"82",X"70",X"00",X"39",
		X"0C",X"0D",X"03",X"02",X"00",X"00",X"00",X"00",X"79",X"89",X"09",X"02",X"62",X"60",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"0F",X"07",X"00",X"39",X"3A",X"00",X"00",X"80",X"80",X"80",X"00",X"1C",X"7C",
		X"3B",X"30",X"00",X"01",X"01",X"01",X"00",X"00",X"7C",X"1C",X"00",X"E0",X"F0",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"07",X"08",X"18",X"20",X"23",X"22",X"00",X"00",X"E0",X"10",X"28",X"24",X"F4",X"74",
		X"20",X"23",X"22",X"10",X"08",X"07",X"00",X"00",X"74",X"F4",X"64",X"28",X"10",X"E0",X"00",X"00",
		X"00",X"00",X"04",X"04",X"04",X"04",X"04",X"0C",X"00",X"80",X"C0",X"40",X"40",X"40",X"40",X"C0",
		X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"00",X"00",X"00",X"00",X"0C",X"0C",X"00",X"C0",X"00",X"00",X"00",X"00",X"C0",X"C0",X"00",
		X"00",X"00",X"00",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"00",X"00",X"00",
		X"0C",X"0C",X"00",X"00",X"00",X"00",X"0C",X"0C",X"C0",X"C0",X"00",X"00",X"00",X"00",X"40",X"C0",
		X"00",X"00",X"00",X"00",X"0C",X"0C",X"00",X"0C",X"C0",X"80",X"00",X"00",X"C0",X"C0",X"00",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"13",X"33",X"20",X"20",X"20",X"20",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"13",X"31",X"21",X"21",X"31",X"13",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"20",X"20",X"33",X"33",X"20",X"20",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"20",X"20",X"20",X"00",X"12",X"32",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"21",X"21",X"21",X"33",X"33",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"32",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"00",X"00",X"00",X"20",X"20",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"E1",X"70",X"7E",X"C7",X"C7",X"00",X"18",X"FC",X"FC",X"F8",X"24",X"20",X"20",
		X"FF",X"C7",X"C7",X"7E",X"70",X"E0",X"00",X"00",X"24",X"20",X"20",X"24",X"FC",X"F8",X"38",X"08",
		X"00",X"00",X"00",X"1C",X"0E",X"1F",X"3E",X"3E",X"00",X"18",X"0C",X"0C",X"5E",X"26",X"20",X"20",
		X"3F",X"3E",X"3E",X"1F",X"0E",X"1C",X"00",X"00",X"A4",X"20",X"20",X"26",X"5E",X"0C",X"0C",X"18",
		X"00",X"18",X"3F",X"3F",X"1F",X"3F",X"1F",X"3F",X"00",X"00",X"00",X"C0",X"E0",X"F0",X"88",X"88",
		X"3F",X"1F",X"3F",X"3F",X"1F",X"3F",X"3F",X"18",X"F8",X"88",X"88",X"F0",X"E0",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"00",X"06",X"07",X"0E",X"1F",X"1F",X"0F",X"1E",
		X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"0F",X"1F",X"1F",X"0E",X"1F",X"0F",X"07",X"02",
		X"00",X"00",X"00",X"70",X"38",X"3D",X"63",X"E3",X"00",X"04",X"1C",X"1C",X"04",X"00",X"A0",X"A0",
		X"FF",X"E3",X"63",X"3D",X"38",X"70",X"00",X"00",X"A0",X"A0",X"A0",X"00",X"04",X"1C",X"3C",X"18",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"0F",X"00",X"00",X"00",X"30",X"7C",X"00",X"C0",X"F0",X"F8",X"3C",X"1C",X"0E",X"0E",
		X"7F",X"7F",X"3F",X"3F",X"1F",X"0F",X"03",X"00",X"06",X"06",X"84",X"84",X"C0",X"C0",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"11",X"09",X"03",X"00",X"00",X"00",X"00",X"80",X"80",X"F8",X"FC",X"E0",X"FE",X"BE",
		X"14",X"16",X"1E",X"0F",X"07",X"01",X"01",X"01",X"BE",X"BE",X"FE",X"C0",X"60",X"78",X"80",X"80",
		X"00",X"00",X"00",X"01",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"FC",X"F0",X"DC",X"BF",
		X"1C",X"1E",X"1E",X"0F",X"07",X"01",X"01",X"00",X"BE",X"FE",X"DC",X"C4",X"60",X"78",X"80",X"00",
		X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"FC",X"E8",X"DC",X"BE",
		X"1C",X"1E",X"1E",X"0F",X"07",X"00",X"00",X"00",X"FF",X"BE",X"DC",X"C8",X"60",X"38",X"00",X"00",
		X"00",X"00",X"01",X"41",X"23",X"10",X"00",X"00",X"00",X"00",X"80",X"F8",X"FC",X"E4",X"DC",X"FE",
		X"1C",X"16",X"16",X"07",X"07",X"01",X"00",X"00",X"BE",X"BF",X"9C",X"D0",X"60",X"78",X"00",X"00",
		X"00",X"00",X"06",X"0E",X"1F",X"1F",X"3F",X"3F",X"00",X"00",X"10",X"18",X"DC",X"FC",X"FE",X"FE",
		X"3F",X"3F",X"1F",X"1F",X"0F",X"07",X"00",X"00",X"FE",X"FE",X"FC",X"FC",X"F8",X"F0",X"00",X"00",
		X"00",X"01",X"04",X"0E",X"1E",X"1E",X"3F",X"3F",X"00",X"C0",X"10",X"18",X"1C",X"1C",X"DE",X"FE",
		X"3F",X"3F",X"1F",X"1F",X"0F",X"07",X"01",X"00",X"FE",X"FE",X"FC",X"FC",X"F8",X"F0",X"C0",X"00",
		X"00",X"01",X"07",X"0F",X"1C",X"1E",X"3E",X"3E",X"00",X"C0",X"F0",X"F8",X"1C",X"1C",X"1E",X"1E",
		X"3F",X"3F",X"1F",X"1F",X"0F",X"07",X"01",X"00",X"DE",X"FE",X"FC",X"FC",X"F8",X"F0",X"C0",X"00",
		X"00",X"01",X"07",X"0F",X"1F",X"1F",X"3C",X"3E",X"00",X"C0",X"F0",X"F8",X"FC",X"FC",X"1E",X"1E",
		X"3E",X"3E",X"1F",X"1F",X"0F",X"07",X"01",X"00",X"1E",X"1E",X"DC",X"FC",X"F8",X"F0",X"C0",X"00",
		X"00",X"01",X"07",X"0F",X"1F",X"1F",X"3F",X"3F",X"00",X"C0",X"F0",X"F8",X"FC",X"FC",X"FE",X"FE",
		X"3C",X"3E",X"1E",X"1E",X"0F",X"07",X"01",X"00",X"1E",X"1E",X"1C",X"1C",X"D8",X"F0",X"C0",X"00",
		X"00",X"01",X"07",X"0F",X"1F",X"1F",X"3F",X"3F",X"00",X"C0",X"F0",X"F8",X"FC",X"FC",X"FE",X"FE",
		X"3F",X"3F",X"1C",X"1E",X"0E",X"06",X"01",X"00",X"FE",X"FE",X"1C",X"1C",X"18",X"10",X"C0",X"00",
		X"00",X"00",X"07",X"0F",X"1F",X"1F",X"3F",X"3F",X"00",X"00",X"D0",X"F8",X"FC",X"FC",X"FE",X"FE",
		X"3F",X"3F",X"1F",X"1F",X"0C",X"06",X"00",X"00",X"FE",X"FE",X"FC",X"FC",X"18",X"10",X"00",X"00",
		X"00",X"00",X"06",X"0E",X"1F",X"1F",X"3F",X"3F",X"00",X"00",X"10",X"18",X"DC",X"FC",X"FE",X"FE",
		X"3F",X"3F",X"1F",X"1F",X"0F",X"07",X"00",X"00",X"FE",X"FE",X"FC",X"FC",X"F8",X"F0",X"00",X"00",
		X"00",X"03",X"0F",X"00",X"00",X"00",X"30",X"7D",X"00",X"C0",X"F0",X"F8",X"3C",X"1C",X"0E",X"8E",
		X"7E",X"7F",X"3F",X"3F",X"1F",X"0F",X"03",X"00",X"86",X"06",X"84",X"84",X"C0",X"C0",X"80",X"00",
		X"00",X"03",X"0F",X"00",X"00",X"00",X"31",X"78",X"00",X"C0",X"F0",X"F8",X"3C",X"1C",X"0E",X"8E",
		X"7C",X"7E",X"3F",X"3F",X"1F",X"0F",X"03",X"00",X"46",X"06",X"84",X"84",X"C0",X"C0",X"80",X"00",
		X"00",X"03",X"0F",X"00",X"00",X"00",X"33",X"7C",X"00",X"C0",X"F0",X"F8",X"3C",X"1C",X"8E",X"4E",
		X"7C",X"7C",X"3F",X"3F",X"1F",X"0F",X"03",X"00",X"46",X"46",X"84",X"84",X"C0",X"C0",X"80",X"00",
		X"00",X"03",X"0F",X"00",X"00",X"02",X"30",X"78",X"00",X"C0",X"F0",X"F8",X"3C",X"9C",X"4E",X"2E",
		X"78",X"78",X"3C",X"3F",X"1F",X"0F",X"03",X"00",X"06",X"26",X"04",X"84",X"C0",X"C0",X"80",X"00",
		X"00",X"01",X"03",X"01",X"01",X"01",X"31",X"39",X"C0",X"C0",X"C0",X"C0",X"C0",X"00",X"00",X"00",
		X"39",X"3B",X"1F",X"1F",X"0B",X"03",X"01",X"00",X"00",X"00",X"00",X"C0",X"D0",X"F0",X"E0",X"C0",
		X"00",X"01",X"03",X"01",X"01",X"01",X"31",X"39",X"C0",X"C0",X"D0",X"F0",X"E0",X"00",X"00",X"00",
		X"3B",X"3F",X"1F",X"1B",X"0B",X"03",X"01",X"00",X"00",X"00",X"00",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"00",X"01",X"03",X"01",X"01",X"01",X"31",X"39",X"C0",X"C0",X"C0",X"C0",X"C0",X"00",X"00",X"10",
		X"3D",X"3F",X"1B",X"1B",X"0B",X"03",X"01",X"00",X"30",X"20",X"00",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"00",X"01",X"03",X"01",X"01",X"01",X"31",X"39",X"C0",X"C0",X"C0",X"C0",X"C0",X"00",X"00",X"00",
		X"3D",X"3B",X"1B",X"1B",X"0B",X"07",X"01",X"00",X"00",X"00",X"00",X"C0",X"D0",X"F0",X"E0",X"C0",
		X"00",X"01",X"03",X"03",X"03",X"01",X"31",X"39",X"C0",X"C0",X"D0",X"F0",X"E0",X"00",X"00",X"00",
		X"39",X"39",X"1B",X"1B",X"0F",X"07",X"01",X"00",X"00",X"00",X"00",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"00",X"01",X"03",X"0B",X"01",X"01",X"31",X"39",X"C0",X"C0",X"C0",X"C0",X"C0",X"00",X"00",X"10",
		X"39",X"3B",X"1B",X"1F",X"0F",X"03",X"01",X"00",X"30",X"20",X"00",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"07",X"04",X"00",X"31",X"32",X"7C",X"00",X"C0",X"C0",X"E0",X"30",X"9C",X"4E",X"2E",
		X"7C",X"7E",X"0F",X"0F",X"07",X"07",X"03",X"00",X"26",X"46",X"8C",X"80",X"E0",X"E0",X"80",X"00",
		X"00",X"03",X"01",X"01",X"12",X"0C",X"70",X"3C",X"00",X"C0",X"F0",X"F0",X"38",X"7C",X"9E",X"0E",
		X"3F",X"7F",X"3B",X"31",X"01",X"01",X"03",X"00",X"06",X"96",X"E4",X"80",X"C0",X"C0",X"80",X"00",
		X"00",X"00",X"08",X"08",X"04",X"23",X"10",X"0C",X"00",X"C0",X"70",X"78",X"3C",X"1C",X"26",X"42",
		X"07",X"1F",X"3F",X"3C",X"18",X"08",X"00",X"00",X"42",X"22",X"9C",X"84",X"40",X"40",X"80",X"00",
		X"00",X"03",X"0E",X"02",X"01",X"30",X"08",X"04",X"00",X"00",X"10",X"18",X"3C",X"DC",X"08",X"10",
		X"07",X"0F",X"3F",X"3F",X"1E",X"0E",X"03",X"00",X"10",X"08",X"44",X"24",X"10",X"10",X"00",X"00",
		X"00",X"03",X"0F",X"00",X"00",X"06",X"39",X"60",X"00",X"C0",X"00",X"88",X"4C",X"3C",X"0C",X"88",
		X"70",X"79",X"3F",X"1F",X"0F",X"0F",X"03",X"00",X"80",X"04",X"B4",X"CC",X"80",X"80",X"C0",X"00",
		X"00",X"03",X"00",X"00",X"18",X"03",X"34",X"7C",X"00",X"C0",X"E0",X"E0",X"20",X"90",X"4E",X"2E",
		X"7C",X"6E",X"07",X"03",X"03",X"03",X"03",X"00",X"22",X"50",X"90",X"A0",X"E0",X"E0",X"80",X"00",
		X"00",X"00",X"00",X"10",X"0C",X"01",X"30",X"7C",X"00",X"C0",X"F0",X"98",X"8C",X"04",X"86",X"8E",
		X"7F",X"47",X"03",X"01",X"01",X"03",X"03",X"00",X"70",X"00",X"90",X"A0",X"E0",X"D0",X"80",X"00",
		X"00",X"03",X"03",X"00",X"00",X"38",X"30",X"7C",X"00",X"C0",X"C0",X"80",X"80",X"40",X"26",X"1E",
		X"73",X"61",X"00",X"00",X"01",X"07",X"03",X"00",X"02",X"08",X"90",X"A0",X"E0",X"E0",X"80",X"00",
		X"00",X"03",X"03",X"00",X"00",X"00",X"70",X"7F",X"00",X"C0",X"C0",X"C0",X"20",X"10",X"0E",X"0E",
		X"70",X"70",X"30",X"18",X"0F",X"07",X"03",X"00",X"86",X"4E",X"54",X"A0",X"C0",X"C0",X"80",X"00",
		X"03",X"07",X"07",X"07",X"03",X"07",X"07",X"07",X"E0",X"E0",X"E0",X"C0",X"E0",X"E0",X"E0",X"C0",
		X"00",X"03",X"07",X"04",X"00",X"00",X"00",X"00",X"20",X"E0",X"E0",X"40",X"00",X"00",X"00",X"00",
		X"03",X"07",X"07",X"07",X"03",X"07",X"07",X"07",X"E0",X"E0",X"E0",X"C0",X"E0",X"E0",X"E0",X"C0",
		X"03",X"07",X"07",X"05",X"00",X"00",X"00",X"00",X"A0",X"E0",X"E0",X"C0",X"00",X"00",X"00",X"00",
		X"03",X"07",X"07",X"07",X"03",X"07",X"07",X"07",X"E0",X"E0",X"E0",X"C0",X"E0",X"E0",X"E0",X"C0",
		X"03",X"07",X"07",X"05",X"00",X"00",X"00",X"00",X"E0",X"E0",X"E0",X"40",X"00",X"00",X"00",X"00",
		X"03",X"07",X"07",X"07",X"03",X"07",X"07",X"07",X"E0",X"E0",X"E0",X"C0",X"E0",X"E0",X"E0",X"C0",
		X"02",X"07",X"07",X"07",X"00",X"00",X"00",X"00",X"E0",X"E0",X"E0",X"40",X"00",X"00",X"00",X"00",
		X"03",X"07",X"07",X"07",X"03",X"07",X"07",X"07",X"E0",X"E0",X"E0",X"C0",X"E0",X"E0",X"E0",X"C0",
		X"02",X"07",X"07",X"07",X"00",X"00",X"00",X"00",X"E0",X"E0",X"E0",X"40",X"00",X"00",X"00",X"00",
		X"03",X"07",X"07",X"07",X"03",X"07",X"07",X"07",X"E0",X"E0",X"E0",X"C0",X"E0",X"E0",X"E0",X"C0",
		X"03",X"07",X"07",X"07",X"00",X"03",X"07",X"04",X"E0",X"E0",X"E0",X"C0",X"20",X"E0",X"E0",X"40",
		X"03",X"07",X"07",X"07",X"03",X"07",X"07",X"07",X"E0",X"E0",X"E0",X"C0",X"E0",X"E0",X"E0",X"C0",
		X"03",X"07",X"07",X"07",X"00",X"00",X"00",X"00",X"E0",X"E0",X"E0",X"C0",X"00",X"00",X"00",X"00",
		X"03",X"07",X"07",X"07",X"03",X"07",X"07",X"07",X"E0",X"E0",X"E0",X"C0",X"E0",X"E0",X"E0",X"C0",
		X"03",X"07",X"07",X"07",X"00",X"03",X"07",X"04",X"E0",X"E0",X"E0",X"C0",X"20",X"E0",X"E0",X"40",
		X"03",X"07",X"07",X"07",X"03",X"07",X"07",X"07",X"E0",X"E0",X"E0",X"C0",X"E0",X"E0",X"E0",X"C0",
		X"03",X"07",X"07",X"05",X"00",X"03",X"07",X"04",X"A0",X"E0",X"E0",X"C0",X"20",X"E0",X"E0",X"40",
		X"03",X"07",X"07",X"07",X"03",X"07",X"07",X"07",X"E0",X"E0",X"E0",X"C0",X"E0",X"E0",X"E0",X"C0",
		X"03",X"07",X"07",X"07",X"03",X"07",X"07",X"05",X"E0",X"E0",X"E0",X"C0",X"E0",X"E0",X"E0",X"40",
		X"03",X"07",X"07",X"07",X"03",X"07",X"07",X"07",X"E0",X"E0",X"E0",X"C0",X"E0",X"E0",X"E0",X"C0",
		X"03",X"07",X"07",X"07",X"03",X"07",X"07",X"05",X"E0",X"E0",X"E0",X"C0",X"A0",X"E0",X"E0",X"C0",
		X"03",X"07",X"07",X"07",X"03",X"07",X"07",X"07",X"E0",X"E0",X"E0",X"C0",X"E0",X"E0",X"E0",X"C0",
		X"03",X"07",X"07",X"07",X"03",X"07",X"07",X"07",X"E0",X"E0",X"E0",X"C0",X"E0",X"E0",X"E0",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"07",X"07",X"05",X"00",X"01",X"00",X"01",X"A0",X"E0",X"E0",X"C0",X"A0",X"40",X"A0",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"07",X"07",X"05",X"00",X"01",X"00",X"01",X"E0",X"E0",X"E0",X"40",X"A0",X"40",X"A0",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"03",X"03",X"07",X"00",X"01",X"00",X"01",X"E0",X"C0",X"C0",X"80",X"A0",X"40",X"A0",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"07",X"07",X"07",X"00",X"01",X"00",X"01",X"E0",X"E0",X"E0",X"40",X"A0",X"40",X"A0",X"40",
		X"00",X"00",X"00",X"00",X"08",X"04",X"02",X"01",X"00",X"00",X"00",X"10",X"11",X"11",X"01",X"01",
		X"00",X"00",X"00",X"1C",X"00",X"00",X"00",X"0F",X"08",X"08",X"25",X"11",X"C9",X"20",X"03",X"3B",
		X"00",X"00",X"00",X"08",X"88",X"88",X"80",X"80",X"00",X"00",X"00",X"00",X"10",X"20",X"40",X"80",
		X"10",X"10",X"A4",X"88",X"93",X"04",X"C0",X"DC",X"00",X"00",X"00",X"38",X"00",X"00",X"00",X"F0",
		X"0F",X"00",X"00",X"00",X"1C",X"00",X"00",X"00",X"3B",X"03",X"20",X"C9",X"11",X"25",X"08",X"08",
		X"01",X"02",X"04",X"08",X"00",X"00",X"00",X"00",X"01",X"01",X"11",X"11",X"10",X"00",X"00",X"00",
		X"DC",X"C0",X"04",X"93",X"88",X"A4",X"10",X"10",X"F0",X"00",X"00",X"00",X"38",X"00",X"00",X"00",
		X"80",X"80",X"88",X"88",X"08",X"00",X"00",X"00",X"80",X"40",X"20",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"20",X"10",X"08",X"04",X"00",X"00",X"00",X"01",X"21",X"21",X"20",X"01",X"01",X"11",
		X"00",X"00",X"1C",X"01",X"00",X"00",X"00",X"73",X"90",X"48",X"20",X"80",X"40",X"00",X"00",X"80",
		X"00",X"80",X"80",X"84",X"04",X"04",X"80",X"88",X"00",X"00",X"04",X"08",X"10",X"20",X"00",X"00",
		X"89",X"12",X"04",X"01",X"02",X"00",X"00",X"00",X"00",X"00",X"1C",X"80",X"00",X"00",X"00",X"EE",
		X"77",X"00",X"00",X"00",X"01",X"38",X"00",X"00",X"00",X"00",X"00",X"40",X"80",X"20",X"48",X"91",
		X"00",X"00",X"04",X"08",X"10",X"20",X"00",X"00",X"11",X"01",X"20",X"20",X"21",X"01",X"01",X"00",
		X"01",X"00",X"00",X"02",X"01",X"04",X"12",X"09",X"CE",X"00",X"00",X"00",X"80",X"38",X"00",X"00",
		X"88",X"80",X"80",X"04",X"84",X"84",X"80",X"00",X"00",X"00",X"20",X"10",X"08",X"04",X"00",X"00",
		X"00",X"40",X"20",X"10",X"00",X"00",X"02",X"01",X"81",X"81",X"01",X"00",X"21",X"21",X"00",X"00",
		X"60",X"00",X"0C",X"00",X"00",X"00",X"00",X"EC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"81",X"81",X"00",X"84",X"84",X"00",X"00",X"00",X"02",X"04",X"08",X"00",X"00",X"40",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"30",X"00",X"00",X"00",X"00",X"37",
		X"EC",X"00",X"00",X"00",X"00",X"0C",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"02",X"00",X"00",X"10",X"20",X"40",X"00",X"00",X"00",X"21",X"21",X"00",X"81",X"81",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"37",X"00",X"00",X"00",X"00",X"30",X"00",X"06",
		X"00",X"00",X"84",X"84",X"00",X"80",X"81",X"81",X"80",X"40",X"00",X"00",X"08",X"04",X"02",X"00",
		X"00",X"40",X"20",X"10",X"00",X"00",X"00",X"00",X"81",X"81",X"01",X"00",X"00",X"00",X"00",X"00",
		X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"81",X"81",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"04",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"07",
		X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"20",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"81",X"81",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"06",
		X"00",X"00",X"00",X"00",X"00",X"80",X"81",X"81",X"00",X"00",X"00",X"00",X"08",X"04",X"02",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"7C",X"7E",X"64",X"04",X"05",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"07",X"0E",X"7E",X"E3",X"63",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"04",X"64",X"7E",X"7B",X"30",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"63",X"E3",X"7E",X"0E",X"07",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"4E",X"47",X"02",X"62",X"72",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"07",X"0E",X"7E",X"E3",X"E3",X"F7",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"72",X"62",X"42",X"07",X"4E",X"60",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E3",X"E3",X"7E",X"0E",X"07",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"71",X"73",X"27",X"1F",X"B9",X"B9",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"B9",X"B9",X"1F",X"27",X"73",X"71",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"71",X"E3",X"C7",X"9F",X"B9",X"B9",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"B9",X"B9",X"9F",X"C7",X"E3",X"71",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"FB",X"FA",X"F2",X"F6",X"F4",X"F4",X"E4",X"E8",
		X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"E8",X"E0",X"E0",X"E0",X"E0",X"E0",X"C0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"3F",X"3F",X"3F",X"1F",X"4F",X"07",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"83",X"F0",X"FE",X"FF",X"FF",X"FF",X"7F",X"7F",
		X"9F",X"9F",X"9F",X"9F",X"9F",X"9E",X"9E",X"9E",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",
		X"9C",X"9C",X"88",X"C0",X"40",X"60",X"38",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"02",X"02",X"02",X"03",X"07",X"07",X"03",X"00",X"7F",X"0F",X"01",X"1C",X"1F",X"1F",X"7F",X"7F",
		X"0F",X"0F",X"0F",X"0F",X"1F",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"C0",X"9C",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"86",X"80",X"00",X"C0",X"C0",X"C0",X"80",X"80",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"07",X"07",X"07",X"87",X"87",X"87",X"C3",X"C3",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C3",X"E3",X"E3",X"E1",X"E1",X"E1",X"F1",X"F1",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"80",X"80",X"80",X"00",X"80",X"F0",X"FE",X"FF",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"C3",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"FF",
		X"F1",X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"78",X"08",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",
		X"9C",X"98",X"90",X"80",X"80",X"80",X"80",X"80",X"03",X"02",X"00",X"00",X"08",X"08",X"1F",X"1F",
		X"80",X"80",X"80",X"80",X"83",X"80",X"89",X"8C",X"0F",X"45",X"01",X"40",X"40",X"50",X"FC",X"78",
		X"03",X"07",X"07",X"0F",X"0F",X"1F",X"0F",X"E1",X"F8",X"F0",X"F0",X"E0",X"E0",X"E0",X"C0",X"C0",
		X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"04",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"BC",X"B8",X"0C",X"EE",X"E8",X"E4",X"E5",X"F7",
		X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"F7",X"FF",X"FF",X"FE",X"FE",X"FC",X"FD",X"F9",
		X"0C",X"1C",X"38",X"98",X"C8",X"60",X"30",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"80",X"00",X"40",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"17",X"17",
		X"3E",X"20",X"00",X"30",X"7E",X"7E",X"7C",X"00",X"00",X"30",X"00",X"00",X"00",X"08",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"7F",X"7F",X"0F",X"0F",X"0F",X"8F",X"8F",X"E0",X"F0",X"F0",X"F8",X"F8",X"F8",X"FC",X"FC",
		X"8F",X"8F",X"8F",X"0F",X"0F",X"0F",X"0F",X"0F",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",X"E0",X"00",X"00",X"00",X"00",X"00",X"04",X"0E",X"0E",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"41",X"49",X"49",X"49",X"7F",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"7F",X"38",X"1C",X"38",X"7F",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"39",X"7B",X"4F",X"46",X"44",X"7F",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"41",X"49",X"49",X"49",X"7F",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"3F",X"64",X"44",X"64",X"3F",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"4F",X"4F",X"49",X"49",X"63",X"3E",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"78",X"7C",X"0E",X"07",X"0E",X"7C",X"78",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3E",X"7F",X"41",X"41",X"41",X"7F",X"3E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"03",X"07",X"0E",X"1C",X"38",X"71",X"E3",X"FF",X"FF",X"00",X"00",X"7F",X"FF",X"C0",X"80",
		X"C7",X"CE",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"FE",X"FF",X"03",X"01",X"80",X"C0",X"E0",X"70",X"38",X"1C",X"8E",X"C7",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E3",X"73",X"33",X"33",X"33",X"33",X"33",X"33",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CE",X"C7",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E3",X"71",X"38",X"1C",X"0E",X"07",X"03",X"01",X"80",X"C0",X"FF",X"7F",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"33",X"33",X"33",X"33",X"33",X"73",X"E3",
		X"01",X"03",X"FF",X"FE",X"00",X"00",X"FF",X"FF",X"C7",X"8E",X"1C",X"38",X"70",X"E0",X"C0",X"80",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"F0",X"F0",X"F1",X"F7",X"F7",X"F3",X"FB",X"F8",
		X"9F",X"9F",X"9E",X"98",X"80",X"80",X"80",X"80",X"F0",X"C0",X"00",X"00",X"02",X"0B",X"3B",X"7B",
		X"04",X"3C",X"FC",X"FC",X"F8",X"E0",X"80",X"00",X"80",X"F0",X"C1",X"07",X"1E",X"3C",X"78",X"11",
		X"06",X"0E",X"06",X"00",X"00",X"F8",X"E0",X"C1",X"03",X"38",X"70",X"00",X"00",X"00",X"F8",X"F8",
		X"81",X"83",X"8F",X"9F",X"9F",X"9F",X"9F",X"9F",X"FB",X"FB",X"F8",X"F8",X"F8",X"FC",X"FF",X"FE",
		X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9E",X"FC",X"F8",X"F0",X"E0",X"C0",X"80",X"03",X"03",
		X"83",X"07",X"0F",X"1F",X"3F",X"7F",X"1F",X"06",X"F0",X"F0",X"E1",X"C3",X"83",X"07",X"0E",X"0F",
		X"00",X"04",X"00",X"00",X"00",X"00",X"81",X"03",X"1F",X"3E",X"3E",X"06",X"3C",X"FC",X"F8",X"F8",
		X"00",X"00",X"80",X"98",X"3F",X"7A",X"F6",X"F6",X"A8",X"28",X"28",X"28",X"68",X"68",X"4C",X"4C",
		X"EC",X"4C",X"08",X"00",X"00",X"00",X"00",X"60",X"CC",X"CC",X"CC",X"CC",X"0C",X"04",X"00",X"00",
		X"4F",X"67",X"73",X"39",X"3C",X"3E",X"3F",X"3F",X"C0",X"F0",X"FC",X"FF",X"7F",X"3F",X"18",X"80",
		X"1F",X"1F",X"2F",X"27",X"27",X"F3",X"31",X"39",X"C0",X"0E",X"0F",X"07",X"43",X"41",X"60",X"70",
		X"E3",X"E3",X"C3",X"C3",X"87",X"87",X"07",X"07",X"80",X"8E",X"8E",X"8E",X"8E",X"8F",X"0F",X"0F",
		X"00",X"08",X"0E",X"0F",X"1F",X"1F",X"1E",X"1E",X"0F",X"00",X"00",X"00",X"00",X"08",X"0E",X"0F",
		X"38",X"38",X"1C",X"1C",X"1E",X"1E",X"1E",X"1F",X"78",X"7C",X"7C",X"3E",X"1F",X"1F",X"00",X"07",
		X"7F",X"7F",X"FF",X"3F",X"0F",X"0F",X"0F",X"BF",X"07",X"83",X"81",X"81",X"C0",X"C0",X"E0",X"E0",
		X"9E",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"01",X"00",X"C0",X"E0",X"F8",X"FC",X"FF",X"FF",
		X"9F",X"9F",X"9F",X"9F",X"87",X"81",X"80",X"80",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"0F",
		X"FF",X"FF",X"7F",X"3F",X"1F",X"0F",X"07",X"83",X"F0",X"F0",X"F8",X"FC",X"FC",X"FE",X"FF",X"FF",
		X"C1",X"E0",X"F8",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"1F",X"8F",X"C7",X"E3",
		X"80",X"80",X"9C",X"9F",X"9F",X"9F",X"9F",X"9F",X"03",X"00",X"00",X"80",X"F0",X"FC",X"FD",X"F9",
		X"9F",X"9F",X"9F",X"9F",X"80",X"80",X"80",X"80",X"FB",X"F8",X"F0",X"F0",X"07",X"07",X"07",X"30",
		X"F0",X"40",X"00",X"04",X"00",X"00",X"C0",X"F8",X"71",X"1C",X"06",X"02",X"00",X"00",X"03",X"01",
		X"FF",X"3F",X"00",X"00",X"FC",X"FC",X"C0",X"00",X"80",X"F8",X"1F",X"00",X"1F",X"00",X"07",X"06",
		X"FF",X"7F",X"7F",X"3F",X"3F",X"3F",X"1F",X"1E",X"10",X"11",X"91",X"91",X"91",X"81",X"81",X"00",
		X"1E",X"8E",X"8E",X"C6",X"C6",X"E6",X"F2",X"F2",X"60",X"70",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"C0",X"E0",X"C0",X"C0",X"C3",X"47",X"F0",X"70",X"F0",X"1E",X"10",X"03",X"01",X"00",
		X"06",X"06",X"00",X"1C",X"07",X"00",X"00",X"00",X"10",X"3C",X"7E",X"7C",X"18",X"01",X"11",X"00",
		X"00",X"00",X"00",X"04",X"62",X"32",X"88",X"E4",X"B2",X"B2",X"96",X"96",X"D4",X"55",X"55",X"54",
		X"7A",X"1C",X"C2",X"00",X"FF",X"02",X"30",X"01",X"55",X"55",X"38",X"17",X"C0",X"21",X"98",X"48",
		X"60",X"EF",X"DE",X"BC",X"F9",X"73",X"E6",X"CC",X"00",X"00",X"20",X"78",X"E0",X"81",X"1F",X"F8",
		X"9B",X"40",X"80",X"C1",X"07",X"C3",X"58",X"1E",X"80",X"03",X"7F",X"07",X"F0",X"FC",X"0E",X"00",
		X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"00",X"00",X"80",X"C0",X"C0",X"E0",X"F0",X"F0",
		X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"F8",X"FC",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",
		X"1F",X"0F",X"0F",X"07",X"07",X"07",X"03",X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"01",X"01",X"01",X"00",X"00",X"00",X"80",X"C0",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",
		X"9F",X"9F",X"9F",X"9F",X"9F",X"8F",X"87",X"83",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"81",X"80",X"80",X"80",X"80",X"80",X"98",X"9C",X"FF",X"FF",X"7F",X"3F",X"1F",X"0F",X"07",X"03",
		X"C0",X"E0",X"E0",X"F0",X"F0",X"F8",X"F8",X"FC",X"3F",X"3F",X"1F",X"1F",X"1F",X"0F",X"0F",X"07",
		X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"07",X"07",X"03",X"03",X"81",X"C1",X"C1",X"E0",
		X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"70",X"70",X"70",X"60",X"00",X"10",X"30",X"70",
		X"F8",X"F8",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"70",X"70",X"70",X"30",X"30",X"10",X"10",X"00",
		X"0F",X"0F",X"1F",X"1F",X"1F",X"03",X"00",X"00",X"E0",X"E0",X"E0",X"E0",X"C0",X"C0",X"00",X"C0",
		X"01",X"13",X"07",X"07",X"01",X"00",X"00",X"30",X"80",X"80",X"80",X"80",X"00",X"00",X"01",X"00",
		X"FC",X"FC",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"00",X"00",X"00",X"08",X"0C",X"0E",X"00",X"00",
		X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"3E",X"3E",X"7E",X"7E",X"7C",X"7C",X"1C",X"04",X"00",X"00",X"07",X"07",X"07",X"0F",X"0F",X"1F",
		X"00",X"78",X"D8",X"C8",X"C0",X"E0",X"F0",X"F0",X"1F",X"1F",X"00",X"3F",X"5E",X"0C",X"28",X"E0",
		X"0F",X"38",X"60",X"40",X"C0",X"80",X"80",X"80",X"FF",X"00",X"00",X"FF",X"FF",X"7F",X"7F",X"7F",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"3F",X"3F",X"1F",X"1F",X"1F",X"0F",X"0F",X"07",
		X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"07",X"07",X"03",X"03",X"01",X"01",X"01",X"00",
		X"90",X"90",X"98",X"98",X"9C",X"9C",X"9E",X"9E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"7F",X"7F",X"7F",X"3F",X"3F",X"1F",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"FF",X"00",X"00",X"0F",X"0F",X"07",X"03",X"01",
		X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"40",X"60",X"70",X"70",X"70",X"70",X"70",X"70",
		X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"7F",X"3F",X"1F",X"0F",X"07",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"C0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"70",X"70",X"10",X"00",X"00",X"00",X"08",X"02",
		X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"60",X"70",X"70",X"70",X"70",X"70",
		X"00",X"00",X"00",X"04",X"06",X"07",X"07",X"07",X"7E",X"3E",X"0E",X"04",X"00",X"80",X"C4",X"EC",
		X"07",X"07",X"07",X"01",X"00",X"0F",X"0F",X"0F",X"F8",X"F8",X"F8",X"F8",X"70",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"60",X"30",X"1C",X"0E",X"07",X"00",X"00",X"20",X"20",X"10",X"10",X"18",X"0C",
		X"03",X"03",X"01",X"00",X"00",X"0F",X"03",X"00",X"8E",X"CF",X"E7",X"F7",X"7F",X"3F",X"FF",X"FF",
		X"00",X"00",X"01",X"02",X"02",X"04",X"0C",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"38",X"78",X"F9",X"FF",X"FF",X"FF",X"FF",X"FE",X"00",X"0F",X"FC",X"F0",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"1E",X"3F",X"1F",X"3F",X"7F",X"FF",X"FF",X"C7",X"07",
		X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"04",X"0C",X"08",X"08",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"7F",X"77",X"80",X"E0",X"F8",X"FC",X"00",X"00",X"00",X"80",
		X"33",X"31",X"30",X"10",X"10",X"10",X"00",X"00",X"C0",X"C0",X"E0",X"60",X"30",X"18",X"08",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"42",X"00",X"40",X"00",
		X"00",X"00",X"09",X"00",X"00",X"02",X"00",X"24",X"00",X"04",X"00",X"00",X"20",X"02",X"00",X"88",
		X"00",X"00",X"00",X"40",X"00",X"00",X"02",X"90",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",
		X"00",X"00",X"10",X"82",X"00",X"00",X"50",X"00",X"00",X"20",X"00",X"00",X"88",X"00",X"00",X"02",
		X"00",X"10",X"00",X"01",X"00",X"10",X"02",X"00",X"02",X"00",X"10",X"00",X"40",X"01",X"00",X"00",
		X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"81",X"08",X"00",X"40",X"08",X"00",X"01",X"00",
		X"04",X"01",X"40",X"00",X"00",X"08",X"00",X"00",X"10",X"00",X"00",X"08",X"00",X"40",X"00",X"00",
		X"10",X"00",X"04",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"10",X"00",X"00",X"00",X"00",
		X"04",X"00",X"11",X"00",X"08",X"00",X"00",X"40",X"01",X"10",X"00",X"00",X"24",X"00",X"00",X"82",
		X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",
		X"00",X"10",X"01",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"12",X"00",X"00",
		X"00",X"08",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"40",X"00",X"00",X"04",X"20",X"00",X"00",
		X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"20",X"00",X"01",X"00",X"00",
		X"00",X"81",X"00",X"10",X"00",X"00",X"80",X"00",X"10",X"00",X"00",X"00",X"90",X"00",X"00",X"10",
		X"01",X"10",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
