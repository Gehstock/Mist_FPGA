library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity e1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of e1 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"18",X"C3",X"95",X"17",X"E5",X"7D",X"C6",X"0E",X"6F",X"7E",X"B7",X"C2",X"36",X"18",X"E1",X"7E",
		X"B8",X"DC",X"40",X"18",X"7E",X"B9",X"D8",X"06",X"00",X"70",X"2B",X"70",X"7D",X"C6",X"0E",X"6F",
		X"70",X"2B",X"2B",X"2B",X"46",X"2B",X"4E",X"7D",X"D6",X"0C",X"6F",X"CD",X"11",X"15",X"1E",X"08",
		X"CD",X"42",X"15",X"C1",X"C1",X"C9",X"7D",X"C6",X"05",X"6F",X"EF",X"E1",X"C0",X"C3",X"17",X"18",
		X"1A",X"FE",X"80",X"D8",X"2F",X"C6",X"05",X"12",X"1B",X"1B",X"1B",X"1A",X"D6",X"02",X"12",X"13",
		X"13",X"13",X"C9",X"3A",X"66",X"20",X"B7",X"CA",X"5F",X"18",X"CD",X"63",X"18",X"2B",X"2B",X"CD",
		X"63",X"18",X"C9",X"7E",X"23",X"35",X"23",X"C0",X"2B",X"77",X"23",X"1A",X"86",X"12",X"C9",X"3A",
		X"CF",X"22",X"B7",X"CA",X"64",X"19",X"21",X"C4",X"22",X"11",X"C2",X"22",X"CD",X"53",X"18",X"23",
		X"13",X"CD",X"53",X"18",X"2A",X"CC",X"22",X"44",X"4D",X"2A",X"CA",X"22",X"1A",X"BC",X"DA",X"38",
		X"19",X"BD",X"D2",X"38",X"19",X"21",X"C0",X"22",X"CD",X"F2",X"18",X"C9",X"3A",X"DF",X"22",X"B7",
		X"C8",X"21",X"D4",X"22",X"11",X"D2",X"22",X"CD",X"53",X"18",X"23",X"13",X"CD",X"53",X"18",X"2A",
		X"DC",X"22",X"44",X"4D",X"2A",X"DA",X"22",X"1A",X"BC",X"DA",X"1E",X"19",X"BD",X"D2",X"1E",X"19",
		X"21",X"D0",X"22",X"CD",X"F2",X"18",X"C9",X"3A",X"EF",X"22",X"B7",X"C8",X"21",X"E4",X"22",X"11",
		X"E2",X"22",X"CD",X"53",X"18",X"23",X"13",X"CD",X"53",X"18",X"2A",X"EC",X"22",X"44",X"4D",X"2A",
		X"EA",X"22",X"1A",X"BC",X"DA",X"1E",X"19",X"BD",X"D2",X"1E",X"19",X"21",X"E0",X"22",X"CD",X"F2",
		X"18",X"C9",X"C5",X"E5",X"CD",X"0E",X"19",X"1E",X"05",X"CD",X"2A",X"15",X"E1",X"C1",X"23",X"23",
		X"E5",X"CD",X"0E",X"19",X"1E",X"05",X"CD",X"B7",X"15",X"E1",X"CD",X"F2",X"15",X"C9",X"7E",X"07",
		X"07",X"07",X"07",X"E6",X"70",X"81",X"D2",X"1A",X"19",X"04",X"4F",X"C3",X"DD",X"14",X"EB",X"2B",
		X"2B",X"2B",X"E5",X"CD",X"0E",X"19",X"1E",X"08",X"CD",X"2A",X"15",X"E1",X"23",X"23",X"CD",X"F2",
		X"15",X"7D",X"C6",X"0F",X"6F",X"36",X"00",X"C9",X"AF",X"32",X"C6",X"22",X"32",X"C9",X"22",X"32",
		X"CF",X"22",X"EB",X"2B",X"2B",X"2B",X"CD",X"0E",X"19",X"1E",X"08",X"CD",X"2A",X"15",X"21",X"88",
		X"43",X"22",X"CC",X"22",X"3E",X"04",X"32",X"F6",X"22",X"2A",X"C0",X"22",X"11",X"FE",X"FF",X"19",
		X"22",X"F7",X"22",X"C9",X"21",X"F6",X"22",X"EF",X"DA",X"73",X"19",X"C8",X"CD",X"80",X"19",X"CD",
		X"B7",X"15",X"C9",X"CD",X"80",X"19",X"CD",X"2A",X"15",X"21",X"00",X"13",X"22",X"CC",X"22",X"C9",
		X"2A",X"CC",X"22",X"44",X"4D",X"21",X"F7",X"22",X"CD",X"8E",X"19",X"1E",X"08",X"C9",X"7E",X"07",
		X"07",X"07",X"E6",X"30",X"81",X"D2",X"99",X"19",X"14",X"4F",X"C3",X"DD",X"14",X"10",X"E0",X"10",
		X"E0",X"10",X"E0",X"5C",X"96",X"50",X"A0",X"46",X"AA",X"3C",X"B4",X"32",X"BE",X"28",X"C8",X"1E",
		X"D2",X"14",X"DC",X"0A",X"E6",X"0A",X"E6",X"0A",X"E6",X"0A",X"E6",X"0A",X"E6",X"3A",X"90",X"22",
		X"B7",X"C8",X"2A",X"8A",X"22",X"44",X"4D",X"21",X"83",X"22",X"11",X"89",X"22",X"CD",X"FE",X"17",
		X"EB",X"2B",X"2B",X"CD",X"53",X"18",X"23",X"13",X"CD",X"53",X"18",X"2A",X"8C",X"22",X"44",X"4D",
		X"21",X"80",X"22",X"CD",X"11",X"1A",X"C9",X"3A",X"B0",X"22",X"B7",X"C8",X"2A",X"AA",X"22",X"44",
		X"4D",X"21",X"A3",X"22",X"11",X"A9",X"22",X"CD",X"FE",X"17",X"EB",X"2B",X"2B",X"CD",X"53",X"18",
		X"23",X"13",X"CD",X"53",X"18",X"2A",X"AC",X"22",X"44",X"4D",X"21",X"A0",X"22",X"CD",X"11",X"1A",
		X"C9",X"C5",X"E5",X"E5",X"7D",X"C6",X"13",X"6F",X"7E",X"B7",X"CA",X"23",X"1A",X"36",X"00",X"23",
		X"4E",X"23",X"46",X"E1",X"CD",X"11",X"15",X"22",X"F1",X"21",X"E1",X"E5",X"1E",X"08",X"CD",X"75",
		X"1A",X"2A",X"F1",X"21",X"CD",X"42",X"15",X"E1",X"C1",X"23",X"23",X"E5",X"CD",X"11",X"15",X"22",
		X"F1",X"21",X"E1",X"E5",X"1E",X"08",X"CD",X"54",X"1A",X"2A",X"F1",X"21",X"CD",X"CD",X"15",X"E1",
		X"CD",X"F2",X"15",X"C9",X"23",X"56",X"7D",X"C6",X"06",X"6F",X"7E",X"FE",X"7F",X"D8",X"7D",X"C6",
		X"0E",X"6F",X"3A",X"0A",X"20",X"77",X"92",X"DA",X"72",X"1A",X"5F",X"1C",X"3E",X"08",X"BB",X"D0",
		X"5F",X"C9",X"1E",X"00",X"C9",X"23",X"56",X"7D",X"C6",X"08",X"6F",X"7E",X"FE",X"7F",X"D8",X"7D",
		X"C6",X"0E",X"6F",X"7E",X"92",X"DA",X"90",X"1A",X"5F",X"1C",X"3E",X"08",X"BB",X"D0",X"5F",X"C9",
		X"1E",X"00",X"C9",X"CD",X"13",X"1B",X"21",X"6A",X"20",X"11",X"6E",X"20",X"3A",X"04",X"20",X"B7",
		X"C2",X"4C",X"1B",X"1A",X"86",X"77",X"3E",X"D0",X"BE",X"DA",X"E5",X"1A",X"3E",X"20",X"BE",X"D2",
		X"E5",X"1A",X"13",X"13",X"13",X"1A",X"23",X"86",X"77",X"3E",X"40",X"BE",X"DA",X"C0",X"1A",X"77",
		X"3E",X"D0",X"BE",X"D0",X"AF",X"32",X"C0",X"21",X"32",X"C3",X"21",X"3E",X"FF",X"32",X"22",X"20",
		X"21",X"7B",X"20",X"BE",X"CA",X"DE",X"1A",X"77",X"2A",X"74",X"20",X"22",X"7C",X"20",X"21",X"80",
		X"11",X"22",X"74",X"20",X"C9",X"77",X"21",X"C2",X"21",X"EF",X"C0",X"1A",X"2F",X"3C",X"12",X"13",
		X"13",X"13",X"3E",X"02",X"12",X"3A",X"C0",X"21",X"2F",X"32",X"C0",X"21",X"AF",X"32",X"D7",X"20",
		X"32",X"62",X"20",X"21",X"90",X"21",X"7E",X"23",X"23",X"B6",X"C2",X"12",X"1B",X"3E",X"FF",X"32",
		X"D9",X"20",X"C9",X"21",X"C1",X"21",X"EF",X"C0",X"36",X"03",X"3E",X"FF",X"21",X"7B",X"20",X"BE",
		X"CA",X"2A",X"1B",X"77",X"2A",X"74",X"20",X"22",X"7C",X"20",X"21",X"C3",X"21",X"34",X"3A",X"C0",
		X"21",X"B7",X"CA",X"37",X"1B",X"35",X"35",X"7E",X"E6",X"03",X"07",X"21",X"80",X"40",X"85",X"D2",
		X"43",X"1B",X"24",X"6F",X"5E",X"23",X"56",X"EB",X"22",X"74",X"20",X"C9",X"1A",X"86",X"77",X"3E",
		X"DF",X"BE",X"DA",X"83",X"1B",X"3E",X"01",X"BE",X"D2",X"83",X"1B",X"13",X"13",X"13",X"1A",X"23",
		X"86",X"77",X"3A",X"C2",X"21",X"B7",X"CA",X"70",X"1B",X"3E",X"40",X"BE",X"DA",X"70",X"1B",X"77",
		X"3E",X"D0",X"BE",X"D0",X"3A",X"89",X"21",X"3D",X"32",X"89",X"21",X"3E",X"FF",X"32",X"D9",X"20",
		X"C3",X"C4",X"1A",X"21",X"FF",X"FF",X"22",X"6A",X"20",X"21",X"A0",X"21",X"7E",X"E6",X"FB",X"77",
		X"21",X"C2",X"21",X"EF",X"C0",X"1A",X"FE",X"80",X"DA",X"9D",X"1B",X"2F",X"3C",X"12",X"13",X"13",
		X"13",X"3E",X"02",X"12",X"3E",X"00",X"32",X"C0",X"21",X"AF",X"32",X"D7",X"20",X"32",X"62",X"20",
		X"CD",X"CE",X"1B",X"3E",X"30",X"32",X"6B",X"20",X"3A",X"89",X"21",X"C6",X"03",X"07",X"07",X"07",
		X"32",X"6A",X"20",X"11",X"00",X"01",X"2A",X"E0",X"21",X"19",X"22",X"E0",X"21",X"C9",X"2A",X"8A",
		X"21",X"2B",X"22",X"8A",X"21",X"23",X"11",X"D0",X"43",X"06",X"08",X"CD",X"0A",X"0E",X"AF",X"32",
		X"F4",X"21",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C3",X"75",X"1C",X"C3",X"C2",X"1C",X"C3",X"12",X"1C",X"C3",X"00",X"5C",X"C3",X"1B",X"1D",X"C3",
		X"24",X"1D",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"FF",X"32",X"4E",X"20",X"21",X"4D",X"20",
		X"7E",X"36",X"FF",X"B7",X"CC",X"12",X"50",X"AF",X"32",X"01",X"20",X"CD",X"C4",X"0C",X"CD",X"22",
		X"14",X"CD",X"55",X"14",X"CD",X"00",X"48",X"CD",X"0A",X"48",X"CD",X"0D",X"48",X"CD",X"77",X"0D",
		X"CD",X"12",X"01",X"CD",X"1A",X"0E",X"CD",X"00",X"44",X"CD",X"07",X"44",X"CD",X"00",X"50",X"CD",
		X"03",X"50",X"CD",X"06",X"50",X"CD",X"09",X"50",X"CD",X"16",X"48",X"CD",X"77",X"1D",X"CD",X"24",
		X"50",X"CD",X"58",X"14",X"CD",X"27",X"50",X"CD",X"48",X"14",X"CD",X"0F",X"14",X"00",X"00",X"00",
		X"00",X"00",X"00",X"E7",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"CD",X"C4",X"0C",X"CD",X"22",
		X"14",X"CD",X"55",X"14",X"CD",X"00",X"48",X"CD",X"0D",X"48",X"CD",X"77",X"0D",X"CD",X"1A",X"0E",
		X"CD",X"07",X"44",X"CD",X"00",X"50",X"CD",X"03",X"50",X"CD",X"06",X"50",X"CD",X"09",X"50",X"CD",
		X"88",X"1D",X"CD",X"58",X"14",X"CD",X"27",X"50",X"CD",X"48",X"14",X"CD",X"0F",X"14",X"CD",X"1A",
		X"5C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CD",X"0C",X"50",
		X"E7",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"CD",X"C4",X"0C",X"CD",X"22",X"14",X"CD",X"55",
		X"14",X"CD",X"00",X"48",X"CD",X"0A",X"48",X"CD",X"0D",X"48",X"CD",X"77",X"0D",X"CD",X"12",X"01",
		X"CD",X"1A",X"0E",X"CD",X"15",X"50",X"CD",X"00",X"44",X"CD",X"07",X"44",X"CD",X"00",X"50",X"CD",
		X"03",X"50",X"CD",X"06",X"50",X"CD",X"09",X"50",X"CD",X"16",X"48",X"CD",X"24",X"50",X"CD",X"58",
		X"14",X"CD",X"27",X"50",X"CD",X"48",X"14",X"CD",X"0F",X"14",X"CD",X"1A",X"5C",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E7",X"C9",X"21",X"02",X"20",X"AF",X"77",
		X"2F",X"23",X"77",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"CD",X"C4",X"0C",X"CD",X"22",X"14",
		X"CD",X"55",X"14",X"CD",X"00",X"48",X"CD",X"0D",X"48",X"CD",X"77",X"0D",X"CD",X"12",X"01",X"CD",
		X"1A",X"0E",X"CD",X"18",X"50",X"CD",X"1B",X"50",X"CD",X"00",X"44",X"CD",X"07",X"44",X"CD",X"00",
		X"50",X"CD",X"03",X"50",X"CD",X"06",X"50",X"CD",X"09",X"50",X"CD",X"16",X"48",X"CD",X"24",X"50",
		X"CD",X"58",X"14",X"CD",X"48",X"14",X"CD",X"0F",X"14",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E7",X"C9",X"21",X"A0",X"21",X"7E",X"E6",X"FB",X"77",X"DB",X"00",
		X"E6",X"80",X"C0",X"7E",X"F6",X"04",X"77",X"C9",X"21",X"5A",X"23",X"3E",X"FF",X"BE",X"C2",X"59",
		X"1E",X"CD",X"DC",X"1F",X"21",X"90",X"21",X"7E",X"23",X"23",X"B6",X"C0",X"CD",X"89",X"5A",X"2A",
		X"5C",X"23",X"CD",X"0F",X"50",X"22",X"5C",X"23",X"CA",X"6B",X"1E",X"CD",X"BE",X"1D",X"CD",X"2F",
		X"1E",X"CD",X"10",X"1E",X"CD",X"4E",X"1E",X"CD",X"64",X"1F",X"CD",X"1C",X"48",X"C9",X"3A",X"12",
		X"20",X"E6",X"1F",X"FE",X"0F",X"C0",X"3A",X"22",X"20",X"B7",X"C8",X"3A",X"12",X"20",X"07",X"07",
		X"07",X"E6",X"06",X"21",X"00",X"1E",X"85",X"D2",X"DB",X"1D",X"24",X"6F",X"5E",X"23",X"56",X"1A",
		X"B7",X"C0",X"7B",X"D6",X"10",X"5F",X"01",X"08",X"1E",X"3A",X"12",X"20",X"07",X"07",X"07",X"E6",
		X"06",X"81",X"D2",X"F6",X"1D",X"04",X"4F",X"0A",X"6F",X"03",X"0A",X"67",X"06",X"20",X"FF",X"C9",
		X"10",X"22",X"30",X"22",X"50",X"22",X"70",X"22",X"74",X"06",X"9C",X"06",X"C4",X"06",X"EC",X"06",
		X"3A",X"12",X"20",X"E6",X"60",X"C0",X"21",X"21",X"20",X"3A",X"12",X"20",X"E6",X"80",X"CA",X"28",
		X"1E",X"3E",X"B0",X"34",X"BE",X"D0",X"77",X"C9",X"3E",X"90",X"35",X"BE",X"D8",X"77",X"C9",X"3A",
		X"12",X"20",X"E6",X"01",X"C0",X"21",X"20",X"20",X"11",X"26",X"20",X"1A",X"86",X"77",X"FE",X"20",
		X"D2",X"47",X"1E",X"3E",X"01",X"12",X"C9",X"FE",X"C0",X"D8",X"3E",X"FF",X"12",X"C9",X"21",X"C5",
		X"21",X"EF",X"C0",X"36",X"FF",X"23",X"36",X"FF",X"C9",X"77",X"3E",X"B0",X"32",X"21",X"20",X"11",
		X"AD",X"59",X"21",X"98",X"28",X"0E",X"05",X"CD",X"EE",X"02",X"C9",X"3E",X"FF",X"32",X"F1",X"22",
		X"32",X"F2",X"22",X"32",X"DE",X"22",X"32",X"EE",X"22",X"CD",X"C3",X"1E",X"CD",X"8C",X"1E",X"CD",
		X"1F",X"1F",X"CD",X"41",X"1F",X"CD",X"64",X"1F",X"CD",X"1C",X"48",X"C9",X"3A",X"5E",X"23",X"B7",
		X"C2",X"9A",X"1E",X"CD",X"2F",X"1E",X"CD",X"10",X"1E",X"C9",X"CD",X"B5",X"1E",X"CD",X"A1",X"1E",
		X"C9",X"3A",X"12",X"20",X"E6",X"01",X"C0",X"21",X"21",X"20",X"3E",X"80",X"BE",X"C8",X"DA",X"B3",
		X"1E",X"34",X"34",X"35",X"C9",X"21",X"20",X"20",X"3E",X"74",X"BE",X"C8",X"DA",X"C1",X"1E",X"34",
		X"34",X"35",X"C9",X"3A",X"F6",X"22",X"21",X"CF",X"22",X"B6",X"C0",X"3A",X"5E",X"23",X"B7",X"C2",
		X"E1",X"1E",X"CD",X"0F",X"1F",X"C8",X"21",X"C5",X"21",X"EF",X"C0",X"36",X"1E",X"23",X"36",X"FF",
		X"C9",X"3A",X"E3",X"21",X"FE",X"03",X"D2",X"02",X"1F",X"3E",X"FF",X"32",X"60",X"23",X"3A",X"B1",
		X"22",X"B7",X"C0",X"3A",X"A2",X"22",X"FE",X"8C",X"D0",X"FE",X"60",X"D8",X"21",X"C6",X"21",X"36",
		X"FF",X"C9",X"21",X"60",X"23",X"EF",X"C0",X"36",X"FF",X"21",X"C6",X"21",X"36",X"FF",X"C9",X"3A",
		X"10",X"22",X"21",X"30",X"22",X"B6",X"21",X"50",X"22",X"B6",X"21",X"70",X"22",X"B6",X"C9",X"3A",
		X"5E",X"23",X"B7",X"C0",X"21",X"FF",X"FF",X"22",X"E0",X"21",X"AF",X"32",X"E3",X"21",X"CD",X"0F",
		X"1F",X"C0",X"21",X"01",X"00",X"22",X"E0",X"21",X"21",X"5E",X"23",X"36",X"FF",X"23",X"36",X"10",
		X"C9",X"21",X"5F",X"23",X"EF",X"C0",X"2B",X"7E",X"B7",X"C8",X"3A",X"E2",X"21",X"B7",X"C0",X"AF",
		X"77",X"32",X"F1",X"22",X"32",X"F2",X"22",X"32",X"DE",X"22",X"32",X"EE",X"22",X"21",X"00",X"06",
		X"22",X"5C",X"23",X"C9",X"2A",X"80",X"21",X"7D",X"B4",X"C0",X"2A",X"61",X"23",X"CD",X"0F",X"50",
		X"22",X"61",X"23",X"C0",X"CD",X"9E",X"1F",X"21",X"63",X"23",X"34",X"7E",X"E6",X"01",X"CA",X"B5",
		X"1F",X"21",X"80",X"00",X"22",X"61",X"23",X"11",X"60",X"59",X"21",X"2C",X"28",X"0E",X"0B",X"CD",
		X"D9",X"02",X"11",X"8C",X"59",X"21",X"30",X"28",X"0E",X"0B",X"CD",X"EE",X"02",X"C9",X"21",X"28",
		X"28",X"11",X"13",X"00",X"0E",X"0B",X"06",X"0D",X"AF",X"77",X"23",X"05",X"C2",X"A8",X"1F",X"19",
		X"0D",X"C2",X"A6",X"1F",X"C9",X"21",X"00",X"04",X"22",X"61",X"23",X"21",X"C8",X"1F",X"22",X"80",
		X"21",X"21",X"42",X"28",X"22",X"82",X"21",X"C9",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"49",X"4E",X"53",X"45",X"52",X"54",X"20",X"43",X"4F",X"49",X"4E",X"FF",X"11",X"BC",X"59",X"21",
		X"3B",X"28",X"0E",X"0B",X"CD",X"EE",X"02",X"3A",X"41",X"20",X"07",X"07",X"07",X"21",X"7C",X"28",
		X"CD",X"31",X"0F",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
