library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity kick_bg_bits_1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of kick_bg_bits_1 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"55",X"55",X"55",X"AA",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"AA",X"AA",X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"FF",X"FF",
		X"AA",X"A0",X"AA",X"A8",X"AA",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"0F",X"55",X"0F",X"55",X"4F",X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"55",X"55",X"55",X"55",X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"FF",X"FF",
		X"00",X"AA",X"00",X"2A",X"00",X"0A",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",
		X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"00",
		X"C2",X"AB",X"C2",X"AB",X"C2",X"AB",X"C2",X"AB",X"C2",X"AB",X"C2",X"AB",X"C2",X"AB",X"C2",X"AB",
		X"C0",X"03",X"C2",X"AB",X"C2",X"AB",X"C2",X"AB",X"C2",X"AB",X"C2",X"AB",X"C2",X"AB",X"C2",X"AB",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"AA",X"AA",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"CA",X"A8",X"CA",X"A8",X"CA",X"A8",X"CA",X"A8",X"CA",X"A8",X"80",X"00",X"FF",X"FF",X"FF",X"FF",
		X"CA",X"A8",X"CA",X"A8",X"CA",X"A8",X"CA",X"A8",X"CA",X"A8",X"CA",X"A8",X"CA",X"A8",X"80",X"00",
		X"00",X"00",X"00",X"00",X"AA",X"A8",X"AA",X"A8",X"AA",X"A8",X"AA",X"A8",X"AA",X"A8",X"AA",X"A8",
		X"55",X"50",X"55",X"50",X"55",X"50",X"00",X"00",X"AA",X"A0",X"AA",X"A8",X"FF",X"FF",X"FF",X"FF",
		X"55",X"50",X"55",X"50",X"55",X"50",X"55",X"50",X"55",X"50",X"55",X"50",X"55",X"50",X"55",X"50",
		X"55",X"50",X"55",X"50",X"55",X"50",X"55",X"50",X"55",X"50",X"55",X"50",X"55",X"50",X"55",X"50",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"FF",X"FF",X"FF",X"FF",
		X"A6",X"6A",X"A6",X"6A",X"AE",X"6A",X"AA",X"EA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"A5",X"5A",X"A6",X"AA",X"A5",X"5A",X"A6",X"AA",X"A5",X"5A",X"AA",X"AA",X"A5",X"5A",
		X"AA",X"AA",X"A5",X"5A",X"A6",X"9A",X"A6",X"9A",X"A9",X"6A",X"AA",X"AA",X"A5",X"5A",X"AA",X"9A",
		X"A5",X"5A",X"AA",X"9A",X"A5",X"5A",X"AA",X"AA",X"A5",X"5A",X"A6",X"6A",X"A5",X"5A",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"05",X"00",X"05",X"00",X"15",X"00",X"15",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"AA",X"95",X"55",X"95",X"55",X"95",X"55",X"95",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"55",X"00",X"55",X"00",
		X"55",X"00",X"55",X"00",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"0F",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",
		X"08",X"00",X"08",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"80",X"0A",X"80",X"02",X"A0",X"02",X"A8",
		X"02",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"2A",X"00",X"0A",X"00",X"02",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"0C",
		X"55",X"5A",X"55",X"5A",X"55",X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"15",X"00",X"00",
		X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"15",X"51",X"95",X"00",X"00",
		X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"15",X"51",X"95",X"59",X"95",X"00",X"00",
		X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"15",X"51",X"95",X"59",X"95",X"59",X"95",X"00",X"00",
		X"00",X"00",X"55",X"15",X"51",X"95",X"59",X"95",X"59",X"95",X"59",X"95",X"6A",X"AA",X"00",X"00",
		X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"57",X"00",X"00",X"00",
		X"00",X"00",X"51",X"95",X"59",X"95",X"59",X"95",X"59",X"95",X"6A",X"AA",X"2A",X"AA",X"00",X"00",
		X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"5C",X"01",X"5C",X"C1",X"5C",X"00",X"00",X"00",
		X"55",X"55",X"50",X"00",X"50",X"00",X"51",X"54",X"51",X"54",X"50",X"00",X"50",X"00",X"55",X"55",
		X"55",X"55",X"51",X"54",X"51",X"54",X"50",X"00",X"50",X"00",X"55",X"54",X"55",X"54",X"55",X"55",
		X"55",X"55",X"51",X"00",X"51",X"00",X"51",X"14",X"51",X"14",X"50",X"14",X"50",X"14",X"55",X"55",
		X"55",X"55",X"51",X"14",X"51",X"14",X"51",X"14",X"51",X"14",X"50",X"00",X"50",X"00",X"55",X"55",
		X"55",X"55",X"54",X"05",X"54",X"05",X"55",X"45",X"55",X"45",X"50",X"00",X"50",X"00",X"55",X"55",
		X"55",X"55",X"50",X"14",X"51",X"14",X"51",X"14",X"51",X"14",X"51",X"00",X"51",X"00",X"55",X"55",
		X"55",X"55",X"50",X"00",X"50",X"00",X"51",X"44",X"51",X"44",X"51",X"40",X"51",X"40",X"55",X"55",
		X"55",X"55",X"55",X"55",X"50",X"55",X"51",X"55",X"51",X"55",X"50",X"00",X"50",X"00",X"55",X"55",
		X"55",X"55",X"50",X"00",X"50",X"00",X"51",X"14",X"51",X"14",X"50",X"00",X"50",X"00",X"55",X"55",
		X"55",X"55",X"50",X"04",X"50",X"04",X"51",X"44",X"51",X"44",X"50",X"00",X"50",X"00",X"55",X"55",
		X"00",X"00",X"59",X"95",X"59",X"95",X"6A",X"AA",X"6A",X"AA",X"2A",X"AA",X"2A",X"AA",X"00",X"00",
		X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"15",X"51",X"95",X"59",X"95",X"00",X"00",
		X"00",X"00",X"55",X"55",X"55",X"55",X"57",X"00",X"57",X"30",X"57",X"00",X"57",X"00",X"00",X"00",
		X"00",X"00",X"6A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"6A",X"AA",X"55",X"55",X"00",X"00",
		X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"15",X"51",X"95",X"59",X"95",X"59",X"95",X"00",X"00",
		X"00",X"00",X"55",X"55",X"57",X"00",X"57",X"30",X"57",X"00",X"57",X"00",X"57",X"FF",X"00",X"00",
		X"00",X"00",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"6A",X"AA",X"55",X"55",X"55",X"55",X"00",X"00",
		X"55",X"55",X"50",X"00",X"50",X"00",X"51",X"45",X"51",X"45",X"50",X"00",X"50",X"00",X"55",X"55",
		X"55",X"55",X"50",X"00",X"50",X"00",X"50",X"44",X"50",X"44",X"50",X"00",X"55",X"40",X"55",X"55",
		X"55",X"55",X"50",X"00",X"50",X"00",X"51",X"54",X"51",X"54",X"51",X"54",X"51",X"54",X"55",X"55",
		X"55",X"55",X"50",X"00",X"50",X"00",X"51",X"54",X"50",X"50",X"50",X"00",X"54",X"01",X"55",X"55",
		X"55",X"55",X"50",X"00",X"50",X"00",X"51",X"14",X"51",X"14",X"51",X"14",X"51",X"54",X"55",X"55",
		X"55",X"55",X"50",X"00",X"50",X"00",X"51",X"45",X"51",X"45",X"51",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"50",X"00",X"50",X"00",X"51",X"54",X"51",X"54",X"51",X"40",X"51",X"40",X"55",X"55",
		X"55",X"55",X"50",X"00",X"50",X"00",X"55",X"45",X"55",X"45",X"50",X"00",X"50",X"00",X"55",X"55",
		X"55",X"55",X"51",X"54",X"51",X"54",X"50",X"00",X"50",X"00",X"51",X"54",X"51",X"54",X"55",X"55",
		X"55",X"55",X"55",X"40",X"55",X"40",X"51",X"54",X"51",X"54",X"50",X"00",X"50",X"00",X"51",X"55",
		X"55",X"55",X"50",X"00",X"50",X"00",X"54",X"05",X"50",X"41",X"51",X"50",X"51",X"54",X"55",X"55",
		X"55",X"55",X"50",X"00",X"50",X"00",X"55",X"54",X"55",X"54",X"55",X"50",X"55",X"50",X"55",X"55",
		X"55",X"55",X"50",X"00",X"50",X"00",X"51",X"55",X"50",X"00",X"51",X"55",X"50",X"00",X"55",X"55",
		X"55",X"55",X"50",X"00",X"50",X"00",X"54",X"15",X"55",X"01",X"50",X"00",X"50",X"00",X"55",X"55",
		X"55",X"55",X"50",X"00",X"50",X"00",X"51",X"54",X"51",X"54",X"50",X"00",X"50",X"00",X"55",X"55",
		X"55",X"55",X"50",X"00",X"50",X"00",X"51",X"45",X"51",X"45",X"50",X"05",X"50",X"05",X"55",X"55",
		X"55",X"55",X"50",X"00",X"50",X"00",X"51",X"54",X"51",X"50",X"50",X"00",X"50",X"00",X"55",X"55",
		X"55",X"55",X"50",X"00",X"50",X"00",X"51",X"15",X"51",X"05",X"50",X"00",X"50",X"10",X"55",X"55",
		X"55",X"55",X"50",X"14",X"51",X"14",X"51",X"14",X"51",X"00",X"51",X"00",X"55",X"55",X"55",X"55",
		X"55",X"55",X"50",X"55",X"51",X"54",X"50",X"00",X"50",X"00",X"51",X"54",X"50",X"55",X"55",X"55",
		X"55",X"55",X"50",X"00",X"50",X"00",X"55",X"54",X"55",X"54",X"50",X"00",X"50",X"00",X"55",X"55",
		X"55",X"55",X"51",X"55",X"50",X"05",X"50",X"00",X"55",X"40",X"50",X"05",X"51",X"55",X"55",X"55",
		X"55",X"55",X"50",X"00",X"50",X"00",X"55",X"54",X"50",X"00",X"55",X"54",X"50",X"00",X"55",X"55",
		X"55",X"55",X"51",X"54",X"50",X"40",X"55",X"05",X"50",X"15",X"50",X"45",X"51",X"50",X"55",X"55",
		X"55",X"55",X"51",X"55",X"50",X"15",X"54",X"00",X"55",X"00",X"50",X"55",X"51",X"55",X"55",X"55",
		X"55",X"55",X"51",X"50",X"51",X"40",X"51",X"04",X"50",X"14",X"50",X"54",X"51",X"54",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"55",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"55",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"6A",X"AA",X"6A",X"AA",X"5A",X"AA",X"5A",X"AA",X"02",X"AA",X"02",X"AA",
		X"55",X"40",X"55",X"40",X"55",X"40",X"55",X"40",X"55",X"40",X"55",X"40",X"55",X"40",X"55",X"40",
		X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",
		X"00",X"55",X"01",X"55",X"01",X"55",X"05",X"55",X"15",X"55",X"15",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"55",X"15",X"51",X"95",X"59",X"95",X"59",X"95",X"59",X"95",X"6A",X"AA",X"00",X"00",
		X"00",X"00",X"57",X"00",X"57",X"00",X"57",X"00",X"57",X"FF",X"55",X"55",X"55",X"55",X"00",X"00",
		X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A9",X"FF",X"00",X"00",
		X"00",X"00",X"51",X"95",X"59",X"95",X"6A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"00",X"00",
		X"00",X"00",X"55",X"55",X"55",X"55",X"57",X"00",X"57",X"30",X"57",X"00",X"57",X"00",X"00",X"00",
		X"00",X"00",X"59",X"95",X"6A",X"AA",X"2A",X"AA",X"2A",X"AA",X"6A",X"AA",X"55",X"55",X"00",X"00",
		X"00",X"00",X"55",X"55",X"57",X"00",X"57",X"30",X"57",X"00",X"57",X"00",X"57",X"FF",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"6A",X"AA",X"6A",X"AA",X"5A",X"AA",
		X"00",X"00",X"2A",X"AA",X"2A",X"AA",X"6A",X"AA",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"00",
		X"00",X"00",X"55",X"C0",X"55",X"C0",X"55",X"FF",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"00",
		X"00",X"00",X"55",X"FF",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"00",
		X"56",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"6A",X"55",X"5A",X"55",X"5A",X"55",X"56",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"20",X"02",X"20",X"02",X"20",X"2A",X"AA",X"2A",X"AA",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"15",X"30",X"15",X"00",X"15",X"00",X"15",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"0A",X"CC",X"0A",X"C0",X"0A",X"C0",X"0A",X"FF",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"33",X"00",X"30",X"00",X"30",X"00",X"3F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0F",X"00",X"00",
		X"55",X"45",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"59",X"95",X"51",X"95",X"55",X"15",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"59",X"95",X"59",X"95",X"59",X"95",X"51",X"95",X"55",X"15",X"55",X"55",X"55",X"55",X"55",X"55",
		X"2A",X"AA",X"6A",X"AA",X"59",X"95",X"59",X"95",X"59",X"95",X"51",X"95",X"55",X"15",X"55",X"55",
		X"56",X"FF",X"56",X"FF",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"2A",X"AA",X"2A",X"AA",X"6A",X"AA",X"59",X"95",X"59",X"95",X"59",X"95",X"51",X"95",X"55",X"15",
		X"5C",X"00",X"5C",X"00",X"5C",X"81",X"5C",X"01",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"6A",X"AA",X"2A",X"AA",X"2A",X"AA",X"6A",X"AA",X"6A",X"AA",X"59",X"95",X"59",X"95",X"51",X"95",
		X"57",X"00",X"57",X"00",X"57",X"00",X"57",X"30",X"57",X"00",X"55",X"55",X"55",X"55",X"55",X"55",
		X"59",X"95",X"59",X"95",X"51",X"95",X"55",X"15",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"6A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"6A",X"AA",X"55",X"55",X"55",X"55",
		X"59",X"95",X"59",X"95",X"59",X"95",X"51",X"95",X"55",X"15",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"57",X"FF",X"57",X"00",X"57",X"00",X"57",X"30",X"57",X"00",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"6A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"6A",X"AA",
		X"2A",X"AA",X"6A",X"AA",X"59",X"95",X"59",X"95",X"59",X"95",X"51",X"95",X"55",X"15",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"57",X"FF",X"57",X"00",X"57",X"00",X"57",X"00",X"57",X"00",
		X"57",X"30",X"57",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"6A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"6A",X"AA",X"59",X"95",X"51",X"95",X"55",X"15",
		X"57",X"FF",X"57",X"00",X"57",X"00",X"57",X"30",X"57",X"00",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"6A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"6A",X"AA",X"59",X"95",X"59",X"95",
		X"55",X"55",X"57",X"FF",X"57",X"00",X"57",X"00",X"57",X"30",X"57",X"00",X"55",X"55",X"55",X"55",
		X"55",X"55",X"FF",X"D5",X"C0",X"1A",X"C0",X"0A",X"CC",X"0A",X"C0",X"1A",X"55",X"55",X"55",X"55",
		X"55",X"55",X"FF",X"D5",X"C0",X"1A",X"C0",X"0A",X"CC",X"0A",X"C0",X"1A",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"7F",X"55",X"70",X"55",X"70",X"55",X"73",X"55",X"70",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"5F",X"55",X"5C",X"55",X"5C",X"55",X"5C",X"55",X"5C",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"A5",X"AA",X"AA",X"5A",X"AA",X"5A",X"A5",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"6A",X"AA",X"6A",X"AA",X"5A",X"AA",X"56",X"AA",X"55",X"AA",X"55",X"6A",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"6A",X"AA",X"5A",X"AA",
		X"56",X"AA",X"56",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"6A",X"55",X"5A",X"55",X"56",X"55",X"56",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"50",X"55",X"50",X"55",X"40",X"55",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"2A",X"AA",X"0A",X"AA",X"5A",X"AA",X"56",X"AA",X"55",X"AA",X"55",X"AA",
		X"54",X"00",X"50",X"00",X"40",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"AA",X"02",X"AA",X"00",X"AA",X"00",X"2A",X"00",X"2A",X"00",X"0A",X"00",X"0A",X"00",X"02",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"2A",X"AA",X"2A",X"AA",X"0A",X"AA",
		X"6A",X"AA",X"6A",X"AA",X"00",X"0A",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"5A",X"55",X"5A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"50",X"55",X"50",X"55",X"40",X"55",X"00",X"55",X"00",X"54",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"5A",X"55",X"5A",X"55",X"5A",X"55",X"5A",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"02",X"AA",X"00",X"AA",X"00",X"2A",X"00",X"2A",X"C0",X"0A",X"FF",X"0A",X"00",X"00",X"C0",X"00",
		X"55",X"57",X"55",X"57",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"AA",X"FF",X"AA",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"2A",X"AA",X"0A",X"AA",X"0A",X"AA",
		X"54",X"00",X"54",X"00",X"54",X"00",X"55",X"00",X"55",X"00",X"55",X"40",X"55",X"40",X"55",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"2A",X"00",X"2A",X"00",X"0A",X"00",X"02",X"00",X"02",X"FF",X"C0",X"C0",X"00",X"C0",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"40",X"55",X"00",X"55",X"00",X"54",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"2A",X"AA",X"0A",X"AA",X"0A",X"AA",X"02",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"2A",
		X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",
		X"0A",X"AA",X"02",X"AA",X"00",X"AA",X"80",X"2A",X"00",X"2A",X"00",X"0A",X"A8",X"0A",X"00",X"00",
		X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"54",X"00",X"54",X"00",X"54",X"00",X"54",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"40",X"55",X"40",X"55",X"40",X"55",X"40",X"55",X"00",
		X"00",X"AA",X"00",X"2A",X"28",X"0A",X"00",X"02",X"00",X"02",X"0C",X"02",X"02",X"A0",X"02",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"0A",X"AA",X"0A",X"AA",X"02",X"AA",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"56",X"55",X"6A",X"55",X"AA",X"5A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"6A",
		X"02",X"AA",X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"AA",X"02",X"AA",X"2A",X"AA",X"AA",X"AA",
		X"55",X"56",X"55",X"6A",X"55",X"AA",X"5A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"55",X"AA",X"56",X"AA",X"5A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"6A",X"56",X"AA",X"5A",X"AA",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"6A",X"55",X"56",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"AA",X"AA",X"AA",X"AA",X"6A",X"AA",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"55",X"FF",X"55",X"FF",
		X"55",X"55",X"55",X"55",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FF",X"FF",X"FF",X"FF",
		X"55",X"55",X"55",X"55",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FF",X"AA",X"FF",X"AA",
		X"55",X"55",X"55",X"55",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"AA",X"FF",X"AA",X"00",X"AA",X"02",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",
		X"55",X"FF",X"55",X"FF",X"55",X"00",X"55",X"40",X"55",X"50",X"55",X"54",X"55",X"55",X"55",X"55",
		X"55",X"6A",X"55",X"5A",X"55",X"56",X"55",X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"57",X"67",X"67",X"67",X"65",X"67",X"66",X"65",X"56",X"67",X"76",X"57",X"75",X"77",X"76",X"77",
		X"AA",X"57",X"AA",X"67",X"AA",X"67",X"AA",X"65",X"AA",X"67",X"AA",X"57",X"AA",X"77",X"AA",X"75",
		X"55",X"55",X"55",X"41",X"41",X"14",X"40",X"04",X"41",X"14",X"51",X"14",X"55",X"41",X"55",X"55",
		X"55",X"55",X"55",X"55",X"51",X"04",X"51",X"15",X"51",X"15",X"50",X"15",X"55",X"55",X"55",X"55",
		X"00",X"00",X"15",X"54",X"14",X"14",X"11",X"44",X"11",X"44",X"11",X"44",X"15",X"54",X"00",X"00",
		X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"56",X"AA",X"56",X"AA",X"55",X"AA",X"55",X"6A",X"55",X"56",
		X"55",X"56",X"55",X"6A",X"55",X"AA",X"56",X"AA",X"56",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",
		X"AA",X"A5",X"AA",X"A5",X"AA",X"A5",X"AA",X"95",X"AA",X"95",X"AA",X"55",X"A9",X"55",X"95",X"55",
		X"95",X"55",X"A9",X"55",X"AA",X"55",X"AA",X"95",X"AA",X"95",X"AA",X"A5",X"AA",X"A5",X"AA",X"A5",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"00",X"C0",X"00",X"0C",X"03",X"0C",X"08",X"38",X"00",X"30",X"00",X"00",X"00",X"00",X"00",
		X"02",X"00",X"00",X"E0",X"00",X"30",X"00",X"0F",X"00",X"00",X"FF",X"FF",X"03",X"03",X"0C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"C0",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"20",X"00",X"C0",X"00",X"CF",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"AA",X"00",X"00",X"A3",X"00",X"80",X"C0",X"00",X"30",X"0F",X"FF",X"00",X"00",X"00",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"A8",X"00",X"2A",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"00",X"00",X"80",X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"28",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0C",X"00",X"0C",X"00",X"0C",X"FF",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",
		X"00",X"0C",X"00",X"0C",X"00",X"0C",X"FF",X"FC",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FC",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"E0",X"00",X"E0",X"00",X"E0",X"00",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",
		X"C0",X"00",X"C0",X"00",X"C0",X"00",X"FF",X"FF",X"C0",X"08",X"C0",X"08",X"C0",X"08",X"C0",X"08",
		X"C0",X"00",X"C0",X"00",X"C0",X"00",X"FF",X"FF",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"08",
		X"30",X"00",X"30",X"00",X"30",X"00",X"3F",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"00",X"30",X"00",X"30",X"00",X"30",X"00",X"30",X"00",X"30",X"00",X"30",X"00",X"30",X"00",
		X"30",X"00",X"30",X"00",X"30",X"00",X"3F",X"FF",X"30",X"00",X"30",X"00",X"30",X"00",X"30",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"FF",X"30",X"00",X"30",X"00",X"30",X"00",X"30",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
