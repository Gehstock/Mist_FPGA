library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity cpu0_rom is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of cpu0_rom is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"F3",X"ED",X"56",X"C3",X"E6",X"00",X"FF",X"FF",X"87",X"30",X"05",X"24",X"C3",X"10",X"00",X"00",
		X"85",X"6F",X"D0",X"24",X"C9",X"00",X"00",X"00",X"C0",X"3E",X"9C",X"77",X"C9",X"00",X"00",X"00",
		X"FE",X"64",X"D8",X"D6",X"64",X"18",X"F9",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C3",X"80",X"02",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"21",X"00",X"60",X"32",X"30",X"68",
		X"2B",X"7D",X"B4",X"20",X"F8",X"C9",X"D9",X"ED",X"A0",X"EA",X"9E",X"00",X"F5",X"2A",X"00",X"89",
		X"7E",X"A7",X"CA",X"98",X"00",X"36",X"00",X"F5",X"2C",X"2C",X"4E",X"2C",X"46",X"2C",X"5E",X"2C",
		X"56",X"2C",X"7E",X"2C",X"2C",X"22",X"00",X"89",X"2D",X"66",X"6F",X"3E",X"10",X"32",X"00",X"71",
		X"F1",X"D9",X"32",X"00",X"71",X"F1",X"ED",X"45",X"3E",X"10",X"32",X"00",X"71",X"F1",X"D9",X"ED",
		X"45",X"08",X"F3",X"3A",X"00",X"71",X"E6",X"E0",X"20",X"07",X"08",X"D9",X"32",X"00",X"71",X"FB",
		X"C9",X"E5",X"D5",X"EB",X"2A",X"02",X"89",X"7D",X"C6",X"08",X"6F",X"22",X"02",X"89",X"2D",X"72",
		X"2D",X"73",X"2D",X"D1",X"72",X"2D",X"73",X"2D",X"70",X"2D",X"71",X"32",X"30",X"68",X"2D",X"2D",
		X"08",X"77",X"3A",X"00",X"71",X"FE",X"10",X"28",X"03",X"E1",X"FB",X"C9",X"7E",X"36",X"00",X"22",
		X"02",X"89",X"E1",X"C3",X"AA",X"00",X"3E",X"10",X"32",X"00",X"71",X"32",X"00",X"70",X"21",X"20",
		X"68",X"77",X"23",X"77",X"23",X"36",X"01",X"23",X"77",X"3C",X"32",X"30",X"68",X"23",X"23",X"3E",
		X"FF",X"77",X"23",X"77",X"23",X"77",X"AF",X"21",X"E0",X"89",X"06",X"0B",X"77",X"23",X"10",X"FC",
		X"21",X"EF",X"89",X"06",X"04",X"77",X"23",X"10",X"FC",X"C3",X"7E",X"38",X"F3",X"AF",X"32",X"20",
		X"68",X"21",X"07",X"A0",X"77",X"21",X"1B",X"9B",X"36",X"10",X"3E",X"88",X"21",X"00",X"84",X"36",
		X"00",X"32",X"30",X"68",X"23",X"BC",X"20",X"F7",X"3E",X"94",X"21",X"00",X"90",X"36",X"00",X"32",
		X"30",X"68",X"23",X"BC",X"20",X"F7",X"21",X"33",X"9B",X"36",X"00",X"21",X"80",X"9A",X"06",X"20",
		X"36",X"00",X"32",X"30",X"68",X"23",X"10",X"F8",X"21",X"00",X"98",X"01",X"80",X"01",X"32",X"30",
		X"68",X"36",X"00",X"23",X"0B",X"78",X"B1",X"20",X"F5",X"3E",X"01",X"32",X"23",X"68",X"3A",X"D0",
		X"89",X"FE",X"00",X"CA",X"00",X"00",X"FE",X"FF",X"20",X"08",X"3E",X"00",X"32",X"C0",X"87",X"C3",
		X"B4",X"01",X"21",X"AA",X"85",X"36",X"00",X"23",X"E6",X"0F",X"77",X"3A",X"D1",X"89",X"FE",X"FF",
		X"20",X"08",X"3E",X"01",X"32",X"C0",X"87",X"C3",X"B4",X"01",X"47",X"21",X"AC",X"85",X"36",X"00",
		X"23",X"E6",X"0F",X"77",X"78",X"E6",X"F0",X"FE",X"10",X"20",X"04",X"3E",X"02",X"18",X"02",X"3E",
		X"03",X"32",X"C0",X"87",X"31",X"00",X"9A",X"CD",X"5A",X"00",X"21",X"00",X"88",X"22",X"00",X"89",
		X"22",X"02",X"89",X"AF",X"21",X"00",X"A0",X"06",X"04",X"36",X"00",X"23",X"10",X"FB",X"CD",X"5A",
		X"00",X"21",X"04",X"89",X"06",X"04",X"36",X"02",X"23",X"10",X"FB",X"21",X"04",X"89",X"11",X"00",
		X"70",X"01",X"04",X"00",X"3E",X"C1",X"CD",X"A1",X"00",X"CD",X"A6",X"15",X"21",X"00",X"80",X"06",
		X"40",X"36",X"7F",X"23",X"32",X"30",X"68",X"10",X"F8",X"21",X"ED",X"83",X"11",X"09",X"00",X"06",
		X"02",X"3E",X"10",X"77",X"23",X"77",X"19",X"10",X"FA",X"CD",X"A3",X"19",X"CD",X"4F",X"14",X"CD",
		X"32",X"14",X"3E",X"FF",X"32",X"87",X"87",X"21",X"27",X"89",X"11",X"AE",X"89",X"06",X"03",X"1A",
		X"77",X"23",X"1B",X"10",X"FA",X"CD",X"DE",X"14",X"3E",X"01",X"21",X"A9",X"87",X"77",X"23",X"77",
		X"23",X"77",X"32",X"05",X"9A",X"32",X"20",X"68",X"FB",X"31",X"00",X"9A",X"21",X"00",X"84",X"CB",
		X"4E",X"20",X"08",X"21",X"14",X"84",X"3A",X"0D",X"84",X"18",X"06",X"21",X"17",X"84",X"3A",X"0E",
		X"84",X"47",X"3A",X"CC",X"87",X"CB",X"4F",X"28",X"19",X"CB",X"57",X"20",X"15",X"78",X"E5",X"F5",
		X"CD",X"F2",X"0B",X"F1",X"E1",X"CD",X"F0",X"32",X"21",X"03",X"A0",X"36",X"00",X"21",X"CC",X"87",
		X"CB",X"8E",X"21",X"CC",X"87",X"CB",X"46",X"28",X"05",X"CB",X"86",X"CD",X"E3",X"35",X"18",X"B8",
		X"DD",X"E5",X"FD",X"E5",X"E5",X"D5",X"C5",X"F5",X"AF",X"32",X"20",X"68",X"32",X"30",X"68",X"3A",
		X"9A",X"87",X"A7",X"20",X"2B",X"21",X"00",X"98",X"11",X"80",X"8B",X"01",X"80",X"00",X"C5",X"ED",
		X"B0",X"C1",X"21",X"00",X"99",X"11",X"80",X"9B",X"ED",X"B0",X"3A",X"CF",X"87",X"CB",X"6F",X"CA",
		X"27",X"0A",X"3A",X"8E",X"89",X"21",X"00",X"84",X"2F",X"E6",X"04",X"B6",X"77",X"CD",X"B1",X"0B",
		X"2A",X"23",X"84",X"23",X"22",X"23",X"84",X"3A",X"9A",X"87",X"A7",X"20",X"06",X"3A",X"A5",X"85",
		X"32",X"A6",X"85",X"21",X"00",X"70",X"11",X"A7",X"85",X"01",X"03",X"00",X"3E",X"71",X"CD",X"A1",
		X"00",X"3A",X"9A",X"87",X"A7",X"C2",X"27",X"0A",X"21",X"A7",X"87",X"CB",X"46",X"28",X"26",X"CB",
		X"86",X"21",X"11",X"84",X"AF",X"77",X"23",X"3A",X"E7",X"87",X"77",X"23",X"AF",X"77",X"CD",X"C8",
		X"2F",X"3A",X"57",X"86",X"CB",X"4F",X"20",X"0D",X"CD",X"6B",X"14",X"3A",X"00",X"84",X"CB",X"5F",
		X"20",X"03",X"CD",X"DF",X"0B",X"21",X"00",X"84",X"CB",X"4E",X"20",X"14",X"3A",X"A8",X"85",X"47",
		X"E6",X"0F",X"FE",X"09",X"38",X"02",X"CB",X"98",X"78",X"CB",X"87",X"32",X"B0",X"85",X"18",X"0C",
		X"CB",X"56",X"28",X"E8",X"3A",X"A9",X"85",X"18",X"E6",X"32",X"B0",X"85",X"21",X"24",X"86",X"11",
		X"B0",X"85",X"1A",X"E6",X"30",X"77",X"21",X"A5",X"85",X"11",X"A6",X"85",X"3A",X"A7",X"85",X"77",
		X"FE",X"B0",X"D2",X"7E",X"38",X"E6",X"0F",X"FE",X"0A",X"D2",X"7E",X"38",X"7E",X"A7",X"20",X"0E",
		X"1A",X"A7",X"20",X"0A",X"3A",X"00",X"84",X"CB",X"77",X"CA",X"80",X"0A",X"18",X"5A",X"3A",X"CC",
		X"87",X"CB",X"4F",X"20",X"16",X"CB",X"47",X"20",X"12",X"1A",X"47",X"7E",X"FE",X"90",X"30",X"0B",
		X"90",X"27",X"4F",X"38",X"06",X"28",X"04",X"79",X"32",X"33",X"9B",X"7E",X"EB",X"BE",X"30",X"30",
		X"1A",X"FE",X"99",X"28",X"0A",X"FE",X"9F",X"28",X"06",X"C6",X"01",X"27",X"BE",X"20",X"14",X"21",
		X"00",X"84",X"CB",X"86",X"CB",X"8E",X"CB",X"F6",X"3E",X"01",X"21",X"E1",X"89",X"CD",X"26",X"12",
		X"C3",X"27",X"0A",X"21",X"00",X"84",X"CB",X"C6",X"CB",X"8E",X"CB",X"F6",X"3E",X"02",X"18",X"EA",
		X"21",X"00",X"84",X"CB",X"76",X"CA",X"03",X"0B",X"21",X"57",X"86",X"CB",X"86",X"CB",X"4E",X"C2",
		X"27",X"0A",X"21",X"F3",X"89",X"34",X"21",X"88",X"9A",X"7E",X"A7",X"C2",X"27",X"0A",X"21",X"00",
		X"84",X"CB",X"5E",X"C2",X"45",X"04",X"CB",X"DE",X"CD",X"A6",X"15",X"CD",X"7C",X"17",X"CD",X"ED",
		X"17",X"CD",X"7F",X"18",X"CD",X"92",X"18",X"CD",X"5A",X"00",X"3A",X"B0",X"85",X"CB",X"6F",X"28",
		X"05",X"21",X"87",X"87",X"36",X"FF",X"CD",X"22",X"0C",X"3A",X"CF",X"87",X"CB",X"5F",X"20",X"19",
		X"3A",X"87",X"87",X"CB",X"4F",X"20",X"12",X"3A",X"0E",X"84",X"6F",X"67",X"32",X"0F",X"84",X"22",
		X"27",X"86",X"21",X"85",X"87",X"36",X"00",X"18",X"10",X"3E",X"01",X"32",X"0F",X"84",X"21",X"01",
		X"01",X"22",X"27",X"86",X"21",X"85",X"87",X"36",X"00",X"CD",X"AC",X"18",X"CD",X"B1",X"12",X"CD",
		X"51",X"0C",X"C3",X"27",X"0A",X"CB",X"7E",X"20",X"47",X"CB",X"FE",X"CD",X"AE",X"17",X"CD",X"15",
		X"0C",X"CD",X"51",X"15",X"21",X"00",X"00",X"3A",X"00",X"84",X"CB",X"4F",X"20",X"09",X"AF",X"32",
		X"DA",X"87",X"22",X"D4",X"87",X"18",X"07",X"AF",X"32",X"D8",X"87",X"22",X"D2",X"87",X"32",X"99",
		X"87",X"32",X"EB",X"87",X"22",X"ED",X"87",X"32",X"6D",X"89",X"32",X"6C",X"89",X"32",X"F0",X"87",
		X"21",X"9E",X"98",X"77",X"23",X"36",X"E0",X"CD",X"A6",X"0B",X"CD",X"B1",X"0B",X"C3",X"27",X"0A",
		X"21",X"00",X"84",X"CB",X"66",X"20",X"33",X"CB",X"E6",X"CD",X"F7",X"19",X"3A",X"27",X"86",X"3D",
		X"4F",X"D6",X"0C",X"30",X"FB",X"79",X"1F",X"1F",X"4F",X"E6",X"01",X"32",X"04",X"A0",X"79",X"1F",
		X"E6",X"01",X"32",X"05",X"A0",X"CD",X"05",X"0C",X"CD",X"0B",X"14",X"CD",X"45",X"18",X"CD",X"51",
		X"15",X"CD",X"A6",X"0B",X"CD",X"B1",X"0B",X"C3",X"27",X"0A",X"E5",X"3A",X"57",X"86",X"CB",X"4F",
		X"20",X"06",X"CD",X"81",X"0C",X"CD",X"6B",X"14",X"E1",X"CB",X"6E",X"C2",X"C7",X"05",X"CB",X"EE",
		X"21",X"68",X"10",X"22",X"25",X"86",X"AF",X"32",X"4A",X"86",X"32",X"53",X"86",X"CD",X"F7",X"19",
		X"CD",X"51",X"15",X"21",X"4B",X"86",X"06",X"08",X"0E",X"02",X"3A",X"57",X"86",X"CB",X"47",X"20",
		X"11",X"3A",X"27",X"86",X"FE",X"14",X"38",X"0A",X"FE",X"20",X"30",X"04",X"0E",X"01",X"18",X"02",
		X"0E",X"00",X"3E",X"02",X"77",X"23",X"91",X"10",X"FB",X"CD",X"EC",X"11",X"CD",X"E0",X"11",X"21",
		X"A1",X"83",X"11",X"20",X"00",X"19",X"3E",X"7F",X"77",X"23",X"77",X"19",X"77",X"2B",X"77",X"21",
		X"9E",X"98",X"AF",X"77",X"23",X"36",X"E0",X"32",X"EF",X"87",X"32",X"F0",X"87",X"21",X"00",X"00",
		X"22",X"D6",X"87",X"32",X"6F",X"89",X"32",X"6C",X"89",X"32",X"A7",X"87",X"32",X"B3",X"85",X"32",
		X"22",X"99",X"21",X"28",X"85",X"11",X"10",X"00",X"0E",X"00",X"06",X"08",X"CB",X"7E",X"28",X"01",
		X"0C",X"19",X"10",X"F8",X"79",X"FE",X"08",X"20",X"0F",X"CD",X"7D",X"1B",X"21",X"6C",X"89",X"CB",
		X"DE",X"21",X"01",X"84",X"CB",X"EE",X"18",X"0E",X"CD",X"2E",X"1B",X"CD",X"7D",X"1B",X"CD",X"45",
		X"18",X"21",X"01",X"84",X"CB",X"AE",X"21",X"93",X"9A",X"36",X"00",X"21",X"87",X"87",X"36",X"FF",
		X"CD",X"A6",X"0B",X"CD",X"B1",X"0B",X"3E",X"02",X"32",X"AE",X"85",X"32",X"AF",X"85",X"21",X"E0",
		X"01",X"22",X"F2",X"85",X"21",X"01",X"84",X"CB",X"B6",X"32",X"30",X"68",X"21",X"00",X"00",X"22",
		X"F4",X"85",X"3A",X"57",X"86",X"CB",X"4F",X"28",X"05",X"3E",X"80",X"32",X"76",X"86",X"CD",X"A6",
		X"0B",X"CD",X"B1",X"0B",X"C3",X"27",X"0A",X"3A",X"6C",X"89",X"CB",X"5F",X"20",X"61",X"21",X"01",
		X"84",X"CB",X"6E",X"20",X"30",X"E5",X"CD",X"94",X"1C",X"3E",X"78",X"32",X"D5",X"85",X"E1",X"CB",
		X"EE",X"21",X"85",X"87",X"3A",X"00",X"84",X"CB",X"4F",X"20",X"0D",X"CB",X"46",X"C2",X"27",X"0A",
		X"3E",X"01",X"32",X"81",X"9A",X"C3",X"27",X"0A",X"CB",X"4E",X"C2",X"27",X"0A",X"3E",X"01",X"32",
		X"81",X"9A",X"C3",X"27",X"0A",X"21",X"81",X"9A",X"7E",X"A7",X"C2",X"27",X"0A",X"3A",X"D5",X"85",
		X"A7",X"28",X"0C",X"FE",X"01",X"CC",X"D3",X"1C",X"21",X"D5",X"85",X"35",X"C3",X"27",X"0A",X"21",
		X"85",X"87",X"3A",X"00",X"84",X"CB",X"4F",X"20",X"04",X"CB",X"C6",X"18",X"02",X"CB",X"CE",X"21",
		X"6C",X"89",X"CB",X"DE",X"3A",X"46",X"86",X"CB",X"4F",X"28",X"19",X"21",X"86",X"9A",X"3E",X"00",
		X"77",X"21",X"89",X"9A",X"77",X"21",X"47",X"86",X"7E",X"A7",X"20",X"07",X"21",X"01",X"84",X"CB",
		X"FE",X"18",X"01",X"35",X"21",X"6F",X"89",X"CB",X"46",X"20",X"15",X"CB",X"C6",X"21",X"00",X"00",
		X"22",X"23",X"84",X"AF",X"21",X"B0",X"85",X"CD",X"64",X"19",X"21",X"F4",X"85",X"77",X"23",X"77",
		X"21",X"F0",X"87",X"CB",X"4E",X"C2",X"49",X"09",X"21",X"01",X"84",X"CB",X"7E",X"CA",X"49",X"09",
		X"AF",X"32",X"92",X"9A",X"23",X"CB",X"46",X"C2",X"98",X"07",X"21",X"1C",X"86",X"35",X"7E",X"FE",
		X"64",X"C2",X"F7",X"06",X"21",X"46",X"86",X"CB",X"4E",X"28",X"02",X"36",X"80",X"21",X"32",X"85",
		X"06",X"08",X"11",X"10",X"00",X"36",X"00",X"19",X"32",X"30",X"68",X"10",X"F8",X"21",X"9E",X"98",
		X"36",X"00",X"23",X"36",X"E0",X"21",X"26",X"85",X"06",X"08",X"11",X"0E",X"00",X"CB",X"B6",X"23",
		X"23",X"CB",X"B6",X"19",X"32",X"30",X"68",X"10",X"F4",X"21",X"2B",X"85",X"11",X"10",X"00",X"06",
		X"08",X"36",X"32",X"19",X"32",X"30",X"68",X"10",X"F8",X"21",X"4A",X"86",X"36",X"00",X"CD",X"51",
		X"15",X"CD",X"89",X"0F",X"AF",X"32",X"A0",X"98",X"32",X"A1",X"98",X"21",X"F4",X"98",X"06",X"0C",
		X"77",X"23",X"10",X"FC",X"C3",X"27",X"0A",X"FE",X"50",X"C2",X"1B",X"07",X"3E",X"01",X"32",X"85",
		X"9A",X"21",X"22",X"98",X"36",X"14",X"21",X"46",X"86",X"CB",X"7E",X"28",X"09",X"CB",X"BE",X"21",
		X"1C",X"86",X"36",X"22",X"18",X"66",X"CD",X"DA",X"11",X"18",X"61",X"FE",X"34",X"20",X"1A",X"21",
		X"22",X"98",X"36",X"15",X"21",X"DA",X"87",X"3A",X"00",X"84",X"CB",X"4F",X"28",X"03",X"21",X"D8",
		X"87",X"7E",X"FE",X"02",X"20",X"46",X"34",X"18",X"43",X"FE",X"20",X"20",X"07",X"21",X"22",X"98",
		X"36",X"16",X"18",X"38",X"FE",X"14",X"20",X"07",X"21",X"22",X"98",X"36",X"17",X"18",X"2D",X"A7",
		X"C2",X"27",X"0A",X"3A",X"57",X"86",X"CB",X"4F",X"C2",X"C7",X"0B",X"AF",X"32",X"80",X"98",X"32",
		X"81",X"98",X"21",X"22",X"98",X"36",X"32",X"21",X"A2",X"98",X"36",X"00",X"23",X"36",X"50",X"21",
		X"02",X"84",X"CB",X"C6",X"21",X"1C",X"86",X"36",X"3C",X"C3",X"27",X"0A",X"3A",X"AE",X"85",X"CB",
		X"4F",X"CA",X"27",X"0A",X"21",X"22",X"98",X"7E",X"C6",X"04",X"77",X"21",X"F4",X"98",X"06",X"0C",
		X"36",X"00",X"23",X"10",X"FB",X"C3",X"27",X"0A",X"21",X"1C",X"86",X"7E",X"A7",X"28",X"04",X"35",
		X"C3",X"27",X"0A",X"21",X"00",X"84",X"CB",X"4E",X"20",X"0C",X"3A",X"0A",X"84",X"A7",X"20",X"13",
		X"23",X"23",X"CB",X"CE",X"18",X"69",X"3A",X"0B",X"84",X"A7",X"20",X"51",X"23",X"23",X"CB",X"D6",
		X"C3",X"66",X"08",X"CB",X"46",X"20",X"21",X"21",X"00",X"84",X"CB",X"AE",X"CB",X"A6",X"23",X"7E",
		X"E6",X"57",X"77",X"23",X"7E",X"E6",X"E6",X"77",X"23",X"CB",X"96",X"CB",X"9E",X"23",X"CB",X"B6",
		X"21",X"46",X"86",X"36",X"00",X"C3",X"27",X"0A",X"23",X"23",X"CB",X"56",X"20",X"D9",X"21",X"00",
		X"84",X"32",X"30",X"68",X"CB",X"56",X"28",X"05",X"21",X"07",X"A0",X"36",X"01",X"21",X"00",X"84",
		X"CB",X"CE",X"CD",X"97",X"12",X"CD",X"A4",X"12",X"CD",X"B1",X"12",X"18",X"BA",X"21",X"02",X"84",
		X"CB",X"4E",X"20",X"B3",X"2B",X"2B",X"CB",X"8E",X"21",X"07",X"A0",X"36",X"00",X"18",X"E3",X"21",
		X"00",X"84",X"CB",X"46",X"CA",X"B0",X"08",X"23",X"23",X"CB",X"56",X"C2",X"B0",X"08",X"21",X"02",
		X"84",X"CB",X"5E",X"20",X"17",X"21",X"1D",X"86",X"36",X"78",X"CD",X"C9",X"12",X"21",X"02",X"84",
		X"CB",X"DE",X"21",X"CC",X"87",X"CB",X"CE",X"CB",X"D6",X"C3",X"27",X"0A",X"21",X"1D",X"86",X"7E",
		X"A7",X"28",X"04",X"35",X"C3",X"27",X"0A",X"21",X"CC",X"87",X"CB",X"96",X"CB",X"4E",X"C2",X"27",
		X"0A",X"CD",X"4B",X"13",X"18",X"88",X"21",X"02",X"84",X"CB",X"4E",X"20",X"43",X"21",X"02",X"84",
		X"CB",X"5E",X"20",X"17",X"21",X"1D",X"86",X"36",X"78",X"CD",X"D3",X"12",X"21",X"02",X"84",X"CB",
		X"DE",X"21",X"CC",X"87",X"CB",X"CE",X"CB",X"D6",X"C3",X"27",X"0A",X"21",X"1D",X"86",X"7E",X"A7",
		X"28",X"04",X"35",X"C3",X"27",X"0A",X"21",X"CC",X"87",X"CB",X"96",X"CB",X"4E",X"C2",X"27",X"0A",
		X"21",X"00",X"84",X"CB",X"8E",X"CD",X"4B",X"13",X"21",X"07",X"A0",X"36",X"00",X"C3",X"02",X"08",
		X"21",X"02",X"84",X"CB",X"66",X"20",X"1D",X"CB",X"E6",X"21",X"83",X"9A",X"CB",X"C6",X"21",X"1E",
		X"86",X"36",X"41",X"21",X"CC",X"87",X"CB",X"CE",X"CB",X"D6",X"AF",X"32",X"58",X"86",X"32",X"57",
		X"86",X"C3",X"27",X"0A",X"21",X"1E",X"86",X"7E",X"A7",X"28",X"1D",X"FE",X"38",X"20",X"0A",X"E5",
		X"21",X"83",X"9A",X"7E",X"E1",X"A7",X"C2",X"27",X"0A",X"E5",X"CD",X"CF",X"12",X"E1",X"35",X"CD",
		X"8D",X"18",X"CD",X"A7",X"18",X"C3",X"27",X"0A",X"21",X"CC",X"87",X"CB",X"96",X"CB",X"4E",X"C2",
		X"27",X"0A",X"CD",X"4B",X"13",X"21",X"00",X"84",X"7E",X"E6",X"01",X"77",X"23",X"06",X"06",X"36",
		X"00",X"23",X"10",X"FB",X"3E",X"90",X"32",X"76",X"86",X"21",X"46",X"86",X"36",X"00",X"3A",X"0D",
		X"84",X"32",X"A9",X"87",X"21",X"04",X"89",X"06",X"04",X"36",X"02",X"23",X"10",X"FB",X"21",X"04",
		X"89",X"11",X"00",X"70",X"01",X"04",X"00",X"3E",X"C1",X"CD",X"A1",X"00",X"21",X"87",X"87",X"36",
		X"00",X"21",X"07",X"A0",X"36",X"00",X"C3",X"27",X"0A",X"3A",X"F5",X"98",X"A7",X"C2",X"E6",X"09",
		X"3A",X"F7",X"98",X"A7",X"C2",X"E6",X"09",X"3A",X"22",X"98",X"FE",X"08",X"CA",X"E6",X"09",X"FE",
		X"09",X"CA",X"E6",X"09",X"FE",X"0C",X"CA",X"E6",X"09",X"FE",X"0D",X"CA",X"E6",X"09",X"3A",X"87",
		X"9A",X"A7",X"C2",X"E6",X"09",X"3A",X"57",X"86",X"CB",X"4F",X"20",X"14",X"21",X"2B",X"85",X"06",
		X"08",X"11",X"10",X"00",X"7E",X"FE",X"82",X"28",X"5D",X"FE",X"85",X"28",X"59",X"19",X"10",X"F4",
		X"21",X"28",X"85",X"06",X"08",X"11",X"10",X"00",X"CB",X"7E",X"28",X"4A",X"CB",X"B6",X"19",X"32",
		X"30",X"68",X"10",X"F4",X"3A",X"46",X"86",X"CB",X"47",X"20",X"3B",X"CD",X"8C",X"12",X"AF",X"32",
		X"A0",X"98",X"32",X"A1",X"98",X"CD",X"89",X"0F",X"21",X"46",X"86",X"36",X"00",X"21",X"88",X"9A",
		X"CB",X"C6",X"21",X"00",X"84",X"7E",X"E6",X"4F",X"77",X"23",X"CB",X"AE",X"CB",X"9E",X"2B",X"CB",
		X"4E",X"20",X"0C",X"21",X"0A",X"84",X"34",X"21",X"4A",X"86",X"36",X"00",X"C3",X"27",X"0A",X"21",
		X"0B",X"84",X"34",X"C3",X"27",X"0A",X"CD",X"A6",X"0B",X"CD",X"B1",X"0B",X"2A",X"D6",X"87",X"23",
		X"22",X"D6",X"87",X"CD",X"32",X"14",X"3A",X"57",X"86",X"CB",X"4F",X"20",X"06",X"3A",X"0D",X"84",
		X"32",X"05",X"9A",X"CD",X"00",X"1F",X"CD",X"25",X"14",X"3A",X"46",X"86",X"CB",X"47",X"28",X"05",
		X"CD",X"89",X"0F",X"18",X"08",X"CD",X"A2",X"0D",X"3E",X"FF",X"32",X"23",X"68",X"3A",X"46",X"86",
		X"CB",X"47",X"20",X"03",X"CD",X"4E",X"13",X"21",X"00",X"70",X"11",X"CE",X"87",X"01",X"02",X"00",
		X"3E",X"D2",X"CD",X"A1",X"00",X"32",X"30",X"68",X"3A",X"9A",X"87",X"A7",X"C2",X"71",X"0A",X"3A",
		X"57",X"86",X"CB",X"47",X"28",X"09",X"3A",X"58",X"86",X"E6",X"0F",X"FE",X"07",X"20",X"22",X"CD",
		X"0D",X"1D",X"21",X"25",X"98",X"06",X"0C",X"36",X"05",X"23",X"23",X"32",X"30",X"68",X"10",X"F7",
		X"3A",X"CC",X"87",X"CB",X"4F",X"C2",X"71",X"0A",X"CD",X"92",X"1B",X"CD",X"AF",X"1B",X"CD",X"E5",
		X"16",X"CB",X"C7",X"32",X"20",X"68",X"F1",X"C1",X"D1",X"E1",X"FD",X"E1",X"DD",X"E1",X"FB",X"C9",
		X"21",X"87",X"87",X"3A",X"57",X"86",X"CB",X"47",X"20",X"0C",X"3A",X"CF",X"87",X"CB",X"5F",X"20",
		X"05",X"CB",X"4E",X"CA",X"EC",X"1D",X"36",X"FF",X"21",X"57",X"86",X"CB",X"C6",X"CB",X"4E",X"CA",
		X"27",X"0A",X"CD",X"CA",X"0B",X"3A",X"58",X"86",X"FE",X"17",X"C2",X"27",X"0A",X"3A",X"76",X"86",
		X"FE",X"10",X"C2",X"FB",X"0A",X"AF",X"32",X"99",X"87",X"32",X"6C",X"89",X"32",X"F0",X"87",X"CD",
		X"22",X"0C",X"CD",X"15",X"0C",X"21",X"00",X"00",X"22",X"D6",X"87",X"21",X"9E",X"98",X"36",X"00",
		X"23",X"36",X"E0",X"CD",X"05",X"0C",X"21",X"23",X"84",X"36",X"FE",X"CD",X"6B",X"14",X"21",X"23",
		X"84",X"36",X"01",X"CD",X"6B",X"14",X"21",X"C0",X"83",X"06",X"3F",X"7E",X"FE",X"0C",X"20",X"02",
		X"36",X"8C",X"32",X"30",X"68",X"23",X"10",X"F3",X"C3",X"E0",X"04",X"FE",X"80",X"CA",X"54",X"06",
		X"C3",X"27",X"0A",X"21",X"87",X"87",X"3A",X"CF",X"87",X"CB",X"5F",X"20",X"05",X"CB",X"4E",X"CA",
		X"EC",X"1D",X"36",X"FF",X"CD",X"9B",X"19",X"21",X"F0",X"87",X"CB",X"9E",X"21",X"93",X"9A",X"36",
		X"00",X"21",X"57",X"86",X"CB",X"86",X"CB",X"4E",X"C2",X"71",X"0A",X"CD",X"CA",X"0B",X"3A",X"01",
		X"84",X"CB",X"4F",X"CA",X"5F",X"0B",X"CD",X"8D",X"18",X"CD",X"A7",X"18",X"CD",X"F2",X"0B",X"21",
		X"00",X"84",X"7E",X"E6",X"07",X"77",X"23",X"7E",X"E6",X"02",X"77",X"06",X"03",X"23",X"36",X"00",
		X"23",X"10",X"FB",X"CD",X"06",X"16",X"CD",X"DB",X"15",X"CD",X"90",X"16",X"C3",X"71",X"0A",X"CB",
		X"CF",X"32",X"01",X"84",X"21",X"80",X"98",X"DD",X"21",X"00",X"99",X"11",X"00",X"98",X"06",X"80",
		X"36",X"00",X"DD",X"36",X"00",X"00",X"32",X"30",X"68",X"3E",X"32",X"12",X"DD",X"23",X"13",X"23",
		X"10",X"EE",X"3E",X"FE",X"32",X"23",X"84",X"CD",X"6B",X"14",X"3E",X"01",X"32",X"23",X"84",X"CD",
		X"6B",X"14",X"CD",X"DF",X"0B",X"CD",X"97",X"15",X"CD",X"25",X"16",X"CD",X"40",X"16",X"21",X"03",
		X"A0",X"CB",X"C6",X"C3",X"71",X"0A",X"21",X"00",X"A0",X"06",X"04",X"36",X"00",X"23",X"10",X"FB",
		X"C9",X"11",X"07",X"A0",X"21",X"00",X"84",X"CB",X"4E",X"28",X"08",X"CB",X"56",X"28",X"04",X"EB",
		X"36",X"01",X"C9",X"EB",X"36",X"00",X"C9",X"C3",X"F8",X"08",X"CD",X"32",X"14",X"CD",X"4F",X"14",
		X"21",X"17",X"84",X"01",X"00",X"03",X"3A",X"00",X"84",X"E6",X"01",X"C2",X"5B",X"14",X"C9",X"21",
		X"C0",X"83",X"06",X"3F",X"7E",X"FE",X"8C",X"20",X"02",X"36",X"0C",X"32",X"30",X"68",X"23",X"10",
		X"F3",X"C9",X"21",X"00",X"98",X"11",X"80",X"98",X"06",X"80",X"32",X"30",X"68",X"AF",X"77",X"12",
		X"23",X"13",X"10",X"F6",X"C9",X"CD",X"39",X"1A",X"CD",X"94",X"1A",X"CD",X"73",X"1A",X"CD",X"C6",
		X"1A",X"CD",X"32",X"14",X"C9",X"CD",X"8D",X"18",X"CD",X"A7",X"18",X"CD",X"A3",X"19",X"CD",X"AC",
		X"18",X"C9",X"CD",X"AE",X"17",X"CD",X"3E",X"18",X"CD",X"45",X"18",X"CD",X"F8",X"17",X"CD",X"51",
		X"15",X"AF",X"32",X"A7",X"87",X"32",X"BF",X"87",X"32",X"9F",X"87",X"32",X"EB",X"87",X"32",X"DA",
		X"87",X"32",X"D8",X"87",X"21",X"00",X"00",X"22",X"ED",X"87",X"22",X"D4",X"87",X"22",X"D2",X"87",
		X"C9",X"DD",X"21",X"2A",X"86",X"21",X"AA",X"85",X"CD",X"6F",X"0C",X"DD",X"21",X"2D",X"86",X"21",
		X"AC",X"85",X"E5",X"CD",X"6F",X"0C",X"E1",X"DD",X"21",X"30",X"86",X"CD",X"6F",X"0C",X"C9",X"DD",
		X"36",X"00",X"00",X"7E",X"87",X"87",X"87",X"87",X"DD",X"77",X"01",X"23",X"7E",X"DD",X"77",X"02",
		X"C9",X"3A",X"00",X"84",X"CB",X"4F",X"20",X"05",X"21",X"16",X"84",X"18",X"03",X"21",X"19",X"84",
		X"7E",X"FE",X"90",X"D0",X"3A",X"57",X"86",X"CB",X"47",X"C0",X"3A",X"C0",X"87",X"A7",X"C8",X"21",
		X"00",X"84",X"CB",X"4E",X"20",X"1A",X"21",X"14",X"84",X"11",X"11",X"84",X"CD",X"54",X"0D",X"21",
		X"2D",X"86",X"11",X"33",X"86",X"CD",X"54",X"0D",X"21",X"02",X"84",X"22",X"F6",X"85",X"18",X"18",
		X"21",X"17",X"84",X"11",X"11",X"84",X"CD",X"54",X"0D",X"21",X"30",X"86",X"11",X"33",X"86",X"CD",
		X"54",X"0D",X"21",X"03",X"84",X"22",X"F6",X"85",X"CB",X"7E",X"20",X"20",X"21",X"11",X"84",X"11",
		X"2A",X"86",X"CD",X"60",X"0D",X"D8",X"2A",X"F6",X"85",X"CB",X"FE",X"21",X"87",X"9A",X"CB",X"C6",
		X"CD",X"6C",X"0D",X"3E",X"01",X"21",X"EA",X"89",X"CD",X"26",X"12",X"C9",X"21",X"11",X"84",X"3A",
		X"00",X"84",X"CB",X"4F",X"20",X"08",X"3A",X"BF",X"87",X"CB",X"47",X"C0",X"18",X"06",X"3A",X"BF",
		X"87",X"CB",X"4F",X"C0",X"3A",X"C0",X"87",X"FE",X"01",X"C8",X"11",X"33",X"86",X"CD",X"60",X"0D",
		X"D8",X"CD",X"6C",X"0D",X"21",X"87",X"9A",X"CB",X"C6",X"3E",X"01",X"21",X"EA",X"89",X"CD",X"26",
		X"12",X"DD",X"21",X"33",X"86",X"21",X"AC",X"85",X"CD",X"6F",X"0C",X"CD",X"84",X"0D",X"3A",X"C0",
		X"87",X"FE",X"02",X"C0",X"21",X"BF",X"87",X"3A",X"00",X"84",X"CB",X"4F",X"20",X"03",X"CB",X"C6",
		X"C9",X"CB",X"CE",X"C9",X"06",X"03",X"7E",X"12",X"23",X"13",X"32",X"30",X"68",X"10",X"F7",X"C9",
		X"06",X"03",X"EB",X"A7",X"1A",X"9E",X"23",X"13",X"10",X"FA",X"EB",X"C9",X"21",X"00",X"84",X"CB",
		X"4E",X"20",X"05",X"21",X"0A",X"84",X"18",X"03",X"21",X"0B",X"84",X"34",X"7E",X"32",X"0C",X"84",
		X"CD",X"45",X"18",X"C9",X"21",X"00",X"84",X"CB",X"4E",X"20",X"05",X"21",X"2D",X"86",X"18",X"03",
		X"21",X"30",X"86",X"11",X"33",X"86",X"06",X"03",X"A7",X"1A",X"8E",X"27",X"77",X"13",X"23",X"10",
		X"F8",X"C9",X"3A",X"01",X"84",X"CB",X"7F",X"20",X"51",X"3A",X"03",X"84",X"CB",X"57",X"C2",X"34",
		X"0E",X"21",X"01",X"84",X"CB",X"5E",X"20",X"36",X"3A",X"57",X"86",X"CB",X"4F",X"28",X"05",X"3A",
		X"70",X"89",X"18",X"03",X"3A",X"B0",X"85",X"CB",X"67",X"C0",X"21",X"01",X"84",X"CB",X"DE",X"3A",
		X"57",X"86",X"CB",X"4F",X"20",X"04",X"3E",X"32",X"18",X"02",X"3E",X"36",X"32",X"3E",X"86",X"CD",
		X"97",X"0F",X"AF",X"32",X"9E",X"87",X"21",X"8F",X"9A",X"36",X"01",X"C9",X"35",X"C9",X"21",X"3E",
		X"86",X"7E",X"FE",X"33",X"30",X"F6",X"FE",X"06",X"30",X"0E",X"CD",X"89",X"0F",X"21",X"01",X"84",
		X"CB",X"9E",X"21",X"3E",X"86",X"36",X"00",X"C9",X"22",X"42",X"86",X"3A",X"87",X"98",X"FE",X"08",
		X"38",X"E8",X"5F",X"3A",X"86",X"98",X"57",X"CD",X"16",X"1C",X"CD",X"3B",X"10",X"79",X"A7",X"28",
		X"D9",X"21",X"04",X"84",X"CB",X"B6",X"CD",X"09",X"12",X"3A",X"87",X"98",X"FE",X"F2",X"30",X"CA",
		X"CD",X"E0",X"10",X"C9",X"21",X"04",X"84",X"CB",X"76",X"C0",X"CB",X"56",X"20",X"1E",X"2B",X"CB",
		X"9E",X"3A",X"57",X"86",X"CB",X"4F",X"28",X"05",X"3A",X"70",X"89",X"18",X"03",X"3A",X"B0",X"85",
		X"CB",X"6F",X"20",X"03",X"23",X"CB",X"D6",X"AF",X"32",X"41",X"86",X"C9",X"21",X"41",X"86",X"34",
		X"7E",X"E6",X"1F",X"FE",X"09",X"30",X"06",X"21",X"03",X"84",X"CB",X"9E",X"C9",X"28",X"2B",X"FE",
		X"12",X"28",X"21",X"D8",X"FE",X"1F",X"20",X"04",X"AF",X"32",X"41",X"86",X"3A",X"57",X"86",X"CB",
		X"4F",X"28",X"05",X"3A",X"70",X"89",X"18",X"03",X"3A",X"B0",X"85",X"CB",X"6F",X"C8",X"21",X"04",
		X"84",X"CB",X"96",X"C9",X"21",X"03",X"84",X"CB",X"9E",X"C9",X"21",X"03",X"84",X"CB",X"DE",X"21",
		X"DF",X"32",X"3A",X"10",X"84",X"3D",X"5F",X"16",X"00",X"19",X"7E",X"2A",X"C8",X"87",X"11",X"0C",
		X"00",X"19",X"77",X"2A",X"C8",X"87",X"23",X"23",X"CB",X"6E",X"C2",X"CD",X"11",X"3E",X"01",X"32",
		X"90",X"9A",X"2B",X"2B",X"7E",X"87",X"D8",X"E6",X"38",X"20",X"03",X"CB",X"D6",X"C9",X"CB",X"56",
		X"28",X"09",X"CB",X"96",X"CB",X"DE",X"23",X"23",X"CB",X"E6",X"C9",X"CB",X"5E",X"28",X"09",X"CB",
		X"9E",X"CB",X"E6",X"23",X"23",X"CB",X"E6",X"C9",X"CB",X"66",X"C8",X"CB",X"A6",X"CB",X"B6",X"CB",
		X"EE",X"23",X"23",X"23",X"CB",X"FE",X"3E",X"01",X"32",X"8B",X"9A",X"21",X"04",X"84",X"CB",X"F6",
		X"2A",X"C8",X"87",X"11",X"0C",X"00",X"19",X"36",X"16",X"2A",X"C8",X"87",X"CB",X"46",X"C2",X"48",
		X"0F",X"CD",X"6C",X"12",X"F5",X"3C",X"6F",X"87",X"85",X"6F",X"CD",X"B5",X"2F",X"F1",X"CD",X"51",
		X"12",X"A7",X"20",X"0F",X"36",X"39",X"3E",X"0A",X"12",X"DD",X"36",X"00",X"00",X"21",X"F7",X"98",
		X"36",X"01",X"C9",X"3D",X"20",X"05",X"36",X"3A",X"C3",X"26",X"0F",X"3D",X"20",X"05",X"36",X"3B",
		X"C3",X"26",X"0F",X"36",X"3C",X"C3",X"26",X"0F",X"3A",X"10",X"84",X"FE",X"0A",X"30",X"04",X"3C",
		X"32",X"10",X"84",X"3A",X"AE",X"85",X"CB",X"4F",X"CA",X"11",X"0F",X"CD",X"6C",X"12",X"F5",X"6F",
		X"87",X"85",X"C6",X"0F",X"6F",X"CD",X"B5",X"2F",X"F1",X"CD",X"51",X"12",X"A7",X"20",X"05",X"36",
		X"3B",X"C3",X"26",X"0F",X"3D",X"20",X"05",X"36",X"3D",X"C3",X"26",X"0F",X"3D",X"20",X"05",X"36",
		X"3E",X"C3",X"26",X"0F",X"36",X"3F",X"C3",X"26",X"0F",X"21",X"82",X"98",X"06",X"08",X"36",X"00",
		X"23",X"32",X"30",X"68",X"10",X"F8",X"C9",X"21",X"08",X"84",X"CB",X"C6",X"11",X"02",X"98",X"DD",
		X"21",X"02",X"99",X"01",X"08",X"00",X"FD",X"21",X"82",X"98",X"3A",X"AE",X"85",X"32",X"E4",X"87",
		X"CB",X"4F",X"28",X"17",X"21",X"BB",X"0F",X"ED",X"B0",X"18",X"15",X"37",X"08",X"37",X"08",X"36",
		X"08",X"13",X"06",X"35",X"08",X"35",X"08",X"34",X"08",X"12",X"06",X"21",X"C3",X"0F",X"ED",X"B0",
		X"DD",X"E5",X"E1",X"3A",X"22",X"99",X"06",X"04",X"77",X"23",X"23",X"10",X"FB",X"FD",X"E5",X"E1",
		X"3A",X"A2",X"98",X"4F",X"3A",X"A3",X"98",X"06",X"04",X"71",X"23",X"77",X"23",X"10",X"FA",X"C9",
		X"21",X"82",X"98",X"FD",X"21",X"83",X"98",X"18",X"10",X"21",X"84",X"98",X"FD",X"21",X"85",X"98",
		X"18",X"07",X"21",X"86",X"98",X"FD",X"21",X"87",X"98",X"3A",X"06",X"98",X"FE",X"34",X"CA",X"1A",
		X"10",X"3A",X"06",X"99",X"E6",X"02",X"28",X"17",X"18",X"09",X"3A",X"06",X"99",X"E6",X"01",X"28",
		X"11",X"18",X"03",X"35",X"35",X"C9",X"FD",X"7E",X"00",X"3C",X"3C",X"FD",X"77",X"00",X"C9",X"34",
		X"34",X"C9",X"FD",X"7E",X"00",X"3D",X"3D",X"FD",X"77",X"00",X"C9",X"3A",X"E4",X"87",X"E6",X"07",
		X"28",X"11",X"FE",X"02",X"28",X"16",X"FE",X"04",X"28",X"1B",X"2A",X"02",X"86",X"ED",X"5B",X"06",
		X"86",X"18",X"5C",X"2A",X"02",X"86",X"ED",X"5B",X"04",X"86",X"18",X"10",X"2A",X"04",X"86",X"ED",
		X"5B",X"08",X"86",X"18",X"4A",X"2A",X"06",X"86",X"ED",X"5B",X"08",X"86",X"3A",X"3E",X"86",X"FE",
		X"2C",X"38",X"08",X"7E",X"FE",X"7F",X"20",X"0A",X"0E",X"00",X"C9",X"CD",X"92",X"10",X"79",X"FE",
		X"00",X"C8",X"EB",X"3A",X"3E",X"86",X"FE",X"2C",X"38",X"08",X"7E",X"FE",X"7F",X"20",X"1D",X"0E",
		X"00",X"C9",X"7E",X"FE",X"02",X"28",X"15",X"FE",X"03",X"28",X"11",X"FE",X"8D",X"28",X"0D",X"FE",
		X"7E",X"28",X"09",X"CB",X"BF",X"FE",X"0C",X"28",X"03",X"0E",X"00",X"C9",X"0E",X"01",X"C9",X"3A",
		X"3E",X"86",X"FE",X"2C",X"38",X"08",X"7E",X"FE",X"7F",X"20",X"0A",X"0E",X"00",X"C9",X"CD",X"D5",
		X"10",X"79",X"FE",X"00",X"C8",X"EB",X"3A",X"3E",X"86",X"FE",X"2C",X"38",X"08",X"7E",X"FE",X"7F",
		X"20",X"DA",X"0E",X"00",X"C9",X"7E",X"FE",X"08",X"28",X"D2",X"FE",X"09",X"28",X"CE",X"18",X"BB",
		X"21",X"25",X"85",X"22",X"F6",X"85",X"06",X"08",X"3A",X"E4",X"87",X"4F",X"DD",X"2A",X"F6",X"85",
		X"DD",X"CB",X"00",X"7E",X"20",X"32",X"DD",X"CB",X"03",X"7E",X"20",X"2C",X"2A",X"86",X"98",X"DD",
		X"5E",X"04",X"DD",X"56",X"05",X"DD",X"7E",X"06",X"FE",X"40",X"30",X"07",X"CD",X"77",X"11",X"30",
		X"17",X"18",X"22",X"3A",X"00",X"84",X"2F",X"E6",X"06",X"20",X"08",X"3E",X"10",X"85",X"6F",X"3E",
		X"10",X"84",X"67",X"CD",X"A1",X"11",X"38",X"0D",X"2A",X"F6",X"85",X"11",X"10",X"00",X"19",X"22",
		X"F6",X"85",X"10",X"B8",X"C9",X"78",X"32",X"9E",X"87",X"DD",X"22",X"C8",X"87",X"21",X"03",X"84",
		X"CB",X"D6",X"21",X"01",X"84",X"CB",X"9E",X"2A",X"F6",X"85",X"CB",X"B6",X"11",X"0C",X"00",X"19",
		X"22",X"F6",X"85",X"21",X"DF",X"32",X"3A",X"10",X"84",X"3D",X"5F",X"16",X"00",X"19",X"7E",X"DD",
		X"77",X"0C",X"21",X"03",X"84",X"CB",X"9E",X"CD",X"9F",X"0E",X"3A",X"03",X"84",X"CB",X"57",X"C8",
		X"CD",X"09",X"12",X"CD",X"09",X"12",X"C9",X"CB",X"49",X"20",X"13",X"7D",X"93",X"C6",X"08",X"FE",
		X"0C",X"D0",X"7C",X"92",X"CB",X"51",X"28",X"01",X"2F",X"D6",X"02",X"FE",X"0C",X"C9",X"7C",X"92",
		X"C6",X"08",X"FE",X"0C",X"D0",X"7D",X"93",X"CB",X"51",X"20",X"01",X"2F",X"D6",X"02",X"FE",X"0C",
		X"C9",X"CB",X"49",X"20",X"14",X"7D",X"93",X"C6",X"03",X"FE",X"12",X"D0",X"7C",X"92",X"CB",X"51",
		X"28",X"02",X"C6",X"10",X"D6",X"03",X"FE",X"12",X"C9",X"7C",X"92",X"C6",X"07",X"FE",X"12",X"D0",
		X"7D",X"93",X"CB",X"51",X"20",X"02",X"C6",X"10",X"D6",X"07",X"FE",X"12",X"C9",X"2A",X"03",X"84",
		X"CB",X"5E",X"C0",X"CB",X"96",X"2B",X"2B",X"CB",X"DE",X"C9",X"21",X"56",X"86",X"CB",X"DE",X"C9",
		X"21",X"24",X"98",X"06",X"0C",X"36",X"32",X"23",X"23",X"10",X"FA",X"C9",X"21",X"00",X"84",X"CB",
		X"4E",X"20",X"0B",X"21",X"0D",X"84",X"7E",X"23",X"23",X"77",X"23",X"77",X"18",X"08",X"21",X"0E",
		X"84",X"7E",X"23",X"77",X"23",X"77",X"C3",X"BD",X"19",X"2A",X"42",X"86",X"7E",X"A7",X"C8",X"35",
		X"35",X"7E",X"FE",X"22",X"D2",X"22",X"12",X"FE",X"12",X"D2",X"1F",X"12",X"CD",X"F0",X"0F",X"CD",
		X"F9",X"0F",X"CD",X"02",X"10",X"C9",X"A7",X"86",X"27",X"77",X"2B",X"7E",X"CE",X"00",X"27",X"77",
		X"C9",X"C5",X"F5",X"3A",X"00",X"84",X"CB",X"4F",X"28",X"14",X"CB",X"57",X"28",X"10",X"2A",X"F6",
		X"85",X"11",X"04",X"00",X"19",X"7E",X"C6",X"10",X"77",X"23",X"7E",X"C6",X"10",X"77",X"F1",X"C1",
		X"C9",X"DD",X"21",X"7E",X"99",X"21",X"7E",X"98",X"36",X"47",X"23",X"36",X"0A",X"DD",X"36",X"00",
		X"00",X"DD",X"21",X"76",X"99",X"21",X"76",X"98",X"11",X"77",X"98",X"C9",X"11",X"05",X"00",X"19",
		X"3A",X"00",X"84",X"CB",X"4F",X"28",X"09",X"CB",X"57",X"28",X"05",X"7E",X"D6",X"10",X"18",X"01",
		X"7E",X"FE",X"20",X"38",X"02",X"D6",X"08",X"07",X"07",X"E6",X"03",X"C9",X"21",X"80",X"9A",X"06",
		X"20",X"36",X"00",X"23",X"10",X"FB",X"C9",X"21",X"25",X"85",X"11",X"A5",X"84",X"01",X"80",X"00",
		X"CD",X"BE",X"12",X"C9",X"21",X"65",X"84",X"11",X"25",X"84",X"01",X"40",X"00",X"CD",X"BE",X"12",
		X"C9",X"21",X"40",X"80",X"11",X"00",X"90",X"01",X"80",X"03",X"CD",X"BE",X"12",X"C9",X"1A",X"ED",
		X"A0",X"2B",X"77",X"23",X"79",X"B0",X"20",X"F6",X"C9",X"CD",X"19",X"13",X"CD",X"33",X"13",X"CD",
		X"DC",X"12",X"C9",X"CD",X"19",X"13",X"CD",X"44",X"13",X"C3",X"CF",X"12",X"21",X"05",X"13",X"11",
		X"F0",X"98",X"01",X"08",X"00",X"C5",X"ED",X"B0",X"C1",X"21",X"FD",X"12",X"11",X"70",X"98",X"ED",
		X"B0",X"21",X"70",X"99",X"06",X"04",X"36",X"00",X"23",X"23",X"10",X"FA",X"C9",X"68",X"0C",X"71",
		X"0C",X"70",X"0C",X"6F",X"0C",X"91",X"98",X"81",X"98",X"69",X"98",X"59",X"98",X"79",X"70",X"69",
		X"70",X"59",X"70",X"68",X"0C",X"67",X"0C",X"66",X"0C",X"21",X"0D",X"13",X"11",X"FA",X"98",X"01",
		X"06",X"00",X"C5",X"ED",X"B0",X"C1",X"21",X"13",X"13",X"11",X"7A",X"98",X"ED",X"B0",X"21",X"78",
		X"99",X"18",X"C1",X"21",X"78",X"98",X"36",X"6A",X"23",X"36",X"0C",X"21",X"F8",X"98",X"36",X"89",
		X"23",X"36",X"70",X"C9",X"21",X"78",X"98",X"36",X"6B",X"18",X"ED",X"C3",X"D3",X"1C",X"21",X"29",
		X"85",X"11",X"10",X"00",X"06",X"08",X"22",X"F6",X"85",X"4E",X"3A",X"A2",X"98",X"B9",X"DA",X"64",
		X"13",X"91",X"18",X"05",X"D5",X"57",X"79",X"92",X"D1",X"32",X"1A",X"86",X"2A",X"F6",X"85",X"23",
		X"4E",X"3A",X"A3",X"98",X"B9",X"DA",X"7B",X"13",X"91",X"18",X"05",X"D5",X"57",X"79",X"92",X"D1",
		X"5F",X"16",X"00",X"3A",X"1A",X"86",X"6F",X"26",X"00",X"19",X"7C",X"A7",X"C2",X"FF",X"13",X"7D",
		X"FE",X"0A",X"D2",X"FF",X"13",X"2A",X"F6",X"85",X"2B",X"2B",X"2B",X"2B",X"7E",X"E6",X"BC",X"C2",
		X"FF",X"13",X"21",X"4A",X"86",X"CB",X"86",X"21",X"01",X"84",X"CB",X"7E",X"C0",X"CB",X"FE",X"23",
		X"CB",X"86",X"21",X"4A",X"86",X"CB",X"46",X"20",X"1F",X"2A",X"F6",X"85",X"2B",X"2B",X"2B",X"2B",
		X"CB",X"8E",X"CB",X"46",X"F5",X"11",X"06",X"00",X"19",X"F1",X"20",X"07",X"36",X"20",X"23",X"36",
		X"01",X"18",X"05",X"36",X"24",X"23",X"36",X"02",X"21",X"1C",X"86",X"36",X"A0",X"CD",X"8C",X"12",
		X"21",X"76",X"98",X"36",X"32",X"21",X"7E",X"98",X"36",X"32",X"3E",X"01",X"32",X"84",X"9A",X"21",
		X"22",X"98",X"3A",X"AE",X"85",X"CB",X"4F",X"28",X"03",X"36",X"4D",X"C9",X"36",X"4C",X"C9",X"2A",
		X"F6",X"85",X"11",X"10",X"00",X"19",X"05",X"C2",X"56",X"13",X"C9",X"21",X"00",X"84",X"CB",X"4E",
		X"20",X"07",X"3A",X"0A",X"84",X"32",X"0C",X"84",X"C9",X"3A",X"0B",X"84",X"32",X"0C",X"84",X"C9",
		X"AF",X"32",X"92",X"9A",X"C9",X"3A",X"46",X"86",X"CB",X"47",X"20",X"F4",X"3E",X"01",X"32",X"92",
		X"9A",X"C9",X"21",X"D4",X"83",X"DD",X"21",X"45",X"14",X"06",X"0A",X"DD",X"7E",X"00",X"77",X"2B",
		X"DD",X"23",X"10",X"F7",X"C9",X"A1",X"A2",X"A0",X"A1",X"7F",X"AC",X"9C",X"A8",X"AB",X"9E",X"21",
		X"DA",X"83",X"DD",X"21",X"65",X"14",X"06",X"03",X"C3",X"3B",X"14",X"21",X"C7",X"83",X"DD",X"21",
		X"68",X"14",X"C3",X"56",X"14",X"91",X"AE",X"A9",X"92",X"AE",X"A9",X"CD",X"32",X"14",X"CD",X"83",
		X"14",X"CD",X"DE",X"14",X"3A",X"00",X"84",X"CB",X"47",X"CA",X"7F",X"14",X"CD",X"F4",X"14",X"CD",
		X"E9",X"14",X"C9",X"3A",X"00",X"84",X"CB",X"47",X"C2",X"9C",X"14",X"CD",X"D8",X"14",X"3A",X"23",
		X"84",X"CB",X"6F",X"F5",X"C4",X"4F",X"14",X"F1",X"CC",X"B8",X"14",X"C9",X"CB",X"4F",X"C2",X"A7",
		X"14",X"CD",X"5B",X"14",X"C3",X"8E",X"14",X"CD",X"4F",X"14",X"3A",X"23",X"84",X"CB",X"6F",X"F5",
		X"C4",X"5B",X"14",X"F1",X"CC",X"D8",X"14",X"C9",X"21",X"DA",X"83",X"3A",X"CC",X"87",X"CB",X"4F",
		X"CA",X"D0",X"14",X"CB",X"57",X"C2",X"D0",X"14",X"3E",X"0C",X"77",X"2B",X"77",X"2B",X"77",X"C9",
		X"3E",X"8C",X"77",X"2B",X"77",X"2B",X"77",X"C9",X"21",X"C7",X"83",X"C3",X"BB",X"14",X"11",X"27",
		X"89",X"DD",X"21",X"F2",X"83",X"CD",X"FF",X"14",X"C9",X"11",X"14",X"84",X"DD",X"21",X"FC",X"83",
		X"CD",X"FF",X"14",X"C9",X"11",X"17",X"84",X"DD",X"21",X"E9",X"83",X"CD",X"FF",X"14",X"C9",X"21",
		X"1D",X"84",X"06",X"03",X"1A",X"E6",X"0F",X"77",X"23",X"1A",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",
		X"CB",X"3F",X"77",X"23",X"13",X"10",X"ED",X"21",X"22",X"84",X"06",X"04",X"7E",X"A7",X"20",X"18",
		X"3A",X"CC",X"87",X"CB",X"4F",X"CA",X"32",X"15",X"CB",X"57",X"C2",X"32",X"15",X"3E",X"0C",X"C3",
		X"34",X"15",X"3E",X"8C",X"77",X"2B",X"10",X"E4",X"21",X"22",X"84",X"06",X"06",X"7E",X"FE",X"8C",
		X"28",X"06",X"FE",X"0C",X"28",X"02",X"C6",X"10",X"DD",X"77",X"00",X"2B",X"DD",X"2B",X"10",X"ED",
		X"C9",X"21",X"A4",X"98",X"06",X"0C",X"36",X"00",X"23",X"36",X"50",X"23",X"10",X"F8",X"C9",X"DD",
		X"4E",X"00",X"3A",X"A2",X"98",X"B9",X"DA",X"6C",X"15",X"91",X"18",X"03",X"57",X"79",X"92",X"FE",
		X"0B",X"D0",X"FD",X"4E",X"00",X"3A",X"A3",X"98",X"B9",X"DA",X"7F",X"15",X"91",X"18",X"03",X"57",
		X"79",X"92",X"FE",X"0B",X"D0",X"2A",X"F6",X"85",X"11",X"04",X"00",X"19",X"22",X"F6",X"85",X"21",
		X"4A",X"86",X"CB",X"C6",X"C3",X"A7",X"13",X"F5",X"21",X"00",X"80",X"01",X"C0",X"03",X"CD",X"BF",
		X"15",X"CD",X"EC",X"11",X"F1",X"C9",X"F5",X"21",X"40",X"80",X"01",X"80",X"03",X"CD",X"BF",X"15",
		X"21",X"C0",X"83",X"06",X"3F",X"36",X"7F",X"32",X"30",X"68",X"23",X"10",X"F8",X"F1",X"C9",X"36",
		X"7F",X"32",X"30",X"68",X"23",X"0B",X"79",X"B0",X"20",X"F5",X"C9",X"F5",X"11",X"20",X"00",X"DD",
		X"7E",X"00",X"77",X"DD",X"23",X"19",X"F1",X"3D",X"20",X"F1",X"C9",X"F5",X"21",X"62",X"30",X"11",
		X"16",X"80",X"01",X"06",X"00",X"ED",X"B0",X"3A",X"A5",X"85",X"47",X"E6",X"0F",X"C6",X"10",X"32",
		X"13",X"80",X"78",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"28",X"04",X"C6",X"10",X"18",X"02",X"3E",
		X"7F",X"32",X"14",X"80",X"F1",X"C9",X"21",X"2D",X"81",X"11",X"20",X"00",X"3A",X"A5",X"85",X"FE",
		X"01",X"20",X"0A",X"DD",X"21",X"6F",X"30",X"3E",X"0D",X"CD",X"CB",X"15",X"C9",X"DD",X"21",X"7C",
		X"30",X"3E",X"0E",X"18",X"F4",X"F5",X"21",X"FA",X"80",X"11",X"20",X"00",X"DD",X"21",X"8A",X"30",
		X"3E",X"11",X"CD",X"CB",X"15",X"21",X"9C",X"81",X"DD",X"21",X"9B",X"30",X"3E",X"08",X"18",X"4B",
		X"F5",X"21",X"EA",X"80",X"11",X"20",X"00",X"DD",X"21",X"A3",X"30",X"3E",X"11",X"CD",X"CB",X"15",
		X"3A",X"C0",X"87",X"A7",X"20",X"02",X"F1",X"C9",X"21",X"B1",X"80",X"DD",X"21",X"B4",X"30",X"3E",
		X"14",X"CD",X"CB",X"15",X"3A",X"C0",X"87",X"FE",X"01",X"20",X"02",X"F1",X"C9",X"21",X"B4",X"80",
		X"DD",X"21",X"C8",X"30",X"3E",X"14",X"CD",X"CB",X"15",X"3A",X"C0",X"87",X"FE",X"02",X"20",X"02",
		X"F1",X"C9",X"21",X"B7",X"80",X"DD",X"21",X"DC",X"30",X"3E",X"14",X"CD",X"CB",X"15",X"F1",X"C9",
		X"F5",X"3A",X"C0",X"87",X"A7",X"20",X"02",X"F1",X"C9",X"11",X"20",X"00",X"21",X"B1",X"81",X"01",
		X"AA",X"85",X"0A",X"C6",X"50",X"77",X"03",X"19",X"0A",X"A7",X"28",X"05",X"C6",X"50",X"77",X"18",
		X"02",X"36",X"7F",X"3A",X"C0",X"87",X"FE",X"01",X"20",X"02",X"F1",X"C9",X"21",X"B4",X"81",X"CD",
		X"D3",X"16",X"3A",X"C0",X"87",X"FE",X"02",X"20",X"02",X"F1",X"C9",X"21",X"B7",X"81",X"CD",X"D3",
		X"16",X"F1",X"C9",X"01",X"AC",X"85",X"11",X"20",X"00",X"0A",X"C6",X"50",X"77",X"03",X"19",X"DD",
		X"19",X"0A",X"C6",X"50",X"77",X"21",X"32",X"85",X"11",X"64",X"99",X"06",X"08",X"7E",X"12",X"13",
		X"13",X"D5",X"11",X"10",X"00",X"19",X"D1",X"10",X"F4",X"C9",X"3A",X"00",X"84",X"CB",X"4F",X"20",
		X"05",X"21",X"0D",X"84",X"18",X"03",X"21",X"0E",X"84",X"7E",X"21",X"E8",X"87",X"FE",X"12",X"DA",
		X"14",X"17",X"3E",X"12",X"77",X"D6",X"01",X"87",X"87",X"5F",X"16",X"00",X"21",X"34",X"17",X"19",
		X"7E",X"32",X"1E",X"98",X"23",X"7E",X"32",X"1F",X"98",X"23",X"7E",X"32",X"E7",X"87",X"23",X"7E",
		X"32",X"E6",X"87",X"C9",X"52",X"0D",X"04",X"5D",X"53",X"0E",X"06",X"5E",X"54",X"0F",X"08",X"5F",
		X"55",X"10",X"10",X"60",X"55",X"10",X"10",X"60",X"56",X"10",X"20",X"4E",X"56",X"10",X"20",X"4E",
		X"57",X"11",X"30",X"4F",X"57",X"11",X"30",X"4F",X"58",X"12",X"40",X"61",X"58",X"12",X"40",X"61",
		X"59",X"13",X"50",X"50",X"59",X"13",X"50",X"50",X"5A",X"14",X"60",X"62",X"5A",X"14",X"60",X"62",
		X"5B",X"15",X"70",X"51",X"5B",X"15",X"70",X"51",X"5C",X"16",X"80",X"63",X"21",X"00",X"90",X"7D",
		X"E6",X"1F",X"FE",X"03",X"DA",X"A2",X"17",X"36",X"7F",X"23",X"32",X"30",X"68",X"7D",X"FE",X"80",
		X"20",X"ED",X"7C",X"FE",X"93",X"20",X"E8",X"3E",X"8F",X"32",X"01",X"90",X"3E",X"8E",X"32",X"61",
		X"93",X"C9",X"FE",X"01",X"20",X"04",X"36",X"8D",X"18",X"DF",X"36",X"7E",X"18",X"DB",X"21",X"40",
		X"80",X"7D",X"E6",X"1F",X"FE",X"03",X"DA",X"E1",X"17",X"36",X"7F",X"23",X"32",X"30",X"68",X"7D",
		X"FE",X"C0",X"20",X"ED",X"7C",X"FE",X"83",X"20",X"E8",X"3E",X"8F",X"32",X"41",X"80",X"36",X"8E",
		X"32",X"A1",X"83",X"21",X"00",X"80",X"06",X"40",X"32",X"30",X"68",X"36",X"0C",X"23",X"10",X"F8",
		X"C9",X"FE",X"01",X"20",X"04",X"36",X"8D",X"18",X"D2",X"36",X"7E",X"18",X"CE",X"21",X"11",X"84",
		X"06",X"09",X"36",X"00",X"23",X"10",X"FB",X"C9",X"3A",X"CF",X"87",X"CB",X"5F",X"20",X"1F",X"3A",
		X"87",X"87",X"CB",X"4F",X"20",X"18",X"21",X"0D",X"84",X"7E",X"FE",X"00",X"28",X"01",X"35",X"4E",
		X"23",X"7E",X"FE",X"00",X"20",X"02",X"36",X"01",X"23",X"71",X"23",X"71",X"18",X"0F",X"21",X"0D",
		X"84",X"06",X"04",X"36",X"00",X"23",X"10",X"FB",X"3E",X"01",X"32",X"0E",X"84",X"3A",X"57",X"86",
		X"CB",X"4F",X"C8",X"06",X"04",X"21",X"0D",X"84",X"36",X"02",X"23",X"10",X"FB",X"C9",X"21",X"09",
		X"84",X"7E",X"C3",X"64",X"19",X"21",X"0C",X"80",X"11",X"2C",X"80",X"06",X"14",X"3E",X"0C",X"77",
		X"32",X"30",X"68",X"12",X"23",X"13",X"10",X"F5",X"3A",X"0C",X"84",X"FE",X"00",X"C8",X"FE",X"0A",
		X"38",X"02",X"3E",X"09",X"47",X"21",X"1D",X"80",X"E5",X"CD",X"72",X"18",X"E1",X"2B",X"2B",X"10",
		X"F7",X"C9",X"11",X"20",X"00",X"3E",X"7F",X"77",X"2B",X"77",X"19",X"77",X"23",X"77",X"C9",X"21",
		X"A5",X"84",X"06",X"80",X"36",X"00",X"23",X"32",X"30",X"68",X"10",X"F8",X"C9",X"21",X"25",X"85",
		X"18",X"F0",X"21",X"25",X"84",X"06",X"08",X"3E",X"00",X"77",X"23",X"36",X"90",X"CD",X"64",X"19",
		X"CD",X"64",X"19",X"23",X"10",X"F1",X"C9",X"21",X"65",X"84",X"18",X"E9",X"21",X"68",X"31",X"CD",
		X"DE",X"1B",X"4F",X"87",X"87",X"87",X"87",X"5F",X"16",X"00",X"19",X"06",X"08",X"E5",X"5E",X"23",
		X"56",X"7A",X"A7",X"28",X"04",X"EB",X"CD",X"28",X"19",X"E1",X"23",X"23",X"32",X"30",X"68",X"10",
		X"EC",X"21",X"D0",X"81",X"3E",X"02",X"4F",X"AF",X"CD",X"28",X"19",X"3A",X"57",X"86",X"CB",X"4F",
		X"20",X"12",X"21",X"85",X"87",X"3A",X"00",X"84",X"CB",X"4F",X"20",X"05",X"CB",X"46",X"C8",X"18",
		X"03",X"CB",X"4E",X"C8",X"21",X"0A",X"19",X"11",X"02",X"82",X"01",X"0F",X"00",X"C5",X"ED",X"B0",
		X"C1",X"21",X"19",X"19",X"11",X"22",X"82",X"ED",X"B0",X"C9",X"8C",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"0C",X"8C",X"03",X"03",X"03",X"03",X"03",X"03",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"0C",X"C5",X"78",X"FE",X"05",X"DA",X"6B",X"19",X"E5",
		X"36",X"00",X"3E",X"02",X"CD",X"64",X"19",X"79",X"FE",X"00",X"20",X"05",X"3E",X"02",X"CD",X"62",
		X"19",X"23",X"36",X"02",X"23",X"36",X"04",X"E1",X"11",X"20",X"00",X"19",X"36",X"01",X"3E",X"03",
		X"CD",X"62",X"19",X"79",X"FE",X"00",X"20",X"05",X"3E",X"03",X"CD",X"62",X"19",X"23",X"36",X"05",
		X"C1",X"C9",X"23",X"77",X"23",X"77",X"23",X"77",X"23",X"77",X"C9",X"11",X"20",X"00",X"36",X"0A",
		X"23",X"36",X"0B",X"2B",X"79",X"FE",X"00",X"20",X"06",X"CD",X"93",X"19",X"CD",X"93",X"19",X"CD",
		X"93",X"19",X"CD",X"93",X"19",X"CD",X"93",X"19",X"CD",X"93",X"19",X"19",X"36",X"06",X"23",X"36",
		X"07",X"C1",X"C9",X"19",X"36",X"08",X"23",X"36",X"09",X"2B",X"C9",X"21",X"05",X"9A",X"7E",X"23",
		X"77",X"18",X"22",X"21",X"00",X"84",X"CB",X"4E",X"20",X"0C",X"21",X"0D",X"84",X"34",X"7E",X"23",
		X"23",X"77",X"23",X"77",X"18",X"07",X"21",X"0E",X"84",X"34",X"7E",X"18",X"F3",X"3A",X"57",X"86",
		X"CB",X"4F",X"20",X"D7",X"2B",X"CD",X"21",X"1A",X"7E",X"E6",X"0F",X"C6",X"10",X"32",X"23",X"80",
		X"7E",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"28",X"07",X"C6",X"10",X"32",X"24",X"80",X"18",X"05",
		X"3E",X"7F",X"32",X"24",X"80",X"21",X"08",X"80",X"06",X"07",X"DD",X"21",X"68",X"30",X"DD",X"7E",
		X"00",X"77",X"2B",X"DD",X"23",X"10",X"F7",X"21",X"00",X"84",X"CB",X"4E",X"20",X"0B",X"21",X"0D",
		X"84",X"7E",X"23",X"23",X"77",X"23",X"77",X"18",X"08",X"21",X"0E",X"84",X"7E",X"23",X"77",X"23",
		X"77",X"21",X"0F",X"84",X"7E",X"32",X"27",X"86",X"FE",X"0F",X"D8",X"3E",X"0F",X"77",X"23",X"77",
		X"C9",X"11",X"01",X"00",X"7E",X"A7",X"28",X"0F",X"1F",X"47",X"30",X"04",X"7A",X"83",X"27",X"57",
		X"7B",X"87",X"27",X"5F",X"78",X"18",X"EE",X"72",X"C9",X"21",X"58",X"32",X"CD",X"DE",X"1B",X"87",
		X"87",X"87",X"5F",X"16",X"00",X"19",X"11",X"10",X"00",X"E5",X"DD",X"E1",X"21",X"29",X"85",X"06",
		X"08",X"E5",X"DD",X"7E",X"00",X"4F",X"A7",X"28",X"10",X"79",X"87",X"87",X"87",X"87",X"3C",X"77",
		X"23",X"79",X"DD",X"23",X"E6",X"F0",X"77",X"18",X"05",X"DD",X"23",X"2B",X"CB",X"FE",X"E1",X"19",
		X"10",X"DF",X"C9",X"11",X"10",X"00",X"21",X"28",X"85",X"06",X"08",X"E5",X"CB",X"7E",X"28",X"06",
		X"23",X"36",X"00",X"23",X"36",X"00",X"E1",X"E5",X"2B",X"2B",X"2B",X"7E",X"E6",X"01",X"77",X"E1",
		X"19",X"10",X"E8",X"C9",X"21",X"2B",X"85",X"11",X"10",X"00",X"06",X"08",X"E5",X"78",X"FE",X"05",
		X"38",X"07",X"36",X"20",X"23",X"36",X"01",X"18",X"15",X"22",X"F6",X"85",X"E1",X"E5",X"2B",X"2B",
		X"2B",X"2B",X"2B",X"2B",X"CB",X"C6",X"2A",X"F6",X"85",X"36",X"24",X"23",X"36",X"02",X"23",X"36",
		X"00",X"E1",X"19",X"10",X"D7",X"C9",X"21",X"F0",X"30",X"CD",X"DE",X"1B",X"87",X"87",X"87",X"5F",
		X"16",X"00",X"19",X"E5",X"DD",X"E1",X"21",X"67",X"84",X"11",X"08",X"00",X"06",X"08",X"FD",X"21",
		X"65",X"84",X"FD",X"E5",X"CB",X"46",X"28",X"10",X"36",X"FF",X"FD",X"36",X"00",X"00",X"FD",X"23",
		X"FD",X"36",X"00",X"60",X"DD",X"23",X"18",X"1A",X"DD",X"7E",X"00",X"A7",X"28",X"EA",X"87",X"87",
		X"87",X"87",X"3C",X"FD",X"77",X"00",X"FD",X"23",X"DD",X"7E",X"00",X"E6",X"F0",X"FD",X"77",X"00",
		X"DD",X"23",X"FD",X"E1",X"FD",X"19",X"19",X"10",X"C9",X"21",X"3C",X"98",X"11",X"3C",X"99",X"06",
		X"08",X"36",X"1E",X"23",X"36",X"04",X"23",X"AF",X"12",X"13",X"13",X"10",X"F4",X"C9",X"3E",X"02",
		X"32",X"22",X"98",X"AF",X"32",X"23",X"98",X"32",X"80",X"98",X"32",X"81",X"98",X"3E",X"38",X"32",
		X"00",X"98",X"3E",X"06",X"32",X"01",X"98",X"3A",X"57",X"86",X"CB",X"4F",X"20",X"1F",X"21",X"85",
		X"87",X"3A",X"00",X"84",X"CB",X"4F",X"20",X"06",X"CB",X"46",X"20",X"11",X"18",X"04",X"CB",X"4E",
		X"20",X"0B",X"3E",X"08",X"32",X"A3",X"98",X"3E",X"B1",X"32",X"A2",X"98",X"C9",X"3E",X"71",X"32",
		X"A2",X"98",X"3E",X"80",X"32",X"A3",X"98",X"21",X"01",X"84",X"CB",X"E6",X"C9",X"21",X"00",X"84",
		X"CB",X"4E",X"20",X"05",X"21",X"0A",X"84",X"18",X"03",X"21",X"0B",X"84",X"35",X"7E",X"32",X"0C",
		X"84",X"C9",X"21",X"65",X"84",X"11",X"07",X"00",X"06",X"08",X"DD",X"21",X"BC",X"98",X"7E",X"DD",
		X"77",X"00",X"23",X"DD",X"23",X"7E",X"DD",X"77",X"00",X"DD",X"23",X"19",X"10",X"F0",X"C9",X"21",
		X"29",X"85",X"06",X"08",X"11",X"0D",X"00",X"DD",X"21",X"64",X"98",X"FD",X"21",X"E4",X"98",X"7E",
		X"FD",X"77",X"00",X"FD",X"23",X"23",X"7E",X"FD",X"77",X"00",X"23",X"FD",X"23",X"7E",X"DD",X"77",
		X"00",X"23",X"DD",X"23",X"7E",X"DD",X"77",X"00",X"DD",X"23",X"19",X"10",X"E2",X"C9",X"3A",X"27",
		X"86",X"FE",X"10",X"38",X"04",X"E6",X"03",X"C6",X"0C",X"3D",X"C9",X"06",X"00",X"2A",X"D6",X"85",
		X"CD",X"8E",X"1C",X"2A",X"D8",X"85",X"CD",X"8E",X"1C",X"2A",X"DA",X"85",X"CD",X"8E",X"1C",X"2A",
		X"DC",X"85",X"CD",X"8E",X"1C",X"78",X"21",X"01",X"84",X"CB",X"A6",X"A7",X"C0",X"CB",X"E6",X"C9",
		X"DD",X"21",X"FA",X"85",X"18",X"23",X"DD",X"21",X"02",X"86",X"18",X"1D",X"DD",X"21",X"0A",X"86",
		X"18",X"17",X"3A",X"AE",X"85",X"E6",X"0F",X"28",X"0C",X"FE",X"06",X"28",X"08",X"3E",X"06",X"82",
		X"57",X"3E",X"06",X"83",X"5F",X"DD",X"21",X"D6",X"85",X"CD",X"5A",X"1C",X"DD",X"75",X"00",X"DD",
		X"74",X"01",X"CD",X"87",X"1C",X"DD",X"73",X"02",X"DD",X"72",X"03",X"23",X"DD",X"75",X"04",X"DD",
		X"74",X"05",X"13",X"DD",X"73",X"06",X"DD",X"72",X"07",X"C9",X"7A",X"D6",X"11",X"CB",X"3F",X"CB",
		X"3F",X"57",X"CB",X"3F",X"87",X"87",X"87",X"87",X"87",X"6F",X"7A",X"CB",X"3F",X"CB",X"3F",X"CB",
		X"3F",X"CB",X"3F",X"67",X"16",X"00",X"CB",X"3B",X"CB",X"3B",X"CB",X"3B",X"A7",X"ED",X"52",X"EB",
		X"21",X"A0",X"83",X"A7",X"ED",X"52",X"C9",X"11",X"E0",X"FF",X"EB",X"19",X"EB",X"C9",X"7E",X"FE",
		X"7F",X"C0",X"04",X"C9",X"CD",X"19",X"13",X"3A",X"00",X"84",X"CB",X"4F",X"20",X"05",X"CD",X"33",
		X"13",X"18",X"03",X"CD",X"44",X"13",X"21",X"C7",X"1C",X"11",X"DE",X"98",X"01",X"06",X"00",X"C5",
		X"ED",X"B0",X"C1",X"21",X"CD",X"1C",X"11",X"5E",X"98",X"ED",X"B0",X"21",X"5E",X"99",X"06",X"03",
		X"36",X"00",X"23",X"23",X"10",X"FA",X"C9",X"81",X"98",X"71",X"98",X"61",X"98",X"6E",X"0C",X"6D",
		X"0C",X"6C",X"0C",X"21",X"F0",X"98",X"06",X"10",X"36",X"00",X"23",X"10",X"FB",X"21",X"70",X"98",
		X"06",X"10",X"36",X"00",X"23",X"10",X"FB",X"21",X"5E",X"98",X"11",X"DE",X"98",X"06",X"06",X"3E",
		X"00",X"77",X"12",X"23",X"13",X"10",X"F8",X"C9",X"E5",X"D5",X"F5",X"2A",X"F4",X"85",X"ED",X"5B",
		X"F4",X"85",X"29",X"29",X"19",X"23",X"22",X"F4",X"85",X"F1",X"D1",X"E1",X"C9",X"DD",X"E5",X"FD",
		X"E5",X"E5",X"D5",X"C5",X"F5",X"21",X"56",X"86",X"CB",X"56",X"28",X"1C",X"CB",X"96",X"21",X"48",
		X"86",X"3A",X"A3",X"98",X"FE",X"18",X"D2",X"2D",X"1D",X"36",X"00",X"18",X"0B",X"34",X"7E",X"FE",
		X"02",X"20",X"05",X"36",X"00",X"CD",X"B3",X"2F",X"F1",X"C1",X"D1",X"E1",X"FD",X"E1",X"DD",X"E1",
		X"C9",X"3A",X"A2",X"98",X"57",X"3A",X"A3",X"98",X"5F",X"3A",X"AF",X"85",X"C3",X"25",X"1C",X"27",
		X"28",X"2D",X"2D",X"2E",X"1B",X"0C",X"29",X"26",X"2E",X"29",X"0C",X"1D",X"25",X"28",X"21",X"0C",
		X"1D",X"27",X"1A",X"0C",X"21",X"2C",X"2E",X"29",X"5E",X"66",X"62",X"6D",X"35",X"10",X"0C",X"2C",
		X"2B",X"1E",X"2D",X"27",X"1E",X"0C",X"2D",X"27",X"2E",X"28",X"1C",X"0C",X"1E",X"26",X"22",X"2D",
		X"27",X"28",X"2D",X"2D",X"2E",X"1B",X"0C",X"2D",X"2B",X"1A",X"2D",X"2C",X"0C",X"21",X"2C",X"2E",
		X"29",X"0C",X"27",X"1E",X"21",X"2D",X"1E",X"2B",X"28",X"1F",X"1E",X"1B",X"0C",X"9E",X"A6",X"9A",
		X"A0",X"0C",X"9E",X"AE",X"A7",X"A2",X"AD",X"A7",X"A8",X"9C",X"0C",X"A8",X"AD",X"0C",X"0C",X"0C",
		X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",
		X"0C",X"0C",X"1D",X"27",X"1A",X"0C",X"27",X"22",X"28",X"1C",X"0C",X"2D",X"2B",X"1E",X"2C",X"27",
		X"22",X"6C",X"6B",X"5E",X"72",X"5A",X"65",X"69",X"0C",X"52",X"0C",X"6B",X"68",X"0C",X"51",X"72",
		X"65",X"67",X"68",X"0C",X"6B",X"5E",X"72",X"5A",X"65",X"69",X"0C",X"51",X"CB",X"56",X"C2",X"17",
		X"1E",X"CB",X"D6",X"26",X"17",X"2E",X"3A",X"22",X"89",X"87",X"3E",X"01",X"32",X"03",X"A0",X"CD",
		X"8D",X"18",X"CD",X"A7",X"18",X"CD",X"F2",X"0B",X"CD",X"97",X"15",X"CD",X"6B",X"14",X"CD",X"CA",
		X"0B",X"CD",X"DF",X"0B",X"C3",X"71",X"0A",X"CD",X"DB",X"15",X"2A",X"89",X"87",X"2C",X"7D",X"FE",
		X"3C",X"20",X"2D",X"2E",X"00",X"A7",X"25",X"7C",X"FE",X"0F",X"20",X"02",X"26",X"09",X"7C",X"FE",
		X"40",X"38",X"08",X"21",X"87",X"87",X"CB",X"CE",X"C3",X"71",X"0A",X"E6",X"0F",X"C6",X"50",X"32",
		X"D7",X"81",X"7C",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"C6",X"50",X"32",X"F7",X"81",
		X"22",X"89",X"87",X"3E",X"04",X"21",X"57",X"82",X"DD",X"21",X"68",X"1D",X"CD",X"CB",X"15",X"3E",
		X"14",X"21",X"D4",X"80",X"DD",X"21",X"6C",X"1D",X"CD",X"CB",X"15",X"3E",X"06",X"21",X"92",X"82",
		X"DD",X"21",X"96",X"1D",X"CD",X"CB",X"15",X"3E",X"16",X"21",X"CE",X"80",X"DD",X"21",X"80",X"1D",
		X"CD",X"CB",X"15",X"3E",X"19",X"21",X"6C",X"80",X"DD",X"21",X"4F",X"1D",X"CD",X"CB",X"15",X"2A",
		X"89",X"87",X"7D",X"FE",X"1E",X"30",X"06",X"DD",X"21",X"AF",X"1D",X"18",X"04",X"DD",X"21",X"9C",
		X"1D",X"21",X"E6",X"80",X"3E",X"13",X"CD",X"CB",X"15",X"3A",X"A5",X"85",X"FE",X"00",X"20",X"06",
		X"CD",X"CC",X"1E",X"C3",X"71",X"0A",X"FE",X"01",X"20",X"09",X"CD",X"CC",X"1E",X"CD",X"D9",X"1E",
		X"C3",X"71",X"0A",X"CD",X"E6",X"1E",X"CD",X"F3",X"1E",X"C3",X"71",X"0A",X"3E",X"0F",X"21",X"2A",
		X"81",X"DD",X"21",X"C2",X"1D",X"CD",X"CB",X"15",X"C9",X"3E",X"0D",X"21",X"30",X"81",X"DD",X"21",
		X"DF",X"1D",X"CD",X"CB",X"15",X"C9",X"3E",X"0E",X"21",X"10",X"81",X"DD",X"21",X"D1",X"1D",X"CD",
		X"CB",X"15",X"C9",X"21",X"2A",X"81",X"3E",X"0F",X"DD",X"21",X"AF",X"1D",X"CD",X"CB",X"15",X"C9",
		X"2A",X"23",X"84",X"7D",X"E6",X"03",X"FE",X"03",X"28",X"10",X"FE",X"02",X"28",X"1A",X"FE",X"01",
		X"28",X"24",X"21",X"6D",X"84",X"CD",X"75",X"1F",X"18",X"24",X"21",X"75",X"84",X"CD",X"75",X"1F",
		X"21",X"7D",X"84",X"CD",X"75",X"1F",X"18",X"1B",X"21",X"85",X"84",X"CD",X"75",X"1F",X"21",X"8D",
		X"84",X"CD",X"75",X"1F",X"18",X"08",X"21",X"95",X"84",X"CD",X"75",X"1F",X"18",X"05",X"21",X"25",
		X"85",X"18",X"03",X"21",X"65",X"85",X"11",X"10",X"00",X"06",X"04",X"78",X"32",X"29",X"86",X"C5",
		X"D5",X"E5",X"A7",X"11",X"25",X"85",X"ED",X"52",X"7D",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",
		X"3F",X"4F",X"3E",X"08",X"A7",X"91",X"32",X"9D",X"87",X"E1",X"E5",X"CD",X"39",X"23",X"E1",X"D1",
		X"C1",X"19",X"10",X"D7",X"C9",X"E5",X"23",X"23",X"CB",X"66",X"20",X"07",X"CB",X"7E",X"C2",X"BC",
		X"21",X"18",X"02",X"E1",X"C9",X"E1",X"E5",X"56",X"7A",X"A7",X"28",X"54",X"23",X"5E",X"7B",X"FE",
		X"F0",X"30",X"4D",X"CD",X"CB",X"22",X"2A",X"EA",X"85",X"7E",X"FE",X"09",X"28",X"1E",X"FE",X"08",
		X"28",X"1A",X"FE",X"0C",X"28",X"16",X"FE",X"03",X"28",X"12",X"FE",X"01",X"28",X"0E",X"FE",X"05",
		X"28",X"0A",X"FE",X"06",X"28",X"06",X"FE",X"07",X"28",X"02",X"20",X"24",X"2A",X"EC",X"85",X"7E",
		X"FE",X"09",X"28",X"24",X"FE",X"08",X"28",X"20",X"FE",X"0C",X"28",X"1C",X"FE",X"02",X"28",X"18",
		X"FE",X"00",X"28",X"14",X"FE",X"04",X"28",X"10",X"FE",X"0A",X"28",X"0C",X"FE",X"0B",X"28",X"08",
		X"E1",X"E5",X"23",X"23",X"CB",X"8E",X"18",X"0D",X"21",X"F0",X"87",X"CB",X"CE",X"E1",X"E5",X"23",
		X"23",X"CB",X"C6",X"CB",X"CE",X"CB",X"46",X"20",X"02",X"E1",X"C9",X"CB",X"4E",X"CA",X"BC",X"21",
		X"CB",X"56",X"20",X"0A",X"23",X"23",X"36",X"0C",X"2B",X"2B",X"CB",X"D6",X"E1",X"C9",X"23",X"23",
		X"7E",X"FE",X"0C",X"28",X"2B",X"FE",X"09",X"28",X"32",X"FE",X"06",X"28",X"23",X"FE",X"03",X"28",
		X"2A",X"FE",X"0A",X"38",X"02",X"18",X"2D",X"F5",X"E5",X"21",X"33",X"85",X"06",X"08",X"11",X"10",
		X"00",X"7E",X"E6",X"07",X"20",X"03",X"C6",X"04",X"77",X"19",X"10",X"F5",X"E1",X"F1",X"18",X"14",
		X"E5",X"F5",X"CD",X"0C",X"29",X"36",X"1F",X"F1",X"E1",X"18",X"09",X"E5",X"F5",X"CD",X"0C",X"29",
		X"36",X"1E",X"F1",X"E1",X"A7",X"28",X"0C",X"FE",X"01",X"20",X"05",X"3E",X"01",X"32",X"8D",X"9A",
		X"35",X"E1",X"C9",X"DD",X"E1",X"DD",X"E5",X"3A",X"46",X"86",X"CB",X"47",X"C2",X"A9",X"20",X"21",
		X"A2",X"98",X"DD",X"7E",X"00",X"BE",X"30",X"05",X"4F",X"7E",X"91",X"18",X"01",X"96",X"FE",X"07",
		X"D2",X"B6",X"20",X"23",X"DD",X"4E",X"01",X"7E",X"91",X"FE",X"12",X"30",X"29",X"AF",X"32",X"22",
		X"99",X"21",X"46",X"86",X"CB",X"C6",X"3E",X"01",X"32",X"8A",X"9A",X"DD",X"36",X"03",X"FF",X"3A",
		X"A3",X"98",X"D6",X"02",X"32",X"A3",X"98",X"18",X"0D",X"21",X"A3",X"98",X"7E",X"C6",X"08",X"77",
		X"FE",X"EE",X"38",X"02",X"36",X"EE",X"21",X"25",X"85",X"22",X"F6",X"85",X"11",X"04",X"00",X"19",
		X"22",X"1A",X"86",X"11",X"10",X"00",X"06",X"08",X"2A",X"F6",X"85",X"CB",X"7E",X"C2",X"9B",X"21",
		X"CB",X"6E",X"C2",X"A3",X"21",X"D5",X"11",X"06",X"00",X"19",X"D1",X"7E",X"FE",X"3F",X"38",X"49",
		X"2A",X"1A",X"86",X"3A",X"00",X"84",X"CB",X"4F",X"28",X"04",X"CB",X"57",X"20",X"03",X"7E",X"18",
		X"03",X"7E",X"D6",X"10",X"4F",X"DD",X"7E",X"00",X"B9",X"30",X"0C",X"79",X"DD",X"4E",X"00",X"91",
		X"FE",X"09",X"D2",X"A3",X"21",X"18",X"06",X"91",X"FE",X"19",X"D2",X"A3",X"21",X"23",X"DD",X"4E",
		X"01",X"3A",X"00",X"84",X"CB",X"4F",X"28",X"04",X"CB",X"57",X"20",X"03",X"7E",X"18",X"03",X"7E",
		X"D6",X"10",X"91",X"FE",X"0C",X"30",X"7C",X"18",X"1F",X"2A",X"1A",X"86",X"DD",X"7E",X"00",X"BE",
		X"30",X"05",X"4F",X"7E",X"91",X"18",X"01",X"96",X"FE",X"0C",X"30",X"67",X"23",X"DD",X"4E",X"01",
		X"7E",X"91",X"FE",X"0C",X"30",X"5D",X"18",X"28",X"DD",X"7E",X"01",X"C6",X"08",X"2A",X"1A",X"86",
		X"23",X"77",X"2B",X"3A",X"00",X"84",X"CB",X"4F",X"28",X"0A",X"CB",X"57",X"28",X"06",X"7E",X"D6",
		X"08",X"77",X"18",X"04",X"7E",X"C6",X"08",X"77",X"D5",X"2A",X"F6",X"85",X"CD",X"F8",X"26",X"D1",
		X"2A",X"F6",X"85",X"3E",X"C3",X"A6",X"77",X"CB",X"FE",X"D5",X"11",X"0D",X"00",X"19",X"D1",X"CB",
		X"9E",X"CB",X"96",X"3E",X"01",X"32",X"8A",X"9A",X"21",X"C5",X"87",X"CB",X"C6",X"DD",X"36",X"03",
		X"FF",X"2A",X"1A",X"86",X"23",X"7E",X"D6",X"02",X"77",X"18",X"08",X"2A",X"1A",X"86",X"23",X"7E",
		X"C6",X"08",X"77",X"2A",X"F6",X"85",X"19",X"22",X"F6",X"85",X"2A",X"1A",X"86",X"19",X"22",X"1A",
		X"86",X"05",X"C2",X"C8",X"20",X"E1",X"23",X"3E",X"08",X"86",X"77",X"C9",X"CB",X"5E",X"C2",X"6B",
		X"22",X"CB",X"DE",X"CB",X"FE",X"23",X"23",X"36",X"14",X"E1",X"11",X"03",X"00",X"19",X"CB",X"46",
		X"28",X"0D",X"2B",X"2B",X"3A",X"46",X"86",X"CB",X"47",X"20",X"04",X"7E",X"D6",X"08",X"77",X"3E",
		X"01",X"32",X"8C",X"9A",X"C9",X"21",X"C5",X"87",X"36",X"00",X"21",X"25",X"85",X"11",X"10",X"00",
		X"0E",X"00",X"06",X"08",X"22",X"F6",X"85",X"CB",X"7E",X"28",X"0E",X"0C",X"36",X"00",X"23",X"23",
		X"23",X"CB",X"FE",X"23",X"36",X"00",X"23",X"36",X"00",X"2A",X"F6",X"85",X"19",X"22",X"F6",X"85",
		X"10",X"E2",X"21",X"47",X"86",X"36",X"3C",X"21",X"1C",X"86",X"36",X"C8",X"21",X"46",X"86",X"CB",
		X"46",X"28",X"02",X"CB",X"CE",X"79",X"A7",X"CA",X"69",X"22",X"06",X"3E",X"80",X"32",X"74",X"98",
		X"3E",X"47",X"32",X"78",X"98",X"3E",X"0A",X"32",X"75",X"98",X"32",X"79",X"98",X"AF",X"32",X"74",
		X"99",X"32",X"78",X"99",X"E1",X"E5",X"7E",X"D6",X"08",X"32",X"F4",X"98",X"C6",X"10",X"32",X"F8",
		X"98",X"36",X"00",X"23",X"7E",X"32",X"F5",X"98",X"32",X"F9",X"98",X"36",X"00",X"E1",X"79",X"87",
		X"C8",X"81",X"C6",X"15",X"6F",X"CD",X"B5",X"2F",X"C9",X"E1",X"C9",X"23",X"23",X"7E",X"A7",X"28",
		X"35",X"35",X"FE",X"04",X"CA",X"E5",X"21",X"E5",X"21",X"C5",X"87",X"CB",X"46",X"28",X"03",X"E1",
		X"E1",X"C9",X"E1",X"FE",X"12",X"28",X"0A",X"FE",X"09",X"28",X"0D",X"FE",X"05",X"28",X"10",X"E1",
		X"C9",X"CD",X"0C",X"29",X"36",X"74",X"E1",X"C9",X"CD",X"0C",X"29",X"36",X"75",X"E1",X"C9",X"CD",
		X"0C",X"29",X"36",X"32",X"E1",X"C9",X"E1",X"AF",X"77",X"23",X"36",X"90",X"23",X"36",X"11",X"CD",
		X"62",X"19",X"23",X"77",X"32",X"F4",X"98",X"32",X"F5",X"98",X"32",X"F8",X"98",X"32",X"F9",X"98",
		X"21",X"99",X"87",X"CB",X"C6",X"21",X"F0",X"87",X"CB",X"8E",X"C9",X"C5",X"E5",X"D5",X"CD",X"10",
		X"1C",X"2A",X"FE",X"85",X"23",X"22",X"EA",X"85",X"2A",X"00",X"86",X"23",X"22",X"EC",X"85",X"2A",
		X"EA",X"85",X"7E",X"FE",X"7F",X"28",X"14",X"2A",X"EC",X"85",X"7E",X"FE",X"7F",X"28",X"0C",X"2A",
		X"FE",X"85",X"CD",X"FF",X"22",X"2A",X"00",X"86",X"CD",X"FF",X"22",X"D1",X"E1",X"C1",X"C9",X"E5",
		X"2B",X"7E",X"FE",X"7F",X"20",X"02",X"E1",X"C9",X"23",X"7E",X"FE",X"00",X"28",X"1F",X"3D",X"28",
		X"20",X"3D",X"3D",X"3D",X"28",X"17",X"3D",X"28",X"18",X"3D",X"28",X"15",X"3D",X"28",X"12",X"3D",
		X"28",X"13",X"3D",X"28",X"10",X"3D",X"28",X"05",X"3D",X"28",X"02",X"E1",X"C9",X"36",X"02",X"E1",
		X"C9",X"36",X"03",X"E1",X"C9",X"36",X"0C",X"E1",X"C9",X"E5",X"CD",X"8E",X"26",X"E1",X"3A",X"01",
		X"84",X"CB",X"7F",X"C0",X"CD",X"48",X"23",X"C9",X"E5",X"7E",X"E6",X"BC",X"C2",X"31",X"25",X"CB",
		X"4E",X"CA",X"1F",X"29",X"22",X"F6",X"85",X"11",X"0B",X"00",X"19",X"7E",X"A7",X"28",X"0E",X"FE",
		X"01",X"20",X"09",X"ED",X"5B",X"F6",X"85",X"EB",X"23",X"CB",X"86",X"EB",X"35",X"2A",X"F6",X"85",
		X"23",X"23",X"23",X"CB",X"7E",X"28",X"02",X"E1",X"C9",X"3A",X"BD",X"87",X"47",X"2A",X"F6",X"85",
		X"11",X"09",X"00",X"19",X"7E",X"90",X"77",X"38",X"02",X"E1",X"C9",X"2A",X"F6",X"85",X"11",X"04",
		X"00",X"19",X"7E",X"FE",X"01",X"20",X"05",X"2B",X"CB",X"FE",X"E1",X"C9",X"CD",X"F8",X"1C",X"2A",
		X"F6",X"85",X"23",X"CB",X"8E",X"2B",X"11",X"04",X"00",X"19",X"46",X"23",X"4E",X"2A",X"F6",X"85",
		X"23",X"23",X"23",X"CB",X"76",X"C2",X"02",X"24",X"3A",X"F0",X"87",X"CB",X"47",X"C2",X"02",X"24",
		X"3A",X"A2",X"98",X"B8",X"DA",X"CA",X"23",X"90",X"18",X"06",X"3A",X"A2",X"98",X"57",X"78",X"92",
		X"FE",X"20",X"D2",X"02",X"24",X"3A",X"A3",X"98",X"B9",X"DA",X"DF",X"23",X"91",X"18",X"06",X"3A",
		X"A3",X"98",X"57",X"79",X"92",X"FE",X"20",X"D2",X"02",X"24",X"2A",X"F6",X"85",X"11",X"0F",X"00",
		X"19",X"3A",X"A3",X"98",X"77",X"2B",X"3A",X"A2",X"98",X"77",X"2A",X"F6",X"85",X"23",X"23",X"23",
		X"CB",X"F6",X"3A",X"F4",X"85",X"CB",X"4F",X"28",X"4A",X"2A",X"F6",X"85",X"23",X"23",X"23",X"CB",
		X"76",X"28",X"0E",X"3A",X"F0",X"87",X"CB",X"47",X"20",X"07",X"11",X"0C",X"00",X"19",X"7E",X"18",
		X"0E",X"3A",X"F0",X"87",X"CB",X"47",X"28",X"04",X"3E",X"08",X"18",X"03",X"3A",X"A3",X"98",X"B9",
		X"DA",X"4A",X"24",X"CA",X"90",X"24",X"CD",X"3F",X"24",X"19",X"34",X"34",X"C3",X"90",X"24",X"2A",
		X"F6",X"85",X"23",X"CB",X"CE",X"2B",X"11",X"05",X"00",X"C9",X"CD",X"3F",X"24",X"19",X"35",X"35",
		X"C3",X"90",X"24",X"2A",X"F6",X"85",X"23",X"23",X"23",X"CB",X"76",X"28",X"0E",X"3A",X"F0",X"87",
		X"CB",X"47",X"20",X"07",X"11",X"0B",X"00",X"19",X"7E",X"18",X"0E",X"3A",X"F0",X"87",X"CB",X"47",
		X"28",X"04",X"3E",X"21",X"18",X"03",X"3A",X"A2",X"98",X"B8",X"DA",X"88",X"24",X"CA",X"90",X"24",
		X"2A",X"F6",X"85",X"11",X"04",X"00",X"18",X"B1",X"2A",X"F6",X"85",X"11",X"04",X"00",X"18",X"BD",
		X"21",X"4A",X"86",X"CB",X"F6",X"2A",X"F6",X"85",X"23",X"CB",X"46",X"C2",X"04",X"25",X"06",X"00",
		X"2A",X"F6",X"85",X"23",X"CB",X"4E",X"CC",X"A1",X"28",X"C4",X"B7",X"28",X"CB",X"40",X"CA",X"04",
		X"25",X"CD",X"DB",X"28",X"CB",X"40",X"CA",X"04",X"25",X"2A",X"F6",X"85",X"CB",X"8E",X"23",X"CB",
		X"4E",X"20",X"28",X"23",X"23",X"23",X"23",X"7E",X"FE",X"20",X"D2",X"D7",X"24",X"FE",X"16",X"D2",
		X"DE",X"24",X"36",X"08",X"C3",X"1F",X"25",X"E6",X"0F",X"FE",X"08",X"DA",X"E7",X"24",X"0E",X"10",
		X"7E",X"E6",X"F0",X"81",X"77",X"E1",X"C9",X"0E",X"00",X"18",X"F5",X"23",X"23",X"23",X"7E",X"E6",
		X"0F",X"FE",X"08",X"DA",X"FF",X"24",X"7E",X"E6",X"F0",X"C6",X"11",X"77",X"C3",X"1F",X"25",X"7E",
		X"E6",X"F0",X"3C",X"77",X"21",X"4A",X"86",X"CB",X"76",X"28",X"14",X"CB",X"B6",X"2A",X"F6",X"85",
		X"23",X"CB",X"4E",X"28",X"05",X"CB",X"8E",X"C3",X"95",X"24",X"CB",X"CE",X"C3",X"95",X"24",X"E1",
		X"C9",X"7E",X"E6",X"7F",X"FE",X"10",X"DA",X"2F",X"25",X"FE",X"7E",X"CA",X"2F",X"25",X"C9",X"0D",
		X"C9",X"22",X"F6",X"85",X"2A",X"F6",X"85",X"23",X"23",X"CB",X"66",X"C2",X"C7",X"25",X"2A",X"F6",
		X"85",X"CB",X"46",X"C2",X"37",X"26",X"2A",X"F6",X"85",X"7E",X"E6",X"3C",X"CA",X"C7",X"25",X"11",
		X"0C",X"00",X"19",X"35",X"7E",X"FE",X"0D",X"C2",X"C9",X"25",X"2A",X"F6",X"85",X"CB",X"6E",X"CA",
		X"C7",X"25",X"11",X"04",X"00",X"19",X"3A",X"00",X"84",X"E6",X"06",X"FE",X"06",X"C2",X"85",X"25",
		X"7E",X"32",X"FE",X"98",X"D6",X"10",X"32",X"F6",X"98",X"23",X"7E",X"D6",X"09",X"32",X"FF",X"98",
		X"32",X"F7",X"98",X"18",X"13",X"7E",X"32",X"F6",X"98",X"C6",X"10",X"32",X"FE",X"98",X"23",X"7E",
		X"C6",X"07",X"32",X"F7",X"98",X"32",X"FF",X"98",X"2A",X"F6",X"85",X"CB",X"EE",X"23",X"23",X"CB",
		X"C6",X"23",X"CB",X"FE",X"2B",X"2B",X"2B",X"11",X"04",X"00",X"19",X"36",X"F1",X"23",X"36",X"00",
		X"23",X"36",X"32",X"11",X"07",X"00",X"19",X"CB",X"96",X"CB",X"9E",X"AF",X"32",X"A0",X"98",X"32",
		X"A1",X"98",X"21",X"03",X"84",X"CB",X"96",X"E1",X"C9",X"A7",X"C2",X"C7",X"25",X"21",X"DF",X"32",
		X"3A",X"10",X"84",X"3D",X"5F",X"16",X"00",X"19",X"7E",X"2A",X"F6",X"85",X"11",X"0C",X"00",X"19",
		X"77",X"2A",X"F6",X"85",X"CB",X"56",X"28",X"1B",X"CB",X"96",X"CB",X"B6",X"21",X"9E",X"87",X"3A",
		X"9D",X"87",X"BE",X"20",X"0C",X"CD",X"89",X"0F",X"21",X"03",X"84",X"CB",X"96",X"2B",X"2B",X"CB",
		X"9E",X"E1",X"C9",X"CB",X"5E",X"28",X"06",X"CB",X"9E",X"CB",X"D6",X"18",X"08",X"CB",X"66",X"28",
		X"0A",X"CB",X"A6",X"CB",X"DE",X"23",X"23",X"CB",X"EE",X"E1",X"C9",X"CB",X"6E",X"20",X"02",X"E1",
		X"C9",X"CB",X"AE",X"21",X"04",X"84",X"CB",X"B6",X"AF",X"32",X"F6",X"98",X"32",X"F7",X"98",X"32",
		X"FE",X"98",X"32",X"FF",X"98",X"E1",X"C9",X"3A",X"29",X"86",X"E5",X"C5",X"3D",X"28",X"10",X"3D",
		X"28",X"12",X"3D",X"20",X"05",X"21",X"A4",X"98",X"18",X"0D",X"21",X"B6",X"98",X"18",X"08",X"21",
		X"AA",X"98",X"18",X"03",X"21",X"B0",X"98",X"06",X"03",X"36",X"00",X"23",X"36",X"50",X"23",X"10",
		X"F8",X"C1",X"E1",X"C3",X"46",X"25",X"11",X"06",X"00",X"19",X"22",X"F6",X"85",X"11",X"04",X"00",
		X"19",X"34",X"7E",X"E6",X"0F",X"FE",X"08",X"DA",X"84",X"26",X"2A",X"F6",X"85",X"36",X"2A",X"23",
		X"36",X"03",X"E1",X"C9",X"2A",X"F6",X"85",X"36",X"2B",X"23",X"36",X"03",X"E1",X"C9",X"E5",X"7E",
		X"E6",X"FC",X"C2",X"C7",X"26",X"CB",X"4E",X"CA",X"2D",X"28",X"CB",X"46",X"C2",X"66",X"26",X"11",
		X"06",X"00",X"19",X"22",X"F6",X"85",X"11",X"04",X"00",X"19",X"34",X"7E",X"E6",X"0F",X"FE",X"08",
		X"DA",X"BD",X"26",X"2A",X"F6",X"85",X"36",X"28",X"23",X"36",X"03",X"E1",X"C9",X"2A",X"F6",X"85",
		X"36",X"29",X"23",X"36",X"03",X"E1",X"C9",X"CB",X"7F",X"28",X"3C",X"3A",X"9E",X"87",X"57",X"3A",
		X"9D",X"87",X"BA",X"20",X"13",X"E5",X"CD",X"89",X"0F",X"21",X"01",X"84",X"CB",X"9E",X"23",X"23",
		X"CB",X"96",X"21",X"3E",X"86",X"36",X"00",X"E1",X"CB",X"46",X"C2",X"FC",X"26",X"11",X"06",X"00",
		X"19",X"36",X"22",X"23",X"36",X"01",X"E1",X"C9",X"E5",X"C3",X"E8",X"26",X"11",X"06",X"00",X"19",
		X"36",X"26",X"23",X"36",X"02",X"E1",X"C9",X"22",X"F6",X"85",X"11",X"07",X"00",X"19",X"E5",X"DD",
		X"E1",X"2B",X"E5",X"FD",X"E1",X"2A",X"F6",X"85",X"23",X"23",X"CB",X"46",X"CA",X"21",X"27",X"E1",
		X"C9",X"2A",X"F6",X"85",X"CB",X"46",X"C2",X"E4",X"27",X"DD",X"36",X"00",X"01",X"CB",X"56",X"28",
		X"21",X"FD",X"36",X"00",X"23",X"23",X"23",X"CB",X"6E",X"C2",X"3E",X"27",X"E1",X"C9",X"CB",X"AE",
		X"3A",X"00",X"84",X"E6",X"06",X"FE",X"06",X"CA",X"8B",X"27",X"CD",X"A9",X"27",X"C6",X"04",X"77",
		X"E1",X"C9",X"CB",X"5E",X"28",X"70",X"FD",X"36",X"00",X"80",X"23",X"23",X"CB",X"6E",X"C2",X"68",
		X"27",X"CB",X"66",X"C2",X"77",X"27",X"E1",X"C9",X"CB",X"AE",X"2A",X"F6",X"85",X"11",X"05",X"00",
		X"19",X"7E",X"C6",X"04",X"77",X"E1",X"C9",X"CB",X"A6",X"3A",X"00",X"84",X"E6",X"06",X"FE",X"06",
		X"CA",X"93",X"27",X"CD",X"9B",X"27",X"D6",X"04",X"77",X"E1",X"C9",X"CD",X"9B",X"27",X"D6",X"0C",
		X"77",X"E1",X"C9",X"CD",X"A9",X"27",X"C6",X"0C",X"77",X"E1",X"C9",X"2A",X"F6",X"85",X"11",X"04",
		X"00",X"19",X"7E",X"D6",X"08",X"77",X"23",X"7E",X"C9",X"2A",X"F6",X"85",X"11",X"04",X"00",X"19",
		X"7E",X"C6",X"08",X"77",X"23",X"7E",X"C9",X"CB",X"A6",X"2A",X"F6",X"85",X"11",X"05",X"00",X"19",
		X"7E",X"D6",X"04",X"77",X"E1",X"C9",X"CB",X"66",X"28",X"0D",X"FD",X"36",X"00",X"81",X"23",X"23",
		X"CB",X"66",X"C2",X"B7",X"27",X"E1",X"C9",X"CB",X"6E",X"28",X"07",X"FD",X"36",X"00",X"82",X"CD",
		X"89",X"0F",X"E1",X"C9",X"DD",X"36",X"00",X"02",X"CB",X"56",X"28",X"0D",X"FD",X"36",X"00",X"27",
		X"23",X"23",X"CB",X"6E",X"C2",X"3E",X"27",X"E1",X"C9",X"CB",X"5E",X"28",X"12",X"FD",X"36",X"00",
		X"83",X"23",X"23",X"CB",X"6E",X"C2",X"68",X"27",X"CB",X"66",X"C2",X"77",X"27",X"E1",X"C9",X"CB",
		X"66",X"28",X"0D",X"FD",X"36",X"00",X"84",X"23",X"23",X"CB",X"66",X"C2",X"B7",X"27",X"E1",X"C9",
		X"CB",X"6E",X"28",X"07",X"FD",X"36",X"00",X"85",X"CD",X"89",X"0F",X"E1",X"C9",X"3A",X"01",X"84",
		X"CB",X"7F",X"28",X"02",X"E1",X"C9",X"11",X"0E",X"00",X"19",X"7E",X"E6",X"07",X"FE",X"02",X"28",
		X"09",X"FE",X"06",X"20",X"08",X"2B",X"36",X"02",X"18",X"03",X"2B",X"36",X"00",X"E1",X"E5",X"CB",
		X"46",X"20",X"1C",X"11",X"06",X"00",X"CD",X"94",X"28",X"FE",X"04",X"DA",X"68",X"28",X"2A",X"F6",
		X"85",X"36",X"21",X"23",X"36",X"01",X"E1",X"C9",X"2A",X"F6",X"85",X"36",X"20",X"18",X"F4",X"23",
		X"CB",X"76",X"28",X"02",X"E1",X"C9",X"11",X"05",X"00",X"CD",X"94",X"28",X"E6",X"07",X"FE",X"04",
		X"DA",X"8D",X"28",X"2A",X"F6",X"85",X"36",X"25",X"23",X"36",X"02",X"E1",X"C9",X"2A",X"F6",X"85",
		X"36",X"24",X"18",X"F4",X"19",X"22",X"F6",X"85",X"11",X"04",X"00",X"19",X"34",X"7E",X"E6",X"0F",
		X"C9",X"E5",X"F5",X"23",X"23",X"23",X"7E",X"E6",X"0F",X"FE",X"01",X"28",X"05",X"CB",X"80",X"F1",
		X"E1",X"C9",X"CB",X"C0",X"F1",X"E1",X"C9",X"E5",X"F5",X"23",X"23",X"23",X"23",X"7E",X"4F",X"E6",
		X"0F",X"57",X"79",X"FE",X"20",X"D2",X"D2",X"28",X"FE",X"08",X"CA",X"D6",X"28",X"CB",X"80",X"F1",
		X"E1",X"C9",X"7A",X"A7",X"20",X"F7",X"CB",X"C0",X"F1",X"E1",X"C9",X"2A",X"F6",X"85",X"11",X"04",
		X"00",X"19",X"56",X"23",X"5E",X"CD",X"10",X"1C",X"0E",X"04",X"2A",X"FA",X"85",X"CD",X"21",X"25",
		X"2A",X"FC",X"85",X"CD",X"21",X"25",X"2A",X"FE",X"85",X"CD",X"21",X"25",X"2A",X"00",X"86",X"CD",
		X"21",X"25",X"79",X"A7",X"28",X"03",X"CB",X"80",X"C9",X"CB",X"C0",X"C9",X"11",X"69",X"84",X"A7",
		X"ED",X"52",X"7D",X"CB",X"3F",X"CB",X"3F",X"5F",X"16",X"00",X"21",X"3C",X"98",X"19",X"C9",X"22",
		X"F6",X"85",X"11",X"04",X"00",X"19",X"7E",X"FE",X"01",X"C2",X"31",X"29",X"2B",X"CB",X"FE",X"E1",
		X"C9",X"11",X"0B",X"00",X"19",X"22",X"1A",X"86",X"2A",X"F6",X"85",X"23",X"23",X"CB",X"A6",X"CB",
		X"AE",X"23",X"CB",X"B6",X"CB",X"7E",X"28",X"02",X"E1",X"C9",X"2A",X"F6",X"85",X"11",X"05",X"00",
		X"19",X"7E",X"FE",X"08",X"C2",X"6A",X"29",X"3A",X"BD",X"87",X"2A",X"F6",X"85",X"CB",X"46",X"28",
		X"06",X"C6",X"0A",X"30",X"02",X"3E",X"FF",X"47",X"18",X"41",X"3A",X"46",X"86",X"CB",X"5F",X"28",
		X"11",X"2A",X"F6",X"85",X"CB",X"46",X"28",X"05",X"21",X"A5",X"87",X"18",X"2C",X"21",X"A2",X"87",
		X"18",X"27",X"3A",X"53",X"86",X"CB",X"4F",X"28",X"11",X"2A",X"F6",X"85",X"CB",X"46",X"28",X"05",
		X"21",X"A4",X"87",X"18",X"14",X"21",X"A1",X"87",X"18",X"0F",X"2A",X"F6",X"85",X"CB",X"46",X"28",
		X"05",X"21",X"A3",X"87",X"18",X"03",X"21",X"A0",X"87",X"00",X"46",X"2A",X"F6",X"85",X"11",X"0E",
		X"00",X"19",X"7E",X"E6",X"07",X"FE",X"04",X"20",X"19",X"3A",X"57",X"86",X"CB",X"4F",X"20",X"07",
		X"3A",X"0F",X"84",X"FE",X"04",X"38",X"0B",X"3A",X"EE",X"32",X"80",X"47",X"FE",X"28",X"30",X"02",
		X"06",X"FF",X"2A",X"F6",X"85",X"11",X"09",X"00",X"19",X"7E",X"90",X"77",X"38",X"02",X"E1",X"C9",
		X"2A",X"F6",X"85",X"23",X"CD",X"A1",X"28",X"CB",X"40",X"20",X"0B",X"CD",X"B7",X"28",X"CB",X"40",
		X"CA",X"71",X"2C",X"C3",X"E2",X"2C",X"CD",X"B7",X"28",X"CB",X"40",X"CA",X"E2",X"2C",X"23",X"23",
		X"23",X"56",X"23",X"5E",X"CD",X"16",X"1C",X"2A",X"F6",X"85",X"CB",X"46",X"CA",X"28",X"2C",X"11",
		X"06",X"00",X"19",X"7E",X"FE",X"2A",X"CA",X"28",X"2C",X"FE",X"2B",X"CA",X"28",X"2C",X"FE",X"27",
		X"C2",X"25",X"2A",X"36",X"24",X"2A",X"1A",X"86",X"2B",X"CB",X"4E",X"CA",X"28",X"2C",X"2A",X"F6",
		X"85",X"11",X"04",X"00",X"19",X"7E",X"FE",X"D1",X"D2",X"28",X"2C",X"FE",X"22",X"DA",X"28",X"2C",
		X"CD",X"D4",X"2E",X"78",X"FE",X"03",X"CA",X"28",X"2C",X"2A",X"F6",X"85",X"23",X"CB",X"76",X"C2",
		X"A4",X"2A",X"21",X"D0",X"32",X"3A",X"0F",X"84",X"3D",X"E6",X"0F",X"5F",X"16",X"00",X"19",X"46",
		X"2A",X"F6",X"85",X"11",X"04",X"00",X"19",X"3A",X"A2",X"98",X"BE",X"38",X"03",X"96",X"18",X"03",
		X"4F",X"7E",X"91",X"FE",X"3C",X"30",X"15",X"3A",X"A3",X"98",X"23",X"BE",X"38",X"03",X"96",X"18",
		X"03",X"4F",X"7E",X"91",X"FE",X"3C",X"30",X"04",X"78",X"87",X"87",X"47",X"CD",X"F8",X"1C",X"3A",
		X"F4",X"85",X"90",X"D2",X"28",X"2C",X"2A",X"F6",X"85",X"23",X"CB",X"F6",X"11",X"0A",X"00",X"19",
		X"36",X"0E",X"E1",X"C9",X"DD",X"21",X"A4",X"98",X"FD",X"21",X"A5",X"98",X"21",X"24",X"98",X"01",
		X"24",X"99",X"3A",X"29",X"86",X"FE",X"01",X"28",X"12",X"FE",X"02",X"28",X"09",X"FE",X"03",X"28",
		X"19",X"11",X"12",X"00",X"18",X"08",X"11",X"0C",X"00",X"18",X"03",X"11",X"06",X"00",X"19",X"E5",
		X"C5",X"E1",X"19",X"E5",X"C1",X"E1",X"DD",X"19",X"FD",X"19",X"EB",X"2A",X"1A",X"86",X"2B",X"7E",
		X"2A",X"F6",X"85",X"23",X"23",X"23",X"23",X"E6",X"07",X"FE",X"02",X"28",X"1C",X"7E",X"D6",X"10",
		X"DD",X"77",X"00",X"DD",X"23",X"DD",X"23",X"D6",X"10",X"DD",X"77",X"00",X"DD",X"23",X"DD",X"23",
		X"D6",X"10",X"DD",X"77",X"00",X"3E",X"02",X"18",X"19",X"7E",X"C6",X"10",X"DD",X"77",X"00",X"DD",
		X"23",X"DD",X"23",X"C6",X"10",X"DD",X"77",X"00",X"DD",X"23",X"DD",X"23",X"C6",X"10",X"DD",X"77",
		X"00",X"AF",X"02",X"03",X"03",X"02",X"03",X"03",X"02",X"23",X"7E",X"FD",X"77",X"00",X"FD",X"23",
		X"FD",X"23",X"FD",X"77",X"00",X"FD",X"23",X"FD",X"23",X"FD",X"77",X"00",X"ED",X"53",X"27",X"86",
		X"2A",X"F6",X"85",X"11",X"0B",X"00",X"19",X"35",X"4E",X"2A",X"F6",X"85",X"11",X"08",X"00",X"19",
		X"7E",X"A7",X"20",X"28",X"79",X"A7",X"28",X"5D",X"3D",X"CA",X"13",X"2C",X"3D",X"CA",X"13",X"2C",
		X"3D",X"CA",X"F8",X"2B",X"3D",X"28",X"68",X"3D",X"28",X"3D",X"3D",X"3D",X"28",X"2E",X"3D",X"3D",
		X"28",X"35",X"3D",X"3D",X"28",X"26",X"3D",X"3D",X"28",X"2D",X"E1",X"C9",X"FE",X"01",X"20",X"0F",
		X"79",X"3D",X"28",X"31",X"3D",X"28",X"71",X"3D",X"28",X"6E",X"3D",X"28",X"42",X"18",X"D8",X"79",
		X"3D",X"3D",X"28",X"21",X"3D",X"28",X"38",X"3D",X"28",X"35",X"18",X"CB",X"2A",X"F6",X"85",X"11",
		X"07",X"00",X"19",X"36",X"02",X"18",X"09",X"2A",X"F6",X"85",X"11",X"07",X"00",X"19",X"36",X"0C",
		X"CD",X"9D",X"2F",X"E1",X"C9",X"2A",X"F6",X"85",X"23",X"CB",X"B6",X"CD",X"9D",X"2F",X"2A",X"27",
		X"86",X"3E",X"32",X"77",X"23",X"23",X"77",X"23",X"23",X"77",X"CD",X"5F",X"15",X"E1",X"C9",X"2A",
		X"27",X"86",X"36",X"2C",X"23",X"36",X"05",X"23",X"36",X"32",X"23",X"23",X"36",X"32",X"DD",X"2B",
		X"DD",X"2B",X"DD",X"2B",X"DD",X"2B",X"FD",X"2B",X"FD",X"2B",X"FD",X"2B",X"FD",X"2B",X"CD",X"5F",
		X"15",X"21",X"8E",X"9A",X"36",X"01",X"E1",X"C9",X"2A",X"27",X"86",X"3E",X"05",X"36",X"2D",X"23",
		X"77",X"23",X"36",X"2E",X"23",X"77",X"23",X"36",X"32",X"DD",X"2B",X"DD",X"2B",X"FD",X"2B",X"FD",
		X"2B",X"18",X"B7",X"2A",X"27",X"86",X"3E",X"05",X"36",X"2F",X"23",X"77",X"23",X"36",X"30",X"23",
		X"77",X"23",X"36",X"31",X"23",X"77",X"18",X"A2",X"CD",X"F8",X"1C",X"3A",X"F4",X"85",X"CB",X"47",
		X"20",X"12",X"CD",X"3A",X"2D",X"CB",X"41",X"C2",X"CE",X"2C",X"CD",X"67",X"2D",X"CB",X"41",X"C2",
		X"CE",X"2C",X"18",X"10",X"CD",X"67",X"2D",X"CB",X"41",X"C2",X"CE",X"2C",X"CD",X"3A",X"2D",X"CB",
		X"41",X"C2",X"CE",X"2C",X"2A",X"1A",X"86",X"2B",X"7E",X"23",X"77",X"CD",X"A8",X"2D",X"CB",X"41",
		X"C2",X"CE",X"2C",X"CD",X"F8",X"1C",X"3A",X"F4",X"85",X"E6",X"0F",X"FE",X"0A",X"38",X"1E",X"18",
		X"44",X"2A",X"F6",X"85",X"CB",X"CE",X"23",X"CB",X"C6",X"11",X"0A",X"00",X"19",X"36",X"28",X"23",
		X"23",X"23",X"7E",X"3C",X"3C",X"77",X"CD",X"7A",X"2F",X"36",X"03",X"E1",X"C9",X"2A",X"1A",X"86",
		X"2B",X"7E",X"23",X"77",X"35",X"35",X"CD",X"A8",X"2D",X"CB",X"41",X"F5",X"C4",X"92",X"2F",X"F1",
		X"20",X"2C",X"2A",X"1A",X"86",X"34",X"34",X"34",X"34",X"CD",X"A8",X"2D",X"CB",X"41",X"F5",X"C4",
		X"98",X"2F",X"F1",X"20",X"19",X"2A",X"1A",X"86",X"2B",X"7E",X"23",X"3C",X"3C",X"3C",X"3C",X"77",
		X"CD",X"A8",X"2D",X"CB",X"41",X"F5",X"C4",X"98",X"2F",X"F1",X"20",X"02",X"18",X"A3",X"CD",X"7A",
		X"2F",X"7E",X"FE",X"06",X"38",X"04",X"FE",X"C0",X"38",X"97",X"2A",X"1A",X"86",X"7E",X"E6",X"07",
		X"2B",X"77",X"2A",X"F6",X"85",X"11",X"05",X"00",X"19",X"7E",X"FE",X"08",X"20",X"0F",X"3A",X"F0",
		X"87",X"CB",X"47",X"28",X"08",X"2A",X"1A",X"86",X"2B",X"36",X"06",X"18",X"11",X"2A",X"1A",X"86",
		X"2B",X"7E",X"E6",X"07",X"28",X"1E",X"FE",X"02",X"28",X"0F",X"FE",X"04",X"28",X"1B",X"11",X"04",
		X"00",X"2A",X"F6",X"85",X"19",X"35",X"35",X"E1",X"C9",X"11",X"04",X"00",X"2A",X"F6",X"85",X"19",
		X"34",X"34",X"E1",X"C9",X"11",X"05",X"00",X"18",X"E8",X"2A",X"F6",X"85",X"11",X"05",X"00",X"19",
		X"3A",X"F0",X"87",X"CB",X"47",X"C2",X"71",X"2C",X"18",X"E6",X"2A",X"F6",X"85",X"CB",X"46",X"C2",
		X"55",X"2F",X"3A",X"A2",X"98",X"21",X"F0",X"87",X"CB",X"46",X"CA",X"4E",X"2D",X"AF",X"2A",X"F6",
		X"85",X"11",X"04",X"00",X"19",X"BE",X"CA",X"A1",X"2D",X"D2",X"61",X"2D",X"3E",X"06",X"C3",X"63",
		X"2D",X"3E",X"02",X"23",X"C3",X"90",X"2D",X"2A",X"F6",X"85",X"CB",X"46",X"C2",X"68",X"2F",X"3A",
		X"A3",X"98",X"21",X"F0",X"87",X"CB",X"46",X"CA",X"7C",X"2D",X"3E",X"08",X"2A",X"F6",X"85",X"11",
		X"05",X"00",X"19",X"BE",X"CA",X"A1",X"2D",X"D2",X"8E",X"2D",X"AF",X"C3",X"90",X"2D",X"3E",X"04",
		X"11",X"0A",X"00",X"19",X"77",X"E6",X"07",X"47",X"2B",X"7E",X"C6",X"04",X"E6",X"07",X"B8",X"20",
		X"03",X"0E",X"00",X"C9",X"CD",X"A8",X"2D",X"C9",X"2A",X"1A",X"86",X"7E",X"E6",X"07",X"28",X"22",
		X"FE",X"02",X"28",X"35",X"FE",X"04",X"28",X"4B",X"2A",X"02",X"86",X"22",X"12",X"86",X"11",X"20",
		X"00",X"19",X"22",X"16",X"86",X"2A",X"06",X"86",X"22",X"14",X"86",X"19",X"22",X"18",X"86",X"C3",
		X"63",X"2E",X"2A",X"02",X"86",X"22",X"12",X"86",X"2B",X"22",X"16",X"86",X"2A",X"04",X"86",X"22",
		X"14",X"86",X"2B",X"22",X"18",X"86",X"C3",X"21",X"2E",X"2A",X"04",X"86",X"22",X"12",X"86",X"11",
		X"E0",X"FF",X"19",X"22",X"16",X"86",X"2A",X"08",X"86",X"22",X"14",X"86",X"19",X"22",X"18",X"86",
		X"C3",X"63",X"2E",X"2A",X"06",X"86",X"22",X"12",X"86",X"23",X"22",X"16",X"86",X"2A",X"08",X"86",
		X"22",X"14",X"86",X"23",X"22",X"18",X"86",X"3A",X"F0",X"87",X"CB",X"47",X"28",X"03",X"0E",X"00",
		X"C9",X"2A",X"12",X"86",X"CD",X"42",X"2E",X"79",X"FE",X"00",X"C8",X"2A",X"14",X"86",X"CD",X"42",
		X"2E",X"79",X"FE",X"00",X"C8",X"2A",X"16",X"86",X"CD",X"42",X"2E",X"79",X"FE",X"00",X"C8",X"2A",
		X"18",X"86",X"7E",X"FE",X"02",X"28",X"19",X"FE",X"03",X"28",X"15",X"FE",X"7E",X"28",X"11",X"FE",
		X"8E",X"28",X"0D",X"FE",X"8F",X"28",X"09",X"CB",X"BF",X"FE",X"0C",X"28",X"03",X"0E",X"00",X"C9",
		X"0E",X"01",X"C9",X"2A",X"12",X"86",X"CD",X"84",X"2E",X"79",X"FE",X"00",X"C8",X"2A",X"14",X"86",
		X"CD",X"84",X"2E",X"79",X"FE",X"00",X"C8",X"2A",X"16",X"86",X"CD",X"84",X"2E",X"79",X"FE",X"00",
		X"C8",X"2A",X"18",X"86",X"7E",X"FE",X"8D",X"CA",X"A3",X"2E",X"FE",X"7E",X"CA",X"A3",X"2E",X"FE",
		X"08",X"CA",X"A3",X"2E",X"FE",X"09",X"CA",X"A3",X"2E",X"CB",X"BF",X"FE",X"0C",X"CA",X"A3",X"2E",
		X"0E",X"00",X"C9",X"0E",X"01",X"C9",X"7E",X"FE",X"8C",X"CA",X"D1",X"2E",X"FE",X"7E",X"CA",X"D1",
		X"2E",X"FE",X"09",X"CA",X"D1",X"2E",X"FE",X"08",X"CA",X"D1",X"2E",X"FE",X"0C",X"CA",X"D1",X"2E",
		X"FE",X"02",X"CA",X"D1",X"2E",X"FE",X"8D",X"CA",X"D1",X"2E",X"FE",X"03",X"CA",X"D1",X"2E",X"AF",
		X"C9",X"3E",X"01",X"C9",X"E5",X"2A",X"1A",X"86",X"2B",X"7E",X"E6",X"07",X"FE",X"02",X"CA",X"EA",
		X"2E",X"FE",X"06",X"CA",X"F8",X"2E",X"06",X"03",X"E1",X"C9",X"2A",X"02",X"86",X"22",X"36",X"86",
		X"2A",X"06",X"86",X"22",X"38",X"86",X"18",X"0C",X"2A",X"04",X"86",X"22",X"36",X"86",X"2A",X"08",
		X"86",X"22",X"38",X"86",X"06",X"03",X"2A",X"1A",X"86",X"2B",X"7E",X"E6",X"07",X"FE",X"02",X"CA",
		X"1A",X"2F",X"FE",X"06",X"CA",X"2E",X"2F",X"AF",X"E1",X"C9",X"11",X"C0",X"FF",X"2A",X"36",X"86",
		X"19",X"22",X"36",X"86",X"2A",X"38",X"86",X"19",X"22",X"38",X"86",X"C3",X"33",X"2F",X"11",X"40",
		X"00",X"18",X"EA",X"2A",X"36",X"86",X"CD",X"A6",X"2E",X"CB",X"47",X"CA",X"4B",X"2F",X"2A",X"38",
		X"86",X"CD",X"A6",X"2E",X"CB",X"47",X"CA",X"4B",X"2F",X"10",X"BB",X"2A",X"F6",X"85",X"11",X"08",
		X"00",X"19",X"70",X"E1",X"C9",X"3A",X"A2",X"98",X"2A",X"F6",X"85",X"11",X"04",X"00",X"19",X"BE",
		X"D2",X"61",X"2D",X"3E",X"06",X"C3",X"63",X"2D",X"3A",X"A3",X"98",X"2A",X"F6",X"85",X"11",X"05",
		X"00",X"19",X"BE",X"D2",X"8E",X"2D",X"AF",X"C3",X"90",X"2D",X"2A",X"F6",X"85",X"11",X"25",X"85",
		X"A7",X"ED",X"52",X"7D",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"5F",X"16",X"00",X"21",X"4B",X"86",
		X"19",X"C9",X"CD",X"7A",X"2F",X"36",X"03",X"C9",X"CD",X"7A",X"2F",X"34",X"C9",X"3E",X"50",X"FD",
		X"77",X"00",X"FD",X"77",X"FE",X"FD",X"77",X"FC",X"AF",X"DD",X"77",X"00",X"DD",X"77",X"FE",X"DD",
		X"77",X"FC",X"C9",X"2E",X"00",X"26",X"00",X"11",X"2B",X"30",X"19",X"11",X"11",X"84",X"7E",X"12",
		X"23",X"13",X"7E",X"12",X"23",X"13",X"7E",X"12",X"3A",X"57",X"86",X"CB",X"4F",X"C0",X"3A",X"81",
		X"9A",X"FE",X"00",X"C0",X"11",X"11",X"84",X"21",X"EF",X"89",X"A7",X"06",X"03",X"1A",X"8E",X"27",
		X"77",X"23",X"13",X"10",X"F8",X"3E",X"00",X"8E",X"27",X"77",X"3A",X"00",X"84",X"CB",X"4F",X"20",
		X"05",X"11",X"14",X"84",X"18",X"03",X"11",X"17",X"84",X"21",X"11",X"84",X"A7",X"06",X"03",X"1A",
		X"8E",X"27",X"12",X"13",X"23",X"10",X"F8",X"1B",X"EB",X"22",X"27",X"86",X"11",X"29",X"89",X"06",
		X"03",X"1A",X"BE",X"20",X"05",X"2B",X"1B",X"10",X"F8",X"C9",X"D0",X"21",X"29",X"89",X"ED",X"5B",
		X"27",X"86",X"06",X"03",X"1A",X"77",X"2B",X"1B",X"10",X"FA",X"C9",X"10",X"00",X"00",X"00",X"02",
		X"00",X"00",X"03",X"00",X"00",X"04",X"00",X"00",X"05",X"00",X"00",X"04",X"00",X"00",X"06",X"00",
		X"00",X"08",X"00",X"00",X"10",X"00",X"00",X"25",X"00",X"00",X"40",X"00",X"00",X"60",X"00",X"00",
		X"80",X"00",X"00",X"00",X"01",X"00",X"20",X"01",X"00",X"50",X"01",X"34",X"7F",X"32",X"1D",X"1A",
		X"1E",X"2B",X"2D",X"22",X"1D",X"1E",X"2B",X"1C",X"7F",X"2B",X"28",X"2E",X"27",X"1D",X"7F",X"32",
		X"25",X"27",X"28",X"7F",X"2B",X"1E",X"32",X"1A",X"25",X"29",X"7F",X"51",X"2C",X"2B",X"1E",X"32",
		X"1A",X"25",X"29",X"7F",X"52",X"7F",X"2B",X"28",X"7F",X"51",X"35",X"1D",X"2D",X"25",X"7F",X"28",
		X"1C",X"26",X"1A",X"27",X"7F",X"12",X"18",X"19",X"11",X"7F",X"38",X"BF",X"BE",X"BD",X"BC",X"BB",
		X"BA",X"B9",X"7F",X"27",X"28",X"2D",X"2D",X"2E",X"1B",X"7F",X"2D",X"2B",X"1A",X"2D",X"2C",X"7F",
		X"21",X"2C",X"2E",X"29",X"35",X"2C",X"2D",X"29",X"7F",X"50",X"50",X"50",X"7F",X"7F",X"7F",X"2C",
		X"2E",X"27",X"28",X"1B",X"7F",X"2D",X"2C",X"11",X"35",X"2C",X"2D",X"29",X"7F",X"50",X"50",X"50",
		X"7F",X"7F",X"7F",X"2C",X"2E",X"27",X"28",X"1B",X"7F",X"1D",X"27",X"12",X"35",X"2C",X"2D",X"29",
		X"7F",X"50",X"50",X"50",X"7F",X"7F",X"7F",X"32",X"2B",X"1E",X"2F",X"1E",X"7F",X"1D",X"27",X"1A",
		X"00",X"45",X"AB",X"C4",X"00",X"00",X"00",X"00",X"00",X"33",X"49",X"9D",X"C5",X"00",X"00",X"00",
		X"00",X"33",X"7C",X"A4",X"CD",X"00",X"00",X"00",X"00",X"53",X"6C",X"CD",X"94",X"3B",X"00",X"00",
		X"00",X"39",X"4D",X"73",X"B6",X"CB",X"00",X"00",X"00",X"A7",X"38",X"7B",X"C3",X"00",X"00",X"00",
		X"00",X"39",X"62",X"7D",X"BC",X"00",X"00",X"00",X"00",X"7D",X"A6",X"64",X"C8",X"00",X"00",X"00",
		X"00",X"4C",X"38",X"8A",X"82",X"C6",X"00",X"00",X"00",X"44",X"9C",X"C8",X"82",X"00",X"00",X"00",
		X"00",X"43",X"4B",X"B6",X"CC",X"00",X"00",X"00",X"00",X"49",X"92",X"8B",X"DA",X"00",X"00",X"00",
		X"00",X"42",X"CA",X"B3",X"39",X"00",X"00",X"00",X"00",X"5B",X"93",X"42",X"C9",X"00",X"00",X"00",
		X"00",X"62",X"C4",X"49",X"AA",X"00",X"00",X"00",X"46",X"83",X"54",X"81",X"00",X"00",X"00",X"00",
		X"86",X"80",X"56",X"82",X"00",X"00",X"00",X"00",X"54",X"83",X"00",X"00",X"00",X"00",X"00",X"00",
		X"94",X"81",X"88",X"80",X"98",X"80",X"CE",X"82",X"C8",X"81",X"54",X"82",X"00",X"00",X"00",X"00",
		X"1A",X"81",X"86",X"80",X"00",X"00",X"CC",X"82",X"D0",X"80",X"C8",X"81",X"00",X"00",X"00",X"00",
		X"48",X"82",X"56",X"82",X"5A",X"81",X"00",X"00",X"48",X"82",X"0E",X"81",X"46",X"81",X"00",X"00",
		X"94",X"82",X"C8",X"82",X"96",X"80",X"00",X"00",X"0C",X"83",X"00",X"00",X"00",X"00",X"00",X"00",
		X"D2",X"80",X"48",X"82",X"D4",X"82",X"D8",X"81",X"46",X"82",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C8",X"80",X"18",X"81",X"94",X"82",X"00",X"00",X"48",X"82",X"12",X"83",X"00",X"00",X"00",X"00",
		X"1A",X"82",X"C8",X"82",X"CA",X"80",X"D6",X"80",X"88",X"82",X"8C",X"80",X"00",X"00",X"00",X"00",
		X"98",X"80",X"0C",X"81",X"D8",X"82",X"D4",X"81",X"C6",X"80",X"4E",X"81",X"CC",X"82",X"00",X"00",
		X"D8",X"80",X"56",X"82",X"4A",X"81",X"00",X"00",X"8E",X"80",X"4A",X"81",X"14",X"83",X"00",X"00",
		X"4A",X"82",X"CE",X"82",X"00",X"00",X"00",X"00",X"8A",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"D6",X"80",X"4C",X"81",X"18",X"82",X"8A",X"82",X"CE",X"80",X"CC",X"82",X"00",X"00",X"00",X"00",
		X"C8",X"80",X"D6",X"81",X"9A",X"80",X"00",X"00",X"C8",X"82",X"8A",X"80",X"00",X"00",X"00",X"00",
		X"D2",X"80",X"48",X"81",X"56",X"82",X"00",X"00",X"D4",X"81",X"48",X"82",X"54",X"82",X"00",X"00",
		X"86",X"80",X"CE",X"80",X"D0",X"82",X"00",X"00",X"32",X"3C",X"DA",X"00",X"00",X"B4",X"00",X"00",
		X"A8",X"73",X"B2",X"00",X"00",X"00",X"4C",X"CC",X"58",X"63",X"B6",X"00",X"00",X"3C",X"DA",X"00",
		X"44",X"D9",X"58",X"00",X"00",X"8C",X"B5",X"00",X"4A",X"56",X"00",X"43",X"BC",X"8B",X"00",X"A4",
		X"45",X"45",X"00",X"00",X"73",X"9B",X"A3",X"C7",X"36",X"4B",X"46",X"A3",X"4C",X"A5",X"00",X"CB",
		X"56",X"56",X"5B",X"D6",X"00",X"BB",X"B3",X"43",X"7D",X"55",X"6A",X"6A",X"C3",X"C3",X"A7",X"CC",
		X"3C",X"59",X"CB",X"3C",X"59",X"74",X"7A",X"B5",X"73",X"73",X"7A",X"55",X"55",X"7D",X"B3",X"7A",
		X"6D",X"54",X"69",X"69",X"BB",X"BB",X"C6",X"54",X"4B",X"4B",X"7C",X"74",X"DB",X"B8",X"DB",X"B8",
		X"6D",X"54",X"49",X"49",X"9A",X"54",X"B5",X"B5",X"46",X"46",X"3C",X"7A",X"83",X"83",X"B6",X"B8",
		X"0C",X"14",X"0C",X"0F",X"11",X"0C",X"11",X"11",X"14",X"11",X"11",X"14",X"0C",X"0C",X"14",X"24",
		X"24",X"20",X"20",X"20",X"20",X"1C",X"1C",X"1C",X"1C",X"1A",X"1A",X"1A",X"18",X"18",X"1E",X"10",
		X"ED",X"73",X"85",X"89",X"32",X"88",X"89",X"3A",X"A7",X"85",X"32",X"87",X"89",X"11",X"82",X"89",
		X"06",X"03",X"7E",X"23",X"12",X"1B",X"10",X"FA",X"3E",X"01",X"32",X"3D",X"9B",X"3A",X"3D",X"9B",
		X"A7",X"20",X"FA",X"21",X"A0",X"89",X"06",X"05",X"11",X"80",X"89",X"0E",X"03",X"1A",X"96",X"38",
		X"14",X"20",X"07",X"23",X"13",X"0D",X"20",X"F5",X"18",X"0B",X"23",X"0D",X"20",X"FC",X"10",X"E8",
		X"CD",X"3B",X"35",X"06",X"00",X"04",X"78",X"32",X"C5",X"89",X"FE",X"06",X"20",X"05",X"ED",X"7B",
		X"85",X"89",X"C9",X"3E",X"05",X"90",X"28",X"1F",X"4F",X"06",X"00",X"21",X"C1",X"89",X"11",X"C0",
		X"89",X"87",X"81",X"ED",X"B0",X"21",X"A3",X"89",X"11",X"A0",X"89",X"4F",X"ED",X"B0",X"4F",X"21",
		X"B3",X"89",X"11",X"B0",X"89",X"ED",X"B0",X"4F",X"21",X"A0",X"89",X"06",X"00",X"09",X"EB",X"21",
		X"80",X"89",X"0E",X"03",X"ED",X"B0",X"21",X"B0",X"89",X"4F",X"09",X"06",X"03",X"36",X"37",X"23",
		X"10",X"FB",X"3A",X"C5",X"89",X"D6",X"05",X"ED",X"44",X"4F",X"21",X"C0",X"89",X"09",X"3A",X"88",
		X"89",X"77",X"21",X"A8",X"85",X"3A",X"00",X"84",X"F6",X"F9",X"3C",X"20",X"01",X"23",X"22",X"C7",
		X"89",X"CD",X"33",X"3E",X"21",X"2D",X"37",X"CD",X"F3",X"36",X"CD",X"F3",X"36",X"CD",X"F3",X"36",
		X"21",X"80",X"89",X"11",X"2F",X"83",X"01",X"00",X"03",X"CD",X"C6",X"36",X"06",X"05",X"CD",X"E9",
		X"36",X"10",X"FB",X"3A",X"88",X"89",X"0E",X"10",X"CD",X"61",X"36",X"21",X"2F",X"81",X"22",X"C9",
		X"89",X"AF",X"32",X"C6",X"89",X"21",X"28",X"F0",X"22",X"CD",X"89",X"CD",X"E7",X"35",X"CD",X"EE",
		X"34",X"3E",X"FF",X"32",X"94",X"9A",X"06",X"02",X"CD",X"DD",X"34",X"3A",X"23",X"84",X"4F",X"CD",
		X"EE",X"34",X"3A",X"23",X"84",X"B9",X"28",X"F7",X"E6",X"0F",X"CC",X"19",X"35",X"2A",X"C7",X"89",
		X"CB",X"66",X"CC",X"82",X"34",X"2A",X"C7",X"89",X"7E",X"E6",X"0E",X"21",X"84",X"89",X"BE",X"77",
		X"28",X"1A",X"FE",X"02",X"28",X"0F",X"FE",X"0C",X"28",X"0B",X"FE",X"06",X"20",X"CD",X"3E",X"FD",
		X"32",X"CB",X"89",X"18",X"3A",X"3E",X"FD",X"32",X"CC",X"89",X"18",X"0C",X"FE",X"06",X"28",X"2F",
		X"FE",X"0C",X"28",X"04",X"FE",X"02",X"20",X"B3",X"21",X"CC",X"89",X"34",X"20",X"AD",X"36",X"F0",
		X"3E",X"28",X"32",X"CD",X"89",X"2A",X"C9",X"89",X"34",X"7E",X"E6",X"3F",X"FE",X"34",X"38",X"05",
		X"FE",X"38",X"30",X"07",X"34",X"CD",X"E7",X"35",X"C3",X"EB",X"33",X"36",X"1A",X"18",X"F6",X"21",
		X"CB",X"89",X"34",X"20",X"F3",X"36",X"F0",X"3E",X"28",X"32",X"CD",X"89",X"2A",X"C9",X"89",X"35",
		X"7E",X"E6",X"3F",X"FE",X"19",X"28",X"07",X"FE",X"34",X"38",X"DA",X"35",X"18",X"D7",X"36",X"37",
		X"18",X"D3",X"2A",X"C9",X"89",X"CB",X"BE",X"4E",X"EB",X"CD",X"E9",X"36",X"ED",X"53",X"C9",X"89",
		X"3E",X"28",X"32",X"CD",X"89",X"3A",X"C6",X"89",X"5F",X"3C",X"32",X"C6",X"89",X"47",X"16",X"00",
		X"3A",X"C5",X"89",X"21",X"2F",X"35",X"CF",X"7E",X"23",X"66",X"6F",X"19",X"71",X"78",X"FE",X"03",
		X"C2",X"E7",X"35",X"ED",X"7B",X"85",X"89",X"CD",X"E7",X"35",X"CD",X"FC",X"34",X"3E",X"01",X"32",
		X"94",X"9A",X"06",X"04",X"CD",X"DD",X"34",X"3A",X"94",X"9A",X"A7",X"20",X"FA",X"3E",X"02",X"32",
		X"3D",X"9B",X"3A",X"3D",X"9B",X"A7",X"20",X"FA",X"ED",X"7B",X"85",X"89",X"C9",X"3A",X"23",X"84",
		X"E6",X"3F",X"20",X"F9",X"3A",X"23",X"84",X"E6",X"3F",X"28",X"F9",X"10",X"F0",X"C9",X"3A",X"A7",
		X"85",X"5F",X"3A",X"87",X"89",X"BB",X"C8",X"CD",X"82",X"34",X"18",X"FB",X"3A",X"A7",X"85",X"5F",
		X"3A",X"87",X"89",X"BB",X"C8",X"3A",X"94",X"9A",X"A7",X"28",X"C2",X"3E",X"01",X"32",X"94",X"9A",
		X"3A",X"94",X"9A",X"A7",X"28",X"FA",X"18",X"B5",X"C9",X"2A",X"C9",X"89",X"7E",X"EE",X"80",X"77",
		X"3A",X"23",X"84",X"E6",X"1F",X"C0",X"21",X"CD",X"89",X"35",X"28",X"CB",X"23",X"35",X"28",X"C7",
		X"C9",X"BC",X"89",X"B9",X"89",X"B6",X"89",X"B3",X"89",X"B0",X"89",X"CD",X"33",X"3E",X"21",X"77",
		X"37",X"CD",X"F3",X"36",X"CD",X"F3",X"36",X"CD",X"F3",X"36",X"CD",X"F3",X"36",X"3E",X"01",X"32",
		X"82",X"9A",X"3A",X"23",X"84",X"E6",X"1F",X"CC",X"75",X"35",X"E6",X"0F",X"CC",X"C9",X"35",X"3A",
		X"82",X"9A",X"A7",X"20",X"ED",X"CD",X"75",X"35",X"3A",X"23",X"84",X"C6",X"3C",X"4F",X"3A",X"23",
		X"84",X"B9",X"20",X"FA",X"C9",X"21",X"80",X"89",X"11",X"6D",X"83",X"06",X"03",X"AF",X"32",X"83",
		X"89",X"7E",X"1F",X"1F",X"1F",X"1F",X"CD",X"93",X"35",X"7E",X"CD",X"93",X"35",X"23",X"10",X"F1",
		X"3E",X"01",X"C9",X"E6",X"0F",X"20",X"0E",X"3A",X"83",X"89",X"A7",X"3E",X"00",X"20",X"06",X"CD",
		X"E9",X"36",X"C3",X"E9",X"36",X"E5",X"C5",X"21",X"CA",X"37",X"CF",X"7E",X"23",X"66",X"6F",X"01",
		X"FF",X"04",X"D5",X"ED",X"A0",X"ED",X"A0",X"ED",X"A0",X"ED",X"A0",X"D1",X"CD",X"E9",X"36",X"10",
		X"F1",X"C1",X"E1",X"3E",X"01",X"32",X"83",X"89",X"C9",X"11",X"6D",X"83",X"CD",X"D5",X"35",X"CD",
		X"D5",X"35",X"CD",X"D5",X"35",X"D5",X"06",X"18",X"3E",X"40",X"12",X"CD",X"E9",X"36",X"10",X"F8",
		X"D1",X"13",X"C9",X"AF",X"32",X"C5",X"89",X"21",X"63",X"37",X"CD",X"F3",X"36",X"11",X"5D",X"83",
		X"06",X"05",X"CD",X"F8",X"35",X"10",X"FB",X"C9",X"0E",X"00",X"3A",X"C5",X"89",X"B8",X"20",X"02",
		X"0E",X"40",X"78",X"21",X"8D",X"36",X"CF",X"7E",X"23",X"66",X"6F",X"D5",X"C5",X"06",X"03",X"7E",
		X"B1",X"12",X"23",X"CD",X"E9",X"36",X"10",X"F7",X"CD",X"E9",X"36",X"CD",X"E9",X"36",X"CD",X"45",
		X"36",X"06",X"04",X"CD",X"E9",X"36",X"10",X"FB",X"CD",X"64",X"36",X"CD",X"E9",X"36",X"CD",X"E9",
		X"36",X"7E",X"23",X"66",X"6F",X"06",X"03",X"7E",X"B1",X"12",X"CD",X"E9",X"36",X"23",X"10",X"F7",
		X"C1",X"D1",X"1B",X"1B",X"C9",X"7E",X"23",X"E5",X"66",X"6F",X"C5",X"D5",X"01",X"00",X"03",X"CD",
		X"C6",X"36",X"D1",X"C1",X"06",X"06",X"1A",X"B1",X"12",X"CD",X"E9",X"36",X"10",X"F8",X"E1",X"23",
		X"C9",X"E5",X"18",X"06",X"7E",X"23",X"E5",X"66",X"6F",X"7E",X"06",X"00",X"D6",X"0A",X"38",X"03",
		X"04",X"18",X"F9",X"F5",X"78",X"CD",X"81",X"36",X"F1",X"C6",X"0A",X"CD",X"87",X"36",X"E1",X"23",
		X"C9",X"E6",X"0F",X"20",X"02",X"3E",X"27",X"C6",X"10",X"B1",X"12",X"CD",X"E9",X"36",X"C9",X"99",
		X"36",X"A2",X"36",X"AB",X"36",X"B4",X"36",X"BD",X"36",X"11",X"2C",X"2D",X"AC",X"89",X"C4",X"89",
		X"BC",X"89",X"12",X"27",X"1D",X"A9",X"89",X"C3",X"89",X"B9",X"89",X"13",X"2B",X"1D",X"A6",X"89",
		X"C2",X"89",X"B6",X"89",X"14",X"2D",X"21",X"A3",X"89",X"C1",X"89",X"B3",X"89",X"15",X"2D",X"21",
		X"A0",X"89",X"C0",X"89",X"B0",X"89",X"7E",X"CD",X"CE",X"36",X"23",X"10",X"F9",X"C9",X"F5",X"1F",
		X"1F",X"1F",X"1F",X"CD",X"DC",X"36",X"F1",X"10",X"02",X"0E",X"FF",X"04",X"E6",X"0F",X"28",X"02",
		X"0E",X"FF",X"F6",X"10",X"A1",X"CC",X"F0",X"36",X"12",X"7B",X"D6",X"20",X"5F",X"D0",X"15",X"C9",
		X"3E",X"37",X"C9",X"4E",X"23",X"46",X"23",X"5E",X"23",X"56",X"23",X"7E",X"CD",X"0C",X"37",X"FE",
		X"FF",X"28",X"05",X"81",X"12",X"CD",X"E9",X"36",X"23",X"10",X"F0",X"C9",X"D6",X"30",X"FE",X"0A",
		X"D8",X"D6",X"07",X"FE",X"23",X"D8",X"C6",X"3E",X"FE",X"27",X"C8",X"C6",X"FC",X"FE",X"24",X"C8",
		X"C6",X"F4",X"FE",X"25",X"C8",X"C6",X"08",X"FE",X"26",X"C8",X"3E",X"FF",X"C9",X"50",X"15",X"2A",
		X"83",X"45",X"4E",X"54",X"45",X"52",X"20",X"59",X"4F",X"55",X"52",X"20",X"49",X"4E",X"49",X"54",
		X"49",X"41",X"4C",X"53",X"20",X"21",X"50",X"12",X"0D",X"83",X"53",X"43",X"4F",X"52",X"45",X"20",
		X"20",X"52",X"4F",X"55",X"4E",X"44",X"20",X"20",X"4E",X"41",X"4D",X"45",X"10",X"03",X"2F",X"81",
		X"41",X"41",X"41",X"10",X"10",X"93",X"82",X"53",X"43",X"4F",X"52",X"45",X"20",X"52",X"4F",X"55",
		X"4E",X"44",X"20",X"4E",X"41",X"4D",X"45",X"90",X"12",X"04",X"83",X"43",X"4F",X"4E",X"47",X"52",
		X"41",X"54",X"55",X"4C",X"41",X"54",X"49",X"4F",X"4E",X"53",X"20",X"21",X"21",X"50",X"15",X"27",
		X"83",X"20",X"20",X"20",X"48",X"49",X"47",X"48",X"45",X"53",X"54",X"20",X"53",X"43",X"4F",X"52",
		X"45",X"20",X"20",X"20",X"20",X"20",X"10",X"17",X"54",X"83",X"47",X"4F",X"20",X"46",X"4F",X"52",
		X"20",X"54",X"48",X"45",X"20",X"57",X"4F",X"52",X"4C",X"44",X"20",X"52",X"45",X"43",X"4F",X"52",
		X"44",X"10",X"05",X"56",X"82",X"4E",X"4F",X"57",X"20",X"21",X"DE",X"37",X"EE",X"37",X"FE",X"37",
		X"0E",X"38",X"1E",X"38",X"2E",X"38",X"3E",X"38",X"4E",X"38",X"5E",X"38",X"6E",X"38",X"40",X"48",
		X"4F",X"40",X"4B",X"46",X"42",X"4F",X"44",X"40",X"40",X"49",X"4D",X"41",X"45",X"40",X"40",X"40",
		X"40",X"40",X"4E",X"40",X"40",X"49",X"41",X"41",X"41",X"49",X"40",X"40",X"40",X"49",X"4E",X"40",
		X"4E",X"4F",X"45",X"4E",X"41",X"49",X"49",X"43",X"49",X"49",X"42",X"45",X"40",X"49",X"40",X"40",
		X"4E",X"40",X"49",X"4E",X"4D",X"49",X"44",X"41",X"40",X"49",X"45",X"4D",X"41",X"4C",X"40",X"4E",
		X"4F",X"40",X"4E",X"45",X"49",X"40",X"41",X"48",X"44",X"4F",X"46",X"46",X"45",X"4C",X"48",X"4F",
		X"4E",X"40",X"45",X"49",X"4D",X"49",X"49",X"49",X"40",X"49",X"4C",X"42",X"41",X"4C",X"40",X"48",
		X"48",X"40",X"43",X"42",X"46",X"49",X"49",X"47",X"40",X"49",X"4C",X"4D",X"41",X"4C",X"48",X"40",
		X"40",X"40",X"45",X"40",X"48",X"4F",X"49",X"43",X"46",X"4C",X"41",X"4C",X"40",X"40",X"4E",X"4F",
		X"48",X"40",X"45",X"41",X"40",X"49",X"49",X"47",X"49",X"49",X"4D",X"4C",X"41",X"4C",X"4E",X"4F",
		X"40",X"40",X"45",X"42",X"40",X"49",X"49",X"47",X"4E",X"49",X"42",X"41",X"45",X"40",X"F3",X"3E",
		X"10",X"32",X"00",X"71",X"AF",X"32",X"23",X"68",X"32",X"02",X"A0",X"32",X"20",X"68",X"3D",X"32",
		X"00",X"70",X"3E",X"04",X"32",X"40",X"B8",X"21",X"00",X"00",X"06",X"10",X"D9",X"21",X"00",X"80",
		X"01",X"00",X"04",X"54",X"5D",X"D9",X"54",X"5D",X"D9",X"D9",X"7C",X"AD",X"2F",X"87",X"87",X"ED",
		X"6A",X"7D",X"D9",X"77",X"23",X"32",X"30",X"68",X"0D",X"20",X"EE",X"10",X"EC",X"06",X"04",X"62",
		X"6B",X"D9",X"EB",X"D9",X"D9",X"7D",X"AC",X"2F",X"87",X"87",X"ED",X"6A",X"7D",X"D9",X"AE",X"C2",
		X"78",X"3D",X"23",X"32",X"30",X"68",X"0D",X"20",X"EB",X"10",X"E9",X"EB",X"D9",X"10",X"BD",X"D9",
		X"01",X"00",X"04",X"36",X"00",X"23",X"0D",X"20",X"FA",X"10",X"F8",X"31",X"00",X"84",X"21",X"E0",
		X"89",X"11",X"00",X"80",X"01",X"20",X"00",X"ED",X"B0",X"21",X"00",X"84",X"CD",X"E3",X"3D",X"21",
		X"00",X"88",X"CD",X"E3",X"3D",X"21",X"00",X"90",X"CD",X"E3",X"3D",X"21",X"00",X"98",X"CD",X"E3",
		X"3D",X"21",X"00",X"80",X"11",X"E0",X"89",X"01",X"20",X"00",X"ED",X"B0",X"31",X"00",X"9A",X"32",
		X"30",X"68",X"21",X"00",X"88",X"22",X"02",X"89",X"22",X"00",X"89",X"CD",X"3B",X"3E",X"21",X"95",
		X"3E",X"CD",X"F3",X"36",X"AF",X"32",X"00",X"8A",X"32",X"01",X"8A",X"3C",X"32",X"9A",X"87",X"32",
		X"22",X"68",X"32",X"25",X"68",X"32",X"26",X"68",X"32",X"27",X"68",X"32",X"23",X"68",X"11",X"FC",
		X"3F",X"21",X"00",X"00",X"01",X"00",X"10",X"AF",X"86",X"32",X"30",X"68",X"23",X"0D",X"20",X"F8",
		X"10",X"F6",X"EB",X"BE",X"C2",X"65",X"3E",X"06",X"10",X"EB",X"13",X"7C",X"FE",X"40",X"20",X"E7",
		X"32",X"30",X"68",X"3A",X"00",X"8A",X"A7",X"28",X"FA",X"3C",X"C2",X"6A",X"3E",X"32",X"30",X"68",
		X"3A",X"01",X"8A",X"A7",X"28",X"FA",X"3C",X"C2",X"6A",X"3E",X"21",X"9F",X"3E",X"CD",X"F3",X"36",
		X"AF",X"32",X"00",X"8A",X"32",X"01",X"8A",X"06",X"10",X"32",X"30",X"68",X"0D",X"20",X"FA",X"10",
		X"F8",X"21",X"E5",X"3F",X"11",X"00",X"70",X"01",X"03",X"00",X"D9",X"3E",X"A1",X"32",X"00",X"71",
		X"3A",X"00",X"71",X"FE",X"10",X"20",X"F9",X"21",X"EC",X"3F",X"11",X"18",X"8A",X"01",X"09",X"00",
		X"ED",X"B0",X"ED",X"56",X"AF",X"32",X"20",X"68",X"3C",X"32",X"20",X"68",X"FB",X"3A",X"23",X"84",
		X"C6",X"04",X"4F",X"3A",X"23",X"84",X"B9",X"20",X"FA",X"3E",X"04",X"32",X"3D",X"9B",X"3A",X"3D",
		X"9B",X"A7",X"20",X"FA",X"3A",X"23",X"84",X"4F",X"3A",X"23",X"84",X"B9",X"28",X"FA",X"CD",X"B8",
		X"3A",X"CD",X"85",X"3A",X"CD",X"F1",X"3A",X"CD",X"4A",X"3B",X"CD",X"C0",X"3B",X"CD",X"DE",X"3B",
		X"CD",X"EC",X"3B",X"CD",X"FC",X"3B",X"CD",X"47",X"3C",X"CD",X"B3",X"3C",X"3A",X"A7",X"85",X"87",
		X"30",X"D2",X"CD",X"85",X"3E",X"3A",X"23",X"84",X"C6",X"64",X"4F",X"3A",X"23",X"84",X"B9",X"20",
		X"FA",X"3A",X"A7",X"85",X"87",X"30",X"FA",X"3E",X"01",X"32",X"3D",X"9B",X"3A",X"3D",X"9B",X"A7",
		X"20",X"FA",X"F3",X"32",X"30",X"68",X"3A",X"00",X"71",X"FE",X"10",X"20",X"F6",X"01",X"00",X"08",
		X"32",X"30",X"68",X"0D",X"20",X"FA",X"10",X"F8",X"21",X"18",X"8A",X"11",X"00",X"70",X"01",X"09",
		X"00",X"D9",X"AF",X"32",X"00",X"70",X"3E",X"C1",X"32",X"00",X"71",X"3A",X"00",X"71",X"FE",X"10",
		X"20",X"F9",X"21",X"00",X"70",X"11",X"10",X"8A",X"01",X"03",X"00",X"D9",X"3E",X"B1",X"32",X"00",
		X"71",X"3A",X"00",X"71",X"FE",X"10",X"20",X"F9",X"3A",X"10",X"8A",X"A7",X"20",X"CA",X"FE",X"A0",
		X"20",X"00",X"C3",X"1C",X"01",X"21",X"CE",X"87",X"11",X"8A",X"89",X"7E",X"17",X"E6",X"0E",X"12",
		X"13",X"7E",X"1F",X"1F",X"E6",X"0E",X"12",X"7E",X"13",X"07",X"07",X"3C",X"E6",X"03",X"12",X"23",
		X"13",X"4E",X"CB",X"19",X"8F",X"CB",X"19",X"8F",X"E6",X"03",X"12",X"7E",X"13",X"E6",X"04",X"12",
		X"7E",X"07",X"07",X"E6",X"03",X"13",X"12",X"C9",X"21",X"8A",X"3F",X"3A",X"CF",X"89",X"A7",X"C4",
		X"F3",X"36",X"21",X"D9",X"89",X"11",X"D8",X"89",X"01",X"07",X"00",X"ED",X"B0",X"3A",X"A8",X"85",
		X"06",X"02",X"5A",X"2B",X"77",X"2B",X"B6",X"2B",X"2F",X"A6",X"2B",X"A6",X"77",X"57",X"3A",X"A7",
		X"85",X"10",X"EF",X"EB",X"29",X"06",X"0F",X"29",X"38",X"02",X"10",X"FB",X"78",X"32",X"88",X"89",
		X"C9",X"3A",X"8F",X"89",X"21",X"9C",X"3F",X"CF",X"E5",X"21",X"BF",X"3E",X"CD",X"F3",X"36",X"CD",
		X"F3",X"36",X"CD",X"F3",X"36",X"CD",X"F3",X"36",X"D1",X"21",X"48",X"83",X"01",X"1A",X"8A",X"CD",
		X"20",X"3B",X"3A",X"8A",X"89",X"21",X"A4",X"3F",X"D7",X"EB",X"21",X"4A",X"83",X"01",X"1C",X"8A",
		X"1A",X"77",X"02",X"03",X"C5",X"D6",X"11",X"3E",X"2C",X"20",X"02",X"3E",X"37",X"01",X"40",X"FF",
		X"09",X"77",X"3E",X"37",X"01",X"E0",X"FF",X"09",X"77",X"13",X"1A",X"09",X"77",X"C1",X"02",X"D6",
		X"11",X"3E",X"2C",X"20",X"02",X"3E",X"37",X"25",X"77",X"C9",X"3A",X"8B",X"89",X"A7",X"20",X"0F",
		X"21",X"FF",X"FF",X"22",X"D0",X"89",X"21",X"6F",X"3F",X"CD",X"F3",X"36",X"C3",X"AC",X"3B",X"21",
		X"B2",X"3F",X"4F",X"3A",X"8C",X"89",X"A7",X"20",X"03",X"21",X"C0",X"3F",X"06",X"00",X"09",X"E5",
		X"21",X"E7",X"3E",X"CD",X"F3",X"36",X"CD",X"F3",X"36",X"E1",X"7E",X"32",X"92",X"81",X"32",X"D0",
		X"89",X"23",X"7E",X"32",X"D1",X"89",X"FE",X"FF",X"28",X"22",X"F5",X"E6",X"1F",X"32",X"94",X"81",
		X"21",X"04",X"3F",X"CD",X"F3",X"36",X"CD",X"F3",X"36",X"F1",X"CB",X"7F",X"28",X"14",X"E6",X"1F",
		X"32",X"96",X"81",X"21",X"21",X"3F",X"CD",X"F3",X"36",X"C3",X"F3",X"36",X"21",X"54",X"83",X"CD",
		X"B5",X"3B",X"21",X"56",X"83",X"11",X"E0",X"FF",X"06",X"18",X"36",X"37",X"19",X"10",X"FB",X"C9",
		X"3A",X"8C",X"89",X"A7",X"20",X"02",X"3E",X"05",X"C6",X"10",X"32",X"6C",X"82",X"D6",X"11",X"3E",
		X"37",X"20",X"02",X"3E",X"37",X"32",X"4C",X"82",X"21",X"3E",X"3F",X"C3",X"F3",X"36",X"3A",X"8D",
		X"89",X"C6",X"1A",X"32",X"AE",X"82",X"21",X"48",X"3F",X"C3",X"F3",X"36",X"3A",X"8E",X"89",X"21",
		X"50",X"3F",X"A7",X"CA",X"F3",X"36",X"21",X"5B",X"3F",X"C3",X"F3",X"36",X"3A",X"89",X"89",X"0E",
		X"00",X"FE",X"0A",X"38",X"05",X"D6",X"0A",X"0C",X"18",X"F7",X"C6",X"10",X"32",X"70",X"82",X"79",
		X"C6",X"10",X"32",X"90",X"82",X"21",X"01",X"84",X"CB",X"EE",X"3A",X"88",X"89",X"A7",X"C4",X"27",
		X"3C",X"21",X"66",X"3F",X"C3",X"F3",X"36",X"3A",X"89",X"89",X"3C",X"FE",X"15",X"38",X"01",X"AF",
		X"32",X"89",X"89",X"21",X"80",X"9A",X"06",X"2C",X"36",X"00",X"23",X"10",X"FB",X"21",X"80",X"9A",
		X"4F",X"06",X"00",X"09",X"36",X"01",X"C9",X"2A",X"91",X"89",X"7C",X"B5",X"28",X"05",X"2B",X"22",
		X"91",X"89",X"C9",X"3A",X"88",X"89",X"FE",X"0F",X"28",X"0C",X"21",X"5A",X"83",X"C3",X"B5",X"3B",
		X"3E",X"03",X"32",X"3D",X"9B",X"C9",X"3A",X"A7",X"85",X"E6",X"01",X"28",X"F3",X"21",X"B0",X"04",
		X"22",X"91",X"89",X"21",X"E0",X"89",X"11",X"5A",X"83",X"01",X"02",X"01",X"CD",X"8B",X"3C",X"06",
		X"03",X"CD",X"8B",X"3C",X"06",X"02",X"CD",X"8B",X"3C",X"06",X"01",X"7E",X"CD",X"A0",X"3C",X"23",
		X"CD",X"97",X"3C",X"23",X"10",X"FA",X"C9",X"7E",X"1F",X"1F",X"1F",X"1F",X"CD",X"A0",X"3C",X"7E",
		X"E6",X"0F",X"2F",X"C6",X"1A",X"12",X"CD",X"E9",X"36",X"0D",X"C0",X"0E",X"04",X"3E",X"35",X"12",
		X"C3",X"E9",X"36",X"3A",X"A7",X"85",X"E6",X"03",X"28",X"02",X"3E",X"01",X"3C",X"32",X"07",X"A0",
		X"3A",X"A7",X"85",X"E6",X"01",X"28",X"05",X"AF",X"32",X"90",X"89",X"C9",X"3A",X"88",X"89",X"3D",
		X"FE",X"04",X"D0",X"3C",X"4F",X"3A",X"90",X"89",X"5F",X"3C",X"32",X"90",X"89",X"16",X"00",X"21",
		X"D0",X"3F",X"19",X"7E",X"3C",X"28",X"07",X"B9",X"C8",X"AF",X"32",X"90",X"89",X"C9",X"CD",X"3B",
		X"3E",X"11",X"24",X"3D",X"21",X"42",X"80",X"06",X"1C",X"CD",X"07",X"3D",X"10",X"FB",X"3A",X"A7",
		X"85",X"87",X"30",X"FA",X"C3",X"12",X"3A",X"CD",X"15",X"3D",X"CD",X"15",X"3D",X"CD",X"15",X"3D",
		X"3E",X"05",X"C3",X"10",X"00",X"1A",X"0E",X"08",X"87",X"30",X"02",X"36",X"18",X"23",X"0D",X"20",
		X"F7",X"13",X"23",X"C9",X"00",X"3E",X"00",X"31",X"41",X"00",X"49",X"41",X"00",X"45",X"41",X"00",
		X"23",X"3E",X"00",X"00",X"00",X"03",X"36",X"22",X"03",X"49",X"41",X"00",X"49",X"41",X"3E",X"36",
		X"3E",X"41",X"00",X"00",X"41",X"3E",X"7F",X"41",X"49",X"20",X"7F",X"49",X"18",X"00",X"32",X"20",
		X"40",X"00",X"7F",X"40",X"01",X"00",X"7F",X"7F",X"3F",X"40",X"21",X"44",X"40",X"00",X"44",X"00",
		X"3C",X"44",X"01",X"42",X"3F",X"01",X"81",X"00",X"01",X"A5",X"7F",X"01",X"A5",X"04",X"7F",X"99",
		X"08",X"00",X"42",X"10",X"00",X"3C",X"7F",X"00",X"E6",X"0F",X"1E",X"21",X"28",X"02",X"1E",X"25",
		X"7C",X"1F",X"1F",X"E6",X"07",X"FE",X"03",X"38",X"06",X"3D",X"FE",X"03",X"28",X"01",X"3D",X"21",
		X"00",X"80",X"01",X"00",X"04",X"36",X"37",X"32",X"30",X"68",X"23",X"0D",X"20",X"F7",X"10",X"F5",
		X"21",X"80",X"8B",X"01",X"80",X"00",X"36",X"00",X"23",X"10",X"FB",X"21",X"80",X"93",X"01",X"80",
		X"00",X"36",X"00",X"23",X"10",X"FB",X"21",X"80",X"9B",X"01",X"80",X"00",X"36",X"00",X"23",X"10",
		X"FB",X"C6",X"10",X"32",X"C2",X"82",X"7B",X"32",X"A2",X"82",X"3E",X"2B",X"32",X"42",X"83",X"3E",
		X"1A",X"32",X"22",X"83",X"3E",X"26",X"32",X"02",X"83",X"3E",X"01",X"32",X"03",X"A0",X"32",X"30",
		X"68",X"18",X"FE",X"D9",X"06",X"10",X"D9",X"01",X"00",X"04",X"54",X"5D",X"D9",X"54",X"5D",X"D9",
		X"D9",X"7C",X"AD",X"2F",X"87",X"87",X"ED",X"6A",X"7D",X"D9",X"77",X"23",X"32",X"30",X"68",X"0D",
		X"20",X"EE",X"10",X"EC",X"06",X"04",X"62",X"6B",X"D9",X"EB",X"D9",X"D9",X"7D",X"AC",X"2F",X"87",
		X"87",X"ED",X"6A",X"7D",X"D9",X"AE",X"C2",X"78",X"3D",X"23",X"32",X"30",X"68",X"0D",X"20",X"EB",
		X"10",X"E9",X"EB",X"D9",X"10",X"C0",X"D9",X"01",X"00",X"04",X"36",X"00",X"23",X"0D",X"20",X"FA",
		X"10",X"F8",X"C9",X"21",X"40",X"80",X"01",X"C0",X"04",X"18",X"06",X"21",X"00",X"80",X"01",X"00",
		X"04",X"36",X"37",X"23",X"0D",X"20",X"FA",X"10",X"F8",X"3E",X"01",X"32",X"03",X"A0",X"21",X"80",
		X"8B",X"CD",X"5D",X"3E",X"21",X"80",X"93",X"CD",X"5D",X"3E",X"21",X"80",X"9B",X"06",X"80",X"AF",
		X"77",X"23",X"10",X"FC",X"C9",X"7A",X"1F",X"1F",X"1F",X"1F",X"E6",X"0F",X"F6",X"10",X"32",X"C4",
		X"82",X"3E",X"2B",X"32",X"44",X"83",X"3E",X"28",X"32",X"24",X"83",X"3E",X"26",X"32",X"04",X"83",
		X"32",X"30",X"68",X"18",X"FB",X"CD",X"3B",X"3E",X"21",X"00",X"A0",X"36",X"01",X"06",X"03",X"23",
		X"36",X"00",X"10",X"FB",X"C9",X"10",X"06",X"42",X"83",X"52",X"41",X"4D",X"20",X"4F",X"4B",X"10",
		X"06",X"44",X"83",X"52",X"4F",X"4D",X"20",X"4F",X"4B",X"10",X"12",X"48",X"83",X"46",X"52",X"45",
		X"45",X"20",X"50",X"4C",X"41",X"59",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"10",
		X"05",X"28",X"83",X"20",X"43",X"4F",X"49",X"4E",X"10",X"07",X"28",X"82",X"20",X"43",X"52",X"45",
		X"44",X"49",X"54",X"10",X"05",X"2A",X"83",X"20",X"43",X"4F",X"49",X"4E",X"10",X"07",X"2A",X"82",
		X"20",X"43",X"52",X"45",X"44",X"49",X"54",X"10",X"0D",X"52",X"83",X"31",X"53",X"54",X"20",X"42",
		X"4F",X"4E",X"55",X"53",X"20",X"46",X"4F",X"52",X"10",X"08",X"72",X"81",X"30",X"30",X"30",X"30",
		X"20",X"50",X"54",X"53",X"10",X"0D",X"54",X"83",X"32",X"4E",X"44",X"20",X"42",X"4F",X"4E",X"55",
		X"53",X"20",X"46",X"4F",X"52",X"10",X"08",X"74",X"81",X"30",X"30",X"30",X"30",X"20",X"50",X"54",
		X"53",X"10",X"0D",X"56",X"83",X"41",X"4E",X"44",X"20",X"46",X"4F",X"52",X"20",X"45",X"56",X"45",
		X"52",X"59",X"10",X"08",X"76",X"81",X"30",X"30",X"30",X"30",X"20",X"50",X"54",X"53",X"10",X"06",
		X"4C",X"83",X"44",X"49",X"47",X"44",X"55",X"47",X"10",X"04",X"4E",X"83",X"52",X"41",X"4E",X"4B",
		X"10",X"07",X"46",X"83",X"54",X"41",X"42",X"4C",X"45",X"20",X"20",X"10",X"07",X"46",X"83",X"55",
		X"50",X"52",X"49",X"47",X"48",X"54",X"10",X"05",X"50",X"83",X"53",X"4F",X"55",X"4E",X"44",X"10",
		X"17",X"52",X"83",X"42",X"4F",X"4E",X"55",X"53",X"20",X"4E",X"4F",X"54",X"48",X"49",X"4E",X"47",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"10",X"0E",X"58",X"83",X"42",X"41",
		X"43",X"4B",X"55",X"50",X"20",X"4E",X"4F",X"54",X"48",X"49",X"4E",X"47",X"11",X"11",X"12",X"11",
		X"11",X"12",X"12",X"13",X"11",X"17",X"11",X"11",X"11",X"13",X"12",X"11",X"11",X"16",X"12",X"13",
		X"11",X"12",X"13",X"11",X"12",X"97",X"11",X"95",X"12",X"16",X"11",X"94",X"11",X"14",X"12",X"96",
		X"11",X"FF",X"12",X"16",X"13",X"98",X"12",X"FF",X"12",X"96",X"13",X"17",X"12",X"15",X"13",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"02",X"02",X"02",X"02",X"03",X"03",X"03",
		X"03",X"03",X"03",X"03",X"FF",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"00",X"01",X"01",X"01",
		X"01",X"01",X"04",X"02",X"02",X"02",X"02",X"FF",X"FF",X"FF",X"FF",X"67",X"24",X"52",X"86",X"AA");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
