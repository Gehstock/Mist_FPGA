library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity cclimber_big_sprite_tile_bit0 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of cclimber_big_sprite_tile_bit0 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"00",X"00",X"00",X"1F",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"60",X"FE",X"FE",X"FE",X"FE",X"FE",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"FF",X"FF",
		X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"1F",X"00",X"00",X"00",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"60",X"00",X"00",X"FF",X"FF",X"F0",X"F0",X"F0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"03",X"03",X"01",X"01",X"01",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"F8",X"FC",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"7F",X"3F",X"3F",X"07",X"03",X"01",X"00",
		X"FF",X"FE",X"FE",X"FE",X"FC",X"F9",X"F9",X"1B",X"7C",X"7C",X"7C",X"FE",X"FF",X"FF",X"FF",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C2",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",
		X"00",X"80",X"C0",X"E0",X"F0",X"FC",X"FC",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"3F",X"1F",X"0F",X"07",X"07",X"01",X"00",
		X"FF",X"FF",X"FE",X"FC",X"F9",X"F3",X"E7",X"CF",X"00",X"00",X"40",X"E0",X"F0",X"E0",X"C0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"3F",X"1D",X"08",X"00",X"00",X"00",X"00",X"F0",X"F8",X"F0",X"E0",X"40",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"80",X"C0",X"F0",X"F0",X"F0",X"F8",X"FC",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"1F",X"1F",X"1F",X"1F",X"0F",X"07",X"07",
		X"FE",X"FE",X"FE",X"FF",X"FF",X"F8",X"F1",X"87",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"01",X"01",X"00",X"00",X"00",X"00",
		X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"0E",X"C0",X"C0",X"00",X"00",X"00",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",
		X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"3F",X"3F",X"1F",X"1F",X"1F",X"1F",X"00",
		X"F8",X"FC",X"FC",X"F8",X"F8",X"F8",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"1F",X"1F",X"1F",X"03",X"03",X"03",X"03",
		X"F8",X"F8",X"F8",X"F8",X"C0",X"C0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",
		X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"02",X"0C",X"08",X"08",X"10",X"20",X"20",X"0F",X"0F",X"0F",X"1F",X"1F",X"1F",X"9F",X"1F",
		X"F0",X"F0",X"F1",X"F8",X"F8",X"F8",X"F8",X"F8",X"60",X"10",X"08",X"C8",X"44",X"42",X"42",X"30",
		X"04",X"08",X"10",X"10",X"10",X"20",X"18",X"07",X"1F",X"3F",X"3F",X"1F",X"1D",X"18",X"00",X"00",
		X"F8",X"FC",X"FC",X"F8",X"F8",X"78",X"00",X"00",X"08",X"0C",X"04",X"04",X"04",X"08",X"10",X"70",
		X"10",X"10",X"0C",X"03",X"00",X"00",X"00",X"00",X"C3",X"3C",X"00",X"0A",X"F5",X"00",X"00",X"00",
		X"E3",X"1C",X"00",X"00",X"01",X"E2",X"00",X"00",X"80",X"00",X"10",X"20",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"02",X"1E",X"20",X"00",X"00",X"01",X"00",X"E0",X"00",X"00",X"18",
		X"00",X"00",X"C1",X"20",X"00",X"78",X"04",X"02",X"00",X"00",X"C0",X"20",X"20",X"40",X"30",X"0C",
		X"20",X"00",X"05",X"04",X"08",X"08",X"08",X"10",X"20",X"C0",X"00",X"00",X"00",X"01",X"03",X"07",
		X"01",X"01",X"00",X"02",X"01",X"80",X"C0",X"E0",X"04",X"E0",X"10",X"10",X"08",X"88",X"88",X"80",
		X"08",X"10",X"10",X"20",X"10",X"00",X"00",X"20",X"0F",X"0F",X"0F",X"1F",X"1F",X"1F",X"0C",X"00",
		X"F0",X"F0",X"F0",X"F8",X"F8",X"08",X"00",X"00",X"40",X"20",X"40",X"00",X"0C",X"04",X"04",X"3C",
		X"12",X"11",X"10",X"18",X"04",X"02",X"01",X"00",X"00",X"00",X"C0",X"38",X"07",X"00",X"00",X"00",
		X"0E",X"30",X"00",X"23",X"C0",X"00",X"00",X"00",X"20",X"20",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"0C",X"1E",X"00",X"00",X"2E",X"FF",X"3E",X"F8",X"99",X"A7",
		X"00",X"00",X"30",X"AE",X"31",X"08",X"88",X"F8",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"20",
		X"1E",X"1C",X"28",X"20",X"33",X"24",X"07",X"0F",X"43",X"07",X"7F",X"85",X"0E",X"0E",X"A1",X"BE",
		X"FC",X"FC",X"F0",X"F1",X"59",X"47",X"C1",X"30",X"30",X"70",X"F8",X"F8",X"E0",X"E0",X"E0",X"B0",
		X"0F",X"0F",X"25",X"25",X"12",X"10",X"10",X"13",X"21",X"D9",X"23",X"3E",X"E1",X"C1",X"43",X"2F",
		X"08",X"08",X"3F",X"DE",X"5F",X"1F",X"9F",X"F7",X"A8",X"98",X"10",X"10",X"20",X"88",X"8C",X"8C",
		X"0B",X"0B",X"09",X"04",X"02",X"00",X"00",X"00",X"13",X"C9",X"E1",X"F9",X"47",X"20",X"3E",X"00",
		X"F0",X"F8",X"F9",X"3B",X"03",X"FE",X"00",X"00",X"14",X"3C",X"F0",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"81",X"41",X"21",X"40",X"40",X"80",X"80",X"98",X"04",X"02",X"02",X"81",X"41",X"21",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"20",X"10",X"00",X"00",X"00",X"00",X"00",X"10",X"20",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"04",X"08",X"04",X"08",X"08",
		X"00",X"00",X"20",X"10",X"10",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"01",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"04",X"08",X"10",X"10",X"20",X"00",X"00",X"00",X"20",X"10",X"08",X"08",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"42",X"42",X"84",X"84",X"82",X"00",X"00",X"00",X"42",X"42",X"21",X"21",X"41",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"04",X"08",X"04",X"08",X"08",
		X"00",X"00",X"00",X"20",X"10",X"08",X"08",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"01",X"00",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"81",X"41",X"21",X"40",X"40",X"80",X"40",X"98",X"04",X"02",X"02",X"81",X"41",X"21",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"20",X"10",X"00",X"00",X"00",X"00",X"00",X"10",X"20",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"08",X"10",X"08",X"04",X"04",X"04",X"02",X"00",X"00",X"20",X"10",X"10",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"84",X"82",X"81",X"80",X"40",X"40",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"41",X"21",X"11",X"80",X"40",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"14",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"28",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"08",X"10",X"20",X"20",X"00",X"00",X"00",X"10",X"10",X"08",X"04",X"04",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"84",X"82",X"81",X"80",X"40",X"40",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"41",X"21",X"11",X"80",X"40",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"08",X"10",X"08",X"04",X"04",X"04",X"02",X"00",X"00",X"20",X"10",X"10",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
