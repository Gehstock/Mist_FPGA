library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity gravitar_pgm_rom5 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of gravitar_pgm_rom5 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"29",X"01",X"D0",X"05",X"A0",X"10",X"4C",X"0B",X"D0",X"A0",X"12",X"84",X"22",X"20",X"C2",X"CF",
		X"C6",X"22",X"4C",X"C2",X"CF",X"58",X"3D",X"5C",X"3D",X"64",X"3D",X"6C",X"3D",X"74",X"3D",X"7C",
		X"3D",X"84",X"3D",X"5E",X"3E",X"62",X"3E",X"B2",X"3E",X"B6",X"3E",X"BA",X"3E",X"BE",X"3E",X"1E",
		X"3F",X"24",X"3F",X"EE",X"3F",X"F8",X"3F",X"DA",X"40",X"DE",X"40",X"E2",X"40",X"6A",X"41",X"6E",
		X"41",X"72",X"41",X"2A",X"42",X"30",X"42",X"32",X"42",X"3A",X"42",X"D0",X"42",X"DA",X"42",X"E4",
		X"42",X"F0",X"40",X"F4",X"40",X"F8",X"40",X"D2",X"43",X"D6",X"43",X"DC",X"43",X"E4",X"43",X"E8",
		X"43",X"EE",X"43",X"F6",X"43",X"2A",X"44",X"E2",X"44",X"E8",X"44",X"40",X"45",X"48",X"45",X"52",
		X"45",X"E2",X"3D",X"E8",X"3D",X"EE",X"3D",X"F6",X"3D",X"02",X"3E",X"0E",X"3E",X"00",X"01",X"02",
		X"03",X"04",X"05",X"06",X"F9",X"07",X"07",X"08",X"08",X"FC",X"09",X"0A",X"0B",X"0C",X"FC",X"0D",
		X"0E",X"FE",X"0F",X"0F",X"10",X"10",X"FC",X"11",X"12",X"13",X"FD",X"14",X"14",X"14",X"15",X"15",
		X"FB",X"16",X"FF",X"17",X"18",X"19",X"1A",X"FC",X"1B",X"1C",X"1D",X"FD",X"1E",X"1F",X"20",X"FD",
		X"21",X"22",X"23",X"24",X"25",X"26",X"FA",X"27",X"27",X"28",X"28",X"FC",X"29",X"2A",X"FE",X"2B",
		X"2C",X"2D",X"FD",X"2E",X"2F",X"30",X"FD",X"31",X"32",X"33",X"FD",X"15",X"08",X"0D",X"12",X"1A",
		X"2B",X"1E",X"26",X"24",X"2F",X"42",X"3A",X"3F",X"33",X"1A",X"00",X"46",X"00",X"4A",X"01",X"0F",
		X"03",X"0F",X"07",X"03",X"0F",X"07",X"07",X"03",X"07",X"05",X"07",X"07",X"07",X"03",X"07",X"01",
		X"03",X"A2",X"0F",X"86",X"21",X"20",X"66",X"E4",X"A6",X"21",X"BD",X"CE",X"03",X"85",X"06",X"BD",
		X"DE",X"03",X"85",X"07",X"BD",X"EE",X"03",X"85",X"04",X"BD",X"FE",X"03",X"85",X"05",X"A9",X"00",
		X"85",X"0A",X"A2",X"04",X"20",X"A9",X"E4",X"20",X"8D",X"D9",X"A6",X"21",X"BD",X"0E",X"04",X"48",
		X"38",X"E9",X"04",X"9D",X"0E",X"04",X"68",X"20",X"86",X"E4",X"C6",X"21",X"10",X"C7",X"60",X"A5",
		X"50",X"D0",X"33",X"A5",X"4F",X"29",X"0F",X"AA",X"AD",X"0A",X"60",X"9D",X"CE",X"03",X"AD",X"0A",
		X"60",X"29",X"03",X"18",X"69",X"FE",X"9D",X"DE",X"03",X"AD",X"0A",X"60",X"9D",X"EE",X"03",X"AD",
		X"0A",X"60",X"29",X"03",X"18",X"69",X"FE",X"9D",X"FE",X"03",X"A9",X"C0",X"9D",X"0E",X"04",X"A9",
		X"02",X"85",X"50",X"4C",X"68",X"D1",X"C6",X"50",X"60",X"20",X"76",X"D9",X"A2",X"0E",X"86",X"21",
		X"BD",X"EC",X"02",X"F0",X"30",X"20",X"66",X"E4",X"A6",X"21",X"BD",X"4D",X"02",X"85",X"05",X"BD",
		X"64",X"02",X"85",X"04",X"BD",X"1F",X"02",X"85",X"06",X"BD",X"08",X"02",X"85",X"07",X"A9",X"00",
		X"85",X"0A",X"A2",X"04",X"20",X"A9",X"E4",X"A5",X"21",X"C9",X"04",X"B0",X"03",X"20",X"82",X"D9",
		X"A9",X"E0",X"20",X"86",X"E4",X"C6",X"21",X"A6",X"21",X"10",X"C5",X"60",X"A6",X"CF",X"B5",X"88",
		X"F0",X"0C",X"20",X"BF",X"D1",X"20",X"6E",X"D9",X"20",X"D5",X"D1",X"20",X"E4",X"D1",X"60",X"20",
		X"66",X"E4",X"A2",X"03",X"B5",X"0D",X"95",X"04",X"CA",X"10",X"F9",X"A2",X"04",X"A9",X"00",X"85",
		X"0A",X"20",X"A9",X"E4",X"60",X"A5",X"11",X"29",X"FE",X"A8",X"B9",X"C7",X"45",X"BE",X"C6",X"45",
		X"20",X"56",X"D9",X"60",X"A5",X"4C",X"F0",X"06",X"20",X"76",X"D9",X"4C",X"F1",X"D1",X"20",X"6A",
		X"D9",X"A5",X"11",X"29",X"FE",X"A8",X"BE",X"26",X"4A",X"B9",X"27",X"4A",X"20",X"53",X"E4",X"A5",
		X"4B",X"F0",X"2A",X"A6",X"CF",X"B4",X"4D",X"B9",X"31",X"C1",X"C9",X"A8",X"F0",X"1F",X"20",X"72",
		X"D9",X"20",X"BF",X"D1",X"A4",X"CF",X"B6",X"4D",X"A0",X"00",X"E0",X"03",X"D0",X"06",X"A5",X"10",
		X"10",X"02",X"A0",X"02",X"BE",X"66",X"4A",X"B9",X"67",X"4A",X"20",X"53",X"E4",X"60",X"20",X"8D",
		X"D9",X"A5",X"D0",X"F0",X"1C",X"A6",X"CF",X"B5",X"88",X"F0",X"13",X"A5",X"1D",X"29",X"01",X"F0",
		X"0D",X"20",X"D7",X"E0",X"20",X"BF",X"D1",X"A9",X"45",X"A2",X"B4",X"20",X"53",X"E4",X"4C",X"55",
		X"D2",X"A5",X"4B",X"D0",X"EF",X"AD",X"6E",X"04",X"F0",X"73",X"A6",X"CF",X"B5",X"88",X"F0",X"6D",
		X"20",X"8D",X"D9",X"A9",X"07",X"85",X"21",X"20",X"66",X"E4",X"AD",X"0A",X"60",X"29",X"3F",X"85",
		X"22",X"AD",X"0A",X"60",X"29",X"0F",X"85",X"23",X"A5",X"0F",X"A6",X"CF",X"B4",X"4D",X"C0",X"03",
		X"D0",X"10",X"24",X"10",X"10",X"0C",X"18",X"65",X"22",X"85",X"06",X"A5",X"10",X"69",X"00",X"4C",
		X"9B",X"D2",X"38",X"E5",X"22",X"85",X"06",X"A5",X"10",X"E9",X"00",X"85",X"07",X"A5",X"0D",X"2C",
		X"0A",X"60",X"10",X"0C",X"38",X"E5",X"23",X"85",X"04",X"A5",X"0E",X"E9",X"00",X"4C",X"B9",X"D2",
		X"18",X"65",X"23",X"85",X"04",X"A5",X"0E",X"69",X"00",X"85",X"05",X"A9",X"00",X"85",X"0A",X"A2",
		X"04",X"20",X"A9",X"E4",X"A9",X"E0",X"20",X"86",X"E4",X"C6",X"21",X"10",X"9A",X"60",X"20",X"66",
		X"E4",X"A9",X"00",X"38",X"E5",X"2D",X"85",X"31",X"D0",X"01",X"38",X"A9",X"F8",X"E9",X"00",X"85",
		X"32",X"A5",X"2B",X"0A",X"A8",X"84",X"21",X"98",X"85",X"22",X"A5",X"66",X"71",X"62",X"85",X"33",
		X"A5",X"67",X"C8",X"71",X"62",X"88",X"85",X"34",X"A6",X"CF",X"B5",X"88",X"F0",X"0C",X"B5",X"F6",
		X"29",X"08",X"F0",X"06",X"20",X"6A",X"D9",X"4C",X"0D",X"D3",X"20",X"72",X"D9",X"A5",X"30",X"D0",
		X"0F",X"A5",X"21",X"38",X"E5",X"22",X"29",X"1F",X"C9",X"06",X"90",X"2C",X"C9",X"1C",X"B0",X"28",
		X"A9",X"00",X"85",X"0A",X"A2",X"03",X"B5",X"31",X"95",X"04",X"CA",X"10",X"F9",X"A2",X"04",X"20",
		X"A9",X"E4",X"A4",X"21",X"B1",X"64",X"AA",X"C8",X"B1",X"64",X"F0",X"09",X"20",X"53",X"E4",X"20",
		X"5A",X"D6",X"20",X"B4",X"D6",X"20",X"66",X"E4",X"A4",X"21",X"E6",X"32",X"A5",X"33",X"18",X"71",
		X"5C",X"85",X"33",X"A5",X"34",X"C8",X"71",X"5C",X"88",X"85",X"34",X"C8",X"C8",X"98",X"29",X"1F",
		X"85",X"21",X"C5",X"22",X"D0",X"92",X"4C",X"62",X"D8",X"00",X"00",X"00",X"FF",X"00",X"FF",X"E0",
		X"00",X"A0",X"FF",X"C0",X"FE",X"C0",X"FE",X"80",X"00",X"C0",X"FF",X"C0",X"FF",X"80",X"00",X"00",
		X"00",X"E0",X"FE",X"E0",X"FE",X"E0",X"FE",X"00",X"01",X"00",X"00",X"80",X"FE",X"A0",X"FD",X"A0",
		X"FD",X"00",X"FE",X"E0",X"FE",X"C0",X"FD",X"00",X"FE",X"00",X"00",X"80",X"FE",X"40",X"FE",X"C0",
		X"FD",X"40",X"FE",X"00",X"00",X"60",X"FE",X"A0",X"FE",X"00",X"00",X"80",X"00",X"40",X"00",X"60",
		X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"C0",X"00",X"C0",X"00",X"40",X"00",X"80",
		X"00",X"20",X"00",X"40",X"00",X"40",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"FE",X"00",X"FE",X"00",X"FF",X"00",
		X"FF",X"00",X"00",X"00",X"FF",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"01",X"00",X"FE",X"00",X"FE",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"02",X"80",
		X"03",X"80",X"05",X"40",X"01",X"40",X"01",X"80",X"FF",X"80",X"FF",X"80",X"00",X"80",X"00",X"80",
		X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"00",X"00",X"00",X"FF",X"00",X"FD",X"00",
		X"FD",X"00",X"FD",X"00",X"FD",X"00",X"FD",X"C0",X"FD",X"C0",X"FD",X"80",X"FE",X"80",X"FE",X"80",
		X"FD",X"80",X"FD",X"40",X"FC",X"C0",X"FC",X"C0",X"FD",X"58",X"38",X"E2",X"39",X"C2",X"39",X"02",
		X"39",X"38",X"3A",X"E4",X"38",X"52",X"3A",X"22",X"39",X"6A",X"38",X"F4",X"39",X"D4",X"39",X"14",
		X"39",X"46",X"3A",X"F4",X"38",X"64",X"3A",X"34",X"39",X"82",X"39",X"A2",X"39",X"42",X"39",X"42",
		X"39",X"C2",X"39",X"42",X"39",X"E2",X"39",X"42",X"39",X"94",X"39",X"B4",X"39",X"54",X"39",X"54",
		X"39",X"D4",X"39",X"54",X"39",X"F4",X"39",X"54",X"39",X"42",X"39",X"62",X"39",X"42",X"39",X"62",
		X"39",X"42",X"39",X"62",X"39",X"42",X"39",X"62",X"39",X"54",X"39",X"74",X"39",X"54",X"39",X"74",
		X"39",X"54",X"39",X"74",X"39",X"54",X"39",X"74",X"39",X"A2",X"39",X"E2",X"39",X"82",X"39",X"E2",
		X"39",X"E2",X"39",X"82",X"39",X"62",X"39",X"82",X"39",X"B4",X"39",X"F4",X"39",X"94",X"39",X"F4",
		X"39",X"F4",X"39",X"94",X"39",X"74",X"39",X"94",X"39",X"C2",X"39",X"82",X"39",X"C2",X"39",X"62",
		X"39",X"C2",X"39",X"42",X"39",X"E2",X"39",X"E2",X"39",X"D4",X"39",X"94",X"39",X"D4",X"39",X"74",
		X"39",X"D4",X"39",X"54",X"39",X"F4",X"39",X"F4",X"39",X"C2",X"39",X"62",X"39",X"C2",X"39",X"C2",
		X"39",X"A2",X"39",X"A2",X"39",X"C2",X"39",X"62",X"39",X"D4",X"39",X"74",X"39",X"D4",X"39",X"D4",
		X"39",X"B4",X"39",X"B4",X"39",X"D4",X"39",X"74",X"39",X"82",X"39",X"C2",X"39",X"A2",X"39",X"E2",
		X"39",X"C2",X"39",X"62",X"39",X"E2",X"39",X"82",X"39",X"94",X"39",X"D4",X"39",X"B4",X"39",X"F4",
		X"39",X"D4",X"39",X"74",X"39",X"F4",X"39",X"94",X"39",X"78",X"38",X"20",X"3A",X"A8",X"38",X"90",
		X"38",X"E2",X"39",X"82",X"39",X"C2",X"39",X"E2",X"39",X"84",X"38",X"2C",X"3A",X"B6",X"38",X"9C",
		X"38",X"F4",X"39",X"94",X"39",X"D4",X"39",X"F4",X"39",X"82",X"39",X"82",X"39",X"E2",X"39",X"C2",
		X"39",X"A2",X"39",X"A2",X"39",X"C2",X"39",X"A2",X"39",X"94",X"39",X"94",X"39",X"F4",X"39",X"D4",
		X"39",X"B4",X"39",X"B4",X"39",X"D4",X"39",X"B4",X"39",X"E2",X"39",X"62",X"39",X"82",X"39",X"E2",
		X"39",X"82",X"39",X"82",X"39",X"E2",X"39",X"E2",X"39",X"F4",X"39",X"74",X"39",X"94",X"39",X"F4",
		X"39",X"94",X"39",X"94",X"39",X"F4",X"39",X"F4",X"39",X"C4",X"38",X"C2",X"39",X"02",X"3A",X"A2",
		X"39",X"C2",X"39",X"C4",X"38",X"C4",X"38",X"E2",X"39",X"D6",X"38",X"D4",X"39",X"12",X"3A",X"B4",
		X"39",X"D4",X"39",X"D6",X"38",X"D6",X"38",X"F4",X"39",X"82",X"39",X"E2",X"39",X"E2",X"39",X"A2",
		X"39",X"E2",X"39",X"E2",X"39",X"C2",X"39",X"E2",X"39",X"94",X"39",X"F4",X"39",X"F4",X"39",X"B4",
		X"39",X"F4",X"39",X"F4",X"39",X"D4",X"39",X"F4",X"39",X"00",X"01",X"02",X"03",X"04",X"00",X"05",
		X"00",X"00",X"06",X"00",X"00",X"07",X"00",X"08",X"00",X"01",X"00",X"00",X"02",X"03",X"00",X"04",
		X"00",X"00",X"00",X"05",X"06",X"07",X"00",X"08",X"00",X"00",X"01",X"00",X"02",X"00",X"03",X"00",
		X"04",X"00",X"05",X"00",X"06",X"00",X"07",X"00",X"08",X"00",X"00",X"00",X"00",X"01",X"02",X"03",
		X"04",X"05",X"06",X"07",X"08",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"02",X"00",X"03",
		X"04",X"00",X"05",X"00",X"06",X"07",X"00",X"00",X"08",X"00",X"01",X"02",X"00",X"03",X"04",X"05",
		X"06",X"00",X"00",X"00",X"07",X"00",X"08",X"00",X"00",X"00",X"01",X"02",X"00",X"03",X"04",X"00",
		X"00",X"05",X"00",X"06",X"07",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"03",X"04",
		X"00",X"05",X"06",X"07",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"03",X"04",
		X"05",X"06",X"00",X"07",X"00",X"08",X"00",X"00",X"00",X"7A",X"20",X"66",X"E4",X"A5",X"21",X"4A",
		X"A8",X"B1",X"6E",X"F0",X"4C",X"A8",X"88",X"84",X"24",X"B9",X"E4",X"02",X"F0",X"43",X"B9",X"17",
		X"02",X"85",X"06",X"B9",X"00",X"02",X"85",X"07",X"B9",X"5C",X"02",X"85",X"04",X"B9",X"45",X"02",
		X"85",X"05",X"A9",X"00",X"85",X"0A",X"A2",X"04",X"20",X"A9",X"E4",X"20",X"76",X"D9",X"A4",X"24",
		X"B9",X"8F",X"04",X"F0",X"09",X"38",X"E9",X"01",X"99",X"8F",X"04",X"4C",X"A4",X"D6",X"98",X"18",
		X"69",X"08",X"85",X"24",X"A5",X"24",X"0A",X"A8",X"B1",X"6C",X"AA",X"C8",X"B1",X"6C",X"20",X"53",
		X"E4",X"A4",X"21",X"60",X"20",X"66",X"E4",X"20",X"6E",X"D9",X"A5",X"21",X"4A",X"A8",X"A9",X"00",
		X"85",X"39",X"B9",X"FB",X"02",X"F0",X"5A",X"A5",X"31",X"18",X"71",X"6A",X"85",X"04",X"A5",X"32",
		X"85",X"05",X"90",X"02",X"E6",X"05",X"B1",X"68",X"85",X"38",X"A2",X"03",X"06",X"38",X"26",X"39",
		X"CA",X"10",X"F9",X"A5",X"39",X"C9",X"08",X"90",X"02",X"09",X"F0",X"85",X"39",X"A5",X"33",X"18",
		X"65",X"38",X"85",X"06",X"A5",X"34",X"65",X"39",X"85",X"07",X"A9",X"00",X"85",X"0A",X"A2",X"04",
		X"20",X"A9",X"E4",X"A6",X"CF",X"B5",X"4D",X"C9",X"03",X"D0",X"0D",X"A5",X"07",X"10",X"09",X"AD",
		X"AD",X"3A",X"AE",X"AC",X"3A",X"4C",X"1E",X"D7",X"AE",X"AA",X"3A",X"AD",X"AB",X"3A",X"20",X"53",
		X"E4",X"60",X"20",X"80",X"80",X"A0",X"20",X"60",X"00",X"00",X"60",X"00",X"00",X"00",X"60",X"60",
		X"00",X"C0",X"00",X"00",X"24",X"EC",X"1A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"24",
		X"00",X"F0",X"00",X"00",X"00",X"00",X"0A",X"EE",X"04",X"00",X"00",X"00",X"F8",X"08",X"08",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"40",X"60",X"C0",X"80",X"00",X"00",X"00",X"C0",X"A0",X"80",X"00",
		X"40",X"40",X"00",X"00",X"02",X"00",X"00",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"04",
		X"04",X"00",X"00",X"20",X"60",X"00",X"00",X"20",X"40",X"00",X"20",X"A0",X"20",X"00",X"00",X"40",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"F0",X"00",X"30",X"30",X"04",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"C0",X"40",X"60",X"20",X"C0",X"60",X"40",X"00",X"00",
		X"00",X"00",X"A0",X"00",X"80",X"00",X"80",X"60",X"00",X"00",X"80",X"00",X"80",X"00",X"00",X"80",
		X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"A0",X"60",X"60",X"80",X"40",X"00",X"80",X"60",X"00",X"60",X"00",X"60",X"00",
		X"60",X"00",X"60",X"00",X"20",X"00",X"00",X"60",X"00",X"60",X"40",X"40",X"40",X"60",X"60",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2C",X"2C",X"12",X"12",X"24",X"00",
		X"00",X"00",X"00",X"00",X"00",X"A0",X"A0",X"60",X"60",X"00",X"00",X"60",X"40",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"40",X"00",X"20",X"00",X"00",X"00",X"00",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"40",X"00",X"00",X"A0",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"80",X"00",X"60",X"60",X"00",
		X"00",X"00",X"C0",X"00",X"00",X"00",X"A0",X"00",X"00",X"80",X"00",X"00",X"00",X"60",X"00",X"A0",
		X"00",X"00",X"16",X"00",X"00",X"00",X"16",X"00",X"00",X"0A",X"00",X"00",X"00",X"0A",X"00",X"26",
		X"00",X"00",X"A6",X"CF",X"B5",X"4D",X"AA",X"BD",X"31",X"C1",X"29",X"20",X"F0",X"15",X"AD",X"43",
		X"01",X"30",X"06",X"20",X"8D",X"D9",X"4C",X"7C",X"D8",X"20",X"7E",X"D9",X"A2",X"EC",X"A9",X"3C",
		X"20",X"53",X"E4",X"60",X"A6",X"CF",X"B5",X"00",X"C9",X"22",X"F0",X"0B",X"C9",X"24",X"F0",X"04",
		X"C9",X"08",X"D0",X"03",X"4C",X"B1",X"D8",X"BC",X"3C",X"01",X"D0",X"14",X"C9",X"1C",X"D0",X"07",
		X"A6",X"86",X"86",X"21",X"4C",X"CB",X"D8",X"A2",X"01",X"86",X"21",X"20",X"CB",X"D8",X"10",X"FB",
		X"60",X"A6",X"CF",X"B5",X"4D",X"AA",X"BD",X"31",X"C1",X"30",X"0F",X"A2",X"01",X"86",X"22",X"A2",
		X"03",X"86",X"21",X"20",X"CB",X"D8",X"C6",X"22",X"10",X"F9",X"60",X"20",X"66",X"E4",X"A6",X"21",
		X"BD",X"34",X"01",X"D0",X"2A",X"BD",X"0C",X"01",X"85",X"07",X"BD",X"08",X"01",X"85",X"06",X"BD",
		X"18",X"01",X"85",X"05",X"BD",X"14",X"01",X"85",X"04",X"A2",X"04",X"A9",X"00",X"85",X"0A",X"20",
		X"A9",X"E4",X"A5",X"21",X"0A",X"A8",X"B9",X"7B",X"4A",X"BE",X"7A",X"4A",X"20",X"53",X"E4",X"C6",
		X"21",X"A6",X"21",X"60",X"A2",X"01",X"86",X"24",X"20",X"99",X"D9",X"20",X"66",X"E4",X"A9",X"A0",
		X"85",X"04",X"A9",X"D0",X"85",X"06",X"A9",X"01",X"85",X"07",X"A6",X"24",X"BD",X"54",X"D9",X"85",
		X"05",X"A9",X"00",X"85",X"0A",X"A2",X"04",X"20",X"A9",X"E4",X"A9",X"04",X"18",X"65",X"24",X"85",
		X"21",X"A5",X"D0",X"F0",X"09",X"A5",X"24",X"C5",X"CF",X"F0",X"03",X"20",X"A0",X"D9",X"38",X"A6",
		X"21",X"BD",X"62",X"01",X"20",X"47",X"DE",X"C6",X"21",X"C6",X"21",X"10",X"F2",X"C6",X"24",X"10",
		X"B7",X"4C",X"99",X"D9",X"FE",X"00",X"A0",X"01",X"91",X"08",X"88",X"8A",X"91",X"08",X"A5",X"08",
		X"18",X"69",X"02",X"85",X"08",X"90",X"02",X"E6",X"09",X"60",X"A0",X"00",X"F0",X"1A",X"A0",X"01",
		X"D0",X"16",X"A0",X"02",X"D0",X"12",X"A0",X"04",X"D0",X"0E",X"A0",X"03",X"D0",X"0A",X"A0",X"05",
		X"D0",X"06",X"A0",X"06",X"D0",X"02",X"A0",X"07",X"A9",X"00",X"4C",X"5F",X"E4",X"AD",X"0A",X"60",
		X"29",X"0C",X"D0",X"02",X"09",X"01",X"A8",X"D0",X"EF",X"A9",X"01",X"A0",X"40",X"4C",X"7F",X"E4",
		X"A0",X"68",X"A9",X"01",X"4C",X"7F",X"E4",X"A9",X"01",X"85",X"24",X"20",X"99",X"D9",X"20",X"66",
		X"E4",X"20",X"72",X"D9",X"A9",X"A0",X"85",X"04",X"85",X"06",X"A9",X"01",X"85",X"07",X"A6",X"24",
		X"BD",X"F6",X"D9",X"85",X"05",X"A9",X"00",X"85",X"0A",X"A2",X"04",X"20",X"A9",X"E4",X"A9",X"04",
		X"18",X"65",X"24",X"85",X"21",X"A5",X"D0",X"F0",X"09",X"A5",X"24",X"C5",X"CF",X"F0",X"03",X"20",
		X"A0",X"D9",X"38",X"A6",X"21",X"BD",X"68",X"01",X"20",X"47",X"DE",X"C6",X"21",X"C6",X"21",X"10",
		X"F2",X"C6",X"24",X"10",X"B6",X"60",X"FE",X"00",X"A8",X"BE",X"4A",X"4D",X"B9",X"4B",X"4D",X"20",
		X"56",X"D9",X"60",X"20",X"6E",X"D9",X"A2",X"01",X"86",X"21",X"B5",X"42",X"F0",X"30",X"30",X"2E",
		X"C9",X"05",X"90",X"02",X"A9",X"05",X"85",X"22",X"BD",X"47",X"DA",X"48",X"BD",X"45",X"DA",X"AA",
		X"68",X"20",X"EE",X"E1",X"AD",X"C7",X"45",X"AE",X"C6",X"45",X"20",X"56",X"D9",X"A4",X"21",X"B9",
		X"49",X"DA",X"BE",X"4B",X"DA",X"A0",X"00",X"20",X"8A",X"E4",X"C6",X"22",X"D0",X"E6",X"C6",X"21",
		X"A6",X"21",X"10",X"C6",X"60",X"74",X"74",X"A0",X"58",X"F8",X"08",X"FB",X"FB",X"A6",X"CF",X"B5",
		X"00",X"C9",X"08",X"D0",X"33",X"B5",X"4D",X"AA",X"BD",X"31",X"C1",X"29",X"A8",X"F0",X"29",X"AD",
		X"3E",X"01",X"30",X"24",X"20",X"86",X"D9",X"20",X"66",X"E4",X"A9",X"E0",X"AA",X"A0",X"00",X"20",
		X"8A",X"E4",X"AD",X"3E",X"01",X"D0",X"0D",X"38",X"20",X"54",X"DE",X"18",X"A9",X"00",X"20",X"54",
		X"DE",X"4C",X"88",X"DA",X"38",X"20",X"47",X"DE",X"60",X"A6",X"CF",X"B5",X"00",X"C9",X"1A",X"D0",
		X"42",X"BD",X"7A",X"01",X"C9",X"01",X"D0",X"3B",X"4A",X"85",X"39",X"B4",X"4D",X"B9",X"D4",X"DA",
		X"85",X"38",X"A0",X"03",X"06",X"38",X"26",X"39",X"88",X"10",X"F9",X"B5",X"E9",X"18",X"65",X"38",
		X"85",X"38",X"90",X"02",X"E6",X"39",X"20",X"66",X"E4",X"A9",X"F8",X"A2",X"04",X"A0",X"00",X"20",
		X"8A",X"E4",X"A5",X"39",X"38",X"20",X"47",X"DE",X"A5",X"38",X"20",X"47",X"DE",X"A9",X"00",X"18",
		X"20",X"47",X"DE",X"60",X"00",X"02",X"06",X"12",X"20",X"A6",X"CF",X"B5",X"00",X"C9",X"08",X"D0",
		X"22",X"20",X"66",X"E4",X"A9",X"6F",X"A2",X"68",X"A0",X"00",X"20",X"8A",X"E4",X"A6",X"CF",X"B5",
		X"E9",X"38",X"20",X"47",X"DE",X"A9",X"00",X"20",X"47",X"DE",X"A9",X"20",X"05",X"F2",X"85",X"F2",
		X"4C",X"09",X"DB",X"A9",X"DF",X"25",X"F2",X"85",X"F2",X"60",X"A5",X"F5",X"29",X"02",X"F0",X"22",
		X"20",X"66",X"E4",X"A0",X"00",X"A2",X"5C",X"A9",X"0C",X"20",X"8A",X"E4",X"A6",X"CF",X"BD",X"16",
		X"05",X"38",X"20",X"47",X"DE",X"A6",X"CF",X"BD",X"14",X"05",X"20",X"47",X"DE",X"A9",X"00",X"20",
		X"47",X"DE",X"60",X"20",X"7A",X"D9",X"A9",X"7F",X"25",X"F4",X"85",X"F4",X"A4",X"CF",X"B9",X"F6",
		X"00",X"48",X"29",X"03",X"AA",X"BD",X"F2",X"DB",X"18",X"65",X"CF",X"85",X"24",X"68",X"29",X"01",
		X"85",X"7B",X"AA",X"BD",X"F2",X"DB",X"85",X"7B",X"A9",X"04",X"85",X"23",X"20",X"66",X"E4",X"A6",
		X"24",X"BD",X"44",X"01",X"30",X"2F",X"A6",X"7B",X"BD",X"A2",X"DB",X"85",X"07",X"BD",X"B6",X"DB",
		X"85",X"06",X"BD",X"CA",X"DB",X"85",X"05",X"BD",X"DE",X"DB",X"85",X"04",X"86",X"22",X"A9",X"00",
		X"85",X"0A",X"A2",X"04",X"20",X"A9",X"E4",X"A6",X"24",X"BD",X"71",X"04",X"38",X"20",X"47",X"DE",
		X"A9",X"00",X"20",X"47",X"DE",X"C6",X"7B",X"C6",X"7B",X"C6",X"24",X"C6",X"24",X"C6",X"23",X"10",
		X"BB",X"60",X"02",X"02",X"FE",X"FE",X"FD",X"FD",X"02",X"02",X"00",X"00",X"02",X"02",X"FF",X"FF",
		X"FD",X"FD",X"FF",X"FF",X"02",X"02",X"20",X"20",X"00",X"00",X"60",X"60",X"00",X"00",X"00",X"00",
		X"00",X"00",X"90",X"90",X"80",X"80",X"30",X"30",X"10",X"10",X"02",X"02",X"02",X"02",X"FD",X"FD",
		X"FD",X"FD",X"FD",X"FD",X"FF",X"FF",X"02",X"02",X"FF",X"FF",X"FD",X"FD",X"02",X"02",X"60",X"60",
		X"80",X"80",X"60",X"60",X"E0",X"E0",X"00",X"00",X"A0",X"A0",X"E0",X"E0",X"FF",X"FF",X"10",X"10",
		X"E0",X"E0",X"08",X"12",X"1C",X"A0",X"1F",X"84",X"23",X"A5",X"F2",X"85",X"38",X"A5",X"F3",X"85",
		X"39",X"A5",X"F4",X"85",X"3A",X"A5",X"F5",X"85",X"3B",X"06",X"38",X"26",X"39",X"26",X"3A",X"26",
		X"3B",X"90",X"14",X"A4",X"23",X"B9",X"48",X"DC",X"BE",X"2C",X"DC",X"20",X"EE",X"E1",X"A4",X"23",
		X"B9",X"64",X"DC",X"A8",X"20",X"FC",X"E1",X"C6",X"23",X"10",X"DE",X"60",X"00",X"00",X"C0",X"C0",
		X"C0",X"60",X"5C",X"1C",X"50",X"44",X"38",X"2C",X"20",X"14",X"00",X"5C",X"34",X"28",X"C8",X"28",
		X"14",X"F0",X"F0",X"F0",X"10",X"5C",X"28",X"28",X"00",X"00",X"D0",X"D0",X"D0",X"6C",X"D0",X"91",
		X"D6",X"CA",X"C7",X"D0",X"D0",X"D9",X"18",X"EC",X"E0",X"DA",X"D0",X"E0",X"08",X"30",X"C0",X"B8",
		X"F0",X"D6",X"D8",X"D8",X"00",X"00",X"0B",X"09",X"09",X"0A",X"08",X"07",X"0C",X"0D",X"0E",X"0F",
		X"10",X"11",X"1A",X"1B",X"1C",X"1D",X"1E",X"1F",X"20",X"21",X"22",X"06",X"23",X"24",X"25",X"26",
		X"AD",X"35",X"04",X"A0",X"07",X"0A",X"B0",X"03",X"88",X"D0",X"FA",X"84",X"23",X"B9",X"A4",X"DC",
		X"A2",X"00",X"20",X"EE",X"E1",X"A4",X"23",X"B9",X"AC",X"DC",X"A8",X"20",X"FC",X"E1",X"A0",X"1A",
		X"20",X"FC",X"E1",X"60",X"E6",X"E6",X"E0",X"E8",X"DC",X"D4",X"CC",X"D0",X"12",X"13",X"14",X"15",
		X"16",X"17",X"18",X"19",X"A6",X"CF",X"B5",X"00",X"C9",X"12",X"F0",X"39",X"C9",X"24",X"F0",X"0E",
		X"C9",X"22",X"F0",X"0A",X"C9",X"16",X"D0",X"5B",X"A5",X"F4",X"29",X"9F",X"85",X"F4",X"A5",X"D6",
		X"F0",X"18",X"20",X"5A",X"DD",X"A9",X"E0",X"A2",X"34",X"20",X"EE",X"E1",X"A0",X"00",X"20",X"FC",
		X"E1",X"A5",X"F4",X"29",X"FE",X"09",X"08",X"4C",X"F3",X"DC",X"20",X"3C",X"DD",X"A9",X"01",X"05",
		X"F4",X"29",X"F7",X"85",X"F4",X"A9",X"E6",X"A2",X"40",X"20",X"EE",X"E1",X"A0",X"01",X"20",X"FC",
		X"E1",X"A6",X"CF",X"BD",X"68",X"01",X"1D",X"6A",X"01",X"1D",X"6C",X"01",X"D0",X"15",X"B5",X"00",
		X"C9",X"12",X"D0",X"0F",X"A9",X"E0",X"A2",X"38",X"20",X"EE",X"E1",X"A0",X"02",X"20",X"FC",X"E1",
		X"4C",X"23",X"DD",X"A2",X"74",X"A9",X"F4",X"20",X"EE",X"E1",X"A0",X"03",X"20",X"FC",X"E1",X"A2",
		X"68",X"A9",X"F8",X"20",X"EE",X"E1",X"A0",X"04",X"20",X"FC",X"E1",X"60",X"A5",X"F1",X"29",X"03",
		X"A8",X"C0",X"02",X"F0",X"0A",X"B9",X"56",X"DD",X"05",X"F5",X"85",X"F5",X"4C",X"55",X"DD",X"A5",
		X"F4",X"09",X"02",X"85",X"F4",X"60",X"00",X"04",X"00",X"08",X"A5",X"F5",X"29",X"F3",X"85",X"F5",
		X"A5",X"F4",X"29",X"FD",X"85",X"F4",X"60",X"A5",X"D0",X"D0",X"3B",X"A6",X"CF",X"B5",X"00",X"C9",
		X"1E",X"F0",X"33",X"A5",X"D6",X"F0",X"19",X"A2",X"29",X"A9",X"08",X"A0",X"00",X"20",X"EE",X"E1",
		X"A5",X"D6",X"20",X"A7",X"DD",X"A5",X"22",X"38",X"20",X"47",X"DE",X"A5",X"23",X"20",X"47",X"DE",
		X"A6",X"CF",X"B5",X"00",X"C9",X"22",X"D0",X"0E",X"A9",X"C4",X"A2",X"C6",X"20",X"EE",X"E1",X"A2",
		X"2E",X"A9",X"56",X"20",X"53",X"E4",X"60",X"85",X"24",X"A0",X"07",X"A9",X"00",X"85",X"23",X"85",
		X"22",X"F8",X"06",X"24",X"A5",X"23",X"65",X"23",X"85",X"23",X"A5",X"22",X"65",X"22",X"85",X"22",
		X"88",X"10",X"EF",X"D8",X"60",X"A9",X"07",X"85",X"21",X"20",X"EB",X"DD",X"20",X"66",X"E4",X"A6",
		X"21",X"BC",X"AA",X"04",X"A9",X"02",X"20",X"7F",X"E4",X"A5",X"21",X"0A",X"A8",X"BE",X"6A",X"4A",
		X"B9",X"6B",X"4A",X"20",X"53",X"E4",X"C6",X"21",X"10",X"E2",X"60",X"AD",X"AA",X"04",X"10",X"0D",
		X"AD",X"7F",X"01",X"30",X"08",X"CE",X"7F",X"01",X"10",X"03",X"20",X"2D",X"DE",X"A2",X"07",X"BD",
		X"AA",X"04",X"18",X"7D",X"B2",X"04",X"9D",X"AA",X"04",X"10",X"0E",X"A9",X"00",X"38",X"FD",X"B2",
		X"04",X"9D",X"B2",X"04",X"30",X"03",X"9D",X"AA",X"04",X"CA",X"10",X"E3",X"60",X"A2",X"07",X"A9",
		X"7F",X"9D",X"AA",X"04",X"A9",X"03",X"9D",X"B2",X"04",X"CA",X"10",X"F3",X"60",X"A2",X"07",X"A9",
		X"7F",X"9D",X"AA",X"04",X"CA",X"10",X"F8",X"A2",X"07",X"AD",X"0A",X"60",X"29",X"07",X"09",X"01",
		X"9D",X"B2",X"04",X"CA",X"10",X"F3",X"60",X"48",X"08",X"4A",X"4A",X"4A",X"4A",X"28",X"20",X"54",
		X"DE",X"68",X"29",X"0F",X"90",X"05",X"29",X"0F",X"F0",X"08",X"18",X"0A",X"08",X"20",X"F8",X"D9",
		X"28",X"60",X"AE",X"48",X"4D",X"AD",X"49",X"4D",X"08",X"20",X"56",X"D9",X"28",X"60",X"A9",X"00",
		X"85",X"1B",X"85",X"1C",X"A0",X"07",X"06",X"1B",X"26",X"1C",X"06",X"19",X"90",X"0B",X"A5",X"1A",
		X"18",X"65",X"1B",X"85",X"1B",X"90",X"02",X"E6",X"1C",X"88",X"10",X"EA",X"60",X"00",X"00",X"01",
		X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"0A",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"15",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"6B",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"73",X"6E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"21",X"26",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"4B",X"5A",X"5D",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"60",X"63",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"3E",X"41",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"79",X"76",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"81",X"7E",X"87",X"84",X"1B",X"1E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"8D",X"8A",X"93",X"90",X"00",X"00",X"00",
		X"00",X"00",X"00",X"9E",X"A9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"96",X"9B",X"00",X"00",X"00",X"00",X"10",X"08",X"BF",
		X"20",X"00",X"00",X"A7",X"20",X"FF",X"08",X"00",X"00",X"10",X"01",X"01",X"60",X"00",X"00",X"A4",
		X"10",X"FF",X"04",X"00",X"00",X"0A",X"FF",X"00",X"10",X"00",X"00",X"4F",X"30",X"FF",X"0A",X"46",
		X"20",X"FF",X"06",X"00",X"00",X"24",X"01",X"03",X"40",X"00",X"00",X"09",X"FF",X"00",X"10",X"00",
		X"00",X"30",X"02",X"00",X"0F",X"00",X"00",X"C0",X"01",X"02",X"0F",X"00",X"00",X"06",X"E0",X"00",
		X"01",X"05",X"E0",X"00",X"01",X"00",X"00",X"AF",X"10",X"00",X"01",X"A0",X"10",X"00",X"01",X"AF",
		X"10",X"00",X"01",X"A0",X"10",X"00",X"01",X"AF",X"10",X"00",X"01",X"A0",X"10",X"00",X"01",X"AF",
		X"10",X"00",X"01",X"A0",X"10",X"00",X"01",X"AF",X"10",X"00",X"01",X"A0",X"10",X"00",X"01",X"AF",
		X"10",X"00",X"01",X"A0",X"10",X"00",X"01",X"10",X"02",X"00",X"0F",X"00",X"00",X"A7",X"10",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
