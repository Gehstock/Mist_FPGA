library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity sol_sp_bits is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of sol_sp_bits is
	type rom is array(0 to  32767) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"6F",X"66",X"00",X"00",X"6F",X"66",X"00",X"00",X"6B",X"66",
		X"00",X"00",X"FF",X"A6",X"00",X"09",X"FF",X"A6",X"00",X"00",X"00",X"A6",X"00",X"00",X"B0",X"A6",
		X"00",X"0F",X"B0",X"66",X"00",X"0F",X"BB",X"66",X"00",X"60",X"FF",X"06",X"00",X"6A",X"6F",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"FF",X"90",X"00",X"00",X"00",X"B9",X"66",X"00",X"06",X"B9",X"66",
		X"00",X"66",X"B0",X"66",X"00",X"6F",X"90",X"66",X"00",X"99",X"9B",X"66",X"00",X"99",X"9B",X"66",
		X"00",X"00",X"BB",X"66",X"00",X"00",X"0F",X"66",X"00",X"00",X"60",X"00",X"00",X"00",X"60",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"B9",
		X"00",X"00",X"99",X"B0",X"00",X"00",X"9B",X"00",X"00",X"0B",X"9B",X"BB",X"00",X"0B",X"90",X"BB",
		X"00",X"0B",X"00",X"BB",X"00",X"0F",X"00",X"BB",X"00",X"B0",X"FF",X"B0",X"00",X"BF",X"FF",X"00",
		X"00",X"BF",X"FF",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"0B",X"00",X"00",X"00",X"B9",X"99",
		X"00",X"00",X"BB",X"B9",X"00",X"00",X"9F",X"B0",X"00",X"FF",X"FF",X"F0",X"00",X"BB",X"F9",X"F0",
		X"00",X"B9",X"F0",X"BB",X"00",X"B5",X"00",X"BB",X"00",X"50",X"99",X"BB",X"00",X"0F",X"90",X"BB",
		X"00",X"0F",X"90",X"BB",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"99",X"00",X"99",X"00",X"A9",
		X"00",X"99",X"99",X"A0",X"00",X"99",X"9B",X"60",X"00",X"9A",X"9B",X"BB",X"00",X"9A",X"90",X"BB",
		X"00",X"AA",X"AA",X"BB",X"00",X"AA",X"AA",X"BB",X"00",X"A0",X"AA",X"B0",X"00",X"AF",X"5A",X"00",
		X"00",X"BA",X"5A",X"00",X"00",X"BA",X"55",X"90",X"00",X"BB",X"55",X"00",X"00",X"9A",X"55",X"99",
		X"00",X"AA",X"AA",X"B9",X"00",X"AA",X"AA",X"B0",X"00",X"AA",X"AA",X"F0",X"00",X"AA",X"AA",X"F0",
		X"00",X"B9",X"F0",X"BB",X"00",X"99",X"00",X"6B",X"00",X"AA",X"99",X"AA",X"00",X"AA",X"90",X"BB",
		X"00",X"0A",X"99",X"BB",X"00",X"AA",X"99",X"00",X"00",X"AA",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"44",X"99",X"94",X"00",X"44",X"11",X"44",X"00",X"00",X"11",X"49",X"00",X"09",X"1F",X"49",
		X"00",X"99",X"BB",X"99",X"00",X"99",X"BB",X"09",X"00",X"99",X"BB",X"00",X"00",X"90",X"BB",X"B0",
		X"00",X"00",X"B0",X"BB",X"00",X"00",X"BB",X"B0",X"04",X"50",X"FF",X"B1",X"09",X"50",X"F0",X"BB",
		X"99",X"55",X"00",X"BB",X"99",X"00",X"00",X"BB",X"99",X"09",X"44",X"BB",X"99",X"00",X"04",X"9B",
		X"99",X"BB",X"04",X"9B",X"99",X"BB",X"04",X"BB",X"99",X"BB",X"BF",X"BB",X"99",X"BB",X"B0",X"BB",
		X"09",X"BB",X"BB",X"BB",X"00",X"1B",X"B0",X"B0",X"04",X"11",X"00",X"B9",X"04",X"91",X"00",X"B9",
		X"00",X"91",X"90",X"11",X"00",X"90",X"00",X"19",X"00",X"91",X"99",X"19",X"00",X"99",X"99",X"99",
		X"00",X"99",X"09",X"99",X"00",X"44",X"99",X"94",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"06",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FB",X"00",
		X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",
		X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",
		X"00",X"00",X"0B",X"00",X"00",X"0B",X"0B",X"00",X"00",X"BB",X"FB",X"00",X"00",X"0B",X"9F",X"00",
		X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",
		X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",
		X"00",X"00",X"0B",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9B",X"00",X"00",X"00",X"9B",X"00",
		X"00",X"00",X"9B",X"00",X"00",X"00",X"9B",X"00",X"00",X"00",X"9B",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",
		X"00",X"00",X"00",X"9F",X"00",X"00",X"00",X"9F",X"00",X"00",X"00",X"9F",X"00",X"00",X"00",X"99",
		X"00",X"FF",X"FF",X"99",X"00",X"99",X"99",X"99",X"0F",X"99",X"99",X"99",X"0F",X"99",X"F9",X"99",
		X"0F",X"9F",X"99",X"99",X"F9",X"99",X"99",X"99",X"F9",X"99",X"99",X"99",X"F9",X"99",X"99",X"99",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"0F",X"9F",X"00",X"00",X"F9",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"CC",X"BC",X"00",X"00",X"CC",X"0C",X"00",X"FF",X"C0",X"00",X"FF",
		X"F9",X"00",X"90",X"99",X"F9",X"00",X"90",X"99",X"F9",X"99",X"99",X"99",X"F9",X"99",X"99",X"99",
		X"F9",X"99",X"B9",X"99",X"F9",X"9B",X"0B",X"99",X"F9",X"B0",X"00",X"99",X"BB",X"00",X"00",X"BB",
		X"BB",X"00",X"00",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"9F",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"FF",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",
		X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",X"F9",X"00",
		X"00",X"00",X"F9",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"F9",X"00",
		X"00",X"00",X"F9",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",
		X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"9F",X"00",X"00",X"99",X"FF",
		X"00",X"00",X"99",X"00",X"00",X"00",X"9F",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"59",X"00",
		X"00",X"00",X"59",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"69",X"00",X"00",X"99",X"99",X"00",
		X"00",X"56",X"59",X"60",X"00",X"56",X"56",X"68",X"00",X"59",X"59",X"68",X"F9",X"99",X"69",X"68",
		X"09",X"99",X"69",X"99",X"00",X"56",X"59",X"99",X"00",X"56",X"59",X"99",X"00",X"59",X"59",X"99",
		X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"F9",X"00",
		X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"0B",X"BB",X"00",X"00",X"00",X"99",X"00",X"00",X"B0",X"BB",X"09",X"00",X"B0",X"CB",X"00",
		X"00",X"F0",X"FC",X"99",X"00",X"F0",X"CB",X"99",X"00",X"99",X"CB",X"00",X"00",X"00",X"0B",X"90",
		X"00",X"00",X"99",X"00",X"00",X"00",X"9F",X"90",X"00",X"00",X"9F",X"00",X"00",X"00",X"0B",X"00",
		X"00",X"00",X"B0",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"F0",X"00",X"00",X"99",X"9F",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",
		X"00",X"00",X"B9",X"99",X"00",X"00",X"0B",X"99",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"F0",X"00",X"00",X"BB",X"BF",
		X"00",X"00",X"BB",X"BF",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"0B",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"FB",X"00",X"00",X"00",X"FB",X"00",
		X"00",X"00",X"FB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"44",X"00",X"04",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"04",X"00",X"44",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"04",X"00",X"44",X"00",X"04",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"44",
		X"00",X"04",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",
		X"00",X"00",X"00",X"44",X"00",X"04",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",
		X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"90",X"90",
		X"00",X"00",X"96",X"9F",X"00",X"00",X"90",X"90",X"00",X"00",X"90",X"90",X"00",X"00",X"90",X"90",
		X"00",X"00",X"96",X"99",X"00",X"00",X"90",X"96",X"00",X"00",X"90",X"66",X"00",X"00",X"96",X"69",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"0F",X"00",X"00",X"BB",X"9F",
		X"00",X"00",X"BB",X"0F",X"00",X"00",X"BB",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FB",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"FB",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",
		X"00",X"00",X"0B",X"00",X"00",X"00",X"FB",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0B",X"00",
		X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",
		X"00",X"0B",X"0B",X"00",X"00",X"BB",X"0B",X"00",X"00",X"BB",X"0B",X"00",X"00",X"0B",X"0B",X"00",
		X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",
		X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",
		X"00",X"00",X"0B",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"FB",X"00",X"00",X"00",X"FB",X"00",X"00",X"00",X"FB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BB",X"0B",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BF",
		X"00",X"00",X"BB",X"BF",X"00",X"00",X"BB",X"F0",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"66",X"00",X"00",X"90",X"66",X"00",X"00",X"90",X"99",X"00",X"00",X"90",X"99",
		X"00",X"00",X"96",X"09",X"00",X"00",X"96",X"09",X"00",X"00",X"90",X"69",X"00",X"00",X"90",X"6F",
		X"00",X"00",X"90",X"00",X"00",X"00",X"96",X"00",X"00",X"00",X"96",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9F",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0B",X"00",
		X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0B",X"00",
		X"00",X"00",X"0B",X"00",X"00",X"00",X"FB",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0B",X"00",
		X"00",X"00",X"0B",X"00",X"00",X"0B",X"0B",X"00",X"00",X"BB",X"0B",X"00",X"00",X"0B",X"0B",X"00",
		X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"FB",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",
		X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"00",X"0B",X"99",X"00",X"00",X"B9",X"99",
		X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"9F",X"00",X"00",X"99",X"F0",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"F0",X"00",X"00",X"BB",X"BF",
		X"00",X"00",X"BB",X"BF",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"0B",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"FB",X"00",X"00",X"00",X"FB",X"00",
		X"00",X"00",X"FB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"FB",X"00",X"00",X"00",X"FB",X"00",X"00",X"00",X"FB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BB",X"0B",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BF",
		X"00",X"00",X"BB",X"BF",X"00",X"00",X"BB",X"F0",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"04",X"00",X"00",
		X"00",X"04",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"44",X"44",X"44",X"00",X"44",X"40",X"44",X"00",X"00",
		X"44",X"40",X"00",X"00",X"04",X"00",X"00",X"44",X"04",X"00",X"00",X"44",X"04",X"00",X"00",X"04",
		X"04",X"44",X"00",X"04",X"00",X"44",X"00",X"04",X"00",X"00",X"00",X"04",X"00",X"40",X"00",X"04",
		X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"04",X"00",X"00",
		X"00",X"04",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",
		X"00",X"00",X"00",X"BF",X"00",X"00",X"00",X"BF",X"00",X"00",X"00",X"BF",X"00",X"00",X"00",X"BB",
		X"00",X"FF",X"FF",X"BB",X"00",X"BB",X"BB",X"BB",X"0F",X"BB",X"BB",X"BB",X"0F",X"BB",X"FB",X"BB",
		X"0F",X"BF",X"BB",X"BB",X"FB",X"BF",X"BB",X"BB",X"FB",X"BB",X"BB",X"BB",X"FB",X"BB",X"BB",X"BB",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"0F",X"BF",X"00",X"00",X"FB",X"BB",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",
		X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"FF",X"BB",X"BB",X"FF",
		X"FB",X"BB",X"BB",X"BB",X"FB",X"BB",X"BB",X"BB",X"FB",X"BB",X"BB",X"BB",X"FB",X"BB",X"BB",X"BB",
		X"FB",X"BB",X"FB",X"BB",X"0F",X"BF",X"0F",X"BF",X"00",X"F0",X"00",X"F0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",
		X"00",X"00",X"00",X"BF",X"00",X"00",X"00",X"BF",X"00",X"00",X"00",X"BF",X"00",X"00",X"00",X"BB",
		X"00",X"FF",X"FF",X"BB",X"00",X"BB",X"BB",X"BB",X"0F",X"BB",X"BB",X"BB",X"0F",X"BB",X"FB",X"BB",
		X"0F",X"BF",X"BB",X"BB",X"FB",X"BF",X"BB",X"BB",X"FB",X"BB",X"BB",X"BB",X"FB",X"BB",X"BB",X"BB",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"11",X"00",X"00",X"16",X"66",X"00",X"00",X"10",X"06",X"00",X"00",X"10",X"06",X"00",
		X"00",X"10",X"06",X"00",X"00",X"10",X"06",X"00",X"00",X"16",X"66",X"00",X"00",X"01",X"11",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"11",X"00",X"00",X"16",X"66",X"00",
		X"00",X"10",X"06",X"00",X"00",X"10",X"06",X"00",X"00",X"10",X"06",X"00",X"00",X"10",X"06",X"00",
		X"00",X"16",X"66",X"00",X"00",X"01",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"11",X"00",X"00",X"16",X"66",X"00",
		X"00",X"10",X"06",X"00",X"00",X"10",X"06",X"00",X"00",X"10",X"06",X"00",X"00",X"10",X"06",X"00",
		X"00",X"16",X"06",X"00",X"00",X"01",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"11",X"00",X"00",X"16",X"66",X"00",X"00",X"10",X"06",X"00",X"00",X"10",X"06",X"00",
		X"00",X"10",X"06",X"00",X"00",X"10",X"06",X"00",X"00",X"16",X"66",X"00",X"00",X"01",X"11",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"11",X"00",X"00",X"16",X"66",X"00",
		X"00",X"10",X"06",X"00",X"00",X"10",X"06",X"00",X"00",X"10",X"06",X"00",X"00",X"10",X"06",X"00",
		X"00",X"16",X"66",X"00",X"00",X"01",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"11",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"66",X"00",
		X"00",X"01",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"11",X"00",X"00",X"16",X"66",X"00",X"00",X"10",X"06",X"00",X"00",X"10",X"06",X"00",
		X"00",X"10",X"06",X"00",X"00",X"10",X"06",X"00",X"00",X"16",X"66",X"00",X"00",X"01",X"11",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"11",X"00",X"00",X"16",X"66",X"00",
		X"00",X"10",X"06",X"00",X"00",X"10",X"06",X"00",X"00",X"10",X"06",X"00",X"00",X"10",X"06",X"00",
		X"00",X"16",X"66",X"00",X"00",X"01",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"1B",X"00",X"00",X"0F",X"1B",X"00",X"00",X"00",X"1B",X"00",X"00",X"00",X"11",X"00",X"00",
		X"00",X"11",X"F0",X"00",X"00",X"11",X"BF",X"00",X"00",X"11",X"BB",X"00",X"00",X"11",X"BB",X"00",
		X"00",X"F1",X"BB",X"00",X"00",X"0F",X"BB",X"00",X"00",X"0F",X"BF",X"00",X"00",X"0F",X"BF",X"00",
		X"00",X"0F",X"F0",X"00",X"00",X"0F",X"F0",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"F0",X"00",X"00",X"0F",X"F0",X"00",
		X"00",X"0F",X"BF",X"00",X"00",X"0F",X"BF",X"00",X"00",X"0F",X"BB",X"00",X"00",X"F1",X"BB",X"00",
		X"00",X"11",X"BB",X"00",X"00",X"11",X"BB",X"00",X"00",X"11",X"BF",X"00",X"00",X"11",X"F0",X"00",
		X"00",X"11",X"00",X"00",X"00",X"1B",X"00",X"00",X"0F",X"1B",X"00",X"00",X"0F",X"1B",X"00",X"00",
		X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"0F",X"11",X"00",X"00",X"FB",X"11",
		X"00",X"00",X"BB",X"1B",X"00",X"00",X"BB",X"1B",X"00",X"00",X"BB",X"1F",X"00",X"00",X"BB",X"F0",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"FB",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"FB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BB",X"F0",X"00",X"00",X"BB",X"1F",X"00",X"00",X"BB",X"1B",X"00",X"00",X"BB",X"1B",
		X"00",X"00",X"FB",X"11",X"00",X"00",X"0F",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"0F",X"BB",X"00",X"00",X"FF",X"BB",X"00",X"00",X"BB",X"BB",X"00",
		X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"0F",X"BB",X"BB",X"00",X"0F",X"00",X"BB",X"00",
		X"0F",X"00",X"BB",X"00",X"0F",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"0F",X"00",X"BB",X"00",X"0F",X"00",X"BB",X"00",
		X"0F",X"00",X"BB",X"00",X"0F",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",
		X"00",X"BB",X"BB",X"00",X"00",X"FF",X"BB",X"00",X"00",X"0F",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",
		X"00",X"00",X"60",X"66",X"00",X"00",X"66",X"66",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",
		X"00",X"60",X"06",X"00",X"00",X"60",X"0F",X"B0",X"00",X"66",X"60",X"00",X"00",X"6F",X"66",X"60",
		X"00",X"66",X"60",X"00",X"00",X"60",X"0F",X"B0",X"00",X"60",X"06",X"00",X"00",X"00",X"66",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"66",X"00",X"00",X"60",X"66",X"00",X"00",X"00",X"66",
		X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"0F",X"BB",X"00",X"00",X"FF",X"BB",X"00",X"00",X"BB",X"BB",X"00",
		X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"0F",X"BB",X"BB",X"00",X"0F",X"00",X"BB",X"00",
		X"0F",X"00",X"BB",X"00",X"0F",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"0F",X"00",X"BB",X"00",X"0F",X"00",X"BB",X"00",
		X"0F",X"00",X"BB",X"00",X"0F",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",
		X"00",X"BB",X"BB",X"00",X"00",X"FF",X"BB",X"00",X"00",X"0F",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",
		X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"40",X"00",X"44",X"00",X"40",X"00",X"44",X"00",X"00",
		X"00",X"00",X"00",X"44",X"00",X"40",X"00",X"44",X"00",X"44",X"00",X"00",X"00",X"04",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"04",X"00",X"04",X"00",X"04",
		X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"04",X"04",X"00",X"00",
		X"00",X"44",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"04",X"00",X"44",X"00",X"00",X"00",X"04",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",
		X"00",X"04",X"00",X"44",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"44",X"00",X"00",X"00",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"44",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"44",
		X"00",X"04",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"BB",X"00",X"00",X"BB",X"BB",X"00",
		X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BF",X"B0",X"00",X"0F",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"F0",X"00",X"00",X"BB",X"BF",X"B0",X"00",X"BB",X"BB",X"00",
		X"00",X"BB",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"50",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"50",X"00",X"00",X"00",X"00",X"00",
		X"00",X"50",X"11",X"0B",X"00",X"00",X"11",X"BB",X"00",X"50",X"11",X"BF",X"00",X"00",X"11",X"F0",
		X"00",X"00",X"1C",X"55",X"00",X"00",X"10",X"00",X"00",X"00",X"1C",X"5C",X"00",X"00",X"11",X"10",
		X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"BF",X"00",X"05",X"50",X"BB",X"00",X"00",X"00",X"0B",
		X"00",X"05",X"00",X"50",X"00",X"00",X"00",X"0B",X"00",X"05",X"05",X"0B",X"00",X"00",X"00",X"00",
		X"00",X"05",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"44",X"00",X"44",
		X"00",X"40",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"44",X"00",X"40",X"00",X"00",X"00",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"04",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"04",X"00",X"44",
		X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"00",X"00",X"00",X"44",X"00",X"04",X"00",X"44",X"00",X"04",X"00",X"04",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",
		X"00",X"BB",X"FB",X"B0",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"BB",X"FB",X"B0",X"00",X"BB",X"BB",X"00",
		X"00",X"BB",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9B",X"00",X"00",X"00",X"9B",X"00",
		X"00",X"00",X"9B",X"00",X"00",X"00",X"9B",X"00",X"00",X"00",X"9B",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",
		X"00",X"00",X"66",X"00",X"00",X"66",X"66",X"60",X"00",X"66",X"6F",X"60",X"00",X"66",X"6F",X"60",
		X"00",X"66",X"6F",X"66",X"00",X"66",X"60",X"66",X"00",X"66",X"66",X"66",X"00",X"06",X"6B",X"00",
		X"00",X"66",X"60",X"66",X"00",X"66",X"60",X"66",X"00",X"66",X"60",X"66",X"00",X"66",X"60",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"66",X"00",
		X"00",X"00",X"06",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"06",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"70",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"CC",X"0C",X"00",X"00",X"CC",X"0C",
		X"00",X"00",X"CC",X"0C",X"00",X"00",X"55",X"0C",X"00",X"CC",X"55",X"07",X"00",X"CC",X"55",X"C7",
		X"00",X"CC",X"55",X"C7",X"00",X"C0",X"55",X"CC",X"00",X"05",X"B5",X"CC",X"00",X"55",X"5B",X"5C",
		X"00",X"55",X"BB",X"50",X"00",X"55",X"5B",X"50",X"00",X"C5",X"B5",X"0C",X"00",X"CC",X"55",X"CC",
		X"00",X"CC",X"55",X"CC",X"00",X"CC",X"55",X"C7",X"00",X"00",X"55",X"C7",X"00",X"00",X"55",X"07",
		X"00",X"00",X"CC",X"0C",X"00",X"00",X"CC",X"0C",X"00",X"00",X"CC",X"0C",X"00",X"00",X"70",X"00",
		X"00",X"00",X"70",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"C0",X"00",X"00",X"00",X"0F",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"F0",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"0C",
		X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"DF",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"22",X"55",X"20",X"00",X"22",X"55",X"22",
		X"00",X"22",X"00",X"22",X"00",X"CC",X"55",X"C2",X"00",X"22",X"55",X"20",X"00",X"22",X"55",X"20",
		X"00",X"22",X"55",X"20",X"00",X"25",X"55",X"20",X"00",X"55",X"55",X"55",X"00",X"55",X"AF",X"55",
		X"00",X"55",X"AA",X"55",X"02",X"55",X"AF",X"52",X"02",X"55",X"5F",X"52",X"02",X"55",X"5A",X"52",
		X"02",X"05",X"55",X"02",X"02",X"55",X"5A",X"02",X"02",X"55",X"5F",X"02",X"02",X"55",X"AF",X"02",
		X"00",X"55",X"AA",X"05",X"00",X"55",X"AF",X"05",X"00",X"55",X"55",X"55",X"00",X"20",X"55",X"20",
		X"00",X"22",X"55",X"20",X"00",X"22",X"00",X"20",X"00",X"22",X"55",X"20",X"00",X"CC",X"55",X"C2",
		X"00",X"22",X"55",X"22",X"00",X"22",X"55",X"22",X"00",X"22",X"55",X"20",X"00",X"02",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"11",X"00",X"00",X"16",X"60",X"00",
		X"00",X"10",X"06",X"00",X"00",X"10",X"06",X"00",X"00",X"10",X"06",X"00",X"00",X"10",X"06",X"00",
		X"00",X"16",X"60",X"00",X"00",X"01",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"11",X"00",X"00",X"16",X"66",X"00",X"00",X"10",X"06",X"00",X"00",X"10",X"06",X"00",
		X"00",X"10",X"06",X"00",X"00",X"10",X"06",X"00",X"00",X"16",X"66",X"00",X"00",X"01",X"11",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"11",X"00",X"00",X"16",X"66",X"00",
		X"00",X"10",X"06",X"00",X"00",X"10",X"06",X"00",X"00",X"10",X"06",X"00",X"00",X"10",X"06",X"00",
		X"00",X"16",X"66",X"00",X"00",X"01",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"11",X"00",X"00",X"16",X"66",X"00",
		X"00",X"16",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"16",X"00",X"00",
		X"00",X"16",X"66",X"00",X"00",X"01",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"11",X"00",X"00",X"16",X"66",X"00",X"00",X"10",X"06",X"00",X"00",X"10",X"06",X"00",
		X"00",X"10",X"06",X"00",X"00",X"10",X"06",X"00",X"00",X"16",X"66",X"00",X"00",X"01",X"11",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"11",X"00",X"00",X"16",X"66",X"00",
		X"00",X"10",X"06",X"00",X"00",X"10",X"06",X"00",X"00",X"10",X"06",X"00",X"00",X"10",X"06",X"00",
		X"00",X"16",X"66",X"00",X"00",X"01",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"66",X"66",
		X"00",X"00",X"66",X"66",X"00",X"00",X"66",X"66",X"00",X"00",X"60",X"00",X"00",X"00",X"66",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"BB",X"00",X"00",X"60",X"00",X"00",X"00",X"66",X"66",
		X"00",X"00",X"60",X"00",X"00",X"00",X"0F",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",
		X"00",X"00",X"60",X"00",X"00",X"00",X"66",X"66",X"00",X"00",X"66",X"66",X"00",X"00",X"66",X"66",
		X"00",X"00",X"66",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"06",X"66",X"00",
		X"00",X"66",X"66",X"00",X"00",X"66",X"66",X"60",X"00",X"66",X"6F",X"60",X"00",X"66",X"6F",X"66",
		X"00",X"66",X"6F",X"66",X"00",X"66",X"60",X"66",X"00",X"66",X"66",X"66",X"00",X"06",X"6B",X"00",
		X"00",X"66",X"60",X"66",X"00",X"66",X"60",X"66",X"00",X"66",X"60",X"66",X"00",X"66",X"60",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"D4",X"00",X"00",X"00",X"FD",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0D",X"00",X"00",X"0F",X"F0",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CB",X"00",X"90",
		X"00",X"CC",X"00",X"99",X"00",X"0C",X"B0",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",
		X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"0C",X"B0",X"99",X"00",X"CC",X"00",X"99",
		X"00",X"CB",X"00",X"90",X"00",X"CB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"05",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"05",X"00",X"00",X"00",X"00",
		X"00",X"50",X"05",X"05",X"00",X"00",X"00",X"00",X"05",X"50",X"05",X"05",X"00",X"B0",X"00",X"00",
		X"55",X"5B",X"C0",X"05",X"00",X"01",X"00",X"00",X"05",X"11",X"CC",X"00",X"00",X"11",X"00",X"00",
		X"05",X"51",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"CC",X"00",X"00",X"10",X"00",X"00",
		X"50",X"15",X"00",X"00",X"00",X"10",X"00",X"00",X"50",X"11",X"00",X"00",X"00",X"01",X"00",X"00",
		X"00",X"B5",X"01",X"50",X"00",X"00",X"00",X"00",X"00",X"05",X"50",X"50",X"00",X"00",X"00",X"00",
		X"00",X"05",X"50",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"50",X"00",X"00",X"00",X"00",
		X"00",X"00",X"50",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"BF",X"00",
		X"00",X"00",X"B0",X"00",X"00",X"00",X"F0",X"00",X"00",X"90",X"00",X"00",X"00",X"FF",X"0B",X"00",
		X"00",X"FF",X"BB",X"00",X"00",X"FF",X"BB",X"00",X"00",X"00",X"9B",X"00",X"00",X"0B",X"B6",X"00",
		X"00",X"6B",X"00",X"00",X"00",X"FF",X"B0",X"00",X"00",X"9B",X"0B",X"00",X"00",X"99",X"00",X"00",
		X"00",X"FF",X"90",X"00",X"00",X"FF",X"90",X"00",X"00",X"FF",X"BB",X"00",X"00",X"99",X"F0",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"99",X"00",
		X"00",X"00",X"9B",X"00",X"99",X"0F",X"BB",X"00",X"BB",X"BB",X"BB",X"B0",X"B0",X"9B",X"BB",X"B9",
		X"B0",X"BB",X"0B",X"B0",X"B0",X"F9",X"00",X"00",X"00",X"F9",X"F9",X"00",X"00",X"FF",X"F9",X"00",
		X"00",X"FF",X"FF",X"00",X"00",X"0F",X"99",X"00",X"00",X"BB",X"9F",X"00",X"00",X"09",X"00",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"0B",X"BB",X"0B",X"00",X"F9",X"BB",X"0B",X"00",X"99",X"9F",X"BB",
		X"00",X"90",X"90",X"9B",X"00",X"99",X"99",X"90",X"B0",X"FF",X"B9",X"00",X"BB",X"FF",X"BB",X"00",
		X"9B",X"F9",X"BB",X"00",X"9B",X"09",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"90",X"00",X"99",X"96",X"00",
		X"00",X"99",X"9A",X"00",X"99",X"AA",X"BB",X"00",X"BB",X"AA",X"BB",X"B0",X"B0",X"AA",X"B9",X"B9",
		X"B0",X"AA",X"0B",X"B0",X"B0",X"A9",X"AA",X"00",X"00",X"F9",X"AA",X"00",X"00",X"FF",X"69",X"00",
		X"00",X"AA",X"6A",X"00",X"00",X"0F",X"5A",X"00",X"00",X"BB",X"5A",X"00",X"00",X"A9",X"59",X"00",
		X"00",X"AA",X"AA",X"00",X"00",X"AB",X"AA",X"0B",X"00",X"A9",X"99",X"0B",X"00",X"A9",X"99",X"BB",
		X"00",X"90",X"99",X"9B",X"00",X"99",X"9A",X"90",X"B0",X"9A",X"9A",X"00",X"BB",X"9A",X"BA",X"00",
		X"9B",X"F9",X"BA",X"00",X"9B",X"09",X"0B",X"00",X"00",X"09",X"0B",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"99",X"44",X"00",X"00",X"B0",X"44",X"00",X"00",X"BB",X"44",X"00",X"00",X"BB",X"99",
		X"00",X"99",X"BB",X"99",X"09",X"99",X"BB",X"99",X"04",X"99",X"99",X"09",X"04",X"0B",X"BB",X"09",
		X"44",X"BB",X"0B",X"00",X"49",X"00",X"BB",X"01",X"49",X"0B",X"F0",X"00",X"99",X"0B",X"00",X"B0",
		X"99",X"5B",X"00",X"B0",X"91",X"BB",X"00",X"B0",X"91",X"BB",X"40",X"B0",X"91",X"BB",X"40",X"B9",
		X"49",X"BB",X"40",X"BB",X"99",X"B0",X"00",X"BB",X"49",X"BB",X"B0",X"B0",X"99",X"B0",X"00",X"00",
		X"99",X"BB",X"B0",X"B0",X"99",X"BB",X"BB",X"BB",X"99",X"BB",X"BB",X"1B",X"44",X"1B",X"0B",X"19",
		X"04",X"10",X"00",X"14",X"04",X"11",X"00",X"94",X"04",X"11",X"90",X"94",X"00",X"9F",X"90",X"94",
		X"00",X"99",X"99",X"44",X"00",X"99",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",
		X"00",X"00",X"6F",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"60",X"00",X"00",X"06",X"60",X"00",
		X"00",X"06",X"66",X"00",X"00",X"06",X"60",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"60",X"00",
		X"00",X"00",X"6F",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",
		X"00",X"00",X"B0",X"00",X"00",X"0B",X"BB",X"00",X"00",X"0B",X"BB",X"00",X"00",X"BB",X"BB",X"00",
		X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",
		X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"0B",X"BB",X"00",X"00",X"0B",X"BB",X"00",
		X"00",X"00",X"B0",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"CB",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"F9",X"00",X"00",X"F0",
		X"F9",X"FF",X"FF",X"F0",X"F9",X"99",X"99",X"F0",X"99",X"99",X"99",X"9F",X"99",X"99",X"99",X"9F",
		X"99",X"F9",X"FF",X"9F",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"F9",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"F0",X"00",X"00",X"99",X"9F",X"00",X"00",X"99",X"99",X"00",
		X"00",X"9B",X"99",X"00",X"00",X"BB",X"C9",X"00",X"0F",X"00",X"C9",X"00",X"F9",X"00",X"C0",X"F0",
		X"99",X"99",X"00",X"F0",X"99",X"99",X"00",X"F0",X"99",X"99",X"99",X"F0",X"99",X"9B",X"99",X"F0",
		X"99",X"B0",X"99",X"F0",X"99",X"00",X"99",X"F0",X"99",X"00",X"B9",X"F0",X"BB",X"00",X"0B",X"B0",
		X"BB",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"FF",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",
		X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"09",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",X"F9",X"00",
		X"00",X"00",X"F9",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"09",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",
		X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"FF",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"95",X"00",
		X"00",X"99",X"95",X"00",X"00",X"99",X"95",X"00",X"00",X"99",X"96",X"00",X"00",X"99",X"96",X"00",
		X"00",X"55",X"95",X"00",X"00",X"55",X"65",X"80",X"00",X"55",X"95",X"88",X"99",X"99",X"99",X"88",
		X"99",X"99",X"96",X"99",X"F9",X"55",X"95",X"99",X"06",X"55",X"95",X"99",X"00",X"55",X"95",X"99",
		X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",X"99",X"00",
		X"00",X"F9",X"90",X"00",X"00",X"99",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"BB",X"0F",X"90",
		X"00",X"BB",X"9F",X"00",X"00",X"B9",X"FF",X"00",X"00",X"B9",X"BB",X"00",X"00",X"B9",X"F9",X"00",
		X"00",X"99",X"C9",X"99",X"00",X"B9",X"99",X"99",X"00",X"B9",X"99",X"99",X"00",X"B0",X"99",X"09",
		X"00",X"00",X"9B",X"09",X"00",X"00",X"FB",X"00",X"00",X"99",X"BB",X"00",X"00",X"00",X"B0",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"F0",X"00",X"00",X"99",X"9F",
		X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"B9",X"B9",X"00",X"00",X"0B",X"BB",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"BF",X"00",
		X"00",X"00",X"BF",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BB",X"FF",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",
		X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"FB",X"00",X"00",X"00",X"FB",X"00",X"00",X"00",X"FB",X"00",
		X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"04",X"44",
		X"00",X"44",X"44",X"44",X"00",X"00",X"40",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"40",X"00",
		X"00",X"00",X"40",X"00",X"00",X"00",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"40",X"00",X"00",
		X"00",X"40",X"00",X"00",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"00",X"40",X"04",
		X"00",X"00",X"40",X"04",X"00",X"44",X"40",X"04",X"00",X"44",X"40",X"04",X"00",X"00",X"44",X"44",
		X"00",X"44",X"44",X"44",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"40",
		X"00",X"04",X"44",X"44",X"00",X"44",X"40",X"04",X"00",X"00",X"40",X"04",X"00",X"44",X"40",X"04",
		X"00",X"44",X"40",X"04",X"00",X"00",X"44",X"44",X"00",X"00",X"04",X"40",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"44",X"04",X"40",X"00",X"44",X"44",X"44",X"00",X"00",X"40",X"04",X"00",X"00",X"40",X"04",
		X"00",X"00",X"40",X"04",X"00",X"00",X"40",X"04",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",
		X"00",X"00",X"40",X"04",X"00",X"00",X"40",X"04",X"00",X"00",X"40",X"04",X"00",X"00",X"40",X"04",
		X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",
		X"00",X"00",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"00",X"00",X"40",X"44",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"69",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"69",X"9F",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"69",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"0F",X"BF",X"00",X"00",X"FF",X"BB",X"0F",
		X"00",X"0F",X"BF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"BF",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BF",X"00",
		X"00",X"00",X"BF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",
		X"00",X"00",X"B0",X"00",X"00",X"0B",X"BB",X"00",X"00",X"0B",X"BB",X"00",X"00",X"BB",X"BB",X"00",
		X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",
		X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"0B",X"BB",X"00",X"00",X"0B",X"BB",X"00",
		X"00",X"00",X"B0",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"FB",X"00",X"00",X"00",X"FB",X"00",X"00",X"00",X"FB",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",
		X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"FF",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BF",X"00",
		X"00",X"00",X"BF",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"66",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"69",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"69",X"00",
		X"00",X"00",X"69",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",
		X"00",X"00",X"B0",X"00",X"00",X"0B",X"BB",X"00",X"00",X"0B",X"BB",X"00",X"00",X"BB",X"FB",X"00",
		X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",
		X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"0B",X"BB",X"00",X"00",X"0B",X"BB",X"00",
		X"00",X"00",X"B0",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0B",X"BB",X"00",X"00",X"B9",X"B9",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",
		X"00",X"00",X"99",X"9F",X"00",X"00",X"99",X"F0",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"BF",X"00",
		X"00",X"00",X"BF",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BB",X"FF",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",
		X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"FB",X"00",X"00",X"00",X"FB",X"00",X"00",X"00",X"FB",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"FB",X"00",X"00",X"00",X"FB",X"00",X"00",X"00",X"FB",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",
		X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"FF",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BF",X"00",
		X"00",X"00",X"BF",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",
		X"00",X"04",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"00",X"00",X"04",X"40",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"44",X"00",X"04",X"00",X"44",X"40",X"00",X"00",X"00",
		X"40",X"44",X"44",X"00",X"04",X"44",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",
		X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"FB",X"00",X"00",X"F0",
		X"FB",X"FF",X"FF",X"F0",X"FB",X"BB",X"BB",X"F0",X"BB",X"BB",X"BB",X"BF",X"BB",X"BB",X"BB",X"BF",
		X"BB",X"FB",X"FF",X"BF",X"BB",X"FB",X"FF",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"FB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"F0",X"00",X"00",X"11",X"1F",X"00",X"00",X"11",X"11",X"00",
		X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"0F",X"1B",X"11",X"00",X"F1",X"BB",X"B1",X"F0",
		X"BB",X"BB",X"BB",X"F0",X"BB",X"BB",X"BB",X"F0",X"BB",X"BB",X"BB",X"F0",X"BB",X"BF",X"BB",X"F0",
		X"BB",X"F0",X"BB",X"F0",X"BB",X"00",X"BB",X"00",X"FB",X"00",X"FB",X"00",X"0F",X"00",X"0F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"FB",X"00",X"00",X"F0",
		X"FB",X"FF",X"FF",X"F0",X"FB",X"BB",X"BB",X"F0",X"BB",X"BB",X"BB",X"BF",X"BB",X"BB",X"BB",X"BF",
		X"BB",X"FB",X"FF",X"BF",X"BB",X"FB",X"FF",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"00",X"00",X"00",X"66",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",
		X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"66",X"10",X"00",X"00",X"11",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"66",X"10",X"00",
		X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",
		X"00",X"66",X"10",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"00",X"00",X"60",X"10",X"00",
		X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",
		X"00",X"66",X"10",X"00",X"00",X"11",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"00",X"00",X"00",X"66",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",
		X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"66",X"10",X"00",X"00",X"11",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"66",X"10",X"00",
		X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",
		X"00",X"66",X"10",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"66",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"60",X"00",
		X"00",X"11",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"00",X"00",X"00",X"66",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",
		X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"66",X"10",X"00",X"00",X"11",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"66",X"10",X"00",
		X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",
		X"00",X"66",X"10",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"FB",X"BB",X"00",X"00",X"0F",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"F0",X"00",X"00",X"1B",X"F0",X"00",
		X"00",X"1B",X"F0",X"00",X"00",X"1B",X"F0",X"00",X"00",X"1B",X"00",X"00",X"00",X"1B",X"00",X"00",
		X"00",X"1B",X"00",X"00",X"00",X"1B",X"00",X"00",X"00",X"1B",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"1B",X"00",X"00",X"00",X"1B",X"00",X"00",X"00",X"1B",X"00",X"00",
		X"00",X"1B",X"00",X"00",X"00",X"1B",X"00",X"00",X"00",X"1B",X"F0",X"00",X"00",X"1B",X"F0",X"00",
		X"00",X"1B",X"F0",X"00",X"00",X"BB",X"F0",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"0F",X"BB",X"00",X"00",X"FB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",
		X"00",X"00",X"0F",X"BB",X"00",X"00",X"FB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",
		X"00",X"00",X"BB",X"BF",X"00",X"00",X"BB",X"F0",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"F0",X"00",X"00",X"BB",X"BF",
		X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"FB",X"BB",X"00",X"00",X"0F",X"BB",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"FF",X"F0",X"00",X"00",X"BB",X"F0",X"00",X"00",X"BB",X"F0",X"00",X"00",X"BB",X"F0",X"00",
		X"00",X"BB",X"F0",X"00",X"0F",X"BB",X"F0",X"00",X"FF",X"BB",X"F0",X"00",X"BB",X"BB",X"F0",X"00",
		X"BB",X"BB",X"F0",X"00",X"BB",X"FB",X"F0",X"00",X"00",X"FB",X"F0",X"00",X"00",X"FB",X"F0",X"00",
		X"00",X"FB",X"F0",X"00",X"00",X"FB",X"F0",X"00",X"00",X"FB",X"F0",X"00",X"00",X"FF",X"F0",X"00",
		X"00",X"BF",X"F0",X"00",X"00",X"FF",X"F0",X"00",X"00",X"FB",X"F0",X"00",X"00",X"FB",X"F0",X"00",
		X"00",X"FB",X"F0",X"00",X"00",X"FB",X"F0",X"00",X"BB",X"FB",X"F0",X"00",X"BB",X"BB",X"F0",X"00",
		X"BB",X"BB",X"F0",X"00",X"FF",X"BB",X"F0",X"00",X"0F",X"BB",X"F0",X"00",X"00",X"BB",X"F0",X"00",
		X"00",X"BB",X"F0",X"00",X"00",X"BB",X"F0",X"00",X"00",X"BB",X"F0",X"00",X"00",X"FF",X"F0",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"60",X"00",X"00",X"66",X"60",X"00",X"00",X"66",X"60",X"00",X"00",X"66",X"60",
		X"00",X"00",X"66",X"60",X"00",X"00",X"66",X"60",X"00",X"00",X"66",X"00",X"00",X"00",X"6B",X"00",
		X"00",X"00",X"6B",X"00",X"00",X"00",X"6B",X"00",X"00",X"66",X"FF",X"00",X"00",X"66",X"66",X"00",
		X"00",X"66",X"FF",X"00",X"00",X"00",X"6B",X"00",X"00",X"00",X"6B",X"00",X"00",X"00",X"6B",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"60",X"00",X"00",X"66",X"60",X"00",X"00",X"66",X"60",
		X"00",X"00",X"66",X"60",X"00",X"00",X"66",X"60",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"FF",X"F0",X"00",X"00",X"BB",X"F0",X"00",X"00",X"BB",X"F0",X"00",X"00",X"BB",X"F0",X"00",
		X"00",X"BB",X"F0",X"00",X"0F",X"BB",X"F0",X"00",X"FF",X"BB",X"F0",X"00",X"BB",X"BB",X"F0",X"00",
		X"BB",X"BB",X"F0",X"00",X"BB",X"FB",X"F0",X"00",X"00",X"FB",X"F0",X"00",X"00",X"FB",X"F0",X"00",
		X"00",X"FB",X"F0",X"00",X"00",X"FB",X"F0",X"00",X"00",X"FB",X"F0",X"00",X"00",X"FF",X"F0",X"00",
		X"00",X"BF",X"F0",X"00",X"00",X"FF",X"F0",X"00",X"00",X"FB",X"F0",X"00",X"00",X"FB",X"F0",X"00",
		X"00",X"FB",X"F0",X"00",X"00",X"FB",X"F0",X"00",X"BB",X"FB",X"F0",X"00",X"BB",X"BB",X"F0",X"00",
		X"BB",X"BB",X"F0",X"00",X"FF",X"BB",X"F0",X"00",X"0F",X"BB",X"F0",X"00",X"00",X"BB",X"F0",X"00",
		X"00",X"BB",X"F0",X"00",X"00",X"BB",X"F0",X"00",X"00",X"BB",X"F0",X"00",X"00",X"FF",X"F0",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"40",X"04",X"00",X"44",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"44",X"40",X"04",
		X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"44",X"00",X"00",X"44",X"44",
		X"00",X"00",X"40",X"00",X"00",X"00",X"40",X"00",X"00",X"44",X"40",X"00",X"00",X"44",X"40",X"00",
		X"00",X"40",X"44",X"44",X"00",X"40",X"44",X"44",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"00",X"00",X"04",X"40",X"00",X"00",X"44",X"40",X"00",X"44",X"04",X"00",X"00",X"44",
		X"00",X"40",X"00",X"04",X"00",X"04",X"00",X"04",X"44",X"04",X"00",X"04",X"00",X"40",X"00",X"04",
		X"44",X"04",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"04",X"00",X"00",X"00",X"40",X"00",X"00",
		X"00",X"04",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"44",X"00",X"04",X"00",X"44",X"00",X"04",
		X"00",X"04",X"44",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"40",X"00",X"00",X"04",X"44",X"44",
		X"00",X"44",X"44",X"44",X"00",X"00",X"40",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"44",X"44",X"00",X"00",X"44",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"44",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"44",X"40",X"04",X"00",X"44",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"40",X"04",
		X"00",X"00",X"40",X"04",X"00",X"44",X"40",X"04",X"00",X"44",X"40",X"04",X"00",X"00",X"44",X"44",
		X"00",X"44",X"44",X"40",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"B0",X"00",X"00",X"BB",X"BB",X"00",
		X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"FB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"BB",X"FB",X"00",X"BB",X"BB",X"00",
		X"00",X"BB",X"BB",X"00",X"00",X"BB",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"BB",
		X"00",X"00",X"50",X"BB",X"00",X"00",X"10",X"FB",X"00",X"00",X"11",X"50",X"00",X"00",X"11",X"00",
		X"00",X"0C",X"11",X"50",X"00",X"00",X"11",X"00",X"00",X"0C",X"10",X"50",X"00",X"00",X"10",X"00",
		X"00",X"0C",X"15",X"00",X"00",X"00",X"10",X"10",X"00",X"CC",X"11",X"11",X"00",X"00",X"10",X"10",
		X"00",X"C0",X"11",X"50",X"00",X"00",X"10",X"00",X"00",X"C0",X"11",X"05",X"00",X"00",X"11",X"00",
		X"00",X"C1",X"11",X"05",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"F5",X"00",X"00",X"10",X"BF",
		X"00",X"00",X"05",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"05",X"BB",X"00",X"00",X"00",X"00",
		X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"40",X"04",
		X"00",X"40",X"40",X"04",X"00",X"44",X"40",X"04",X"00",X"44",X"44",X"44",X"00",X"40",X"44",X"44",
		X"00",X"00",X"44",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"44",
		X"00",X"04",X"44",X"44",X"00",X"44",X"40",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"40",X"00",
		X"00",X"00",X"40",X"04",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"44",X"00",X"00",
		X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"04",X"40",
		X"00",X"04",X"44",X"44",X"00",X"00",X"40",X"04",X"00",X"00",X"40",X"04",X"00",X"04",X"40",X"04",
		X"00",X"44",X"40",X"04",X"00",X"00",X"44",X"44",X"00",X"00",X"04",X"40",X"00",X"44",X"00",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0B",X"00",X"00",X"00",X"9B",X"B9",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",
		X"00",X"BB",X"BB",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"BB",X"B0",X"00",X"BB",X"BB",X"00",
		X"00",X"BB",X"BB",X"00",X"00",X"9B",X"B9",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"CB",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"66",X"F0",X"00",X"00",X"66",X"66",X"00",X"00",X"66",X"BB",X"00",
		X"00",X"B6",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"60",X"66",X"00",X"00",X"00",X"0B",X"00",
		X"00",X"66",X"B0",X"00",X"00",X"66",X"B0",X"00",X"00",X"6F",X"B0",X"00",X"00",X"66",X"B0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",
		X"00",X"00",X"6F",X"00",X"00",X"00",X"60",X"00",X"00",X"06",X"60",X"00",X"00",X"06",X"66",X"00",
		X"00",X"06",X"60",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"6F",X"00",
		X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",
		X"00",X"00",X"6F",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"60",X"00",X"00",X"06",X"60",X"00",
		X"00",X"06",X"66",X"00",X"00",X"06",X"60",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"60",X"00",
		X"00",X"00",X"6F",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",
		X"00",X"05",X"CC",X"CC",X"00",X"00",X"55",X"CC",X"0C",X"CC",X"55",X"CC",X"00",X"C0",X"55",X"CC",
		X"00",X"05",X"55",X"00",X"00",X"55",X"55",X"00",X"00",X"55",X"55",X"00",X"00",X"55",X"55",X"00",
		X"00",X"55",X"B5",X"00",X"00",X"55",X"55",X"00",X"00",X"55",X"55",X"00",X"00",X"55",X"55",X"00",
		X"00",X"C5",X"55",X"00",X"0C",X"CC",X"55",X"00",X"00",X"00",X"55",X"CC",X"00",X"55",X"55",X"CC",
		X"00",X"05",X"CC",X"CC",X"00",X"00",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"0D",X"00",X"80",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",
		X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"F0",X"00",X"C0",X"00",X"00",
		X"00",X"0F",X"00",X"D0",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"00",X"20",X"00",X"22",X"55",X"22",X"00",X"22",X"55",X"00",X"00",X"25",X"55",X"55",
		X"00",X"50",X"55",X"55",X"00",X"55",X"55",X"55",X"05",X"55",X"55",X"55",X"05",X"55",X"55",X"55",
		X"55",X"55",X"F5",X"55",X"00",X"55",X"AF",X"00",X"20",X"55",X"FA",X"20",X"22",X"55",X"FF",X"22",
		X"22",X"55",X"FA",X"22",X"22",X"55",X"FF",X"22",X"20",X"55",X"FA",X"20",X"00",X"55",X"AF",X"00",
		X"55",X"55",X"F5",X"55",X"05",X"55",X"55",X"55",X"05",X"55",X"55",X"55",X"00",X"55",X"55",X"55",
		X"00",X"50",X"55",X"55",X"00",X"20",X"00",X"05",X"00",X"22",X"55",X"00",X"00",X"22",X"55",X"22",
		X"00",X"00",X"55",X"20",X"00",X"05",X"55",X"00",X"00",X"05",X"55",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"66",X"10",X"00",
		X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",
		X"00",X"60",X"10",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"00",X"00",X"00",X"66",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",
		X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"66",X"10",X"00",X"00",X"11",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"66",X"10",X"00",
		X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",
		X"00",X"66",X"10",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"66",X"10",X"00",
		X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",
		X"00",X"66",X"10",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"00",X"00",X"00",X"66",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",
		X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"66",X"10",X"00",X"00",X"11",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"66",X"10",X"00",
		X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",
		X"00",X"66",X"10",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"60",X"00",X"00",X"06",X"60",X"00",X"00",X"06",X"60",X"00",X"00",X"66",X"60",
		X"00",X"00",X"66",X"60",X"00",X"00",X"66",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"6B",X"00",
		X"00",X"66",X"6B",X"00",X"00",X"66",X"6B",X"00",X"00",X"66",X"FF",X"00",X"00",X"66",X"66",X"00",
		X"00",X"66",X"FF",X"00",X"00",X"66",X"6B",X"00",X"00",X"66",X"6B",X"00",X"00",X"00",X"6B",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"60",X"00",X"00",X"66",X"60",X"00",X"00",X"66",X"60",
		X"00",X"00",X"66",X"60",X"00",X"00",X"06",X"60",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"66",X"00",X"00",X"66",X"B0",X"00",
		X"00",X"B6",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"60",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"66",X"B0",X"00",X"00",X"66",X"B0",X"00",X"00",X"6F",X"B0",X"00",X"00",X"66",X"B0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"4F",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"CB",X"00",X"90",X"00",X"CC",X"99",X"99",X"00",X"0C",X"99",X"99",
		X"00",X"0C",X"99",X"99",X"00",X"CC",X"99",X"99",X"00",X"CB",X"00",X"90",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"05",X"05",X"05",X"00",X"00",X"00",X"00",X"00",X"05",X"05",X"05",X"00",X"00",X"00",X"00",
		X"0B",X"55",X"05",X"05",X"BB",X"00",X"00",X"00",X"BB",X"50",X"05",X"05",X"00",X"01",X"00",X"00",
		X"05",X"11",X"CC",X"05",X"00",X"11",X"00",X"00",X"05",X"11",X"CC",X"05",X"00",X"01",X"C0",X"00",
		X"00",X"51",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"CC",X"00",X"00",X"00",X"00",X"00",
		X"50",X"10",X"0C",X"00",X"00",X"00",X"00",X"00",X"50",X"11",X"0C",X"50",X"00",X"11",X"00",X"00",
		X"50",X"11",X"11",X"50",X"00",X"01",X"00",X"00",X"50",X"05",X"50",X"50",X"00",X"00",X"00",X"00",
		X"0B",X"55",X"50",X"50",X"0B",X"00",X"00",X"00",X"05",X"50",X"50",X"50",X"00",X"00",X"00",X"00",
		X"00",X"50",X"50",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"66",X"00",
		X"00",X"AA",X"AA",X"00",X"00",X"0A",X"AB",X"00",X"06",X"00",X"B9",X"00",X"06",X"0F",X"96",X"00",
		X"06",X"90",X"B9",X"00",X"06",X"09",X"BA",X"00",X"00",X"FF",X"BB",X"00",X"00",X"0B",X"AA",X"00",
		X"00",X"BB",X"0F",X"00",X"00",X"FB",X"B5",X"00",X"00",X"BB",X"06",X"00",X"00",X"BB",X"96",X"00",
		X"00",X"FF",X"6B",X"00",X"00",X"F0",X"66",X"00",X"00",X"F9",X"66",X"00",X"00",X"00",X"66",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"06",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"9B",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",
		X"BB",X"00",X"00",X"00",X"BB",X"F0",X"00",X"00",X"B0",X"B0",X"B0",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"09",X"00",
		X"00",X"00",X"99",X"00",X"00",X"0B",X"00",X"00",X"BB",X"9B",X"00",X"00",X"0B",X"90",X"0F",X"00",
		X"BB",X"9B",X"FF",X"00",X"BB",X"9B",X"F9",X"00",X"00",X"90",X"FF",X"BB",X"FF",X"90",X"B9",X"9B",
		X"00",X"00",X"99",X"00",X"00",X"0F",X"F9",X"00",X"BB",X"BB",X"FF",X"00",X"B0",X"BB",X"9F",X"00",
		X"B0",X"BB",X"FF",X"00",X"90",X"9B",X"FF",X"90",X"00",X"0B",X"BB",X"00",X"00",X"0B",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"9B",X"0A",X"00",X"00",X"00",X"06",X"00",X"0B",X"00",X"66",X"00",
		X"BB",X"99",X"AA",X"00",X"BB",X"A9",X"9A",X"00",X"B0",X"A9",X"9A",X"00",X"00",X"AB",X"99",X"00",
		X"00",X"BB",X"99",X"00",X"09",X"90",X"0A",X"00",X"99",X"99",X"AA",X"00",X"09",X"AA",X"0A",X"00",
		X"00",X"A5",X"AA",X"00",X"00",X"AA",X"00",X"00",X"BB",X"AA",X"99",X"00",X"0B",X"A5",X"09",X"00",
		X"BB",X"A5",X"A9",X"00",X"BB",X"AA",X"96",X"00",X"00",X"9A",X"96",X"BB",X"FF",X"9A",X"B9",X"9B",
		X"00",X"00",X"AA",X"00",X"00",X"0F",X"AA",X"00",X"BB",X"AA",X"AA",X"00",X"B0",X"AA",X"AA",X"00",
		X"B0",X"AA",X"AA",X"00",X"90",X"9B",X"F6",X"90",X"00",X"99",X"BB",X"00",X"00",X"0B",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"99",X"40",X"04",X"99",X"99",X"40",X"04",X"99",X"99",X"40",X"04",X"99",X"99",X"40",
		X"94",X"90",X"9B",X"44",X"94",X"90",X"99",X"99",X"90",X"00",X"0B",X"94",X"99",X"90",X"BB",X"94",
		X"49",X"B0",X"FF",X"99",X"99",X"BB",X"F0",X"09",X"91",X"BB",X"00",X"99",X"99",X"BB",X"0F",X"99",
		X"11",X"BB",X"0F",X"99",X"10",X"55",X"00",X"99",X"09",X"F0",X"00",X"00",X"10",X"F0",X"50",X"09",
		X"00",X"F5",X"00",X"B0",X"00",X"00",X"50",X"00",X"00",X"99",X"00",X"00",X"0B",X"90",X"00",X"09",
		X"9B",X"9B",X"FF",X"00",X"9B",X"BB",X"BB",X"B9",X"99",X"BB",X"BB",X"B4",X"BB",X"BB",X"BB",X"99",
		X"BB",X"00",X"BB",X"94",X"99",X"11",X"B0",X"94",X"99",X"91",X"00",X"44",X"99",X"99",X"00",X"00",
		X"00",X"F9",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"86",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"60",X"00",X"00",X"60",X"60",X"00",
		X"00",X"B0",X"66",X"00",X"00",X"60",X"60",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"60",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",
		X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"B0",X"00",
		X"00",X"BB",X"B0",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BF",X"BB",X"00",
		X"00",X"BB",X"B0",X"00",X"00",X"BB",X"B0",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",
		X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",
		X"00",X"BB",X"B0",X"00",X"00",X"BB",X"B0",X"00",X"00",X"BB",X"B0",X"00",X"00",X"BB",X"B0",X"00",
		X"00",X"BB",X"B0",X"00",X"00",X"BC",X"B0",X"00",X"00",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"09",X"00",X"0F",X"00",X"09",X"00",
		X"0F",X"00",X"09",X"00",X"F9",X"00",X"09",X"00",X"F9",X"00",X"09",X"00",X"F9",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"09",X"00",X"99",X"00",X"09",X"00",
		X"99",X"FF",X"F9",X"00",X"99",X"9F",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"FF",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"F0",X"99",X"99",X"99",X"F0",X"99",X"99",X"99",X"F0",
		X"FF",X"FF",X"FF",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"9B",X"00",X"00",X"00",X"9B",X"00",X"00",
		X"00",X"9B",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"B0",X"F0",X"00",
		X"0F",X"B0",X"9F",X"00",X"F9",X"B0",X"99",X"00",X"99",X"00",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"9B",X"99",X"00",X"99",X"B0",X"99",X"00",X"99",X"00",X"99",X"00",
		X"99",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"BB",X"00",X"BB",X"00",
		X"BB",X"00",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"FF",X"00",
		X"00",X"0F",X"99",X"00",X"00",X"0F",X"99",X"F0",X"00",X"0F",X"99",X"9F",X"00",X"0F",X"99",X"99",
		X"00",X"0F",X"99",X"99",X"00",X"0F",X"99",X"99",X"00",X"0F",X"99",X"99",X"00",X"0F",X"9F",X"00",
		X"00",X"0F",X"9F",X"00",X"00",X"0F",X"9F",X"00",X"00",X"0F",X"9F",X"00",X"00",X"0F",X"9F",X"00",
		X"00",X"0F",X"9F",X"00",X"00",X"0F",X"9F",X"00",X"00",X"0F",X"9F",X"00",X"00",X"0F",X"FF",X"00",
		X"00",X"0F",X"FF",X"00",X"00",X"0F",X"9F",X"00",X"00",X"0F",X"9F",X"00",X"00",X"0F",X"9F",X"00",
		X"00",X"0F",X"9F",X"00",X"00",X"0F",X"9F",X"00",X"00",X"0F",X"9F",X"00",X"00",X"0F",X"9F",X"00",
		X"00",X"0F",X"9F",X"00",X"00",X"0F",X"99",X"99",X"00",X"0F",X"99",X"99",X"00",X"0F",X"99",X"99",
		X"00",X"0F",X"99",X"99",X"00",X"0F",X"99",X"FF",X"00",X"0F",X"99",X"F0",X"00",X"0F",X"99",X"00",
		X"00",X"0F",X"FF",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"F0",X"00",
		X"00",X"99",X"59",X"00",X"00",X"99",X"59",X"00",X"00",X"99",X"99",X"00",X"09",X"99",X"69",X"00",
		X"09",X"59",X"55",X"00",X"66",X"56",X"55",X"00",X"66",X"56",X"55",X"00",X"99",X"99",X"69",X"88",
		X"99",X"99",X"69",X"98",X"99",X"59",X"55",X"98",X"66",X"59",X"55",X"99",X"F6",X"56",X"55",X"99",
		X"0F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"9B",X"00",
		X"00",X"99",X"BB",X"00",X"00",X"99",X"BB",X"00",X"00",X"9B",X"99",X"00",X"00",X"BC",X"99",X"00",
		X"00",X"BC",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BF",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"99",X"00",X"90",X"00",X"99",X"B0",X"00",X"00",X"9B",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0B",X"FF",X"00",X"00",X"0B",X"99",X"00",X"00",X"0B",X"99",X"00",X"00",X"0B",X"99",X"00",
		X"00",X"0B",X"99",X"00",X"00",X"0B",X"99",X"00",X"00",X"0B",X"99",X"00",X"00",X"0B",X"99",X"00",
		X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"F0",X"00",X"00",X"90",X"9F",X"00",X"00",X"90",X"99",X"00",X"00",X"99",X"BB",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"0F",X"FF",X"00",X"00",X"0F",X"BB",X"00",X"00",X"0F",X"BB",X"00",X"00",X"0F",X"BB",X"00",
		X"00",X"0F",X"BB",X"00",X"00",X"0F",X"BB",X"F0",X"00",X"0F",X"BB",X"FF",X"00",X"0F",X"BB",X"BB",
		X"00",X"0F",X"BB",X"BB",X"00",X"0F",X"BF",X"BB",X"00",X"0F",X"BF",X"00",X"00",X"0F",X"BF",X"00",
		X"00",X"0F",X"BF",X"00",X"00",X"0F",X"BF",X"00",X"00",X"0F",X"BF",X"00",X"00",X"0F",X"FF",X"00",
		X"04",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"04",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",
		X"04",X"00",X"00",X"00",X"04",X"00",X"44",X"00",X"04",X"00",X"44",X"00",X"04",X"00",X"00",X"00",
		X"04",X"00",X"00",X"00",X"04",X"44",X"40",X"00",X"04",X"44",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"44",X"00",X"00",X"04",X"44",X"00",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"44",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"04",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"44",X"00",X"00",
		X"04",X"44",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"44",X"44",X"00",X"04",X"44",X"44",X"00",X"04",X"00",X"00",X"00",X"04",X"00",X"00",X"00",
		X"04",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"04",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"40",X"00",X"04",X"44",X"40",X"00",
		X"04",X"04",X"00",X"00",X"04",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"04",X"00",X"00",X"00",
		X"04",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"40",X"00",X"00",X"00",X"44",X"00",X"00",X"04",X"04",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"04",X"44",X"04",X"00",X"04",X"00",X"44",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"96",X"00",
		X"00",X"00",X"96",X"00",X"00",X"00",X"96",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"96",X"00",X"00",X"00",X"66",X"F0",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",
		X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",X"0F",X"FF",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",
		X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"B0",X"00",
		X"00",X"BB",X"B0",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",
		X"00",X"BB",X"B0",X"00",X"00",X"BB",X"B0",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",
		X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"0F",X"FB",X"00",X"00",X"0F",X"FF",X"00",X"00",X"0F",X"BF",X"00",X"00",X"0F",X"BF",X"00",
		X"00",X"0F",X"BF",X"00",X"00",X"0F",X"BF",X"00",X"00",X"0F",X"BF",X"BB",X"00",X"0F",X"BB",X"BB",
		X"00",X"0F",X"BB",X"BB",X"00",X"0F",X"BB",X"FF",X"00",X"0F",X"BB",X"F0",X"00",X"0F",X"BB",X"00",
		X"00",X"0F",X"BB",X"00",X"00",X"0F",X"BB",X"00",X"00",X"0F",X"BB",X"00",X"00",X"0F",X"FF",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"96",X"F0",X"00",X"00",X"66",X"F0",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"96",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0B",X"00",X"00",
		X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BF",X"00",X"00",X"00",X"FB",X"B0",X"00",
		X"00",X"BB",X"B0",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",
		X"00",X"BB",X"B0",X"00",X"00",X"BB",X"B0",X"00",X"00",X"BB",X"00",X"00",X"00",X"BF",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",
		X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"00",X"99",X"BB",X"00",X"00",X"90",X"99",X"00",X"00",X"90",X"9F",X"00",X"00",X"00",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",
		X"00",X"0B",X"99",X"00",X"00",X"0B",X"99",X"00",X"00",X"0B",X"99",X"00",X"00",X"0B",X"99",X"00",
		X"00",X"0B",X"99",X"00",X"00",X"0B",X"99",X"00",X"00",X"0B",X"99",X"00",X"00",X"0B",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"0F",X"FF",X"00",X"00",X"0F",X"BB",X"00",X"00",X"0F",X"BB",X"00",X"00",X"0F",X"BB",X"00",
		X"00",X"0F",X"BB",X"00",X"00",X"0F",X"BB",X"F0",X"00",X"0F",X"BB",X"FF",X"00",X"0F",X"BB",X"BB",
		X"00",X"0F",X"BB",X"BB",X"00",X"0F",X"BF",X"BB",X"00",X"0F",X"BF",X"00",X"00",X"0F",X"BF",X"00",
		X"00",X"0F",X"BF",X"00",X"00",X"0F",X"BF",X"00",X"00",X"0F",X"BF",X"00",X"00",X"0F",X"FF",X"00",
		X"00",X"0F",X"FB",X"00",X"00",X"0F",X"FF",X"00",X"00",X"0F",X"BF",X"00",X"00",X"0F",X"BF",X"00",
		X"00",X"0F",X"BF",X"00",X"00",X"0F",X"BF",X"00",X"00",X"0F",X"BF",X"BB",X"00",X"0F",X"BB",X"BB",
		X"00",X"0F",X"BB",X"BB",X"00",X"0F",X"BB",X"FF",X"00",X"0F",X"BB",X"F0",X"00",X"0F",X"BB",X"00",
		X"00",X"0F",X"BB",X"00",X"00",X"0F",X"BB",X"00",X"00",X"0F",X"BB",X"00",X"00",X"0F",X"FF",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"04",X"44",X"00",X"00",X"04",X"00",X"00",X"00",
		X"04",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"04",X"04",X"00",X"00",
		X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"44",X"00",X"00",
		X"04",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"00",X"00",X"00",X"04",X"00",X"00",X"04",X"00",X"00",X"00",X"04",X"00",X"00",X"00",
		X"04",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"04",X"00",X"00",X"00",
		X"00",X"04",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"00",X"00",X"00",X"04",X"40",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"04",X"00",X"00",
		X"00",X"04",X"00",X"00",X"00",X"44",X"00",X"00",X"04",X"40",X"00",X"00",X"00",X"00",X"44",X"00",
		X"00",X"40",X"40",X"00",X"40",X"44",X"00",X"00",X"40",X"04",X"40",X"00",X"04",X"04",X"44",X"00",
		X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"44",X"00",X"00",X"04",X"44",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",
		X"04",X"44",X"00",X"00",X"04",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"04",X"00",X"00",X"00",
		X"04",X"00",X"00",X"00",X"04",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0B",X"00",X"0F",X"00",X"0B",X"00",
		X"0F",X"00",X"0B",X"00",X"FB",X"00",X"0B",X"00",X"FB",X"00",X"0B",X"00",X"FB",X"00",X"00",X"00",
		X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"0B",X"00",X"BB",X"00",X"0B",X"00",
		X"BB",X"FF",X"FB",X"00",X"BB",X"BF",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"FF",X"BB",X"00",
		X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"F0",X"BB",X"BB",X"BB",X"F0",X"BB",X"BB",X"BB",X"F0",
		X"FF",X"FF",X"FF",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"F0",X"00",
		X"0F",X"11",X"1F",X"00",X"F1",X"11",X"11",X"00",X"11",X"BB",X"11",X"00",X"11",X"BB",X"11",X"00",
		X"BB",X"BB",X"BB",X"00",X"BB",X"BF",X"BB",X"00",X"BB",X"F0",X"BB",X"00",X"BB",X"00",X"BB",X"00",
		X"BB",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"00",
		X"FF",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0B",X"00",X"0F",X"00",X"0B",X"00",
		X"0F",X"00",X"0B",X"00",X"FB",X"00",X"0B",X"00",X"FB",X"00",X"0B",X"00",X"FB",X"00",X"00",X"00",
		X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"0B",X"00",X"BB",X"00",X"0B",X"00",
		X"BB",X"FF",X"FB",X"00",X"BB",X"BF",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"FF",X"BB",X"00",
		X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"F0",X"BB",X"BB",X"BB",X"F0",X"BB",X"BB",X"BB",X"F0",
		X"FF",X"FF",X"FF",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"11",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"66",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",
		X"00",X"61",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"11",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"66",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"66",X"00",X"00",
		X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"61",X"00",X"00",
		X"00",X"11",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"11",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"66",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"BB",X"F0",X"00",X"00",X"BB",X"BF",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",
		X"FB",X"BB",X"00",X"00",X"0F",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"0F",X"BB",X"00",X"00",X"FB",X"BB",X"00",X"00",
		X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BF",X"00",X"00",X"BB",X"F0",X"00",X"00",
		X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BF",X"00",X"00",X"BB",X"F0",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"0F",X"BB",X"00",X"00",X"0F",X"B1",X"00",
		X"00",X"0F",X"B1",X"00",X"00",X"0F",X"B1",X"00",X"00",X"00",X"B1",X"00",X"00",X"00",X"B1",X"00",
		X"00",X"00",X"B1",X"00",X"00",X"00",X"B1",X"00",X"00",X"00",X"B1",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"B1",X"00",X"00",X"00",X"B1",X"00",X"00",X"00",X"B1",X"00",
		X"00",X"00",X"B1",X"00",X"00",X"00",X"B1",X"00",X"00",X"0F",X"B1",X"00",X"00",X"0F",X"B1",X"00",
		X"00",X"0F",X"B1",X"00",X"00",X"0F",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BB",X"F0",X"00",X"00",X"BB",X"BF",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"FB",X"00",X"00",
		X"00",X"FB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"FF",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",
		X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BF",X"00",X"00",X"00",X"BF",X"00",X"00",X"00",X"BF",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"BF",X"00",X"00",X"00",X"BF",X"00",X"00",X"00",X"BF",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",
		X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"FF",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"FB",X"00",X"00",
		X"00",X"FB",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"B6",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",
		X"66",X"00",X"00",X"00",X"66",X"F0",X"00",X"00",X"66",X"66",X"F0",X"00",X"66",X"F6",X"66",X"00",
		X"66",X"66",X"F0",X"00",X"66",X"F0",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"60",X"00",X"00",X"00",X"B6",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"FB",X"00",X"00",
		X"00",X"FB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"FF",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",
		X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BF",X"00",X"00",X"00",X"BF",X"00",X"00",X"00",X"BF",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"BF",X"00",X"00",X"00",X"BF",X"00",X"00",X"00",X"BF",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",
		X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"FF",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"FB",X"00",X"00",
		X"00",X"FB",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"04",X"44",X"00",X"00",
		X"04",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"44",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",
		X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"00",X"44",X"00",X"44",X"40",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"44",X"44",X"00",
		X"00",X"00",X"44",X"00",X"04",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"04",X"44",X"44",X"00",X"04",X"00",X"44",X"00",
		X"04",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"04",X"44",X"00",X"00",
		X"04",X"44",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",
		X"04",X"44",X"00",X"00",X"04",X"44",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"44",X"00",X"00",X"04",X"44",X"00",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"44",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"04",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0B",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"B0",X"00",
		X"00",X"BB",X"BB",X"00",X"0B",X"BB",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",
		X"00",X"BB",X"B0",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"0B",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"50",X"50",X"50",X"00",X"00",X"00",X"00",X"00",X"50",X"50",X"50",X"00",X"00",X"00",X"00",X"00",
		X"50",X"50",X"55",X"B0",X"00",X"00",X"00",X"BB",X"50",X"50",X"05",X"BB",X"00",X"00",X"1B",X"00",
		X"50",X"CC",X"11",X"50",X"00",X"00",X"11",X"00",X"50",X"CC",X"11",X"50",X"00",X"0C",X"10",X"00",
		X"00",X"CC",X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"11",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"01",X"05",X"00",X"00",X"00",X"00",X"05",X"C0",X"11",X"05",X"00",X"00",X"11",X"00",
		X"05",X"11",X"11",X"05",X"00",X"00",X"10",X"00",X"05",X"05",X"50",X"05",X"00",X"00",X"00",X"00",
		X"05",X"05",X"55",X"B0",X"00",X"00",X"00",X"B0",X"05",X"05",X"05",X"50",X"00",X"00",X"00",X"00",
		X"05",X"05",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"44",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"44",X"00",X"04",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"00",X"00",X"00",X"40",X"00",X"00",X"04",X"40",X"00",X"00",
		X"04",X"40",X"00",X"00",X"04",X"40",X"44",X"00",X"00",X"40",X"44",X"00",X"00",X"44",X"00",X"00",
		X"00",X"44",X"00",X"00",X"04",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"40",X"00",
		X"00",X"44",X"40",X"00",X"00",X"04",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"00",X"44",X"00",X"04",X"00",X"44",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",
		X"BB",X"BB",X"BB",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"0F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"BB",X"BB",X"B0",X"00",X"BB",X"BB",X"00",
		X"00",X"BB",X"BB",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",
		X"00",X"BB",X"B0",X"00",X"00",X"BB",X"B0",X"00",X"00",X"BB",X"B0",X"00",X"00",X"BB",X"B0",X"00",
		X"00",X"BB",X"B0",X"00",X"00",X"BC",X"B0",X"00",X"00",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"66",X"00",
		X"00",X"60",X"66",X"00",X"00",X"60",X"66",X"00",X"00",X"66",X"66",X"00",X"00",X"BB",X"B6",X"00",
		X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"60",X"00",X"00",X"6B",X"60",X"00",
		X"00",X"00",X"06",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"06",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",
		X"00",X"00",X"60",X"00",X"00",X"00",X"60",X"00",X"00",X"60",X"60",X"00",X"00",X"B0",X"66",X"00",
		X"00",X"60",X"60",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"66",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"60",X"00",X"00",X"60",X"60",X"00",
		X"00",X"B0",X"66",X"00",X"00",X"60",X"60",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"60",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",
		X"0C",X"5C",X"55",X"00",X"CC",X"05",X"55",X"00",X"CC",X"55",X"55",X"C0",X"00",X"55",X"5C",X"CC",
		X"00",X"55",X"55",X"00",X"00",X"55",X"55",X"00",X"00",X"55",X"55",X"00",X"00",X"55",X"55",X"00",
		X"00",X"55",X"55",X"00",X"00",X"55",X"55",X"00",X"00",X"55",X"55",X"00",X"00",X"55",X"55",X"00",
		X"00",X"55",X"55",X"00",X"CC",X"55",X"00",X"00",X"CC",X"05",X"0C",X"CC",X"0C",X"05",X"50",X"C0",
		X"00",X"0C",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"04",X"F0",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"40",
		X"00",X"F0",X"00",X"F0",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"F0",X"00",X"0F",X"00",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"00",X"00",X"05",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"25",X"22",X"00",X"00",X"55",X"52",X"00",X"05",X"55",X"50",X"00",
		X"55",X"55",X"50",X"50",X"55",X"55",X"55",X"50",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"00",X"5F",X"55",X"00",X"00",X"5A",X"55",X"00",X"02",X"5F",X"55",X"02",
		X"C2",X"5A",X"55",X"C2",X"02",X"5F",X"55",X"02",X"00",X"5A",X"55",X"00",X"00",X"5F",X"55",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"50",X"50",
		X"55",X"55",X"50",X"50",X"00",X"00",X"00",X"00",X"00",X"55",X"02",X"00",X"02",X"25",X"22",X"00",
		X"00",X"05",X"50",X"00",X"00",X"55",X"55",X"00",X"00",X"55",X"55",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"61",X"00",X"00",
		X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",
		X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"11",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"66",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"61",X"00",X"00",
		X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",
		X"00",X"61",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"11",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"66",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"B6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"F0",X"00",X"00",X"F6",X"66",X"00",
		X"00",X"66",X"F0",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"B6",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"06",X"00",
		X"00",X"66",X"66",X"00",X"00",X"66",X"66",X"00",X"00",X"60",X"66",X"00",X"00",X"B0",X"B6",X"00",
		X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"60",X"00",X"00",X"60",X"60",X"00",
		X"00",X"00",X"06",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"06",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"F0",X"00",X"00",X"F0",X"0F",X"00",
		X"00",X"04",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"90",
		X"00",X"99",X"99",X"90",X"00",X"BB",X"99",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",
		X"BB",X"05",X"00",X"00",X"B0",X"01",X"00",X"00",X"05",X"11",X"00",X"00",X"00",X"11",X"00",X"00",
		X"05",X"11",X"C0",X"00",X"00",X"11",X"00",X"00",X"05",X"01",X"C0",X"00",X"00",X"01",X"00",X"00",
		X"00",X"51",X"C0",X"00",X"01",X"01",X"00",X"00",X"11",X"11",X"CC",X"00",X"01",X"01",X"00",X"00",
		X"05",X"11",X"0C",X"00",X"00",X"01",X"00",X"00",X"50",X"11",X"0C",X"00",X"00",X"11",X"00",X"00",
		X"50",X"11",X"1C",X"00",X"00",X"11",X"00",X"00",X"50",X"11",X"00",X"00",X"0B",X"01",X"00",X"00",
		X"B0",X"50",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"50",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"06",X"00",X"00",
		X"00",X"06",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"66",X"00",X"00",X"A6",X"06",X"00",
		X"00",X"AA",X"09",X"00",X"00",X"AB",X"99",X"00",X"66",X"BB",X"9A",X"00",X"06",X"FB",X"0A",X"00",
		X"66",X"0F",X"5A",X"00",X"66",X"9B",X"06",X"00",X"06",X"FF",X"00",X"00",X"00",X"B6",X"6F",X"00",
		X"00",X"BF",X"FB",X"00",X"00",X"FF",X"FB",X"00",X"00",X"BF",X"BB",X"00",X"00",X"BF",X"06",X"00",
		X"00",X"BF",X"06",X"00",X"00",X"99",X"BA",X"00",X"00",X"09",X"0A",X"00",X"00",X"6B",X"0A",X"00",
		X"00",X"6B",X"0A",X"00",X"00",X"60",X"0A",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"B0",X"00",
		X"B0",X"00",X"BB",X"00",X"B0",X"99",X"BB",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"09",X"9B",X"00",X"00",X"09",X"9B",X"00",X"BB",X"09",X"90",X"00",X"BB",X"99",X"90",X"00",
		X"00",X"55",X"90",X"00",X"00",X"0B",X"00",X"00",X"BB",X"BB",X"00",X"00",X"00",X"FF",X"FB",X"00",
		X"B0",X"FF",X"FB",X"00",X"00",X"BB",X"99",X"00",X"0F",X"FB",X"FF",X"B0",X"FF",X"FB",X"FF",X"B0",
		X"0B",X"FB",X"0B",X"00",X"0B",X"FB",X"5B",X"00",X"00",X"99",X"BB",X"00",X"00",X"B9",X"00",X"00",
		X"00",X"B9",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"99",X"00",X"AA",X"00",
		X"B9",X"99",X"A6",X"00",X"B9",X"99",X"A6",X"00",X"09",X"99",X"A6",X"00",X"09",X"09",X"90",X"00",
		X"9A",X"09",X"9B",X"00",X"9A",X"06",X"9B",X"00",X"99",X"06",X"A9",X"00",X"9B",X"A5",X"A9",X"00",
		X"90",X"55",X"A9",X"00",X"00",X"55",X"99",X"00",X"99",X"55",X"09",X"00",X"99",X"55",X"F9",X"00",
		X"B9",X"55",X"F6",X"00",X"99",X"A5",X"66",X"00",X"9A",X"AA",X"AA",X"B0",X"99",X"AA",X"AA",X"B0",
		X"0B",X"FA",X"AA",X"00",X"0B",X"FB",X"AA",X"00",X"0A",X"99",X"AA",X"00",X"0A",X"B9",X"A6",X"00",
		X"00",X"AA",X"66",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"09",X"99",X"00",X"04",X"11",X"19",X"00",X"44",X"19",X"B9",X"00",X"00",X"11",X"B9",X"00",
		X"99",X"BB",X"B9",X"00",X"99",X"BB",X"BB",X"00",X"99",X"BB",X"BB",X"00",X"99",X"BB",X"0B",X"00",
		X"90",X"BB",X"FB",X"90",X"90",X"BB",X"FB",X"40",X"10",X"BB",X"BB",X"40",X"15",X"0B",X"BB",X"90",
		X"10",X"00",X"F0",X"90",X"00",X"50",X"00",X"99",X"00",X"00",X"0F",X"99",X"00",X"04",X"0F",X"99",
		X"00",X"55",X"99",X"09",X"0B",X"95",X"99",X"09",X"BB",X"0B",X"5F",X"99",X"BB",X"FB",X"0F",X"99",
		X"FB",X"BB",X"0B",X"09",X"BB",X"BB",X"0B",X"99",X"BB",X"BB",X"BB",X"44",X"B9",X"00",X"BB",X"44",
		X"BB",X"00",X"BB",X"44",X"99",X"99",X"00",X"00",X"99",X"19",X"01",X"00",X"99",X"99",X"09",X"00",
		X"05",X"90",X"99",X"00",X"04",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"60",X"00",
		X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"66",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"60",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"F0",X"B0",X"00",X"00",X"90",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"B9",X"00",X"00",X"00",X"B9",X"00",X"00",
		X"00",X"B9",X"00",X"00",X"00",X"B9",X"00",X"00",X"00",X"B9",X"00",X"00",X"00",X"BC",X"00",X"00",
		X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"FF",X"00",X"99",X"00",X"9F",X"00",X"99",X"00",X"9F",X"00",
		X"99",X"00",X"9F",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"90",X"00",X"99",X"00",
		X"90",X"00",X"99",X"00",X"90",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"99",X"00",
		X"99",X"9F",X"99",X"00",X"99",X"FF",X"99",X"00",X"99",X"F9",X"99",X"00",X"99",X"FF",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"9F",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"B9",X"00",X"00",X"0F",X"B9",X"00",X"00",X"F9",X"B9",X"00",X"00",
		X"99",X"BB",X"00",X"00",X"99",X"BB",X"F0",X"00",X"99",X"00",X"9F",X"00",X"90",X"90",X"99",X"00",
		X"90",X"99",X"99",X"00",X"90",X"99",X"99",X"00",X"99",X"B9",X"99",X"00",X"99",X"0B",X"99",X"00",
		X"99",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"BB",X"00",X"BB",X"00",
		X"B0",X"00",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"F0",X"00",
		X"00",X"99",X"9F",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"F0",X"00",X"99",X"99",X"F0",
		X"00",X"99",X"99",X"F0",X"00",X"99",X"99",X"F0",X"00",X"99",X"99",X"F0",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"99",X"F0",X"00",X"99",X"99",X"F0",X"00",X"99",X"99",X"F0",
		X"00",X"99",X"99",X"F0",X"00",X"99",X"99",X"F0",X"00",X"99",X"99",X"00",X"00",X"99",X"9F",X"00",
		X"00",X"99",X"F0",X"00",X"00",X"99",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"55",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"96",X"00",X"00",X"99",X"96",X"99",X"00",
		X"55",X"55",X"96",X"00",X"55",X"55",X"96",X"00",X"55",X"55",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"55",X"55",X"99",X"80",X"55",X"55",X"96",X"99",X"55",X"55",X"96",X"99",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",
		X"00",X"0B",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"99",X"00",
		X"00",X"BB",X"B0",X"00",X"0F",X"9C",X"00",X"00",X"FF",X"BC",X"90",X"00",X"9F",X"FF",X"00",X"00",
		X"0F",X"FF",X"BB",X"00",X"09",X"BB",X"BB",X"00",X"00",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"9B",X"00",X"00",X"00",X"0B",X"09",X"00",X"00",X"99",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"F0",X"00",X"00",X"99",X"F0",X"00",X"00",X"99",X"F0",X"00",X"00",X"99",X"F0",X"00",
		X"00",X"99",X"F0",X"00",X"00",X"99",X"F0",X"00",X"00",X"99",X"F0",X"00",X"00",X"99",X"9F",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"B9",X"CC",X"00",X"00",X"0B",X"CC",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"0B",X"F0",X"00",X"00",X"00",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"F0",X"00",X"00",X"BB",X"FF",X"00",X"00",X"BB",X"BB",X"00",
		X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"F0",X"00",X"BB",X"00",X"F0",
		X"00",X"BB",X"00",X"F0",X"00",X"BB",X"00",X"F0",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"40",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"40",X"00",X"00",X"44",X"40",X"40",X"00",
		X"44",X"00",X"44",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"04",X"00",X"44",X"00",X"04",X"00",
		X"44",X"00",X"04",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"44",X"40",X"00",X"00",X"44",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"04",X"00",X"44",X"40",X"04",X"00",X"44",X"40",X"04",X"00",X"04",X"00",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"40",X"04",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"40",X"00",X"04",X"00",X"40",X"00",X"44",X"40",X"40",X"00",
		X"44",X"40",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"00",X"44",X"00",X"44",X"40",X"44",X"00",X"00",X"40",X"00",X"00",X"00",X"40",X"00",X"00",
		X"00",X"40",X"00",X"00",X"00",X"40",X"00",X"00",X"44",X"40",X"44",X"00",X"44",X"00",X"44",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"40",X"00",X"00",
		X"00",X"40",X"04",X"00",X"00",X"40",X"04",X"00",X"00",X"40",X"04",X"00",X"00",X"40",X"04",X"00",
		X"44",X"40",X"44",X"00",X"44",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"44",X"00",X"00",X"00",X"04",X"00",
		X"00",X"00",X"00",X"00",X"40",X"00",X"04",X"00",X"40",X"40",X"44",X"00",X"00",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"69",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"99",X"00",
		X"00",X"0F",X"99",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"96",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"FB",X"00",X"00",X"00",X"BB",X"FF",X"00",X"00",X"BB",X"FF",X"00",
		X"00",X"BB",X"FF",X"00",X"00",X"FB",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"FB",X"00",X"00",X"00",X"FB",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"F0",X"00",X"BB",X"00",X"F0",
		X"00",X"BB",X"00",X"F0",X"00",X"BB",X"BB",X"F0",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",
		X"00",X"BB",X"BB",X"00",X"00",X"BB",X"FF",X"00",X"00",X"BB",X"F0",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"66",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"66",X"00",X"00",X"0F",X"69",X"00",
		X"00",X"0F",X"60",X"00",X"00",X"0F",X"60",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"0F",X"F0",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"F0",X"00",X"00",X"0B",X"F0",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"0B",X"CC",X"00",X"00",X"B9",X"CC",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"9F",X"00",X"00",X"99",X"F0",X"00",X"00",X"99",X"F0",X"00",X"00",X"99",X"F0",X"00",
		X"00",X"99",X"F0",X"00",X"00",X"99",X"F0",X"00",X"00",X"99",X"F0",X"00",X"00",X"FF",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"F0",X"00",X"00",X"BB",X"FF",X"00",X"00",X"BB",X"BB",X"00",
		X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"F0",X"00",X"BB",X"00",X"F0",
		X"00",X"BB",X"00",X"F0",X"00",X"BB",X"00",X"F0",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"F0",X"00",X"BB",X"00",X"F0",
		X"00",X"BB",X"00",X"F0",X"00",X"BB",X"BB",X"F0",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",
		X"00",X"BB",X"BB",X"00",X"00",X"BB",X"FF",X"00",X"00",X"BB",X"F0",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"40",X"00",X"00",X"00",X"40",X"00",X"00",
		X"00",X"40",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"40",X"00",X"00",X"44",X"40",X"00",X"00",
		X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"40",X"00",X"00",
		X"44",X"40",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"04",X"40",X"00",X"00",
		X"04",X"40",X"00",X"00",X"04",X"40",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"40",X"00",X"00",
		X"40",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"00",X"00",X"00",X"44",X"00",X"44",X"00",X"04",X"00",X"44",X"00",X"00",X"40",X"00",X"00",
		X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"40",X"00",X"40",X"00",
		X"44",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"44",X"40",X"40",X"00",
		X"44",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"40",X"00",X"00",X"44",X"40",X"00",X"00",
		X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",
		X"44",X"40",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"40",X"00",X"00",
		X"00",X"40",X"00",X"00",X"44",X"40",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"FF",X"00",X"BB",X"00",X"BF",X"00",X"BB",X"00",X"BF",X"00",
		X"BB",X"00",X"BF",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"B0",X"00",X"BB",X"00",
		X"B0",X"00",X"BB",X"00",X"B0",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"00",
		X"BB",X"BF",X"BB",X"00",X"BB",X"FF",X"BB",X"00",X"BB",X"FB",X"BB",X"00",X"BB",X"FF",X"BB",X"00",
		X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",
		X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"BF",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"0F",X"11",X"00",X"00",X"F1",X"11",X"00",X"00",
		X"11",X"11",X"00",X"00",X"11",X"11",X"F0",X"00",X"11",X"BB",X"1F",X"00",X"11",X"BB",X"11",X"00",
		X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"FB",X"BB",X"00",X"BB",X"0F",X"BB",X"00",
		X"BB",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"BF",X"00",X"BF",X"00",
		X"F0",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"FF",X"00",X"BB",X"00",X"BF",X"00",X"BB",X"00",X"BF",X"00",
		X"BB",X"00",X"BF",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"B0",X"00",X"BB",X"00",
		X"B0",X"00",X"BB",X"00",X"B0",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"00",
		X"BB",X"BF",X"BB",X"00",X"BB",X"FF",X"BB",X"00",X"BB",X"FB",X"BB",X"00",X"BB",X"FF",X"BB",X"00",
		X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",
		X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"11",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"66",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"16",X"00",X"00",
		X"00",X"60",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"11",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"66",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"60",X"00",X"00",
		X"00",X"60",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"66",X"00",X"00",
		X"00",X"11",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"11",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"66",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"F0",X"00",X"00",X"11",X"BF",X"00",X"00",
		X"B1",X"BB",X"00",X"00",X"B1",X"BB",X"00",X"00",X"F1",X"BB",X"00",X"00",X"0F",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BF",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"BF",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"0F",X"BB",X"00",X"00",X"F1",X"BB",X"00",X"00",X"B1",X"BB",X"00",X"00",X"B1",X"BB",X"00",X"00",
		X"11",X"BF",X"00",X"00",X"11",X"F0",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",
		X"00",X"00",X"B1",X"F0",X"00",X"00",X"B1",X"F0",X"00",X"00",X"B1",X"00",X"00",X"00",X"11",X"00",
		X"00",X"0F",X"11",X"00",X"00",X"FB",X"11",X"00",X"00",X"BB",X"11",X"00",X"00",X"BB",X"11",X"00",
		X"00",X"BB",X"1F",X"00",X"00",X"BB",X"F0",X"00",X"00",X"FB",X"F0",X"00",X"00",X"FB",X"F0",X"00",
		X"00",X"0F",X"F0",X"00",X"00",X"0F",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",X"0F",X"F0",X"00",X"00",X"0F",X"F0",X"00",
		X"00",X"FB",X"F0",X"00",X"00",X"FB",X"F0",X"00",X"00",X"BB",X"F0",X"00",X"00",X"BB",X"1F",X"00",
		X"00",X"BB",X"11",X"00",X"00",X"BB",X"11",X"00",X"00",X"FB",X"11",X"00",X"00",X"0F",X"11",X"00",
		X"00",X"00",X"11",X"00",X"00",X"00",X"B1",X"00",X"00",X"00",X"B1",X"F0",X"00",X"00",X"B1",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"0F",X"BB",X"00",X"00",X"FB",X"BB",X"00",X"00",
		X"FB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"B0",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BF",X"00",X"00",X"00",X"BF",X"00",X"00",
		X"00",X"BF",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BF",X"00",X"00",X"00",X"BF",X"00",X"00",X"00",X"BF",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"B0",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"FB",X"BB",X"00",X"00",
		X"FB",X"BB",X"00",X"00",X"0F",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"06",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"06",X"00",
		X"00",X"06",X"06",X"00",X"00",X"06",X"06",X"00",X"00",X"06",X"06",X"00",X"00",X"00",X"66",X"00",
		X"66",X"00",X"6B",X"00",X"66",X"00",X"60",X"00",X"66",X"66",X"6B",X"00",X"66",X"66",X"66",X"00",
		X"66",X"66",X"6B",X"00",X"66",X"00",X"60",X"00",X"66",X"00",X"6B",X"00",X"00",X"00",X"66",X"00",
		X"00",X"06",X"06",X"00",X"00",X"06",X"06",X"00",X"00",X"06",X"06",X"00",X"00",X"00",X"06",X"00",
		X"00",X"00",X"06",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"0F",X"BB",X"00",X"00",X"FB",X"BB",X"00",X"00",
		X"FB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"B0",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BF",X"00",X"00",X"00",X"BF",X"00",X"00",
		X"00",X"BF",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BF",X"00",X"00",X"00",X"BF",X"00",X"00",X"00",X"BF",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"B0",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"FB",X"BB",X"00",X"00",
		X"FB",X"BB",X"00",X"00",X"0F",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"04",X"00",X"44",X"00",X"44",X"40",X"00",X"00",
		X"44",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"04",X"00",X"44",X"00",X"04",X"00",X"44",X"00",X"04",X"00",X"00",X"40",X"04",X"00",
		X"00",X"40",X"44",X"00",X"04",X"40",X"44",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",
		X"40",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"44",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"40",X"44",X"00",X"00",X"40",X"44",X"00",
		X"00",X"40",X"04",X"00",X"00",X"40",X"04",X"00",X"00",X"40",X"04",X"00",X"44",X"40",X"04",X"00",
		X"44",X"40",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",
		X"44",X"40",X"00",X"00",X"44",X"40",X"04",X"00",X"00",X"40",X"04",X"00",X"00",X"00",X"04",X"00",
		X"00",X"00",X"04",X"00",X"44",X"40",X"00",X"00",X"44",X"40",X"00",X"00",X"04",X"00",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"BB",X"BB",X"B0",X"00",X"BB",X"BB",X"BB",X"BB",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"00",
		X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"B0",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"50",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"50",X"00",X"00",X"00",X"00",X"00",X"00",
		X"50",X"50",X"05",X"00",X"00",X"00",X"00",X"00",X"50",X"50",X"0B",X"50",X"00",X"00",X"BB",X"00",
		X"50",X"0C",X"BF",X"55",X"00",X"00",X"10",X"00",X"00",X"CC",X"11",X"50",X"00",X"00",X"11",X"00",
		X"00",X"CC",X"15",X"50",X"00",X"00",X"00",X"00",X"00",X"CC",X"11",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"01",X"05",X"00",X"00",X"01",X"00",X"00",X"00",X"11",X"05",X"00",X"00",X"1F",X"00",
		X"05",X"10",X"BB",X"00",X"00",X"00",X"0B",X"00",X"05",X"05",X"50",X"00",X"00",X"00",X"00",X"00",
		X"05",X"05",X"50",X"00",X"00",X"00",X"00",X"00",X"05",X"05",X"00",X"00",X"00",X"00",X"00",X"00",
		X"05",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"04",X"00",X"00",X"00",
		X"00",X"00",X"04",X"00",X"00",X"40",X"04",X"00",X"00",X"40",X"44",X"00",X"00",X"00",X"44",X"00",
		X"04",X"00",X"44",X"00",X"44",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"40",X"00",
		X"00",X"40",X"44",X"00",X"00",X"40",X"04",X"00",X"04",X"00",X"04",X"00",X"44",X"00",X"04",X"00",
		X"40",X"00",X"04",X"00",X"44",X"00",X"44",X"00",X"04",X"00",X"44",X"00",X"00",X"40",X"00",X"00",
		X"00",X"40",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"04",X"00",
		X"00",X"00",X"44",X"00",X"00",X"40",X"40",X"00",X"00",X"40",X"40",X"00",X"00",X"00",X"40",X"00",
		X"00",X"00",X"40",X"00",X"44",X"00",X"40",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"BB",X"BB",X"BB",X"0B",
		X"BB",X"BB",X"BB",X"B0",X"F0",X"0F",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"F0",X"00",X"00",X"F0",X"0F",X"00",X"00",X"BB",X"BB",X"BB",X"B0",X"BB",X"BB",X"BB",X"0B",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"B9",X"00",X"00",X"00",X"B9",X"00",X"00",
		X"00",X"B9",X"00",X"00",X"00",X"B9",X"00",X"00",X"00",X"B9",X"00",X"00",X"00",X"BC",X"00",X"00",
		X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"60",X"00",X"00",X"F0",X"66",X"00",X"00",X"6F",X"66",X"00",X"00",X"BF",X"66",X"00",
		X"06",X"0F",X"B6",X"00",X"06",X"00",X"F6",X"00",X"06",X"66",X"66",X"00",X"00",X"0B",X"06",X"00",
		X"06",X"B0",X"66",X"00",X"06",X"B0",X"66",X"00",X"06",X"B0",X"66",X"00",X"06",X"B0",X"66",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"60",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"60",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",
		X"00",X"00",X"60",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"60",X"00",
		X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"66",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"60",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"0C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0C",X"00",X"00",X"CC",X"CC",X"00",X"00",
		X"CC",X"CC",X"00",X"00",X"C7",X"55",X"00",X"00",X"C7",X"55",X"00",X"00",X"07",X"55",X"CC",X"00",
		X"0C",X"55",X"CC",X"00",X"0C",X"55",X"5C",X"00",X"0C",X"55",X"55",X"00",X"00",X"5B",X"55",X"00",
		X"00",X"BB",X"55",X"00",X"0C",X"5B",X"55",X"00",X"0C",X"55",X"55",X"00",X"0C",X"55",X"00",X"00",
		X"07",X"55",X"0C",X"00",X"C7",X"55",X"CC",X"00",X"C7",X"55",X"CC",X"00",X"CC",X"55",X"00",X"00",
		X"CC",X"CC",X"00",X"00",X"0C",X"CC",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"F0",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"0F",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"55",X"02",X"00",X"02",X"55",X"02",X"00",
		X"22",X"00",X"02",X"00",X"22",X"55",X"2C",X"00",X"00",X"55",X"22",X"00",X"00",X"55",X"22",X"00",
		X"00",X"55",X"52",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"5F",X"55",X"00",
		X"55",X"FA",X"55",X"50",X"02",X"AF",X"55",X"02",X"22",X"FF",X"55",X"22",X"22",X"FA",X"55",X"22",
		X"22",X"F5",X"55",X"22",X"22",X"FA",X"00",X"22",X"22",X"FF",X"55",X"22",X"02",X"AF",X"55",X"02",
		X"55",X"FA",X"55",X"50",X"55",X"5F",X"00",X"00",X"55",X"55",X"05",X"00",X"50",X"55",X"05",X"00",
		X"50",X"55",X"52",X"00",X"00",X"00",X"22",X"00",X"00",X"55",X"22",X"00",X"22",X"55",X"2C",X"00",
		X"22",X"55",X"02",X"00",X"02",X"55",X"02",X"00",X"00",X"55",X"02",X"00",X"00",X"00",X"02",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"66",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"11",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"66",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"66",X"00",X"00",
		X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"11",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"66",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"06",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"06",X"00",X"00",X"06",X"06",X"00",
		X"00",X"06",X"06",X"00",X"00",X"06",X"06",X"00",X"00",X"06",X"06",X"00",X"00",X"00",X"66",X"00",
		X"00",X"00",X"6B",X"00",X"00",X"00",X"60",X"00",X"00",X"66",X"6B",X"00",X"00",X"66",X"66",X"00",
		X"00",X"66",X"6B",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"6B",X"00",X"00",X"00",X"66",X"00",
		X"00",X"06",X"06",X"00",X"00",X"06",X"06",X"00",X"00",X"06",X"06",X"00",X"00",X"06",X"06",X"00",
		X"00",X"06",X"06",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"6F",X"66",X"00",X"06",X"BF",X"66",X"00",
		X"06",X"0F",X"B6",X"00",X"06",X"00",X"F6",X"00",X"06",X"66",X"66",X"00",X"00",X"0B",X"06",X"00",
		X"06",X"B0",X"66",X"00",X"06",X"B0",X"66",X"00",X"06",X"B0",X"66",X"00",X"06",X"B0",X"66",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"44",X"D0",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"F0",X"00",X"00",X"00",X"CD",X"0F",X"00",
		X"00",X"04",X"F0",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"B0",X"09",X"00",
		X"00",X"BB",X"09",X"00",X"00",X"BB",X"09",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"BB",X"09",X"00",X"00",X"BB",X"09",X"00",
		X"00",X"B0",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"05",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"05",X"00",X"00",X"00",X"00",X"00",
		X"50",X"11",X"05",X"00",X"B0",X"11",X"00",X"00",X"5B",X"11",X"05",X"00",X"00",X"11",X"00",X"00",
		X"55",X"C1",X"00",X"00",X"00",X"01",X"00",X"00",X"C5",X"C1",X"00",X"00",X"01",X"11",X"00",X"00",
		X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"00",X"00",X"00",
		X"11",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"B5",X"05",X"50",X"00",X"00",X"00",X"00",X"00",
		X"05",X"00",X"50",X"00",X"B0",X"00",X"00",X"00",X"B0",X"50",X"50",X"00",X"00",X"00",X"00",X"00",
		X"00",X"50",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
