library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_8E is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_8E is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"70",X"38",X"3C",X"7C",X"F0",X"00",X"00",X"00",X"40",X"E0",X"FC",X"7E",X"3E",
		X"F8",X"F0",X"7C",X"3C",X"38",X"70",X"00",X"00",X"7C",X"3E",X"7E",X"FC",X"E0",X"40",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"82",X"C6",X"7C",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"7C",X"C6",X"82",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"38",X"7C",X"C2",X"82",X"86",X"7C",X"38",X"00",X"00",X"02",X"02",X"FE",X"FE",X"42",X"02",X"00",
		X"62",X"F2",X"BA",X"9A",X"9E",X"CE",X"46",X"00",X"8C",X"DE",X"F2",X"B2",X"92",X"86",X"04",X"00",
		X"08",X"FE",X"FE",X"C8",X"68",X"38",X"18",X"00",X"9C",X"BE",X"A2",X"A2",X"A2",X"E6",X"E4",X"00",
		X"0C",X"9E",X"92",X"92",X"D2",X"7E",X"3C",X"00",X"C0",X"E0",X"B0",X"9E",X"8E",X"C0",X"C0",X"00",
		X"6C",X"FE",X"92",X"92",X"92",X"FE",X"6C",X"00",X"78",X"FC",X"96",X"92",X"92",X"F2",X"60",X"00",
		X"7C",X"82",X"AA",X"AA",X"BA",X"82",X"7C",X"00",X"7C",X"82",X"BA",X"AA",X"BE",X"82",X"7C",X"00",
		X"2E",X"2E",X"3A",X"3A",X"00",X"20",X"7E",X"7E",X"00",X"00",X"00",X"E0",X"C0",X"00",X"00",X"00",
		X"20",X"00",X"70",X"50",X"50",X"7E",X"7E",X"00",X"00",X"00",X"00",X"F0",X"FA",X"FA",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"7E",X"C8",X"88",X"C8",X"7E",X"3E",X"00",
		X"6C",X"FE",X"92",X"92",X"92",X"FE",X"FE",X"00",X"44",X"C6",X"82",X"82",X"C6",X"7C",X"38",X"00",
		X"38",X"7C",X"C6",X"82",X"82",X"FE",X"FE",X"00",X"00",X"82",X"92",X"92",X"92",X"FE",X"FE",X"00",
		X"80",X"90",X"90",X"90",X"90",X"FE",X"FE",X"00",X"9E",X"9E",X"92",X"82",X"C6",X"7C",X"38",X"00",
		X"FE",X"FE",X"10",X"10",X"10",X"FE",X"FE",X"00",X"00",X"82",X"82",X"FE",X"FE",X"82",X"82",X"00",
		X"FC",X"FE",X"02",X"02",X"02",X"06",X"04",X"00",X"82",X"C6",X"6E",X"3C",X"18",X"FE",X"FE",X"00",
		X"00",X"02",X"02",X"02",X"02",X"FE",X"FE",X"00",X"FE",X"FE",X"70",X"38",X"70",X"FE",X"FE",X"00",
		X"FE",X"FE",X"1C",X"38",X"70",X"FE",X"FE",X"00",X"7C",X"FE",X"82",X"82",X"82",X"FE",X"7C",X"00",
		X"70",X"88",X"88",X"88",X"88",X"FE",X"FE",X"00",X"7A",X"FC",X"8E",X"8A",X"82",X"FE",X"7C",X"00",
		X"72",X"F6",X"9E",X"8C",X"88",X"FE",X"FE",X"00",X"4C",X"DE",X"92",X"92",X"92",X"F6",X"64",X"00",
		X"00",X"80",X"80",X"FE",X"FE",X"80",X"80",X"00",X"FC",X"FE",X"02",X"02",X"02",X"FE",X"FC",X"00",
		X"F0",X"F8",X"1C",X"0E",X"1C",X"F8",X"F0",X"00",X"FC",X"FE",X"1C",X"38",X"1C",X"FE",X"FC",X"00",
		X"C6",X"EE",X"7C",X"38",X"7C",X"EE",X"C6",X"00",X"00",X"C0",X"F0",X"1E",X"1E",X"F0",X"C0",X"00",
		X"C2",X"E2",X"F2",X"BA",X"9E",X"8E",X"86",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"FF",
		X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"78",X"78",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"7F",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FE",
		X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F8",X"F8",X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"80",X"C0",X"E0",X"FF",X"FF",X"FB",X"F9",X"F8",
		X"78",X"38",X"18",X"F8",X"F8",X"FC",X"FE",X"FF",X"00",X"00",X"00",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"F8",X"78",X"38",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FB",X"F9",X"F8",
		X"F8",X"F8",X"F8",X"FF",X"FF",X"FF",X"FB",X"F9",X"78",X"38",X"18",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"78",X"78",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"7F",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FE",
		X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F8",X"F8",X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"80",X"C0",X"E0",X"FF",X"FF",X"FB",X"F9",X"F8",
		X"78",X"38",X"18",X"F8",X"F8",X"FC",X"FE",X"FF",X"00",X"00",X"00",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"F8",X"78",X"38",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FB",X"F9",X"F8",
		X"F8",X"F8",X"F8",X"FF",X"FF",X"FF",X"FB",X"F9",X"78",X"38",X"18",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"E0",X"20",X"18",
		X"08",X"04",X"03",X"00",X"00",X"00",X"00",X"00",X"18",X"00",X"C0",X"20",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",X"E0",
		X"07",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"07",X"0F",X"1C",X"38",X"38",X"00",X"00",X"C0",X"E0",X"F0",X"38",X"1C",X"1C",
		X"38",X"38",X"1C",X"0F",X"07",X"03",X"00",X"00",X"1C",X"1C",X"38",X"F0",X"E0",X"C0",X"00",X"00",
		X"07",X"0F",X"1F",X"38",X"70",X"E0",X"E0",X"E0",X"E0",X"F0",X"F8",X"1C",X"0E",X"07",X"07",X"07",
		X"E0",X"E0",X"E0",X"70",X"38",X"1F",X"0F",X"07",X"07",X"07",X"07",X"0E",X"1C",X"F8",X"F0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"1F",X"00",X"00",X"00",X"00",X"00",X"FE",X"FF",X"FF",
		X"1F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FE",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"03",X"00",X"00",X"30",X"1C",X"06",X"C2",X"F1",X"F9",
		X"07",X"05",X"03",X"03",X"01",X"00",X"00",X"00",X"FC",X"FC",X"FE",X"FE",X"FC",X"70",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"1F",X"00",X"00",X"30",X"1C",X"06",X"C2",X"F1",X"F9",
		X"1F",X"07",X"03",X"03",X"01",X"00",X"00",X"00",X"FC",X"FC",X"FE",X"FE",X"FC",X"70",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"78",X"78",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"7F",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FE",
		X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F8",X"F8",X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"80",X"C0",X"E0",X"FF",X"FF",X"FB",X"F9",X"F8",
		X"78",X"38",X"18",X"F8",X"F8",X"FC",X"FE",X"FF",X"00",X"00",X"00",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"F8",X"78",X"38",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FB",X"F9",X"F8",
		X"F8",X"F8",X"F8",X"FF",X"FF",X"FF",X"FB",X"F9",X"78",X"38",X"18",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"78",X"78",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"7F",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FE",
		X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F8",X"F8",X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"80",X"C0",X"E0",X"FF",X"FF",X"FB",X"F9",X"F8",
		X"78",X"38",X"18",X"F8",X"F8",X"FC",X"FE",X"FF",X"00",X"00",X"00",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"F8",X"78",X"38",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FB",X"F9",X"F8",
		X"F8",X"F8",X"F8",X"FF",X"FF",X"FF",X"FB",X"F9",X"78",X"38",X"18",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"C0",X"C0",X"C0",X"C0",X"FF",X"FF",X"FF",X"FF",X"03",X"03",X"03",X"03",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"C0",X"C0",X"C0",X"C0",X"FF",X"FF",X"FF",X"FF",X"03",X"03",X"03",X"03",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"FF",X"FF",X"FF",X"FF",X"C0",X"C0",X"C0",X"C0",X"FF",X"FF",X"FF",X"FF",X"03",X"03",X"03",X"03",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"FF",X"FF",X"FF",X"FF",X"C0",X"C0",X"C0",X"C0",X"FF",X"FF",X"FF",X"FF",X"03",X"03",X"03",X"03",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"FF",X"FF",X"FF",X"FF",X"C0",X"C0",X"C0",X"C0",X"FF",X"FF",X"FF",X"FF",X"03",X"03",X"03",X"03",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"FF",X"FF",X"FF",X"FF",X"C0",X"C0",X"C0",X"C0",X"FF",X"FF",X"FF",X"FF",X"03",X"03",X"03",X"03",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"0F",X"07",X"03",X"00",X"00",X"00",X"00",X"1E",X"1E",X"1E",X"1E",X"1E",X"1E",X"1E",X"1E",
		X"00",X"00",X"00",X"03",X"07",X"0F",X"1F",X"1E",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"F0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"80",X"C0",X"E0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"40",X"60",X"20",X"30",X"18",X"0C",
		X"18",X"30",X"30",X"60",X"60",X"C0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"06",X"06",X"06",X"04",X"04",X"00",X"18",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"00",X"FA",X"FA",X"F2",X"E4",X"CC",X"18",X"E0",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",
		X"C0",X"E0",X"F1",X"F3",X"E7",X"0F",X"7F",X"FF",X"7A",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",
		X"20",X"BC",X"BF",X"BF",X"1F",X"07",X"01",X"C0",X"02",X"02",X"82",X"E2",X"E2",X"E2",X"E2",X"62",
		X"F0",X"F8",X"FE",X"7F",X"1F",X"0F",X"07",X"83",X"02",X"02",X"02",X"02",X"CA",X"8A",X"9A",X"3A",
		X"1F",X"07",X"00",X"00",X"80",X"00",X"70",X"F8",X"8A",X"0A",X"0A",X"3A",X"3A",X"7A",X"3A",X"1A",
		X"FC",X"00",X"00",X"00",X"FF",X"FF",X"7F",X"00",X"0A",X"0A",X"02",X"02",X"82",X"C2",X"C2",X"02",
		X"80",X"00",X"00",X"00",X"00",X"08",X"18",X"38",X"3A",X"3A",X"FA",X"FA",X"FA",X"3A",X"0A",X"0A",
		X"7E",X"78",X"60",X"40",X"00",X"01",X"07",X"1F",X"0A",X"0A",X"0A",X"0A",X"0A",X"8A",X"8A",X"8A",
		X"03",X"07",X"07",X"0F",X"0F",X"1F",X"1F",X"3E",X"C2",X"C2",X"C2",X"CA",X"8A",X"8A",X"0A",X"0A",
		X"38",X"62",X"0C",X"F8",X"F0",X"F0",X"E0",X"C0",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",
		X"F0",X"F0",X"F0",X"E0",X"E0",X"E0",X"C0",X"40",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"00",X"00",X"80",X"00",X"00",X"00",X"01",X"03",X"1A",X"0A",X"0A",X"02",X"82",X"82",X"C2",X"C2",
		X"C0",X"8B",X"1B",X"7B",X"FF",X"FF",X"FF",X"FF",X"02",X"C2",X"C2",X"C2",X"82",X"82",X"82",X"1A",
		X"FF",X"FC",X"F1",X"C7",X"1F",X"01",X"00",X"00",X"1A",X"7A",X"FA",X"FA",X"FA",X"FA",X"1A",X"02",
		X"00",X"FF",X"00",X"FF",X"FF",X"F8",X"FC",X"FE",X"00",X"E0",X"18",X"CC",X"E4",X"12",X"FA",X"7A",
		X"FF",X"FE",X"FC",X"F8",X"FF",X"FA",X"F8",X"F1",X"3A",X"7A",X"FA",X"02",X"02",X"02",X"42",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"78",X"78",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"7F",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FE",
		X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F8",X"F8",X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"80",X"C0",X"E0",X"FF",X"FF",X"FB",X"F9",X"F8",
		X"78",X"38",X"18",X"F8",X"F8",X"FC",X"FE",X"FF",X"00",X"00",X"00",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"F8",X"78",X"38",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FB",X"F9",X"F8",
		X"F8",X"F8",X"F8",X"FF",X"FF",X"FF",X"FB",X"F9",X"78",X"38",X"18",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"78",X"78",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"7F",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FE",
		X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F8",X"F8",X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"80",X"C0",X"E0",X"FF",X"FF",X"FB",X"F9",X"F8",
		X"78",X"38",X"18",X"F8",X"F8",X"FC",X"FE",X"FF",X"00",X"00",X"00",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"F8",X"78",X"38",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FB",X"F9",X"F8",
		X"F8",X"F8",X"F8",X"FF",X"FF",X"FF",X"FB",X"F9",X"78",X"38",X"18",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"00",X"00",X"03",X"07",X"07",X"07",X"03",X"07",X"00",X"00",X"E0",X"E0",X"E0",X"C0",X"E0",X"E0",
		X"07",X"07",X"03",X"07",X"07",X"05",X"00",X"00",X"E0",X"C0",X"A0",X"E0",X"E0",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"07",X"0F",X"0F",X"00",X"00",X"00",X"00",X"C0",X"E0",X"F0",X"F0",
		X"0F",X"0F",X"07",X"03",X"00",X"00",X"00",X"00",X"F0",X"F0",X"E0",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"07",X"0F",X"1C",X"38",X"38",X"00",X"00",X"C0",X"E0",X"F0",X"38",X"1C",X"1C",
		X"38",X"38",X"1C",X"0F",X"07",X"03",X"00",X"00",X"1C",X"1C",X"38",X"F0",X"E0",X"C0",X"00",X"00",
		X"07",X"0F",X"1F",X"38",X"70",X"E0",X"E0",X"E0",X"E0",X"F0",X"F8",X"1C",X"0E",X"07",X"07",X"07",
		X"E0",X"E0",X"E0",X"70",X"38",X"1F",X"0F",X"07",X"07",X"07",X"07",X"0E",X"1C",X"F8",X"F0",X"E0",
		X"00",X"00",X"1F",X"3F",X"3F",X"3E",X"1F",X"3F",X"00",X"00",X"00",X"3A",X"7E",X"7E",X"5C",X"00",
		X"3F",X"3E",X"1D",X"3F",X"3F",X"2E",X"00",X"00",X"0A",X"14",X"0A",X"14",X"00",X"00",X"00",X"00",
		X"00",X"00",X"1F",X"3F",X"3F",X"3E",X"1F",X"3F",X"00",X"00",X"00",X"3E",X"7E",X"7E",X"54",X"00",
		X"3F",X"3E",X"1D",X"3F",X"3F",X"2E",X"00",X"00",X"0A",X"14",X"0A",X"14",X"00",X"00",X"00",X"00",
		X"00",X"00",X"1F",X"3F",X"3F",X"3E",X"1F",X"3F",X"00",X"00",X"00",X"3E",X"7C",X"38",X"70",X"00",
		X"3F",X"3E",X"1D",X"3F",X"3F",X"2E",X"00",X"00",X"0A",X"14",X"0A",X"14",X"00",X"00",X"00",X"00",
		X"00",X"00",X"1F",X"3F",X"3F",X"3E",X"1F",X"3F",X"00",X"00",X"00",X"2E",X"7E",X"7E",X"74",X"00",
		X"3F",X"3E",X"1D",X"3F",X"3F",X"2E",X"00",X"00",X"0A",X"14",X"0A",X"14",X"00",X"00",X"00",X"00",
		X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FE",X"FF",X"80",X"C0",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"FF",X"81",X"85",X"9F",X"85",X"FD",X"81",X"FF",X"FF",X"81",X"DF",X"D3",X"D3",X"F3",X"81",X"FF",
		X"FF",X"81",X"DF",X"D3",X"D3",X"FF",X"81",X"FF",X"FF",X"81",X"FF",X"C1",X"C1",X"C1",X"81",X"FF",
		X"FF",X"81",X"FF",X"D3",X"D3",X"FF",X"81",X"FF",X"FF",X"81",X"FF",X"D3",X"D3",X"F3",X"81",X"FF",
		X"FF",X"81",X"FF",X"D1",X"D1",X"FF",X"81",X"FF",X"FF",X"81",X"9F",X"93",X"93",X"FF",X"81",X"FF",
		X"FF",X"81",X"E7",X"C3",X"C3",X"FF",X"81",X"FF",X"FF",X"81",X"FF",X"93",X"93",X"9F",X"81",X"FF",
		X"FF",X"81",X"C3",X"D3",X"D3",X"FF",X"81",X"FF",X"FF",X"81",X"C1",X"D1",X"D1",X"FF",X"81",X"FF",
		X"00",X"00",X"7E",X"42",X"42",X"7E",X"00",X"00",X"00",X"00",X"02",X"7E",X"22",X"00",X"00",X"00",
		X"00",X"00",X"7A",X"4A",X"4A",X"6E",X"00",X"00",X"00",X"00",X"7E",X"52",X"42",X"66",X"00",X"00",
		X"00",X"00",X"04",X"1E",X"04",X"7C",X"00",X"00",X"00",X"00",X"5E",X"52",X"52",X"72",X"00",X"00",
		X"00",X"00",X"5E",X"52",X"52",X"7E",X"00",X"00",X"00",X"00",X"7E",X"40",X"40",X"40",X"00",X"00",
		X"00",X"00",X"7E",X"52",X"52",X"7E",X"00",X"00",X"00",X"00",X"7E",X"52",X"52",X"72",X"00",X"00",
		X"00",X"00",X"7E",X"50",X"50",X"7E",X"00",X"00",X"00",X"00",X"1E",X"12",X"12",X"7E",X"00",X"00",
		X"00",X"00",X"66",X"42",X"42",X"7E",X"00",X"00",X"00",X"00",X"7E",X"12",X"12",X"1E",X"00",X"00",
		X"00",X"00",X"42",X"52",X"52",X"7E",X"00",X"00",X"00",X"00",X"40",X"50",X"50",X"7E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"1F",X"7F",X"00",X"00",X"00",X"00",X"00",X"FE",X"FF",X"FF",
		X"7F",X"1F",X"0F",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FE",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"07",X"00",X"00",X"00",X"60",X"18",X"8C",X"C4",X"F2",
		X"07",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"FA",X"FC",X"FC",X"F8",X"60",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"07",X"00",X"00",X"30",X"1C",X"06",X"C2",X"F1",X"F9",
		X"07",X"07",X"03",X"03",X"01",X"00",X"00",X"00",X"FC",X"FC",X"FE",X"FE",X"FC",X"70",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"03",X"00",X"00",X"30",X"1C",X"06",X"C2",X"F1",X"F9",
		X"07",X"07",X"03",X"03",X"01",X"00",X"00",X"00",X"FC",X"FC",X"FE",X"FE",X"FC",X"70",X"00",X"00",
		X"00",X"00",X"00",X"07",X"07",X"0F",X"3F",X"4F",X"00",X"00",X"00",X"AC",X"AC",X"AE",X"AE",X"AE",
		X"87",X"87",X"80",X"47",X"38",X"00",X"00",X"00",X"AC",X"AC",X"00",X"00",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"21",X"13",X"00",X"00",X"00",X"30",X"FC",X"FE",X"FE",X"FF",
		X"0F",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FE",X"FE",X"FC",X"30",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"21",X"13",X"00",X"00",X"00",X"30",X"FC",X"FE",X"FE",X"FF",
		X"0F",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FE",X"FE",X"FC",X"30",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"21",X"13",X"00",X"00",X"00",X"30",X"FC",X"FE",X"FE",X"FF",
		X"0F",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FE",X"FE",X"FC",X"30",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
