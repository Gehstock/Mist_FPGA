library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_PGM is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_PGM is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"AF",X"32",X"01",X"68",X"C3",X"71",X"00",X"FF",X"77",X"3C",X"23",X"77",X"3C",X"19",X"C9",X"FF",
		X"77",X"23",X"10",X"FC",X"C9",X"FF",X"FF",X"FF",X"77",X"23",X"10",X"FC",X"0D",X"20",X"F9",X"C9",
		X"85",X"6F",X"3E",X"00",X"8C",X"67",X"7E",X"C9",X"87",X"E1",X"5F",X"16",X"00",X"19",X"5E",X"23",
		X"56",X"EB",X"E9",X"FF",X"FF",X"FF",X"FF",X"FF",X"E5",X"26",X"40",X"3A",X"A0",X"40",X"6F",X"CB",
		X"7E",X"28",X"0E",X"72",X"2C",X"73",X"2C",X"7D",X"FE",X"C0",X"30",X"02",X"3E",X"C0",X"32",X"A0",
		X"40",X"E1",X"C9",X"0F",X"11",X"22",X"04",X"31",X"06",X"15",X"02",X"33",X"07",X"21",X"03",X"24",
		X"05",X"13",X"01",X"FF",X"FF",X"FF",X"C3",X"A3",X"04",X"80",X"40",X"20",X"10",X"08",X"04",X"02",
		X"01",X"21",X"00",X"40",X"11",X"01",X"40",X"01",X"00",X"08",X"36",X"00",X"ED",X"B0",X"3E",X"9B",
		X"32",X"03",X"81",X"3E",X"89",X"32",X"03",X"82",X"3E",X"08",X"32",X"42",X"42",X"32",X"01",X"82",
		X"C3",X"F6",X"3F",X"21",X"C0",X"40",X"06",X"40",X"3E",X"FF",X"D7",X"21",X"43",X"42",X"06",X"1C",
		X"D7",X"21",X"43",X"43",X"22",X"40",X"42",X"3A",X"00",X"70",X"AF",X"32",X"01",X"68",X"32",X"07",
		X"68",X"32",X"06",X"68",X"21",X"C0",X"C0",X"22",X"A0",X"40",X"21",X"00",X"48",X"CD",X"1C",X"0D",
		X"3E",X"10",X"32",X"17",X"40",X"3A",X"02",X"81",X"2F",X"0F",X"47",X"E6",X"02",X"32",X"00",X"40",
		X"78",X"0F",X"0F",X"E6",X"01",X"32",X"0F",X"40",X"3A",X"01",X"81",X"2F",X"E6",X"03",X"FE",X"03",
		X"28",X"07",X"C6",X"03",X"32",X"07",X"40",X"18",X"05",X"3E",X"FF",X"32",X"07",X"40",X"CD",X"B1",
		X"3F",X"47",X"E6",X"F0",X"0F",X"0F",X"0F",X"0F",X"21",X"53",X"00",X"85",X"6F",X"7E",X"32",X"0F",
		X"41",X"78",X"E6",X"0F",X"21",X"53",X"00",X"85",X"6F",X"7E",X"32",X"0C",X"41",X"CD",X"97",X"0A",
		X"AF",X"3D",X"20",X"FD",X"CD",X"A6",X"0A",X"21",X"00",X"50",X"01",X"00",X"01",X"16",X"00",X"72",
		X"23",X"0B",X"78",X"B1",X"20",X"F9",X"16",X"3F",X"21",X"00",X"48",X"01",X"00",X"08",X"72",X"3A",
		X"00",X"70",X"23",X"0B",X"78",X"B1",X"20",X"F6",X"CD",X"72",X"01",X"00",X"00",X"CD",X"72",X"01",
		X"00",X"00",X"CD",X"F1",X"0A",X"3E",X"01",X"32",X"01",X"68",X"21",X"00",X"42",X"06",X"0A",X"36",
		X"00",X"2C",X"36",X"00",X"2C",X"36",X"01",X"2C",X"10",X"F5",X"21",X"AA",X"40",X"36",X"01",X"21",
		X"C0",X"41",X"3E",X"0F",X"06",X"1E",X"D7",X"CD",X"93",X"3F",X"C3",X"81",X"01",X"3A",X"00",X"70",
		X"18",X"FB",X"0B",X"3A",X"00",X"70",X"3A",X"01",X"81",X"07",X"D0",X"78",X"B1",X"20",X"F3",X"37",
		X"C9",X"26",X"40",X"3A",X"A1",X"40",X"6F",X"7E",X"87",X"30",X"08",X"CD",X"85",X"36",X"CD",X"C9",
		X"01",X"18",X"EE",X"E6",X"1F",X"4F",X"06",X"00",X"36",X"FF",X"23",X"5E",X"36",X"FF",X"2C",X"7D",
		X"FE",X"C0",X"30",X"02",X"3E",X"C0",X"32",X"A1",X"40",X"7B",X"21",X"B7",X"01",X"09",X"5E",X"23",
		X"56",X"21",X"81",X"01",X"E5",X"EB",X"E9",X"2B",X"02",X"52",X"02",X"79",X"02",X"F9",X"02",X"B2",
		X"03",X"CB",X"03",X"12",X"04",X"41",X"04",X"7F",X"04",X"3A",X"80",X"41",X"47",X"E6",X"0F",X"CA",
		X"D3",X"01",X"C9",X"3A",X"06",X"40",X"A7",X"C8",X"11",X"E0",X"FF",X"21",X"E0",X"48",X"3A",X"0E",
		X"40",X"A7",X"28",X"22",X"36",X"02",X"CD",X"1C",X"02",X"21",X"40",X"4B",X"CD",X"1A",X"02",X"3A",
		X"BD",X"40",X"A7",X"21",X"40",X"4B",X"28",X"03",X"21",X"E0",X"48",X"CB",X"60",X"C8",X"3A",X"06",
		X"40",X"0F",X"D0",X"C3",X"23",X"02",X"21",X"E0",X"48",X"CD",X"23",X"02",X"21",X"21",X"49",X"CD",
		X"23",X"02",X"CD",X"23",X"02",X"CD",X"23",X"02",X"18",X"CF",X"36",X"01",X"19",X"36",X"25",X"19",
		X"36",X"20",X"C9",X"3E",X"10",X"77",X"19",X"77",X"19",X"77",X"C9",X"3A",X"06",X"40",X"A7",X"C8",
		X"21",X"82",X"48",X"11",X"20",X"00",X"3A",X"80",X"42",X"3C",X"FE",X"10",X"38",X"02",X"3E",X"10",
		X"4F",X"47",X"36",X"0C",X"19",X"10",X"FB",X"3E",X"10",X"91",X"C8",X"47",X"36",X"10",X"19",X"10",
		X"FB",X"C9",X"21",X"82",X"4B",X"11",X"E0",X"FF",X"3A",X"88",X"42",X"A7",X"C8",X"3D",X"4F",X"28",
		X"0D",X"FE",X"08",X"38",X"02",X"3E",X"08",X"4F",X"47",X"36",X"5F",X"19",X"10",X"FB",X"3E",X"08",
		X"91",X"C8",X"47",X"36",X"10",X"19",X"10",X"FB",X"C9",X"3E",X"1A",X"06",X"0B",X"F5",X"C5",X"CD",
		X"12",X"04",X"C1",X"F1",X"3C",X"10",X"F6",X"21",X"C7",X"49",X"11",X"20",X"00",X"06",X"0A",X"DD",
		X"21",X"00",X"42",X"DD",X"7E",X"00",X"4F",X"E6",X"0F",X"77",X"19",X"79",X"0F",X"0F",X"0F",X"0F",
		X"E6",X"0F",X"77",X"19",X"DD",X"23",X"DD",X"7E",X"00",X"4F",X"E6",X"0F",X"77",X"19",X"79",X"0F",
		X"0F",X"0F",X"0F",X"E6",X"0F",X"77",X"19",X"DD",X"23",X"DD",X"7E",X"00",X"4F",X"E6",X"0F",X"77",
		X"19",X"79",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"28",X"01",X"77",X"11",X"62",X"FF",X"19",X"11",
		X"20",X"00",X"DD",X"23",X"10",X"BD",X"CD",X"DA",X"02",X"C9",X"DD",X"21",X"C0",X"41",X"21",X"A7",
		X"48",X"0E",X"0A",X"11",X"20",X"00",X"06",X"03",X"DD",X"7E",X"00",X"77",X"19",X"DD",X"23",X"10",
		X"F7",X"11",X"A2",X"FF",X"19",X"0D",X"20",X"EB",X"C9",X"4F",X"3A",X"06",X"40",X"0F",X"D0",X"79",
		X"A7",X"28",X"47",X"CD",X"55",X"03",X"87",X"81",X"4F",X"06",X"00",X"21",X"64",X"03",X"09",X"A7",
		X"06",X"03",X"1A",X"8E",X"27",X"12",X"13",X"23",X"10",X"F8",X"D5",X"3A",X"0D",X"40",X"0F",X"30",
		X"02",X"3E",X"01",X"CD",X"CB",X"03",X"D1",X"1B",X"21",X"AA",X"40",X"06",X"03",X"1A",X"BE",X"D8",
		X"20",X"05",X"1B",X"2B",X"10",X"F7",X"C9",X"CD",X"55",X"03",X"21",X"A8",X"40",X"06",X"03",X"1A",
		X"77",X"13",X"23",X"10",X"FA",X"3E",X"02",X"C3",X"CB",X"03",X"CD",X"55",X"03",X"21",X"AB",X"40",
		X"A7",X"06",X"03",X"18",X"BD",X"F5",X"3A",X"0D",X"40",X"11",X"A2",X"40",X"0F",X"30",X"03",X"11",
		X"A5",X"40",X"F1",X"C9",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"07",X"00",X"00",X"05",X"00",
		X"50",X"04",X"00",X"00",X"04",X"00",X"80",X"03",X"00",X"50",X"03",X"00",X"30",X"03",X"00",X"00",
		X"03",X"00",X"80",X"02",X"00",X"50",X"02",X"00",X"30",X"02",X"00",X"00",X"02",X"00",X"80",X"01",
		X"00",X"50",X"01",X"00",X"30",X"01",X"00",X"00",X"01",X"00",X"00",X"01",X"00",X"00",X"02",X"00",
		X"00",X"04",X"00",X"00",X"08",X"00",X"00",X"16",X"00",X"00",X"32",X"00",X"00",X"64",X"00",X"00",
		X"50",X"00",X"F5",X"21",X"A2",X"40",X"A7",X"28",X"09",X"21",X"A5",X"40",X"3D",X"28",X"03",X"21",
		X"A8",X"40",X"36",X"00",X"23",X"36",X"00",X"23",X"36",X"00",X"F1",X"21",X"A4",X"40",X"DD",X"21",
		X"81",X"4B",X"A7",X"28",X"11",X"21",X"A7",X"40",X"DD",X"21",X"21",X"49",X"3D",X"28",X"07",X"21",
		X"AA",X"40",X"DD",X"21",X"41",X"4A",X"11",X"E0",X"FF",X"06",X"03",X"0E",X"04",X"7E",X"0F",X"0F",
		X"0F",X"0F",X"CD",X"FD",X"03",X"7E",X"CD",X"FD",X"03",X"2B",X"10",X"F1",X"C9",X"E6",X"0F",X"28",
		X"08",X"0E",X"00",X"DD",X"77",X"00",X"DD",X"19",X"C9",X"79",X"A7",X"28",X"F6",X"3E",X"10",X"0D",
		X"18",X"F1",X"87",X"F5",X"21",X"6E",X"21",X"E6",X"7F",X"5F",X"16",X"00",X"19",X"5E",X"23",X"56",
		X"EB",X"5E",X"23",X"56",X"23",X"EB",X"01",X"E0",X"FF",X"F1",X"38",X"0B",X"1A",X"FE",X"3F",X"C8",
		X"D6",X"30",X"77",X"13",X"09",X"18",X"F5",X"1A",X"FE",X"3F",X"C8",X"36",X"10",X"13",X"09",X"18",
		X"F6",X"3E",X"05",X"CD",X"12",X"04",X"3A",X"02",X"40",X"FE",X"63",X"38",X"02",X"3E",X"63",X"CD",
		X"65",X"04",X"47",X"E6",X"F0",X"28",X"07",X"0F",X"0F",X"0F",X"0F",X"32",X"9F",X"4A",X"78",X"E6",
		X"0F",X"32",X"7F",X"4A",X"C9",X"47",X"E6",X"0F",X"C6",X"00",X"27",X"4F",X"78",X"E6",X"F0",X"28",
		X"0B",X"0F",X"0F",X"0F",X"0F",X"47",X"AF",X"C6",X"16",X"27",X"10",X"FB",X"81",X"27",X"C9",X"21",
		X"FF",X"48",X"11",X"E0",X"FF",X"3A",X"85",X"42",X"FE",X"04",X"38",X"02",X"3E",X"04",X"4F",X"47",
		X"A7",X"28",X"05",X"36",X"2A",X"19",X"10",X"FB",X"3E",X"04",X"91",X"C8",X"47",X"36",X"10",X"19",
		X"10",X"FB",X"C9",X"F5",X"C5",X"D5",X"E5",X"08",X"D9",X"F5",X"C5",X"D5",X"E5",X"DD",X"E5",X"FD",
		X"E5",X"AF",X"32",X"01",X"68",X"21",X"20",X"40",X"11",X"00",X"50",X"01",X"40",X"00",X"ED",X"B0",
		X"11",X"5C",X"50",X"0E",X"04",X"ED",X"B0",X"11",X"40",X"50",X"0E",X"1C",X"ED",X"B0",X"3A",X"00",
		X"70",X"3A",X"15",X"40",X"32",X"16",X"40",X"3A",X"13",X"40",X"32",X"15",X"40",X"2A",X"10",X"40",
		X"22",X"13",X"40",X"21",X"12",X"40",X"3A",X"02",X"81",X"2F",X"77",X"2B",X"3A",X"01",X"81",X"2F",
		X"77",X"2B",X"3A",X"00",X"81",X"2F",X"77",X"21",X"80",X"41",X"35",X"21",X"5F",X"42",X"35",X"CD",
		X"3E",X"35",X"CD",X"6C",X"0A",X"21",X"17",X"05",X"E5",X"3A",X"05",X"40",X"EF",X"49",X"05",X"41",
		X"06",X"07",X"09",X"0E",X"0C",X"5B",X"0A",X"3A",X"1E",X"40",X"32",X"06",X"68",X"32",X"07",X"68",
		X"3A",X"80",X"41",X"E6",X"3F",X"20",X"0E",X"21",X"26",X"41",X"7E",X"A7",X"28",X"01",X"35",X"23",
		X"7E",X"A7",X"28",X"01",X"35",X"FD",X"E1",X"DD",X"E1",X"E1",X"D1",X"C1",X"F1",X"D9",X"08",X"E1",
		X"D1",X"C1",X"3E",X"01",X"32",X"01",X"68",X"F1",X"C9",X"06",X"20",X"CD",X"04",X"0D",X"C0",X"21",
		X"06",X"40",X"36",X"00",X"2B",X"36",X"01",X"AF",X"32",X"0A",X"40",X"21",X"81",X"05",X"CD",X"71",
		X"05",X"11",X"04",X"06",X"FF",X"11",X"00",X"05",X"FF",X"1E",X"02",X"FF",X"AF",X"32",X"51",X"46",
		X"C9",X"11",X"20",X"40",X"06",X"20",X"EB",X"36",X"00",X"2C",X"1A",X"77",X"2C",X"13",X"10",X"F7",
		X"C9",X"07",X"06",X"06",X"00",X"01",X"01",X"06",X"03",X"03",X"04",X"04",X"04",X"04",X"01",X"01",
		X"01",X"00",X"00",X"00",X"07",X"07",X"07",X"07",X"07",X"06",X"06",X"06",X"06",X"06",X"06",X"06",
		X"01",X"07",X"06",X"06",X"02",X"02",X"02",X"02",X"03",X"03",X"04",X"04",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"06",X"06",X"04",
		X"01",X"07",X"06",X"06",X"06",X"06",X"06",X"06",X"02",X"07",X"07",X"07",X"07",X"07",X"07",X"07",
		X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"04",X"06",X"06",X"04",
		X"01",X"07",X"06",X"06",X"04",X"01",X"07",X"07",X"07",X"07",X"07",X"07",X"06",X"06",X"06",X"06",
		X"04",X"04",X"04",X"04",X"01",X"01",X"01",X"01",X"03",X"03",X"03",X"03",X"06",X"06",X"06",X"04",
		X"01",X"07",X"06",X"06",X"01",X"01",X"01",X"01",X"01",X"02",X"02",X"03",X"03",X"04",X"04",X"05",
		X"05",X"06",X"06",X"07",X"07",X"01",X"01",X"02",X"02",X"01",X"01",X"01",X"04",X"06",X"06",X"04",
		X"01",X"07",X"06",X"06",X"04",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"04",
		X"01",X"21",X"D9",X"08",X"E5",X"3A",X"51",X"46",X"EF",X"65",X"06",X"88",X"06",X"C7",X"06",X"E1",
		X"06",X"F1",X"06",X"CB",X"07",X"F7",X"07",X"1B",X"08",X"63",X"08",X"63",X"08",X"69",X"08",X"A5",
		X"08",X"E1",X"06",X"CA",X"08",X"AF",X"32",X"03",X"68",X"32",X"19",X"40",X"21",X"60",X"40",X"11",
		X"61",X"40",X"01",X"3F",X"00",X"36",X"00",X"ED",X"B0",X"CD",X"19",X"0D",X"21",X"51",X"46",X"34",
		X"AF",X"32",X"06",X"40",X"CD",X"EB",X"0C",X"C9",X"06",X"1D",X"CD",X"04",X"0D",X"C0",X"21",X"A1",
		X"05",X"CD",X"71",X"05",X"AF",X"32",X"07",X"68",X"32",X"06",X"68",X"CD",X"5C",X"0A",X"11",X"11",
		X"06",X"FF",X"11",X"0B",X"06",X"FF",X"1E",X"0C",X"FF",X"3E",X"0C",X"32",X"40",X"46",X"3E",X"03",
		X"32",X"80",X"42",X"21",X"6E",X"19",X"22",X"BB",X"40",X"21",X"C0",X"42",X"06",X"80",X"3E",X"FF",
		X"D7",X"21",X"51",X"46",X"36",X"0A",X"C9",X"21",X"50",X"46",X"35",X"C0",X"2C",X"34",X"21",X"E1",
		X"05",X"CD",X"71",X"05",X"11",X"8B",X"06",X"FF",X"11",X"8C",X"06",X"FF",X"11",X"00",X"02",X"FF",
		X"C9",X"21",X"50",X"46",X"35",X"C0",X"CD",X"EB",X"0C",X"CD",X"19",X"0D",X"21",X"51",X"46",X"34",
		X"C9",X"06",X"19",X"CD",X"04",X"0D",X"C0",X"21",X"C1",X"05",X"CD",X"71",X"05",X"11",X"0D",X"06",
		X"FF",X"21",X"80",X"45",X"AF",X"06",X"C0",X"D7",X"21",X"64",X"07",X"11",X"70",X"07",X"DD",X"21",
		X"98",X"45",X"CD",X"4B",X"07",X"01",X"18",X"00",X"DD",X"09",X"1A",X"3C",X"20",X"F4",X"21",X"7D",
		X"07",X"22",X"54",X"46",X"21",X"4A",X"4A",X"22",X"56",X"46",X"21",X"50",X"46",X"36",X"32",X"2C",
		X"34",X"2C",X"36",X"0D",X"2C",X"36",X"06",X"DD",X"21",X"98",X"45",X"06",X"06",X"11",X"18",X"00",
		X"CD",X"1B",X"32",X"DD",X"19",X"10",X"F9",X"CD",X"1E",X"11",X"C9",X"1A",X"DD",X"77",X"06",X"13",
		X"1A",X"13",X"DD",X"77",X"04",X"7E",X"DD",X"77",X"0C",X"23",X"7E",X"DD",X"77",X"0D",X"DD",X"36",
		X"0E",X"00",X"23",X"C9",X"E3",X"17",X"E6",X"33",X"6B",X"18",X"27",X"18",X"2A",X"34",X"AF",X"18",
		X"0A",X"0A",X"0A",X"0D",X"0A",X"10",X"0A",X"13",X"0A",X"16",X"0A",X"19",X"FF",X"0F",X"0F",X"0F",
		X"10",X"10",X"13",X"1F",X"20",X"19",X"15",X"22",X"10",X"10",X"0F",X"0F",X"0F",X"10",X"10",X"20",
		X"1F",X"1C",X"19",X"13",X"15",X"10",X"10",X"0F",X"0F",X"0F",X"10",X"10",X"24",X"18",X"19",X"15",
		X"16",X"10",X"10",X"10",X"0F",X"0F",X"0F",X"10",X"10",X"22",X"25",X"23",X"24",X"1C",X"15",X"22",
		X"10",X"0F",X"0F",X"0F",X"10",X"10",X"13",X"11",X"24",X"24",X"1C",X"15",X"10",X"10",X"0F",X"0F",
		X"0F",X"10",X"10",X"24",X"18",X"19",X"15",X"16",X"10",X"10",X"10",X"CD",X"37",X"07",X"21",X"50",
		X"46",X"35",X"C0",X"36",X"05",X"2A",X"54",X"46",X"7E",X"23",X"22",X"54",X"46",X"2A",X"56",X"46",
		X"77",X"11",X"E0",X"FF",X"19",X"22",X"56",X"46",X"21",X"52",X"46",X"35",X"C0",X"36",X"0D",X"21",
		X"50",X"46",X"36",X"14",X"2C",X"34",X"C9",X"CD",X"37",X"07",X"21",X"50",X"46",X"35",X"C0",X"36",
		X"01",X"2C",X"35",X"2A",X"56",X"46",X"11",X"A3",X"01",X"19",X"22",X"56",X"46",X"21",X"53",X"46",
		X"35",X"C0",X"21",X"50",X"46",X"36",X"96",X"2C",X"34",X"34",X"C9",X"21",X"00",X"00",X"22",X"0D",
		X"40",X"AF",X"32",X"0A",X"40",X"3E",X"03",X"32",X"05",X"40",X"3E",X"00",X"32",X"06",X"40",X"CD",
		X"16",X"0A",X"3E",X"03",X"32",X"05",X"40",X"21",X"7F",X"41",X"34",X"7E",X"E6",X"01",X"20",X"06",
		X"3E",X"00",X"32",X"0A",X"40",X"C9",X"CD",X"62",X"0C",X"3E",X"01",X"32",X"80",X"43",X"32",X"83",
		X"43",X"32",X"0A",X"40",X"21",X"C0",X"43",X"06",X"80",X"3E",X"FF",X"D7",X"21",X"F7",X"43",X"CD",
		X"4E",X"0A",X"C9",X"21",X"51",X"46",X"36",X"00",X"C9",X"3E",X"1D",X"32",X"48",X"46",X"21",X"40",
		X"46",X"4E",X"3E",X"10",X"32",X"0A",X"40",X"CD",X"94",X"24",X"21",X"48",X"46",X"35",X"20",X"F7",
		X"21",X"40",X"46",X"34",X"7E",X"FE",X"1A",X"D8",X"21",X"51",X"46",X"34",X"2B",X"36",X"3C",X"CD",
		X"77",X"3F",X"E6",X"07",X"FE",X"06",X"38",X"02",X"D6",X"06",X"CD",X"24",X"14",X"21",X"CC",X"45",
		X"7E",X"C6",X"07",X"77",X"C9",X"21",X"50",X"46",X"7E",X"A7",X"28",X"03",X"35",X"18",X"0A",X"DD",
		X"21",X"C8",X"45",X"CD",X"F9",X"2D",X"CD",X"0D",X"28",X"CD",X"1E",X"11",X"3A",X"6F",X"40",X"FE",
		X"CD",X"D8",X"21",X"51",X"46",X"34",X"2B",X"36",X"3C",X"C9",X"06",X"19",X"CD",X"04",X"0D",X"C0",
		X"21",X"51",X"46",X"36",X"02",X"2B",X"36",X"1E",X"C9",X"3A",X"0C",X"41",X"FE",X"0F",X"20",X"19",
		X"3A",X"11",X"40",X"CB",X"7F",X"28",X"09",X"CD",X"F1",X"0A",X"21",X"00",X"00",X"C3",X"D6",X"09",
		X"CB",X"77",X"C8",X"CD",X"F1",X"0A",X"C3",X"D3",X"09",X"3A",X"02",X"40",X"A7",X"C8",X"21",X"05",
		X"40",X"34",X"AF",X"32",X"0A",X"40",X"C9",X"21",X"BD",X"09",X"E5",X"3A",X"0A",X"40",X"EF",X"15",
		X"09",X"41",X"09",X"A6",X"09",X"AF",X"32",X"19",X"40",X"32",X"03",X"68",X"21",X"40",X"50",X"06",
		X"40",X"AF",X"D7",X"32",X"06",X"40",X"21",X"02",X"48",X"22",X"0B",X"40",X"21",X"09",X"40",X"36",
		X"10",X"23",X"34",X"21",X"60",X"40",X"11",X"61",X"40",X"01",X"1F",X"00",X"36",X"00",X"ED",X"B0",
		X"C9",X"2A",X"0B",X"40",X"06",X"1D",X"3E",X"10",X"D7",X"11",X"03",X"00",X"19",X"06",X"1D",X"D7",
		X"19",X"22",X"0B",X"40",X"21",X"09",X"40",X"35",X"C0",X"2C",X"34",X"21",X"81",X"05",X"CD",X"71",
		X"05",X"AF",X"32",X"07",X"68",X"32",X"06",X"68",X"32",X"0D",X"40",X"CD",X"5C",X"0A",X"11",X"01",
		X"06",X"FF",X"1E",X"11",X"FF",X"1E",X"0C",X"FF",X"1E",X"16",X"FF",X"1C",X"3A",X"00",X"40",X"E6",
		X"02",X"28",X"02",X"1E",X"28",X"FF",X"1E",X"2A",X"3A",X"00",X"40",X"E6",X"02",X"28",X"01",X"1D",
		X"FF",X"3A",X"17",X"40",X"47",X"E6",X"0F",X"32",X"78",X"49",X"78",X"E6",X"F0",X"C8",X"0F",X"0F",
		X"0F",X"0F",X"32",X"98",X"49",X"C9",X"3A",X"02",X"40",X"A7",X"C8",X"3D",X"11",X"18",X"06",X"28",
		X"01",X"1C",X"FF",X"11",X"00",X"03",X"FF",X"3E",X"02",X"32",X"05",X"40",X"C9",X"3A",X"11",X"40",
		X"CB",X"7F",X"C2",X"00",X"0A",X"CB",X"77",X"C8",X"3A",X"02",X"40",X"FE",X"02",X"D8",X"D6",X"02",
		X"32",X"02",X"40",X"21",X"00",X"01",X"22",X"0D",X"40",X"CD",X"5C",X"0A",X"AF",X"32",X"0A",X"40",
		X"3E",X"03",X"32",X"05",X"40",X"3E",X"01",X"32",X"06",X"40",X"11",X"04",X"06",X"FF",X"CD",X"16",
		X"0A",X"CD",X"E1",X"0B",X"11",X"00",X"04",X"FF",X"3A",X"0E",X"40",X"0F",X"D0",X"1C",X"FF",X"C9",
		X"3A",X"02",X"40",X"A7",X"28",X"0A",X"3D",X"32",X"02",X"40",X"21",X"00",X"00",X"C3",X"D6",X"09",
		X"3E",X"01",X"32",X"05",X"40",X"C9",X"21",X"80",X"42",X"AF",X"06",X"40",X"D7",X"21",X"6E",X"19",
		X"11",X"C0",X"43",X"0E",X"80",X"ED",X"B0",X"21",X"F7",X"43",X"CD",X"4E",X"0A",X"21",X"6E",X"19",
		X"11",X"C0",X"44",X"0E",X"80",X"ED",X"B0",X"21",X"F7",X"44",X"CD",X"4E",X"0A",X"21",X"60",X"40",
		X"06",X"20",X"AF",X"D7",X"3A",X"07",X"40",X"32",X"88",X"43",X"32",X"88",X"44",X"C9",X"11",X"04",
		X"00",X"06",X"06",X"3E",X"FB",X"A6",X"77",X"19",X"10",X"F9",X"C9",X"C9",X"11",X"01",X"07",X"FF",
		X"3A",X"0C",X"41",X"FE",X"0F",X"20",X"04",X"11",X"06",X"06",X"FF",X"C9",X"11",X"41",X"42",X"1A",
		X"6F",X"26",X"42",X"7E",X"FE",X"FF",X"C8",X"47",X"3A",X"00",X"40",X"E6",X"01",X"20",X"06",X"3A",
		X"06",X"40",X"A7",X"28",X"04",X"78",X"CD",X"B6",X"0A",X"36",X"FF",X"7D",X"FE",X"5E",X"28",X"03",
		X"3C",X"12",X"C9",X"3E",X"43",X"12",X"C9",X"3A",X"42",X"42",X"F6",X"10",X"32",X"42",X"42",X"32",
		X"01",X"82",X"AF",X"C3",X"B6",X"0A",X"AF",X"CD",X"B6",X"0A",X"3A",X"42",X"42",X"E6",X"EF",X"32",
		X"42",X"42",X"32",X"01",X"82",X"C9",X"32",X"00",X"82",X"3A",X"42",X"42",X"E6",X"F7",X"32",X"01",
		X"82",X"00",X"00",X"00",X"00",X"3A",X"42",X"42",X"F6",X"08",X"32",X"01",X"82",X"C9",X"47",X"3A",
		X"06",X"40",X"A7",X"C8",X"78",X"C5",X"D5",X"E5",X"47",X"11",X"40",X"42",X"1A",X"6F",X"26",X"42",
		X"70",X"7D",X"FE",X"5E",X"28",X"04",X"3C",X"12",X"18",X"03",X"3E",X"43",X"12",X"E1",X"D1",X"C1",
		X"C9",X"AF",X"18",X"C2",X"3E",X"10",X"18",X"BE",X"3A",X"80",X"42",X"E6",X"01",X"28",X"09",X"3E",
		X"01",X"CD",X"CE",X"0A",X"3E",X"02",X"18",X"C6",X"3E",X"06",X"18",X"C2",X"3E",X"04",X"18",X"BE",
		X"3E",X"05",X"18",X"C1",X"3E",X"07",X"CD",X"CE",X"0A",X"3E",X"08",X"18",X"B1",X"3E",X"25",X"CD",
		X"CE",X"0A",X"3E",X"26",X"CD",X"CE",X"0A",X"3E",X"27",X"C3",X"CE",X"0A",X"3E",X"09",X"C3",X"CE",
		X"0A",X"3E",X"28",X"CD",X"CE",X"0A",X"3E",X"29",X"CD",X"CE",X"0A",X"3E",X"2A",X"C3",X"CE",X"0A",
		X"3E",X"22",X"CD",X"CE",X"0A",X"3E",X"23",X"CD",X"CE",X"0A",X"3E",X"24",X"C3",X"CE",X"0A",X"DD",
		X"7E",X"04",X"FE",X"10",X"06",X"03",X"38",X"08",X"FE",X"18",X"06",X"0E",X"38",X"02",X"06",X"0F",
		X"78",X"C3",X"D5",X"0A",X"3E",X"0A",X"C3",X"D5",X"0A",X"3E",X"0D",X"C3",X"CE",X"0A",X"3E",X"2B",
		X"CD",X"CE",X"0A",X"3E",X"2C",X"CD",X"CE",X"0A",X"3E",X"2D",X"C3",X"CE",X"0A",X"3E",X"0C",X"C3",
		X"CE",X"0A",X"3E",X"1C",X"CD",X"CE",X"0A",X"3E",X"1D",X"CD",X"CE",X"0A",X"3E",X"1E",X"C3",X"CE",
		X"0A",X"3E",X"1F",X"CD",X"CE",X"0A",X"3E",X"20",X"CD",X"CE",X"0A",X"3E",X"21",X"C3",X"CE",X"0A",
		X"3E",X"A5",X"CD",X"CE",X"0A",X"3E",X"A6",X"CD",X"CE",X"0A",X"3E",X"A7",X"C3",X"CE",X"0A",X"3E",
		X"A8",X"CD",X"CE",X"0A",X"3E",X"A9",X"CD",X"CE",X"0A",X"3E",X"AA",X"C3",X"CE",X"0A",X"3E",X"A2",
		X"CD",X"CE",X"0A",X"3E",X"A3",X"CD",X"CE",X"0A",X"3E",X"A4",X"C3",X"CE",X"0A",X"3E",X"AB",X"CD",
		X"CE",X"0A",X"3E",X"AC",X"CD",X"CE",X"0A",X"3E",X"AD",X"C3",X"CE",X"0A",X"3E",X"0B",X"C3",X"D5",
		X"0A",X"3E",X"13",X"CD",X"CE",X"0A",X"3E",X"14",X"CD",X"CE",X"0A",X"3E",X"15",X"C3",X"CE",X"0A",
		X"3E",X"16",X"CD",X"CE",X"0A",X"3E",X"17",X"CD",X"CE",X"0A",X"3E",X"18",X"C3",X"CE",X"0A",X"3E",
		X"19",X"CD",X"CE",X"0A",X"3E",X"1A",X"CD",X"CE",X"0A",X"3E",X"1B",X"C3",X"CE",X"0A",X"21",X"45",
		X"0C",X"E5",X"3A",X"0A",X"40",X"EF",X"62",X"0C",X"D5",X"0C",X"25",X"0D",X"F0",X"0D",X"F4",X"0D",
		X"48",X"0E",X"55",X"0E",X"99",X"0E",X"15",X"0F",X"1E",X"0F",X"27",X"0F",X"50",X"0F",X"AA",X"0F",
		X"B9",X"0F",X"50",X"0F",X"CD",X"0F",X"E8",X"0F",X"24",X"10",X"48",X"10",X"85",X"10",X"BA",X"10",
		X"0A",X"11",X"FF",X"FF",X"FF",X"3A",X"06",X"40",X"A7",X"C0",X"3A",X"0C",X"41",X"FE",X"0F",X"CA",
		X"D9",X"08",X"3A",X"02",X"40",X"A7",X"C8",X"21",X"05",X"40",X"36",X"02",X"21",X"0A",X"40",X"36",
		X"00",X"C9",X"21",X"39",X"19",X"7E",X"D6",X"06",X"32",X"81",X"43",X"32",X"81",X"44",X"23",X"7E",
		X"32",X"82",X"43",X"32",X"82",X"44",X"3E",X"03",X"32",X"85",X"43",X"32",X"85",X"44",X"AF",X"32",
		X"80",X"43",X"32",X"80",X"44",X"32",X"83",X"43",X"32",X"83",X"44",X"21",X"80",X"45",X"11",X"81",
		X"45",X"01",X"C0",X"00",X"77",X"ED",X"B0",X"32",X"BD",X"40",X"CD",X"1E",X"11",X"06",X"0E",X"3A",
		X"0E",X"40",X"A7",X"20",X"02",X"06",X"1C",X"78",X"32",X"10",X"41",X"21",X"0A",X"40",X"34",X"C9",
		X"21",X"C0",X"42",X"11",X"42",X"0C",X"06",X"20",X"CD",X"C2",X"0C",X"21",X"F7",X"42",X"CD",X"4E",
		X"0A",X"C9",X"1A",X"77",X"13",X"23",X"1A",X"77",X"23",X"1A",X"77",X"13",X"23",X"1A",X"77",X"1B",
		X"1B",X"23",X"10",X"EE",X"C9",X"CD",X"19",X"0D",X"CD",X"C4",X"11",X"CD",X"D9",X"11",X"3E",X"02",
		X"32",X"0A",X"40",X"21",X"F0",X"41",X"06",X"10",X"AF",X"D7",X"C9",X"21",X"60",X"40",X"06",X"20",
		X"AF",X"77",X"23",X"10",X"FC",X"21",X"80",X"45",X"06",X"C0",X"77",X"23",X"10",X"FC",X"C9",X"CD",
		X"EB",X"0C",X"06",X"1C",X"3E",X"20",X"90",X"5F",X"16",X"00",X"2A",X"0B",X"40",X"3E",X"10",X"D7",
		X"19",X"22",X"0B",X"40",X"21",X"09",X"40",X"35",X"C9",X"21",X"03",X"48",X"22",X"0B",X"40",X"3E",
		X"20",X"32",X"09",X"40",X"C9",X"3A",X"1A",X"40",X"A7",X"20",X"07",X"CD",X"FF",X"0C",X"C0",X"CD",
		X"19",X"0D",X"3A",X"0E",X"40",X"A7",X"28",X"2F",X"21",X"1A",X"40",X"7E",X"A7",X"28",X"06",X"34",
		X"FE",X"80",X"28",X"23",X"C9",X"4F",X"11",X"02",X"06",X"3A",X"0D",X"40",X"A7",X"28",X"02",X"0C",
		X"1C",X"FF",X"3A",X"0F",X"40",X"A7",X"20",X"04",X"79",X"32",X"1E",X"40",X"21",X"1A",X"40",X"34",
		X"3A",X"0D",X"40",X"32",X"BD",X"40",X"C9",X"AF",X"32",X"1A",X"40",X"11",X"82",X"06",X"FF",X"1C",
		X"FF",X"11",X"0A",X"06",X"FF",X"16",X"08",X"FF",X"11",X"80",X"42",X"21",X"80",X"43",X"3A",X"0D",
		X"40",X"A7",X"28",X"03",X"21",X"80",X"44",X"01",X"C0",X"00",X"ED",X"B0",X"21",X"49",X"19",X"3A",
		X"80",X"42",X"E6",X"07",X"47",X"CD",X"2B",X"2C",X"ED",X"53",X"BB",X"40",X"78",X"21",X"E8",X"0D",
		X"85",X"30",X"01",X"24",X"6F",X"7E",X"21",X"25",X"40",X"36",X"06",X"2C",X"2C",X"06",X"1C",X"77",
		X"2C",X"2C",X"10",X"FB",X"CD",X"5C",X"0A",X"3E",X"1D",X"32",X"48",X"46",X"3E",X"03",X"32",X"0A",
		X"40",X"CD",X"1E",X"11",X"16",X"00",X"FF",X"16",X"01",X"FF",X"3A",X"80",X"42",X"FE",X"01",X"D0",
		X"3A",X"83",X"42",X"A7",X"C0",X"CD",X"B0",X"0C",X"3E",X"01",X"32",X"83",X"42",X"21",X"89",X"42",
		X"06",X"04",X"36",X"00",X"23",X"10",X"FB",X"C9",X"00",X"02",X"01",X"03",X"00",X"02",X"01",X"03",
		X"CD",X"8B",X"13",X"C9",X"CD",X"31",X"13",X"CD",X"C0",X"25",X"3A",X"F1",X"41",X"A7",X"20",X"06",
		X"CD",X"7A",X"2D",X"CD",X"69",X"3C",X"CD",X"67",X"12",X"CD",X"1E",X"11",X"CD",X"16",X"2D",X"2A",
		X"81",X"42",X"7D",X"B4",X"28",X"11",X"3A",X"4F",X"43",X"A7",X"C8",X"3E",X"07",X"32",X"0A",X"40",
		X"CD",X"AF",X"0B",X"CD",X"A0",X"0B",X"C9",X"32",X"5F",X"42",X"3C",X"32",X"10",X"41",X"21",X"0A",
		X"40",X"34",X"3A",X"80",X"42",X"E6",X"01",X"28",X"0A",X"CD",X"AF",X"0B",X"CD",X"CD",X"0B",X"CD",
		X"F0",X"0B",X"C9",X"CD",X"A0",X"0B",X"18",X"F4",X"CD",X"31",X"13",X"3A",X"5F",X"42",X"A7",X"C0",
		X"21",X"0A",X"40",X"34",X"C9",X"CD",X"DD",X"0D",X"21",X"80",X"42",X"34",X"7E",X"E6",X"07",X"11",
		X"39",X"19",X"87",X"83",X"5F",X"30",X"01",X"14",X"1A",X"23",X"D6",X"06",X"77",X"23",X"13",X"1A",
		X"77",X"3E",X"03",X"32",X"85",X"42",X"3A",X"80",X"42",X"21",X"49",X"19",X"E6",X"07",X"87",X"5F",
		X"16",X"00",X"19",X"5E",X"23",X"56",X"ED",X"53",X"6E",X"43",X"CD",X"B0",X"0C",X"CD",X"AF",X"11",
		X"3E",X"10",X"32",X"0A",X"40",X"CD",X"19",X"0D",X"C9",X"CD",X"7A",X"2D",X"CD",X"C0",X"25",X"CD",
		X"69",X"3C",X"CD",X"1E",X"11",X"21",X"91",X"45",X"35",X"C0",X"3A",X"06",X"40",X"A7",X"28",X"3B",
		X"CD",X"CD",X"0B",X"3E",X"01",X"32",X"10",X"41",X"21",X"88",X"42",X"35",X"3E",X"03",X"32",X"85",
		X"42",X"CD",X"AF",X"11",X"3A",X"0D",X"40",X"A7",X"20",X"2D",X"3A",X"88",X"43",X"A7",X"28",X"12",
		X"3A",X"0E",X"40",X"A7",X"28",X"2D",X"3A",X"88",X"44",X"A7",X"28",X"27",X"3E",X"09",X"32",X"0A",
		X"40",X"C9",X"3E",X"0A",X"32",X"0A",X"40",X"CD",X"FF",X"0B",X"C9",X"AF",X"32",X"51",X"46",X"32",
		X"0A",X"40",X"3C",X"32",X"05",X"40",X"C9",X"3A",X"88",X"44",X"A7",X"28",X"0F",X"3A",X"88",X"43",
		X"A7",X"28",X"D9",X"3E",X"08",X"32",X"0A",X"40",X"CD",X"CD",X"0B",X"C9",X"3E",X"0D",X"32",X"0A",
		X"40",X"CD",X"FF",X"0B",X"C9",X"AF",X"32",X"0D",X"40",X"3C",X"32",X"0A",X"40",X"C9",X"3E",X"01",
		X"32",X"0D",X"40",X"32",X"0A",X"40",X"C9",X"CD",X"FF",X"0C",X"C0",X"CD",X"19",X"0D",X"CD",X"E1",
		X"11",X"11",X"02",X"06",X"FF",X"1E",X"00",X"FF",X"3E",X"78",X"32",X"5F",X"42",X"3E",X"FF",X"32",
		X"BE",X"40",X"CD",X"A0",X"0B",X"CD",X"AF",X"0B",X"CD",X"BE",X"0B",X"21",X"0A",X"40",X"34",X"C9",
		X"3A",X"5F",X"42",X"A7",X"20",X"33",X"3A",X"BF",X"40",X"A7",X"28",X"E6",X"3E",X"82",X"CD",X"12",
		X"04",X"3E",X"80",X"CD",X"12",X"04",X"CD",X"79",X"02",X"21",X"E1",X"05",X"CD",X"71",X"05",X"21",
		X"2B",X"40",X"3A",X"BF",X"40",X"47",X"2C",X"2C",X"2C",X"2C",X"10",X"FA",X"36",X"04",X"22",X"FD",
		X"41",X"AF",X"32",X"BF",X"40",X"32",X"FF",X"41",X"C9",X"21",X"BE",X"40",X"7E",X"FE",X"80",X"30",
		X"15",X"E6",X"07",X"20",X"11",X"3A",X"FF",X"41",X"ED",X"5B",X"FD",X"41",X"12",X"3C",X"FE",X"08",
		X"38",X"01",X"AF",X"32",X"FF",X"41",X"35",X"C0",X"18",X"98",X"3A",X"0E",X"40",X"A7",X"28",X"26",
		X"3A",X"88",X"44",X"A7",X"28",X"20",X"C3",X"DC",X"0E",X"CD",X"FF",X"0C",X"C0",X"CD",X"19",X"0D",
		X"CD",X"E1",X"11",X"11",X"03",X"06",X"FF",X"1E",X"00",X"FF",X"C3",X"35",X"0F",X"3A",X"88",X"43",
		X"A7",X"28",X"03",X"C3",X"03",X"0F",X"AF",X"32",X"06",X"40",X"32",X"1E",X"40",X"32",X"0A",X"40",
		X"32",X"51",X"46",X"3C",X"32",X"05",X"40",X"C9",X"CD",X"FF",X"0C",X"C0",X"16",X"01",X"FF",X"AF",
		X"32",X"F1",X"41",X"3E",X"05",X"32",X"40",X"46",X"3E",X"01",X"32",X"80",X"42",X"21",X"6C",X"43",
		X"36",X"78",X"21",X"E1",X"05",X"CD",X"71",X"05",X"11",X"25",X"06",X"FF",X"1C",X"FF",X"1C",X"FF",
		X"1E",X"11",X"FF",X"21",X"6C",X"40",X"36",X"48",X"23",X"36",X"21",X"23",X"36",X"05",X"23",X"36",
		X"75",X"C3",X"4B",X"0F",X"21",X"6C",X"43",X"35",X"7E",X"FE",X"02",X"28",X"0F",X"A7",X"C0",X"21",
		X"21",X"06",X"CD",X"71",X"05",X"AF",X"32",X"6C",X"40",X"C3",X"4B",X"0F",X"11",X"A5",X"06",X"FF",
		X"1C",X"FF",X"1C",X"FF",X"1E",X"91",X"FF",X"C9",X"3E",X"1D",X"32",X"48",X"46",X"21",X"40",X"46",
		X"4E",X"CD",X"94",X"24",X"21",X"48",X"46",X"35",X"20",X"F7",X"21",X"40",X"46",X"34",X"7E",X"FE",
		X"1D",X"D8",X"21",X"6C",X"43",X"36",X"00",X"23",X"36",X"3C",X"AF",X"CD",X"24",X"14",X"CD",X"77",
		X"3F",X"E6",X"07",X"FE",X"06",X"38",X"02",X"D6",X"06",X"CD",X"6F",X"14",X"CD",X"7D",X"0B",X"CD",
		X"1E",X"11",X"C3",X"4B",X"0F",X"3A",X"1E",X"40",X"A7",X"3A",X"10",X"40",X"28",X"03",X"3A",X"11",
		X"40",X"E6",X"08",X"C2",X"4B",X"0F",X"21",X"6C",X"43",X"34",X"7E",X"E6",X"07",X"20",X"17",X"7E",
		X"0F",X"0F",X"0F",X"E6",X"07",X"FE",X"06",X"38",X"02",X"AF",X"77",X"23",X"35",X"CA",X"4B",X"0F",
		X"CD",X"24",X"14",X"CD",X"7D",X"0B",X"CD",X"1E",X"11",X"C9",X"DD",X"21",X"C8",X"45",X"CD",X"F9",
		X"2D",X"CD",X"0D",X"28",X"CD",X"1E",X"11",X"3A",X"6F",X"40",X"21",X"6B",X"40",X"BE",X"D8",X"3A",
		X"6C",X"40",X"21",X"68",X"40",X"96",X"30",X"02",X"ED",X"44",X"FE",X"03",X"38",X"0D",X"CD",X"42",
		X"0F",X"3E",X"1F",X"32",X"6D",X"40",X"CD",X"91",X"0B",X"18",X"19",X"CD",X"42",X"0F",X"3E",X"1E",
		X"32",X"6D",X"40",X"3E",X"3C",X"32",X"69",X"40",X"3E",X"06",X"32",X"6A",X"40",X"11",X"19",X"03",
		X"FF",X"CD",X"82",X"0B",X"21",X"6C",X"43",X"36",X"78",X"C9",X"21",X"6C",X"43",X"35",X"C0",X"2A",
		X"6E",X"43",X"22",X"BB",X"40",X"3E",X"01",X"32",X"0A",X"40",X"32",X"10",X"41",X"C9",X"21",X"60",
		X"40",X"DD",X"21",X"80",X"45",X"11",X"18",X"00",X"DD",X"7E",X"06",X"D6",X"0B",X"77",X"DD",X"7E",
		X"0F",X"2C",X"77",X"DD",X"7E",X"10",X"2C",X"77",X"DD",X"7E",X"04",X"2C",X"D6",X"06",X"77",X"2C",
		X"DD",X"19",X"3A",X"F1",X"41",X"A7",X"C2",X"3B",X"12",X"06",X"07",X"DD",X"4E",X"05",X"DD",X"7E",
		X"06",X"CB",X"01",X"17",X"CB",X"01",X"17",X"CB",X"01",X"17",X"D6",X"08",X"77",X"2C",X"DD",X"7E",
		X"0F",X"77",X"2C",X"DD",X"7E",X"10",X"77",X"2C",X"DD",X"7E",X"04",X"DD",X"4E",X"03",X"CB",X"01",
		X"17",X"CB",X"01",X"17",X"CB",X"01",X"17",X"D6",X"08",X"77",X"2C",X"DD",X"19",X"10",X"CC",X"CD",
		X"94",X"11",X"3A",X"1E",X"40",X"A7",X"C0",X"21",X"64",X"40",X"11",X"04",X"00",X"06",X"03",X"34",
		X"19",X"10",X"FC",X"C9",X"21",X"63",X"40",X"3A",X"61",X"40",X"47",X"E6",X"3F",X"FE",X"34",X"28",
		X"06",X"FE",X"35",X"28",X"02",X"34",X"C9",X"CB",X"70",X"C0",X"7E",X"C6",X"02",X"77",X"C9",X"21",
		X"80",X"42",X"11",X"80",X"43",X"3A",X"0D",X"40",X"A7",X"28",X"03",X"11",X"80",X"44",X"01",X"C0",
		X"00",X"ED",X"B0",X"C9",X"21",X"40",X"43",X"06",X"40",X"AF",X"D7",X"AF",X"21",X"40",X"44",X"06",
		X"40",X"D7",X"21",X"40",X"45",X"06",X"40",X"D7",X"C9",X"21",X"B0",X"45",X"06",X"90",X"AF",X"D7",
		X"C9",X"01",X"1E",X"00",X"11",X"03",X"00",X"6A",X"DD",X"21",X"A2",X"40",X"3A",X"0D",X"40",X"0F",
		X"30",X"02",X"DD",X"19",X"FD",X"21",X"00",X"42",X"DD",X"7E",X"02",X"FD",X"BE",X"02",X"20",X"0E",
		X"DD",X"7E",X"01",X"FD",X"BE",X"01",X"20",X"06",X"DD",X"7E",X"00",X"FD",X"BE",X"00",X"30",X"09",
		X"FD",X"19",X"2C",X"0D",X"0D",X"0D",X"C8",X"18",X"DF",X"7D",X"3C",X"32",X"BF",X"40",X"3D",X"21",
		X"1D",X"42",X"11",X"20",X"42",X"ED",X"B8",X"6F",X"DD",X"7E",X"00",X"FD",X"77",X"00",X"DD",X"7E",
		X"01",X"FD",X"77",X"01",X"DD",X"7E",X"02",X"FD",X"77",X"02",X"C9",X"21",X"67",X"40",X"06",X"07",
		X"ED",X"5B",X"F2",X"41",X"1A",X"4F",X"FE",X"80",X"20",X"09",X"AF",X"21",X"F0",X"41",X"77",X"2C",
		X"77",X"18",X"10",X"11",X"04",X"00",X"79",X"86",X"77",X"19",X"10",X"FA",X"2A",X"F2",X"41",X"23",
		X"22",X"F2",X"41",X"CD",X"94",X"11",X"C9",X"CD",X"6B",X"12",X"C9",X"3A",X"F9",X"41",X"A7",X"20",
		X"37",X"3A",X"F5",X"41",X"A7",X"C0",X"21",X"F1",X"41",X"7E",X"A7",X"C0",X"3A",X"85",X"42",X"A7",
		X"C8",X"2B",X"7E",X"A7",X"28",X"02",X"35",X"C9",X"3A",X"06",X"40",X"A7",X"C8",X"3A",X"10",X"40",
		X"47",X"AF",X"21",X"0F",X"40",X"B6",X"20",X"0D",X"2D",X"B6",X"28",X"09",X"2D",X"7E",X"A7",X"28",
		X"04",X"3A",X"11",X"40",X"47",X"CB",X"58",X"C8",X"21",X"86",X"42",X"7E",X"4F",X"FE",X"0C",X"38",
		X"02",X"36",X"00",X"34",X"21",X"17",X"13",X"3A",X"80",X"42",X"E6",X"01",X"20",X"03",X"21",X"24",
		X"13",X"79",X"E7",X"21",X"65",X"40",X"11",X"04",X"00",X"06",X"07",X"77",X"19",X"10",X"FC",X"3E",
		X"80",X"32",X"F0",X"41",X"3E",X"01",X"32",X"F1",X"41",X"21",X"F2",X"12",X"22",X"F2",X"41",X"CD",
		X"DC",X"0B",X"AF",X"32",X"F9",X"41",X"21",X"85",X"42",X"7E",X"A7",X"28",X"01",X"35",X"16",X"08",
		X"FF",X"C9",X"FA",X"FC",X"FD",X"FE",X"FE",X"FF",X"FF",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"01",X"00",X"01",X"01",X"01",
		X"01",X"02",X"02",X"03",X"04",X"06",X"80",X"1D",X"9D",X"1F",X"9F",X"1E",X"5E",X"20",X"A0",X"1E",
		X"9F",X"1D",X"9D",X"5E",X"27",X"29",X"26",X"76",X"27",X"29",X"26",X"27",X"28",X"A8",X"76",X"36",
		X"26",X"11",X"A4",X"40",X"3A",X"0D",X"40",X"A7",X"28",X"03",X"11",X"A7",X"40",X"DD",X"21",X"87",
		X"42",X"21",X"6F",X"13",X"3A",X"00",X"40",X"E6",X"02",X"20",X"03",X"21",X"7E",X"13",X"4E",X"06",
		X"00",X"23",X"1A",X"ED",X"B1",X"28",X"04",X"DD",X"70",X"00",X"C9",X"DD",X"7E",X"00",X"A7",X"C0",
		X"DD",X"36",X"00",X"FF",X"21",X"88",X"42",X"34",X"CD",X"14",X"0B",X"16",X"01",X"FF",X"C9",X"0E",
		X"03",X"10",X"17",X"24",X"31",X"38",X"45",X"52",X"59",X"66",X"73",X"80",X"87",X"94",X"0C",X"05",
		X"13",X"21",X"29",X"37",X"45",X"53",X"61",X"69",X"77",X"85",X"93",X"3A",X"5F",X"42",X"E6",X"01",
		X"C0",X"CD",X"AB",X"13",X"21",X"48",X"46",X"35",X"C0",X"3E",X"04",X"32",X"0A",X"40",X"CD",X"B6",
		X"13",X"CD",X"8D",X"14",X"CD",X"1E",X"11",X"CD",X"53",X"15",X"C9",X"06",X"1C",X"0E",X"03",X"CD",
		X"94",X"24",X"0C",X"10",X"FA",X"C9",X"DD",X"21",X"B0",X"45",X"3A",X"80",X"42",X"FE",X"03",X"38",
		X"02",X"3E",X"03",X"21",X"E4",X"13",X"E7",X"47",X"21",X"14",X"16",X"3A",X"80",X"42",X"E6",X"0F",
		X"87",X"5F",X"16",X"00",X"19",X"5E",X"23",X"56",X"EB",X"11",X"18",X"00",X"CD",X"E8",X"13",X"DD",
		X"19",X"10",X"F9",X"C9",X"04",X"04",X"05",X"06",X"7E",X"DD",X"77",X"06",X"23",X"7E",X"DD",X"77",
		X"05",X"23",X"7E",X"DD",X"77",X"04",X"23",X"7E",X"DD",X"77",X"03",X"23",X"DD",X"36",X"00",X"01",
		X"D9",X"21",X"57",X"34",X"3A",X"80",X"42",X"E6",X"01",X"20",X"03",X"21",X"13",X"34",X"DD",X"75",
		X"0C",X"DD",X"74",X"0D",X"DD",X"36",X"0E",X"00",X"CD",X"1B",X"32",X"D9",X"AF",X"DD",X"77",X"01",
		X"DD",X"77",X"02",X"C9",X"DD",X"21",X"C8",X"45",X"21",X"34",X"16",X"87",X"87",X"E7",X"CD",X"E8",
		X"13",X"CD",X"B9",X"2D",X"DD",X"36",X"09",X"20",X"DD",X"36",X"0A",X"E0",X"C9",X"7E",X"DD",X"77",
		X"06",X"23",X"7E",X"DD",X"77",X"05",X"23",X"7E",X"DD",X"77",X"04",X"23",X"7E",X"DD",X"77",X"03",
		X"23",X"DD",X"36",X"00",X"01",X"D9",X"21",X"2A",X"19",X"DD",X"75",X"0C",X"DD",X"74",X"0D",X"DD",
		X"36",X"0E",X"00",X"CD",X"1B",X"32",X"D9",X"AF",X"DD",X"77",X"01",X"DD",X"77",X"02",X"C9",X"DD",
		X"21",X"B0",X"45",X"21",X"B4",X"17",X"87",X"87",X"E7",X"CD",X"3D",X"14",X"C9",X"5A",X"4D",X"40",
		X"33",X"26",X"19",X"0C",X"0A",X"08",X"06",X"04",X"02",X"02",X"02",X"02",X"02",X"3A",X"80",X"42",
		X"FE",X"10",X"38",X"02",X"3E",X"0F",X"21",X"7D",X"14",X"E7",X"32",X"26",X"41",X"AF",X"32",X"81",
		X"41",X"3E",X"84",X"32",X"86",X"45",X"3E",X"EC",X"32",X"84",X"45",X"DD",X"21",X"80",X"45",X"3A",
		X"80",X"42",X"E6",X"01",X"21",X"D4",X"17",X"28",X"03",X"21",X"18",X"18",X"DD",X"75",X"0C",X"DD",
		X"74",X"0D",X"AF",X"DD",X"77",X"0E",X"CD",X"1B",X"32",X"3E",X"01",X"32",X"9A",X"45",X"32",X"99",
		X"45",X"3E",X"E4",X"32",X"AA",X"45",X"3E",X"EC",X"32",X"AB",X"45",X"3E",X"01",X"32",X"50",X"43",
		X"DD",X"21",X"98",X"45",X"3A",X"80",X"42",X"E6",X"01",X"21",X"89",X"18",X"28",X"03",X"21",X"CD",
		X"18",X"DD",X"75",X"0C",X"DD",X"74",X"0D",X"AF",X"DD",X"77",X"0E",X"CD",X"1B",X"32",X"C9",X"A7",
		X"C8",X"08",X"21",X"CC",X"17",X"3A",X"80",X"42",X"E6",X"01",X"28",X"03",X"21",X"10",X"18",X"08",
		X"1E",X"FF",X"0F",X"1C",X"30",X"FC",X"7B",X"DD",X"21",X"80",X"45",X"CD",X"2B",X"2C",X"DD",X"73",
		X"0C",X"DD",X"72",X"0D",X"AF",X"DD",X"77",X"0E",X"C9",X"A7",X"C8",X"08",X"21",X"54",X"18",X"3A",
		X"80",X"42",X"E6",X"01",X"28",X"03",X"21",X"98",X"18",X"08",X"1E",X"FF",X"0F",X"1C",X"30",X"FC",
		X"7B",X"DD",X"21",X"98",X"45",X"CD",X"2B",X"2C",X"DD",X"73",X"0C",X"DD",X"72",X"0D",X"AF",X"DD",
		X"77",X"0E",X"C9",X"3A",X"80",X"42",X"E6",X"07",X"21",X"59",X"19",X"CD",X"2B",X"2C",X"ED",X"53",
		X"12",X"41",X"3A",X"80",X"42",X"E6",X"01",X"C8",X"DD",X"21",X"60",X"4B",X"3E",X"07",X"32",X"44",
		X"43",X"AF",X"32",X"45",X"43",X"CD",X"97",X"15",X"DD",X"23",X"21",X"45",X"43",X"34",X"7E",X"FE",
		X"20",X"38",X"F2",X"36",X"00",X"01",X"40",X"FF",X"DD",X"09",X"3A",X"44",X"43",X"C6",X"05",X"32",
		X"44",X"43",X"FE",X"1E",X"38",X"DF",X"C9",X"CD",X"A1",X"15",X"3C",X"C8",X"3D",X"CD",X"ED",X"15",
		X"C9",X"CD",X"72",X"24",X"2A",X"12",X"41",X"3A",X"47",X"43",X"E7",X"3A",X"46",X"43",X"A6",X"EB",
		X"3E",X"FF",X"C8",X"21",X"C0",X"42",X"3A",X"47",X"43",X"E7",X"3A",X"46",X"43",X"4F",X"A6",X"3E",
		X"FF",X"C8",X"06",X"00",X"D5",X"FD",X"E1",X"79",X"FD",X"A6",X"FC",X"28",X"02",X"CB",X"D8",X"79",
		X"FD",X"A6",X"F8",X"28",X"02",X"CB",X"D0",X"79",X"FD",X"A6",X"F4",X"28",X"02",X"CB",X"C8",X"79",
		X"FD",X"A6",X"F0",X"28",X"02",X"CB",X"C0",X"78",X"21",X"04",X"16",X"E7",X"C9",X"ED",X"47",X"E6",
		X"F0",X"0F",X"0F",X"0F",X"0F",X"DD",X"77",X"00",X"ED",X"57",X"E6",X"0F",X"DD",X"77",X"E0",X"AF",
		X"DD",X"77",X"C0",X"C9",X"70",X"50",X"45",X"40",X"38",X"35",X"33",X"30",X"28",X"25",X"23",X"20",
		X"18",X"15",X"13",X"10",X"34",X"16",X"4C",X"16",X"64",X"16",X"7C",X"16",X"94",X"16",X"AC",X"16",
		X"C4",X"16",X"DC",X"16",X"F4",X"16",X"0C",X"17",X"24",X"17",X"3C",X"17",X"54",X"17",X"6C",X"17",
		X"84",X"17",X"9C",X"17",X"03",X"00",X"04",X"00",X"08",X"00",X"04",X"00",X"0D",X"00",X"04",X"00",
		X"12",X"00",X"04",X"00",X"17",X"00",X"04",X"00",X"1C",X"00",X"04",X"00",X"03",X"00",X"04",X"00",
		X"08",X"00",X"08",X"00",X"0D",X"00",X"0B",X"00",X"12",X"00",X"0E",X"00",X"17",X"00",X"10",X"00",
		X"03",X"00",X"0D",X"00",X"12",X"00",X"04",X"00",X"12",X"00",X"08",X"00",X"12",X"00",X"0B",X"00",
		X"12",X"00",X"11",X"00",X"12",X"00",X"17",X"00",X"03",X"00",X"10",X"00",X"03",X"00",X"04",X"00",
		X"08",X"00",X"04",X"00",X"0D",X"00",X"04",X"00",X"12",X"00",X"04",X"00",X"17",X"00",X"04",X"00",
		X"1C",X"00",X"04",X"00",X"03",X"00",X"04",X"00",X"08",X"00",X"04",X"00",X"0D",X"00",X"04",X"00",
		X"12",X"00",X"04",X"00",X"17",X"00",X"04",X"00",X"1C",X"00",X"04",X"00",X"03",X"00",X"04",X"00",
		X"08",X"00",X"04",X"00",X"0D",X"00",X"04",X"00",X"12",X"00",X"04",X"00",X"17",X"00",X"04",X"00",
		X"1C",X"00",X"04",X"00",X"03",X"00",X"04",X"00",X"08",X"00",X"04",X"00",X"0D",X"00",X"04",X"00",
		X"12",X"00",X"04",X"00",X"17",X"00",X"04",X"00",X"1C",X"00",X"04",X"00",X"03",X"00",X"04",X"00",
		X"08",X"00",X"04",X"00",X"0D",X"00",X"04",X"00",X"12",X"00",X"04",X"00",X"17",X"00",X"04",X"00",
		X"1C",X"00",X"04",X"00",X"03",X"00",X"04",X"00",X"08",X"00",X"04",X"00",X"0D",X"00",X"04",X"00",
		X"12",X"00",X"04",X"00",X"17",X"00",X"04",X"00",X"1C",X"00",X"04",X"00",X"03",X"00",X"04",X"00",
		X"08",X"00",X"04",X"00",X"0D",X"00",X"04",X"00",X"12",X"00",X"04",X"00",X"17",X"00",X"04",X"00",
		X"1C",X"00",X"04",X"00",X"03",X"00",X"04",X"00",X"08",X"00",X"04",X"00",X"0D",X"00",X"04",X"00",
		X"12",X"00",X"04",X"00",X"17",X"00",X"04",X"00",X"1C",X"00",X"04",X"00",X"03",X"00",X"04",X"00",
		X"08",X"00",X"04",X"00",X"0D",X"00",X"04",X"00",X"12",X"00",X"04",X"00",X"17",X"00",X"04",X"00",
		X"1C",X"00",X"04",X"00",X"03",X"00",X"04",X"00",X"08",X"00",X"04",X"00",X"0D",X"00",X"04",X"00",
		X"12",X"00",X"04",X"00",X"17",X"00",X"04",X"00",X"1C",X"00",X"04",X"00",X"03",X"00",X"04",X"00",
		X"08",X"00",X"04",X"00",X"0D",X"00",X"04",X"00",X"12",X"00",X"04",X"00",X"17",X"00",X"04",X"00",
		X"1C",X"00",X"04",X"00",X"03",X"00",X"04",X"00",X"08",X"00",X"04",X"00",X"0D",X"00",X"04",X"00",
		X"12",X"00",X"04",X"00",X"17",X"00",X"04",X"00",X"1C",X"00",X"04",X"00",X"03",X"00",X"04",X"00",
		X"08",X"00",X"04",X"00",X"0D",X"00",X"04",X"00",X"12",X"00",X"04",X"00",X"17",X"00",X"04",X"00",
		X"1C",X"00",X"04",X"00",X"03",X"00",X"1D",X"00",X"08",X"00",X"1D",X"00",X"0D",X"00",X"1D",X"00",
		X"12",X"00",X"1D",X"00",X"17",X"00",X"1D",X"00",X"1C",X"00",X"1D",X"00",X"01",X"18",X"F2",X"17",
		X"E3",X"17",X"D4",X"17",X"04",X"30",X"08",X"04",X"31",X"08",X"04",X"32",X"08",X"04",X"33",X"08",
		X"FF",X"D4",X"17",X"04",X"B0",X"08",X"04",X"B1",X"08",X"04",X"B2",X"08",X"04",X"B3",X"08",X"FF",
		X"E3",X"17",X"04",X"2E",X"08",X"04",X"2F",X"08",X"04",X"2E",X"08",X"04",X"2F",X"08",X"FF",X"F2",
		X"17",X"04",X"2E",X"08",X"04",X"2F",X"08",X"04",X"2E",X"08",X"04",X"2F",X"08",X"FF",X"01",X"18",
		X"45",X"18",X"36",X"18",X"27",X"18",X"18",X"18",X"07",X"F4",X"08",X"07",X"F5",X"08",X"07",X"F4",
		X"08",X"07",X"F5",X"08",X"FF",X"18",X"18",X"07",X"34",X"08",X"07",X"35",X"08",X"07",X"34",X"08",
		X"07",X"35",X"08",X"FF",X"27",X"18",X"07",X"E4",X"08",X"07",X"E5",X"08",X"07",X"E4",X"08",X"07",
		X"E5",X"08",X"FF",X"36",X"18",X"07",X"24",X"08",X"07",X"25",X"08",X"07",X"24",X"08",X"07",X"25",
		X"08",X"FF",X"45",X"18",X"89",X"18",X"7A",X"18",X"6B",X"18",X"5C",X"18",X"07",X"2A",X"08",X"07",
		X"2B",X"08",X"07",X"2C",X"08",X"07",X"2D",X"08",X"FF",X"5C",X"18",X"07",X"2A",X"08",X"07",X"2B",
		X"08",X"07",X"2C",X"08",X"07",X"2D",X"08",X"FF",X"6B",X"18",X"07",X"2A",X"08",X"07",X"2B",X"08",
		X"07",X"2C",X"08",X"07",X"2D",X"08",X"FF",X"7A",X"18",X"07",X"2A",X"08",X"07",X"2B",X"08",X"07",
		X"2C",X"08",X"07",X"2D",X"08",X"FF",X"89",X"18",X"CD",X"18",X"BE",X"18",X"AF",X"18",X"A0",X"18",
		X"07",X"22",X"08",X"07",X"23",X"08",X"07",X"22",X"08",X"07",X"23",X"08",X"FF",X"A0",X"18",X"07",
		X"22",X"08",X"07",X"23",X"08",X"07",X"22",X"08",X"07",X"23",X"08",X"FF",X"AF",X"18",X"07",X"22",
		X"08",X"07",X"23",X"08",X"07",X"22",X"08",X"07",X"23",X"08",X"FF",X"BE",X"18",X"07",X"22",X"08",
		X"07",X"23",X"08",X"07",X"22",X"08",X"07",X"23",X"08",X"FF",X"CD",X"18",X"11",X"09",X"19",X"3A",
		X"80",X"42",X"E6",X"01",X"28",X"03",X"11",X"15",X"19",X"DD",X"21",X"80",X"45",X"DD",X"73",X"0C",
		X"DD",X"72",X"0D",X"DD",X"36",X"0E",X"00",X"DD",X"36",X"11",X"35",X"3E",X"FF",X"32",X"4F",X"43",
		X"36",X"00",X"2C",X"36",X"01",X"2C",X"36",X"09",X"C9",X"04",X"39",X"10",X"04",X"3A",X"10",X"04",
		X"3B",X"20",X"FF",X"09",X"19",X"07",X"3D",X"07",X"07",X"3E",X"07",X"07",X"3F",X"07",X"07",X"7D",
		X"07",X"07",X"7E",X"07",X"07",X"7F",X"07",X"FF",X"15",X"19",X"05",X"21",X"08",X"05",X"21",X"08",
		X"05",X"21",X"08",X"05",X"21",X"08",X"FF",X"2A",X"19",X"52",X"01",X"4A",X"01",X"52",X"01",X"46",
		X"01",X"5A",X"01",X"42",X"01",X"66",X"01",X"4A",X"01",X"6E",X"1A",X"EE",X"19",X"6E",X"1A",X"EE",
		X"1A",X"6E",X"1B",X"EE",X"1B",X"6E",X"1C",X"EE",X"1C",X"6E",X"1E",X"EE",X"1D",X"6E",X"1E",X"EE",
		X"1E",X"6E",X"1F",X"EE",X"1F",X"6E",X"20",X"EE",X"20",X"20",X"48",X"70",X"98",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"FF",X"FF",X"FC",X"10",X"84",
		X"44",X"24",X"10",X"84",X"44",X"24",X"10",X"84",X"44",X"24",X"10",X"84",X"44",X"24",X"1F",X"FF",
		X"FF",X"FC",X"12",X"21",X"00",X"44",X"12",X"21",X"00",X"44",X"12",X"21",X"00",X"44",X"12",X"21",
		X"00",X"44",X"1F",X"FF",X"FF",X"FC",X"10",X"84",X"48",X"24",X"10",X"84",X"48",X"24",X"10",X"84",
		X"48",X"24",X"10",X"84",X"48",X"24",X"1F",X"FF",X"FF",X"FC",X"12",X"21",X"04",X"44",X"12",X"21",
		X"04",X"44",X"12",X"21",X"04",X"44",X"12",X"21",X"04",X"44",X"1F",X"FF",X"FF",X"FC",X"10",X"84",
		X"10",X"24",X"10",X"84",X"10",X"24",X"10",X"84",X"10",X"24",X"10",X"84",X"10",X"24",X"1F",X"FF",
		X"FF",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"FF",X"FF",X"FC",X"10",X"92",
		X"41",X"24",X"10",X"92",X"41",X"24",X"10",X"92",X"41",X"24",X"10",X"92",X"41",X"24",X"1F",X"FF",
		X"FF",X"FC",X"12",X"41",X"24",X"84",X"12",X"41",X"24",X"84",X"12",X"41",X"24",X"84",X"12",X"41",
		X"24",X"84",X"1F",X"FF",X"FF",X"FC",X"10",X"82",X"49",X"24",X"10",X"82",X"49",X"24",X"10",X"82",
		X"49",X"24",X"10",X"82",X"49",X"24",X"1F",X"FF",X"FF",X"FC",X"12",X"49",X"24",X"84",X"12",X"49",
		X"24",X"84",X"12",X"49",X"24",X"84",X"12",X"49",X"24",X"84",X"1F",X"FF",X"FF",X"FC",X"10",X"92",
		X"49",X"24",X"10",X"92",X"49",X"24",X"10",X"92",X"49",X"24",X"10",X"92",X"49",X"24",X"1F",X"FF",
		X"FF",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"FF",X"FF",X"FC",X"14",X"94",
		X"41",X"24",X"14",X"94",X"41",X"24",X"14",X"94",X"41",X"24",X"14",X"94",X"41",X"24",X"1F",X"FF",
		X"FF",X"FC",X"12",X"41",X"24",X"84",X"12",X"41",X"24",X"84",X"12",X"41",X"24",X"84",X"12",X"41",
		X"24",X"84",X"1F",X"FF",X"FF",X"FC",X"10",X"82",X"49",X"24",X"10",X"82",X"49",X"24",X"10",X"82",
		X"49",X"24",X"10",X"82",X"49",X"24",X"1F",X"FF",X"FF",X"FC",X"12",X"49",X"24",X"84",X"12",X"49",
		X"24",X"84",X"12",X"49",X"24",X"84",X"12",X"49",X"24",X"84",X"1F",X"FF",X"FF",X"FC",X"14",X"92",
		X"49",X"24",X"14",X"92",X"49",X"24",X"14",X"92",X"49",X"24",X"14",X"92",X"49",X"24",X"1F",X"FF",
		X"FF",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"FF",X"FF",X"FC",X"11",X"12",
		X"42",X"44",X"11",X"12",X"42",X"44",X"11",X"12",X"42",X"44",X"11",X"12",X"42",X"44",X"1F",X"FF",
		X"FF",X"FC",X"12",X"41",X"24",X"84",X"12",X"41",X"24",X"84",X"12",X"41",X"24",X"84",X"12",X"41",
		X"24",X"84",X"1F",X"FF",X"FF",X"FC",X"10",X"92",X"48",X"44",X"10",X"92",X"48",X"44",X"10",X"92",
		X"48",X"44",X"10",X"92",X"48",X"44",X"1F",X"FF",X"FF",X"FC",X"12",X"49",X"24",X"84",X"12",X"49",
		X"24",X"84",X"12",X"49",X"24",X"84",X"12",X"49",X"24",X"84",X"1F",X"FF",X"FF",X"FC",X"11",X"12",
		X"11",X"24",X"11",X"12",X"11",X"24",X"11",X"12",X"11",X"24",X"11",X"12",X"11",X"24",X"1F",X"FF",
		X"FF",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"FF",X"FF",X"FC",X"12",X"94",
		X"41",X"24",X"12",X"94",X"41",X"24",X"12",X"94",X"41",X"24",X"12",X"94",X"41",X"24",X"1F",X"FF",
		X"FF",X"FC",X"14",X"41",X"24",X"84",X"14",X"41",X"24",X"84",X"14",X"41",X"24",X"84",X"14",X"41",
		X"24",X"84",X"1F",X"FF",X"FF",X"FC",X"11",X"22",X"49",X"24",X"11",X"22",X"49",X"24",X"11",X"22",
		X"49",X"24",X"11",X"22",X"49",X"24",X"1F",X"FF",X"FF",X"FC",X"12",X"89",X"24",X"84",X"12",X"89",
		X"24",X"84",X"12",X"89",X"24",X"84",X"12",X"89",X"24",X"84",X"1F",X"FF",X"FF",X"FC",X"15",X"52",
		X"48",X"54",X"15",X"52",X"48",X"54",X"15",X"52",X"48",X"54",X"15",X"52",X"48",X"54",X"1F",X"FF",
		X"FF",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"FF",X"FF",X"FC",X"12",X"12",
		X"41",X"24",X"12",X"12",X"41",X"24",X"12",X"12",X"41",X"24",X"12",X"12",X"41",X"24",X"1F",X"FF",
		X"FF",X"FC",X"10",X"89",X"24",X"84",X"10",X"89",X"24",X"84",X"10",X"89",X"24",X"84",X"10",X"89",
		X"24",X"84",X"1F",X"FF",X"FF",X"FC",X"11",X"22",X"41",X"24",X"11",X"22",X"41",X"24",X"11",X"22",
		X"41",X"24",X"11",X"22",X"41",X"24",X"1F",X"FF",X"FF",X"FC",X"10",X"89",X"24",X"84",X"10",X"89",
		X"24",X"84",X"10",X"89",X"24",X"84",X"10",X"89",X"24",X"84",X"1F",X"FF",X"FF",X"FC",X"12",X"12",
		X"41",X"24",X"12",X"12",X"41",X"24",X"12",X"12",X"41",X"24",X"12",X"12",X"41",X"24",X"1F",X"FF",
		X"FF",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"FF",X"FF",X"FC",X"14",X"94",
		X"51",X"24",X"14",X"94",X"51",X"24",X"14",X"94",X"51",X"24",X"14",X"94",X"51",X"24",X"1F",X"FF",
		X"FF",X"FC",X"12",X"41",X"2A",X"94",X"12",X"41",X"2A",X"94",X"12",X"41",X"2A",X"94",X"12",X"41",
		X"2A",X"94",X"1F",X"FF",X"FF",X"FC",X"14",X"8A",X"41",X"24",X"14",X"8A",X"41",X"24",X"14",X"8A",
		X"41",X"24",X"14",X"8A",X"41",X"24",X"1F",X"FF",X"FF",X"FC",X"12",X"45",X"24",X"94",X"12",X"45",
		X"24",X"94",X"12",X"45",X"24",X"94",X"12",X"45",X"24",X"94",X"1F",X"FF",X"FF",X"FC",X"14",X"92",
		X"49",X"24",X"14",X"92",X"49",X"24",X"14",X"92",X"49",X"24",X"14",X"92",X"49",X"24",X"1F",X"FF",
		X"FF",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"FF",X"FF",X"FC",X"10",X"92",
		X"42",X"44",X"10",X"92",X"42",X"44",X"10",X"92",X"42",X"44",X"10",X"92",X"42",X"44",X"1F",X"FF",
		X"FF",X"FC",X"12",X"48",X"89",X"24",X"12",X"48",X"89",X"24",X"12",X"48",X"89",X"24",X"12",X"48",
		X"89",X"24",X"1F",X"FF",X"FF",X"FC",X"10",X"92",X"42",X"44",X"10",X"92",X"42",X"44",X"10",X"92",
		X"42",X"44",X"10",X"92",X"42",X"44",X"1F",X"FF",X"FF",X"FC",X"12",X"48",X"89",X"24",X"12",X"48",
		X"89",X"24",X"12",X"48",X"89",X"24",X"12",X"48",X"89",X"24",X"1F",X"FF",X"FF",X"FC",X"10",X"92",
		X"42",X"44",X"10",X"92",X"42",X"44",X"10",X"92",X"42",X"44",X"10",X"92",X"42",X"44",X"1F",X"FF",
		X"FF",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"08",X"88",X"48",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"42",
		X"01",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"08",X"90",X"48",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"42",X"09",X"08",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"08",X"20",X"48",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"24",X"80",X"48",X"00",X"04",
		X"00",X"08",X"00",X"24",X"00",X"48",X"00",X"00",X"84",X"48",X"02",X"24",X"84",X"48",X"00",X"80",
		X"01",X"10",X"04",X"84",X"09",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"49",X"00",X"04",X"84",
		X"49",X"10",X"00",X"00",X"02",X"48",X"00",X"08",X"12",X"08",X"00",X"00",X"00",X"48",X"00",X"00",
		X"92",X"48",X"02",X"08",X"92",X"48",X"00",X"82",X"01",X"10",X"04",X"90",X"08",X"10",X"00",X"10",
		X"01",X"10",X"00",X"02",X"49",X"00",X"04",X"92",X"49",X"10",X"02",X"20",X"80",X"48",X"00",X"24",
		X"10",X"08",X"00",X"24",X"02",X"48",X"00",X"00",X"92",X"48",X"02",X"24",X"92",X"48",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"28",X"82",X"48",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"82",
		X"49",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"04",X"92",X"48",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"92",X"49",X"08",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"24",X"92",X"48",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"24",X"80",X"88",X"00",X"04",
		X"00",X"08",X"00",X"24",X"08",X"08",X"00",X"00",X"80",X"88",X"02",X"24",X"88",X"88",X"00",X"80",
		X"01",X"00",X"04",X"80",X"09",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"49",X"00",X"04",X"84",
		X"49",X"10",X"00",X"00",X"00",X"08",X"00",X"20",X"10",X"08",X"02",X"00",X"00",X"00",X"00",X"00",
		X"91",X"08",X"02",X"24",X"91",X"08",X"00",X"82",X"01",X"10",X"04",X"90",X"08",X"10",X"00",X"10",
		X"01",X"10",X"00",X"02",X"49",X"00",X"04",X"92",X"49",X"10",X"02",X"20",X"00",X"48",X"00",X"24",
		X"40",X"08",X"00",X"24",X"02",X"48",X"00",X"00",X"02",X"48",X"02",X"24",X"42",X"48",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"28",X"82",X"48",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"82",
		X"49",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"44",X"92",X"48",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"12",X"49",X"08",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"A4",X"90",X"A8",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"20",X"80",X"48",X"04",X"00",
		X"00",X"08",X"00",X"20",X"00",X"48",X"00",X"04",X"84",X"48",X"04",X"24",X"84",X"48",X"02",X"12",
		X"09",X"10",X"00",X"10",X"48",X"10",X"00",X"10",X"01",X"10",X"00",X"02",X"49",X"00",X"02",X"12",
		X"49",X"10",X"00",X"00",X"04",X"48",X"02",X"40",X"84",X"08",X"00",X"40",X"00",X"48",X"00",X"04",
		X"80",X"48",X"02",X"44",X"84",X"48",X"02",X"12",X"09",X"10",X"00",X"10",X"48",X"10",X"00",X"10",
		X"01",X"10",X"00",X"02",X"49",X"00",X"02",X"12",X"49",X"10",X"04",X"20",X"80",X"48",X"04",X"00",
		X"00",X"08",X"00",X"20",X"00",X"48",X"00",X"04",X"84",X"48",X"04",X"24",X"84",X"48",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"28",X"A2",X"48",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"82",
		X"55",X"28",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"14",X"82",X"48",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"8A",X"49",X"28",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"24",X"92",X"48",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"24",X"80",X"80",X"00",X"04",
		X"08",X"00",X"00",X"24",X"00",X"88",X"00",X"00",X"88",X"88",X"02",X"24",X"88",X"88",X"00",X"80",
		X"10",X"08",X"04",X"90",X"00",X"48",X"00",X"10",X"02",X"48",X"00",X"01",X"12",X"48",X"04",X"91",
		X"12",X"48",X"00",X"24",X"08",X"08",X"00",X"24",X"00",X"08",X"00",X"04",X"00",X"80",X"00",X"00",
		X"88",X"88",X"02",X"24",X"88",X"88",X"00",X"82",X"10",X"08",X"04",X"90",X"00",X"48",X"00",X"10",
		X"02",X"48",X"00",X"01",X"12",X"48",X"04",X"91",X"12",X"48",X"02",X"24",X"80",X"80",X"00",X"04",
		X"08",X"00",X"00",X"24",X"00",X"88",X"00",X"00",X"88",X"88",X"02",X"24",X"88",X"88",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C4",X"21",
		X"D1",X"21",X"E5",X"21",X"F2",X"21",X"FF",X"21",X"0C",X"22",X"1B",X"22",X"2D",X"22",X"34",X"22",
		X"46",X"22",X"4C",X"22",X"53",X"22",X"5A",X"22",X"69",X"22",X"7B",X"22",X"7B",X"22",X"7B",X"22",
		X"7B",X"22",X"8C",X"22",X"A5",X"22",X"AA",X"22",X"AF",X"22",X"B4",X"22",X"C7",X"22",X"D3",X"22",
		X"E5",X"22",X"FA",X"22",X"0E",X"23",X"21",X"23",X"34",X"23",X"47",X"23",X"5A",X"23",X"6D",X"23",
		X"80",X"23",X"93",X"23",X"A6",X"23",X"B9",X"23",X"CC",X"23",X"E0",X"23",X"F1",X"23",X"02",X"24",
		X"0E",X"24",X"2A",X"24",X"96",X"4A",X"47",X"41",X"4D",X"45",X"40",X"40",X"4F",X"56",X"45",X"52",
		X"3F",X"EE",X"4A",X"50",X"55",X"53",X"48",X"40",X"53",X"54",X"41",X"52",X"54",X"40",X"42",X"55",
		X"54",X"54",X"4F",X"4E",X"3F",X"94",X"4A",X"50",X"4C",X"41",X"59",X"45",X"52",X"40",X"4F",X"4E",
		X"45",X"3F",X"94",X"4A",X"50",X"4C",X"41",X"59",X"45",X"52",X"40",X"54",X"57",X"4F",X"3F",X"80",
		X"4A",X"48",X"49",X"47",X"48",X"40",X"53",X"43",X"4F",X"52",X"45",X"3F",X"9F",X"4B",X"40",X"43",
		X"52",X"45",X"44",X"49",X"54",X"40",X"40",X"40",X"40",X"40",X"3F",X"9F",X"4B",X"40",X"40",X"46",
		X"52",X"45",X"45",X"40",X"50",X"4C",X"41",X"59",X"40",X"40",X"40",X"40",X"3F",X"5E",X"4B",X"46",
		X"55",X"45",X"4C",X"3F",X"CC",X"4A",X"43",X"4F",X"4E",X"47",X"52",X"41",X"54",X"55",X"4C",X"41",
		X"54",X"49",X"4F",X"4E",X"53",X"3F",X"6E",X"4B",X"59",X"4F",X"55",X"3F",X"9F",X"49",X"4A",X"55",
		X"4D",X"50",X"3F",X"26",X"4A",X"50",X"4C",X"41",X"59",X"3F",X"A9",X"4A",X"5B",X"40",X"40",X"41",
		X"4D",X"49",X"44",X"41",X"52",X"40",X"40",X"5B",X"3F",X"C7",X"4A",X"5B",X"40",X"40",X"43",X"48",
		X"41",X"52",X"41",X"43",X"54",X"45",X"52",X"40",X"40",X"5B",X"3F",X"BC",X"4A",X"3A",X"40",X"4B",
		X"4F",X"4E",X"41",X"4D",X"49",X"40",X"40",X"31",X"39",X"38",X"32",X"3F",X"54",X"4B",X"40",X"54",
		X"48",X"45",X"40",X"40",X"41",X"4D",X"49",X"44",X"41",X"52",X"40",X"40",X"53",X"59",X"53",X"54",
		X"45",X"4D",X"40",X"3B",X"3F",X"D5",X"4A",X"32",X"40",X"3F",X"D5",X"4A",X"33",X"40",X"3F",X"D5",
		X"4A",X"31",X"40",X"3F",X"75",X"4B",X"31",X"53",X"54",X"40",X"42",X"4F",X"4E",X"55",X"53",X"40",
		X"41",X"46",X"54",X"45",X"52",X"40",X"3F",X"75",X"49",X"35",X"30",X"30",X"30",X"30",X"40",X"50",
		X"54",X"53",X"3F",X"D1",X"4A",X"4F",X"4E",X"45",X"40",X"50",X"4C",X"41",X"59",X"45",X"52",X"40",
		X"4F",X"4E",X"4C",X"59",X"3F",X"F1",X"4A",X"4F",X"4E",X"45",X"40",X"4F",X"52",X"40",X"54",X"57",
		X"4F",X"40",X"50",X"4C",X"41",X"59",X"45",X"52",X"53",X"3F",X"04",X"4B",X"5B",X"40",X"53",X"43",
		X"4F",X"52",X"45",X"40",X"52",X"41",X"4E",X"4B",X"49",X"4E",X"47",X"40",X"5B",X"3F",X"27",X"4B",
		X"31",X"53",X"54",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"50",X"54",X"53",
		X"3F",X"29",X"4B",X"32",X"4E",X"44",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",
		X"50",X"54",X"53",X"3F",X"2B",X"4B",X"33",X"52",X"44",X"40",X"40",X"40",X"40",X"40",X"40",X"40",
		X"40",X"40",X"40",X"50",X"54",X"53",X"3F",X"2D",X"4B",X"34",X"54",X"48",X"40",X"40",X"40",X"40",
		X"40",X"40",X"40",X"40",X"40",X"40",X"50",X"54",X"53",X"3F",X"2F",X"4B",X"35",X"54",X"48",X"40",
		X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"50",X"54",X"53",X"3F",X"31",X"4B",X"36",
		X"54",X"48",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"50",X"54",X"53",X"3F",
		X"33",X"4B",X"37",X"54",X"48",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"50",
		X"54",X"53",X"3F",X"35",X"4B",X"38",X"54",X"48",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",
		X"40",X"40",X"50",X"54",X"53",X"3F",X"37",X"4B",X"39",X"54",X"48",X"40",X"40",X"40",X"40",X"40",
		X"40",X"40",X"40",X"40",X"40",X"50",X"54",X"53",X"3F",X"39",X"4B",X"31",X"30",X"54",X"48",X"40",
		X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"50",X"54",X"53",X"3F",X"F4",X"4A",X"50",X"55",
		X"53",X"48",X"40",X"4A",X"55",X"4D",X"50",X"40",X"40",X"42",X"55",X"54",X"54",X"4F",X"4E",X"3F",
		X"A8",X"4A",X"40",X"42",X"4F",X"4E",X"55",X"53",X"40",X"40",X"53",X"54",X"41",X"47",X"45",X"40",
		X"3F",X"6F",X"4A",X"3E",X"3E",X"3E",X"3E",X"40",X"35",X"30",X"30",X"30",X"40",X"50",X"54",X"53",
		X"40",X"3F",X"75",X"49",X"33",X"30",X"30",X"30",X"30",X"40",X"50",X"54",X"53",X"3F",X"78",X"4B",
		X"41",X"4E",X"44",X"40",X"42",X"4F",X"4E",X"55",X"53",X"40",X"45",X"56",X"45",X"52",X"59",X"40",
		X"37",X"30",X"30",X"30",X"30",X"40",X"50",X"54",X"53",X"3F",X"78",X"4B",X"41",X"4E",X"44",X"40",
		X"42",X"4F",X"4E",X"55",X"53",X"40",X"45",X"56",X"45",X"52",X"59",X"40",X"38",X"30",X"30",X"30",
		X"30",X"40",X"50",X"54",X"53",X"3F",X"3A",X"40",X"43",X"0F",X"0F",X"0F",X"E6",X"1F",X"67",X"32",
		X"44",X"43",X"3A",X"41",X"43",X"6F",X"0F",X"0F",X"0F",X"E6",X"1F",X"32",X"45",X"43",X"E6",X"07",
		X"D9",X"21",X"69",X"00",X"85",X"6F",X"7E",X"D9",X"32",X"46",X"43",X"29",X"29",X"7C",X"32",X"47",
		X"43",X"C9",X"3A",X"44",X"43",X"87",X"87",X"67",X"3A",X"45",X"43",X"6F",X"E6",X"07",X"D9",X"21",
		X"69",X"00",X"85",X"6F",X"7E",X"D9",X"32",X"46",X"43",X"7D",X"0F",X"0F",X"0F",X"E6",X"03",X"84",
		X"32",X"47",X"43",X"C9",X"3A",X"80",X"42",X"E6",X"01",X"CA",X"2A",X"25",X"C5",X"CD",X"A2",X"24",
		X"C1",X"C9",X"3A",X"48",X"46",X"32",X"44",X"43",X"79",X"E6",X"1F",X"32",X"45",X"43",X"CD",X"72",
		X"24",X"2A",X"BB",X"40",X"3A",X"47",X"43",X"E7",X"E5",X"DD",X"E1",X"21",X"C0",X"42",X"3A",X"47",
		X"43",X"E7",X"E5",X"FD",X"E1",X"06",X"00",X"3A",X"46",X"43",X"4F",X"DD",X"A6",X"00",X"28",X"02",
		X"CB",X"F0",X"79",X"FD",X"A6",X"00",X"28",X"02",X"CB",X"D0",X"79",X"DD",X"A6",X"04",X"28",X"02",
		X"CB",X"E0",X"79",X"FD",X"A6",X"04",X"28",X"02",X"CB",X"C0",X"79",X"07",X"4F",X"30",X"04",X"DD",
		X"2B",X"FD",X"2B",X"DD",X"A6",X"00",X"28",X"02",X"CB",X"E8",X"79",X"FD",X"A6",X"00",X"28",X"02",
		X"CB",X"C8",X"79",X"FD",X"A6",X"04",X"28",X"02",X"CB",X"D8",X"21",X"22",X"3B",X"78",X"E7",X"47",
		X"3A",X"44",X"43",X"2F",X"E6",X"1F",X"87",X"87",X"87",X"6F",X"26",X"00",X"29",X"29",X"3A",X"45",
		X"43",X"85",X"6F",X"78",X"01",X"00",X"48",X"09",X"77",X"C9",X"C5",X"CD",X"30",X"25",X"C1",X"C9",
		X"3A",X"48",X"46",X"32",X"44",X"43",X"79",X"E6",X"1F",X"32",X"45",X"43",X"CD",X"72",X"24",X"2A",
		X"BB",X"40",X"3A",X"47",X"43",X"E7",X"E5",X"DD",X"E1",X"21",X"C0",X"42",X"3A",X"47",X"43",X"E7",
		X"E5",X"FD",X"E1",X"06",X"00",X"3A",X"46",X"43",X"4F",X"DD",X"A6",X"00",X"28",X"02",X"CB",X"F0",
		X"79",X"FD",X"A6",X"00",X"28",X"02",X"CB",X"D0",X"79",X"DD",X"A6",X"04",X"28",X"02",X"CB",X"E0",
		X"79",X"FD",X"A6",X"04",X"28",X"02",X"CB",X"C0",X"79",X"07",X"4F",X"30",X"04",X"DD",X"2B",X"FD",
		X"2B",X"DD",X"A6",X"00",X"28",X"02",X"CB",X"E8",X"79",X"FD",X"A6",X"00",X"28",X"02",X"CB",X"C8",
		X"79",X"DD",X"A6",X"04",X"28",X"02",X"CB",X"F8",X"79",X"FD",X"A6",X"04",X"28",X"02",X"CB",X"D8",
		X"78",X"21",X"22",X"3A",X"E7",X"47",X"3A",X"44",X"43",X"2F",X"E6",X"1F",X"87",X"87",X"87",X"6F",
		X"26",X"00",X"29",X"29",X"3A",X"45",X"43",X"85",X"6F",X"78",X"01",X"00",X"48",X"09",X"77",X"C9",
		X"21",X"33",X"3F",X"E5",X"3A",X"4F",X"43",X"A7",X"C2",X"94",X"26",X"3A",X"06",X"40",X"A7",X"CA",
		X"AE",X"3D",X"AF",X"32",X"53",X"43",X"CD",X"36",X"2C",X"CA",X"9C",X"26",X"3A",X"4A",X"43",X"4F",
		X"E6",X"03",X"20",X"46",X"AF",X"32",X"53",X"43",X"3A",X"86",X"45",X"E6",X"07",X"FE",X"04",X"20",
		X"03",X"32",X"53",X"43",X"78",X"B9",X"28",X"20",X"78",X"B1",X"FE",X"0C",X"28",X"1A",X"3A",X"53",
		X"43",X"A7",X"20",X"1D",X"78",X"CD",X"E4",X"26",X"28",X"04",X"3E",X"04",X"18",X"57",X"78",X"CD",
		X"0A",X"27",X"28",X"4A",X"3E",X"08",X"18",X"4D",X"3A",X"53",X"43",X"A7",X"20",X"03",X"78",X"18",
		X"44",X"78",X"CD",X"C8",X"26",X"28",X"37",X"78",X"18",X"3B",X"AF",X"32",X"53",X"43",X"3A",X"84",
		X"45",X"E6",X"07",X"FE",X"04",X"20",X"03",X"32",X"53",X"43",X"78",X"B9",X"28",X"DA",X"78",X"B1",
		X"FE",X"03",X"28",X"D4",X"3A",X"53",X"43",X"A7",X"20",X"D7",X"78",X"CD",X"2E",X"27",X"28",X"04",
		X"3E",X"02",X"18",X"11",X"78",X"CD",X"54",X"27",X"28",X"04",X"3E",X"01",X"18",X"07",X"79",X"CD",
		X"C8",X"26",X"28",X"38",X"79",X"5F",X"21",X"4A",X"43",X"BE",X"D9",X"C4",X"FF",X"14",X"D9",X"7E",
		X"A7",X"20",X"01",X"7B",X"32",X"54",X"43",X"73",X"7B",X"CD",X"A0",X"26",X"E5",X"D5",X"C5",X"CD",
		X"C4",X"3B",X"C1",X"D1",X"E1",X"3A",X"40",X"43",X"32",X"86",X"45",X"3A",X"41",X"43",X"32",X"84",
		X"45",X"CD",X"5D",X"28",X"DD",X"21",X"80",X"45",X"CD",X"1B",X"32",X"C9",X"CD",X"C4",X"3B",X"C9",
		X"CD",X"76",X"2C",X"3A",X"86",X"45",X"5F",X"3A",X"4B",X"43",X"83",X"32",X"40",X"43",X"3A",X"84",
		X"45",X"5F",X"3A",X"4C",X"43",X"83",X"32",X"41",X"43",X"CD",X"46",X"24",X"2A",X"BB",X"40",X"3A",
		X"47",X"43",X"E7",X"3A",X"46",X"43",X"A6",X"C9",X"CD",X"A6",X"2C",X"3A",X"86",X"45",X"5F",X"3A",
		X"4B",X"43",X"83",X"32",X"40",X"43",X"3A",X"84",X"45",X"5F",X"3A",X"4C",X"43",X"83",X"32",X"41",
		X"43",X"C3",X"B9",X"26",X"CD",X"A6",X"2C",X"3A",X"86",X"45",X"E6",X"FC",X"C6",X"04",X"CB",X"57",
		X"20",X"02",X"C6",X"04",X"5F",X"3A",X"4B",X"43",X"83",X"32",X"40",X"43",X"3A",X"84",X"45",X"5F",
		X"3A",X"4C",X"43",X"83",X"32",X"41",X"43",X"C3",X"B9",X"26",X"CD",X"A6",X"2C",X"3A",X"86",X"45",
		X"E6",X"FC",X"CB",X"57",X"20",X"02",X"D6",X"04",X"5F",X"3A",X"4B",X"43",X"83",X"32",X"40",X"43",
		X"3A",X"84",X"45",X"5F",X"3A",X"4C",X"43",X"83",X"32",X"41",X"43",X"C3",X"B9",X"26",X"CD",X"A6",
		X"2C",X"3A",X"86",X"45",X"5F",X"3A",X"4B",X"43",X"83",X"32",X"40",X"43",X"3A",X"84",X"45",X"E6",
		X"FC",X"C6",X"04",X"CB",X"57",X"20",X"02",X"C6",X"04",X"5F",X"3A",X"4C",X"43",X"83",X"32",X"41",
		X"43",X"C3",X"B9",X"26",X"CD",X"A6",X"2C",X"3A",X"86",X"45",X"5F",X"3A",X"4B",X"43",X"83",X"32",
		X"40",X"43",X"3A",X"84",X"45",X"E6",X"FC",X"CB",X"57",X"20",X"02",X"D6",X"04",X"5F",X"3A",X"4C",
		X"43",X"83",X"32",X"41",X"43",X"C3",X"B9",X"26",X"3A",X"52",X"43",X"3C",X"C0",X"3A",X"53",X"43",
		X"A7",X"C8",X"3A",X"86",X"45",X"32",X"40",X"43",X"3A",X"84",X"45",X"32",X"41",X"43",X"CD",X"46",
		X"24",X"21",X"C0",X"42",X"3A",X"47",X"43",X"E7",X"3A",X"46",X"43",X"A6",X"C8",X"2F",X"A6",X"77",
		X"CD",X"AE",X"24",X"21",X"45",X"43",X"34",X"CD",X"AE",X"24",X"21",X"45",X"43",X"35",X"2B",X"35",
		X"CD",X"AE",X"24",X"2A",X"81",X"42",X"7C",X"B5",X"C8",X"2B",X"22",X"81",X"42",X"11",X"01",X"03",
		X"FF",X"CD",X"F8",X"0A",X"C9",X"3A",X"53",X"43",X"A7",X"C8",X"3A",X"86",X"45",X"32",X"40",X"43",
		X"3A",X"84",X"45",X"32",X"41",X"43",X"CD",X"46",X"24",X"21",X"C0",X"42",X"3A",X"47",X"43",X"E7",
		X"3A",X"46",X"43",X"A6",X"C8",X"2F",X"A6",X"77",X"CD",X"3C",X"25",X"21",X"45",X"43",X"34",X"CD",
		X"3C",X"25",X"21",X"45",X"43",X"35",X"2B",X"35",X"CD",X"3C",X"25",X"2A",X"81",X"42",X"7C",X"B5",
		X"C8",X"2B",X"22",X"81",X"42",X"11",X"01",X"03",X"FF",X"CD",X"F8",X"0A",X"C9",X"3A",X"CE",X"45",
		X"32",X"44",X"43",X"3A",X"CC",X"45",X"32",X"45",X"43",X"CD",X"72",X"24",X"21",X"C0",X"42",X"3A",
		X"47",X"43",X"E7",X"3A",X"46",X"43",X"A6",X"C8",X"2F",X"A6",X"77",X"CD",X"3F",X"28",X"21",X"45",
		X"43",X"34",X"CD",X"3F",X"28",X"21",X"45",X"43",X"35",X"2B",X"35",X"CD",X"3F",X"28",X"C9",X"3A",
		X"06",X"40",X"A7",X"28",X"0C",X"3A",X"45",X"43",X"FE",X"05",X"D8",X"FE",X"1D",X"D0",X"C3",X"AE",
		X"24",X"3A",X"45",X"43",X"FE",X"0C",X"D8",X"FE",X"1A",X"D0",X"C3",X"AE",X"24",X"3A",X"80",X"42",
		X"E6",X"01",X"CA",X"C5",X"27",X"21",X"78",X"27",X"E5",X"3A",X"53",X"43",X"A7",X"C8",X"21",X"C0",
		X"42",X"3A",X"47",X"43",X"CD",X"24",X"2C",X"3A",X"46",X"43",X"A6",X"28",X"62",X"3A",X"52",X"43",
		X"FE",X"01",X"38",X"6A",X"C8",X"CD",X"BD",X"29",X"21",X"41",X"44",X"7E",X"23",X"BE",X"38",X"01",
		X"77",X"CD",X"2D",X"2A",X"21",X"41",X"45",X"7E",X"23",X"BE",X"38",X"01",X"77",X"3A",X"40",X"44",
		X"3C",X"C0",X"3A",X"40",X"45",X"3C",X"C0",X"3A",X"80",X"42",X"E6",X"01",X"C8",X"3A",X"42",X"44",
		X"21",X"42",X"45",X"BE",X"30",X"11",X"CD",X"9D",X"29",X"3A",X"42",X"45",X"2A",X"81",X"42",X"CD",
		X"24",X"2C",X"22",X"81",X"42",X"18",X"0F",X"CD",X"7D",X"29",X"3A",X"42",X"44",X"2A",X"81",X"42",
		X"CD",X"24",X"2C",X"22",X"81",X"42",X"3E",X"01",X"32",X"52",X"43",X"CD",X"CB",X"11",X"C9",X"3A",
		X"52",X"43",X"FE",X"01",X"D8",X"28",X"02",X"18",X"9C",X"AF",X"32",X"52",X"43",X"C9",X"3A",X"54",
		X"43",X"A7",X"C8",X"06",X"FF",X"04",X"0F",X"30",X"FC",X"78",X"E6",X"03",X"21",X"2D",X"29",X"CD",
		X"2B",X"2C",X"EB",X"22",X"60",X"43",X"23",X"23",X"23",X"23",X"23",X"22",X"62",X"43",X"CD",X"CB",
		X"11",X"CD",X"9D",X"2A",X"CD",X"23",X"2B",X"3E",X"FF",X"32",X"52",X"43",X"3A",X"40",X"44",X"FE",
		X"01",X"CA",X"1F",X"2A",X"3A",X"40",X"45",X"FE",X"01",X"CA",X"8F",X"2A",X"C9",X"49",X"29",X"53",
		X"29",X"3F",X"29",X"35",X"29",X"08",X"02",X"04",X"01",X"08",X"08",X"01",X"04",X"02",X"08",X"04",
		X"01",X"08",X"02",X"04",X"04",X"02",X"08",X"01",X"04",X"01",X"08",X"02",X"04",X"01",X"01",X"04",
		X"02",X"08",X"01",X"02",X"04",X"01",X"08",X"02",X"02",X"08",X"01",X"04",X"02",X"21",X"C0",X"42",
		X"3A",X"47",X"43",X"E7",X"3A",X"46",X"43",X"B6",X"77",X"CD",X"AE",X"24",X"21",X"45",X"43",X"34",
		X"CD",X"AE",X"24",X"21",X"45",X"43",X"35",X"2B",X"35",X"CD",X"AE",X"24",X"C9",X"21",X"42",X"44",
		X"7E",X"A7",X"C8",X"47",X"23",X"23",X"C5",X"7E",X"32",X"40",X"43",X"23",X"7E",X"32",X"41",X"43",
		X"23",X"E5",X"CD",X"46",X"24",X"CD",X"5D",X"29",X"E1",X"C1",X"10",X"EA",X"C9",X"21",X"42",X"45",
		X"7E",X"A7",X"C8",X"47",X"23",X"23",X"C5",X"7E",X"32",X"40",X"43",X"23",X"7E",X"32",X"41",X"43",
		X"23",X"E5",X"CD",X"46",X"24",X"CD",X"5D",X"29",X"E1",X"C1",X"10",X"EA",X"C9",X"21",X"40",X"44",
		X"7E",X"A7",X"C8",X"3C",X"C8",X"23",X"34",X"7E",X"3C",X"CD",X"23",X"2C",X"3A",X"84",X"45",X"E6",
		X"F8",X"BE",X"2B",X"20",X"11",X"3A",X"86",X"45",X"E6",X"F8",X"BE",X"20",X"09",X"21",X"40",X"44",
		X"7E",X"23",X"BE",X"C0",X"18",X"39",X"3A",X"41",X"44",X"3D",X"32",X"41",X"44",X"2B",X"3A",X"84",
		X"45",X"E6",X"F8",X"BE",X"2B",X"20",X"07",X"3A",X"86",X"45",X"E6",X"F8",X"BE",X"C8",X"3A",X"41",
		X"44",X"D6",X"01",X"38",X"14",X"32",X"41",X"44",X"2B",X"3A",X"84",X"45",X"E6",X"F8",X"BE",X"2B",
		X"20",X"07",X"3A",X"86",X"45",X"E6",X"F8",X"BE",X"C8",X"21",X"40",X"44",X"36",X"FF",X"C9",X"CD",
		X"CB",X"11",X"CD",X"5D",X"28",X"AF",X"32",X"52",X"43",X"CD",X"2C",X"0B",X"C9",X"21",X"40",X"45",
		X"7E",X"A7",X"C8",X"3C",X"C8",X"23",X"34",X"7E",X"3C",X"CD",X"23",X"2C",X"3A",X"84",X"45",X"E6",
		X"F8",X"BE",X"2B",X"20",X"11",X"3A",X"86",X"45",X"E6",X"F8",X"BE",X"20",X"09",X"21",X"40",X"45",
		X"7E",X"23",X"BE",X"C0",X"18",X"39",X"3A",X"41",X"45",X"3D",X"32",X"41",X"45",X"2B",X"3A",X"84",
		X"45",X"E6",X"F8",X"BE",X"2B",X"20",X"07",X"3A",X"86",X"45",X"E6",X"F8",X"BE",X"C8",X"3A",X"41",
		X"45",X"D6",X"01",X"38",X"14",X"32",X"41",X"45",X"2B",X"3A",X"84",X"45",X"E6",X"F8",X"BE",X"2B",
		X"20",X"07",X"3A",X"86",X"45",X"E6",X"F8",X"BE",X"C8",X"21",X"40",X"45",X"36",X"FF",X"C9",X"CD",
		X"CB",X"11",X"CD",X"5D",X"28",X"AF",X"32",X"52",X"43",X"CD",X"2C",X"0B",X"C9",X"3A",X"86",X"45",
		X"E6",X"F8",X"32",X"64",X"43",X"3A",X"84",X"45",X"E6",X"F8",X"32",X"65",X"43",X"DD",X"2A",X"60",
		X"43",X"01",X"00",X"00",X"DD",X"7E",X"00",X"CD",X"D6",X"2C",X"DD",X"7E",X"01",X"CD",X"E6",X"2C",
		X"21",X"44",X"44",X"22",X"68",X"43",X"2A",X"68",X"43",X"0C",X"3A",X"64",X"43",X"77",X"23",X"3A",
		X"65",X"43",X"77",X"23",X"22",X"68",X"43",X"CD",X"E6",X"2B",X"20",X"1E",X"CD",X"A9",X"2B",X"28",
		X"2B",X"04",X"78",X"FE",X"08",X"30",X"25",X"2A",X"40",X"43",X"22",X"64",X"43",X"21",X"C0",X"42",
		X"7A",X"CD",X"24",X"2C",X"7B",X"A6",X"28",X"20",X"18",X"CC",X"06",X"00",X"DD",X"23",X"2A",X"6A",
		X"43",X"22",X"4B",X"43",X"DD",X"7E",X"01",X"CD",X"E6",X"2C",X"18",X"DB",X"21",X"40",X"44",X"36",
		X"FF",X"23",X"36",X"00",X"23",X"36",X"00",X"C9",X"21",X"40",X"44",X"71",X"23",X"36",X"01",X"23",
		X"36",X"01",X"C9",X"3A",X"86",X"45",X"E6",X"F8",X"32",X"64",X"43",X"3A",X"84",X"45",X"E6",X"F8",
		X"32",X"65",X"43",X"DD",X"2A",X"62",X"43",X"01",X"00",X"00",X"DD",X"7E",X"00",X"CD",X"D6",X"2C",
		X"DD",X"7E",X"01",X"CD",X"E6",X"2C",X"21",X"44",X"45",X"22",X"68",X"43",X"2A",X"68",X"43",X"0C",
		X"3A",X"64",X"43",X"77",X"23",X"3A",X"65",X"43",X"77",X"23",X"22",X"68",X"43",X"CD",X"E6",X"2B",
		X"20",X"1E",X"CD",X"A9",X"2B",X"28",X"2B",X"04",X"78",X"FE",X"08",X"30",X"25",X"2A",X"40",X"43",
		X"22",X"64",X"43",X"21",X"C0",X"42",X"7A",X"CD",X"24",X"2C",X"7B",X"A6",X"28",X"20",X"18",X"CC",
		X"06",X"00",X"DD",X"23",X"2A",X"6A",X"43",X"22",X"4B",X"43",X"DD",X"7E",X"01",X"CD",X"E6",X"2C",
		X"18",X"DB",X"21",X"40",X"45",X"36",X"FF",X"23",X"36",X"00",X"23",X"36",X"00",X"C9",X"21",X"40",
		X"45",X"71",X"23",X"36",X"01",X"23",X"36",X"01",X"C9",X"3A",X"65",X"43",X"57",X"3A",X"4C",X"43",
		X"82",X"57",X"32",X"41",X"43",X"3A",X"64",X"43",X"5F",X"3A",X"4B",X"43",X"83",X"32",X"40",X"43",
		X"0F",X"0F",X"0F",X"E6",X"1F",X"67",X"7A",X"6F",X"0F",X"0F",X"0F",X"E6",X"07",X"D9",X"21",X"69",
		X"00",X"85",X"6F",X"7E",X"D9",X"5F",X"29",X"29",X"7C",X"57",X"2A",X"BB",X"40",X"85",X"6F",X"3E",
		X"00",X"8C",X"67",X"7B",X"A6",X"C9",X"3A",X"65",X"43",X"57",X"3A",X"6B",X"43",X"82",X"57",X"32",
		X"41",X"43",X"3A",X"64",X"43",X"5F",X"3A",X"6A",X"43",X"83",X"32",X"40",X"43",X"0F",X"0F",X"0F",
		X"E6",X"1F",X"67",X"7A",X"6F",X"0F",X"0F",X"0F",X"E6",X"07",X"D9",X"21",X"69",X"00",X"85",X"6F",
		X"7E",X"D9",X"5F",X"29",X"29",X"7C",X"57",X"2A",X"BB",X"40",X"85",X"6F",X"3E",X"00",X"8C",X"67",
		X"7B",X"A6",X"C9",X"87",X"85",X"6F",X"3E",X"00",X"8C",X"67",X"C9",X"87",X"85",X"6F",X"3E",X"00",
		X"8C",X"67",X"5E",X"23",X"56",X"C9",X"3A",X"1E",X"40",X"A7",X"20",X"22",X"3A",X"10",X"40",X"0F",
		X"0F",X"0F",X"0F",X"E6",X"03",X"47",X"3A",X"12",X"40",X"07",X"07",X"CB",X"10",X"07",X"07",X"CB",
		X"10",X"78",X"E6",X"0C",X"20",X"03",X"78",X"E6",X"03",X"47",X"32",X"48",X"43",X"C9",X"3A",X"11",
		X"40",X"0F",X"0F",X"0F",X"0F",X"E6",X"03",X"47",X"3A",X"12",X"40",X"0F",X"CB",X"10",X"3A",X"10",
		X"40",X"0F",X"CB",X"10",X"18",X"DB",X"21",X"86",X"2C",X"CD",X"23",X"2C",X"7E",X"32",X"4B",X"43",
		X"23",X"7E",X"32",X"4C",X"43",X"C9",X"00",X"00",X"00",X"FF",X"00",X"01",X"00",X"00",X"01",X"00",
		X"01",X"FF",X"01",X"01",X"00",X"00",X"FF",X"00",X"FF",X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"21",X"B6",X"2C",X"CD",X"23",X"2C",X"7E",X"32",X"4B",X"43",
		X"23",X"7E",X"32",X"4C",X"43",X"C9",X"00",X"00",X"00",X"FB",X"00",X"05",X"00",X"00",X"05",X"00",
		X"05",X"FB",X"05",X"05",X"00",X"00",X"FB",X"00",X"FB",X"FB",X"FB",X"05",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"21",X"F6",X"2C",X"CD",X"23",X"2C",X"7E",X"32",X"4B",X"43",
		X"23",X"7E",X"32",X"4C",X"43",X"C9",X"21",X"F6",X"2C",X"CD",X"23",X"2C",X"7E",X"32",X"6A",X"43",
		X"23",X"7E",X"32",X"6B",X"43",X"C9",X"00",X"00",X"00",X"F8",X"00",X"08",X"00",X"00",X"08",X"00",
		X"08",X"F8",X"08",X"08",X"00",X"00",X"F8",X"00",X"F8",X"F8",X"F8",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"3A",X"F1",X"41",X"A7",X"C0",X"06",X"07",X"DD",X"21",X"64",
		X"40",X"3A",X"60",X"40",X"6F",X"3A",X"63",X"40",X"67",X"DD",X"7E",X"00",X"95",X"30",X"02",X"ED",
		X"44",X"FE",X"07",X"30",X"3D",X"DD",X"7E",X"03",X"94",X"30",X"02",X"ED",X"44",X"FE",X"07",X"30",
		X"31",X"48",X"3E",X"08",X"90",X"47",X"21",X"82",X"45",X"11",X"18",X"00",X"19",X"10",X"FD",X"41",
		X"4F",X"7E",X"FE",X"01",X"20",X"1C",X"3A",X"F5",X"41",X"A7",X"20",X"0F",X"2B",X"2B",X"CD",X"DC",
		X"18",X"CD",X"A0",X"0B",X"CD",X"0C",X"0B",X"CD",X"A7",X"28",X"C9",X"79",X"32",X"F4",X"41",X"CD",
		X"10",X"0B",X"11",X"04",X"00",X"DD",X"19",X"10",X"A8",X"C9",X"DD",X"21",X"98",X"45",X"11",X"18",
		X"00",X"06",X"07",X"D9",X"CD",X"93",X"2D",X"D9",X"DD",X"19",X"10",X"F7",X"CD",X"51",X"32",X"CD",
		X"55",X"33",X"C9",X"DD",X"7E",X"00",X"DD",X"B6",X"01",X"0F",X"D0",X"DD",X"7E",X"02",X"E6",X"1F",
		X"EF",X"E0",X"2D",X"F9",X"2D",X"30",X"30",X"31",X"30",X"6D",X"30",X"25",X"31",X"26",X"31",X"7A",
		X"31",X"8F",X"31",X"8F",X"31",X"AD",X"31",X"E9",X"31",X"21",X"CD",X"33",X"3A",X"80",X"42",X"FE",
		X"10",X"38",X"02",X"3E",X"10",X"85",X"30",X"01",X"24",X"6F",X"7E",X"DD",X"77",X"09",X"ED",X"44",
		X"DD",X"77",X"0A",X"AF",X"DD",X"77",X"0E",X"DD",X"77",X"0B",X"3E",X"03",X"DD",X"77",X"07",X"C9",
		X"21",X"57",X"34",X"3A",X"80",X"42",X"E6",X"01",X"20",X"03",X"21",X"13",X"34",X"DD",X"75",X"0C",
		X"DD",X"74",X"0D",X"CD",X"B9",X"2D",X"DD",X"34",X"02",X"DD",X"CB",X"01",X"46",X"C0",X"CD",X"1B",
		X"32",X"CD",X"EA",X"31",X"DD",X"7E",X"07",X"EF",X"10",X"2E",X"3C",X"2E",X"71",X"2E",X"A4",X"2E",
		X"DD",X"7E",X"05",X"DD",X"86",X"09",X"30",X"03",X"DD",X"34",X"06",X"DD",X"77",X"05",X"47",X"DD",
		X"7E",X"0B",X"A7",X"28",X"04",X"DD",X"35",X"0B",X"C9",X"78",X"E6",X"E0",X"28",X"03",X"FE",X"20",
		X"C0",X"DD",X"36",X"0B",X"03",X"CD",X"BE",X"34",X"CD",X"C3",X"2F",X"C9",X"DD",X"7E",X"0A",X"ED",
		X"44",X"47",X"DD",X"7E",X"03",X"B8",X"30",X"03",X"DD",X"35",X"04",X"DD",X"86",X"0A",X"DD",X"77",
		X"03",X"47",X"DD",X"7E",X"0B",X"A7",X"28",X"04",X"DD",X"35",X"0B",X"C9",X"78",X"E6",X"E0",X"FE",
		X"C0",X"28",X"03",X"FE",X"E0",X"C0",X"DD",X"36",X"0B",X"03",X"CD",X"BE",X"34",X"CD",X"82",X"2F",
		X"C9",X"DD",X"7E",X"0A",X"ED",X"44",X"47",X"DD",X"7E",X"05",X"B8",X"30",X"03",X"DD",X"35",X"06",
		X"DD",X"86",X"0A",X"DD",X"77",X"05",X"47",X"DD",X"7E",X"0B",X"A7",X"28",X"04",X"DD",X"35",X"0B",
		X"C9",X"78",X"E6",X"E0",X"28",X"03",X"FE",X"20",X"C0",X"DD",X"36",X"0B",X"03",X"CD",X"BE",X"34",
		X"CD",X"FC",X"2F",X"C9",X"DD",X"7E",X"03",X"DD",X"86",X"09",X"30",X"03",X"DD",X"34",X"04",X"DD",
		X"77",X"03",X"47",X"DD",X"7E",X"0B",X"A7",X"28",X"04",X"DD",X"35",X"0B",X"C9",X"78",X"E6",X"E0",
		X"FE",X"C0",X"28",X"03",X"FE",X"E0",X"C0",X"DD",X"36",X"0B",X"03",X"CD",X"BE",X"34",X"CD",X"D2",
		X"2E",X"C9",X"78",X"21",X"66",X"34",X"85",X"6F",X"30",X"01",X"24",X"7E",X"A7",X"C8",X"3D",X"21",
		X"11",X"2F",X"E5",X"EF",X"EE",X"2E",X"F2",X"2E",X"F7",X"2E",X"FB",X"2E",X"FF",X"2E",X"AF",X"06",
		X"03",X"C9",X"3E",X"02",X"06",X"03",X"C9",X"3E",X"02",X"47",X"C9",X"AF",X"06",X"02",X"C9",X"DD",
		X"36",X"12",X"01",X"DD",X"CB",X"06",X"46",X"28",X"04",X"3E",X"02",X"47",X"C9",X"AF",X"06",X"02",
		X"C9",X"DD",X"77",X"07",X"DD",X"70",X"08",X"C9",X"4F",X"DD",X"CB",X"01",X"46",X"20",X"1C",X"21",
		X"22",X"34",X"3A",X"80",X"42",X"E6",X"01",X"20",X"03",X"21",X"DE",X"33",X"79",X"CD",X"2B",X"2C",
		X"DD",X"73",X"0C",X"DD",X"72",X"0D",X"DD",X"36",X"0E",X"00",X"C9",X"21",X"6B",X"18",X"3A",X"80",
		X"42",X"E6",X"01",X"28",X"03",X"21",X"AF",X"18",X"DD",X"75",X"0C",X"DD",X"74",X"0D",X"DD",X"36",
		X"0E",X"00",X"DD",X"6E",X"03",X"DD",X"66",X"04",X"29",X"29",X"29",X"7C",X"D6",X"02",X"32",X"AB",
		X"45",X"DD",X"6E",X"05",X"DD",X"66",X"06",X"29",X"29",X"29",X"7C",X"C6",X"03",X"32",X"AA",X"45",
		X"21",X"AB",X"45",X"7E",X"FE",X"EC",X"D8",X"36",X"EC",X"21",X"50",X"43",X"36",X"04",X"23",X"36",
		X"03",X"C9",X"78",X"21",X"75",X"34",X"85",X"6F",X"30",X"01",X"24",X"7E",X"A7",X"C8",X"3D",X"21",
		X"11",X"2F",X"E5",X"EF",X"9E",X"2F",X"A2",X"2F",X"A7",X"2F",X"AC",X"2F",X"B0",X"2F",X"AF",X"06",
		X"01",X"C9",X"3E",X"02",X"06",X"01",X"C9",X"3E",X"02",X"06",X"03",X"C9",X"AF",X"06",X"03",X"C9",
		X"DD",X"36",X"12",X"01",X"DD",X"CB",X"06",X"46",X"28",X"05",X"3E",X"02",X"06",X"03",X"C9",X"AF",
		X"06",X"03",X"C9",X"78",X"21",X"84",X"34",X"85",X"6F",X"30",X"01",X"24",X"7E",X"A7",X"C8",X"3D",
		X"21",X"11",X"2F",X"E5",X"EF",X"DB",X"2F",X"E1",X"2F",X"F1",X"2F",X"DD",X"7E",X"08",X"06",X"00",
		X"C9",X"DD",X"7E",X"12",X"A7",X"20",X"05",X"3E",X"03",X"06",X"00",X"C9",X"DD",X"35",X"12",X"F1",
		X"C9",X"DD",X"7E",X"12",X"A7",X"20",X"F5",X"3E",X"01",X"06",X"00",X"C9",X"78",X"21",X"93",X"34",
		X"85",X"6F",X"30",X"01",X"24",X"7E",X"A7",X"C8",X"3D",X"21",X"11",X"2F",X"E5",X"EF",X"14",X"30",
		X"1A",X"30",X"25",X"30",X"DD",X"7E",X"08",X"06",X"02",X"C9",X"DD",X"7E",X"12",X"A7",X"20",X"CC",
		X"3E",X"03",X"06",X"02",X"C9",X"DD",X"7E",X"12",X"A7",X"20",X"C1",X"3E",X"01",X"06",X"02",X"C9",
		X"C9",X"CD",X"1B",X"32",X"DD",X"35",X"11",X"C0",X"DD",X"7E",X"06",X"21",X"CA",X"30",X"06",X"06",
		X"BE",X"28",X"5A",X"23",X"10",X"FA",X"21",X"D0",X"30",X"3A",X"80",X"42",X"E6",X"01",X"28",X"03",
		X"21",X"DF",X"30",X"DD",X"75",X"0C",X"DD",X"74",X"0D",X"DD",X"36",X"0E",X"00",X"DD",X"36",X"11",
		X"68",X"DD",X"36",X"02",X"04",X"3E",X"01",X"DD",X"86",X"04",X"DD",X"77",X"04",X"CD",X"1B",X"32",
		X"3A",X"F6",X"41",X"A7",X"C0",X"DD",X"7E",X"04",X"D6",X"01",X"DD",X"77",X"04",X"DD",X"7E",X"07",
		X"CD",X"18",X"2F",X"CD",X"1B",X"32",X"DD",X"36",X"02",X"01",X"DD",X"CB",X"01",X"46",X"C8",X"21",
		X"26",X"41",X"7E",X"FE",X"02",X"D0",X"36",X"02",X"AF",X"32",X"81",X"41",X"C9",X"DD",X"7E",X"04",
		X"FE",X"1D",X"38",X"07",X"DD",X"7E",X"03",X"FE",X"80",X"30",X"9B",X"21",X"EE",X"30",X"3A",X"80",
		X"42",X"E6",X"01",X"28",X"03",X"21",X"FD",X"30",X"DD",X"75",X"0C",X"DD",X"74",X"0D",X"DD",X"36",
		X"0E",X"00",X"DD",X"36",X"02",X"06",X"CD",X"4F",X"0B",X"C9",X"03",X"08",X"0D",X"12",X"17",X"1C",
		X"05",X"28",X"0A",X"05",X"29",X"0A",X"05",X"28",X"0A",X"05",X"29",X"0A",X"FF",X"D0",X"30",X"06",
		X"0B",X"0A",X"06",X"1D",X"0A",X"06",X"0B",X"0A",X"06",X"1D",X"0A",X"FF",X"DF",X"30",X"05",X"66",
		X"0A",X"05",X"67",X"0A",X"05",X"66",X"0A",X"05",X"67",X"0A",X"FF",X"EE",X"30",X"06",X"20",X"0A",
		X"06",X"20",X"0A",X"06",X"20",X"0A",X"06",X"20",X"0A",X"FF",X"FD",X"30",X"05",X"36",X"0D",X"05",
		X"37",X"0D",X"FF",X"0C",X"31",X"06",X"5E",X"0D",X"06",X"38",X"0D",X"FF",X"15",X"31",X"01",X"40",
		X"80",X"C0",X"FF",X"20",X"60",X"C9",X"CD",X"1B",X"32",X"3E",X"30",X"DD",X"86",X"03",X"DD",X"77",
		X"03",X"30",X"03",X"DD",X"34",X"04",X"DD",X"7E",X"04",X"FE",X"1D",X"D8",X"DD",X"7E",X"03",X"E6",
		X"E0",X"FE",X"C0",X"D8",X"DD",X"36",X"03",X"C0",X"21",X"0C",X"31",X"3A",X"80",X"42",X"E6",X"01",
		X"28",X"03",X"21",X"15",X"31",X"DD",X"75",X"0C",X"DD",X"74",X"0D",X"DD",X"36",X"0E",X"00",X"21",
		X"1E",X"31",X"3A",X"F8",X"41",X"85",X"6F",X"30",X"01",X"24",X"7E",X"DD",X"77",X"11",X"DD",X"36",
		X"02",X"07",X"CD",X"64",X"0B",X"21",X"F8",X"41",X"34",X"C9",X"CD",X"1B",X"32",X"3A",X"F6",X"41",
		X"A7",X"C0",X"DD",X"35",X"11",X"C0",X"DD",X"7E",X"07",X"CD",X"18",X"2F",X"C3",X"86",X"30",X"21",
		X"CB",X"31",X"3A",X"80",X"42",X"E6",X"01",X"20",X"03",X"21",X"DA",X"31",X"DD",X"75",X"0C",X"DD",
		X"74",X"0D",X"DD",X"36",X"0E",X"00",X"DD",X"36",X"11",X"35",X"DD",X"34",X"02",X"CD",X"1B",X"32",
		X"DD",X"35",X"11",X"C0",X"AF",X"DD",X"77",X"00",X"DD",X"77",X"01",X"DD",X"77",X"07",X"DD",X"77",
		X"0A",X"DD",X"77",X"14",X"DD",X"77",X"06",X"DD",X"77",X"05",X"C9",X"06",X"A0",X"09",X"06",X"1D",
		X"09",X"06",X"1E",X"09",X"06",X"1F",X"09",X"FF",X"CB",X"31",X"05",X"66",X"09",X"05",X"68",X"09",
		X"05",X"66",X"09",X"05",X"68",X"09",X"FF",X"DA",X"31",X"C9",X"3A",X"5F",X"42",X"E6",X"1F",X"C0",
		X"21",X"10",X"41",X"7E",X"A7",X"C8",X"FE",X"01",X"28",X"02",X"35",X"C9",X"36",X"00",X"3A",X"0A",
		X"40",X"FE",X"04",X"28",X"07",X"FE",X"14",X"C0",X"CD",X"40",X"0B",X"C9",X"3A",X"80",X"42",X"E6",
		X"01",X"20",X"04",X"CD",X"1D",X"0B",X"C9",X"CD",X"31",X"0B",X"C9",X"DD",X"7E",X"0E",X"A7",X"28",
		X"04",X"DD",X"35",X"0E",X"C9",X"DD",X"6E",X"0C",X"DD",X"66",X"0D",X"7E",X"FE",X"FF",X"28",X"15",
		X"DD",X"77",X"10",X"23",X"7E",X"DD",X"77",X"0F",X"23",X"7E",X"DD",X"77",X"0E",X"23",X"DD",X"75",
		X"0C",X"DD",X"74",X"0D",X"C9",X"23",X"7E",X"DD",X"77",X"0C",X"23",X"7E",X"DD",X"77",X"0D",X"18",
		X"D4",X"3A",X"F5",X"41",X"A7",X"C8",X"3A",X"F4",X"41",X"A7",X"C8",X"47",X"AF",X"32",X"F4",X"41",
		X"DD",X"21",X"80",X"45",X"11",X"18",X"00",X"DD",X"19",X"10",X"FC",X"21",X"F7",X"41",X"34",X"7E",
		X"FE",X"07",X"28",X"2D",X"FE",X"05",X"38",X"02",X"3E",X"04",X"11",X"12",X"03",X"83",X"5F",X"FF",
		X"7E",X"3D",X"FE",X"06",X"38",X"02",X"36",X"00",X"21",X"FC",X"32",X"CD",X"2B",X"2C",X"DD",X"73",
		X"0C",X"DD",X"72",X"0D",X"DD",X"36",X"0E",X"00",X"DD",X"36",X"11",X"4F",X"DD",X"36",X"02",X"03",
		X"C9",X"3E",X"05",X"18",X"D5",X"DD",X"21",X"98",X"45",X"11",X"18",X"00",X"06",X"07",X"21",X"37",
		X"33",X"3A",X"80",X"42",X"E6",X"01",X"28",X"03",X"21",X"46",X"33",X"DD",X"75",X"0C",X"DD",X"74",
		X"0D",X"DD",X"36",X"0E",X"00",X"CD",X"1B",X"32",X"DD",X"19",X"10",X"E2",X"C9",X"DD",X"21",X"98",
		X"45",X"11",X"18",X"00",X"06",X"07",X"DD",X"7E",X"02",X"FE",X"01",X"20",X"1A",X"21",X"19",X"33",
		X"3A",X"80",X"42",X"E6",X"01",X"28",X"03",X"21",X"28",X"33",X"DD",X"75",X"0C",X"DD",X"74",X"0D",
		X"DD",X"36",X"0E",X"00",X"CD",X"1B",X"32",X"DD",X"19",X"10",X"DB",X"C9",X"0A",X"33",X"0D",X"33",
		X"10",X"33",X"13",X"33",X"13",X"33",X"13",X"33",X"16",X"33",X"06",X"18",X"60",X"06",X"19",X"60",
		X"06",X"1A",X"60",X"06",X"1B",X"60",X"06",X"1C",X"60",X"03",X"2A",X"09",X"03",X"2B",X"09",X"03",
		X"2C",X"09",X"06",X"2D",X"09",X"FF",X"19",X"33",X"01",X"22",X"09",X"01",X"23",X"09",X"01",X"22",
		X"09",X"07",X"23",X"09",X"FF",X"28",X"33",X"03",X"2A",X"09",X"03",X"2B",X"09",X"03",X"2C",X"09",
		X"03",X"2D",X"09",X"FF",X"37",X"33",X"01",X"22",X"09",X"01",X"23",X"09",X"01",X"22",X"09",X"01",
		X"23",X"09",X"FF",X"46",X"33",X"3A",X"F5",X"41",X"A7",X"C8",X"3A",X"5F",X"42",X"E6",X"3F",X"C0",
		X"3A",X"F6",X"41",X"A7",X"28",X"0C",X"3D",X"32",X"F6",X"41",X"28",X"06",X"FE",X"02",X"CA",X"CD",
		X"32",X"C9",X"AF",X"32",X"F5",X"41",X"32",X"F4",X"41",X"32",X"F7",X"41",X"32",X"F8",X"41",X"CD",
		X"CD",X"0B",X"CD",X"86",X"31",X"CD",X"FE",X"31",X"DD",X"21",X"98",X"45",X"11",X"18",X"00",X"06",
		X"07",X"DD",X"7E",X"02",X"FE",X"01",X"20",X"23",X"FE",X"0A",X"28",X"1F",X"3A",X"80",X"42",X"E6",
		X"01",X"20",X"1D",X"21",X"E6",X"33",X"78",X"FE",X"07",X"20",X"03",X"21",X"6B",X"18",X"DD",X"75",
		X"0C",X"DD",X"74",X"0D",X"DD",X"36",X"0E",X"00",X"CD",X"1B",X"32",X"DD",X"19",X"10",X"D2",X"C9",
		X"21",X"2A",X"34",X"78",X"FE",X"07",X"20",X"03",X"21",X"AF",X"18",X"18",X"E1",X"20",X"20",X"22",
		X"22",X"24",X"24",X"26",X"26",X"28",X"28",X"2A",X"2A",X"2C",X"2C",X"2E",X"2E",X"30",X"E6",X"33",
		X"F5",X"33",X"04",X"34",X"13",X"34",X"05",X"2A",X"09",X"05",X"2B",X"09",X"05",X"2C",X"09",X"05",
		X"2D",X"09",X"FF",X"E6",X"33",X"05",X"2A",X"09",X"05",X"2B",X"09",X"05",X"2C",X"09",X"05",X"2D",
		X"09",X"FF",X"F5",X"33",X"05",X"2A",X"09",X"05",X"2B",X"09",X"05",X"2C",X"09",X"05",X"2D",X"09",
		X"FF",X"04",X"34",X"05",X"2A",X"09",X"05",X"2B",X"09",X"05",X"2C",X"09",X"05",X"2D",X"09",X"FF",
		X"13",X"34",X"2A",X"34",X"39",X"34",X"48",X"34",X"57",X"34",X"06",X"22",X"09",X"06",X"23",X"09",
		X"06",X"22",X"09",X"06",X"23",X"09",X"FF",X"2A",X"34",X"06",X"22",X"09",X"06",X"23",X"09",X"06",
		X"22",X"09",X"06",X"23",X"09",X"FF",X"39",X"34",X"06",X"22",X"09",X"06",X"23",X"09",X"06",X"22",
		X"09",X"06",X"23",X"09",X"FF",X"48",X"34",X"06",X"22",X"09",X"06",X"23",X"09",X"06",X"22",X"09",
		X"06",X"23",X"09",X"FF",X"57",X"34",X"00",X"00",X"00",X"04",X"00",X"00",X"03",X"05",X"00",X"00",
		X"00",X"01",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",
		X"01",X"03",X"05",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"00",X"00",X"00",X"00",
		X"02",X"02",X"01",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"03",X"00",X"02",X"00",X"01",X"00",
		X"02",X"00",X"DD",X"7E",X"06",X"87",X"87",X"67",X"DD",X"7E",X"04",X"6F",X"E6",X"07",X"11",X"69",
		X"00",X"83",X"5F",X"1A",X"57",X"7D",X"0F",X"0F",X"0F",X"E6",X"03",X"84",X"5F",X"C9",X"CD",X"A2",
		X"34",X"2A",X"BB",X"40",X"7B",X"85",X"6F",X"30",X"01",X"24",X"E5",X"FD",X"E1",X"06",X"00",X"7A",
		X"FE",X"01",X"28",X"49",X"FE",X"80",X"28",X"24",X"4F",X"79",X"FD",X"A6",X"04",X"28",X"02",X"CB",
		X"C0",X"79",X"FD",X"A6",X"FC",X"28",X"02",X"CB",X"D0",X"79",X"07",X"FD",X"A6",X"00",X"28",X"02",
		X"CB",X"C8",X"79",X"0F",X"FD",X"A6",X"00",X"28",X"02",X"CB",X"D8",X"C9",X"FD",X"CB",X"04",X"7E",
		X"28",X"02",X"CB",X"C0",X"FD",X"CB",X"FC",X"7E",X"28",X"02",X"CB",X"D0",X"FD",X"CB",X"FF",X"46",
		X"28",X"02",X"CB",X"C8",X"FD",X"CB",X"00",X"76",X"28",X"02",X"CB",X"D8",X"C9",X"FD",X"CB",X"04",
		X"46",X"28",X"02",X"CB",X"C0",X"FD",X"CB",X"FC",X"46",X"28",X"02",X"CB",X"D0",X"FD",X"CB",X"00",
		X"4E",X"28",X"02",X"CB",X"C8",X"FD",X"CB",X"01",X"7E",X"28",X"02",X"CB",X"D8",X"C9",X"3A",X"0C",
		X"41",X"FE",X"0F",X"C8",X"3A",X"0F",X"41",X"FE",X"0F",X"C8",X"CD",X"5A",X"35",X"CD",X"AA",X"35",
		X"CD",X"73",X"35",X"CD",X"F0",X"35",X"CD",X"14",X"36",X"C9",X"3A",X"10",X"40",X"0F",X"0F",X"0F",
		X"21",X"09",X"41",X"CB",X"16",X"7E",X"E6",X"07",X"FE",X"01",X"C0",X"CD",X"F4",X"0A",X"3E",X"01",
		X"C3",X"E0",X"35",X"3A",X"10",X"40",X"21",X"0D",X"41",X"07",X"07",X"CB",X"16",X"7E",X"E6",X"07",
		X"FE",X"01",X"C0",X"EB",X"CD",X"F4",X"0A",X"21",X"06",X"41",X"34",X"EB",X"23",X"7E",X"C6",X"10",
		X"77",X"47",X"23",X"7E",X"90",X"D0",X"7E",X"4F",X"E6",X"F0",X"C6",X"10",X"2B",X"ED",X"44",X"86",
		X"77",X"79",X"E6",X"0F",X"FE",X"0F",X"20",X"38",X"18",X"34",X"3A",X"10",X"40",X"21",X"0A",X"41",
		X"07",X"CB",X"16",X"7E",X"E6",X"07",X"FE",X"01",X"C0",X"EB",X"CD",X"F4",X"0A",X"21",X"04",X"41",
		X"34",X"EB",X"23",X"7E",X"C6",X"10",X"77",X"47",X"23",X"7E",X"90",X"D0",X"7E",X"4F",X"E6",X"F0",
		X"C6",X"10",X"2B",X"ED",X"44",X"86",X"77",X"79",X"E6",X"0F",X"FE",X"0F",X"20",X"02",X"3E",X"63",
		X"21",X"02",X"40",X"86",X"77",X"FE",X"63",X"38",X"02",X"36",X"63",X"11",X"01",X"07",X"FF",X"C9",
		X"3A",X"04",X"41",X"A7",X"C8",X"21",X"05",X"41",X"7E",X"A7",X"20",X"07",X"36",X"30",X"3C",X"32",
		X"02",X"68",X"C9",X"35",X"28",X"09",X"7E",X"FE",X"18",X"C0",X"AF",X"32",X"02",X"68",X"C9",X"21",
		X"04",X"41",X"35",X"C9",X"3A",X"06",X"41",X"A7",X"C8",X"21",X"07",X"41",X"7E",X"A7",X"20",X"07",
		X"36",X"30",X"3C",X"32",X"02",X"68",X"C9",X"35",X"28",X"09",X"7E",X"FE",X"18",X"C0",X"AF",X"32",
		X"02",X"68",X"C9",X"21",X"06",X"41",X"35",X"C9",X"7B",X"0F",X"0F",X"0F",X"E6",X"1F",X"67",X"7A",
		X"6F",X"0F",X"0F",X"0F",X"E6",X"07",X"11",X"69",X"00",X"83",X"5F",X"1A",X"57",X"29",X"29",X"7C",
		X"21",X"6E",X"1D",X"CD",X"24",X"2C",X"7A",X"A6",X"20",X"04",X"07",X"30",X"01",X"2B",X"1E",X"00",
		X"E5",X"DD",X"E1",X"7A",X"DD",X"A6",X"FC",X"28",X"02",X"CB",X"DB",X"7A",X"DD",X"A6",X"F8",X"28",
		X"02",X"CB",X"D3",X"7A",X"DD",X"A6",X"F4",X"28",X"02",X"CB",X"CB",X"7A",X"DD",X"A6",X"F0",X"28",
		X"02",X"CB",X"C3",X"7B",X"C9",X"3A",X"05",X"40",X"FE",X"03",X"C0",X"3A",X"0A",X"40",X"FE",X"04",
		X"D8",X"FE",X"06",X"D0",X"21",X"23",X"41",X"34",X"7E",X"FE",X"05",X"38",X"02",X"36",X"00",X"7E",
		X"FE",X"01",X"38",X"0D",X"28",X"10",X"FE",X"03",X"38",X"11",X"28",X"14",X"16",X"6C",X"C3",X"83",
		X"38",X"16",X"1C",X"C3",X"83",X"38",X"16",X"30",X"C3",X"83",X"38",X"16",X"44",X"C3",X"83",X"38",
		X"16",X"58",X"C3",X"83",X"38",X"C9",X"2A",X"28",X"41",X"22",X"2A",X"41",X"DD",X"2A",X"32",X"41",
		X"01",X"00",X"00",X"DD",X"7E",X"00",X"CD",X"63",X"38",X"DD",X"7E",X"01",X"CD",X"73",X"38",X"ED",
		X"5B",X"2A",X"41",X"18",X"0C",X"A7",X"2A",X"28",X"41",X"ED",X"5B",X"2A",X"41",X"ED",X"52",X"28",
		X"32",X"CD",X"26",X"38",X"20",X"1B",X"CD",X"E9",X"37",X"C8",X"04",X"78",X"FE",X"0A",X"D0",X"2A",
		X"30",X"41",X"22",X"2A",X"41",X"21",X"C0",X"42",X"7A",X"CD",X"24",X"2C",X"7B",X"A6",X"C0",X"18",
		X"D4",X"06",X"00",X"DD",X"23",X"2A",X"2E",X"41",X"22",X"2C",X"41",X"DD",X"7E",X"01",X"CD",X"73",
		X"38",X"18",X"DC",X"3A",X"80",X"42",X"E6",X"01",X"28",X"71",X"AF",X"2A",X"34",X"41",X"54",X"5D",
		X"01",X"C0",X"42",X"ED",X"42",X"22",X"34",X"41",X"ED",X"4B",X"BB",X"40",X"09",X"3A",X"20",X"41",
		X"0F",X"4F",X"30",X"02",X"23",X"13",X"A6",X"28",X"07",X"79",X"07",X"4F",X"30",X"02",X"2B",X"1B",
		X"D5",X"DD",X"E1",X"1E",X"00",X"79",X"2F",X"47",X"78",X"DD",X"A6",X"00",X"DD",X"77",X"00",X"78",
		X"DD",X"A6",X"FC",X"DD",X"77",X"FC",X"78",X"DD",X"A6",X"F8",X"DD",X"77",X"F8",X"78",X"DD",X"A6",
		X"F4",X"DD",X"77",X"F4",X"79",X"07",X"4F",X"30",X"03",X"2B",X"DD",X"2B",X"1C",X"A6",X"28",X"D5",
		X"7B",X"C6",X"02",X"CD",X"E6",X"38",X"2A",X"34",X"41",X"ED",X"5B",X"12",X"41",X"19",X"3A",X"20",
		X"41",X"57",X"CD",X"5E",X"36",X"C6",X"02",X"CD",X"F9",X"02",X"C9",X"AF",X"2A",X"34",X"41",X"54",
		X"5D",X"01",X"C0",X"42",X"ED",X"42",X"22",X"34",X"41",X"ED",X"4B",X"BB",X"40",X"09",X"3A",X"20",
		X"41",X"4F",X"D5",X"DD",X"E1",X"1E",X"00",X"79",X"2F",X"47",X"78",X"DD",X"A6",X"00",X"DD",X"77",
		X"00",X"78",X"DD",X"A6",X"FC",X"DD",X"77",X"FC",X"78",X"DD",X"A6",X"F8",X"DD",X"77",X"F8",X"78",
		X"DD",X"A6",X"F4",X"DD",X"77",X"F4",X"79",X"07",X"4F",X"30",X"03",X"2B",X"DD",X"2B",X"1C",X"A6",
		X"28",X"D5",X"7B",X"C6",X"02",X"CD",X"E6",X"38",X"C9",X"3A",X"2B",X"41",X"57",X"3A",X"2D",X"41",
		X"82",X"57",X"32",X"31",X"41",X"3A",X"2A",X"41",X"5F",X"3A",X"2C",X"41",X"83",X"32",X"30",X"41",
		X"0F",X"0F",X"0F",X"E6",X"1F",X"67",X"7A",X"6F",X"0F",X"0F",X"0F",X"E6",X"07",X"D9",X"21",X"69",
		X"00",X"85",X"6F",X"7E",X"D9",X"5F",X"29",X"29",X"7C",X"57",X"2A",X"BB",X"40",X"85",X"6F",X"3E",
		X"00",X"8C",X"67",X"7B",X"A6",X"C9",X"3A",X"2B",X"41",X"57",X"3A",X"2F",X"41",X"82",X"57",X"32",
		X"31",X"41",X"3A",X"2A",X"41",X"5F",X"3A",X"2E",X"41",X"83",X"32",X"30",X"41",X"0F",X"0F",X"0F",
		X"E6",X"1F",X"67",X"7A",X"6F",X"0F",X"0F",X"0F",X"E6",X"07",X"D9",X"21",X"69",X"00",X"85",X"6F",
		X"7E",X"D9",X"5F",X"29",X"29",X"7C",X"57",X"2A",X"BB",X"40",X"85",X"6F",X"3E",X"00",X"8C",X"67",
		X"7B",X"A6",X"C9",X"21",X"F6",X"2C",X"CD",X"23",X"2C",X"7E",X"32",X"2C",X"41",X"23",X"7E",X"32",
		X"2D",X"41",X"C9",X"21",X"F6",X"2C",X"CD",X"23",X"2C",X"7E",X"32",X"2E",X"41",X"23",X"7E",X"32",
		X"2F",X"41",X"C9",X"2A",X"12",X"41",X"7A",X"E7",X"1E",X"00",X"0E",X"80",X"06",X"20",X"79",X"A6",
		X"E5",X"D5",X"C5",X"C4",X"A3",X"38",X"C1",X"D1",X"E1",X"79",X"0F",X"4F",X"30",X"01",X"23",X"1C",
		X"10",X"EC",X"C9",X"7B",X"0F",X"0F",X"0F",X"E6",X"03",X"82",X"21",X"C0",X"42",X"E7",X"79",X"A6",
		X"C8",X"32",X"20",X"41",X"22",X"34",X"41",X"7A",X"87",X"C6",X"08",X"E6",X"F8",X"32",X"28",X"41",
		X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"32",X"21",X"41",X"7B",X"C6",X"02",X"32",X"22",X"41",X"7B",
		X"87",X"87",X"87",X"32",X"29",X"41",X"3E",X"00",X"21",X"2D",X"29",X"CD",X"2B",X"2C",X"EB",X"22",
		X"32",X"41",X"CD",X"C6",X"36",X"C9",X"47",X"3A",X"80",X"42",X"E6",X"01",X"20",X"1A",X"C5",X"06",
		X"06",X"C5",X"CD",X"9E",X"39",X"C1",X"21",X"21",X"41",X"35",X"10",X"F5",X"7E",X"C6",X"06",X"77",
		X"21",X"22",X"41",X"35",X"C1",X"10",X"E7",X"C9",X"C5",X"06",X"06",X"C5",X"CD",X"22",X"39",X"C1",
		X"21",X"21",X"41",X"35",X"10",X"F5",X"7E",X"C6",X"06",X"77",X"21",X"22",X"41",X"35",X"C1",X"10",
		X"E7",X"C9",X"CD",X"A2",X"3B",X"2A",X"BB",X"40",X"3A",X"25",X"41",X"E7",X"E5",X"DD",X"E1",X"21",
		X"C0",X"42",X"3A",X"25",X"41",X"E7",X"E5",X"FD",X"E1",X"06",X"00",X"3A",X"24",X"41",X"4F",X"DD",
		X"A6",X"00",X"28",X"02",X"CB",X"F0",X"79",X"FD",X"A6",X"00",X"28",X"02",X"CB",X"D0",X"79",X"DD",
		X"A6",X"04",X"28",X"02",X"CB",X"E0",X"79",X"FD",X"A6",X"04",X"28",X"02",X"CB",X"C0",X"79",X"07",
		X"4F",X"30",X"04",X"DD",X"2B",X"FD",X"2B",X"DD",X"A6",X"00",X"28",X"02",X"CB",X"E8",X"79",X"FD",
		X"A6",X"00",X"28",X"02",X"CB",X"C8",X"79",X"FD",X"A6",X"04",X"28",X"02",X"CB",X"D8",X"21",X"22",
		X"3B",X"78",X"E7",X"47",X"3A",X"21",X"41",X"2F",X"E6",X"1F",X"87",X"87",X"87",X"6F",X"26",X"00",
		X"29",X"29",X"3A",X"22",X"41",X"85",X"6F",X"78",X"01",X"00",X"48",X"09",X"77",X"C9",X"CD",X"A2",
		X"3B",X"2A",X"BB",X"40",X"3A",X"25",X"41",X"E7",X"E5",X"DD",X"E1",X"21",X"C0",X"42",X"3A",X"25",
		X"41",X"E7",X"E5",X"FD",X"E1",X"06",X"00",X"3A",X"24",X"41",X"4F",X"DD",X"A6",X"00",X"28",X"02",
		X"CB",X"F0",X"79",X"FD",X"A6",X"00",X"28",X"02",X"CB",X"D0",X"79",X"DD",X"A6",X"04",X"28",X"02",
		X"CB",X"E0",X"79",X"FD",X"A6",X"04",X"28",X"02",X"CB",X"C0",X"79",X"07",X"4F",X"30",X"04",X"DD",
		X"2B",X"FD",X"2B",X"DD",X"A6",X"00",X"28",X"02",X"CB",X"E8",X"79",X"FD",X"A6",X"00",X"28",X"02",
		X"CB",X"C8",X"79",X"DD",X"A6",X"04",X"28",X"02",X"CB",X"F8",X"79",X"FD",X"A6",X"04",X"28",X"02",
		X"CB",X"D8",X"78",X"21",X"22",X"3A",X"E7",X"47",X"3A",X"21",X"41",X"2F",X"E6",X"1F",X"87",X"87",
		X"87",X"6F",X"26",X"00",X"29",X"29",X"3A",X"22",X"41",X"85",X"6F",X"78",X"01",X"00",X"48",X"09",
		X"77",X"C9",X"0D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",
		X"00",X"41",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"31",X"00",X"00",
		X"00",X"43",X"5C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"34",X"47",X"00",X"00",
		X"4A",X"4B",X"5D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"00",X"4F",X"00",X"51",
		X"00",X"53",X"5E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"55",X"56",X"57",X"58",X"59",
		X"5A",X"5B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"10",X"0D",X"00",X"00",X"00",X"00",X"00",X"10",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"40",X"0D",X"00",X"00",X"00",X"00",X"10",X"00",X"41",X"00",X"00",X"00",X"00",X"00",X"10",
		X"00",X"41",X"0D",X"00",X"00",X"00",X"10",X"40",X"41",X"42",X"00",X"00",X"00",X"00",X"10",X"40",
		X"41",X"42",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"5C",X"00",X"34",X"47",X"00",X"00",X"4A",X"4B",X"00",X"00",X"34",X"47",X"00",X"00",
		X"4A",X"4B",X"5D",X"38",X"00",X"4F",X"00",X"51",X"00",X"53",X"00",X"38",X"00",X"4F",X"00",X"51",
		X"00",X"53",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0D",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"0D",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"0D",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"0D",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"30",X"30",X"30",X"30",X"31",X"31",X"31",X"31",X"30",X"30",X"30",X"30",X"31",X"31",
		X"31",X"31",X"35",X"33",X"32",X"33",X"34",X"34",X"34",X"34",X"32",X"33",X"32",X"33",X"34",X"34",
		X"34",X"34",X"39",X"36",X"37",X"37",X"38",X"38",X"38",X"38",X"36",X"36",X"37",X"37",X"38",X"38",
		X"38",X"38",X"3F",X"3B",X"3C",X"3D",X"3E",X"3E",X"3E",X"3E",X"3A",X"3B",X"3C",X"3D",X"3E",X"3E",
		X"3E",X"3E",X"3A",X"21",X"41",X"87",X"87",X"67",X"3A",X"22",X"41",X"6F",X"E6",X"07",X"D9",X"21",
		X"69",X"00",X"85",X"6F",X"7E",X"D9",X"32",X"24",X"41",X"7D",X"0F",X"0F",X"0F",X"E6",X"03",X"84",
		X"32",X"25",X"41",X"C9",X"3A",X"26",X"41",X"FE",X"01",X"28",X"26",X"D0",X"3A",X"53",X"43",X"A7",
		X"C8",X"3A",X"3C",X"41",X"A7",X"28",X"79",X"3A",X"86",X"45",X"E6",X"F8",X"6F",X"3A",X"84",X"45",
		X"E6",X"F8",X"67",X"3A",X"42",X"43",X"95",X"28",X"3B",X"06",X"04",X"38",X"42",X"06",X"08",X"18",
		X"3E",X"21",X"38",X"41",X"36",X"00",X"23",X"36",X"00",X"23",X"3A",X"86",X"45",X"77",X"E6",X"F8",
		X"4F",X"23",X"3A",X"84",X"45",X"77",X"E6",X"F8",X"47",X"ED",X"43",X"42",X"43",X"23",X"36",X"00",
		X"23",X"36",X"00",X"21",X"59",X"3C",X"3A",X"80",X"42",X"FE",X"10",X"38",X"02",X"3E",X"0F",X"E7",
		X"32",X"27",X"41",X"C9",X"3A",X"43",X"43",X"94",X"C8",X"06",X"02",X"38",X"02",X"06",X"01",X"0E",
		X"00",X"22",X"42",X"43",X"21",X"38",X"41",X"34",X"7E",X"E6",X"7F",X"CB",X"3F",X"CB",X"11",X"C6",
		X"05",X"E7",X"79",X"A7",X"20",X"02",X"70",X"C9",X"78",X"87",X"87",X"87",X"87",X"B6",X"77",X"C9",
		X"CD",X"F1",X"3B",X"21",X"3C",X"41",X"36",X"FF",X"C9",X"06",X"06",X"05",X"04",X"03",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"3A",X"9A",X"45",X"FE",X"01",X"C0",X"21",
		X"81",X"3D",X"E5",X"3A",X"4F",X"43",X"A7",X"C0",X"DD",X"21",X"98",X"45",X"CD",X"1B",X"32",X"3A",
		X"26",X"41",X"FE",X"01",X"28",X"52",X"38",X"47",X"3A",X"50",X"43",X"E6",X"03",X"20",X"0B",X"3A",
		X"AA",X"45",X"E6",X"07",X"FE",X"04",X"20",X"24",X"18",X"09",X"3A",X"AB",X"45",X"E6",X"07",X"FE",
		X"04",X"20",X"19",X"3A",X"50",X"43",X"CD",X"0B",X"3F",X"20",X"11",X"21",X"51",X"43",X"7E",X"3C",
		X"E6",X"03",X"77",X"21",X"ED",X"3E",X"E7",X"32",X"50",X"43",X"18",X"E7",X"3A",X"50",X"43",X"CD",
		X"F1",X"3E",X"2A",X"40",X"43",X"22",X"AA",X"45",X"2A",X"41",X"43",X"22",X"AB",X"45",X"C9",X"3A",
		X"81",X"41",X"A7",X"C2",X"9B",X"3E",X"18",X"10",X"AF",X"32",X"51",X"43",X"3A",X"80",X"41",X"E6",
		X"3F",X"FE",X"3F",X"C0",X"CD",X"69",X"0B",X"C9",X"2A",X"3A",X"41",X"3A",X"AB",X"45",X"94",X"06",
		X"01",X"30",X"04",X"06",X"02",X"ED",X"44",X"67",X"3A",X"AA",X"45",X"95",X"0E",X"08",X"30",X"04",
		X"0E",X"04",X"ED",X"44",X"6F",X"B4",X"28",X"62",X"3A",X"50",X"43",X"E6",X"03",X"20",X"0B",X"3A",
		X"AA",X"45",X"E6",X"07",X"FE",X"04",X"20",X"A4",X"18",X"0A",X"3A",X"AB",X"45",X"E6",X"07",X"FE",
		X"04",X"C2",X"BC",X"3C",X"3A",X"51",X"43",X"A7",X"20",X"2C",X"7D",X"BC",X"30",X"14",X"78",X"32",
		X"51",X"43",X"CD",X"0B",X"3F",X"20",X"28",X"79",X"32",X"50",X"43",X"CD",X"0B",X"3F",X"C2",X"BC",
		X"3C",X"C9",X"79",X"32",X"51",X"43",X"CD",X"0B",X"3F",X"20",X"14",X"78",X"32",X"50",X"43",X"CD",
		X"0B",X"3F",X"C2",X"BC",X"3C",X"C9",X"3A",X"51",X"43",X"CD",X"0B",X"3F",X"CA",X"BC",X"3C",X"21",
		X"51",X"43",X"7E",X"36",X"00",X"2B",X"77",X"C3",X"BC",X"3C",X"3A",X"27",X"41",X"A7",X"C0",X"3E",
		X"FF",X"32",X"81",X"41",X"3A",X"3D",X"41",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"32",X"50",X"43",
		X"C9",X"3A",X"AA",X"45",X"2E",X"00",X"D6",X"03",X"0F",X"CB",X"1D",X"0F",X"CB",X"1D",X"0F",X"CB",
		X"1D",X"E6",X"1F",X"67",X"22",X"9D",X"45",X"3A",X"AB",X"45",X"C6",X"02",X"2E",X"00",X"0F",X"CB",
		X"1D",X"0F",X"CB",X"1D",X"0F",X"CB",X"1D",X"E6",X"1F",X"67",X"22",X"9B",X"45",X"C9",X"3A",X"48",
		X"43",X"E6",X"03",X"20",X"0E",X"3A",X"86",X"45",X"E6",X"07",X"FE",X"04",X"20",X"1A",X"CD",X"E1",
		X"3D",X"18",X"0C",X"3A",X"84",X"45",X"E6",X"07",X"FE",X"04",X"20",X"0C",X"CD",X"E1",X"3D",X"3A",
		X"48",X"43",X"CD",X"C8",X"26",X"20",X"01",X"C9",X"3A",X"48",X"43",X"32",X"49",X"43",X"C3",X"65",
		X"26",X"3E",X"FF",X"32",X"53",X"43",X"21",X"55",X"43",X"7E",X"3C",X"E6",X"03",X"77",X"23",X"20",
		X"01",X"34",X"3C",X"87",X"47",X"4E",X"21",X"28",X"3E",X"3A",X"80",X"42",X"E6",X"01",X"28",X"03",
		X"21",X"67",X"3E",X"79",X"E7",X"3A",X"55",X"43",X"A7",X"CC",X"1A",X"3E",X"7E",X"07",X"10",X"FD",
		X"E6",X"03",X"21",X"ED",X"3E",X"E7",X"32",X"48",X"43",X"C9",X"7E",X"FE",X"D2",X"C0",X"3A",X"F1",
		X"41",X"A7",X"C0",X"2F",X"32",X"F9",X"41",X"C9",X"FF",X"FF",X"FF",X"C0",X"55",X"6A",X"FF",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"01",X"55",X"AA",X"BF",X"F0",X"01",X"55",X"55",X"55",X"55",X"55",
		X"55",X"AA",X"BF",X"F0",X"01",X"55",X"2A",X"D2",X"AA",X"0A",X"D2",X"AA",X"AA",X"AA",X"AA",X"FF",
		X"EA",X"55",X"40",X"00",X"00",X"3F",X"F0",X"FF",X"EA",X"AF",X"FE",X"AB",X"FF",X"AA",X"80",X"FF",
		X"C0",X"00",X"55",X"6A",X"AA",X"A9",X"55",X"55",X"03",X"FF",X"AB",X"FF",X"00",X"00",X"AA",X"AA",
		X"55",X"5F",X"FF",X"00",X"15",X"5A",X"01",X"55",X"A8",X"00",X"3F",X"FA",X"00",X"00",X"00",X"05",
		X"56",X"55",X"69",X"55",X"AA",X"AF",X"FE",X"FF",X"EA",X"55",X"6A",X"FF",X"EA",X"A5",X"54",X"00",
		X"15",X"5A",X"BF",X"FA",X"A9",X"D2",X"55",X"00",X"00",X"00",X"FF",X"3A",X"50",X"43",X"E6",X"03",
		X"20",X"0B",X"3A",X"AA",X"45",X"E6",X"07",X"FE",X"04",X"20",X"2F",X"18",X"09",X"3A",X"AB",X"45",
		X"E6",X"07",X"FE",X"04",X"20",X"24",X"0E",X"00",X"21",X"39",X"41",X"34",X"7E",X"E6",X"7F",X"CB",
		X"3F",X"CB",X"11",X"C6",X"04",X"E7",X"CB",X"19",X"38",X"07",X"E6",X"0F",X"32",X"50",X"43",X"18",
		X"09",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"32",X"50",X"43",X"3A",X"50",X"43",X"CD",X"F1",X"3E",
		X"3A",X"40",X"43",X"32",X"AA",X"45",X"3A",X"41",X"43",X"32",X"AB",X"45",X"C9",X"01",X"08",X"02",
		X"04",X"CD",X"76",X"2C",X"3A",X"AA",X"45",X"5F",X"3A",X"4B",X"43",X"83",X"32",X"40",X"43",X"3A",
		X"AB",X"45",X"5F",X"3A",X"4C",X"43",X"83",X"32",X"41",X"43",X"C9",X"CD",X"A6",X"2C",X"3A",X"AA",
		X"45",X"5F",X"3A",X"4B",X"43",X"83",X"32",X"40",X"43",X"3A",X"AB",X"45",X"5F",X"3A",X"4C",X"43",
		X"83",X"32",X"41",X"43",X"CD",X"46",X"24",X"2A",X"BB",X"40",X"3A",X"47",X"43",X"E7",X"3A",X"46",
		X"43",X"A6",X"C9",X"3A",X"F1",X"41",X"A7",X"C0",X"3A",X"4F",X"43",X"A7",X"C0",X"3A",X"10",X"41",
		X"A7",X"C0",X"21",X"89",X"42",X"7E",X"A7",X"C0",X"3A",X"2C",X"43",X"E6",X"08",X"C0",X"3A",X"2F",
		X"43",X"E6",X"08",X"C0",X"3A",X"D0",X"42",X"E6",X"08",X"C0",X"3A",X"D3",X"42",X"E6",X"08",X"C0",
		X"36",X"FF",X"21",X"F5",X"41",X"36",X"FF",X"23",X"36",X"0A",X"CD",X"A0",X"0B",X"CD",X"AF",X"0B",
		X"CD",X"6E",X"0B",X"CD",X"A5",X"32",X"C9",X"D9",X"21",X"BE",X"41",X"11",X"BF",X"41",X"01",X"10",
		X"00",X"ED",X"B8",X"21",X"BF",X"41",X"3A",X"B6",X"41",X"AE",X"32",X"AF",X"41",X"21",X"80",X"41",
		X"86",X"D9",X"C9",X"21",X"9F",X"3F",X"11",X"AF",X"41",X"01",X"11",X"00",X"ED",X"B0",X"C9",X"FF",
		X"05",X"F6",X"80",X"32",X"17",X"9C",X"C9",X"DD",X"21",X"74",X"98",X"FD",X"BF",X"24",X"AE",X"46",
		X"FF",X"3A",X"02",X"81",X"E6",X"02",X"28",X"03",X"3E",X"B1",X"C9",X"3E",X"5F",X"C9",X"3A",X"80",
		X"42",X"F5",X"21",X"02",X"82",X"7E",X"E6",X"80",X"28",X"0F",X"F1",X"C9",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F1",X"21",X"FF",X"47",X"FE",X"03",X"28",
		X"05",X"F5",X"AF",X"77",X"F1",X"C9",X"F5",X"7E",X"A7",X"20",X"09",X"3A",X"02",X"40",X"C6",X"04",
		X"32",X"02",X"40",X"77",X"F1",X"C9",X"31",X"FE",X"47",X"C3",X"93",X"00",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
