library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity moon_patrol_sound_prog is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of moon_patrol_sound_prog is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"88",X"08",X"14",X"3F",X"8D",X"51",X"0C",X"24",X"E0",X"91",X"00",X"F9",X"3A",X"1A",X"80",X"C2",
		X"F1",X"35",X"00",X"D1",X"59",X"88",X"89",X"D4",X"2B",X"B0",X"52",X"8D",X"84",X"A1",X"2B",X"84",
		X"A9",X"03",X"F0",X"88",X"21",X"30",X"BF",X"02",X"B9",X"B3",X"40",X"42",X"1D",X"98",X"B2",X"0C",
		X"8A",X"02",X"80",X"09",X"7F",X"91",X"12",X"88",X"23",X"23",X"98",X"D9",X"C3",X"42",X"3B",X"8E",
		X"C2",X"00",X"0A",X"A1",X"9C",X"33",X"38",X"89",X"C7",X"8A",X"10",X"02",X"F9",X"12",X"81",X"22",
		X"2A",X"9B",X"E9",X"B2",X"0F",X"19",X"B9",X"63",X"9A",X"20",X"A0",X"08",X"9A",X"88",X"2F",X"A4",
		X"35",X"20",X"A8",X"83",X"40",X"AA",X"C9",X"89",X"8B",X"90",X"BD",X"92",X"35",X"18",X"C9",X"52",
		X"33",X"29",X"03",X"38",X"9B",X"FD",X"82",X"AA",X"18",X"11",X"0B",X"F9",X"13",X"19",X"92",X"62",
		X"3A",X"CB",X"D8",X"32",X"1A",X"AB",X"83",X"49",X"B4",X"39",X"B9",X"AD",X"CC",X"A2",X"72",X"89",
		X"11",X"09",X"82",X"28",X"88",X"99",X"0E",X"05",X"21",X"89",X"BC",X"CA",X"02",X"99",X"80",X"2A",
		X"EB",X"13",X"33",X"25",X"42",X"43",X"10",X"36",X"09",X"B9",X"CE",X"90",X"14",X"31",X"10",X"9D",
		X"D9",X"80",X"99",X"B8",X"8A",X"AB",X"A8",X"9B",X"B2",X"76",X"34",X"22",X"18",X"09",X"BB",X"98",
		X"33",X"1B",X"DA",X"89",X"92",X"0A",X"BA",X"BD",X"47",X"20",X"9B",X"E9",X"01",X"18",X"88",X"25",
		X"41",X"32",X"33",X"52",X"CD",X"98",X"08",X"09",X"82",X"31",X"AF",X"99",X"90",X"89",X"9C",X"CB",
		X"CA",X"00",X"A0",X"11",X"10",X"B8",X"44",X"64",X"23",X"10",X"9C",X"99",X"C9",X"01",X"20",X"05",
		X"28",X"26",X"22",X"00",X"38",X"DB",X"B0",X"8A",X"A0",X"43",X"53",X"18",X"CD",X"D8",X"03",X"19",
		X"AA",X"9A",X"A9",X"AC",X"B2",X"76",X"22",X"AA",X"99",X"9A",X"90",X"0C",X"CA",X"AB",X"99",X"37",
		X"61",X"00",X"89",X"02",X"09",X"22",X"81",X"BD",X"CB",X"C9",X"05",X"54",X"20",X"08",X"99",X"A9",
		X"22",X"18",X"01",X"18",X"AE",X"B9",X"04",X"48",X"BC",X"88",X"8A",X"EC",X"80",X"11",X"9A",X"99",
		X"93",X"75",X"08",X"98",X"88",X"91",X"89",X"12",X"02",X"9A",X"DB",X"04",X"33",X"82",X"39",X"FA",
		X"24",X"10",X"9A",X"DD",X"91",X"35",X"33",X"10",X"19",X"A1",X"99",X"AB",X"C3",X"77",X"1A",X"AB",
		X"CC",X"90",X"08",X"AC",X"A0",X"23",X"33",X"22",X"05",X"31",X"31",X"13",X"09",X"BA",X"91",X"24",
		X"10",X"2C",X"FC",X"DC",X"A8",X"99",X"99",X"88",X"BE",X"92",X"43",X"14",X"31",X"12",X"34",X"35",
		X"31",X"13",X"42",X"AA",X"CC",X"BD",X"CA",X"BA",X"01",X"00",X"99",X"9B",X"A0",X"82",X"34",X"63",
		X"20",X"81",X"17",X"52",X"00",X"8A",X"9A",X"03",X"32",X"8C",X"CB",X"CD",X"BC",X"AB",X"DA",X"8A",
		X"04",X"53",X"21",X"8A",X"81",X"45",X"42",X"28",X"AD",X"BB",X"A9",X"82",X"62",X"21",X"21",X"88",
		X"88",X"02",X"00",X"AD",X"AA",X"92",X"70",X"8A",X"CC",X"CB",X"BA",X"A8",X"37",X"42",X"00",X"8A",
		X"99",X"AA",X"B8",X"02",X"11",X"0A",X"CA",X"13",X"23",X"75",X"41",X"08",X"99",X"82",X"54",X"32",
		X"98",X"A9",X"9A",X"A9",X"9A",X"82",X"54",X"1D",X"EB",X"CB",X"99",X"03",X"53",X"10",X"99",X"89",
		X"BC",X"92",X"10",X"33",X"65",X"20",X"99",X"AA",X"A1",X"00",X"32",X"1B",X"EE",X"BA",X"01",X"44",
		X"32",X"80",X"13",X"36",X"89",X"A9",X"ED",X"B9",X"88",X"09",X"A0",X"31",X"18",X"07",X"31",X"14",
		X"08",X"80",X"31",X"20",X"09",X"DB",X"98",X"89",X"DD",X"90",X"03",X"82",X"50",X"9C",X"A9",X"12",
		X"9C",X"D8",X"88",X"34",X"83",X"63",X"32",X"12",X"08",X"32",X"AF",X"BB",X"FC",X"9A",X"CC",X"A0",
		X"13",X"42",X"08",X"81",X"11",X"35",X"32",X"42",X"22",X"0C",X"CD",X"98",X"98",X"02",X"08",X"22",
		X"2A",X"DA",X"8A",X"11",X"89",X"DC",X"99",X"B0",X"34",X"9D",X"C8",X"12",X"1A",X"EA",X"99",X"01",
		X"00",X"9A",X"37",X"42",X"36",X"23",X"21",X"98",X"10",X"9A",X"CB",X"AB",X"B3",X"73",X"53",X"10",
		X"AA",X"FA",X"01",X"28",X"AA",X"88",X"90",X"9E",X"DA",X"A0",X"98",X"AC",X"E9",X"82",X"11",X"10",
		X"22",X"81",X"47",X"53",X"22",X"09",X"90",X"89",X"12",X"8C",X"FB",X"AA",X"98",X"9A",X"AB",X"90",
		X"32",X"1B",X"D9",X"45",X"22",X"62",X"22",X"42",X"9C",X"BB",X"BB",X"99",X"02",X"45",X"34",X"23",
		X"9B",X"B9",X"9C",X"BB",X"C8",X"02",X"63",X"39",X"91",X"44",X"30",X"01",X"48",X"BB",X"FC",X"BA",
		X"CC",X"A8",X"10",X"11",X"11",X"89",X"11",X"9D",X"B8",X"03",X"74",X"34",X"20",X"88",X"01",X"23",
		X"20",X"88",X"BF",X"B9",X"9A",X"01",X"08",X"AD",X"05",X"38",X"9B",X"DA",X"93",X"48",X"AB",X"AB",
		X"8B",X"DB",X"99",X"82",X"37",X"29",X"CB",X"A0",X"41",X"53",X"23",X"48",X"12",X"22",X"DD",X"C9",
		X"81",X"34",X"32",X"28",X"9A",X"98",X"39",X"D9",X"8B",X"83",X"53",X"0F",X"A9",X"9E",X"B9",X"8A",
		X"88",X"88",X"25",X"12",X"32",X"BA",X"09",X"27",X"3A",X"9A",X"14",X"53",X"01",X"41",X"10",X"89",
		X"DC",X"BB",X"83",X"52",X"9B",X"DC",X"90",X"10",X"10",X"13",X"12",X"11",X"25",X"40",X"00",X"C8",
		X"8A",X"B1",X"18",X"BC",X"B4",X"34",X"09",X"9D",X"CC",X"BA",X"AC",X"82",X"26",X"32",X"89",X"BC",
		X"DA",X"98",X"21",X"32",X"37",X"31",X"00",X"11",X"A9",X"01",X"8F",X"98",X"00",X"23",X"1A",X"A9",
		X"34",X"03",X"53",X"43",X"32",X"AD",X"DB",X"CB",X"A9",X"BC",X"98",X"0B",X"00",X"61",X"24",X"20",
		X"88",X"35",X"23",X"50",X"08",X"CD",X"B9",X"82",X"64",X"20",X"9A",X"BB",X"B9",X"9D",X"DB",X"90",
		X"10",X"24",X"31",X"31",X"18",X"03",X"38",X"10",X"1A",X"1B",X"FD",X"CA",X"80",X"12",X"33",X"64",
		X"20",X"9A",X"88",X"88",X"98",X"03",X"30",X"BE",X"90",X"09",X"98",X"40",X"0A",X"A4",X"53",X"19",
		X"13",X"9C",X"FD",X"AA",X"A8",X"80",X"19",X"82",X"24",X"22",X"AD",X"90",X"56",X"20",X"99",X"20",
		X"8B",X"BB",X"12",X"1B",X"85",X"30",X"EE",X"B9",X"02",X"42",X"12",X"15",X"22",X"20",X"88",X"11",
		X"88",X"90",X"09",X"BF",X"BC",X"EA",X"A8",X"88",X"9A",X"90",X"09",X"00",X"11",X"32",X"36",X"08",
		X"00",X"05",X"08",X"12",X"33",X"95",X"33",X"13",X"10",X"BC",X"EC",X"99",X"21",X"11",X"33",X"63",
		X"31",X"00",X"AA",X"FC",X"AA",X"80",X"00",X"23",X"40",X"AC",X"B9",X"90",X"92",X"53",X"89",X"FA",
		X"A0",X"02",X"8A",X"91",X"2B",X"DE",X"99",X"81",X"23",X"62",X"30",X"21",X"23",X"28",X"DC",X"BC",
		X"81",X"10",X"99",X"08",X"14",X"72",X"20",X"9A",X"A9",X"99",X"BE",X"B9",X"24",X"18",X"AC",X"03",
		X"10",X"AB",X"A9",X"02",X"34",X"35",X"42",X"00",X"08",X"88",X"29",X"9D",X"A0",X"53",X"2A",X"FB",
		X"BB",X"01",X"00",X"8A",X"A8",X"01",X"90",X"00",X"A1",X"36",X"32",X"02",X"3A",X"AB",X"9C",X"BB",
		X"89",X"8A",X"CC",X"AA",X"32",X"32",X"28",X"32",X"21",X"00",X"25",X"52",X"18",X"8A",X"AA",X"11",
		X"28",X"08",X"20",X"32",X"AD",X"EB",X"A9",X"81",X"42",X"89",X"08",X"99",X"01",X"99",X"99",X"88",
		X"80",X"0A",X"08",X"33",X"52",X"37",X"10",X"AB",X"D9",X"00",X"98",X"01",X"08",X"A8",X"03",X"42",
		X"00",X"00",X"00",X"01",X"F0",X"00",X"04",X"00",X"F0",X"04",X"00",X"E0",X"F0",X"04",X"03",X"FC",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"01",X"F7",X"E1",X"F7",X"B9",X"F7",X"AB",X"F7",X"F1",X"F8",X"03",X"F4",X"F2",
		X"F4",X"F5",X"F5",X"16",X"F5",X"6C",X"F4",X"A7",X"F4",X"A7",X"F4",X"64",X"F8",X"4D",X"F4",X"A8",
		X"F8",X"EC",X"F9",X"5F",X"66",X"F8",X"48",X"10",X"49",X"10",X"4A",X"10",X"4B",X"00",X"4C",X"10",
		X"20",X"EE",X"00",X"28",X"20",X"BD",X"00",X"28",X"20",X"9F",X"00",X"28",X"20",X"86",X"00",X"28",
		X"27",X"07",X"28",X"66",X"F8",X"20",X"86",X"00",X"28",X"20",X"8E",X"00",X"28",X"20",X"9F",X"00",
		X"28",X"20",X"0C",X"01",X"28",X"20",X"86",X"00",X"28",X"20",X"FD",X"00",X"28",X"20",X"7E",X"00",
		X"28",X"20",X"EE",X"00",X"A0",X"67",X"07",X"FF",X"66",X"F8",X"48",X"10",X"49",X"10",X"4A",X"10",
		X"4B",X"00",X"4C",X"10",X"FE",X"F4",X"CD",X"20",X"77",X"00",X"24",X"20",X"7E",X"00",X"24",X"20",
		X"9F",X"00",X"24",X"FE",X"F4",X"CD",X"20",X"EE",X"00",X"60",X"67",X"07",X"FF",X"20",X"EE",X"00",
		X"24",X"20",X"9F",X"00",X"24",X"20",X"77",X"00",X"24",X"20",X"B3",X"00",X"24",X"20",X"8E",X"00",
		X"24",X"20",X"77",X"00",X"24",X"20",X"9F",X"00",X"24",X"20",X"7E",X"00",X"24",X"20",X"6A",X"00",
		X"24",X"FD",X"67",X"01",X"FF",X"66",X"FE",X"48",X"0F",X"41",X"02",X"00",X"CE",X"24",X"00",X"A7",
		X"24",X"00",X"7D",X"24",X"00",X"A7",X"24",X"00",X"58",X"24",X"00",X"A7",X"24",X"00",X"7D",X"24",
		X"00",X"A7",X"24",X"FE",X"F4",X"FB",X"66",X"FE",X"41",X"00",X"48",X"0D",X"C0",X"10",X"30",X"01",
		X"06",X"48",X"0D",X"C0",X"18",X"40",X"01",X"04",X"C0",X"14",X"58",X"FF",X"04",X"48",X"0C",X"C0",
		X"18",X"44",X"01",X"04",X"C0",X"14",X"5C",X"FF",X"04",X"48",X"0B",X"C0",X"18",X"48",X"01",X"04",
		X"C0",X"14",X"60",X"FF",X"04",X"48",X"0A",X"C0",X"14",X"4C",X"01",X"04",X"C0",X"18",X"60",X"FF",
		X"04",X"48",X"0B",X"C0",X"14",X"48",X"01",X"04",X"C0",X"18",X"5C",X"FF",X"04",X"48",X"0C",X"C0",
		X"14",X"44",X"01",X"04",X"C0",X"18",X"58",X"FF",X"04",X"FE",X"F5",X"21",X"6D",X"10",X"46",X"00",
		X"4B",X"00",X"4C",X"02",X"4A",X"10",X"66",X"DD",X"FE",X"F5",X"9F",X"FE",X"F5",X"F4",X"FE",X"F5",
		X"9F",X"FE",X"F5",X"F4",X"FE",X"F6",X"A2",X"FE",X"F6",X"F9",X"FE",X"F5",X"9F",X"FE",X"F5",X"F4",
		X"FE",X"F7",X"54",X"FE",X"F6",X"A2",X"FE",X"F5",X"9F",X"FE",X"F6",X"4B",X"FE",X"F5",X"6C",X"42",
		X"A7",X"43",X"02",X"69",X"0E",X"0D",X"09",X"20",X"0D",X"09",X"20",X"69",X"0E",X"0D",X"09",X"20",
		X"0D",X"09",X"20",X"42",X"51",X"43",X"01",X"69",X"0E",X"0D",X"09",X"20",X"0D",X"09",X"20",X"69",
		X"0E",X"0D",X"09",X"20",X"42",X"7A",X"69",X"0E",X"0D",X"09",X"20",X"0D",X"09",X"20",X"69",X"0E",
		X"0D",X"09",X"20",X"42",X"C1",X"69",X"0E",X"0D",X"09",X"20",X"0D",X"09",X"20",X"42",X"7A",X"69",
		X"0E",X"0D",X"09",X"20",X"0D",X"09",X"20",X"42",X"51",X"43",X"01",X"69",X"0E",X"0D",X"09",X"20",
		X"0D",X"09",X"20",X"FD",X"42",X"A7",X"43",X"02",X"69",X"0E",X"0D",X"09",X"20",X"0D",X"09",X"20",
		X"69",X"0E",X"0D",X"09",X"20",X"0D",X"09",X"20",X"42",X"51",X"43",X"01",X"69",X"0E",X"0D",X"09",
		X"20",X"0D",X"09",X"20",X"69",X"0E",X"0D",X"09",X"20",X"42",X"7A",X"69",X"0E",X"0D",X"09",X"20",
		X"0D",X"09",X"20",X"69",X"0E",X"0D",X"09",X"20",X"42",X"C1",X"69",X"0E",X"0D",X"09",X"20",X"0D",
		X"09",X"20",X"42",X"FC",X"69",X"0E",X"0D",X"09",X"20",X"42",X"DD",X"69",X"0E",X"0D",X"09",X"20",
		X"42",X"C1",X"69",X"0E",X"0D",X"09",X"20",X"0D",X"09",X"20",X"FD",X"42",X"A7",X"43",X"02",X"69",
		X"0E",X"0D",X"09",X"20",X"69",X"0E",X"0D",X"09",X"20",X"0D",X"09",X"20",X"69",X"0E",X"0D",X"09",
		X"20",X"42",X"16",X"69",X"0E",X"0D",X"09",X"20",X"69",X"0E",X"0D",X"09",X"20",X"0D",X"09",X"20",
		X"69",X"0E",X"0D",X"09",X"20",X"42",X"FC",X"43",X"01",X"69",X"0E",X"0D",X"09",X"20",X"69",X"0E",
		X"0D",X"09",X"20",X"0D",X"09",X"20",X"69",X"0E",X"0D",X"09",X"20",X"42",X"DD",X"69",X"0E",X"0D",
		X"09",X"20",X"69",X"0E",X"0D",X"09",X"20",X"0D",X"09",X"20",X"42",X"C1",X"69",X"0E",X"0D",X"09",
		X"20",X"FD",X"42",X"FC",X"43",X"01",X"69",X"0E",X"0D",X"09",X"20",X"0D",X"09",X"20",X"69",X"0E",
		X"0D",X"09",X"20",X"0D",X"09",X"20",X"42",X"FD",X"43",X"00",X"69",X"0E",X"0D",X"09",X"20",X"0D",
		X"09",X"20",X"69",X"0E",X"0D",X"09",X"20",X"42",X"1C",X"43",X"01",X"69",X"0E",X"0D",X"09",X"20",
		X"0D",X"09",X"20",X"69",X"0E",X"0D",X"09",X"20",X"42",X"51",X"69",X"0E",X"0D",X"09",X"20",X"0D",
		X"09",X"20",X"42",X"1C",X"69",X"0E",X"0D",X"09",X"20",X"0D",X"09",X"20",X"42",X"FD",X"43",X"00",
		X"69",X"0E",X"0D",X"09",X"20",X"0D",X"09",X"20",X"FD",X"42",X"FC",X"43",X"01",X"69",X"0E",X"0D",
		X"09",X"20",X"0D",X"09",X"20",X"69",X"0E",X"0D",X"09",X"20",X"0D",X"09",X"20",X"42",X"FD",X"43",
		X"00",X"69",X"0E",X"0D",X"09",X"20",X"0D",X"09",X"20",X"69",X"0E",X"0D",X"09",X"20",X"42",X"1C",
		X"43",X"01",X"69",X"0E",X"0D",X"09",X"20",X"0D",X"09",X"20",X"69",X"0E",X"0D",X"09",X"20",X"42",
		X"51",X"69",X"0E",X"0D",X"09",X"20",X"0D",X"09",X"20",X"42",X"7A",X"43",X"01",X"69",X"0E",X"0D",
		X"09",X"20",X"42",X"65",X"69",X"0E",X"0D",X"09",X"20",X"42",X"51",X"69",X"0E",X"0D",X"09",X"20",
		X"0D",X"09",X"20",X"FD",X"42",X"C1",X"43",X"01",X"69",X"0E",X"0D",X"09",X"20",X"0D",X"09",X"20",
		X"69",X"0E",X"0D",X"09",X"20",X"0D",X"09",X"20",X"42",X"E1",X"43",X"00",X"69",X"0E",X"0D",X"09",
		X"20",X"0D",X"09",X"20",X"69",X"0E",X"0D",X"09",X"20",X"42",X"FD",X"69",X"0E",X"0D",X"09",X"20",
		X"0D",X"09",X"20",X"69",X"0E",X"0D",X"09",X"20",X"42",X"2C",X"43",X"01",X"69",X"0E",X"0D",X"09",
		X"20",X"0D",X"09",X"20",X"42",X"FD",X"43",X"00",X"69",X"0E",X"0D",X"09",X"20",X"0D",X"09",X"20",
		X"42",X"E1",X"69",X"0E",X"0D",X"09",X"20",X"0D",X"09",X"20",X"FD",X"76",X"FE",X"51",X"00",X"58",
		X"0D",X"D0",X"0B",X"20",X"FF",X"04",X"77",X"01",X"FF",X"76",X"FE",X"58",X"10",X"51",X"00",X"5C",
		X"18",X"5D",X"09",X"90",X"18",X"0E",X"60",X"50",X"60",X"72",X"60",X"50",X"60",X"72",X"60",X"50",
		X"60",X"72",X"60",X"50",X"60",X"72",X"60",X"50",X"60",X"72",X"60",X"50",X"60",X"72",X"77",X"01",
		X"FF",X"76",X"FE",X"58",X"10",X"50",X"4C",X"51",X"00",X"5C",X"14",X"1D",X"09",X"E0",X"77",X"01",
		X"FF",X"50",X"70",X"51",X"00",X"76",X"FE",X"58",X"10",X"5B",X"00",X"5C",X"10",X"1D",X"09",X"E0",
		X"77",X"01",X"FF",X"52",X"00",X"53",X"05",X"55",X"00",X"76",X"F9",X"59",X"0F",X"5A",X"0F",X"D4",
		X"08",X"60",X"01",X"04",X"59",X"0E",X"5A",X"0E",X"D4",X"08",X"68",X"01",X"04",X"59",X"0D",X"5A",
		X"0D",X"D4",X"08",X"70",X"01",X"04",X"59",X"0C",X"5A",X"0C",X"D4",X"08",X"78",X"01",X"04",X"59",
		X"0B",X"5A",X"0B",X"D4",X"08",X"80",X"01",X"04",X"59",X"0A",X"5A",X"0A",X"D4",X"08",X"88",X"01",
		X"04",X"59",X"09",X"5A",X"09",X"D4",X"08",X"90",X"01",X"04",X"77",X"06",X"FF",X"6C",X"14",X"6D",
		X"14",X"6E",X"0A",X"42",X"DD",X"43",X"01",X"4A",X"10",X"46",X"00",X"4B",X"00",X"4C",X"04",X"47",
		X"9C",X"FE",X"F8",X"79",X"FE",X"F8",X"79",X"47",X"B8",X"40",X"EE",X"44",X"77",X"45",X"00",X"68",
		X"0F",X"69",X"0F",X"2A",X"0F",X"40",X"47",X"BF",X"FF",X"40",X"EE",X"41",X"00",X"68",X"0F",X"49",
		X"00",X"0D",X"09",X"20",X"0D",X"09",X"20",X"68",X"0F",X"0D",X"09",X"20",X"0D",X"09",X"20",X"40",
		X"86",X"68",X"0F",X"69",X"0F",X"0D",X"09",X"20",X"68",X"0F",X"0D",X"09",X"20",X"48",X"00",X"49",
		X"00",X"0D",X"09",X"20",X"40",X"9F",X"69",X"0F",X"68",X"0F",X"0D",X"09",X"20",X"48",X"00",X"0D",
		X"09",X"20",X"49",X"00",X"0D",X"09",X"20",X"40",X"1C",X"41",X"01",X"68",X"0F",X"0D",X"09",X"20",
		X"40",X"86",X"41",X"00",X"0D",X"09",X"20",X"40",X"0C",X"41",X"01",X"68",X"0F",X"69",X"0F",X"0D",
		X"09",X"20",X"40",X"86",X"41",X"00",X"68",X"0F",X"0D",X"09",X"20",X"40",X"FD",X"68",X"0F",X"49",
		X"00",X"0D",X"09",X"20",X"40",X"7E",X"68",X"0F",X"0D",X"09",X"20",X"FD",X"66",X"F8",X"48",X"10",
		X"49",X"10",X"4A",X"10",X"4B",X"00",X"4C",X"10",X"FE",X"F9",X"2D",X"FE",X"F9",X"46",X"FE",X"F9",
		X"2D",X"20",X"77",X"00",X"28",X"20",X"7E",X"00",X"28",X"20",X"8E",X"00",X"28",X"20",X"9F",X"00",
		X"78",X"FE",X"F9",X"2D",X"FE",X"F9",X"46",X"FE",X"F9",X"2D",X"20",X"3E",X"01",X"28",X"20",X"1C",
		X"01",X"28",X"20",X"FD",X"00",X"28",X"20",X"EE",X"00",X"78",X"67",X"07",X"FF",X"20",X"EE",X"00",
		X"28",X"20",X"9F",X"00",X"28",X"20",X"77",X"00",X"28",X"20",X"5E",X"00",X"28",X"20",X"77",X"00",
		X"28",X"20",X"9F",X"00",X"28",X"FD",X"20",X"59",X"00",X"28",X"20",X"77",X"00",X"28",X"20",X"9F",
		X"00",X"28",X"20",X"4F",X"00",X"28",X"20",X"6A",X"00",X"28",X"20",X"9F",X"00",X"28",X"FD",X"46",
		X"10",X"66",X"C7",X"48",X"10",X"49",X"10",X"4A",X"10",X"4B",X"00",X"4C",X"0A",X"0D",X"09",X"20",
		X"0D",X"09",X"20",X"0D",X"09",X"20",X"4C",X"20",X"0D",X"09",X"FE",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"00",X"00",X"FE",X"67",X"38",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"8E",X"00",X"FF",X"BD",X"FC",X"98",X"86",X"BF",X"C6",X"07",X"BD",X"FC",X"D8",X"86",X"13",
		X"C6",X"0F",X"BD",X"FC",X"D8",X"BD",X"FC",X"AD",X"7F",X"90",X"00",X"0F",X"BD",X"FC",X"48",X"96",
		X"BC",X"2B",X"07",X"BD",X"FE",X"E1",X"86",X"FF",X"97",X"BC",X"0E",X"CE",X"00",X"00",X"DF",X"D1",
		X"96",X"80",X"26",X"0B",X"DE",X"84",X"D6",X"8C",X"BD",X"FD",X"DC",X"DF",X"84",X"97",X"80",X"7C",
		X"00",X"D2",X"96",X"81",X"26",X"0B",X"DE",X"86",X"D6",X"8D",X"BD",X"FD",X"DC",X"DF",X"86",X"97",
		X"81",X"7C",X"00",X"D2",X"96",X"82",X"26",X"0B",X"DE",X"88",X"D6",X"8E",X"BD",X"FD",X"DC",X"DF",
		X"88",X"97",X"82",X"7C",X"00",X"D2",X"96",X"83",X"26",X"0B",X"DE",X"8A",X"D6",X"8F",X"BD",X"FD",
		X"DC",X"DF",X"8A",X"97",X"83",X"96",X"A8",X"27",X"08",X"7F",X"00",X"A8",X"C6",X"08",X"BD",X"FD",
		X"3A",X"96",X"A9",X"27",X"08",X"7F",X"00",X"A9",X"C6",X"09",X"BD",X"FD",X"3A",X"96",X"AA",X"27",
		X"08",X"7F",X"00",X"AA",X"C6",X"0A",X"BD",X"FD",X"3A",X"96",X"AB",X"27",X"08",X"7F",X"00",X"AB",
		X"C6",X"18",X"BD",X"FD",X"53",X"96",X"AC",X"27",X"08",X"7F",X"00",X"AC",X"C6",X"19",X"BD",X"FD",
		X"53",X"96",X"AD",X"27",X"08",X"7F",X"00",X"AD",X"C6",X"1A",X"BD",X"FD",X"53",X"96",X"BE",X"16",
		X"9A",X"D8",X"0F",X"97",X"D8",X"54",X"24",X"09",X"D6",X"CB",X"C1",X"02",X"26",X"03",X"5C",X"D7",
		X"BC",X"C6",X"0F",X"BD",X"FC",X"DE",X"7E",X"FB",X"1B",X"96",X"C1",X"B7",X"08",X"01",X"96",X"C2",
		X"B7",X"08",X"02",X"7C",X"00",X"BD",X"96",X"BF",X"4C",X"97",X"BF",X"44",X"24",X"32",X"DE",X"C3",
		X"09",X"27",X"1E",X"DF",X"C3",X"DE",X"C7",X"A6",X"00",X"44",X"44",X"44",X"44",X"97",X"C1",X"DE",
		X"C5",X"09",X"27",X"15",X"DF",X"C5",X"DE",X"C9",X"A6",X"00",X"44",X"44",X"44",X"44",X"97",X"C2",
		X"3B",X"86",X"01",X"9A",X"BE",X"97",X"BE",X"20",X"E6",X"86",X"02",X"9A",X"BE",X"97",X"BE",X"3B",
		X"96",X"C7",X"81",X"A0",X"25",X"09",X"DE",X"C7",X"A6",X"00",X"97",X"C1",X"08",X"DF",X"C7",X"96",
		X"C9",X"81",X"A0",X"25",X"09",X"DE",X"C9",X"A6",X"00",X"97",X"C2",X"08",X"DF",X"C9",X"96",X"BF",
		X"84",X"0E",X"26",X"CC",X"7C",X"00",X"C0",X"3B",X"96",X"C0",X"27",X"3E",X"7A",X"00",X"C0",X"96",
		X"80",X"27",X"06",X"4C",X"27",X"03",X"7A",X"00",X"80",X"96",X"81",X"27",X"06",X"4C",X"27",X"03",
		X"7A",X"00",X"81",X"96",X"82",X"27",X"06",X"4C",X"27",X"03",X"7A",X"00",X"82",X"96",X"83",X"27",
		X"06",X"4C",X"27",X"03",X"7A",X"00",X"83",X"CE",X"00",X"06",X"A6",X"AD",X"27",X"09",X"4A",X"26",
		X"04",X"6C",X"A7",X"A6",X"B3",X"A7",X"AD",X"09",X"26",X"F0",X"39",X"B7",X"90",X"00",X"C6",X"0E",
		X"BD",X"FD",X"20",X"84",X"1F",X"97",X"BC",X"3B",X"CE",X"FF",X"FF",X"DF",X"00",X"C6",X"4F",X"08",
		X"86",X"00",X"A7",X"80",X"08",X"5A",X"26",X"FA",X"86",X"13",X"97",X"D8",X"39",X"BD",X"FC",X"C3",
		X"86",X"BF",X"97",X"BB",X"C6",X"FF",X"D7",X"82",X"D7",X"B1",X"D7",X"B2",X"D7",X"B3",X"C6",X"17",
		X"7E",X"FC",X"DE",X"86",X"BF",X"97",X"BA",X"C6",X"FF",X"D7",X"80",X"D7",X"81",X"D7",X"AE",X"D7",
		X"AF",X"D7",X"B0",X"C6",X"07",X"7E",X"FC",X"DE",X"7C",X"00",X"BD",X"20",X"04",X"0F",X"7F",X"00",
		X"BD",X"37",X"36",X"C1",X"10",X"2A",X"19",X"86",X"0D",X"97",X"03",X"D7",X"02",X"C6",X"08",X"D7",
		X"03",X"5C",X"32",X"97",X"02",X"96",X"BD",X"27",X"FC",X"D7",X"03",X"5A",X"D7",X"03",X"33",X"39",
		X"86",X"15",X"97",X"03",X"C4",X"0F",X"D7",X"02",X"C6",X"10",X"20",X"E3",X"37",X"20",X"E4",X"37",
		X"86",X"15",X"97",X"03",X"C4",X"0F",X"D7",X"02",X"C6",X"14",X"20",X"0D",X"C1",X"10",X"2A",X"EF",
		X"37",X"86",X"0D",X"97",X"03",X"D7",X"02",X"C6",X"0C",X"4F",X"97",X"03",X"97",X"00",X"D7",X"03",
		X"96",X"02",X"5F",X"D7",X"03",X"5A",X"D7",X"00",X"33",X"39",X"0F",X"BD",X"FD",X"20",X"C6",X"09",
		X"7F",X"00",X"BD",X"84",X"1F",X"81",X"10",X"2A",X"08",X"4A",X"81",X"07",X"2B",X"03",X"BD",X"FD",
		X"0C",X"0E",X"39",X"0F",X"BD",X"FD",X"0F",X"C6",X"11",X"20",X"E5",X"17",X"84",X"0F",X"81",X"08",
		X"2A",X"08",X"A6",X"94",X"AB",X"98",X"A7",X"94",X"20",X"67",X"CB",X"38",X"DE",X"CD",X"A6",X"05",
		X"36",X"DE",X"D1",X"AB",X"94",X"A7",X"94",X"32",X"2B",X"0C",X"24",X"02",X"6C",X"98",X"BD",X"FC",
		X"DD",X"5C",X"A6",X"94",X"20",X"4B",X"25",X"F6",X"6A",X"98",X"20",X"F2",X"6F",X"8C",X"DE",X"CD",
		X"C1",X"A0",X"2B",X"02",X"08",X"08",X"08",X"08",X"08",X"C1",X"C0",X"2B",X"08",X"17",X"84",X"0F",
		X"81",X"08",X"2B",X"01",X"08",X"86",X"01",X"39",X"DF",X"CD",X"DE",X"D1",X"6A",X"90",X"27",X"DC",
		X"C1",X"A0",X"2A",X"10",X"C4",X"1F",X"A6",X"94",X"36",X"DE",X"CD",X"A6",X"03",X"BD",X"FC",X"DD",
		X"0E",X"32",X"08",X"39",X"C1",X"C0",X"2A",X"93",X"A6",X"90",X"44",X"A6",X"94",X"25",X"02",X"A6",
		X"98",X"C4",X"1F",X"BD",X"FC",X"DD",X"0E",X"DE",X"CD",X"A6",X"04",X"39",X"26",X"CA",X"DF",X"CD",
		X"E6",X"00",X"2A",X"03",X"7E",X"FE",X"93",X"C4",X"3F",X"C1",X"20",X"2A",X"11",X"A6",X"01",X"BD",
		X"FC",X"DD",X"0E",X"E6",X"00",X"08",X"08",X"58",X"2B",X"E4",X"A6",X"00",X"08",X"39",X"C4",X"1F",
		X"17",X"84",X"0F",X"26",X"31",X"A6",X"01",X"97",X"CE",X"A6",X"02",X"97",X"CD",X"BD",X"FE",X"D4",
		X"DC",X"CD",X"04",X"DD",X"CD",X"E6",X"00",X"C4",X"1F",X"5C",X"5C",X"BD",X"FE",X"D4",X"7C",X"00",
		X"CE",X"26",X"03",X"7C",X"00",X"CD",X"BD",X"FE",X"D4",X"CB",X"07",X"86",X"09",X"BD",X"FC",X"DE",
		X"0E",X"E6",X"00",X"08",X"20",X"BF",X"80",X"08",X"2B",X"29",X"DD",X"CF",X"84",X"03",X"C1",X"30",
		X"2B",X"02",X"8B",X"03",X"16",X"A6",X"01",X"CE",X"00",X"00",X"3A",X"D6",X"CF",X"C1",X"04",X"2A",
		X"0B",X"A6",X"B4",X"A7",X"AE",X"DE",X"CD",X"D6",X"D0",X"7E",X"FD",X"ED",X"A7",X"B4",X"DE",X"CD",
		X"7E",X"FD",X"F3",X"4C",X"27",X"17",X"5C",X"C1",X"10",X"2A",X"09",X"96",X"BA",X"A4",X"01",X"97",
		X"BA",X"7E",X"FD",X"EF",X"96",X"BB",X"A4",X"01",X"97",X"BB",X"7E",X"FD",X"EF",X"C1",X"10",X"2A",
		X"09",X"96",X"BA",X"AA",X"01",X"97",X"BA",X"7E",X"FD",X"EF",X"96",X"BB",X"AA",X"01",X"97",X"BB",
		X"7E",X"FD",X"EF",X"C1",X"F0",X"2A",X"17",X"A6",X"01",X"EE",X"02",X"3C",X"DE",X"D1",X"E7",X"8C",
		X"4C",X"A7",X"90",X"32",X"A7",X"94",X"32",X"A7",X"98",X"DE",X"CD",X"86",X"01",X"39",X"5C",X"27",
		X"12",X"DE",X"D1",X"5C",X"26",X"10",X"DC",X"CD",X"A7",X"9C",X"E7",X"A0",X"DE",X"CD",X"EE",X"01",
		X"86",X"01",X"39",X"86",X"FF",X"39",X"A6",X"9C",X"E6",X"A0",X"DD",X"CD",X"DE",X"CD",X"08",X"08",
		X"08",X"86",X"01",X"39",X"96",X"CE",X"BD",X"FC",X"DD",X"5C",X"96",X"CD",X"BD",X"FC",X"DE",X"5C",
		X"39",X"26",X"06",X"BD",X"FC",X"98",X"7E",X"FC",X"AD",X"81",X"10",X"2B",X"03",X"7E",X"FF",X"25",
		X"97",X"CB",X"96",X"D8",X"8A",X"01",X"16",X"C4",X"FE",X"D7",X"D8",X"C6",X"0F",X"BD",X"FC",X"DE",
		X"86",X"05",X"7F",X"00",X"BD",X"D6",X"BD",X"27",X"FC",X"4A",X"26",X"F6",X"D6",X"CB",X"58",X"58",
		X"CE",X"F4",X"00",X"3A",X"3C",X"EE",X"00",X"DF",X"C7",X"38",X"EE",X"02",X"DF",X"C3",X"96",X"BE",
		X"84",X"02",X"97",X"BE",X"39",X"16",X"58",X"CE",X"F4",X"24",X"3A",X"EE",X"00",X"81",X"14",X"2A",
		X"1C",X"D6",X"82",X"5C",X"27",X"06",X"91",X"A6",X"27",X"02",X"2A",X"10",X"97",X"A6",X"DF",X"88",
		X"7F",X"00",X"82",X"7F",X"00",X"8E",X"C6",X"89",X"DA",X"BB",X"D7",X"BB",X"39",X"26",X"11",X"DF",
		X"8A",X"97",X"A7",X"7F",X"00",X"83",X"7F",X"00",X"8F",X"86",X"B6",X"9A",X"BB",X"97",X"BB",X"39",
		X"81",X"18",X"2A",X"0B",X"DF",X"86",X"97",X"A5",X"7F",X"00",X"81",X"7F",X"00",X"8D",X"39",X"3C",
		X"36",X"BD",X"FC",X"98",X"BD",X"FC",X"AD",X"32",X"38",X"DF",X"84",X"97",X"A4",X"7F",X"00",X"80",
		X"7F",X"00",X"8C",X"86",X"BE",X"9A",X"BA",X"97",X"BA",X"39",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FB",X"00",X"FB",X"00",X"FB",X"00",X"FB",X"00",X"FC",X"8B",X"FB",X"00",X"FB",X"D9",X"FB",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
