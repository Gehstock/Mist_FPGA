library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity GFX1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of GFX1 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"9C",X"63",X"41",X"9C",X"BE",X"BE",X"41",X"00",X"41",X"14",X"36",X"41",X"63",X"63",X"14",X"00",
		X"41",X"41",X"FF",X"00",X"41",X"41",X"FF",X"00",X"00",X"22",X"77",X"00",X"00",X"00",X"77",X"00",
		X"41",X"FF",X"DD",X"63",X"C9",X"77",X"DD",X"00",X"63",X"14",X"55",X"22",X"77",X"36",X"14",X"00",
		X"36",X"C9",X"C9",X"22",X"FF",X"63",X"C9",X"00",X"14",X"14",X"77",X"00",X"36",X"14",X"55",X"00",
		X"14",X"14",X"FF",X"9C",X"FF",X"9C",X"14",X"00",X"00",X"63",X"77",X"00",X"77",X"41",X"36",X"00",
		X"BE",X"41",X"41",X"22",X"FF",X"63",X"41",X"00",X"00",X"55",X"55",X"77",X"55",X"77",X"55",X"00",
		X"36",X"C9",X"C9",X"BE",X"FF",X"FF",X"C9",X"00",X"00",X"36",X"14",X"41",X"14",X"63",X"14",X"00",
		X"00",X"77",X"88",X"00",X"00",X"00",X"FF",X"00",X"36",X"14",X"55",X"36",X"77",X"36",X"14",X"00",
		X"36",X"C9",X"DD",X"36",X"77",X"C9",X"DD",X"00",X"00",X"55",X"14",X"63",X"63",X"77",X"14",X"00",
		X"9C",X"C9",X"EB",X"00",X"BE",X"C9",X"C9",X"00",X"63",X"14",X"14",X"63",X"77",X"77",X"14",X"00",
		X"F0",X"FF",X"F0",X"F0",X"F0",X"F0",X"FF",X"F0",X"F1",X"FF",X"F1",X"F1",X"F1",X"F1",X"FF",X"F1",
		X"F0",X"FF",X"F0",X"F0",X"F0",X"F0",X"FF",X"F0",X"F0",X"F1",X"F0",X"F1",X"F0",X"F1",X"F1",X"F1",
		X"F0",X"FF",X"F0",X"F0",X"F0",X"F0",X"FF",X"F0",X"F1",X"F1",X"F1",X"F0",X"F1",X"F0",X"F1",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"FF",X"F0",X"F1",X"F0",X"F1",X"FF",X"F1",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F1",X"FF",X"F1",X"F0",X"F1",X"F0",X"FF",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",
		X"F0",X"FF",X"F0",X"F0",X"F0",X"F0",X"FF",X"F0",X"F0",X"FF",X"F0",X"F0",X"F0",X"F0",X"FF",X"F0",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"90",X"F0",X"F8",X"B8",X"B8",X"F8",X"F0",X"90",X"60",X"F0",X"B2",X"32",X"32",X"B2",X"F0",X"60",
		X"00",X"00",X"36",X"36",X"36",X"36",X"00",X"00",X"00",X"00",X"36",X"36",X"36",X"36",X"00",X"00",
		X"FC",X"F5",X"F1",X"F2",X"F2",X"F9",X"F5",X"FC",X"F3",X"FA",X"F8",X"F4",X"F4",X"F9",X"FA",X"F3",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"BF",X"FF",X"BF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"BF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"BF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"BF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"88",X"36",X"22",X"88",X"9C",X"9C",X"22",X"00",X"63",X"88",X"9C",X"63",X"77",X"77",X"88",X"00",
		X"22",X"22",X"BE",X"00",X"22",X"22",X"BE",X"00",X"00",X"14",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"22",X"BE",X"AA",X"36",X"22",X"BE",X"AA",X"00",X"36",X"C9",X"EB",X"14",X"FF",X"9C",X"C9",X"00",
		X"9C",X"22",X"22",X"14",X"BE",X"36",X"22",X"00",X"88",X"C9",X"FF",X"00",X"DD",X"88",X"EB",X"00",
		X"88",X"88",X"BE",X"88",X"BE",X"88",X"88",X"00",X"00",X"36",X"FF",X"41",X"FF",X"63",X"9C",X"00",
		X"9C",X"22",X"22",X"14",X"BE",X"36",X"22",X"00",X"41",X"AA",X"AA",X"BE",X"EB",X"BE",X"AA",X"00",
		X"9C",X"22",X"22",X"9C",X"BE",X"BE",X"22",X"00",X"00",X"DD",X"C9",X"63",X"C9",X"77",X"C9",X"00",
		X"00",X"BE",X"00",X"00",X"00",X"00",X"BE",X"00",X"9C",X"88",X"EB",X"9C",X"BE",X"9C",X"C9",X"00",
		X"9C",X"22",X"AA",X"9C",X"BE",X"22",X"AA",X"00",X"00",X"EB",X"C9",X"36",X"36",X"FF",X"C9",X"00",
		X"88",X"22",X"36",X"00",X"9C",X"22",X"22",X"00",X"77",X"C9",X"C9",X"36",X"FF",X"FF",X"C9",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"BE",X"88",X"88",X"BE",X"BE",X"BE",X"88",X"00",X"63",X"9C",X"9C",X"63",X"77",X"77",X"88",X"00",
		X"9C",X"22",X"22",X"BE",X"BE",X"BE",X"22",X"00",X"36",X"C9",X"C9",X"FF",X"FF",X"FF",X"C9",X"00",
		X"14",X"36",X"22",X"88",X"36",X"9C",X"22",X"00",X"14",X"9C",X"88",X"63",X"9C",X"77",X"88",X"00",
		X"88",X"22",X"36",X"BE",X"9C",X"BE",X"22",X"00",X"63",X"88",X"9C",X"FF",X"77",X"FF",X"88",X"00",
		X"22",X"BE",X"22",X"00",X"22",X"BE",X"22",X"00",X"88",X"FF",X"C9",X"00",X"C9",X"FF",X"C9",X"00",
		X"00",X"00",X"00",X"BE",X"00",X"BE",X"00",X"00",X"88",X"C9",X"C9",X"FF",X"C9",X"FF",X"C9",X"00",
		X"BE",X"36",X"22",X"88",X"BE",X"9C",X"22",X"00",X"C9",X"9C",X"C9",X"63",X"C9",X"77",X"88",X"00",
		X"BE",X"00",X"00",X"BE",X"BE",X"BE",X"00",X"00",X"FF",X"41",X"41",X"FF",X"FF",X"FF",X"41",X"00",
		X"22",X"22",X"BE",X"00",X"22",X"22",X"BE",X"00",X"88",X"88",X"FF",X"00",X"88",X"88",X"FF",X"00",
		X"9C",X"22",X"22",X"14",X"BE",X"36",X"22",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"22",X"88",X"BE",X"BE",X"36",X"BE",X"9C",X"00",X"88",X"41",X"36",X"FF",X"9C",X"FF",X"63",X"00",
		X"22",X"BE",X"22",X"00",X"22",X"BE",X"22",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"BE",X"00",X"00",X"BE",X"BE",X"BE",X"88",X"00",X"FF",X"77",X"77",X"FF",X"FF",X"FF",X"63",X"00",
		X"BE",X"00",X"9C",X"BE",X"BE",X"BE",X"88",X"00",X"FF",X"77",X"41",X"FF",X"FF",X"FF",X"63",X"00",
		X"9C",X"22",X"22",X"9C",X"BE",X"BE",X"22",X"00",X"77",X"88",X"88",X"77",X"FF",X"FF",X"88",X"00",
		X"00",X"88",X"88",X"BE",X"88",X"BE",X"88",X"00",X"77",X"88",X"88",X"FF",X"FF",X"FF",X"88",X"00",
		X"AA",X"22",X"BE",X"9C",X"9C",X"BE",X"AA",X"00",X"77",X"88",X"88",X"77",X"FF",X"FF",X"88",X"00",
		X"22",X"88",X"BE",X"BE",X"36",X"BE",X"9C",X"00",X"77",X"88",X"C9",X"FF",X"FF",X"FF",X"88",X"00",
		X"9C",X"22",X"22",X"14",X"BE",X"36",X"22",X"00",X"00",X"C9",X"DD",X"36",X"55",X"FF",X"C9",X"00",
		X"00",X"00",X"BE",X"00",X"00",X"00",X"BE",X"00",X"88",X"88",X"FF",X"00",X"88",X"88",X"FF",X"00",
		X"9C",X"22",X"22",X"9C",X"BE",X"BE",X"22",X"00",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"9C",X"9C",X"00",X"88",X"88",X"BE",X"00",X"FF",X"41",X"41",X"FF",X"FF",X"FF",X"00",X"00",
		X"BE",X"9C",X"9C",X"BE",X"BE",X"BE",X"88",X"00",X"FF",X"41",X"41",X"FF",X"FF",X"FF",X"63",X"00",
		X"36",X"9C",X"9C",X"36",X"BE",X"BE",X"88",X"00",X"9C",X"77",X"77",X"9C",X"BE",X"BE",X"63",X"00",
		X"00",X"00",X"BE",X"00",X"00",X"00",X"BE",X"00",X"BE",X"FF",X"41",X"00",X"FF",X"BE",X"41",X"00",
		X"22",X"BE",X"22",X"36",X"22",X"BE",X"AA",X"00",X"9C",X"C9",X"FF",X"88",X"BE",X"88",X"EB",X"00",
		X"C0",X"50",X"09",X"48",X"50",X"11",X"49",X"50",X"01",X"27",X"00",X"1E",X"00",X"ED",X"98",X"1A",
		X"C0",X"50",X"09",X"D8",X"67",X"11",X"D9",X"67",X"01",X"27",X"00",X"1E",X"00",X"ED",X"98",X"1A",
		X"C0",X"50",X"09",X"40",X"50",X"11",X"41",X"50",X"01",X"37",X"00",X"1E",X"00",X"ED",X"98",X"09",
		X"24",X"64",X"11",X"25",X"64",X"01",X"67",X"00",X"1E",X"FF",X"ED",X"98",X"09",X"7B",X"38",X"0A",
		X"6C",X"3F",X"BF",X"DE",X"DE",X"BF",X"3F",X"6C",X"93",X"3F",X"7F",X"E7",X"E7",X"7F",X"3F",X"93",
		X"6C",X"2F",X"2F",X"DE",X"DE",X"2F",X"2F",X"6C",X"93",X"1F",X"1F",X"E7",X"E7",X"1F",X"1F",X"93",
		X"6C",X"0F",X"0F",X"4E",X"4E",X"0F",X"0F",X"6C",X"93",X"0F",X"0F",X"87",X"87",X"0F",X"0F",X"93",
		X"F0",X"7F",X"FC",X"F8",X"F8",X"FC",X"7F",X"F0",X"F1",X"9F",X"B7",X"F3",X"F3",X"B7",X"9F",X"F1",
		X"F0",X"FF",X"F0",X"F0",X"F0",X"F0",X"FF",X"F0",X"F1",X"FF",X"F1",X"F1",X"F1",X"F1",X"FF",X"F1",
		X"F0",X"2D",X"F0",X"F0",X"F0",X"F0",X"2D",X"F0",X"F0",X"78",X"39",X"E4",X"C6",X"78",X"78",X"F0",
		X"6C",X"01",X"01",X"82",X"82",X"01",X"01",X"6C",X"93",X"08",X"08",X"84",X"84",X"08",X"08",X"93",
		X"F0",X"78",X"F0",X"F0",X"F0",X"F0",X"78",X"78",X"93",X"93",X"B1",X"B1",X"B1",X"B1",X"93",X"B1",
		X"E4",X"78",X"E4",X"F0",X"D2",X"F0",X"78",X"F0",X"F0",X"B1",X"F0",X"E4",X"F0",X"D2",X"B1",X"D2",
		X"F0",X"78",X"F0",X"D2",X"F0",X"A5",X"78",X"F0",X"F0",X"B1",X"5A",X"F0",X"E4",X"F0",X"B1",X"F0",
		X"F0",X"78",X"F0",X"F0",X"F0",X"F0",X"78",X"F0",X"F0",X"D2",X"B1",X"F0",X"F0",X"B1",X"D2",X"F0",
		X"F0",X"E4",X"78",X"F0",X"F0",X"78",X"E4",X"F0",X"F0",X"E4",X"D2",X"B1",X"B1",X"D2",X"E4",X"F0",
		X"F0",X"D2",X"E4",X"78",X"78",X"E4",X"D2",X"F0",X"B1",X"78",X"E4",X"D2",X"D2",X"E4",X"78",X"B1",
		X"E4",X"F0",X"93",X"E4",X"E4",X"93",X"F0",X"E4",X"D2",X"F0",X"6C",X"D2",X"D2",X"6C",X"F0",X"D2",
		X"78",X"93",X"E4",X"78",X"78",X"E4",X"93",X"78",X"B1",X"6C",X"D2",X"B1",X"B1",X"D2",X"6C",X"B1",
		X"78",X"87",X"78",X"78",X"78",X"78",X"87",X"78",X"B1",X"4E",X"B1",X"B1",X"B1",X"B1",X"4E",X"B1",
		X"F0",X"6C",X"78",X"F0",X"F0",X"78",X"6C",X"F0",X"4E",X"B1",X"93",X"87",X"87",X"93",X"B1",X"4E",
		X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"B1",X"B1",X"B1",X"B1",X"B1",X"B1",X"B1",X"B1",
		X"87",X"78",X"6C",X"4E",X"4E",X"6C",X"78",X"87",X"F0",X"93",X"B1",X"F0",X"F0",X"B1",X"93",X"F0",
		X"6C",X"B1",X"B1",X"D2",X"D2",X"B1",X"B1",X"6C",X"93",X"78",X"78",X"E4",X"E4",X"78",X"78",X"93",
		X"F0",X"B1",X"4E",X"F0",X"F0",X"4E",X"B1",X"F0",X"F0",X"78",X"87",X"F0",X"F0",X"87",X"78",X"F0",
		X"F0",X"2D",X"93",X"F0",X"F0",X"93",X"2D",X"F0",X"F0",X"1B",X"6C",X"F0",X"F0",X"6C",X"1B",X"F0",
		X"F0",X"6C",X"E4",X"78",X"78",X"E4",X"6C",X"F0",X"F0",X"93",X"D2",X"B1",X"B1",X"D2",X"93",X"F0",
		X"F0",X"5A",X"D2",X"E4",X"E4",X"D2",X"5A",X"F0",X"F0",X"A5",X"E4",X"D2",X"D2",X"E4",X"A5",X"F0",
		X"C6",X"39",X"B1",X"B1",X"B1",X"B1",X"39",X"C6",X"C6",X"39",X"78",X"78",X"78",X"78",X"39",X"C6",
		X"78",X"B1",X"D2",X"78",X"78",X"D2",X"B1",X"78",X"B1",X"78",X"E4",X"B1",X"B1",X"E4",X"78",X"B1",
		X"C6",X"F0",X"39",X"78",X"39",X"78",X"F0",X"F0",X"F0",X"F0",X"B1",X"39",X"B1",X"39",X"F0",X"C6",
		X"F0",X"78",X"78",X"B1",X"F0",X"39",X"78",X"C6",X"C6",X"B1",X"39",X"F0",X"78",X"B1",X"B1",X"F0",
		X"F0",X"B1",X"4E",X"F0",X"F0",X"4E",X"B1",X"F0",X"F0",X"78",X"87",X"F0",X"F0",X"87",X"78",X"F0",
		X"F0",X"B1",X"B1",X"4E",X"4E",X"B1",X"B1",X"F0",X"F0",X"78",X"78",X"87",X"87",X"78",X"78",X"F0",
		X"4E",X"B1",X"B1",X"B1",X"B1",X"B1",X"B1",X"4E",X"87",X"78",X"78",X"78",X"78",X"78",X"78",X"87",
		X"F0",X"6C",X"78",X"F0",X"F0",X"78",X"6C",X"F0",X"F0",X"93",X"B1",X"F0",X"F0",X"B1",X"93",X"F0",
		X"F0",X"4E",X"6C",X"78",X"78",X"6C",X"4E",X"F0",X"F0",X"87",X"93",X"B1",X"B1",X"93",X"87",X"F0",
		X"78",X"0F",X"4E",X"6C",X"6C",X"4E",X"0F",X"78",X"B1",X"0F",X"87",X"93",X"93",X"87",X"0F",X"B1",
		X"C6",X"F0",X"B1",X"93",X"93",X"B1",X"F0",X"C6",X"C6",X"F0",X"78",X"6C",X"6C",X"78",X"F0",X"C6",
		X"4E",X"B1",X"93",X"87",X"87",X"93",X"B1",X"4E",X"87",X"78",X"6C",X"4E",X"4E",X"6C",X"78",X"87",
		X"6C",X"93",X"87",X"0F",X"0F",X"87",X"93",X"6C",X"87",X"6C",X"4E",X"0F",X"0F",X"4E",X"6C",X"87",
		X"93",X"F0",X"E4",X"B1",X"B1",X"E4",X"F0",X"93",X"6C",X"F0",X"D2",X"78",X"78",X"D2",X"F0",X"6C",
		X"F0",X"78",X"D2",X"C6",X"C6",X"D2",X"78",X"F0",X"F0",X"B1",X"E4",X"C6",X"C6",X"E4",X"B1",X"F0",
		X"F0",X"6C",X"6C",X"F0",X"F0",X"6C",X"6C",X"F0",X"F0",X"93",X"93",X"F0",X"F0",X"93",X"93",X"F0",
		X"F0",X"0F",X"D2",X"F0",X"F0",X"D2",X"0F",X"F0",X"F0",X"0F",X"E4",X"F0",X"F0",X"E4",X"0F",X"F0",
		X"F0",X"78",X"F0",X"87",X"F0",X"87",X"78",X"C6",X"C6",X"B1",X"4E",X"F0",X"4E",X"F0",X"B1",X"F0",
		X"C6",X"78",X"87",X"F0",X"87",X"F0",X"78",X"F0",X"F0",X"B1",X"F0",X"4E",X"F0",X"4E",X"B1",X"C6",
		X"B0",X"F0",X"E0",X"F0",X"D0",X"F0",X"70",X"F0",X"F0",X"B0",X"F0",X"E0",X"F0",X"D0",X"F0",X"70",
		X"F1",X"FF",X"F7",X"FF",X"F3",X"FF",X"FF",X"FF",X"F0",X"F1",X"F0",X"F7",X"F0",X"F3",X"F0",X"FF",
		X"F0",X"F8",X"F0",X"FE",X"F0",X"FC",X"F0",X"FF",X"F8",X"FF",X"FE",X"FF",X"FC",X"FF",X"FF",X"FF",
		X"F0",X"00",X"F0",X"F0",X"F0",X"F0",X"00",X"F0",X"F0",X"00",X"F0",X"F0",X"F0",X"F0",X"00",X"F0",
		X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"B0",X"B0",X"B0",X"B0",X"B0",X"B0",X"B0",X"B0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"F3",X"FF",X"F7",X"FF",X"F1",X"FF",X"F0",X"F3",X"F0",X"F7",X"F0",X"F1",X"F0",
		X"FF",X"F0",X"FC",X"F0",X"FE",X"F0",X"F8",X"F0",X"FF",X"FF",X"FF",X"FC",X"FF",X"FE",X"FF",X"F8",
		X"1D",X"1E",X"20",X"2C",X"52",X"54",X"54",X"13",X"1F",X"19",X"59",X"18",X"50",X"17",X"52",X"54",
		X"20",X"63",X"69",X"15",X"61",X"54",X"68",X"1C",X"1B",X"1E",X"20",X"16",X"1F",X"13",X"19",X"E3",
		X"CE",X"E3",X"AE",X"09",X"96",X"64",X"E3",X"A6",X"E3",X"96",X"E3",X"B6",X"09",X"97",X"64",X"E3",
		X"96",X"09",X"96",X"64",X"E3",X"C6",X"09",X"24",X"64",X"11",X"25",X"64",X"01",X"67",X"00",X"1E",
		X"FF",X"ED",X"98",X"3E",X"FF",X"1A",X"01",X"50",X"09",X"97",X"64",X"E3",X"56",X"08",X"27",X"3A",
		X"FD",X"64",X"3C",X"1A",X"FD",X"64",X"FE",X"14",X"08",X"04",X"E3",X"D6",X"E3",X"F6",X"00",X"1A",
		X"C0",X"50",X"3E",X"40",X"E5",X"FD",X"14",X"3E",X"03",X"E5",X"25",X"15",X"3A",X"B3",X"64",X"FE",
		X"00",X"E2",X"14",X"22",X"3A",X"B2",X"64",X"FE",X"02",X"18",X"64",X"11",X"58",X"41",X"09",X"9C",
		X"30",X"3E",X"01",X"06",X"23",X"E5",X"D5",X"15",X"3A",X"40",X"50",X"E3",X"6F",X"08",X"5C",X"3A",
		X"B3",X"64",X"FE",X"00",X"28",X"15",X"3A",X"B2",X"64",X"FE",X"02",X"38",X"4E",X"D6",X"02",X"1A",
		X"B2",X"64",X"3A",X"B5",X"64",X"D6",X"01",X"0F",X"1A",X"B5",X"64",X"09",X"96",X"64",X"E3",X"CE",
		X"3A",X"8A",X"64",X"1A",X"8E",X"64",X"E5",X"13",X"00",X"3A",X"B3",X"64",X"FE",X"00",X"E2",X"6F",
		X"22",X"E5",X"35",X"15",X"C3",X"6F",X"22",X"FE",X"04",X"18",X"29",X"11",X"26",X"41",X"09",X"BF",
		X"30",X"3E",X"01",X"06",X"11",X"E5",X"D5",X"15",X"11",X"10",X"42",X"09",X"D0",X"30",X"3E",X"01",
		X"06",X"02",X"E5",X"D5",X"15",X"11",X"5A",X"41",X"09",X"9C",X"30",X"3E",X"01",X"06",X"23",X"E5",
		X"D5",X"15",X"30",X"94",X"11",X"90",X"40",X"09",X"D2",X"30",X"3E",X"01",X"06",X"31",X"E5",X"D5",
		X"15",X"30",X"85",X"3A",X"40",X"50",X"E3",X"5F",X"08",X"1B",X"3A",X"B3",X"64",X"FE",X"00",X"28",
		X"15",X"3A",X"B2",X"64",X"FE",X"04",X"38",X"0D",X"D6",X"04",X"1A",X"B2",X"64",X"3A",X"B5",X"64",
		X"D6",X"02",X"0F",X"1A",X"B5",X"64",X"09",X"96",X"64",X"E3",X"8E",X"3A",X"8A",X"64",X"1A",X"8E",
		X"64",X"1A",X"8F",X"64",X"E5",X"13",X"00",X"E5",X"0C",X"00",X"C3",X"F1",X"21",X"1A",X"C0",X"50",
		X"09",X"95",X"64",X"E3",X"5E",X"08",X"03",X"C3",X"A8",X"21",X"E3",X"9E",X"C3",X"7F",X"21",X"AF",
		X"09",X"A8",X"64",X"11",X"A9",X"64",X"01",X"05",X"00",X"5F",X"ED",X"98",X"1A",X"99",X"64",X"1A",
		X"9A",X"64",X"3E",X"40",X"09",X"CC",X"43",X"11",X"CD",X"43",X"01",X"05",X"00",X"5F",X"ED",X"98",
		X"09",X"DE",X"43",X"11",X"DF",X"43",X"01",X"05",X"00",X"5F",X"ED",X"98",X"AF",X"1A",X"CC",X"43",
		X"1A",X"DE",X"43",X"AF",X"1A",X"FF",X"64",X"1A",X"01",X"65",X"1A",X"03",X"65",X"1A",X"00",X"65",
		X"1A",X"02",X"65",X"1A",X"04",X"65",X"E5",X"ED",X"1A",X"E5",X"FA",X"1A",X"09",X"97",X"64",X"E3",
		X"E6",X"09",X"96",X"64",X"E3",X"4E",X"28",X"02",X"30",X"32",X"3E",X"00",X"1A",X"03",X"50",X"E5",
		X"44",X"15",X"11",X"50",X"41",X"09",X"EB",X"30",X"3E",X"01",X"06",X"25",X"E5",X"D5",X"15",X"3E",
		X"03",X"E5",X"67",X"15",X"09",X"96",X"64",X"E3",X"EE",X"3A",X"8E",X"64",X"3D",X"1A",X"8E",X"64",
		X"3E",X"40",X"09",X"16",X"40",X"11",X"17",X"40",X"01",X"20",X"00",X"5F",X"ED",X"98",X"E5",X"13",
		X"00",X"3A",X"FF",X"64",X"1A",X"03",X"65",X"3A",X"00",X"65",X"1A",X"04",X"65",X"E5",X"39",X"1B",
		X"C3",X"B3",X"23",X"09",X"96",X"64",X"E3",X"4E",X"08",X"E2",X"E3",X"6E",X"28",X"AC",X"3A",X"96",
		X"64",X"E3",X"7F",X"08",X"43",X"E5",X"44",X"15",X"11",X"50",X"41",X"09",X"F8",X"30",X"3E",X"01",
		X"06",X"25",X"E5",X"D5",X"15",X"3E",X"03",X"E5",X"67",X"15",X"09",X"96",X"64",X"E3",X"AE",X"3A",
		X"8F",X"64",X"3D",X"1A",X"8F",X"64",X"3E",X"40",X"09",X"02",X"40",X"11",X"03",X"40",X"01",X"20",
		X"00",X"5F",X"ED",X"98",X"E5",X"0C",X"00",X"3A",X"01",X"65",X"1A",X"03",X"65",X"3A",X"02",X"65",
		X"1A",X"04",X"65",X"E5",X"3B",X"1B",X"30",X"1B",X"3E",X"01",X"1A",X"03",X"50",X"30",X"9E",X"E5",
		X"44",X"15",X"09",X"96",X"64",X"E3",X"4E",X"C2",X"E9",X"22",X"11",X"10",X"41",X"09",X"05",X"31",
		X"3E",X"01",X"06",X"11",X"E5",X"D5",X"15",X"09",X"08",X"65",X"E3",X"C6",X"3E",X"01",X"E5",X"67",
		X"15",X"09",X"96",X"64",X"E3",X"6E",X"28",X"8F",X"C3",X"E9",X"22",X"E5",X"FA",X"26",X"09",X"97",
		X"64",X"E3",X"66",X"28",X"13",X"E3",X"A6",X"09",X"C2",X"65",X"E3",X"C6",X"1A",X"C0",X"50",X"3A",
		X"C2",X"65",X"FE",X"00",X"08",X"DE",X"30",X"05",X"3E",X"02",X"E5",X"67",X"15",X"09",X"8F",X"65",
		X"E3",X"C6",X"09",X"59",X"65",X"E3",X"C6",X"E5",X"BC",X"33",X"ED",X"73",X"AE",X"64",X"7B",X"9A",
		X"28",X"21",X"09",X"00",X"00",X"0A",X"AE",X"64",X"E5",X"4E",X"27",X"1A",X"C0",X"50",X"E5",X"15",
		X"16",X"09",X"96",X"64",X"E3",X"66",X"28",X"F7",X"E3",X"A6",X"E5",X"22",X"16",X"09",X"96",X"64",
		X"E3",X"56",X"08",X"27",X"E5",X"3F",X"1B",X"E5",X"22",X"16",X"09",X"96",X"64",X"E3",X"76",X"08",
		X"21",X"30",X"4F",X"E3",X"96",X"E5",X"3E",X"1B",X"30",X"EA",X"E3",X"B6",X"09",X"97",X"64",X"E3",
		X"E6",X"09",X"96",X"64",X"E3",X"6E",X"08",X"29",X"3A",X"01",X"65",X"3C",X"FE",X"24",X"08",X"02",
		X"3E",X"23",X"1A",X"01",X"65",X"1A",X"03",X"65",X"3A",X"02",X"65",X"3C",X"FE",X"31",X"08",X"02",
		X"3E",X"30",X"1A",X"02",X"65",X"1A",X"04",X"65",X"E5",X"40",X"1B",X"E5",X"3D",X"1B",X"C3",X"B3",
		X"23",X"3A",X"FF",X"64",X"3C",X"FE",X"24",X"08",X"02",X"3E",X"23",X"1A",X"FF",X"64",X"1A",X"03",
		X"65",X"3A",X"00",X"65",X"3C",X"FE",X"31",X"08",X"02",X"3E",X"30",X"1A",X"00",X"65",X"1A",X"04",
		X"65",X"E5",X"40",X"1B",X"E5",X"3C",X"1B",X"C3",X"B3",X"23",X"3A",X"98",X"64",X"FE",X"00",X"08",
		X"2E",X"09",X"96",X"64",X"E3",X"6E",X"08",X"2F",X"3A",X"8F",X"64",X"FE",X"00",X"08",X"66",X"E5",
		X"44",X"15",X"11",X"90",X"41",X"09",X"16",X"31",X"3E",X"01",X"06",X"21",X"E5",X"D5",X"15",X"3E",
		X"02",X"E5",X"67",X"15",X"E5",X"EE",X"11",X"09",X"95",X"64",X"E3",X"DE",X"C3",X"79",X"07",X"D6",
		X"01",X"1A",X"98",X"64",X"C3",X"6F",X"23",X"3A",X"8E",X"64",X"FE",X"00",X"08",X"0D",X"09",X"96",
		X"64",X"E3",X"4E",X"08",X"E2",X"E5",X"44",X"15",X"11",X"D8",X"40",X"09",X"37",X"31",X"3E",X"01",
		X"06",X"14",X"E5",X"D5",X"15",X"3E",X"03",X"E5",X"67",X"15",X"C3",X"36",X"23",X"E5",X"3A",X"1B",
		X"C3",X"13",X"23",X"E5",X"38",X"1B",X"C3",X"13",X"23",X"2A",X"91",X"64",X"EB",X"F5",X"09",X"00",
		X"00",X"F5",X"31",X"F5",X"7E",X"01",X"F5",X"86",X"02",X"47",X"CE",X"27",X"F5",X"5F",X"02",X"E3",
		X"38",X"E3",X"38",X"E3",X"38",X"E3",X"38",X"F5",X"7E",X"00",X"09",X"07",X"25",X"E3",X"0F",X"E5",
		X"98",X"15",X"76",X"0B",X"56",X"EB",X"E9",X"13",X"25",X"13",X"25",X"14",X"25",X"34",X"25",X"0C",
		X"25",X"2C",X"25",X"E1",X"F5",X"7E",X"04",X"90",X"F5",X"5F",X"04",X"E1",X"F5",X"7E",X"04",X"80",
		X"F5",X"5F",X"04",X"E1",X"F5",X"7E",X"03",X"80",X"F5",X"5F",X"03",X"E1",X"F5",X"7E",X"03",X"90",
		X"F5",X"5F",X"03",X"E1",X"2A",X"76",X"64",X"EB",X"F5",X"09",X"00",X"00",X"F5",X"31",X"EB",X"01",
		X"00",X"64",X"1F",X"3F",X"ED",X"42",X"CD",X"F5",X"7E",X"00",X"09",X"57",X"25",X"E3",X"0F",X"E5",
		X"98",X"15",X"76",X"0B",X"56",X"EB",X"E9",X"0F",X"26",X"4B",X"25",X"8E",X"25",X"1E",X"26",X"40",
		X"26",X"53",X"26",X"F5",X"7E",X"03",X"1A",X"74",X"64",X"F5",X"7E",X"04",X"1A",X"75",X"64",X"E5",
		X"BD",X"26",X"F5",X"7E",X"06",X"12",X"3A",X"22",X"64",X"FE",X"00",X"08",X"17",X"3A",X"23",X"64",
		X"FE",X"00",X"08",X"17",X"C1",X"09",X"24",X"64",X"21",X"CD",X"D1",X"13",X"01",X"05",X"00",X"1E",
		X"FF",X"ED",X"98",X"E1",X"F5",X"7E",X"06",X"13",X"12",X"30",X"E9",X"F5",X"7E",X"06",X"09",X"08",
		X"00",X"31",X"EB",X"12",X"30",X"F6",X"E5",X"CD",X"26",X"F5",X"7E",X"03",X"90",X"1A",X"74",X"64",
		X"F5",X"7E",X"04",X"1A",X"75",X"64",X"E5",X"BD",X"26",X"3A",X"22",X"64",X"FE",X"00",X"28",X"1A",
		X"3A",X"22",X"64",X"E3",X"0F",X"F5",X"46",X"05",X"80",X"3D",X"C1",X"FD",X"09",X"24",X"64",X"FD",
		X"21",X"FD",X"5B",X"00",X"FD",X"5A",X"01",X"FD",X"5F",X"02",X"3C",X"13",X"FD",X"5B",X"03",X"FD",
		X"5A",X"04",X"FD",X"5F",X"05",X"3A",X"74",X"64",X"F5",X"5F",X"03",X"3A",X"75",X"64",X"F5",X"5F",
		X"04",X"E1",X"3A",X"23",X"64",X"FE",X"00",X"E2",X"74",X"26",X"3A",X"23",X"64",X"E3",X"0F",X"C6",
		X"27",X"F5",X"46",X"05",X"80",X"C1",X"FD",X"09",X"24",X"64",X"FD",X"21",X"FD",X"5B",X"00",X"FD",
		X"5A",X"01",X"FD",X"5F",X"02",X"3C",X"09",X"08",X"00",X"31",X"EB",X"FD",X"5B",X"03",X"FD",X"5A",
		X"04",X"FD",X"5F",X"05",X"C3",X"CD",X"25",X"F5",X"7E",X"03",X"1A",X"74",X"64",X"F5",X"7E",X"04",
		X"1A",X"75",X"64",X"C3",X"9E",X"25",X"E5",X"CD",X"26",X"F5",X"7E",X"03",X"80",X"C3",X"AD",X"25",
		X"E5",X"CD",X"26",X"F5",X"7E",X"04",X"90",X"1A",X"75",X"64",X"F5",X"7E",X"03",X"1A",X"74",X"64",
		X"C3",X"9E",X"25",X"E5",X"CD",X"26",X"F5",X"7E",X"04",X"80",X"30",X"EB",X"F5",X"7E",X"05",X"C1",
		X"FD",X"09",X"24",X"64",X"FD",X"21",X"FD",X"5B",X"00",X"FD",X"5A",X"01",X"FD",X"5F",X"02",X"3A",
		X"74",X"64",X"F5",X"5F",X"03",X"3A",X"75",X"64",X"F5",X"5F",X"04",X"F5",X"7E",X"00",X"09",X"90",
		X"26",X"E3",X"0F",X"E5",X"98",X"15",X"D5",X"76",X"0B",X"56",X"EB",X"D1",X"F5",X"7E",X"06",X"E9",
		X"B4",X"26",X"B4",X"26",X"B5",X"26",X"A8",X"26",X"AB",X"26",X"9A",X"26",X"E1",X"13",X"FD",X"5B",
		X"03",X"FD",X"5A",X"04",X"FD",X"5F",X"05",X"E1",X"33",X"30",X"DB",X"09",X"08",X"00",X"31",X"EB",
		X"30",X"EC",X"EB",X"11",X"08",X"00",X"1F",X"3F",X"ED",X"52",X"EB",X"30",X"C9",X"3A",X"74",X"64",
		X"CE",X"07",X"1A",X"22",X"64",X"3A",X"75",X"64",X"CE",X"07",X"1A",X"23",X"64",X"3A",X"74",X"64",
		X"E3",X"3F",X"E3",X"3F",X"E3",X"3F",X"57",X"3A",X"75",X"64",X"E3",X"3F",X"E3",X"3F",X"E3",X"3F",
		X"77",X"E5",X"F7",X"14",X"E1",X"F5",X"7E",X"01",X"F5",X"86",X"02",X"47",X"CE",X"27",X"F5",X"5F",
		X"02",X"E3",X"38",X"E3",X"38",X"E3",X"38",X"E3",X"38",X"E1",X"3A",X"03",X"65",X"09",X"20",X"27",
		X"E3",X"0F",X"E3",X"0F",X"E5",X"98",X"15",X"E9",X"E5",X"12",X"0F",X"E1",X"E5",X"64",X"0F",X"E1",
		X"E5",X"86",X"0F",X"E1",X"E5",X"C0",X"0F",X"E1",X"E5",X"FA",X"0F",X"E1",X"E5",X"1C",X"28",X"E1",
		X"E5",X"6E",X"28",X"E1",X"E5",X"A8",X"28",X"E1",X"E5",X"CA",X"28",X"E1",X"E5",X"34",X"29",X"E1",
		X"E5",X"56",X"29",X"E1",X"E5",X"90",X"29",X"E1",X"E5",X"E2",X"29",X"E1",X"E5",X"E3",X"29",X"E1",
		X"E5",X"E4",X"29",X"E1",X"E5",X"E5",X"29",X"E1",X"D5",X"1F",X"3F",X"09",X"26",X"01",X"16",X"00",
		X"ED",X"52",X"7D",X"1F",X"3F",X"09",X"10",X"01",X"D1",X"72",X"16",X"00",X"ED",X"52",X"55",X"77",
		X"E1",X"7D",X"EE",X"03",X"6F",X"E1",X"09",X"96",X"64",X"E3",X"46",X"E0",X"E3",X"6E",X"28",X"43",
		X"09",X"A8",X"64",X"7B",X"86",X"0F",X"5F",X"0B",X"7A",X"A6",X"0F",X"5F",X"0B",X"3E",X"00",X"A6",
		X"0F",X"5F",X"38",X"02",X"30",X"1A",X"09",X"96",X"64",X"E3",X"6E",X"28",X"13",X"09",X"DE",X"43",
		X"11",X"DF",X"43",X"01",X"05",X"00",X"1E",X"40",X"ED",X"98",X"AF",X"1A",X"DE",X"43",X"30",X"30",
		X"09",X"CC",X"43",X"11",X"CD",X"43",X"01",X"05",X"00",X"1E",X"40",X"ED",X"98",X"AF",X"1A",X"CC",
		X"43",X"30",X"05",X"09",X"AB",X"64",X"30",X"BB",X"09",X"96",X"64",X"E3",X"6E",X"28",X"74",X"09",
		X"AA",X"64",X"11",X"FB",X"43",X"3A",X"99",X"64",X"DD",X"E5",X"0E",X"10",X"0B",X"0B",X"0B",X"EB",
		X"2A",X"8B",X"64",X"D9",X"FE",X"04",X"D0",X"E3",X"0F",X"E3",X"0F",X"3C",X"3C",X"E5",X"98",X"15",
		X"E5",X"AA",X"11",X"D0",X"3A",X"98",X"64",X"3C",X"1A",X"98",X"64",X"09",X"08",X"65",X"E3",X"C6",
		X"09",X"96",X"64",X"E3",X"6E",X"28",X"12",X"3A",X"99",X"64",X"3C",X"1A",X"99",X"64",X"3A",X"8E",
		X"DB",X"09",X"06",X"50",X"AF",X"00",X"20",X"5F",X"0B",X"56",X"FC",X"D9",X"40",X"49",X"BD",X"37",
		X"93",X"8E",X"02",X"FE",X"97",X"34",X"6A",X"00",X"B0",X"09",X"6E",X"10",X"17",X"65",X"60",X"5F",
		X"2B",X"6A",X"FC",X"34",X"40",X"8F",X"B1",X"FE",X"00",X"60",X"17",X"02",X"B0",X"09",X"6E",X"10",
		X"5F",X"B1",X"40",X"00",X"0B",X"9B",X"FC",X"00",X"20",X"FD",X"F5",X"AF",X"F1",X"9D",X"9D",X"4A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"63",X"00",X"00",X"00",X"FF",X"00",X"63",X"00",X"9C",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"63",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"9C",X"00",X"63",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"41",X"00",X"63",X"00",X"41",X"00",X"63",X"00",X"88",X"00",X"9C",X"00",X"88",X"00",X"9C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"36",X"00",X"9C",X"00",X"36",X"00",X"9C",X"00",X"36",X"00",X"63",X"00",X"36",X"00",X"63",X"00",
		X"00",X"00",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"00",X"00",X"40",X"00",X"40",X"00",X"40",
		X"00",X"F0",X"00",X"F0",X"00",X"F0",X"60",X"F0",X"00",X"76",X"00",X"F0",X"00",X"F0",X"22",X"62",
		X"80",X"00",X"80",X"00",X"80",X"00",X"00",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"00",X"00",
		X"F0",X"60",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"76",X"90",X"F0",X"00",X"F0",X"00",X"F0",X"00",
		X"00",X"00",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"00",X"00",X"40",X"00",X"40",X"00",X"40",
		X"00",X"F0",X"00",X"F0",X"00",X"F0",X"60",X"F0",X"00",X"F0",X"00",X"B6",X"00",X"94",X"90",X"F0",
		X"80",X"00",X"80",X"00",X"80",X"00",X"00",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"00",X"00",
		X"F0",X"60",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"90",X"B6",X"00",X"94",X"00",X"F0",X"00",
		X"00",X"00",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"00",X"00",X"40",X"00",X"40",X"00",X"40",
		X"00",X"F0",X"00",X"F0",X"00",X"F0",X"60",X"F0",X"00",X"F0",X"00",X"76",X"00",X"62",X"90",X"F0",
		X"80",X"00",X"80",X"00",X"80",X"00",X"00",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"00",X"00",
		X"F0",X"60",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"90",X"62",X"00",X"76",X"00",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"41",X"00",X"00",X"00",X"63",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"9C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"63",X"00",X"00",X"00",X"41",X"00",X"00",X"00",X"9C",X"00",X"00",X"00",X"88",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"41",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"41",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"70",X"00",X"10",X"00",X"70",X"90",X"F3",X"90",X"F1",X"90",X"F3",X"B2",X"F0",
		X"00",X"63",X"00",X"FE",X"00",X"FF",X"41",X"F0",X"00",X"F0",X"00",X"E0",X"00",X"F0",X"90",X"E0",
		X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"40",X"B0",X"70",X"90",X"60",X"90",X"F0",X"90",
		X"70",X"40",X"F0",X"00",X"70",X"00",X"F0",X"00",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"B2",X"F0",X"F1",X"F0",X"F3",X"F0",X"F0",X"F0",
		X"41",X"F0",X"FE",X"70",X"63",X"70",X"F0",X"70",X"F0",X"E0",X"E0",X"F0",X"F0",X"F0",X"E0",X"F0",
		X"70",X"00",X"10",X"00",X"70",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"70",X"70",X"70",X"10",X"70",X"70",X"70",X"00",X"F0",X"90",X"F0",X"00",X"F0",X"00",X"F0",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"B0",X"00",X"20",X"00",X"B0",
		X"00",X"F0",X"00",X"F0",X"00",X"F0",X"60",X"F0",X"00",X"B0",X"B0",X"B0",X"20",X"B0",X"B0",X"B0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"B0",X"B0",X"B0",X"B0",X"B0",X"B0",X"B0",X"B0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"B0",X"B0",X"B0",X"B0",X"B0",X"B0",X"B0",X"B0",
		X"78",X"6C",X"4E",X"F0",X"6C",X"78",X"6C",X"F0",X"B0",X"B0",X"B0",X"B0",X"B0",X"B0",X"B0",X"B0",
		X"F0",X"F0",X"F0",X"B1",X"F0",X"F0",X"F0",X"B1",X"B1",X"0F",X"87",X"0F",X"93",X"0F",X"87",X"0E",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"B0",X"03",X"20",X"0F",X"B0",X"0F",X"01",X"0E",
		X"93",X"6C",X"0F",X"00",X"87",X"08",X"4E",X"00",X"2C",X"B0",X"B0",X"20",X"38",X"B0",X"B0",X"00",
		X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"01",X"00",X"03",X"00",X"03",X"00",X"03",
		X"00",X"0E",X"00",X"0F",X"00",X"0E",X"06",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"70",X"00",X"10",X"00",X"70",X"90",X"F0",X"40",X"F0",X"F0",X"90",X"F0",X"F0",
		X"00",X"70",X"70",X"40",X"10",X"70",X"70",X"00",X"00",X"90",X"00",X"90",X"00",X"00",X"90",X"D0",
		X"70",X"40",X"60",X"00",X"00",X"60",X"60",X"40",X"00",X"F0",X"10",X"F3",X"F0",X"F1",X"F0",X"B2",
		X"00",X"F0",X"70",X"63",X"30",X"FE",X"F0",X"41",X"70",X"80",X"F0",X"F0",X"70",X"80",X"00",X"F0",
		X"70",X"40",X"70",X"70",X"60",X"60",X"00",X"70",X"90",X"F0",X"90",X"60",X"90",X"70",X"0E",X"40",
		X"00",X"F0",X"00",X"F0",X"00",X"F0",X"40",X"F0",X"F0",X"F0",X"B0",X"B0",X"B0",X"B0",X"90",X"A0",
		X"50",X"00",X"10",X"00",X"50",X"00",X"00",X"00",X"F0",X"B2",X"F3",X"90",X"F1",X"90",X"F3",X"00",
		X"F0",X"41",X"FF",X"00",X"FE",X"00",X"63",X"00",X"E0",X"90",X"F0",X"00",X"E0",X"00",X"F0",X"00",
		X"D0",X"F0",X"F0",X"F0",X"F0",X"90",X"60",X"60",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"D0",
		X"00",X"B0",X"00",X"F0",X"00",X"90",X"60",X"F0",X"00",X"00",X"F0",X"F0",X"60",X"60",X"90",X"F0",
		X"60",X"C0",X"B0",X"F0",X"F0",X"B0",X"40",X"F0",X"00",X"60",X"90",X"F0",X"F0",X"B0",X"F0",X"B0",
		X"60",X"F0",X"00",X"F0",X"F0",X"90",X"F0",X"00",X"B0",X"F0",X"F0",X"60",X"00",X"F0",X"B0",X"00",
		X"60",X"70",X"00",X"F0",X"40",X"60",X"F0",X"F0",X"60",X"B0",X"F0",X"40",X"F0",X"F0",X"00",X"B0",
		X"F0",X"60",X"F0",X"B0",X"80",X"80",X"70",X"70",X"00",X"80",X"00",X"00",X"00",X"00",X"80",X"F0",
		X"00",X"60",X"B0",X"90",X"90",X"F0",X"F0",X"90",X"70",X"00",X"60",X"00",X"90",X"00",X"00",X"00",
		X"C0",X"60",X"F0",X"00",X"B0",X"00",X"40",X"00",X"F0",X"90",X"B0",X"60",X"70",X"F0",X"F0",X"00",
		X"00",X"88",X"88",X"9C",X"00",X"9C",X"88",X"9C",X"00",X"41",X"41",X"63",X"00",X"63",X"41",X"63",
		X"FB",X"FC",X"FB",X"FC",X"F8",X"FB",X"FF",X"FF",X"FB",X"F3",X"FF",X"F3",X"F1",X"FD",X"FF",X"FF",
		X"9C",X"88",X"88",X"00",X"9C",X"00",X"88",X"00",X"63",X"41",X"41",X"00",X"63",X"00",X"41",X"00",
		X"FC",X"FC",X"FC",X"FC",X"FB",X"FB",X"FF",X"00",X"F3",X"F3",X"F3",X"F3",X"FD",X"FD",X"FF",X"00",
		X"00",X"88",X"88",X"9C",X"00",X"9C",X"88",X"9C",X"00",X"41",X"41",X"63",X"00",X"63",X"41",X"63",
		X"F9",X"FF",X"FB",X"FB",X"FA",X"FC",X"FB",X"FC",X"FB",X"FF",X"F5",X"FD",X"FD",X"F3",X"FB",X"F3",
		X"9C",X"88",X"9C",X"00",X"9C",X"88",X"88",X"00",X"63",X"41",X"63",X"00",X"63",X"41",X"41",X"00",
		X"FF",X"FF",X"FB",X"FB",X"FC",X"FC",X"FC",X"FC",X"FF",X"FF",X"FD",X"FD",X"F3",X"F3",X"F3",X"F3",
		X"00",X"88",X"88",X"9C",X"00",X"9C",X"88",X"9C",X"00",X"41",X"41",X"63",X"00",X"63",X"41",X"63",
		X"FF",X"FE",X"FE",X"FB",X"FE",X"FC",X"F8",X"FC",X"FF",X"FF",X"FB",X"FD",X"F7",X"F3",X"F1",X"F3",
		X"9C",X"88",X"9C",X"00",X"9C",X"88",X"88",X"00",X"63",X"41",X"63",X"00",X"63",X"41",X"41",X"00",
		X"FF",X"FF",X"FB",X"FB",X"FC",X"FC",X"FC",X"FC",X"FF",X"FF",X"FD",X"FD",X"F3",X"F3",X"F3",X"F3",
		X"00",X"88",X"88",X"9C",X"00",X"9C",X"88",X"9C",X"00",X"41",X"41",X"63",X"00",X"63",X"41",X"63",
		X"FC",X"FF",X"FB",X"FB",X"FB",X"FC",X"FC",X"FC",X"FB",X"FF",X"F5",X"FD",X"F5",X"F3",X"FB",X"F3",
		X"9C",X"88",X"9C",X"00",X"9C",X"88",X"88",X"00",X"63",X"41",X"63",X"00",X"63",X"41",X"41",X"00",
		X"FF",X"FF",X"FB",X"FB",X"FC",X"FC",X"FC",X"FC",X"FF",X"FF",X"FD",X"FD",X"F3",X"F3",X"F3",X"F3",
		X"1D",X"1E",X"20",X"2C",X"52",X"54",X"54",X"13",X"1F",X"19",X"59",X"18",X"50",X"17",X"52",X"54",
		X"20",X"63",X"69",X"15",X"61",X"54",X"68",X"1C",X"1B",X"1E",X"20",X"20",X"1F",X"13",X"19",X"B3",
		X"B7",X"D8",X"7E",X"7B",X"20",X"57",X"9E",X"9E",X"D8",X"B3",X"B0",X"20",X"EA",X"97",X"20",X"7B",
		X"B1",X"54",X"52",X"54",X"35",X"36",X"08",X"2C",X"13",X"52",X"50",X"17",X"37",X"31",X"71",X"30",
		X"54",X"68",X"49",X"54",X"08",X"4B",X"69",X"15",X"34",X"31",X"37",X"13",X"33",X"36",X"08",X"4A",
		X"90",X"10",X"09",X"01",X"50",X"41",X"00",X"10",X"01",X"10",X"07",X"C8",X"FE",X"BD",X"4E",X"4A",
		X"90",X"34",X"09",X"01",X"50",X"41",X"00",X"34",X"01",X"00",X"03",X"C8",X"FE",X"BD",X"4E",X"4A",
		X"90",X"50",X"09",X"19",X"50",X"41",X"18",X"50",X"01",X"00",X"00",X"C8",X"27",X"BD",X"4E",X"4A",
		X"90",X"37",X"09",X"D9",X"50",X"41",X"D8",X"37",X"01",X"00",X"00",X"C8",X"27",X"BD",X"4E",X"4A",
		X"90",X"50",X"09",X"11",X"50",X"41",X"10",X"50",X"01",X"00",X"00",X"C8",X"67",X"BD",X"4E",X"09",
		X"24",X"34",X"41",X"37",X"34",X"01",X"25",X"00",X"4E",X"09",X"BD",X"68",X"FF",X"7B",X"C8",X"0A",
		X"C3",X"50",X"6A",X"9E",X"34",X"17",X"80",X"03",X"4A",X"E4",X"34",X"B5",X"E3",X"63",X"09",X"C8",
		X"45",X"34",X"4A",X"9E",X"7E",X"78",X"E4",X"24",X"B3",X"09",X"B3",X"68",X"6F",X"5F",X"6F",X"B5",
		X"C8",X"8A",X"7E",X"78",X"45",X"34",X"4A",X"9E",X"48",X"B5",X"4F",X"45",X"09",X"C8",X"68",X"0A",
		X"8B",X"48",X"78",X"6F",X"34",X"B3",X"9E",X"B3",X"6F",X"6F",X"6F",X"8D",X"B3",X"4A",X"B3",X"34",
		X"78",X"05",X"5F",X"C6",X"B3",X"09",X"08",X"34",X"B3",X"01",X"FB",X"00",X"FE",X"4A",X"6E",X"50",
		X"B5",X"92",X"4A",X"41",X"BB",X"13",X"09",X"93",X"13",X"4E",X"6C",X"BD",X"01",X"10",X"00",X"C8",
		X"09",X"93",X"17",X"01",X"92",X"17",X"41",X"64",X"00",X"C8",X"05",X"90",X"4E",X"4A",X"BD",X"50",
		X"09",X"9B",X"17",X"01",X"9A",X"17",X"41",X"64",X"00",X"C8",X"21",X"90",X"4E",X"4A",X"BD",X"50",
		X"09",X"93",X"60",X"01",X"A3",X"13",X"41",X"62",X"00",X"4A",X"C8",X"13",X"BD",X"9C",X"AF",X"4A",
		X"BD",X"13",X"4A",X"C0",X"13",X"09",X"DE",X"68",X"41",X"6C",X"34",X"BD",X"CB",X"00",X"01",X"C8",
		X"09",X"DA",X"34",X"B5",X"E8",X"13",X"41",X"0E",X"40",X"41",X"02",X"10",X"09",X"03",X"10",X"01",
		X"6C",X"BD",X"4E",X"4A",X"00",X"C8",X"10",X"90",X"50",X"41",X"02",X"14",X"09",X"03",X"14",X"01",
		X"64",X"BD",X"4E",X"09",X"00",X"C8",X"21",X"0A",X"14",X"01",X"0B",X"00",X"41",X"64",X"14",X"4E",
		X"41",X"90",X"C8",X"09",X"BD",X"50",X"4A",X"8D",X"60",X"01",X"27",X"00",X"41",X"06",X"10",X"BD",
		X"C8",X"10",X"4A",X"E3",X"AF",X"6A",X"24",X"34",X"FE",X"09",X"08",X"60",X"00",X"AB",X"23",X"41",
		X"24",X"00",X"01",X"C8",X"10",X"BD",X"21",X"4A",X"90",X"35",X"09",X"06",X"50",X"41",X"05",X"35",
		X"01",X"00",X"00",X"C8",X"FF",X"BD",X"4E",X"09",X"12",X"35",X"0A",X"06",X"4C",X"0A",X"66",X"35",
		X"09",X"25",X"35",X"09",X"65",X"35",X"0A",X"58",X"4C",X"0A",X"69",X"35",X"0A",X"09",X"35",X"09",
		X"68",X"35",X"0A",X"87",X"35",X"09",X"28",X"4C",X"0A",X"6C",X"35",X"09",X"54",X"35",X"0A",X"53",
		X"35",X"09",X"13",X"4C",X"0A",X"E9",X"35",X"0A",X"3F",X"35",X"0A",X"3E",X"35",X"09",X"57",X"35",
		X"0A",X"1E",X"35",X"0A",X"76",X"4D",X"09",X"A2",X"35",X"09",X"5A",X"35",X"0A",X"A1",X"35",X"0A",
		X"79",X"4D",X"09",X"8D",X"35",X"0A",X"E0",X"35",X"0A",X"8C",X"35",X"0A",X"A5",X"35",X"09",X"C4",
		X"35",X"0A",X"D2",X"35",X"09",X"90",X"4E",X"0A",X"A8",X"35",X"09",X"AF",X"35",X"0A",X"EF",X"35",
		X"09",X"F3",X"4E",X"0A",X"9F",X"35",X"0A",X"93",X"35",X"0A",X"F2",X"35",X"09",X"B2",X"35",X"06",
		X"08",X"4E",X"10",X"0B",X"09",X"00",X"50",X"40",X"FB",X"03",X"00",X"09",X"6E",X"50",X"4A",X"C6",
		X"34",X"E3",X"BE",X"FE",X"B3",X"34",X"6A",X"00",X"B2",X"E2",X"21",X"FE",X"69",X"34",X"6A",X"00",
		X"92",X"C5",X"21",X"B3",X"69",X"34",X"09",X"8E",X"AF",X"09",X"01",X"34",X"4A",X"C6",X"50",X"B3",
		X"86",X"4A",X"22",X"50",X"B5",X"90",X"46",X"B5",X"E8",X"B5",X"6E",X"45",X"48",X"37",X"01",X"09",
		X"C5",X"92",X"B3",X"21",X"34",X"69",X"3E",X"B5",X"7C",X"B5",X"6E",X"45",X"40",X"37",X"07",X"09",
		X"C5",X"92",X"B3",X"21",X"34",X"69",X"3E",X"6E",X"10",X"41",X"FD",X"14",X"B5",X"14",X"44",X"09",
		X"B4",X"06",X"6E",X"B5",X"68",X"64",X"01",X"BB",X"45",X"09",X"31",X"68",X"41",X"B6",X"14",X"6E",
		X"03",X"BB",X"64",X"41",X"06",X"45",X"B5",X"50",X"14",X"6E",X"B5",X"06",X"09",X"03",X"68",X"64",
		X"B5",X"70",X"45",X"09",X"BB",X"14",X"41",X"B6",X"68",X"64",X"03",X"BB",X"6E",X"B5",X"06",X"45",
		X"41",X"B7",X"14",X"6E",X"73",X"68",X"09",X"03",X"06",X"45",X"B5",X"94",X"64",X"41",X"BB",X"10",
		X"09",X"01",X"61",X"44",X"C6",X"06",X"6E",X"B5",X"D5",X"10",X"41",X"AB",X"45",X"09",X"B1",X"61",
		X"6E",X"B5",X"06",X"45",X"01",X"D5",X"44",X"41",X"A3",X"61",X"09",X"01",X"10",X"6E",X"EF",X"06",
		X"60",X"41",X"D5",X"10",X"B5",X"C8",X"45",X"09",X"D7",X"06",X"6E",X"B5",X"61",X"46",X"01",X"D5",
		X"45",X"09",X"52",X"61",X"41",X"BD",X"11",X"6E",X"01",X"D5",X"24",X"6A",X"06",X"45",X"B5",X"E3",
		X"34",X"27",X"01",X"61",X"FE",X"41",X"08",X"11",X"09",X"01",X"61",X"27",X"F9",X"06",X"6E",X"B5",
		X"D5",X"FE",X"60",X"08",X"45",X"02",X"08",X"27",X"41",X"20",X"11",X"6E",X"61",X"62",X"09",X"01",
		X"06",X"45",X"B5",X"25",X"27",X"60",X"D5",X"41",X"61",X"62",X"09",X"01",X"11",X"6E",X"47",X"06",
		X"27",X"41",X"D5",X"10",X"B5",X"E4",X"45",X"09",X"0E",X"06",X"6E",X"B5",X"62",X"61",X"01",X"D5",
		X"45",X"FE",X"8D",X"08",X"6A",X"00",X"34",X"27",X"41",X"6F",X"11",X"6E",X"7C",X"62",X"09",X"01",
		X"06",X"45",X"B5",X"4B",X"06",X"60",X"D5",X"FE",X"01",X"7C",X"27",X"09",X"08",X"11",X"41",X"15",
		X"62",X"06",X"01",X"D5",X"6E",X"B5",X"06",X"45",X"60",X"08",X"FE",X"41",X"08",X"27",X"02",X"7C",
		X"11",X"6E",X"33",X"06",X"09",X"01",X"62",X"06",X"B5",X"25",X"45",X"7C",X"D5",X"41",X"60",X"11",
		X"09",X"01",X"62",X"06",X"51",X"06",X"6E",X"B5",X"D5",X"B5",X"6E",X"45",X"45",X"37",X"04",X"09",
		X"C5",X"08",X"B3",X"B5",X"34",X"53",X"3E",X"BC",X"4A",X"34",X"4A",X"01",X"AF",X"4A",X"FF",X"35",
		X"4A",X"00",X"35",X"4A",X"03",X"35",X"4A",X"02",X"35",X"B5",X"04",X"4A",X"4A",X"BE",X"35",X"B5",
		X"FA",X"4A",X"B5",X"EC",X"26",X"B5",X"FB",X"63",X"AF",X"4A",X"08",X"35",X"4A",X"6B",X"35",X"4A",
		X"56",X"35",X"4A",X"A4",X"35",X"4A",X"59",X"35",X"4A",X"92",X"35",X"B5",X"8F",X"35",X"4A",X"45",
		X"46",X"09",X"90",X"34",X"4A",X"C5",X"50",X"B3",X"3E",X"C6",X"26",X"B3",X"08",X"34",X"09",X"36",
		X"08",X"B3",X"60",X"93",X"02",X"A6",X"B6",X"89",X"07",X"09",X"22",X"34",X"B5",X"C5",X"46",X"B3",
		X"9E",X"C6",X"AE",X"B3",X"B3",X"34",X"09",X"A6",X"B3",X"09",X"B3",X"34",X"C6",X"C7",X"E6",X"B3",
		X"C6",X"B3",X"C6",X"09",X"09",X"96",X"34",X"24",X"34",X"01",X"25",X"00",X"41",X"37",X"34",X"4E",
		X"FF",X"FF",X"C8",X"01",X"BD",X"4A",X"6E",X"50",X"09",X"56",X"34",X"27",X"C7",X"08",X"B3",X"6A",
		X"FD",X"FD",X"6C",X"FE",X"34",X"34",X"4A",X"44",X"08",X"B3",X"B3",X"00",X"04",X"F6",X"D6",X"4A",
		X"90",X"B5",X"6E",X"44",X"50",X"FD",X"10",X"6E",X"03",X"6A",X"25",X"34",X"B5",X"E3",X"45",X"FE",
		X"00",X"6A",X"44",X"34",X"B2",X"E2",X"22",X"FE",X"02",X"58",X"34",X"09",X"48",X"11",X"41",X"CC",
		X"60",X"23",X"01",X"D5",X"6E",X"B5",X"06",X"45",X"6A",X"3F",X"50",X"5C",X"10",X"08",X"B3",X"6A",
		X"E3",X"28",X"FE",X"6A",X"34",X"45",X"00",X"E2",X"34",X"1E",X"02",X"02",X"FE",X"D6",X"68",X"4A",
		X"E2",X"34",X"6A",X"01",X"34",X"D6",X"E5",X"0F",X"4A",X"C6",X"34",X"B3",X"E5",X"34",X"09",X"9E",
		X"6A",X"8E",X"34",X"B5",X"8A",X"34",X"4A",X"43",X"00",X"FE",X"E3",X"B2",X"6A",X"00",X"34",X"3F",
		X"22",X"93",X"65",X"22",X"B5",X"3F",X"45",X"FE",X"04",X"26",X"29",X"09",X"48",X"11",X"41",X"EF",
		X"60",X"41",X"01",X"D5",X"6E",X"B5",X"06",X"45",X"41",X"D0",X"12",X"6E",X"40",X"60",X"09",X"01",
		X"06",X"45",X"B5",X"5A",X"02",X"41",X"D5",X"11",X"09",X"01",X"60",X"23",X"CC",X"06",X"6E",X"B5",
		X"D5",X"41",X"60",X"10",X"45",X"C0",X"C4",X"09",X"D2",X"06",X"6E",X"B5",X"60",X"61",X"01",X"D5",
		X"45",X"10",X"85",X"B3",X"60",X"50",X"6A",X"5F",X"08",X"34",X"6A",X"00",X"4B",X"FE",X"E3",X"28",
		X"45",X"FE",X"E2",X"68",X"6A",X"04",X"34",X"0D",X"D6",X"34",X"4A",X"E5",X"04",X"6A",X"E2",X"34",
		X"D6",X"E5",X"0F",X"09",X"02",X"34",X"4A",X"C6",X"34",X"8A",X"8E",X"4A",X"B3",X"34",X"6A",X"8E",
		X"34",X"B5",X"8F",X"00",X"4A",X"43",X"34",X"B5",X"0C",X"21",X"93",X"90",X"00",X"4A",X"F1",X"50",
		X"09",X"5E",X"34",X"03",X"C5",X"08",X"B3",X"93",X"A8",X"93",X"B3",X"21",X"21",X"7F",X"CE",X"AF",
		X"09",X"A9",X"34",X"01",X"A8",X"34",X"41",X"05",X"00",X"4A",X"BD",X"34",X"5F",X"C9",X"C8",X"4A",
		X"CA",X"09",X"6E",X"13",X"34",X"9C",X"10",X"41",X"9D",X"00",X"01",X"BD",X"13",X"5F",X"05",X"C8",
		X"09",X"DF",X"13",X"01",X"DE",X"13",X"41",X"05",X"00",X"AF",X"BD",X"9C",X"5F",X"4A",X"C8",X"13",
		X"4A",X"4A",X"13",X"34",X"DE",X"FF",X"AF",X"4A",X"01",X"35",X"4A",X"00",X"35",X"4A",X"03",X"35",
		X"4A",X"04",X"35",X"B5",X"02",X"35",X"4A",X"BD",X"4A",X"09",X"FA",X"34",X"B5",X"C7",X"4A",X"B3",
		X"B6",X"B3",X"C6",X"28",X"09",X"1E",X"34",X"02",X"60",X"4A",X"6E",X"50",X"62",X"03",X"00",X"B5",
		X"14",X"11",X"41",X"BB",X"45",X"09",X"50",X"60",X"6E",X"B5",X"06",X"45",X"01",X"D5",X"25",X"6E",
		X"03",X"09",X"37",X"34",X"B5",X"C6",X"45",X"B3",X"BE",X"6D",X"8E",X"8E",X"6A",X"4A",X"34",X"34",
		X"6E",X"10",X"09",X"47",X"10",X"41",X"46",X"10",X"01",X"BD",X"00",X"B5",X"20",X"C8",X"5F",X"43",
		X"00",X"4A",X"FF",X"35",X"6A",X"03",X"34",X"6A",X"00",X"35",X"4A",X"69",X"35",X"B5",X"04",X"4B",
		X"93",X"C6",X"23",X"B3",X"E3",X"34",X"09",X"1E",X"08",X"28",X"B3",X"6A",X"B2",X"AC",X"3E",X"C6",
		X"34",X"13",X"7F",X"14",X"B3",X"B5",X"08",X"45",X"41",X"F8",X"11",X"6E",X"50",X"60",X"09",X"01",
		X"06",X"45",X"B5",X"03",X"25",X"6E",X"D5",X"B5",X"37",X"34",X"09",X"AE",X"45",X"B3",X"C6",X"6A",
		X"8F",X"8F",X"6D",X"6E",X"34",X"34",X"4A",X"10",X"09",X"03",X"10",X"01",X"02",X"10",X"41",X"20",
		X"00",X"B5",X"BD",X"00",X"5F",X"0C",X"C8",X"6A",X"01",X"35",X"4A",X"02",X"35",X"6A",X"03",X"35",
		X"4A",X"6B",X"35",X"60",X"04",X"4B",X"B5",X"4B",X"6E",X"50",X"4A",X"CE",X"01",X"60",X"03",X"B5",
		X"14",X"34",X"09",X"1E",X"45",X"B3",X"C6",X"92",X"B9",X"11",X"41",X"05",X"22",X"09",X"40",X"61",
		X"6E",X"B5",X"06",X"45",X"01",X"D5",X"41",X"09",X"08",X"6E",X"B3",X"B5",X"35",X"01",X"96",X"37",
		X"45",X"B3",X"C6",X"28",X"09",X"3E",X"34",X"8F",X"93",X"FA",X"22",X"09",X"B9",X"26",X"B5",X"C7",
		X"34",X"43",X"36",X"A6",X"B3",X"B3",X"28",X"09",X"92",X"4A",X"B3",X"50",X"35",X"90",X"96",X"6A",
		X"92",X"08",X"FE",X"60",X"35",X"DE",X"00",X"05",X"6E",X"45",X"B5",X"8F",X"02",X"09",X"37",X"35",
		X"B3",X"35",X"09",X"96",X"96",X"B3",X"59",X"B5",X"EC",X"AE",X"BD",X"7B",X"63",X"34",X"73",X"CA",
		X"28",X"00",X"09",X"AE",X"21",X"0A",X"00",X"34",X"B5",X"90",X"27",X"B5",X"1E",X"50",X"4A",X"45",
		X"46",X"B3",X"C6",X"28",X"09",X"36",X"34",X"F7",X"B3",X"46",X"B5",X"C6",X"A6",X"09",X"22",X"34",
		X"B3",X"B5",X"08",X"4B",X"56",X"6F",X"27",X"B5",X"22",X"34",X"09",X"76",X"46",X"B3",X"C6",X"08",
		X"21",X"C6",X"1F",X"6E",X"60",X"B5",X"B3",X"4B",X"60",X"09",X"B3",X"34",X"BA",X"C7",X"E6",X"B3",
		X"B6",X"B3",X"C6",X"08",X"09",X"3E",X"34",X"29",X"6A",X"FE",X"35",X"08",X"01",X"24",X"6C",X"02",
		X"6E",X"35",X"4A",X"03",X"23",X"4A",X"01",X"35",X"6A",X"FE",X"35",X"08",X"02",X"61",X"6C",X"02",
		X"6E",X"35",X"4A",X"04",X"60",X"4A",X"02",X"35",X"B5",X"6D",X"4B",X"93",X"10",X"4B",X"B5",X"E3",
		X"23",X"6C",X"FF",X"24",X"6A",X"FE",X"34",X"08",X"02",X"FF",X"23",X"4A",X"6E",X"34",X"4A",X"03",
		X"35",X"6C",X"00",X"61",X"6A",X"FE",X"35",X"08",X"02",X"00",X"60",X"4A",X"6E",X"35",X"4A",X"04",
		X"35",X"B5",X"10",X"4B",X"B5",X"6C",X"4B",X"93",X"E3",X"34",X"6A",X"00",X"23",X"FE",X"C8",X"08",
		X"2E",X"B3",X"C6",X"08",X"09",X"3E",X"34",X"2F",X"6A",X"00",X"34",X"36",X"8F",X"08",X"FE",X"B5",
		X"14",X"11",X"41",X"46",X"45",X"09",X"C0",X"61",X"6E",X"B5",X"06",X"45",X"01",X"D5",X"21",X"6E",
		X"02",X"B5",X"37",X"41",X"B5",X"BE",X"45",X"09",X"C5",X"93",X"B3",X"07",X"34",X"79",X"DE",X"D6",
		X"01",X"93",X"C8",X"23",X"4A",X"3F",X"34",X"6A",X"8E",X"08",X"FE",X"09",X"34",X"0D",X"00",X"C6",
		X"34",X"B2",X"1E",X"14",X"B3",X"B5",X"08",X"45",X"41",X"67",X"10",X"6E",X"D8",X"61",X"09",X"01",
		X"06",X"45",X"B5",X"03",X"44",X"6E",X"D5",X"B5",X"37",X"23",X"93",X"6A",X"45",X"B5",X"66",X"4B",
		X"93",X"68",X"23",X"93",X"43",X"4B",X"B5",X"43",X"23",X"BB",X"C1",X"09",X"2A",X"F5",X"34",X"00",
		X"00",X"7E",X"61",X"F5",X"F5",X"01",X"F5",X"86",X"02",X"F5",X"9E",X"02",X"17",X"5F",X"27",X"B3",
		X"68",X"68",X"68",X"68",X"B3",X"B3",X"B3",X"F5",X"7E",X"25",X"09",X"0F",X"00",X"B3",X"07",X"B5",
		X"C8",X"56",X"76",X"B9",X"45",X"BB",X"0B",X"43",X"25",X"25",X"25",X"25",X"43",X"64",X"44",X"0C",
		X"25",X"F5",X"25",X"04",X"2C",X"7E",X"B1",X"C0",X"F5",X"F5",X"04",X"04",X"5F",X"7E",X"B1",X"80",
		X"F5",X"F5",X"04",X"03",X"5F",X"7E",X"B1",X"80",X"F5",X"F5",X"03",X"03",X"5F",X"7E",X"B1",X"C0",
		X"F5",X"2A",X"03",X"34",X"5F",X"76",X"B1",X"BB",X"F5",X"F5",X"00",X"BB",X"09",X"61",X"00",X"01",
		X"00",X"BD",X"4F",X"9D",X"34",X"12",X"6F",X"F5",X"7E",X"25",X"09",X"0F",X"00",X"B3",X"57",X"B5",
		X"C8",X"56",X"76",X"B9",X"45",X"BB",X"0B",X"0F",X"26",X"25",X"25",X"26",X"1B",X"4E",X"8E",X"10",
		X"26",X"7E",X"26",X"4A",X"53",X"03",X"F5",X"74",X"34",X"4A",X"7E",X"34",X"F5",X"75",X"04",X"B5",
		X"ED",X"06",X"F5",X"6A",X"26",X"42",X"7E",X"22",X"34",X"47",X"00",X"23",X"FE",X"6A",X"08",X"34",
		X"FE",X"91",X"08",X"24",X"00",X"09",X"47",X"34",X"21",X"01",X"D1",X"00",X"9D",X"05",X"43",X"4E",
		X"FF",X"F5",X"C8",X"06",X"BD",X"7E",X"B1",X"43",X"42",X"7E",X"B9",X"09",X"60",X"06",X"F5",X"08",
		X"00",X"60",X"BB",X"B5",X"61",X"F6",X"42",X"9D",X"26",X"C0",X"7E",X"74",X"F5",X"4A",X"03",X"34",
		X"F5",X"75",X"04",X"B5",X"7E",X"34",X"4A",X"ED",X"26",X"FE",X"22",X"28",X"6A",X"00",X"34",X"4A",
		X"6A",X"0F",X"34",X"16",X"22",X"F5",X"B3",X"05",X"80",X"09",X"91",X"34",X"6D",X"24",X"FD",X"FD",
		X"21",X"FD",X"5B",X"01",X"FD",X"5A",X"00",X"FD",X"5F",X"FD",X"6C",X"03",X"02",X"5B",X"43",X"FD",
		X"5A",X"05",X"FD",X"74",X"04",X"6A",X"5F",X"34",X"F5",X"75",X"03",X"F5",X"5F",X"34",X"6A",X"5F",
		X"04",X"34",X"6A",X"00",X"B1",X"FE",X"23",X"B2",X"74",X"34",X"6A",X"0F",X"26",X"B3",X"23",X"96",
		X"27",X"80",X"16",X"FD",X"F5",X"91",X"05",X"09",X"24",X"FD",X"FD",X"00",X"34",X"5B",X"21",X"FD",
		X"5A",X"02",X"FD",X"09",X"01",X"6C",X"5F",X"08",X"00",X"5B",X"BB",X"FD",X"61",X"03",X"FD",X"5A",
		X"04",X"93",X"5F",X"25",X"FD",X"9D",X"05",X"F5",X"7E",X"34",X"4A",X"7E",X"03",X"F5",X"74",X"04",
		X"4A",X"CE",X"34",X"B5",X"75",X"25",X"93",X"9D",X"26",X"80",X"7E",X"AD",X"F5",X"93",X"03",X"25",
		X"B5",X"7E",X"26",X"C0",X"9D",X"04",X"F5",X"4A",X"75",X"03",X"F5",X"74",X"34",X"4A",X"7E",X"34",
		X"93",X"9D",X"25",X"F5",X"CE",X"26",X"B5",X"7E",X"04",X"F5",X"60",X"05",X"80",X"7E",X"BB",X"91",
		X"FD",X"FD",X"24",X"FD",X"09",X"21",X"34",X"5B",X"00",X"FD",X"5A",X"02",X"FD",X"5F",X"01",X"6A",
		X"74",X"03",X"F5",X"75",X"34",X"6A",X"5F",X"34",X"F5",X"7E",X"04",X"09",X"5F",X"00",X"F5",X"C0",
		X"26",X"C8",X"0F",X"D5",X"B3",X"45",X"B5",X"76",X"0B",X"F5",X"BB",X"06",X"56",X"7E",X"D1",X"B9",
		X"E4",X"E5",X"E4",X"A8",X"26",X"26",X"26",X"26",X"AB",X"B1",X"CA",X"FD",X"26",X"43",X"26",X"5B",
		X"03",X"FD",X"5A",X"05",X"FD",X"5F",X"04",X"B1",X"63",X"08",X"DB",X"61",X"60",X"00",X"09",X"BB",
		X"60",X"08",X"BB",X"4F",X"BC",X"00",X"41",X"6F",X"BD",X"99",X"BB",X"74",X"52",X"6A",X"60",X"34",
		X"9E",X"34",X"4A",X"75",X"07",X"6A",X"22",X"34",X"9E",X"34",X"4A",X"74",X"07",X"6A",X"23",X"34",
		X"B3",X"B3",X"B3",X"57",X"6F",X"6F",X"6F",X"6A",X"75",X"B3",X"B3",X"B3",X"34",X"6F",X"6F",X"6F",
		X"77",X"B1",X"F7",X"7E",X"B5",X"F5",X"44",X"01",X"F5",X"9E",X"02",X"F5",X"86",X"27",X"17",X"5F",
		X"02",X"68",X"68",X"68",X"B3",X"B3",X"B3",X"B3",X"68",X"35",X"6A",X"20",X"B1",X"09",X"03",X"27",
		X"B3",X"B5",X"B3",X"45",X"0F",X"C8",X"0F",X"B9",X"B5",X"B5",X"0F",X"0F",X"42",X"34",X"B1",X"B1",
		X"B5",X"B5",X"0F",X"0F",X"86",X"90",X"B1",X"B1",X"B5",X"B5",X"0F",X"28",X"FA",X"4C",X"B1",X"B1",
		X"B5",X"B5",X"28",X"28",X"3E",X"A8",X"B1",X"B1",X"B5",X"B5",X"28",X"29",X"9A",X"64",X"B1",X"B1",
		X"B5",X"B5",X"29",X"29",X"56",X"C0",X"B1",X"B1",X"B5",X"B5",X"29",X"29",X"B2",X"B3",X"B1",X"B1",
		X"B5",X"B5",X"29",X"29",X"B4",X"B5",X"B1",X"B1",X"D5",X"26",X"6F",X"46",X"4F",X"01",X"09",X"00",
		X"BD",X"6F",X"7D",X"40",X"52",X"09",X"4F",X"01",X"D1",X"BD",X"46",X"55",X"72",X"52",X"00",X"77",
		X"B1",X"3F",X"BE",X"09",X"7D",X"B1",X"03",X"C6",X"34",X"B3",X"16",X"28",X"B3",X"3E",X"B0",X"13",
		X"09",X"86",X"34",X"5F",X"A8",X"0F",X"7B",X"0B",X"7A",X"0B",X"0F",X"00",X"A6",X"6E",X"5F",X"A6",
		X"0F",X"60",X"68",X"09",X"5F",X"4A",X"02",X"C6",X"34",X"43",X"3E",X"DE",X"B3",X"09",X"28",X"13",
		X"41",X"05",X"13",X"4E",X"DF",X"00",X"01",X"10",X"BD",X"DE",X"AF",X"60",X"C8",X"13",X"4A",X"60",
		X"09",X"9D",X"13",X"01",X"9C",X"13",X"41",X"05",X"00",X"C8",X"10",X"4A",X"4E",X"AF",X"BD",X"9C",
		X"13",X"AB",X"05",X"60",X"60",X"34",X"09",X"EB",X"09",X"3E",X"34",X"74",X"C6",X"28",X"B3",X"09",
		X"AA",X"13",X"41",X"C9",X"34",X"6A",X"FB",X"34",X"DD",X"0B",X"0E",X"0B",X"B5",X"0B",X"40",X"BB",
		X"2A",X"FE",X"34",X"D0",X"8B",X"04",X"D9",X"B3",X"0F",X"6C",X"0F",X"C8",X"B3",X"B5",X"6C",X"45",
		X"B5",X"6A",X"41",X"34",X"AA",X"C8",X"D0",X"6C",X"4A",X"08",X"34",X"B3",X"C8",X"35",X"09",X"96",
		X"09",X"3E",X"34",X"42",X"C6",X"28",X"B3",X"6A",X"C9",X"C9",X"6C",X"6A",X"34",X"34",X"4A",X"8E");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
