library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity terrain_2c is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of terrain_2c is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"50",X"50",X"00",X"00",X"00",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"08",X"08",X"08",X"08",X"04",X"04",X"04",X"04",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"00",X"04",X"00",X"04",X"04",X"04",X"04",X"04",
		X"00",X"10",X"10",X"10",X"90",X"00",X"90",X"00",X"10",X"04",X"10",X"04",X"10",X"50",X"10",X"90",
		X"50",X"44",X"00",X"04",X"84",X"C4",X"04",X"44",X"00",X"10",X"00",X"10",X"00",X"10",X"00",X"10",
		X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"00",X"10",X"00",X"10",
		X"00",X"10",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"5C",X"D0",X"00",X"C0",X"5C",X"10",X"90",X"9C",X"9C",X"80",X"C0",
		X"00",X"50",X"40",X"10",X"10",X"5C",X"5C",X"40",X"1C",X"C0",X"5C",X"40",X"5C",X"50",X"00",X"C0",
		X"DC",X"10",X"DC",X"10",X"9C",X"50",X"40",X"00",X"80",X"80",X"1C",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"9C",X"10",X"9C",X"10",X"00",X"50",X"00",X"00",X"02",X"30",X"30",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"02",X"00",
		X"00",X"00",X"00",X"00",X"02",X"06",X"02",X"06",X"00",X"80",X"00",X"80",X"00",X"00",X"00",X"00",
		X"02",X"00",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"00",X"00",X"00",X"00",X"02",X"00",
		X"02",X"02",X"C2",X"02",X"02",X"02",X"02",X"00",X"02",X"02",X"02",X"02",X"02",X"02",X"00",X"00",
		X"00",X"00",X"02",X"00",X"02",X"02",X"00",X"00",X"02",X"00",X"C2",X"02",X"02",X"00",X"C2",X"02",
		X"02",X"02",X"00",X"82",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"02",X"02",X"02",X"02",
		X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"02",X"02",X"04",X"04",X"02",X"04",X"02",X"04",
		X"04",X"04",X"04",X"04",X"06",X"04",X"06",X"04",X"04",X"06",X"04",X"06",X"04",X"04",X"04",X"04",
		X"04",X"04",X"0A",X"0A",X"04",X"06",X"04",X"06",X"04",X"06",X"06",X"04",X"04",X"04",X"06",X"06",
		X"06",X"06",X"04",X"04",X"02",X"02",X"02",X"02",X"00",X"02",X"02",X"02",X"00",X"00",X"08",X"08",
		X"08",X"08",X"04",X"04",X"00",X"08",X"08",X"04",X"8C",X"8C",X"04",X"04",X"10",X"10",X"8C",X"8C",
		X"10",X"10",X"0C",X"8C",X"8C",X"0C",X"04",X"04",X"10",X"10",X"D0",X"D0",X"D0",X"D0",X"00",X"00",
		X"90",X"0C",X"08",X"90",X"00",X"00",X"90",X"00",X"00",X"00",X"10",X"10",X"90",X"00",X"10",X"10",
		X"10",X"10",X"50",X"10",X"10",X"10",X"50",X"10",X"D0",X"D0",X"90",X"00",X"10",X"10",X"D0",X"D0",
		X"90",X"00",X"50",X"90",X"10",X"90",X"50",X"90",X"10",X"10",X"10",X"D0",X"50",X"90",X"50",X"90",
		X"08",X"08",X"D0",X"D0",X"12",X"12",X"50",X"50",X"D0",X"D0",X"50",X"50",X"C6",X"C6",X"90",X"90",
		X"00",X"00",X"1C",X"1C",X"1C",X"9C",X"50",X"50",X"1C",X"1C",X"50",X"50",X"1C",X"9C",X"10",X"10",
		X"9C",X"9C",X"10",X"10",X"00",X"00",X"1C",X"00",X"1C",X"1C",X"DC",X"DC",X"10",X"5C",X"1C",X"00",
		X"00",X"9C",X"9C",X"5C",X"DC",X"1C",X"DC",X"1C",X"9C",X"10",X"9C",X"5C",X"9C",X"10",X"10",X"5C",
		X"5C",X"10",X"1C",X"10",X"1C",X"00",X"10",X"1C",X"50",X"1C",X"00",X"1C",X"10",X"1C",X"50",X"1C",
		X"00",X"C0",X"5C",X"C0",X"5C",X"40",X"1C",X"40",X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"20",
		X"40",X"20",X"00",X"20",X"00",X"00",X"40",X"20",X"20",X"20",X"40",X"40",X"00",X"00",X"20",X"20",
		X"20",X"20",X"00",X"40",X"00",X"00",X"20",X"20",X"20",X"40",X"40",X"40",X"20",X"C0",X"20",X"00",
		X"20",X"00",X"20",X"80",X"40",X"C0",X"20",X"A0",X"00",X"82",X"00",X"82",X"02",X"82",X"02",X"82",
		X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",
		X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",
		X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",
		X"06",X"06",X"06",X"06",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"00",X"0A",X"00",X"0A",
		X"01",X"01",X"01",X"01",X"A8",X"01",X"A8",X"01",X"28",X"A8",X"00",X"A8",X"A8",X"01",X"A8",X"01",
		X"00",X"E8",X"E8",X"01",X"00",X"00",X"68",X"68",X"68",X"68",X"01",X"01",X"68",X"68",X"01",X"01",
		X"00",X"00",X"E8",X"E8",X"00",X"00",X"E8",X"E8",X"E8",X"E8",X"01",X"01",X"E8",X"E8",X"01",X"01",
		X"00",X"00",X"1C",X"1C",X"00",X"00",X"1C",X"1C",X"00",X"00",X"1C",X"1C",X"00",X"00",X"1C",X"1C",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"C1",X"01",X"01",X"01",X"C1",X"01",X"01",X"01",X"C1",
		X"C1",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"C1",X"01",X"01",X"01",X"C1",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"41",X"01",X"01",X"01",X"01",X"01",X"01",X"C1",X"01",X"01",
		X"01",X"01",X"01",X"01",X"C1",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"41",X"01",X"01",X"01",X"41",X"01",
		X"41",X"41",X"01",X"01",X"01",X"81",X"01",X"81",X"01",X"01",X"01",X"81",X"41",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"C1",X"01",X"01",X"01",X"C1",X"01",X"01",X"C1",X"01",X"01",X"01",X"C1",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"C1",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"81",X"01",X"81",X"81",X"81",X"01",X"01",X"81",X"81",X"01",X"01",X"01",X"01",
		X"81",X"01",X"81",X"81",X"81",X"81",X"81",X"81",X"41",X"81",X"01",X"41",X"81",X"01",X"81",X"01",
		X"00",X"80",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"00",X"00",X"40",X"00",X"00",
		X"00",X"C0",X"00",X"00",X"00",X"80",X"00",X"80",X"C0",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",
		X"00",X"80",X"00",X"00",X"00",X"40",X"00",X"40",X"00",X"40",X"40",X"00",X"00",X"40",X"40",X"00",
		X"00",X"00",X"00",X"40",X"00",X"1C",X"10",X"5C",X"1C",X"50",X"00",X"1C",X"D0",X"D0",X"1C",X"1C",
		X"00",X"44",X"00",X"04",X"04",X"04",X"04",X"04",X"00",X"04",X"00",X"04",X"04",X"04",X"04",X"04",
		X"04",X"C4",X"04",X"C4",X"44",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"00",X"04",X"00",X"04",
		X"00",X"04",X"00",X"04",X"04",X"04",X"00",X"04",X"04",X"04",X"04",X"04",X"00",X"04",X"00",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"14",X"54",X"04",X"04",X"14",X"54",X"04",X"04",X"00",X"94",X"54",X"04",X"14",X"14",X"04",X"04",
		X"04",X"14",X"04",X"14",X"14",X"00",X"94",X"00",X"14",X"00",X"14",X"00",X"D4",X"00",X"94",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"20",X"20",X"C0",X"20",X"20",X"00",X"40",X"20",X"20",X"00",X"40",X"04",X"04",X"20",X"20",
		X"04",X"04",X"20",X"20",X"20",X"20",X"40",X"00",X"04",X"04",X"20",X"20",X"04",X"04",X"20",X"A0",
		X"20",X"A0",X"00",X"40",X"04",X"04",X"04",X"20",X"C4",X"20",X"20",X"C0",X"04",X"60",X"04",X"20",
		X"20",X"00",X"60",X"00",X"20",X"40",X"00",X"C0",X"A0",X"04",X"E0",X"04",X"00",X"00",X"00",X"00",
		X"00",X"00",X"1C",X"9C",X"50",X"50",X"00",X"9C",X"D0",X"00",X"9C",X"00",X"9C",X"10",X"10",X"10",
		X"00",X"DC",X"1C",X"9C",X"10",X"5C",X"90",X"00",X"9C",X"1C",X"00",X"9C",X"5C",X"1C",X"5C",X"1C",
		X"00",X"2C",X"02",X"02",X"00",X"00",X"AC",X"2C",X"0E",X"0E",X"04",X"04",X"02",X"02",X"04",X"44",
		X"02",X"02",X"0E",X"0E",X"00",X"00",X"18",X"18",X"50",X"10",X"9C",X"DC",X"5C",X"00",X"9C",X"9C",
		X"04",X"16",X"16",X"00",X"44",X"44",X"96",X"16",X"44",X"44",X"16",X"00",X"16",X"16",X"16",X"16",
		X"16",X"96",X"16",X"16",X"00",X"84",X"16",X"04",X"16",X"16",X"16",X"16",X"26",X"26",X"1A",X"1A",
		X"16",X"16",X"00",X"00",X"1A",X"1A",X"1A",X"1A",X"00",X"00",X"1A",X"16",X"1A",X"1A",X"1A",X"1A",
		X"9A",X"1A",X"1A",X"16",X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",
		X"00",X"16",X"D6",X"84",X"16",X"00",X"1A",X"1A",X"1A",X"16",X"16",X"16",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"05",X"01",X"01",X"01",X"05",X"05",X"05",X"01",
		X"05",X"01",X"01",X"01",X"05",X"05",X"01",X"05",X"01",X"01",X"01",X"01",X"05",X"05",X"01",X"05",
		X"01",X"01",X"09",X"01",X"01",X"01",X"01",X"01",X"41",X"01",X"45",X"01",X"09",X"01",X"09",X"01",
		X"41",X"41",X"41",X"45",X"01",X"01",X"01",X"01",X"4D",X"01",X"4D",X"01",X"0D",X"0D",X"11",X"01",
		X"01",X"01",X"0D",X"01",X"89",X"11",X"89",X"11",X"01",X"0D",X"11",X"0D",X"01",X"01",X"01",X"4D",
		X"41",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"11",X"01",X"01",X"01",X"15",X"15",X"0D",X"C1",
		X"09",X"01",X"09",X"41",X"09",X"01",X"09",X"01",X"01",X"01",X"01",X"41",X"01",X"01",X"09",X"09",
		X"C5",X"C5",X"11",X"11",X"01",X"01",X"01",X"01",X"01",X"09",X"01",X"09",X"09",X"01",X"09",X"09",
		X"01",X"41",X"09",X"41",X"01",X"01",X"01",X"01",X"81",X"05",X"41",X"81",X"01",X"05",X"01",X"09",
		X"01",X"01",X"01",X"01",X"81",X"05",X"01",X"01",X"01",X"CD",X"C5",X"01",X"01",X"01",X"C5",X"15",
		X"01",X"01",X"15",X"01",X"41",X"01",X"01",X"01",X"01",X"01",X"81",X"01",X"01",X"81",X"01",X"C1",
		X"01",X"01",X"01",X"41",X"01",X"41",X"01",X"01",X"01",X"01",X"05",X"01",X"01",X"01",X"C1",X"01",
		X"05",X"01",X"01",X"05",X"81",X"01",X"01",X"C1",X"01",X"01",X"01",X"41",X"41",X"01",X"41",X"01",
		X"01",X"01",X"0D",X"01",X"01",X"01",X"11",X"01",X"01",X"15",X"01",X"91",X"01",X"41",X"41",X"01",
		X"01",X"01",X"11",X"01",X"C1",X"01",X"01",X"81",X"01",X"01",X"41",X"41",X"01",X"01",X"01",X"01",
		X"01",X"41",X"01",X"01",X"41",X"41",X"11",X"41",X"41",X"41",X"8D",X"11",X"41",X"51",X"11",X"C5",
		X"81",X"05",X"01",X"81",X"01",X"01",X"01",X"41",X"15",X"C1",X"09",X"01",X"01",X"41",X"01",X"01",
		X"41",X"01",X"41",X"01",X"41",X"01",X"01",X"01",X"01",X"01",X"01",X"41",X"09",X"01",X"09",X"01",
		X"01",X"01",X"01",X"01",X"05",X"05",X"01",X"01",X"41",X"01",X"41",X"01",X"01",X"01",X"01",X"01",
		X"01",X"CD",X"01",X"01",X"01",X"01",X"01",X"CD",X"01",X"01",X"01",X"01",X"01",X"CD",X"01",X"01",
		X"05",X"05",X"01",X"01",X"01",X"01",X"4D",X"81",X"0D",X"4D",X"01",X"01",X"01",X"01",X"4D",X"01",
		X"01",X"01",X"05",X"0D",X"4D",X"01",X"0D",X"11",X"01",X"09",X"01",X"01",X"01",X"01",X"CD",X"CD",
		X"01",X"01",X"01",X"0D",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"41",X"01",X"01",X"01",X"01",X"01",X"09",X"01",X"01",X"09",X"01",X"01",X"01",X"01",
		X"01",X"01",X"09",X"01",X"01",X"01",X"01",X"01",X"09",X"01",X"09",X"01",X"01",X"01",X"01",X"41",
		X"15",X"41",X"09",X"01",X"01",X"01",X"01",X"01",X"01",X"41",X"09",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"09",X"01",X"01",X"01",X"41",X"01",X"01",X"09",X"01",X"09",X"01",X"01",X"01",X"41",
		X"01",X"09",X"01",X"09",X"09",X"01",X"09",X"01",X"C1",X"C1",X"01",X"09",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"09",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"09",X"01",
		X"09",X"01",X"09",X"41",X"CD",X"CD",X"01",X"01",X"01",X"01",X"19",X"19",X"CD",X"01",X"19",X"01",
		X"01",X"01",X"01",X"09",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"81",X"01",X"01",X"81",
		X"01",X"01",X"01",X"01",X"05",X"05",X"01",X"81",X"01",X"01",X"09",X"41",X"09",X"09",X"01",X"09",
		X"09",X"01",X"09",X"01",X"09",X"09",X"01",X"09",X"C1",X"01",X"41",X"01",X"41",X"01",X"41",X"41",
		X"41",X"01",X"81",X"01",X"01",X"01",X"09",X"01",X"01",X"01",X"41",X"01",X"41",X"01",X"41",X"01",
		X"00",X"01",X"02",X"03",X"2A",X"2A",X"24",X"24",X"2A",X"2A",X"02",X"03",X"00",X"28",X"28",X"24",
		X"24",X"24",X"24",X"24",X"10",X"11",X"12",X"13",X"10",X"11",X"12",X"13",X"81",X"83",X"80",X"82",
		X"85",X"87",X"84",X"86",X"25",X"24",X"25",X"24",X"00",X"3B",X"02",X"3B",X"44",X"44",X"44",X"44",
		X"00",X"28",X"2A",X"24",X"25",X"01",X"25",X"03",X"2A",X"39",X"24",X"3A",X"24",X"2A",X"24",X"28",
		X"2A",X"39",X"02",X"3B",X"44",X"44",X"44",X"44",X"00",X"26",X"02",X"25",X"00",X"25",X"02",X"25",
		X"00",X"01",X"2A",X"2A",X"27",X"24",X"2F",X"24",X"27",X"24",X"26",X"24",X"00",X"27",X"02",X"26",
		X"00",X"25",X"28",X"24",X"89",X"8B",X"88",X"8A",X"8D",X"8F",X"8C",X"8E",X"91",X"93",X"90",X"92",
		X"95",X"97",X"94",X"96",X"99",X"9B",X"98",X"9A",X"9D",X"9F",X"9C",X"9E",X"A1",X"A3",X"A0",X"A2",
		X"A5",X"A7",X"A4",X"A6",X"24",X"4A",X"28",X"A9",X"03",X"50",X"28",X"32",X"52",X"49",X"A8",X"03",
		X"AD",X"26",X"AD",X"31",X"2A",X"4A",X"4A",X"A8",X"49",X"AD",X"48",X"AE",X"58",X"2A",X"AD",X"03",
		X"49",X"2A",X"53",X"24",X"53",X"2A",X"AD",X"02",X"A9",X"A8",X"58",X"2A",X"2A",X"24",X"24",X"24",
		X"25",X"24",X"24",X"24",X"4A",X"2A",X"49",X"24",X"00",X"27",X"02",X"03",X"C8",X"D0",X"D0",X"24",
		X"01",X"05",X"03",X"04",X"01",X"05",X"03",X"05",X"07",X"07",X"06",X"06",X"0A",X"07",X"0A",X"07",
		X"07",X"07",X"07",X"07",X"0C",X"0D",X"0C",X"0D",X"07",X"05",X"07",X"05",X"05",X"07",X"04",X"06",
		X"0E",X"07",X"0C",X"0E",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"06",X"06",X"07",X"07",X"0B",X"07",
		X"0A",X"0B",X"0B",X"0A",X"0A",X"0A",X"0A",X"07",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"07",X"07",
		X"07",X"07",X"0A",X"07",X"0A",X"0A",X"06",X"06",X"0A",X"07",X"0B",X"0B",X"0B",X"07",X"0B",X"0A",
		X"0A",X"0A",X"07",X"0B",X"C0",X"C1",X"C2",X"C3",X"C4",X"C5",X"C6",X"C7",X"C8",X"C8",X"C8",X"C8",
		X"C9",X"C2",X"C9",X"C0",X"C0",X"C4",X"CA",X"CA",X"C8",X"C8",X"C2",X"C5",X"C8",X"C9",X"C8",X"CB",
		X"C9",X"C0",X"CB",X"CA",X"CD",X"C0",X"CC",X"C5",X"C8",X"CD",X"C8",X"CC",X"C8",X"C8",X"C8",X"C8",
		X"C8",X"C8",X"CE",X"CE",X"C8",X"CF",X"C8",X"CF",X"C8",X"D0",X"D0",X"C0",X"C8",X"C8",X"D1",X"D2",
		X"D1",X"D2",X"C2",X"C4",X"D3",X"D4",X"C8",X"C8",X"90",X"D5",X"D5",X"C8",X"98",X"A0",X"D3",X"D4",
		X"D3",X"D4",X"C8",X"C8",X"93",X"D5",X"D5",X"C8",X"D2",X"D1",X"C0",X"C2",X"24",X"24",X"D2",X"D1",
		X"24",X"24",X"D6",X"D6",X"D6",X"D6",X"C2",X"C5",X"24",X"24",X"2C",X"2B",X"2C",X"2B",X"00",X"00",
		X"D0",X"C8",X"C8",X"D0",X"00",X"02",X"28",X"01",X"00",X"02",X"28",X"2A",X"25",X"02",X"24",X"2A",
		X"24",X"24",X"28",X"24",X"2B",X"2C",X"28",X"24",X"2C",X"2B",X"28",X"00",X"2B",X"2C",X"2C",X"2B",
		X"28",X"00",X"28",X"28",X"24",X"27",X"28",X"26",X"28",X"24",X"24",X"28",X"26",X"27",X"27",X"26",
		X"C8",X"C8",X"D2",X"D1",X"D6",X"D6",X"2A",X"2A",X"D2",X"D1",X"2B",X"2C",X"D2",X"D1",X"2C",X"2B",
		X"88",X"8A",X"45",X"46",X"47",X"47",X"24",X"24",X"45",X"46",X"2B",X"2C",X"47",X"47",X"24",X"24",
		X"46",X"45",X"24",X"24",X"89",X"8B",X"48",X"8A",X"45",X"46",X"46",X"45",X"24",X"48",X"47",X"8E",
		X"8D",X"48",X"48",X"48",X"49",X"4A",X"4A",X"49",X"4A",X"24",X"49",X"48",X"48",X"24",X"24",X"48",
		X"4B",X"24",X"4B",X"24",X"48",X"8B",X"24",X"48",X"28",X"51",X"00",X"50",X"24",X"53",X"2A",X"52",
		X"A9",X"9F",X"50",X"B3",X"49",X"A9",X"50",X"AE",X"91",X"DC",X"95",X"90",X"A1",X"DE",X"95",X"DD",
		X"95",X"E0",X"8F",X"DF",X"8E",X"90",X"93",X"E1",X"E2",X"E4",X"9A",X"9F",X"9F",X"A5",X"E3",X"E5",
		X"E6",X"E8",X"90",X"92",X"9A",X"9B",X"E7",X"E9",X"EA",X"95",X"A5",X"9B",X"EC",X"95",X"EB",X"93",
		X"EE",X"93",X"ED",X"8F",X"A0",X"A1",X"EF",X"9D",X"01",X"12",X"00",X"11",X"12",X"00",X"11",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"0D",X"00",X"10",X"00",X"0F",X"12",X"13",X"11",X"13",
		X"01",X"13",X"00",X"01",X"13",X"13",X"13",X"13",X"09",X"09",X"09",X"09",X"14",X"14",X"14",X"14",
		X"13",X"15",X"15",X"14",X"13",X"17",X"13",X"16",X"17",X"14",X"16",X"14",X"00",X"00",X"0A",X"00",
		X"0A",X"00",X"09",X"0A",X"00",X"12",X"00",X"11",X"12",X"13",X"11",X"13",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"19",X"00",X"18",X"00",X"01",X"19",X"00",X"18",X"1A",X"00",X"1A",X"00",
		X"03",X"10",X"10",X"00",X"00",X"01",X"15",X"16",X"15",X"16",X"00",X"00",X"17",X"17",X"00",X"00",
		X"03",X"01",X"14",X"13",X"03",X"00",X"12",X"11",X"14",X"13",X"00",X"00",X"12",X"11",X"00",X"00",
		X"91",X"92",X"B4",X"B5",X"93",X"94",X"B6",X"B7",X"9B",X"9A",X"B8",X"B9",X"99",X"9F",X"BA",X"BB",
		X"00",X"01",X"00",X"00",X"02",X"03",X"03",X"02",X"04",X"05",X"06",X"04",X"07",X"00",X"08",X"07",
		X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"09",X"0A",X"00",X"00",X"00",X"0B",X"00",X"0C",
		X"0D",X"0E",X"0B",X"00",X"00",X"0E",X"0A",X"0F",X"00",X"00",X"0E",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"10",X"0E",X"11",X"11",X"12",X"0E",X"00",X"13",X"14",X"0E",X"15",X"16",X"17",X"0E",X"18",
		X"14",X"14",X"15",X"15",X"16",X"17",X"16",X"17",X"19",X"1B",X"15",X"1A",X"1C",X"1D",X"16",X"1E",
		X"00",X"1F",X"00",X"00",X"22",X"15",X"20",X"21",X"00",X"23",X"00",X"00",X"24",X"16",X"25",X"26",
		X"15",X"15",X"27",X"21",X"24",X"16",X"28",X"16",X"29",X"21",X"00",X"2A",X"2B",X"24",X"00",X"2C",
		X"15",X"15",X"21",X"21",X"24",X"16",X"24",X"16",X"15",X"1A",X"21",X"21",X"24",X"1C",X"24",X"16",
		X"00",X"00",X"2D",X"00",X"00",X"00",X"2E",X"00",X"2D",X"00",X"19",X"1B",X"1D",X"00",X"1E",X"2E",
		X"21",X"21",X"14",X"14",X"17",X"24",X"17",X"24",X"14",X"14",X"2F",X"15",X"16",X"17",X"30",X"17",
		X"00",X"00",X"21",X"21",X"00",X"00",X"47",X"00",X"21",X"21",X"00",X"00",X"00",X"1D",X"00",X"00",
		X"07",X"00",X"08",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"2D",X"00",X"00",X"00",X"2E",X"00",
		X"00",X"31",X"32",X"15",X"16",X"33",X"34",X"00",X"00",X"35",X"0E",X"00",X"00",X"36",X"0E",X"00",
		X"14",X"14",X"15",X"15",X"16",X"17",X"16",X"17",X"37",X"38",X"00",X"16",X"15",X"39",X"00",X"3A",
		X"3B",X"3C",X"15",X"3D",X"3E",X"3F",X"16",X"40",X"41",X"00",X"42",X"43",X"44",X"00",X"45",X"46",
		X"47",X"00",X"47",X"00",X"00",X"00",X"48",X"48",X"00",X"00",X"47",X"00",X"00",X"00",X"48",X"00",
		X"49",X"4A",X"4B",X"4C",X"4D",X"4E",X"4F",X"50",X"51",X"52",X"53",X"54",X"55",X"56",X"57",X"58",
		X"59",X"5A",X"35",X"00",X"00",X"5B",X"36",X"5C",X"37",X"35",X"00",X"00",X"00",X"36",X"00",X"3A",
		X"5D",X"5E",X"5F",X"60",X"61",X"62",X"63",X"64",X"65",X"66",X"67",X"68",X"69",X"6A",X"6B",X"6C",
		X"6D",X"6E",X"6F",X"70",X"71",X"72",X"73",X"74",X"75",X"76",X"77",X"78",X"79",X"7A",X"7B",X"7C",
		X"7D",X"7E",X"7F",X"80",X"81",X"82",X"83",X"84",X"85",X"86",X"87",X"88",X"89",X"8A",X"8B",X"8C",
		X"8D",X"8E",X"8F",X"90",X"91",X"92",X"92",X"93",X"94",X"95",X"95",X"94",X"96",X"97",X"98",X"99",
		X"00",X"1B",X"9A",X"17",X"9A",X"17",X"17",X"17",X"00",X"9A",X"16",X"17",X"00",X"00",X"1B",X"00",
		X"24",X"1B",X"17",X"24",X"17",X"17",X"17",X"17",X"48",X"17",X"00",X"48",X"24",X"1B",X"17",X"9B",
		X"90",X"B2",X"94",X"A8",X"00",X"AA",X"00",X"AA",X"8C",X"A9",X"B3",X"00",X"00",X"A9",X"00",X"A8",
		X"00",X"AD",X"00",X"A9",X"00",X"AD",X"00",X"AD",X"AC",X"00",X"A0",X"B0",X"00",X"00",X"A8",X"00",
		X"00",X"AD",X"00",X"AC",X"00",X"A8",X"00",X"AE",X"92",X"B3",X"AD",X"00",X"00",X"B1",X"A8",X"89",
		X"00",X"00",X"B0",X"B1",X"00",X"54",X"2A",X"53",X"55",X"28",X"88",X"55",X"2C",X"2B",X"56",X"57",
		X"01",X"3B",X"00",X"3C",X"3D",X"44",X"3C",X"44",X"01",X"3D",X"00",X"3C",X"4D",X"44",X"4C",X"44",
		X"44",X"4E",X"44",X"4F",X"39",X"44",X"3B",X"44",X"39",X"44",X"3A",X"44",X"01",X"4D",X"00",X"4C",
		X"01",X"4F",X"00",X"4E",X"3F",X"43",X"01",X"3F",X"43",X"43",X"43",X"43",X"00",X"3E",X"02",X"3E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AC",X"B0",X"C0",X"C1",X"B1",X"B0",X"C0",X"C1",X"88",X"A8",X"B3",X"C1",X"B1",X"B1",X"C0",X"C1",
		X"C2",X"A9",X"C0",X"AA",X"AB",X"94",X"AD",X"90",X"AE",X"99",X"B2",X"98",X"B3",X"9B",X"AD",X"9A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C4",X"10",X"10",X"03",X"11",X"12",X"00",X"03",X"13",X"14",X"02",X"01",X"C0",X"C3",X"11",X"12",
		X"C0",X"C3",X"13",X"14",X"15",X"16",X"03",X"00",X"C3",X"C0",X"15",X"16",X"C1",X"C2",X"15",X"15",
		X"15",X"15",X"00",X"03",X"C1",X"C2",X"C0",X"10",X"C2",X"10",X"10",X"03",X"C1",X"1A",X"C0",X"1A",
		X"1A",X"01",X"1A",X"02",X"10",X"02",X"01",X"03",X"1A",X"C7",X"10",X"C0",X"00",X"00",X"00",X"00",
		X"88",X"8A",X"47",X"47",X"28",X"2A",X"02",X"57",X"28",X"03",X"56",X"8A",X"48",X"24",X"24",X"24",
		X"89",X"48",X"47",X"48",X"24",X"48",X"25",X"8A",X"56",X"58",X"88",X"49",X"49",X"55",X"4A",X"59",
		X"8C",X"82",X"C8",X"C8",X"8D",X"8C",X"80",X"B1",X"D8",X"D9",X"C5",X"C0",X"C8",X"C8",X"C2",X"C0",
		X"C8",X"C8",X"D8",X"D9",X"01",X"02",X"DA",X"DB",X"2A",X"24",X"55",X"48",X"59",X"8B",X"46",X"45",
		X"C0",X"1D",X"1E",X"00",X"C0",X"C2",X"1E",X"1F",X"C2",X"C0",X"20",X"01",X"22",X"21",X"09",X"09",
		X"23",X"1D",X"24",X"23",X"01",X"C2",X"20",X"C0",X"23",X"09",X"24",X"23",X"26",X"25",X"0B",X"0C",
		X"26",X"25",X"00",X"00",X"29",X"27",X"28",X"27",X"01",X"03",X"00",X"20",X"2A",X"2B",X"00",X"00",
		X"2A",X"2C",X"00",X"2D",X"27",X"27",X"2E",X"27",X"27",X"27",X"30",X"2F",X"00",X"31",X"0B",X"0C",
		X"00",X"32",X"1D",X"C0",X"33",X"01",X"0B",X"0C",X"00",X"33",X"2D",X"34",X"80",X"80",X"81",X"80",
		X"80",X"82",X"81",X"80",X"83",X"81",X"82",X"83",X"80",X"82",X"80",X"80",X"85",X"84",X"82",X"83",
		X"88",X"87",X"86",X"80",X"8A",X"89",X"80",X"80",X"80",X"8D",X"8B",X"8C",X"80",X"80",X"80",X"8B",
		X"80",X"8A",X"8E",X"80",X"80",X"80",X"8F",X"80",X"92",X"93",X"90",X"91",X"80",X"80",X"93",X"80",
		X"83",X"94",X"80",X"83",X"96",X"93",X"89",X"95",X"90",X"98",X"91",X"97",X"80",X"9A",X"80",X"99",
		X"89",X"90",X"8C",X"91",X"80",X"9C",X"80",X"9B",X"8A",X"80",X"8B",X"80",X"83",X"8F",X"80",X"9D",
		X"9E",X"80",X"94",X"9E",X"8B",X"80",X"8A",X"80",X"9F",X"94",X"80",X"83",X"A1",X"80",X"A0",X"8E",
		X"98",X"80",X"A1",X"80",X"80",X"80",X"A2",X"80",X"80",X"AA",X"A4",X"A9",X"80",X"80",X"83",X"9F",
		X"80",X"90",X"80",X"83",X"80",X"A1",X"80",X"A3",X"81",X"80",X"83",X"98",X"A4",X"A5",X"80",X"80",
		X"A5",X"A4",X"80",X"80",X"80",X"A7",X"A6",X"A8",X"82",X"80",X"80",X"80",X"80",X"90",X"80",X"80",
		X"90",X"98",X"80",X"99",X"A1",X"80",X"A3",X"80",X"8E",X"80",X"98",X"8E",X"80",X"AB",X"80",X"80",
		X"80",X"AD",X"80",X"AC",X"8E",X"80",X"80",X"AE",X"AF",X"88",X"A5",X"B0",X"B2",X"B1",X"A4",X"80",
		X"B3",X"80",X"80",X"B4",X"A1",X"80",X"A1",X"80",X"80",X"B5",X"81",X"98",X"80",X"98",X"80",X"98",
		X"80",X"B6",X"80",X"B6",X"B7",X"98",X"80",X"B8",X"81",X"80",X"94",X"81",X"80",X"80",X"B7",X"B9",
		X"94",X"81",X"BA",X"94",X"B5",X"80",X"B6",X"B6",X"80",X"A3",X"80",X"9B",X"97",X"89",X"98",X"80",
		X"A1",X"80",X"9D",X"80",X"9F",X"98",X"80",X"A1",X"BB",X"80",X"9F",X"BB",X"BC",X"98",X"9F",X"BD",
		X"9F",X"C1",X"80",X"C0",X"B7",X"B9",X"BE",X"BE",X"80",X"89",X"B9",X"B1",X"C3",X"C2",X"80",X"80",
		X"C4",X"BE",X"A5",X"BF",X"BE",X"BE",X"80",X"9F",X"BE",X"BE",X"83",X"80",X"BE",X"BB",X"80",X"A5",
		X"8E",X"80",X"C5",X"8E",X"AD",X"80",X"AC",X"97",X"B3",X"B6",X"80",X"A1",X"A3",X"BD",X"AC",X"A1",
		X"BD",X"80",X"99",X"80",X"AC",X"80",X"AC",X"80",X"81",X"80",X"83",X"BD",X"80",X"AD",X"80",X"AC",
		X"88",X"87",X"80",X"80",X"80",X"80",X"80",X"80",X"99",X"80",X"9A",X"80",X"80",X"80",X"C6",X"C7",
		X"C9",X"88",X"C8",X"CA",X"80",X"80",X"CC",X"88",X"80",X"80",X"CB",X"AF",X"AF",X"88",X"CD",X"B0",
		X"80",X"80",X"88",X"87",X"80",X"80",X"88",X"AF",X"94",X"8E",X"CD",X"A6",X"80",X"80",X"8E",X"80",
		X"AC",X"CE",X"AB",X"91",X"8E",X"89",X"94",X"8D",X"89",X"80",X"80",X"BA",X"80",X"80",X"87",X"88",
		X"D0",X"9E",X"CF",X"94",X"82",X"90",X"80",X"D1",X"D2",X"80",X"90",X"D0",X"D3",X"80",X"90",X"D2",
		X"A2",X"80",X"98",X"80",X"84",X"80",X"85",X"D2",X"80",X"D4",X"82",X"80",X"D5",X"D6",X"80",X"80",
		X"90",X"84",X"80",X"85",X"80",X"BA",X"D2",X"89",X"80",X"AD",X"80",X"85",X"81",X"80",X"83",X"BD",
		X"B1",X"BD",X"80",X"AD",X"80",X"80",X"D2",X"80",X"AC",X"BD",X"80",X"AD",X"D7",X"88",X"AD",X"80",
		X"D4",X"D2",X"80",X"AC",X"80",X"BA",X"98",X"89",X"D8",X"80",X"BA",X"80",X"AD",X"80",X"AC",X"BD",
		X"89",X"80",X"D9",X"80",X"80",X"AD",X"80",X"85",X"06",X"D5",X"82",X"80",X"80",X"82",X"DA",X"80",
		X"D4",X"DB",X"82",X"80",X"AD",X"80",X"90",X"D2",X"DA",X"80",X"AD",X"80",X"85",X"D2",X"80",X"AC",
		X"80",X"AD",X"80",X"AC",X"87",X"88",X"A6",X"CA",X"80",X"80",X"80",X"80",X"88",X"80",X"80",X"DC",
		X"BA",X"AC",X"89",X"80",X"88",X"87",X"D2",X"80",X"DD",X"D2",X"89",X"90",X"8E",X"80",X"D2",X"8E",
		X"DE",X"E0",X"98",X"DF",X"80",X"80",X"E1",X"8E",X"E2",X"E1",X"80",X"AC",X"80",X"80",X"E3",X"80",
		X"80",X"9A",X"80",X"99",X"80",X"80",X"82",X"80",X"B6",X"82",X"98",X"80",X"AC",X"98",X"AC",X"A2",
		X"AD",X"80",X"B6",X"80",X"E4",X"B9",X"80",X"A3",X"A2",X"80",X"98",X"80",X"99",X"80",X"9A",X"80");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
