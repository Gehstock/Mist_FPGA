library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity a32a is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(9 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of a32a is
	type rom is array(0 to  1023) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"38",X"44",X"64",X"54",X"4C",X"44",X"38",X"01",X"10",X"18",X"10",X"10",X"10",X"10",X"38",
		X"02",X"38",X"44",X"40",X"20",X"10",X"08",X"7C",X"03",X"7C",X"20",X"10",X"20",X"40",X"44",X"38",
		X"04",X"30",X"28",X"24",X"7C",X"20",X"20",X"20",X"05",X"7C",X"04",X"3C",X"40",X"40",X"44",X"38",
		X"06",X"30",X"08",X"04",X"3C",X"44",X"44",X"38",X"07",X"7C",X"40",X"20",X"10",X"08",X"08",X"08",
		X"08",X"38",X"44",X"44",X"38",X"44",X"44",X"38",X"09",X"38",X"44",X"44",X"78",X"40",X"20",X"18",
		X"0A",X"38",X"44",X"44",X"7C",X"44",X"44",X"44",X"0B",X"3C",X"44",X"44",X"3C",X"44",X"44",X"3C",
		X"0C",X"38",X"44",X"04",X"04",X"04",X"44",X"38",X"0D",X"1C",X"24",X"44",X"44",X"44",X"24",X"1C",
		X"0E",X"7C",X"04",X"04",X"3C",X"04",X"04",X"7C",X"0F",X"7C",X"04",X"04",X"1C",X"04",X"04",X"04",
		X"10",X"78",X"04",X"04",X"64",X"44",X"44",X"78",X"11",X"44",X"44",X"44",X"7C",X"44",X"44",X"44",
		X"12",X"38",X"10",X"10",X"10",X"10",X"10",X"38",X"13",X"70",X"20",X"20",X"20",X"20",X"24",X"18",
		X"14",X"44",X"24",X"14",X"0C",X"14",X"24",X"44",X"15",X"04",X"04",X"04",X"04",X"04",X"04",X"7C",
		X"16",X"44",X"6C",X"54",X"54",X"44",X"44",X"44",X"17",X"44",X"44",X"4C",X"54",X"64",X"44",X"44",
		X"18",X"38",X"44",X"44",X"44",X"44",X"44",X"38",X"19",X"3C",X"44",X"44",X"3C",X"04",X"04",X"04",
		X"1A",X"38",X"44",X"44",X"44",X"54",X"24",X"58",X"1B",X"3C",X"44",X"44",X"3C",X"14",X"24",X"44",
		X"1C",X"78",X"04",X"04",X"38",X"40",X"40",X"3C",X"1D",X"7C",X"10",X"10",X"10",X"10",X"10",X"10",
		X"1E",X"44",X"44",X"44",X"44",X"44",X"44",X"38",X"1F",X"44",X"44",X"44",X"44",X"44",X"28",X"10",
		X"05",X"3D",X"C2",X"F7",X"11",X"C9",X"21",X"08",X"2D",X"11",X"82",X"20",X"CD",X"34",X"12",X"21",
		X"08",X"2F",X"11",X"92",X"20",X"CD",X"34",X"12",X"21",X"08",X"31",X"11",X"A2",X"20",X"CD",X"34",
		X"12",X"21",X"08",X"33",X"11",X"B2",X"20",X"CD",X"34",X"12",X"21",X"08",X"35",X"11",X"C2",X"20",
		X"CD",X"34",X"12",X"C9",X"1A",X"D5",X"E5",X"CD",X"40",X"11",X"E1",X"23",X"D1",X"13",X"7B",X"E6",
		X"0F",X"FE",X"00",X"C8",X"C3",X"34",X"12",X"21",X"08",X"2D",X"AF",X"77",X"23",X"7D",X"E6",X"1F",
		X"FE",X"16",X"CA",X"58",X"12",X"C3",X"4A",X"12",X"11",X"12",X"00",X"19",X"7C",X"FE",X"36",X"C8",
		X"C3",X"4A",X"12",X"CD",X"8A",X"11",X"21",X"22",X"36",X"22",X"E0",X"20",X"3E",X"0A",X"32",X"E2",
		X"20",X"CD",X"D9",X"11",X"21",X"D5",X"20",X"22",X"E3",X"20",X"21",X"0D",X"2D",X"22",X"E5",X"20",
		X"21",X"FF",X"01",X"22",X"E7",X"20",X"DB",X"00",X"1F",X"D2",X"B3",X"12",X"1F",X"D2",X"D4",X"12",
		X"DB",X"00",X"1F",X"1F",X"1F",X"D2",X"F0",X"12",X"CD",X"EB",X"11",X"3A",X"01",X"21",X"B7",X"C0",
		X"3E",X"05",X"CD",X"F7",X"11",X"2A",X"E7",X"20",X"2B",X"22",X"E7",X"20",X"7C",X"FE",X"00",X"C8",
		X"C3",X"86",X"12",X"3A",X"E0",X"20",X"FE",X"3D",X"CA",X"90",X"12",X"2A",X"E0",X"20",X"CD",X"E6",
		X"11",X"23",X"22",X"E0",X"20",X"CD",X"D9",X"11",X"21",X"E2",X"20",X"34",X"3E",X"02",X"CD",X"F7",
		X"11",X"C3",X"90",X"12",X"3A",X"E0",X"20",X"FE",X"22",X"CA",X"90",X"12",X"2A",X"E0",X"20",X"CD",
		X"E6",X"11",X"2B",X"22",X"E0",X"20",X"CD",X"D9",X"11",X"21",X"E2",X"20",X"35",X"C3",X"CC",X"12",
		X"2A",X"E3",X"20",X"3A",X"E2",X"20",X"77",X"23",X"22",X"E3",X"20",X"2A",X"E5",X"20",X"CD",X"40",
		X"20",X"44",X"44",X"44",X"54",X"54",X"54",X"28",X"21",X"44",X"44",X"28",X"10",X"28",X"44",X"44",
		X"22",X"44",X"44",X"44",X"28",X"10",X"10",X"10",X"23",X"7C",X"40",X"20",X"10",X"08",X"04",X"7C",
		X"24",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"25",X"00",X"00",X"00",X"00",X"00",X"18",X"18",
		X"0E",X"07",X"1A",X"77",X"13",X"0D",X"C8",X"D5",X"11",X"20",X"00",X"19",X"D1",X"C3",X"32",X"11",
		X"E5",X"21",X"00",X"10",X"01",X"08",X"00",X"BE",X"CA",X"4F",X"11",X"09",X"C3",X"47",X"11",X"23",
		X"EB",X"E1",X"CD",X"30",X"11",X"C9",X"F5",X"C5",X"D5",X"E5",X"EB",X"01",X"F0",X"D8",X"CD",X"7A",
		X"11",X"01",X"18",X"FC",X"CD",X"7A",X"11",X"01",X"9C",X"FF",X"CD",X"7A",X"11",X"01",X"F6",X"FF",
		X"CD",X"7A",X"11",X"7D",X"12",X"E1",X"D1",X"C1",X"F1",X"C9",X"AF",X"D5",X"5D",X"54",X"3C",X"09",
		X"DA",X"7C",X"11",X"3D",X"6B",X"62",X"D1",X"12",X"13",X"C9",X"3E",X"0A",X"21",X"02",X"35",X"E5",
		X"F5",X"CD",X"40",X"11",X"F1",X"E1",X"23",X"3C",X"FE",X"26",X"C2",X"8F",X"11",X"C9",X"21",X"82",
		X"20",X"3E",X"01",X"CD",X"C7",X"11",X"21",X"92",X"20",X"3E",X"02",X"CD",X"C7",X"11",X"21",X"A2",
		X"20",X"3E",X"03",X"CD",X"C7",X"11",X"21",X"B2",X"20",X"3E",X"04",X"CD",X"C7",X"11",X"21",X"C2",
		X"20",X"3E",X"05",X"C3",X"F0",X"13",X"C9",X"77",X"23",X"3E",X"25",X"77",X"23",X"3E",X"24",X"77",
		X"7D",X"E6",X"0F",X"FE",X"0F",X"C8",X"C3",X"CC",X"11",X"E5",X"3E",X"7C",X"77",X"11",X"20",X"00",
		X"19",X"77",X"00",X"00",X"E1",X"C9",X"E5",X"AF",X"C3",X"DC",X"11",X"DB",X"00",X"17",X"D8",X"3E",
		X"01",X"32",X"01",X"21",X"C9",X"3E",X"FF",X"F5",X"CD",X"B2",X"19",X"CD",X"23",X"00",X"F1",X"D3",
		X"11",X"2A",X"E5",X"20",X"23",X"22",X"E5",X"20",X"3E",X"20",X"CD",X"F7",X"11",X"2A",X"E3",X"20",
		X"7D",X"FE",X"D8",X"C2",X"98",X"12",X"CD",X"FA",X"13",X"C9",X"7E",X"12",X"7D",X"E6",X"0F",X"FE",
		X"01",X"CA",X"2C",X"13",X"FE",X"0F",X"C8",X"23",X"13",X"C3",X"1A",X"13",X"23",X"13",X"23",X"13",
		X"23",X"13",X"C3",X"1A",X"13",X"EB",X"2A",X"D0",X"20",X"7D",X"93",X"7C",X"9A",X"C9",X"21",X"DB",
		X"20",X"7E",X"B7",X"CA",X"47",X"13",X"C9",X"3E",X"24",X"77",X"23",X"C3",X"41",X"13",X"21",X"B0",
		X"20",X"11",X"C0",X"20",X"CD",X"1A",X"13",X"2A",X"C0",X"20",X"CD",X"35",X"13",X"FA",X"A0",X"13",
		X"21",X"A0",X"20",X"11",X"B0",X"20",X"CD",X"1A",X"13",X"2A",X"B0",X"20",X"CD",X"35",X"13",X"FA",
		X"A6",X"13",X"21",X"90",X"20",X"11",X"A0",X"20",X"CD",X"1A",X"13",X"2A",X"A0",X"20",X"CD",X"35",
		X"13",X"FA",X"AC",X"13",X"21",X"80",X"20",X"11",X"90",X"20",X"CD",X"1A",X"13",X"2A",X"90",X"20",
		X"CD",X"35",X"13",X"FA",X"B2",X"13",X"11",X"80",X"20",X"21",X"D0",X"20",X"CD",X"1A",X"13",X"C9",
		X"11",X"C0",X"20",X"CB",X"99",X"13",X"11",X"B0",X"20",X"C3",X"99",X"13",X"11",X"A0",X"20",X"C3",
		X"99",X"13",X"11",X"90",X"20",X"C3",X"99",X"13",X"2A",X"C0",X"20",X"EB",X"2A",X"45",X"20",X"CD",
		X"39",X"13",X"D8",X"CD",X"63",X"12",X"CD",X"65",X"00",X"3A",X"01",X"21",X"B7",X"C0",X"2A",X"45",
		X"20",X"22",X"D0",X"20",X"EB",X"21",X"DB",X"20",X"CD",X"56",X"11",X"CD",X"3E",X"13",X"CD",X"4E",
		X"13",X"CD",X"06",X"12",X"CD",X"F5",X"11",X"CD",X"F5",X"11",X"CD",X"47",X"12",X"C9",X"FF",X"FF",
		X"CD",X"C7",X"11",X"21",X"D4",X"20",X"CD",X"CD",X"11",X"C9",X"3E",X"2F",X"CD",X"F7",X"11",X"C9");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
