library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_7J is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_7J is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"18",X"12",X"7D",X"7D",X"00",X"00",X"00",X"00",X"12",X"E2",X"72",X"2E",X"FE",
		X"00",X"6F",X"2F",X"31",X"0A",X"00",X"00",X"00",X"FC",X"4C",X"4E",X"A2",X"72",X"30",X"00",X"00",
		X"00",X"00",X"00",X"30",X"24",X"FA",X"FA",X"00",X"00",X"08",X"2C",X"46",X"E1",X"70",X"38",X"F8",
		X"00",X"DE",X"5E",X"62",X"34",X"00",X"00",X"00",X"F8",X"4C",X"42",X"B5",X"76",X"30",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"3C",X"00",X"00",X"00",X"00",X"10",X"30",X"30",X"62",
		X"6C",X"0D",X"13",X"67",X"33",X"39",X"0A",X"00",X"74",X"F0",X"F4",X"38",X"6E",X"38",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"3C",X"00",X"00",X"00",X"00",X"10",X"3C",X"36",X"66",
		X"6C",X"0D",X"13",X"67",X"33",X"39",X"0A",X"00",X"76",X"F6",X"B3",X"34",X"6E",X"1E",X"07",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"3C",X"00",X"00",X"00",X"00",X"14",X"39",X"37",X"67",
		X"6C",X"0D",X"13",X"67",X"33",X"39",X"0A",X"00",X"7F",X"F8",X"F8",X"38",X"6C",X"37",X"0B",X"0E",
		X"00",X"0A",X"39",X"33",X"67",X"13",X"0D",X"6C",X"00",X"00",X"38",X"6E",X"38",X"F4",X"F0",X"74",
		X"20",X"1C",X"0C",X"00",X"00",X"00",X"00",X"00",X"62",X"30",X"30",X"10",X"00",X"00",X"00",X"00",
		X"00",X"0A",X"39",X"33",X"67",X"13",X"0D",X"6C",X"00",X"07",X"1E",X"6E",X"34",X"B3",X"F6",X"76",
		X"20",X"1C",X"0C",X"00",X"00",X"00",X"00",X"00",X"66",X"36",X"3C",X"10",X"00",X"00",X"00",X"00",
		X"00",X"0A",X"39",X"33",X"67",X"13",X"0D",X"6C",X"0E",X"0B",X"37",X"6C",X"38",X"FC",X"7C",X"78",
		X"20",X"1C",X"0C",X"00",X"00",X"00",X"00",X"00",X"22",X"36",X"3A",X"16",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"07",X"04",X"04",X"00",X"00",X"00",X"00",X"60",X"F0",X"90",X"90",
		X"04",X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"90",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"1F",X"3F",X"3C",X"34",X"00",X"00",X"00",X"08",X"FC",X"FE",X"9E",X"96",
		X"34",X"3F",X"3F",X"18",X"0F",X"07",X"00",X"00",X"96",X"FE",X"FE",X"0C",X"F8",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"07",X"38",X"38",X"00",X"00",X"00",X"00",X"60",X"F0",X"00",X"00",
		X"38",X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"0F",X"0C",X"04",X"00",X"00",X"00",X"00",X"F0",X"F0",X"90",X"90",
		X"04",X"07",X"00",X"00",X"07",X"07",X"00",X"00",X"90",X"F2",X"06",X"0C",X"F8",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"04",X"04",X"04",X"00",X"00",X"00",X"00",X"10",X"90",X"90",X"90",
		X"04",X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"90",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"1F",X"3F",X"3C",X"34",X"00",X"00",X"00",X"08",X"FC",X"FE",X"9E",X"96",
		X"34",X"3F",X"3F",X"18",X"0F",X"07",X"00",X"00",X"96",X"FE",X"FE",X"0C",X"F8",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"04",X"38",X"38",X"00",X"00",X"00",X"00",X"10",X"90",X"00",X"00",
		X"38",X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"0F",X"0C",X"04",X"00",X"00",X"00",X"00",X"F0",X"F0",X"90",X"90",
		X"04",X"07",X"00",X"00",X"07",X"07",X"00",X"00",X"90",X"F2",X"06",X"0C",X"F8",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"06",X"04",X"04",X"00",X"00",X"00",X"00",X"60",X"F0",X"90",X"90",
		X"04",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"90",X"B0",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"1F",X"3F",X"3C",X"34",X"00",X"00",X"00",X"08",X"FC",X"FE",X"9E",X"96",
		X"34",X"3F",X"3B",X"18",X"0F",X"07",X"00",X"00",X"96",X"BE",X"2E",X"0C",X"F8",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"06",X"38",X"38",X"00",X"00",X"00",X"00",X"60",X"F0",X"00",X"00",
		X"38",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"0F",X"0C",X"04",X"00",X"00",X"00",X"00",X"F0",X"F0",X"90",X"90",
		X"04",X"07",X"00",X"00",X"07",X"07",X"00",X"00",X"90",X"B2",X"06",X"0C",X"F8",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"06",X"1E",X"00",X"00",X"60",X"E0",X"C0",X"DA",X"DE",X"DE",
		X"06",X"1E",X"06",X"01",X"01",X"00",X"00",X"00",X"F8",X"DE",X"DE",X"DA",X"C0",X"E0",X"60",X"00",
		X"00",X"00",X"0C",X"0E",X"07",X"05",X"06",X"36",X"00",X"00",X"00",X"00",X"00",X"D9",X"DF",X"DE",
		X"0E",X"36",X"06",X"05",X"07",X"0E",X"0C",X"00",X"F8",X"DE",X"DF",X"D9",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"38",X"78",X"FC",X"6E",X"AE",X"AA",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"B8",X"AA",X"AE",X"6E",X"FC",X"78",X"38",X"00",
		X"00",X"00",X"00",X"04",X"1E",X"06",X"00",X"0E",X"00",X"C2",X"C2",X"CE",X"DE",X"FC",X"D8",X"D0",
		X"0C",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"DA",X"DE",X"DE",X"CE",X"C4",X"E0",X"60",X"00",
		X"00",X"00",X"00",X"04",X"1E",X"06",X"00",X"0E",X"00",X"04",X"04",X"7C",X"FC",X"DA",X"5E",X"DE",
		X"0C",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"DE",X"FC",X"F8",X"78",X"00",X"00",X"00",X"00",
		X"00",X"01",X"01",X"04",X"1E",X"06",X"00",X"0E",X"00",X"82",X"C2",X"CE",X"DE",X"FC",X"58",X"D0",
		X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DA",X"5E",X"1E",X"04",X"C0",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"04",X"1E",X"06",X"00",X"0E",X"00",X"04",X"C4",X"DC",X"FC",X"DA",X"DE",X"DE",
		X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"F8",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"0C",X"00",X"60",X"E0",X"C4",X"CE",X"DE",X"DE",X"DA",
		X"0E",X"00",X"06",X"1E",X"04",X"00",X"00",X"00",X"D0",X"D8",X"FC",X"DE",X"CE",X"C2",X"C2",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"0C",X"00",X"00",X"00",X"00",X"78",X"F8",X"FC",X"DE",
		X"0E",X"00",X"06",X"1E",X"04",X"00",X"00",X"00",X"DE",X"DE",X"DA",X"FC",X"7C",X"04",X"04",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"C0",X"C0",X"04",X"1E",X"5E",X"DA",
		X"0E",X"00",X"06",X"1E",X"04",X"01",X"01",X"00",X"D0",X"D8",X"FC",X"DE",X"CE",X"C2",X"82",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"60",X"60",X"F8",X"FE",
		X"0E",X"00",X"06",X"1E",X"04",X"00",X"00",X"00",X"DE",X"DE",X"DE",X"FC",X"DC",X"C4",X"04",X"00",
		X"00",X"00",X"06",X"07",X"03",X"02",X"03",X"1B",X"00",X"00",X"00",X"00",X"80",X"ED",X"6F",X"6F",
		X"07",X"1B",X"03",X"02",X"03",X"07",X"06",X"00",X"7C",X"6F",X"6F",X"ED",X"80",X"00",X"00",X"00",
		X"00",X"00",X"03",X"03",X"01",X"01",X"01",X"03",X"00",X"00",X"00",X"80",X"C0",X"75",X"B7",X"B7",
		X"03",X"03",X"01",X"01",X"01",X"03",X"03",X"00",X"BC",X"B7",X"B7",X"75",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"04",X"36",X"04",X"01",X"07",X"06",X"40",X"E0",X"F0",X"F9",X"7D",X"EF",X"4F",X"5E",
		X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"5C",X"DC",X"9C",X"CC",X"C6",X"E3",X"C0",X"00",
		X"00",X"00",X"01",X"03",X"03",X"03",X"05",X"1F",X"04",X"C6",X"CF",X"9F",X"BE",X"BC",X"B8",X"DC",
		X"06",X"0E",X"02",X"02",X"03",X"00",X"00",X"00",X"DE",X"DE",X"DE",X"D8",X"D8",X"F8",X"78",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"C0",X"E3",X"C6",X"CC",X"9C",X"DC",X"5C",
		X"06",X"07",X"01",X"04",X"36",X"04",X"00",X"00",X"5E",X"4F",X"EF",X"7D",X"F9",X"F0",X"E0",X"40",
		X"00",X"00",X"00",X"0D",X"02",X"02",X"0E",X"07",X"00",X"78",X"F8",X"D0",X"D8",X"DE",X"DE",X"DE",
		X"1E",X"05",X"03",X"03",X"03",X"01",X"00",X"00",X"DC",X"B8",X"BC",X"BE",X"9F",X"CF",X"C6",X"04",
		X"40",X"40",X"40",X"66",X"65",X"65",X"75",X"74",X"F4",X"70",X"C0",X"00",X"80",X"00",X"00",X"00",
		X"78",X"7C",X"7D",X"7E",X"1F",X"00",X"03",X"07",X"00",X"80",X"00",X"00",X"00",X"80",X"60",X"D0",
		X"03",X"25",X"24",X"34",X"35",X"3F",X"3F",X"3F",X"E0",X"D8",X"70",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"3F",X"3E",X"1C",X"07",X"00",X"03",X"07",X"00",X"00",X"00",X"00",X"00",X"80",X"60",X"D0",
		X"03",X"01",X"00",X"02",X"00",X"00",X"00",X"00",X"80",X"C0",X"60",X"18",X"84",X"80",X"00",X"00",
		X"00",X"00",X"03",X"0C",X"07",X"00",X"03",X"07",X"00",X"00",X"00",X"00",X"00",X"80",X"20",X"D0",
		X"00",X"00",X"00",X"00",X"68",X"17",X"07",X"0F",X"00",X"00",X"00",X"00",X"00",X"80",X"FC",X"D7",
		X"07",X"1B",X"6F",X"40",X"20",X"20",X"10",X"00",X"38",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"08",X"08",X"10",X"03",X"07",X"0F",X"00",X"00",X"00",X"00",X"00",X"80",X"F8",X"D6",
		X"07",X"0B",X"07",X"00",X"10",X"08",X"04",X"00",X"38",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"00",X"00",X"10",X"03",X"07",X"0F",X"00",X"00",X"00",X"00",X"00",X"80",X"F0",X"D4",
		X"07",X"0B",X"07",X"08",X"08",X"0E",X"00",X"00",X"30",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"40",X"40",X"61",X"63",X"73",X"7B",X"7D",X"7D",X"00",X"82",X"70",X"00",X"00",X"00",X"00",X"00",
		X"59",X"7C",X"79",X"71",X"23",X"03",X"07",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"E0",X"00",
		X"00",X"07",X"03",X"23",X"71",X"79",X"7C",X"59",X"00",X"E0",X"E0",X"C0",X"80",X"00",X"00",X"00",
		X"7D",X"7D",X"7B",X"73",X"63",X"61",X"40",X"40",X"00",X"00",X"00",X"00",X"00",X"70",X"82",X"00",
		X"00",X"00",X"00",X"00",X"01",X"05",X"06",X"1E",X"00",X"00",X"40",X"E0",X"E0",X"FA",X"DE",X"DE",
		X"0E",X"1E",X"06",X"05",X"01",X"00",X"00",X"00",X"F8",X"DE",X"DE",X"FA",X"E0",X"E0",X"40",X"00",
		X"00",X"00",X"07",X"07",X"01",X"01",X"01",X"06",X"00",X"00",X"80",X"8E",X"8E",X"DC",X"DC",X"D8",
		X"06",X"1E",X"0E",X"1C",X"00",X"03",X"03",X"00",X"D8",X"F8",X"DE",X"DE",X"CE",X"C2",X"C0",X"00",
		X"00",X"00",X"0C",X"0E",X"07",X"05",X"06",X"36",X"00",X"00",X"00",X"00",X"00",X"DA",X"DE",X"DE",
		X"0E",X"36",X"06",X"05",X"07",X"0E",X"0C",X"00",X"F8",X"DE",X"DE",X"DA",X"00",X"00",X"00",X"00",
		X"00",X"03",X"01",X"01",X"18",X"7D",X"7C",X"41",X"00",X"E0",X"80",X"38",X"A0",X"58",X"C0",X"30",
		X"01",X"12",X"1A",X"0D",X"01",X"00",X"01",X"00",X"30",X"A0",X"BC",X"5C",X"28",X"E0",X"C0",X"00",
		X"00",X"03",X"01",X"01",X"18",X"7D",X"7C",X"41",X"00",X"E0",X"80",X"3F",X"A0",X"59",X"C0",X"30",
		X"01",X"12",X"1A",X"0D",X"01",X"00",X"01",X"00",X"30",X"A0",X"BC",X"5C",X"2F",X"E0",X"C0",X"00",
		X"00",X"03",X"01",X"00",X"18",X"7E",X"7F",X"47",X"00",X"E0",X"F0",X"78",X"3C",X"3C",X"18",X"90",
		X"03",X"11",X"19",X"0C",X"00",X"00",X"01",X"00",X"D0",X"F8",X"FC",X"EC",X"E8",X"C0",X"C0",X"00",
		X"00",X"07",X"1B",X"22",X"2D",X"72",X"F9",X"82",X"00",X"CA",X"04",X"78",X"40",X"B0",X"80",X"60",
		X"02",X"25",X"35",X"1A",X"02",X"01",X"03",X"00",X"68",X"44",X"7C",X"BA",X"50",X"C0",X"80",X"00",
		X"80",X"E0",X"7C",X"5E",X"2C",X"3F",X"17",X"1B",X"04",X"06",X"06",X"0F",X"8F",X"76",X"24",X"8C",
		X"0B",X"0C",X"04",X"04",X"01",X"01",X"00",X"00",X"BC",X"6C",X"34",X"DA",X"EA",X"2C",X"08",X"00",
		X"80",X"E0",X"38",X"56",X"2D",X"2E",X"17",X"1F",X"00",X"02",X"06",X"0F",X"8F",X"66",X"44",X"CC",
		X"0B",X"0C",X"04",X"04",X"00",X"00",X"00",X"00",X"BC",X"6C",X"24",X"D2",X"6A",X"6C",X"C8",X"00",
		X"80",X"E0",X"38",X"77",X"2F",X"2C",X"17",X"1B",X"00",X"00",X"02",X"06",X"8F",X"66",X"84",X"8C",
		X"0B",X"0F",X"06",X"05",X"01",X"01",X"00",X"00",X"8C",X"7C",X"14",X"2A",X"2A",X"EC",X"E8",X"00",
		X"80",X"F0",X"28",X"72",X"2D",X"28",X"1B",X"13",X"00",X"00",X"00",X"02",X"C6",X"E6",X"04",X"8C",
		X"0B",X"0E",X"04",X"04",X"01",X"01",X"00",X"00",X"BC",X"6C",X"24",X"D2",X"8A",X"8C",X"C8",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"01",X"19",X"18",X"3A",X"3A",X"00",X"00",X"80",X"80",X"98",X"38",X"60",X"00",
		X"01",X"08",X"18",X"19",X"01",X"01",X"00",X"00",X"7C",X"1C",X"18",X"98",X"80",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"07",X"0F",X"13",X"27",X"2F",X"2F",X"00",X"00",X"E0",X"10",X"88",X"C4",X"C4",X"E4",
		X"2F",X"2F",X"27",X"13",X"0F",X"07",X"00",X"00",X"E4",X"E4",X"C4",X"88",X"10",X"E0",X"00",X"00",
		X"CC",X"CC",X"C8",X"C8",X"C8",X"C8",X"C8",X"C0",X"C0",X"40",X"00",X"80",X"80",X"80",X"80",X"00",
		X"C4",X"CC",X"CC",X"4C",X"00",X"00",X"00",X"00",X"40",X"C0",X"C0",X"C0",X"00",X"00",X"00",X"00",
		X"C0",X"CC",X"CC",X"CC",X"CC",X"C0",X"C0",X"CC",X"00",X"C0",X"C0",X"C0",X"C0",X"00",X"00",X"C0",
		X"CC",X"CC",X"CC",X"C0",X"C0",X"CC",X"CC",X"CC",X"C0",X"C0",X"C0",X"00",X"00",X"C0",X"C0",X"C0",
		X"C0",X"C0",X"CC",X"CC",X"CC",X"CC",X"C0",X"C0",X"00",X"00",X"C0",X"C0",X"C0",X"C0",X"80",X"00",
		X"CC",X"CC",X"CC",X"CC",X"C0",X"C0",X"CC",X"C0",X"00",X"40",X"C0",X"C0",X"00",X"00",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"4C",X"CC",X"CC",X"C0",X"00",X"00",X"00",X"00",X"C0",X"C0",X"C0",X"C0",
		X"C0",X"C0",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"33",X"20",X"00",X"13",X"13",X"13",X"13",X"03",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",
		X"23",X"33",X"33",X"33",X"00",X"00",X"00",X"00",X"30",X"30",X"30",X"20",X"00",X"00",X"00",X"00",
		X"20",X"02",X"12",X"12",X"02",X"20",X"30",X"33",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",
		X"13",X"13",X"13",X"00",X"00",X"13",X"13",X"13",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",
		X"00",X"00",X"13",X"13",X"13",X"33",X"21",X"01",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",
		X"00",X"12",X"12",X"12",X"00",X"00",X"33",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",
		X"00",X"00",X"00",X"00",X"33",X"33",X"33",X"01",X"00",X"00",X"00",X"00",X"20",X"30",X"30",X"30",
		X"00",X"00",X"33",X"33",X"33",X"13",X"13",X"13",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",
		X"00",X"00",X"0C",X"0E",X"07",X"05",X"06",X"36",X"00",X"00",X"00",X"00",X"00",X"D9",X"DF",X"DE",
		X"0E",X"36",X"06",X"05",X"07",X"0E",X"0C",X"00",X"F8",X"DE",X"DF",X"D9",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"A0",X"D9",X"5F",X"DE",
		X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"F8",X"DE",X"5F",X"D9",X"A0",X"F0",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"1C",X"0E",X"0F",X"1B",
		X"00",X"E0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"18",X"1B",X"0F",X"0E",X"1C",X"00",X"00",X"00",
		X"00",X"00",X"01",X"01",X"00",X"16",X"1E",X"1E",X"00",X"00",X"80",X"C0",X"E0",X"E0",X"F0",X"E0",
		X"02",X"1E",X"1E",X"16",X"00",X"01",X"01",X"00",X"F0",X"E0",X"E0",X"F0",X"E0",X"C0",X"80",X"00",
		X"00",X"00",X"03",X"03",X"03",X"02",X"03",X"13",X"00",X"00",X"40",X"E0",X"F8",X"FC",X"5E",X"5E",
		X"07",X"13",X"03",X"02",X"03",X"03",X"03",X"00",X"7E",X"5E",X"5E",X"FC",X"F8",X"E0",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"00",X"3C",X"3E",X"4F",X"03",X"00",X"00",X"80",X"E0",X"30",X"18",X"88",X"CC",
		X"00",X"1C",X"1E",X"0E",X"06",X"00",X"00",X"00",X"C4",X"E4",X"74",X"74",X"30",X"30",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"20",X"11",X"09",X"03",X"08",X"1C",X"1E",X"00",X"00",X"80",X"80",X"3C",X"60",X"62",X"80",
		X"0B",X"09",X"01",X"00",X"00",X"00",X"00",X"21",X"90",X"98",X"62",X"20",X"9C",X"80",X"00",X"80",
		X"00",X"00",X"00",X"01",X"43",X"28",X"1C",X"1E",X"00",X"00",X"00",X"80",X"BC",X"30",X"40",X"81",
		X"03",X"01",X"01",X"10",X"20",X"40",X"00",X"00",X"90",X"D8",X"40",X"24",X"9C",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"08",X"1C",X"1E",X"00",X"00",X"00",X"00",X"BC",X"28",X"40",X"80",
		X"E3",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"D1",X"98",X"40",X"28",X"9C",X"00",X"00",X"00",
		X"00",X"00",X"80",X"01",X"03",X"08",X"1C",X"1E",X"00",X"00",X"00",X"80",X"BC",X"24",X"40",X"C0",
		X"03",X"09",X"09",X"28",X"40",X"00",X"00",X"00",X"90",X"99",X"00",X"30",X"9C",X"80",X"00",X"00",
		X"00",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"C0",X"20",X"00",X"00",X"00",
		X"00",X"08",X"0C",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"C0",X"20",X"00",
		X"00",X"08",X"0C",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"C0",
		X"00",X"08",X"0C",X"06",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",
		X"01",X"09",X"0C",X"06",X"00",X"00",X"00",X"00",X"C0",X"C0",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"09",X"0D",X"05",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"C0",X"20",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"0E",X"05",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"C0",X"00",X"00",
		X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"0C",X"06",X"02",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"00",
		X"00",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"C0",X"20",X"00",X"00",X"00",
		X"00",X"08",X"0C",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"00",X"3C",X"3E",X"4F",X"01",X"00",X"00",X"80",X"E0",X"30",X"18",X"88",X"4C",
		X"01",X"1C",X"1E",X"0E",X"06",X"00",X"00",X"00",X"C4",X"64",X"74",X"74",X"30",X"30",X"40",X"00",
		X"00",X"00",X"0F",X"00",X"3C",X"3E",X"4F",X"05",X"00",X"00",X"80",X"E0",X"30",X"18",X"88",X"CC",
		X"03",X"1D",X"1E",X"0E",X"06",X"00",X"00",X"00",X"C4",X"64",X"74",X"74",X"30",X"30",X"40",X"00",
		X"00",X"00",X"0F",X"00",X"3C",X"3E",X"4C",X"07",X"00",X"00",X"80",X"E0",X"30",X"18",X"88",X"CC",
		X"07",X"1B",X"1D",X"0E",X"06",X"00",X"00",X"00",X"84",X"A4",X"F4",X"74",X"30",X"30",X"40",X"00",
		X"00",X"00",X"0F",X"00",X"3C",X"3D",X"4F",X"0F",X"00",X"00",X"80",X"E0",X"30",X"98",X"C8",X"EC",
		X"07",X"17",X"1B",X"0C",X"06",X"00",X"00",X"00",X"E4",X"C4",X"F4",X"F4",X"30",X"30",X"40",X"00",
		X"00",X"00",X"06",X"04",X"18",X"1C",X"0E",X"06",X"00",X"20",X"F0",X"F0",X"E0",X"00",X"20",X"30",
		X"26",X"34",X"18",X"1C",X"0E",X"06",X"00",X"00",X"F0",X"E0",X"C0",X"20",X"20",X"10",X"E0",X"C0",
		X"00",X"00",X"06",X"08",X"18",X"1C",X"0E",X"06",X"00",X"20",X"E0",X"D0",X"E0",X"00",X"20",X"30",
		X"34",X"38",X"1C",X"1E",X"0E",X"06",X"00",X"00",X"F0",X"E0",X"C0",X"20",X"30",X"30",X"E0",X"C0",
		X"00",X"00",X"02",X"00",X"1C",X"1C",X"0E",X"26",X"00",X"20",X"F0",X"F0",X"E0",X"00",X"20",X"20",
		X"32",X"38",X"1C",X"1E",X"0E",X"06",X"00",X"00",X"D0",X"E0",X"C0",X"20",X"30",X"30",X"E0",X"C0",
		X"00",X"00",X"02",X"04",X"1C",X"1C",X"0E",X"06",X"00",X"20",X"F0",X"F0",X"E0",X"00",X"20",X"30",
		X"22",X"34",X"1C",X"1C",X"0E",X"06",X"00",X"00",X"F0",X"E0",X"C0",X"20",X"20",X"10",X"E0",X"C0",
		X"00",X"00",X"06",X"06",X"1E",X"1C",X"0C",X"26",X"00",X"20",X"E0",X"D0",X"E0",X"00",X"20",X"30",
		X"36",X"3E",X"1C",X"1C",X"0E",X"06",X"00",X"00",X"F0",X"E0",X"C0",X"20",X"30",X"30",X"E0",X"C0",
		X"00",X"00",X"06",X"0E",X"0C",X"1C",X"2E",X"26",X"00",X"20",X"F0",X"F0",X"E0",X"00",X"20",X"20",
		X"36",X"3C",X"1C",X"1C",X"0E",X"06",X"00",X"00",X"D0",X"E0",X"C0",X"20",X"30",X"30",X"E0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"07",X"0C",X"14",X"0F",X"4F",X"07",X"00",X"00",X"80",X"D0",X"28",X"90",X"C8",X"EC",
		X"03",X"1D",X"0E",X"1E",X"0E",X"04",X"00",X"00",X"C4",X"A4",X"70",X"68",X"10",X"00",X"40",X"00",
		X"00",X"00",X"0E",X"1E",X"2C",X"32",X"0F",X"62",X"00",X"00",X"80",X"E8",X"34",X"18",X"68",X"F4",
		X"60",X"1C",X"16",X"0E",X"1F",X"0F",X"02",X"00",X"F4",X"64",X"14",X"74",X"38",X"30",X"40",X"00",
		X"00",X"03",X"07",X"07",X"3B",X"3C",X"7F",X"73",X"00",X"00",X"80",X"A0",X"B0",X"00",X"98",X"BC",
		X"78",X"6C",X"1F",X"0B",X"07",X"07",X"03",X"00",X"BC",X"D8",X"64",X"F4",X"F0",X"F0",X"C0",X"00",
		X"00",X"00",X"0D",X"01",X"3C",X"3E",X"7F",X"7B",X"00",X"C0",X"E0",X"E0",X"D0",X"18",X"86",X"DE",
		X"78",X"74",X"0E",X"0E",X"05",X"01",X"00",X"00",X"CE",X"E6",X"30",X"F4",X"F0",X"F0",X"C0",X"00",
		X"00",X"00",X"0F",X"10",X"3C",X"3E",X"4F",X"0F",X"00",X"00",X"E0",X"70",X"30",X"08",X"88",X"CC",
		X"1F",X"16",X"18",X"2E",X"16",X"00",X"00",X"00",X"C4",X"E4",X"74",X"3C",X"78",X"70",X"00",X"00",
		X"00",X"00",X"07",X"0E",X"38",X"3C",X"4F",X"07",X"00",X"00",X"80",X"D0",X"18",X"0C",X"80",X"CC",
		X"07",X"1F",X"1F",X"1E",X"0E",X"04",X"00",X"00",X"CC",X"FC",X"F8",X"78",X"30",X"20",X"40",X"00",
		X"00",X"01",X"07",X"0E",X"30",X"3E",X"4F",X"03",X"00",X"00",X"80",X"E0",X"70",X"F8",X"78",X"74",
		X"1C",X"1E",X"1F",X"1F",X"0E",X"00",X"00",X"00",X"86",X"EC",X"6C",X"58",X"10",X"20",X"40",X"00",
		X"00",X"00",X"05",X"0E",X"1E",X"04",X"4F",X"03",X"00",X"00",X"B0",X"78",X"7C",X"3C",X"98",X"C4",
		X"1E",X"3F",X"1F",X"2F",X"17",X"0E",X"00",X"00",X"C4",X"E6",X"EC",X"D8",X"10",X"00",X"40",X"00",
		X"00",X"00",X"05",X"0C",X"18",X"16",X"0F",X"07",X"00",X"40",X"B0",X"B8",X"1C",X"0C",X"84",X"CC",
		X"1F",X"1F",X"1F",X"0F",X"07",X"00",X"00",X"00",X"C4",X"E4",X"E8",X"D8",X"30",X"00",X"40",X"00",
		X"00",X"07",X"04",X"07",X"00",X"07",X"04",X"07",X"00",X"C0",X"40",X"C0",X"00",X"C0",X"40",X"C0",
		X"00",X"00",X"07",X"04",X"00",X"00",X"00",X"00",X"00",X"40",X"C0",X"40",X"00",X"00",X"00",X"00",
		X"00",X"07",X"04",X"07",X"00",X"07",X"04",X"07",X"00",X"C0",X"40",X"C0",X"00",X"C0",X"40",X"C0",
		X"00",X"07",X"05",X"05",X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"07",X"04",X"07",X"00",X"07",X"04",X"07",X"00",X"C0",X"40",X"C0",X"00",X"C0",X"40",X"C0",
		X"00",X"07",X"05",X"05",X"00",X"00",X"00",X"00",X"00",X"C0",X"40",X"40",X"00",X"00",X"00",X"00",
		X"00",X"07",X"04",X"07",X"00",X"07",X"04",X"07",X"00",X"C0",X"40",X"C0",X"00",X"C0",X"40",X"C0",
		X"00",X"05",X"05",X"07",X"00",X"00",X"00",X"00",X"00",X"C0",X"40",X"40",X"00",X"00",X"00",X"00",
		X"00",X"07",X"04",X"07",X"00",X"07",X"04",X"07",X"00",X"C0",X"40",X"C0",X"00",X"C0",X"40",X"C0",
		X"00",X"05",X"05",X"07",X"00",X"00",X"00",X"00",X"00",X"C0",X"40",X"40",X"00",X"00",X"00",X"00",
		X"00",X"07",X"04",X"07",X"00",X"07",X"04",X"07",X"00",X"C0",X"40",X"C0",X"00",X"C0",X"40",X"C0",
		X"00",X"07",X"04",X"07",X"00",X"00",X"07",X"04",X"00",X"C0",X"40",X"C0",X"00",X"40",X"C0",X"40",
		X"00",X"07",X"04",X"07",X"00",X"07",X"04",X"07",X"00",X"C0",X"40",X"C0",X"00",X"C0",X"40",X"C0",
		X"00",X"07",X"05",X"07",X"00",X"00",X"00",X"00",X"00",X"C0",X"40",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"07",X"04",X"07",X"00",X"07",X"04",X"07",X"00",X"C0",X"40",X"C0",X"00",X"C0",X"40",X"C0",
		X"00",X"07",X"04",X"07",X"00",X"00",X"07",X"04",X"00",X"C0",X"40",X"C0",X"00",X"40",X"C0",X"40",
		X"00",X"07",X"04",X"07",X"00",X"07",X"04",X"07",X"00",X"C0",X"40",X"C0",X"00",X"C0",X"40",X"C0",
		X"00",X"07",X"05",X"05",X"00",X"00",X"07",X"04",X"00",X"40",X"40",X"C0",X"00",X"40",X"C0",X"40",
		X"00",X"07",X"04",X"07",X"00",X"07",X"04",X"07",X"00",X"C0",X"40",X"C0",X"00",X"C0",X"40",X"C0",
		X"00",X"07",X"04",X"07",X"00",X"07",X"05",X"05",X"00",X"C0",X"40",X"C0",X"00",X"C0",X"40",X"40",
		X"00",X"07",X"04",X"07",X"00",X"07",X"04",X"07",X"00",X"C0",X"40",X"C0",X"00",X"C0",X"40",X"C0",
		X"00",X"07",X"04",X"07",X"00",X"07",X"05",X"05",X"00",X"C0",X"40",X"C0",X"00",X"40",X"40",X"C0",
		X"00",X"07",X"04",X"07",X"00",X"07",X"04",X"07",X"00",X"C0",X"40",X"C0",X"00",X"C0",X"40",X"C0",
		X"00",X"07",X"04",X"07",X"00",X"05",X"05",X"07",X"00",X"C0",X"40",X"C0",X"00",X"C0",X"40",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"05",X"05",X"00",X"01",X"00",X"01",X"00",X"40",X"40",X"C0",X"00",X"40",X"80",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"05",X"05",X"00",X"01",X"00",X"01",X"00",X"C0",X"40",X"40",X"00",X"40",X"80",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"00",X"07",X"00",X"01",X"00",X"01",X"00",X"C0",X"80",X"80",X"00",X"40",X"80",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"05",X"05",X"07",X"00",X"01",X"00",X"01",X"00",X"C0",X"40",X"40",X"00",X"40",X"80",X"40",
		X"00",X"00",X"00",X"00",X"08",X"04",X"02",X"01",X"00",X"00",X"00",X"10",X"11",X"11",X"01",X"01",
		X"00",X"00",X"00",X"1C",X"00",X"00",X"00",X"0F",X"08",X"08",X"25",X"11",X"C9",X"20",X"03",X"3B",
		X"00",X"00",X"00",X"08",X"88",X"88",X"80",X"80",X"00",X"00",X"00",X"00",X"10",X"20",X"40",X"80",
		X"10",X"10",X"A4",X"88",X"93",X"04",X"C0",X"DC",X"00",X"00",X"00",X"38",X"00",X"00",X"00",X"F0",
		X"0F",X"00",X"00",X"00",X"1C",X"00",X"00",X"00",X"3B",X"03",X"20",X"C9",X"11",X"25",X"08",X"08",
		X"01",X"02",X"04",X"08",X"00",X"00",X"00",X"00",X"01",X"01",X"11",X"11",X"10",X"00",X"00",X"00",
		X"DC",X"C0",X"04",X"93",X"88",X"A4",X"10",X"10",X"F0",X"00",X"00",X"00",X"38",X"00",X"00",X"00",
		X"80",X"80",X"88",X"88",X"08",X"00",X"00",X"00",X"80",X"40",X"20",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"20",X"10",X"08",X"04",X"00",X"00",X"00",X"01",X"21",X"21",X"20",X"01",X"01",X"11",
		X"00",X"00",X"1C",X"01",X"00",X"00",X"00",X"73",X"90",X"48",X"20",X"80",X"40",X"00",X"00",X"80",
		X"00",X"80",X"80",X"84",X"04",X"04",X"80",X"88",X"00",X"00",X"04",X"08",X"10",X"20",X"00",X"00",
		X"89",X"12",X"04",X"01",X"02",X"00",X"00",X"00",X"00",X"00",X"1C",X"80",X"00",X"00",X"00",X"EE",
		X"77",X"00",X"00",X"00",X"01",X"38",X"00",X"00",X"00",X"00",X"00",X"40",X"80",X"20",X"48",X"91",
		X"00",X"00",X"04",X"08",X"10",X"20",X"00",X"00",X"11",X"01",X"20",X"20",X"21",X"01",X"01",X"00",
		X"01",X"00",X"00",X"02",X"01",X"04",X"12",X"09",X"CE",X"00",X"00",X"00",X"80",X"38",X"00",X"00",
		X"88",X"80",X"80",X"04",X"84",X"84",X"80",X"00",X"00",X"00",X"20",X"10",X"08",X"04",X"00",X"00",
		X"00",X"40",X"20",X"10",X"00",X"00",X"02",X"01",X"81",X"81",X"01",X"00",X"21",X"21",X"00",X"00",
		X"60",X"00",X"0C",X"00",X"00",X"00",X"00",X"EC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"81",X"81",X"00",X"84",X"84",X"00",X"00",X"00",X"02",X"04",X"08",X"00",X"00",X"40",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"30",X"00",X"00",X"00",X"00",X"37",
		X"EC",X"00",X"00",X"00",X"00",X"0C",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"02",X"00",X"00",X"10",X"20",X"40",X"00",X"00",X"00",X"21",X"21",X"00",X"81",X"81",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"37",X"00",X"00",X"00",X"00",X"30",X"00",X"06",
		X"00",X"00",X"84",X"84",X"00",X"80",X"81",X"81",X"80",X"40",X"00",X"00",X"08",X"04",X"02",X"00",
		X"00",X"40",X"20",X"10",X"00",X"00",X"00",X"00",X"81",X"81",X"01",X"00",X"00",X"00",X"00",X"00",
		X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"81",X"81",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"04",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"07",
		X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"20",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"81",X"81",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"06",
		X"00",X"00",X"00",X"00",X"00",X"80",X"81",X"81",X"00",X"00",X"00",X"00",X"08",X"04",X"02",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"9B",X"FB",X"7A",X"1B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"70",X"E0",X"C0",X"A0",X"60",X"E0",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"7A",X"FB",X"9B",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"60",X"A0",X"C0",X"E0",X"70",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"19",X"31",X"38",X"3D",X"1D",X"0D",X"0D",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"C0",X"E0",X"A0",X"60",X"60",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"1D",X"3D",X"38",X"31",X"19",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"60",X"60",X"A0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"07",X"07",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"0C",X"8C",X"D8",X"F0",X"70",X"70",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"07",X"07",X"03",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"70",X"70",X"F0",X"D8",X"8C",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"18",X"1E",X"0F",X"07",X"03",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"0E",X"1C",X"38",X"70",X"70",X"70",X"B8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"0F",X"1E",X"18",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"70",X"70",X"70",X"38",X"1C",X"0E",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"03",X"02",X"02",X"06",X"04",X"04",X"04",X"08",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"08",X"00",X"00",X"00",X"00",X"00",X"20",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"3F",X"3F",X"3F",X"1F",X"4F",X"07",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"83",X"F0",X"FE",X"FF",X"FF",X"FF",X"7F",X"7F",
		X"80",X"80",X"80",X"80",X"80",X"81",X"81",X"81",X"70",X"70",X"70",X"F8",X"FE",X"FF",X"FF",X"FF",
		X"83",X"83",X"87",X"C7",X"43",X"60",X"38",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",
		X"02",X"02",X"02",X"03",X"07",X"87",X"E3",X"F8",X"7F",X"0F",X"01",X"1C",X"1F",X"1F",X"7F",X"7F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"C0",X"80",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"80",X"80",X"00",X"C0",X"C0",X"C0",X"80",X"80",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"87",X"87",X"87",X"C3",X"C3",X"FC",X"FC",X"FC",X"FC",X"FE",X"FE",X"FE",X"FE",
		X"C3",X"E3",X"E3",X"E1",X"E1",X"E1",X"F1",X"F1",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"08",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"FF",
		X"F1",X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"78",X"0B",X"C3",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",
		X"83",X"87",X"8E",X"9E",X"9A",X"9B",X"99",X"9C",X"FB",X"FA",X"F8",X"F8",X"78",X"38",X"3F",X"9F",
		X"9C",X"9E",X"98",X"9E",X"9F",X"80",X"98",X"9C",X"8F",X"45",X"01",X"00",X"00",X"00",X"00",X"00",
		X"03",X"07",X"07",X"0F",X"0F",X"1F",X"0F",X"C1",X"F8",X"F0",X"F0",X"E0",X"E0",X"E0",X"C0",X"C0",
		X"C0",X"80",X"00",X"30",X"4C",X"46",X"43",X"40",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",
		X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"80",X"81",X"00",X"C0",X"C0",X"80",X"00",X"00",
		X"9E",X"9E",X"9C",X"9C",X"98",X"98",X"90",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
		X"42",X"82",X"06",X"06",X"07",X"0F",X"0F",X"18",X"00",X"00",X"00",X"00",X"00",X"08",X"8E",X"07",
		X"00",X"00",X"00",X"40",X"80",X"80",X"80",X"00",X"03",X"00",X"00",X"00",X"01",X"03",X"17",X"17",
		X"3E",X"20",X"00",X"30",X"7E",X"7E",X"7C",X"00",X"00",X"0F",X"00",X"00",X"00",X"08",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3C",X"FC",X"FC",X"0C",X"0E",X"0E",X"8E",X"8E",X"1F",X"0F",X"0F",X"07",X"07",X"07",X"03",X"03",
		X"8F",X"8F",X"8F",X"0F",X"0F",X"0F",X"0F",X"0F",X"01",X"01",X"01",X"00",X"80",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"60",X"78",X"0F",X"00",X"00",X"C0",X"E0",X"E0",X"00",X"00",X"00",X"00",X"00",X"04",X"0E",X"0E",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"C0",X"C0",X"C0",X"C0",X"E0",X"E0",X"E0",X"E0",
		X"0F",X"1F",X"1F",X"3F",X"3F",X"1F",X"1F",X"1F",X"F0",X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",
		X"00",X"41",X"49",X"49",X"49",X"7F",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"7F",X"38",X"1C",X"38",X"7F",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"39",X"7B",X"4F",X"46",X"44",X"7F",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"41",X"49",X"49",X"49",X"7F",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"3F",X"64",X"44",X"64",X"3F",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"4F",X"4F",X"49",X"49",X"63",X"3E",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"78",X"7C",X"0E",X"07",X"0E",X"7C",X"78",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3E",X"7F",X"41",X"41",X"41",X"7F",X"3E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"02",X"04",X"09",X"12",X"24",X"49",X"92",X"FF",X"00",X"FF",X"00",X"7F",X"80",X"3F",X"40",
		X"A4",X"A9",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"FF",X"00",X"FE",X"01",X"FC",X"02",X"80",X"40",X"20",X"90",X"48",X"24",X"92",X"49",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"25",X"95",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A9",X"A4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"92",X"49",X"24",X"12",X"09",X"04",X"02",X"01",X"40",X"3F",X"80",X"7F",X"00",X"FF",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"55",X"55",X"55",X"55",X"55",X"55",X"95",X"25",
		X"02",X"FC",X"01",X"FE",X"00",X"FF",X"00",X"FF",X"49",X"92",X"24",X"48",X"90",X"20",X"40",X"80",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"30",X"30",X"3F",X"3F",X"00",X"00",
		X"33",X"33",X"30",X"30",X"3F",X"3F",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"3F",X"3F",X"30",X"30",X"33",X"33",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"00",X"00",X"3F",X"3F",X"30",X"30",X"33",X"33",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"CC",X"CC",X"0C",X"0C",X"FC",X"FC",X"00",X"00",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"CC",X"CC",X"0C",X"0C",X"FC",X"FC",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FC",X"FC",X"0C",X"0C",X"CC",X"CC",
		X"00",X"00",X"FC",X"FC",X"0C",X"0C",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"9F",X"9F",X"9F",X"9F",X"9F",X"9C",X"80",X"80",X"F0",X"F0",X"F1",X"F7",X"87",X"03",X"03",X"00",
		X"80",X"80",X"81",X"87",X"9F",X"9F",X"9F",X"9F",X"0C",X"3E",X"FE",X"F8",X"FA",X"FB",X"FB",X"FB",
		X"04",X"3C",X"FC",X"FC",X"F8",X"E0",X"80",X"00",X"80",X"F0",X"C1",X"07",X"1E",X"3C",X"78",X"11",
		X"06",X"0E",X"06",X"00",X"00",X"F8",X"E0",X"C1",X"03",X"00",X"0F",X"00",X"00",X"00",X"F8",X"F8",
		X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"FB",X"FB",X"F8",X"F8",X"E0",X"C0",X"80",X"01",
		X"9C",X"98",X"80",X"80",X"80",X"80",X"80",X"81",X"03",X"07",X"0F",X"1E",X"3E",X"78",X"FB",X"FB",
		X"83",X"07",X"0F",X"1F",X"3F",X"7F",X"1F",X"C6",X"F0",X"F0",X"E1",X"C3",X"83",X"07",X"0E",X"0F",
		X"F0",X"FC",X"E0",X"00",X"00",X"00",X"81",X"03",X"1F",X"3E",X"3E",X"06",X"3C",X"FC",X"F8",X"F8",
		X"00",X"00",X"80",X"98",X"3F",X"7A",X"F6",X"F6",X"A8",X"28",X"28",X"28",X"68",X"68",X"4C",X"4C",
		X"EC",X"4C",X"08",X"00",X"00",X"00",X"00",X"60",X"CC",X"CC",X"CC",X"CC",X"0C",X"04",X"00",X"00",
		X"3C",X"1F",X"4F",X"27",X"23",X"31",X"38",X"3C",X"3F",X"0F",X"C3",X"F0",X"FC",X"FE",X"F8",X"40",
		X"3C",X"3E",X"1F",X"1F",X"1F",X"0F",X"0F",X"07",X"00",X"0E",X"0F",X"07",X"43",X"41",X"60",X"70",
		X"E3",X"E3",X"C3",X"C3",X"87",X"87",X"07",X"07",X"80",X"8E",X"8E",X"8E",X"8E",X"8F",X"0F",X"0F",
		X"00",X"08",X"0E",X"0F",X"1F",X"1F",X"1E",X"1E",X"0F",X"00",X"00",X"00",X"00",X"08",X"0E",X"0F",
		X"07",X"07",X"03",X"03",X"01",X"01",X"01",X"00",X"78",X"7C",X"7C",X"3E",X"1F",X"1F",X"00",X"FF",
		X"70",X"70",X"F0",X"30",X"08",X"08",X"08",X"B8",X"FF",X"7F",X"7F",X"7F",X"3F",X"3F",X"1F",X"1F",
		X"9F",X"9F",X"9F",X"9F",X"9F",X"8F",X"83",X"81",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"80",X"80",X"80",X"80",X"98",X"9E",X"9F",X"9F",X"7F",X"3F",X"0F",X"03",X"00",X"00",X"C0",X"F0",
		X"01",X"00",X"80",X"C0",X"E0",X"F0",X"F8",X"FC",X"FF",X"FF",X"FF",X"7F",X"3F",X"1F",X"1F",X"0F",
		X"FE",X"FF",X"FF",X"FF",X"FF",X"3F",X"0F",X"07",X"07",X"03",X"81",X"C1",X"E0",X"F0",X"F8",X"FC",
		X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"FC",X"FF",X"FF",X"FF",X"FE",X"FC",X"FD",X"F9",
		X"80",X"80",X"80",X"80",X"9F",X"9F",X"9F",X"9F",X"7B",X"00",X"00",X"00",X"F7",X"F7",X"F7",X"F0",
		X"00",X"80",X"80",X"04",X"00",X"00",X"C0",X"F8",X"7E",X"1F",X"07",X"02",X"00",X"00",X"03",X"01",
		X"FF",X"3F",X"00",X"00",X"FC",X"FC",X"C0",X"00",X"80",X"F8",X"1F",X"00",X"9F",X"00",X"07",X"06",
		X"07",X"87",X"87",X"C7",X"C3",X"C3",X"E3",X"E2",X"D0",X"D1",X"D1",X"D1",X"D1",X"81",X"81",X"00",
		X"E0",X"F0",X"F0",X"F8",X"F8",X"78",X"7C",X"3C",X"60",X"70",X"33",X"33",X"33",X"33",X"33",X"33",
		X"03",X"00",X"C0",X"E0",X"C0",X"C0",X"C3",X"47",X"00",X"00",X"10",X"1E",X"10",X"03",X"01",X"00",
		X"06",X"06",X"10",X"00",X"07",X"00",X"00",X"00",X"10",X"3C",X"7E",X"7C",X"18",X"C1",X"01",X"00",
		X"E0",X"80",X"00",X"04",X"62",X"32",X"88",X"E4",X"B2",X"B2",X"96",X"96",X"D4",X"55",X"55",X"54",
		X"7A",X"1C",X"C2",X"00",X"FF",X"02",X"00",X"09",X"55",X"55",X"38",X"17",X"C0",X"21",X"98",X"48",
		X"60",X"EF",X"DE",X"BC",X"F9",X"73",X"E6",X"CC",X"00",X"00",X"20",X"78",X"E0",X"81",X"1F",X"F8",
		X"9B",X"40",X"80",X"C6",X"00",X"C7",X"47",X"11",X"80",X"03",X"7F",X"07",X"00",X"FC",X"FE",X"FF",
		X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"8F",X"8F",X"87",X"83",X"81",X"80",X"80",X"80",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",
		X"E0",X"F0",X"F0",X"F8",X"F8",X"F8",X"FC",X"FC",X"07",X"07",X"07",X"07",X"03",X"03",X"03",X"03",
		X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"01",X"01",X"01",X"00",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"90",X"98",X"9C",X"3F",X"1F",X"0F",X"0F",X"07",X"03",X"01",X"00",
		X"9E",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"00",X"00",X"80",X"C0",X"E0",X"F0",X"F8",X"FC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C0",X"C0",X"E0",X"E0",X"E0",X"F0",X"F0",X"F8",
		X"FF",X"7F",X"3F",X"1F",X"0F",X"0F",X"07",X"03",X"F8",X"F8",X"FC",X"FC",X"FE",X"FE",X"FE",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"70",X"70",X"70",X"60",X"00",X"90",X"30",X"70",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"70",X"70",X"70",X"30",X"B0",X"90",X"D0",X"C0",
		X"0F",X"0F",X"1F",X"1F",X"1F",X"03",X"00",X"00",X"E0",X"E0",X"E0",X"E0",X"C0",X"C0",X"00",X"C0",
		X"01",X"13",X"07",X"07",X"01",X"00",X"00",X"30",X"FF",X"FE",X"F8",X"F0",X"F8",X"3C",X"02",X"00",
		X"7F",X"7F",X"7F",X"7F",X"3F",X"3F",X"3F",X"3F",X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"1F",X"1F",X"1F",X"1F",X"0F",X"0F",X"0F",X"0F",X"C0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",
		X"3E",X"3E",X"7E",X"7E",X"7C",X"7C",X"1C",X"04",X"00",X"00",X"07",X"07",X"07",X"0F",X"0F",X"1F",
		X"00",X"78",X"D8",X"C8",X"C0",X"E0",X"F0",X"F6",X"1F",X"1F",X"00",X"3F",X"5E",X"0C",X"08",X"00",
		X"0F",X"38",X"60",X"43",X"C7",X"8F",X"9F",X"9F",X"FF",X"00",X"00",X"00",X"00",X"80",X"80",X"80",
		X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"C0",X"C0",X"E0",X"E0",X"E0",X"F0",X"F0",X"F8",
		X"FF",X"00",X"00",X"07",X"03",X"03",X"03",X"03",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"F8",X"F8",X"FC",X"FC",X"FE",X"FE",X"FE",X"FF",
		X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"7F",X"7F",X"7F",X"3F",X"3F",X"3F",X"3F",
		X"00",X"80",X"80",X"80",X"C0",X"C0",X"E0",X"E0",X"1F",X"1F",X"1F",X"1F",X"0F",X"0F",X"0F",X"0F",
		X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"F0",X"F0",X"C0",X"C0",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"40",X"60",X"70",X"70",X"70",X"70",X"70",X"70",
		X"FF",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"01",X"01",X"03",X"03",X"03",X"03",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"70",X"70",X"10",X"C0",X"E0",X"F0",X"F0",X"C0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C0",X"00",X"60",X"70",X"70",X"70",X"70",X"70",
		X"00",X"00",X"00",X"04",X"06",X"07",X"07",X"07",X"7F",X"3F",X"0E",X"04",X"00",X"80",X"C4",X"EC",
		X"07",X"07",X"07",X"01",X"00",X"0F",X"0F",X"0F",X"F8",X"F8",X"F8",X"F8",X"70",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"0D",X"00",X"00",X"78",X"E4",X"92",X"86",X"09",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"60",X"F0",X"96",X"8B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"14",X"28",X"28",X"24",X"02",X"03",X"05",X"06",X"90",X"01",X"40",X"88",X"88",X"45",X"37",X"87",
		X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CD",X"38",X"01",X"03",X"00",X"00",X"00",X"00",
		X"91",X"05",X"0A",X"26",X"98",X"80",X"08",X"18",X"08",X"A0",X"60",X"00",X"00",X"00",X"00",X"00",
		X"A0",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"04",X"02",X"42",X"23",X"1F",X"0C",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"10",X"30",X"E0",X"BF",X"06",X"0C",X"18",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"06",X"0C",X"19",X"3F",X"02",X"02",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"03",X"8F",X"DC",X"78",X"34",X"22",X"01",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"42",X"00",X"40",X"00",
		X"00",X"00",X"09",X"00",X"00",X"02",X"00",X"24",X"00",X"04",X"00",X"00",X"20",X"02",X"00",X"88",
		X"00",X"00",X"00",X"40",X"00",X"00",X"02",X"90",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",
		X"00",X"00",X"10",X"82",X"00",X"00",X"50",X"00",X"00",X"20",X"00",X"00",X"88",X"00",X"00",X"02",
		X"00",X"10",X"00",X"01",X"00",X"10",X"02",X"00",X"02",X"00",X"10",X"00",X"40",X"01",X"00",X"00",
		X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"81",X"08",X"00",X"40",X"08",X"00",X"01",X"00",
		X"04",X"01",X"40",X"00",X"00",X"08",X"00",X"00",X"10",X"00",X"00",X"08",X"00",X"40",X"00",X"00",
		X"10",X"00",X"04",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
