`define BUILD_DATE "180915"
`define BUILD_TIME "160403"
