library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_PGM_1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_PGM_1 is
	type rom is array(0 to  12287) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"53",X"22",X"00",X"10",X"5B",X"74",X"89",X"44",X"95",X"5A",X"53",X"17",X"F0",X"AC",X"E4",X"00",
		X"5C",X"A8",X"53",X"17",X"D8",X"EC",X"3F",X"DE",X"17",X"AA",X"A8",X"3F",X"C4",X"22",X"10",X"22",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E4",X"68",X"5A",X"5B",X"32",X"8B",X"5B",X"3C",
		X"5C",X"AC",X"00",X"EC",X"EC",X"82",X"D2",X"02",X"22",X"00",X"10",X"17",X"F8",X"89",X"5C",X"FB",
		X"C0",X"BD",X"B5",X"9E",X"B1",X"91",X"00",X"42",X"89",X"B7",X"CA",X"0D",X"B5",X"D0",X"B1",X"A0",
		X"B5",X"FE",X"BD",X"B5",X"60",X"BD",X"B3",X"00",X"00",X"42",X"B5",X"FE",X"BD",X"B5",X"28",X"BD",
		X"A9",X"B7",X"E0",X"0D",X"B5",X"80",X"BD",X"B5",X"FF",X"B5",X"D4",X"BD",X"B3",X"00",X"30",X"B7",
		X"28",X"B1",X"81",X"00",X"42",X"B5",X"FE",X"BD",X"4B",X"0D",X"B5",X"FE",X"B1",X"44",X"00",X"8C",
		X"66",X"0B",X"54",X"0B",X"72",X"0B",X"F8",X"0B",X"43",X"09",X"F8",X"0B",X"89",X"0B",X"90",X"05",
		X"92",X"09",X"7A",X"09",X"5F",X"09",X"FB",X"09",X"90",X"05",X"90",X"05",X"90",X"05",X"90",X"05",
		X"90",X"05",X"90",X"05",X"90",X"05",X"90",X"05",X"FF",X"B3",X"00",X"00",X"B7",X"BA",X"0D",X"B5",
		X"90",X"05",X"90",X"05",X"08",X"0D",X"90",X"05",X"02",X"B1",X"00",X"00",X"8C",X"B3",X"EB",X"94",
		X"00",X"B1",X"0E",X"FF",X"B3",X"00",X"89",X"B7",X"B5",X"FE",X"BD",X"FF",X"C6",X"C6",X"C2",X"C2",
		X"12",X"0D",X"B5",X"B4",X"B1",X"80",X"00",X"42",X"C6",X"C6",X"A4",X"A4",X"FF",X"C7",X"C7",X"C3",
		X"FF",X"AF",X"AF",X"6B",X"6B",X"AF",X"AF",X"6F",X"B7",X"B7",X"FF",X"A8",X"A8",X"A2",X"A2",X"A8",
		X"6F",X"FF",X"AC",X"AC",X"B3",X"B3",X"AC",X"AC",X"A8",X"A6",X"A6",X"FF",X"29",X"29",X"29",X"2B",
		X"6F",X"A4",X"99",X"5A",X"53",X"00",X"00",X"24",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"64",X"80",X"5A",X"5B",X"DC",X"8B",X"82",X"10",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"B3",X"FF",X"FE",X"B7",X"E0",X"0D",X"B5",X"D0",X"20",X"BD",X"B3",X"00",X"98",X"B7",X"CA",X"0D",
		X"B1",X"91",X"00",X"42",X"B5",X"FE",X"BD",X"B5",X"B5",X"20",X"B1",X"B0",X"00",X"42",X"B3",X"FF",
		X"B5",X"FE",X"B1",X"80",X"00",X"8C",X"B5",X"A0",X"B3",X"00",X"30",X"B7",X"4F",X"0D",X"B5",X"74",
		X"B1",X"80",X"00",X"8C",X"FF",X"B5",X"7E",X"BD",X"B1",X"44",X"00",X"8C",X"B5",X"FE",X"B1",X"80",
		X"90",X"05",X"A1",X"0B",X"90",X"05",X"90",X"05",X"59",X"0B",X"90",X"05",X"90",X"05",X"90",X"05",
		X"90",X"05",X"90",X"05",X"90",X"05",X"90",X"05",X"90",X"05",X"90",X"05",X"90",X"05",X"71",X"0B",
		X"B5",X"60",X"BD",X"B5",X"8C",X"B1",X"00",X"00",X"88",X"0D",X"B5",X"FE",X"B1",X"B1",X"00",X"42",
		X"8C",X"B5",X"8C",X"BD",X"B3",X"FF",X"98",X"B7",X"B5",X"FE",X"B1",X"B1",X"00",X"42",X"B3",X"00",
		X"C3",X"C7",X"C7",X"A5",X"A5",X"FF",X"7C",X"7C",X"7D",X"D5",X"D5",X"7D",X"7D",X"B5",X"B5",X"FF",
		X"D4",X"D4",X"7C",X"7C",X"B4",X"B4",X"FF",X"7D",X"AE",X"AE",X"6A",X"6A",X"AE",X"AE",X"6E",X"6E",
		X"2B",X"2B",X"FF",X"28",X"28",X"28",X"2A",X"2A",X"FF",X"CE",X"FF",X"CC",X"FF",X"80",X"80",X"80",
		X"2A",X"FF",X"2C",X"2C",X"2C",X"2E",X"2E",X"2E",X"88",X"88",X"88",X"8C",X"8C",X"8C",X"FF",X"82",
		X"00",X"10",X"17",X"03",X"89",X"5C",X"FB",X"22",X"5A",X"5B",X"32",X"8B",X"5B",X"3C",X"62",X"24",
		X"AC",X"4A",X"CC",X"53",X"17",X"C9",X"0D",X"53",X"A4",X"93",X"5A",X"22",X"69",X"5C",X"57",X"BD",
		X"F0",X"FD",X"04",X"EC",X"CE",X"17",X"01",X"8B",X"95",X"17",X"8F",X"8F",X"DB",X"22",X"59",X"5C",
		X"5A",X"17",X"1B",X"0D",X"53",X"E0",X"40",X"CC",X"42",X"0E",X"FB",X"AA",X"00",X"53",X"0C",X"C2",
		X"00",X"8C",X"B5",X"E4",X"B1",X"80",X"00",X"8C",X"00",X"8C",X"B3",X"EB",X"34",X"B5",X"D4",X"BD",
		X"FF",X"B7",X"43",X"0D",X"B5",X"02",X"B1",X"00",X"B3",X"0A",X"30",X"B7",X"C1",X"0D",X"B5",X"FE",
		X"06",X"8C",X"B7",X"C5",X"0D",X"B5",X"02",X"B1",X"00",X"00",X"B7",X"BA",X"0D",X"B5",X"02",X"B1",
		X"00",X"00",X"8C",X"B5",X"20",X"BD",X"FF",X"B3",X"00",X"00",X"8C",X"B3",X"EB",X"94",X"B5",X"60",
		X"FE",X"B7",X"CA",X"0D",X"B5",X"BA",X"B1",X"80",X"B7",X"2C",X"0D",X"B5",X"A0",X"B1",X"00",X"B1",
		X"00",X"42",X"B5",X"08",X"B1",X"80",X"B1",X"42",X"42",X"B7",X"CA",X"0D",X"B5",X"80",X"B1",X"00",
		X"98",X"B7",X"D8",X"0D",X"B5",X"6E",X"BD",X"B5",X"79",X"00",X"0A",X"B3",X"00",X"FE",X"B7",X"36",
		X"B0",X"B1",X"7F",X"00",X"0A",X"B5",X"B8",X"B1",X"0D",X"B5",X"C8",X"BD",X"B5",X"D0",X"B1",X"8C",
		X"82",X"82",X"8A",X"8A",X"8A",X"8E",X"8E",X"8E",X"C0",X"C0",X"C0",X"68",X"68",X"68",X"68",X"FF",
		X"FF",X"84",X"FF",X"86",X"FF",X"A0",X"FF",X"C0",X"0E",X"FF",X"4E",X"FF",X"E4",X"42",X"5A",X"3D",
		X"A8",X"A4",X"44",X"58",X"53",X"E4",X"42",X"5A",X"1E",X"20",X"04",X"EC",X"AA",X"A4",X"44",X"58",
		X"3D",X"0E",X"57",X"EE",X"CC",X"69",X"07",X"57",X"53",X"E4",X"40",X"5A",X"3D",X"0E",X"57",X"EE",
		X"40",X"5C",X"17",X"72",X"A8",X"ED",X"24",X"48",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"40",X"5A",X"82",X"89",X"01",X"17",X"C0",X"41",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"83",X"5C",X"22",X"FA",X"8D",X"DB",X"22",X"D9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"37",X"8B",X"23",X"66",X"BA",X"2C",X"A5",X"2C",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"B1",X"44",X"00",X"8C",X"B5",X"FE",X"B1",X"0C",X"B5",X"48",X"B1",X"06",X"42",X"8C",X"B5",X"0A",
		X"48",X"8C",X"B5",X"0C",X"B1",X"0C",X"B1",X"8C",X"B1",X"0A",X"BD",X"8C",X"B5",X"44",X"B1",X"08",
		X"BD",X"B5",X"8C",X"B1",X"00",X"00",X"8C",X"B5",X"B5",X"02",X"B1",X"00",X"00",X"42",X"B3",X"11",
		X"8C",X"BD",X"B3",X"00",X"00",X"B7",X"E0",X"0D",X"11",X"B5",X"A0",X"BD",X"FF",X"B3",X"00",X"00",
		X"00",X"42",X"FF",X"B3",X"00",X"00",X"B7",X"FE",X"6B",X"94",X"B5",X"60",X"BD",X"B5",X"8C",X"B1",
		X"0D",X"B5",X"02",X"B1",X"00",X"00",X"8C",X"B3",X"00",X"00",X"8C",X"B5",X"8C",X"BD",X"B3",X"FF",
		X"00",X"0A",X"BB",X"80",X"B5",X"0C",X"B1",X"F1",X"B5",X"0C",X"B1",X"F1",X"F1",X"0A",X"B5",X"0C",
		X"F1",X"0A",X"B5",X"0C",X"B1",X"F1",X"40",X"0A",X"B1",X"F1",X"40",X"0A",X"B3",X"00",X"00",X"B7",
		X"0E",X"57",X"EE",X"6E",X"CC",X"A0",X"07",X"57",X"53",X"E4",X"40",X"5A",X"3D",X"0E",X"57",X"EE",
		X"1E",X"20",X"04",X"EC",X"AE",X"A4",X"44",X"58",X"CC",X"A0",X"07",X"57",X"1E",X"20",X"04",X"EC",
		X"6E",X"CC",X"B9",X"07",X"57",X"1E",X"20",X"04",X"5A",X"2F",X"11",X"E4",X"99",X"5A",X"2F",X"55",
		X"EC",X"AC",X"A4",X"44",X"58",X"53",X"E4",X"29",X"1E",X"0F",X"E4",X"95",X"5A",X"2F",X"55",X"1E",
		X"40",X"00",X"8C",X"00",X"02",X"00",X"04",X"00",X"90",X"00",X"90",X"86",X"76",X"34",X"C6",X"57",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"A4",X"E9",X"5C",X"C0",X"0C",X"A4",X"59",X"5C",
		X"A8",X"5C",X"17",X"79",X"89",X"7B",X"21",X"82",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"17",X"7E",X"AC",X"00",X"04",X"53",X"6F",X"04",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"B7",X"FE",X"0D",X"B5",X"02",X"B1",X"00",X"00",X"8C",X"B1",X"00",X"00",X"8C",X"B5",X"8C",X"BD",
		X"8C",X"B3",X"6B",X"94",X"B5",X"60",X"BD",X"B5",X"B3",X"00",X"00",X"B7",X"88",X"0D",X"B5",X"02",
		X"00",X"00",X"8C",X"B5",X"8C",X"BD",X"B3",X"00",X"B5",X"02",X"B1",X"00",X"00",X"8C",X"B3",X"6B",
		X"00",X"FF",X"B3",X"00",X"00",X"B7",X"FE",X"0D",X"94",X"B5",X"60",X"BD",X"B5",X"8C",X"B1",X"00",
		X"B6",X"0D",X"B5",X"02",X"B1",X"00",X"00",X"06",X"06",X"FF",X"B5",X"D4",X"BD",X"B3",X"00",X"29",
		X"B3",X"FE",X"E4",X"B5",X"10",X"B1",X"00",X"00",X"B7",X"12",X"0D",X"B5",X"FE",X"B1",X"80",X"00",
		X"B1",X"42",X"B7",X"E0",X"0D",X"B5",X"80",X"B1",X"02",X"29",X"B7",X"36",X"0D",X"B5",X"6E",X"BD",
		X"00",X"00",X"42",X"FF",X"B5",X"DE",X"BD",X"B3",X"B5",X"B0",X"B1",X"82",X"00",X"06",X"B5",X"B8",
		X"0F",X"E4",X"12",X"58",X"1E",X"22",X"12",X"41",X"5A",X"22",X"12",X"58",X"A8",X"FC",X"3D",X"4E",
		X"DF",X"7B",X"D6",X"95",X"5A",X"C2",X"24",X"95",X"11",X"22",X"10",X"58",X"AA",X"F5",X"AB",X"0F",
		X"0E",X"0E",X"0E",X"A4",X"12",X"58",X"53",X"E4",X"A1",X"11",X"22",X"4A",X"5C",X"17",X"D6",X"0F",
		X"4C",X"5C",X"FD",X"10",X"55",X"D0",X"0F",X"FD",X"22",X"48",X"5C",X"FC",X"2F",X"11",X"A8",X"E4",
		X"18",X"17",X"28",X"8B",X"20",X"04",X"EC",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"B6",X"04",X"17",X"5C",X"AC",X"48",X"DB",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"2F",X"7B",X"94",X"11",X"6F",X"00",X"E8",X"A4",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"B1",X"00",X"00",X"42",X"B3",X"91",X"11",X"B5",X"0D",X"B5",X"02",X"B1",X"00",X"00",X"8C",X"B3",
		X"A0",X"BD",X"FF",X"B3",X"00",X"00",X"B7",X"BA",X"EB",X"94",X"B5",X"60",X"BD",X"B5",X"8C",X"B1",
		X"00",X"8C",X"B5",X"8C",X"BD",X"B3",X"00",X"00",X"00",X"8C",X"B3",X"EB",X"34",X"B5",X"D4",X"BD",
		X"FF",X"B7",X"43",X"0D",X"B5",X"02",X"B1",X"00",X"B3",X"00",X"00",X"FF",X"B7",X"47",X"0D",X"B5",
		X"42",X"B5",X"FE",X"B1",X"80",X"00",X"42",X"B3",X"B1",X"00",X"42",X"B5",X"08",X"B1",X"B1",X"B1",
		X"FF",X"FE",X"B7",X"E0",X"0D",X"B5",X"BC",X"B1",X"42",X"B7",X"54",X"0D",X"B5",X"A0",X"B1",X"00",
		X"B1",X"88",X"00",X"06",X"B3",X"FF",X"FE",X"B7",X"75",X"00",X"06",X"B5",X"0C",X"B1",X"40",X"F1",
		X"D8",X"0D",X"B5",X"C8",X"BD",X"B5",X"D0",X"B1",X"06",X"B5",X"0C",X"B1",X"40",X"40",X"06",X"B5",
		X"FC",X"9E",X"57",X"EE",X"57",X"EE",X"22",X"E9",X"EC",X"06",X"25",X"60",X"0E",X"57",X"E2",X"57",
		X"5C",X"57",X"7D",X"64",X"14",X"58",X"9F",X"5E",X"E2",X"EA",X"20",X"F3",X"EC",X"06",X"23",X"0E",
		X"86",X"5C",X"FD",X"0E",X"E0",X"44",X"0C",X"0E",X"22",X"CB",X"0F",X"1E",X"0F",X"01",X"9F",X"A4",
		X"7B",X"DE",X"3D",X"CE",X"81",X"A0",X"FB",X"01",X"48",X"58",X"26",X"FC",X"A4",X"4A",X"58",X"26",
		X"3B",X"22",X"38",X"10",X"17",X"08",X"8B",X"7B",X"64",X"4C",X"5A",X"5B",X"D2",X"8B",X"82",X"10",
		X"53",X"17",X"A3",X"0D",X"53",X"0E",X"FD",X"0C",X"2D",X"57",X"1F",X"BE",X"53",X"17",X"7D",X"0D",
		X"C4",X"17",X"17",X"8B",X"0C",X"0C",X"DB",X"22",X"E4",X"86",X"5C",X"E8",X"17",X"87",X"0F",X"6C",
		X"40",X"5A",X"17",X"D3",X"0D",X"53",X"E0",X"0A",X"5C",X"17",X"23",X"89",X"00",X"22",X"08",X"5C",
		X"02",X"B1",X"00",X"00",X"8C",X"B3",X"6B",X"34",X"B3",X"00",X"00",X"FF",X"B3",X"00",X"89",X"B7",
		X"B5",X"E2",X"BD",X"BF",X"B5",X"CC",X"BD",X"F1",X"36",X"0D",X"B5",X"B0",X"B1",X"80",X"00",X"02",
		X"00",X"06",X"B7",X"74",X"0D",X"B5",X"E0",X"B1",X"36",X"0D",X"B5",X"B0",X"B1",X"80",X"00",X"0A",
		X"00",X"B1",X"06",X"FF",X"B3",X"00",X"89",X"B7",X"B5",X"90",X"B1",X"80",X"00",X"0A",X"B7",X"74",
		X"0C",X"B1",X"40",X"F1",X"06",X"B5",X"0C",X"B1",X"B1",X"00",X"00",X"8C",X"FF",X"B5",X"D4",X"BD",
		X"40",X"40",X"06",X"B7",X"B2",X"0D",X"B5",X"80",X"B3",X"FF",X"A8",X"B7",X"88",X"0D",X"B5",X"FE",
		X"F9",X"FE",X"B7",X"88",X"0D",X"B5",X"C0",X"BD",X"BD",X"B5",X"C0",X"BD",X"B3",X"00",X"98",X"B7",
		X"B5",X"70",X"B1",X"D1",X"00",X"42",X"B5",X"FE",X"12",X"0D",X"B5",X"20",X"B1",X"B0",X"00",X"42",
		X"FC",X"A4",X"99",X"5A",X"22",X"F1",X"0F",X"5B",X"95",X"5A",X"53",X"FD",X"40",X"D5",X"F3",X"66",
		X"5B",X"0F",X"26",X"DC",X"26",X"9C",X"7B",X"96",X"EC",X"0E",X"17",X"F3",X"66",X"00",X"88",X"0C",
		X"58",X"82",X"40",X"41",X"AE",X"EE",X"7B",X"94",X"72",X"30",X"7B",X"DE",X"3D",X"06",X"1E",X"0F",
		X"20",X"26",X"22",X"00",X"41",X"5B",X"EB",X"89",X"0F",X"01",X"9F",X"DE",X"26",X"9C",X"7B",X"96",
		X"5C",X"17",X"5E",X"A8",X"12",X"3F",X"15",X"22",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"5B",X"00",X"80",X"C0",X"0E",X"C8",X"5B",X"14",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"A4",X"8D",X"5C",X"22",X"4B",X"8D",X"DB",X"22",X"92",X"05",X"27",X"05",X"84",X"07",X"58",X"07",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"72",X"0B",X"F8",X"0B",X"8B",X"07",X"B1",X"07",
		X"B5",X"90",X"B1",X"80",X"00",X"02",X"B7",X"74",X"B3",X"00",X"89",X"B7",X"36",X"0D",X"B5",X"B0",
		X"0D",X"B5",X"50",X"B1",X"00",X"B1",X"02",X"FF",X"B1",X"80",X"00",X"06",X"B5",X"90",X"B1",X"80",
		X"0D",X"B5",X"60",X"B1",X"00",X"B1",X"0A",X"FF",X"B1",X"80",X"00",X"0E",X"B5",X"90",X"B1",X"80",
		X"B3",X"00",X"89",X"B7",X"36",X"0D",X"B5",X"B0",X"00",X"0E",X"B7",X"74",X"0D",X"B5",X"C0",X"B1",
		X"BD",X"B5",X"28",X"BD",X"B5",X"70",X"B1",X"D1",X"B3",X"00",X"89",X"B7",X"12",X"0D",X"B5",X"70",
		X"00",X"42",X"B5",X"FE",X"BD",X"B5",X"C0",X"BD",X"B1",X"60",X"00",X"42",X"B5",X"FE",X"BD",X"B3",
		X"B3",X"FF",X"A9",X"B7",X"88",X"0D",X"B5",X"80",X"B5",X"36",X"BD",X"B3",X"FF",X"A8",X"B7",X"E0",
		X"BD",X"B5",X"28",X"B1",X"81",X"00",X"42",X"FF",X"0D",X"B5",X"28",X"BD",X"B5",X"FE",X"BD",X"B5",
		X"02",X"4E",X"0E",X"04",X"8A",X"40",X"06",X"0E",X"8C",X"48",X"0E",X"00",X"4A",X"E4",X"97",X"5A",
		X"42",X"08",X"88",X"44",X"0A",X"8A",X"46",X"0C",X"1D",X"20",X"FD",X"10",X"E0",X"94",X"64",X"14",
		X"14",X"58",X"26",X"FC",X"A4",X"10",X"58",X"EC",X"24",X"14",X"58",X"EC",X"CA",X"17",X"39",X"0F",
		X"CE",X"A4",X"12",X"58",X"53",X"22",X"40",X"41",X"5E",X"47",X"10",X"4D",X"C4",X"83",X"44",X"89",
		X"53",X"22",X"00",X"10",X"5B",X"74",X"89",X"44",X"95",X"5A",X"53",X"17",X"F0",X"AC",X"E4",X"00",
		X"5C",X"A8",X"53",X"17",X"D8",X"EC",X"3F",X"DE",X"17",X"AA",X"A8",X"3F",X"C4",X"22",X"10",X"22",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E4",X"68",X"5A",X"5B",X"32",X"8B",X"5B",X"3C",
		X"5C",X"AC",X"00",X"EC",X"EC",X"82",X"D2",X"02",X"22",X"00",X"10",X"17",X"F8",X"89",X"5C",X"FB",
		X"C0",X"BD",X"B5",X"9E",X"B1",X"91",X"00",X"42",X"89",X"B7",X"CA",X"0D",X"B5",X"D0",X"B1",X"A0",
		X"B5",X"FE",X"BD",X"B5",X"60",X"BD",X"B3",X"00",X"00",X"42",X"B5",X"FE",X"BD",X"B5",X"28",X"BD",
		X"A9",X"B7",X"E0",X"0D",X"B5",X"80",X"BD",X"B5",X"FF",X"B5",X"D4",X"BD",X"B3",X"00",X"30",X"B7",
		X"28",X"B1",X"81",X"00",X"42",X"B5",X"FE",X"BD",X"4B",X"0D",X"B5",X"FE",X"B1",X"44",X"00",X"8C",
		X"66",X"0B",X"54",X"0B",X"72",X"0B",X"F8",X"0B",X"43",X"09",X"F8",X"0B",X"89",X"0B",X"90",X"05",
		X"92",X"09",X"7A",X"09",X"5F",X"09",X"FB",X"09",X"90",X"05",X"90",X"05",X"90",X"05",X"90",X"05",
		X"90",X"05",X"90",X"05",X"90",X"05",X"90",X"05",X"FF",X"B3",X"00",X"00",X"B7",X"BA",X"0D",X"B5",
		X"90",X"05",X"90",X"05",X"08",X"0D",X"90",X"05",X"02",X"B1",X"00",X"00",X"8C",X"B3",X"EB",X"94",
		X"00",X"B1",X"0E",X"FF",X"B3",X"00",X"89",X"B7",X"B5",X"FE",X"BD",X"FF",X"C6",X"C6",X"C2",X"C2",
		X"12",X"0D",X"B5",X"B4",X"B1",X"80",X"00",X"42",X"C6",X"C6",X"A4",X"A4",X"FF",X"C7",X"C7",X"C3",
		X"FF",X"AF",X"AF",X"6B",X"6B",X"AF",X"AF",X"6F",X"B7",X"B7",X"FF",X"A8",X"A8",X"A2",X"A2",X"A8",
		X"6F",X"FF",X"AC",X"AC",X"B3",X"B3",X"AC",X"AC",X"A8",X"A6",X"A6",X"FF",X"29",X"29",X"29",X"2B",
		X"6F",X"A4",X"99",X"5A",X"53",X"00",X"00",X"24",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"64",X"80",X"5A",X"5B",X"DC",X"8B",X"82",X"10",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"B3",X"FF",X"FE",X"B7",X"E0",X"0D",X"B5",X"D0",X"20",X"BD",X"B3",X"00",X"98",X"B7",X"CA",X"0D",
		X"B1",X"91",X"00",X"42",X"B5",X"FE",X"BD",X"B5",X"B5",X"20",X"B1",X"B0",X"00",X"42",X"B3",X"FF",
		X"B5",X"FE",X"B1",X"80",X"00",X"8C",X"B5",X"A0",X"B3",X"00",X"30",X"B7",X"4F",X"0D",X"B5",X"74",
		X"B1",X"80",X"00",X"8C",X"FF",X"B5",X"7E",X"BD",X"B1",X"44",X"00",X"8C",X"B5",X"FE",X"B1",X"80",
		X"90",X"05",X"A1",X"0B",X"90",X"05",X"90",X"05",X"59",X"0B",X"90",X"05",X"90",X"05",X"90",X"05",
		X"90",X"05",X"90",X"05",X"90",X"05",X"90",X"05",X"90",X"05",X"90",X"05",X"90",X"05",X"71",X"0B",
		X"B5",X"60",X"BD",X"B5",X"8C",X"B1",X"00",X"00",X"88",X"0D",X"B5",X"FE",X"B1",X"B1",X"00",X"42",
		X"8C",X"B5",X"8C",X"BD",X"B3",X"FF",X"98",X"B7",X"B5",X"FE",X"B1",X"B1",X"00",X"42",X"B3",X"00",
		X"C3",X"C7",X"C7",X"A5",X"A5",X"FF",X"7C",X"7C",X"7D",X"D5",X"D5",X"7D",X"7D",X"B5",X"B5",X"FF",
		X"D4",X"D4",X"7C",X"7C",X"B4",X"B4",X"FF",X"7D",X"AE",X"AE",X"6A",X"6A",X"AE",X"AE",X"6E",X"6E",
		X"2B",X"2B",X"FF",X"28",X"28",X"28",X"2A",X"2A",X"FF",X"CE",X"FF",X"CC",X"FF",X"80",X"80",X"80",
		X"2A",X"FF",X"2C",X"2C",X"2C",X"2E",X"2E",X"2E",X"88",X"88",X"88",X"8C",X"8C",X"8C",X"FF",X"82",
		X"00",X"10",X"17",X"03",X"89",X"5C",X"FB",X"22",X"5A",X"5B",X"32",X"8B",X"5B",X"3C",X"62",X"24",
		X"AC",X"4A",X"CC",X"53",X"17",X"C9",X"0D",X"53",X"A4",X"93",X"5A",X"22",X"69",X"5C",X"57",X"BD",
		X"F0",X"FD",X"04",X"EC",X"CE",X"17",X"01",X"8B",X"95",X"17",X"8F",X"8F",X"DB",X"22",X"59",X"5C",
		X"5A",X"17",X"1B",X"0D",X"53",X"E0",X"40",X"CC",X"42",X"0E",X"FB",X"AA",X"00",X"53",X"0C",X"C2",
		X"00",X"8C",X"B5",X"E4",X"B1",X"80",X"00",X"8C",X"00",X"8C",X"B3",X"EB",X"34",X"B5",X"D4",X"BD",
		X"FF",X"B7",X"43",X"0D",X"B5",X"02",X"B1",X"00",X"B3",X"0A",X"30",X"B7",X"C1",X"0D",X"B5",X"FE",
		X"06",X"8C",X"B7",X"C5",X"0D",X"B5",X"02",X"B1",X"00",X"00",X"B7",X"BA",X"0D",X"B5",X"02",X"B1",
		X"00",X"00",X"8C",X"B5",X"20",X"BD",X"FF",X"B3",X"00",X"00",X"8C",X"B3",X"EB",X"94",X"B5",X"60",
		X"FE",X"B7",X"CA",X"0D",X"B5",X"BA",X"B1",X"80",X"B7",X"2C",X"0D",X"B5",X"A0",X"B1",X"00",X"B1",
		X"00",X"42",X"B5",X"08",X"B1",X"80",X"B1",X"42",X"42",X"B7",X"CA",X"0D",X"B5",X"80",X"B1",X"00",
		X"98",X"B7",X"D8",X"0D",X"B5",X"6E",X"BD",X"B5",X"79",X"00",X"0A",X"B3",X"00",X"FE",X"B7",X"36",
		X"B0",X"B1",X"7F",X"00",X"0A",X"B5",X"B8",X"B1",X"0D",X"B5",X"C8",X"BD",X"B5",X"D0",X"B1",X"8C",
		X"82",X"82",X"8A",X"8A",X"8A",X"8E",X"8E",X"8E",X"C0",X"C0",X"C0",X"68",X"68",X"68",X"68",X"FF",
		X"FF",X"84",X"FF",X"86",X"FF",X"A0",X"FF",X"C0",X"0E",X"FF",X"4E",X"FF",X"E4",X"42",X"5A",X"3D",
		X"A8",X"A4",X"44",X"58",X"53",X"E4",X"42",X"5A",X"1E",X"20",X"04",X"EC",X"AA",X"A4",X"44",X"58",
		X"3D",X"0E",X"57",X"EE",X"CC",X"69",X"07",X"57",X"53",X"E4",X"40",X"5A",X"3D",X"0E",X"57",X"EE",
		X"40",X"5C",X"17",X"72",X"A8",X"ED",X"24",X"48",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"40",X"5A",X"82",X"89",X"01",X"17",X"C0",X"41",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"83",X"5C",X"22",X"FA",X"8D",X"DB",X"22",X"D9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"37",X"8B",X"23",X"66",X"BA",X"2C",X"A5",X"2C",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"B1",X"44",X"00",X"8C",X"B5",X"FE",X"B1",X"0C",X"B5",X"48",X"B1",X"06",X"42",X"8C",X"B5",X"0A",
		X"48",X"8C",X"B5",X"0C",X"B1",X"0C",X"B1",X"8C",X"B1",X"0A",X"BD",X"8C",X"B5",X"44",X"B1",X"08",
		X"BD",X"B5",X"8C",X"B1",X"00",X"00",X"8C",X"B5",X"B5",X"02",X"B1",X"00",X"00",X"42",X"B3",X"11",
		X"8C",X"BD",X"B3",X"00",X"00",X"B7",X"E0",X"0D",X"11",X"B5",X"A0",X"BD",X"FF",X"B3",X"00",X"00",
		X"00",X"42",X"FF",X"B3",X"00",X"00",X"B7",X"FE",X"6B",X"94",X"B5",X"60",X"BD",X"B5",X"8C",X"B1",
		X"0D",X"B5",X"02",X"B1",X"00",X"00",X"8C",X"B3",X"00",X"00",X"8C",X"B5",X"8C",X"BD",X"B3",X"FF",
		X"00",X"0A",X"BB",X"80",X"B5",X"0C",X"B1",X"F1",X"B5",X"0C",X"B1",X"F1",X"F1",X"0A",X"B5",X"0C",
		X"F1",X"0A",X"B5",X"0C",X"B1",X"F1",X"40",X"0A",X"B1",X"F1",X"40",X"0A",X"B3",X"00",X"00",X"B7",
		X"0E",X"57",X"EE",X"6E",X"CC",X"A0",X"07",X"57",X"53",X"E4",X"40",X"5A",X"3D",X"0E",X"57",X"EE",
		X"1E",X"20",X"04",X"EC",X"AE",X"A4",X"44",X"58",X"CC",X"A0",X"07",X"57",X"1E",X"20",X"04",X"EC",
		X"6E",X"CC",X"B9",X"07",X"57",X"1E",X"20",X"04",X"5A",X"2F",X"11",X"E4",X"99",X"5A",X"2F",X"55",
		X"EC",X"AC",X"A4",X"44",X"58",X"53",X"E4",X"29",X"1E",X"0F",X"E4",X"95",X"5A",X"2F",X"55",X"1E",
		X"40",X"00",X"8C",X"00",X"02",X"00",X"04",X"00",X"90",X"00",X"90",X"86",X"76",X"34",X"C6",X"57",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"A4",X"E9",X"5C",X"C0",X"0C",X"A4",X"59",X"5C",
		X"A8",X"5C",X"17",X"79",X"89",X"7B",X"21",X"82",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"17",X"7E",X"AC",X"00",X"04",X"53",X"6F",X"04",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"B7",X"FE",X"0D",X"B5",X"02",X"B1",X"00",X"00",X"8C",X"B1",X"00",X"00",X"8C",X"B5",X"8C",X"BD",
		X"8C",X"B3",X"6B",X"94",X"B5",X"60",X"BD",X"B5",X"B3",X"00",X"00",X"B7",X"88",X"0D",X"B5",X"02",
		X"00",X"00",X"8C",X"B5",X"8C",X"BD",X"B3",X"00",X"B5",X"02",X"B1",X"00",X"00",X"8C",X"B3",X"6B",
		X"00",X"FF",X"B3",X"00",X"00",X"B7",X"FE",X"0D",X"94",X"B5",X"60",X"BD",X"B5",X"8C",X"B1",X"00",
		X"B6",X"0D",X"B5",X"02",X"B1",X"00",X"00",X"06",X"06",X"FF",X"B5",X"D4",X"BD",X"B3",X"00",X"29",
		X"B3",X"FE",X"E4",X"B5",X"10",X"B1",X"00",X"00",X"B7",X"12",X"0D",X"B5",X"FE",X"B1",X"80",X"00",
		X"B1",X"42",X"B7",X"E0",X"0D",X"B5",X"80",X"B1",X"02",X"29",X"B7",X"36",X"0D",X"B5",X"6E",X"BD",
		X"00",X"00",X"42",X"FF",X"B5",X"DE",X"BD",X"B3",X"B5",X"B0",X"B1",X"82",X"00",X"06",X"B5",X"B8",
		X"0F",X"E4",X"12",X"58",X"1E",X"22",X"12",X"41",X"5A",X"22",X"12",X"58",X"A8",X"FC",X"3D",X"4E",
		X"DF",X"7B",X"D6",X"95",X"5A",X"C2",X"24",X"95",X"11",X"22",X"10",X"58",X"AA",X"F5",X"AB",X"0F",
		X"0E",X"0E",X"0E",X"A4",X"12",X"58",X"53",X"E4",X"A1",X"11",X"22",X"4A",X"5C",X"17",X"D6",X"0F",
		X"4C",X"5C",X"FD",X"10",X"55",X"D0",X"0F",X"FD",X"22",X"48",X"5C",X"FC",X"2F",X"11",X"A8",X"E4",
		X"18",X"17",X"28",X"8B",X"20",X"04",X"EC",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"B6",X"04",X"17",X"5C",X"AC",X"48",X"DB",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"2F",X"7B",X"94",X"11",X"6F",X"00",X"E8",X"A4",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"B1",X"00",X"00",X"42",X"B3",X"91",X"11",X"B5",X"0D",X"B5",X"02",X"B1",X"00",X"00",X"8C",X"B3",
		X"A0",X"BD",X"FF",X"B3",X"00",X"00",X"B7",X"BA",X"EB",X"94",X"B5",X"60",X"BD",X"B5",X"8C",X"B1",
		X"00",X"8C",X"B5",X"8C",X"BD",X"B3",X"00",X"00",X"00",X"8C",X"B3",X"EB",X"34",X"B5",X"D4",X"BD",
		X"FF",X"B7",X"43",X"0D",X"B5",X"02",X"B1",X"00",X"B3",X"00",X"00",X"FF",X"B7",X"47",X"0D",X"B5",
		X"42",X"B5",X"FE",X"B1",X"80",X"00",X"42",X"B3",X"B1",X"00",X"42",X"B5",X"08",X"B1",X"B1",X"B1",
		X"FF",X"FE",X"B7",X"E0",X"0D",X"B5",X"BC",X"B1",X"42",X"B7",X"54",X"0D",X"B5",X"A0",X"B1",X"00",
		X"B1",X"88",X"00",X"06",X"B3",X"FF",X"FE",X"B7",X"75",X"00",X"06",X"B5",X"0C",X"B1",X"40",X"F1",
		X"D8",X"0D",X"B5",X"C8",X"BD",X"B5",X"D0",X"B1",X"06",X"B5",X"0C",X"B1",X"40",X"40",X"06",X"B5",
		X"FC",X"9E",X"57",X"EE",X"57",X"EE",X"22",X"E9",X"EC",X"06",X"25",X"60",X"0E",X"57",X"E2",X"57",
		X"5C",X"57",X"7D",X"64",X"14",X"58",X"9F",X"5E",X"E2",X"EA",X"20",X"F3",X"EC",X"06",X"23",X"0E",
		X"86",X"5C",X"FD",X"0E",X"E0",X"44",X"0C",X"0E",X"22",X"CB",X"0F",X"1E",X"0F",X"01",X"9F",X"A4",
		X"7B",X"DE",X"3D",X"CE",X"81",X"A0",X"FB",X"01",X"48",X"58",X"26",X"FC",X"A4",X"4A",X"58",X"26",
		X"3B",X"22",X"38",X"10",X"17",X"08",X"8B",X"7B",X"64",X"4C",X"5A",X"5B",X"D2",X"8B",X"82",X"10",
		X"53",X"17",X"A3",X"0D",X"53",X"0E",X"FD",X"0C",X"2D",X"57",X"1F",X"BE",X"53",X"17",X"7D",X"0D",
		X"C4",X"17",X"17",X"8B",X"0C",X"0C",X"DB",X"22",X"E4",X"86",X"5C",X"E8",X"17",X"87",X"0F",X"6C",
		X"40",X"5A",X"17",X"D3",X"0D",X"53",X"E0",X"0A",X"5C",X"17",X"23",X"89",X"00",X"22",X"08",X"5C",
		X"02",X"B1",X"00",X"00",X"8C",X"B3",X"6B",X"34",X"B3",X"00",X"00",X"FF",X"B3",X"00",X"89",X"B7",
		X"B5",X"E2",X"BD",X"BF",X"B5",X"CC",X"BD",X"F1",X"36",X"0D",X"B5",X"B0",X"B1",X"80",X"00",X"02",
		X"00",X"06",X"B7",X"74",X"0D",X"B5",X"E0",X"B1",X"36",X"0D",X"B5",X"B0",X"B1",X"80",X"00",X"0A",
		X"00",X"B1",X"06",X"FF",X"B3",X"00",X"89",X"B7",X"B5",X"90",X"B1",X"80",X"00",X"0A",X"B7",X"74",
		X"0C",X"B1",X"40",X"F1",X"06",X"B5",X"0C",X"B1",X"B1",X"00",X"00",X"8C",X"FF",X"B5",X"D4",X"BD",
		X"40",X"40",X"06",X"B7",X"B2",X"0D",X"B5",X"80",X"B3",X"FF",X"A8",X"B7",X"88",X"0D",X"B5",X"FE",
		X"F9",X"FE",X"B7",X"88",X"0D",X"B5",X"C0",X"BD",X"BD",X"B5",X"C0",X"BD",X"B3",X"00",X"98",X"B7",
		X"B5",X"70",X"B1",X"D1",X"00",X"42",X"B5",X"FE",X"12",X"0D",X"B5",X"20",X"B1",X"B0",X"00",X"42",
		X"FC",X"A4",X"99",X"5A",X"22",X"F1",X"0F",X"5B",X"95",X"5A",X"53",X"FD",X"40",X"D5",X"F3",X"66",
		X"5B",X"0F",X"26",X"DC",X"26",X"9C",X"7B",X"96",X"EC",X"0E",X"17",X"F3",X"66",X"00",X"88",X"0C",
		X"58",X"82",X"40",X"41",X"AE",X"EE",X"7B",X"94",X"72",X"30",X"7B",X"DE",X"3D",X"06",X"1E",X"0F",
		X"20",X"26",X"22",X"00",X"41",X"5B",X"EB",X"89",X"0F",X"01",X"9F",X"DE",X"26",X"9C",X"7B",X"96",
		X"5C",X"17",X"5E",X"A8",X"12",X"3F",X"15",X"22",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"5B",X"00",X"80",X"C0",X"0E",X"C8",X"5B",X"14",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"A4",X"8D",X"5C",X"22",X"4B",X"8D",X"DB",X"22",X"92",X"05",X"27",X"05",X"84",X"07",X"58",X"07",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"72",X"0B",X"F8",X"0B",X"8B",X"07",X"B1",X"07",
		X"B5",X"90",X"B1",X"80",X"00",X"02",X"B7",X"74",X"B3",X"00",X"89",X"B7",X"36",X"0D",X"B5",X"B0",
		X"0D",X"B5",X"50",X"B1",X"00",X"B1",X"02",X"FF",X"B1",X"80",X"00",X"06",X"B5",X"90",X"B1",X"80",
		X"0D",X"B5",X"60",X"B1",X"00",X"B1",X"0A",X"FF",X"B1",X"80",X"00",X"0E",X"B5",X"90",X"B1",X"80",
		X"B3",X"00",X"89",X"B7",X"36",X"0D",X"B5",X"B0",X"00",X"0E",X"B7",X"74",X"0D",X"B5",X"C0",X"B1",
		X"BD",X"B5",X"28",X"BD",X"B5",X"70",X"B1",X"D1",X"B3",X"00",X"89",X"B7",X"12",X"0D",X"B5",X"70",
		X"00",X"42",X"B5",X"FE",X"BD",X"B5",X"C0",X"BD",X"B1",X"60",X"00",X"42",X"B5",X"FE",X"BD",X"B3",
		X"B3",X"FF",X"A9",X"B7",X"88",X"0D",X"B5",X"80",X"B5",X"36",X"BD",X"B3",X"FF",X"A8",X"B7",X"E0",
		X"BD",X"B5",X"28",X"B1",X"81",X"00",X"42",X"FF",X"0D",X"B5",X"28",X"BD",X"B5",X"FE",X"BD",X"B5",
		X"02",X"4E",X"0E",X"04",X"8A",X"40",X"06",X"0E",X"8C",X"48",X"0E",X"00",X"4A",X"E4",X"97",X"5A",
		X"42",X"08",X"88",X"44",X"0A",X"8A",X"46",X"0C",X"1D",X"20",X"FD",X"10",X"E0",X"94",X"64",X"14",
		X"14",X"58",X"26",X"FC",X"A4",X"10",X"58",X"EC",X"24",X"14",X"58",X"EC",X"CA",X"17",X"39",X"0F",
		X"CE",X"A4",X"12",X"58",X"53",X"22",X"40",X"41",X"5E",X"47",X"10",X"4D",X"C4",X"83",X"44",X"89",
		X"04",X"5D",X"F9",X"F9",X"F9",X"D5",X"04",X"3D",X"B9",X"39",X"04",X"D9",X"00",X"00",X"00",X"00",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"0A",X"06",X"46",X"06",X"06",X"06",X"08",X"0A",
		X"06",X"02",X"02",X"02",X"02",X"02",X"46",X"0C",X"80",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"4E",X"44",X"06",X"08",X"4E",X"44",X"02",X"02",X"02",X"02",X"0E",X"08",X"48",X"06",X"06",X"06",
		X"08",X"02",X"02",X"02",X"02",X"02",X"00",X"00",X"10",X"20",X"38",X"10",X"F0",X"10",X"09",X"16",
		X"83",X"CC",X"98",X"B9",X"A8",X"83",X"CC",X"98",X"67",X"F5",X"65",X"65",X"75",X"FF",X"9E",X"9A",
		X"EF",X"65",X"9C",X"83",X"24",X"00",X"00",X"DE",X"00",X"7E",X"83",X"60",X"00",X"00",X"0A",X"00",
		X"00",X"00",X"61",X"44",X"61",X"EF",X"F5",X"67",X"12",X"9A",X"00",X"21",X"04",X"10",X"BB",X"9E",
		X"C9",X"16",X"CA",X"24",X"10",X"20",X"CA",X"E2",X"89",X"CA",X"49",X"B9",X"66",X"89",X"64",X"B8",
		X"ED",X"F5",X"65",X"00",X"90",X"FB",X"9A",X"BB",X"FB",X"8A",X"90",X"02",X"90",X"9A",X"75",X"6F",
		X"00",X"9C",X"89",X"C0",X"00",X"00",X"D8",X"89",X"9A",X"90",X"12",X"9A",X"FB",X"65",X"65",X"21",
		X"21",X"65",X"65",X"9A",X"DE",X"02",X"00",X"90",X"22",X"00",X"10",X"53",X"13",X"41",X"6D",X"47",
		X"27",X"20",X"B9",X"53",X"22",X"C8",X"8B",X"5B",X"26",X"1C",X"26",X"44",X"84",X"86",X"EC",X"06",
		X"84",X"83",X"F5",X"87",X"1B",X"9B",X"22",X"C8",X"9C",X"77",X"57",X"99",X"E4",X"FC",X"18",X"ED",
		X"26",X"9C",X"57",X"95",X"84",X"26",X"DC",X"26",X"57",X"95",X"84",X"93",X"13",X"EC",X"80",X"ED",
		X"5A",X"BB",X"1B",X"3B",X"22",X"F0",X"8B",X"5B",X"9F",X"DE",X"26",X"9C",X"33",X"13",X"B3",X"53",
		X"04",X"3F",X"77",X"04",X"DD",X"39",X"04",X"3F",X"BB",X"39",X"04",X"3F",X"77",X"04",X"3D",X"75",
		X"0A",X"DD",X"39",X"46",X"DD",X"39",X"0A",X"DD",X"39",X"04",X"3D",X"71",X"71",X"B9",X"B5",X"71",
		X"04",X"DD",X"39",X"04",X"3D",X"71",X"71",X"B9",X"77",X"04",X"3F",X"73",X"73",X"BB",X"B7",X"73",
		X"04",X"3F",X"77",X"04",X"3F",X"73",X"73",X"BB",X"40",X"DD",X"39",X"40",X"DD",X"39",X"04",X"D9",
		X"02",X"02",X"0E",X"02",X"02",X"02",X"02",X"02",X"0E",X"0A",X"06",X"02",X"02",X"02",X"08",X"08",
		X"02",X"02",X"02",X"06",X"02",X"02",X"02",X"02",X"02",X"06",X"08",X"08",X"4E",X"06",X"0C",X"08",
		X"02",X"02",X"02",X"02",X"48",X"02",X"02",X"02",X"08",X"0E",X"84",X"06",X"08",X"06",X"02",X"02",
		X"8C",X"0E",X"06",X"8C",X"0E",X"06",X"02",X"02",X"84",X"06",X"08",X"0E",X"84",X"06",X"08",X"02",
		X"3D",X"A0",X"FD",X"A0",X"F0",X"11",X"EC",X"20",X"5B",X"2E",X"8D",X"33",X"13",X"53",X"42",X"20",
		X"BD",X"12",X"42",X"26",X"8C",X"14",X"FF",X"FC",X"DC",X"26",X"9C",X"84",X"F0",X"57",X"95",X"84",
		X"5E",X"53",X"7F",X"C8",X"86",X"7F",X"C8",X"AA",X"00",X"02",X"00",X"08",X"BE",X"42",X"AC",X"02",
		X"02",X"7B",X"14",X"26",X"9D",X"08",X"BE",X"42",X"42",X"AC",X"02",X"7B",X"14",X"C2",X"1D",X"46",
		X"9C",X"98",X"92",X"76",X"72",X"76",X"72",X"76",X"B8",X"B2",X"B8",X"B2",X"76",X"72",X"2D",X"2D",
		X"04",X"B0",X"3C",X"B0",X"1C",X"90",X"0D",X"81",X"3C",X"B0",X"1C",X"90",X"0D",X"81",X"B0",X"32",
		X"29",X"25",X"23",X"B9",X"02",X"0D",X"43",X"47",X"00",X"B5",X"04",X"B7",X"44",X"B9",X"00",X"3A",
		X"0B",X"38",X"0B",X"74",X"72",X"74",X"49",X"BA",X"B2",X"FF",X"B3",X"04",X"B5",X"06",X"B7",X"44",
		X"02",X"02",X"02",X"02",X"02",X"02",X"48",X"06",X"0E",X"8A",X"08",X"02",X"02",X"02",X"02",X"02",
		X"0E",X"08",X"48",X"06",X"06",X"06",X"0E",X"08",X"08",X"48",X"02",X"02",X"02",X"06",X"02",X"02",
		X"02",X"02",X"02",X"4E",X"44",X"06",X"80",X"02",X"08",X"06",X"80",X"0C",X"06",X"08",X"06",X"02",
		X"0A",X"06",X"46",X"02",X"02",X"02",X"06",X"06",X"02",X"04",X"02",X"02",X"06",X"02",X"02",X"02",
		X"95",X"95",X"95",X"95",X"99",X"F9",X"F9",X"D5",X"F9",X"91",X"95",X"95",X"95",X"95",X"95",X"95",
		X"D5",X"04",X"DD",X"39",X"04",X"D9",X"F9",X"F9",X"3D",X"71",X"71",X"71",X"71",X"75",X"04",X"3F",
		X"95",X"95",X"95",X"95",X"77",X"04",X"3D",X"71",X"3F",X"73",X"73",X"73",X"BB",X"39",X"0E",X"DD",
		X"D9",X"F9",X"D5",X"0C",X"DD",X"39",X"04",X"3D",X"04",X"3D",X"71",X"71",X"75",X"04",X"DD",X"39",
		X"06",X"22",X"85",X"28",X"3B",X"22",X"C3",X"89",X"42",X"22",X"00",X"10",X"DB",X"22",X"8C",X"5C",
		X"85",X"1B",X"22",X"AB",X"89",X"5B",X"EB",X"89",X"77",X"40",X"17",X"3B",X"40",X"68",X"47",X"8E",
		X"3B",X"FD",X"4A",X"B5",X"99",X"89",X"22",X"DF",X"5C",X"26",X"1C",X"53",X"9D",X"4A",X"9D",X"40",
		X"00",X"02",X"02",X"02",X"04",X"04",X"04",X"04",X"EB",X"89",X"82",X"A8",X"5C",X"72",X"30",X"5C",
		X"55",X"33",X"28",X"E4",X"04",X"5C",X"2F",X"60",X"E4",X"86",X"5C",X"FD",X"8A",X"B5",X"27",X"8B",
		X"17",X"33",X"28",X"9D",X"8A",X"9D",X"80",X"B5",X"8C",X"8C",X"8C",X"88",X"88",X"88",X"88",X"0E",
		X"CA",X"CA",X"CA",X"E4",X"86",X"5C",X"FD",X"06",X"89",X"22",X"00",X"18",X"44",X"06",X"2F",X"55",
		X"47",X"60",X"4D",X"F0",X"FD",X"44",X"59",X"46",X"59",X"E8",X"8D",X"17",X"DC",X"68",X"1B",X"3B",
		X"75",X"04",X"DD",X"39",X"04",X"79",X"97",X"97",X"71",X"71",X"75",X"04",X"DD",X"39",X"04",X"D9",
		X"77",X"04",X"3F",X"77",X"04",X"D9",X"F9",X"F9",X"73",X"BB",X"39",X"04",X"3F",X"77",X"04",X"D9",
		X"F9",X"F9",X"D5",X"40",X"DD",X"39",X"0A",X"D9",X"71",X"71",X"71",X"75",X"04",X"5D",X"F9",X"F9",
		X"04",X"DD",X"39",X"04",X"3D",X"71",X"71",X"B9",X"02",X"02",X"02",X"4E",X"02",X"02",X"02",X"04",
		X"02",X"02",X"02",X"02",X"02",X"06",X"08",X"08",X"08",X"08",X"02",X"02",X"02",X"06",X"02",X"02",
		X"02",X"02",X"02",X"06",X"08",X"08",X"06",X"06",X"02",X"06",X"06",X"0E",X"0A",X"06",X"02",X"02",
		X"02",X"02",X"02",X"02",X"0C",X"08",X"0E",X"4E",X"4E",X"02",X"02",X"02",X"04",X"02",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"8D",X"D0",X"E8",X"5E",X"8F",X"AD",X"8D",X"C2",X"8F",X"8D",X"8F",X"8D",X"8F",X"B3",X"00",X"B5",
		X"0D",X"45",X"41",X"47",X"74",X"76",X"B2",X"74",X"B6",X"BA",X"8D",X"8B",X"8D",X"FF",X"B3",X"04",
		X"0D",X"81",X"03",X"81",X"0D",X"81",X"70",X"74",X"3A",X"70",X"0D",X"03",X"0D",X"FF",X"B3",X"00",
		X"72",X"0D",X"32",X"38",X"3A",X"0D",X"0D",X"38",X"38",X"38",X"23",X"B0",X"B2",X"B8",X"BA",X"AA",
		X"3C",X"3A",X"81",X"32",X"B0",X"32",X"3A",X"70",X"0B",X"B0",X"0D",X"70",X"3A",X"FF",X"FF",X"E4",
		X"58",X"22",X"90",X"5E",X"02",X"48",X"00",X"7B",X"60",X"48",X"E4",X"44",X"58",X"FD",X"EE",X"20",
		X"8D",X"17",X"19",X"68",X"FF",X"FF",X"FF",X"FF",X"1E",X"1A",X"5C",X"1A",X"94",X"12",X"58",X"20",
		X"20",X"20",X"16",X"5E",X"94",X"90",X"5E",X"94",X"50",X"3A",X"78",X"78",X"7E",X"68",X"20",X"5C",
		X"71",X"71",X"B9",X"39",X"04",X"3D",X"71",X"71",X"34",X"02",X"04",X"02",X"02",X"06",X"02",X"02",
		X"02",X"08",X"02",X"02",X"02",X"02",X"02",X"08",X"06",X"46",X"02",X"02",X"02",X"06",X"06",X"08",
		X"06",X"08",X"06",X"80",X"0C",X"06",X"08",X"06",X"02",X"02",X"08",X"06",X"02",X"02",X"02",X"02",
		X"02",X"08",X"48",X"02",X"02",X"02",X"06",X"02",X"0E",X"08",X"48",X"06",X"06",X"06",X"08",X"02",
		X"00",X"B5",X"10",X"6A",X"CA",X"24",X"CA",X"E2",X"C1",X"16",X"6C",X"83",X"8A",X"98",X"48",X"A8",
		X"B9",X"E8",X"83",X"8A",X"98",X"48",X"75",X"FF",X"9A",X"9B",X"9E",X"9A",X"65",X"65",X"EF",X"F5",
		X"83",X"2A",X"00",X"00",X"DE",X"83",X"2A",X"00",X"00",X"98",X"0A",X"98",X"FE",X"BB",X"46",X"44",
		X"65",X"65",X"05",X"65",X"00",X"21",X"65",X"9A",X"EF",X"10",X"F9",X"91",X"95",X"95",X"95",X"95",
		X"10",X"E6",X"CC",X"89",X"88",X"49",X"48",X"26",X"B9",X"AC",X"89",X"8A",X"B8",X"48",X"01",X"65",
		X"9B",X"9E",X"9A",X"75",X"FF",X"9E",X"9B",X"DE",X"FD",X"64",X"61",X"65",X"90",X"89",X"8A",X"00",
		X"C2",X"00",X"00",X"36",X"89",X"C8",X"00",X"00",X"05",X"65",X"FD",X"65",X"65",X"6F",X"04",X"64",
		X"9A",X"EF",X"22",X"B8",X"89",X"5B",X"EB",X"89",X"61",X"4D",X"F2",X"83",X"22",X"96",X"28",X"C0",
		X"EB",X"89",X"82",X"A8",X"5C",X"72",X"30",X"5C",X"27",X"20",X"B9",X"53",X"AA",X"47",X"20",X"4D",
		X"8B",X"5B",X"EB",X"89",X"30",X"72",X"DC",X"26",X"20",X"04",X"EC",X"00",X"BE",X"77",X"26",X"DC",
		X"9C",X"57",X"95",X"84",X"26",X"DC",X"26",X"9C",X"53",X"E4",X"6C",X"5A",X"C0",X"06",X"E4",X"6E",
		X"EB",X"89",X"72",X"30",X"7B",X"DE",X"3D",X"0C",X"6A",X"47",X"C0",X"4D",X"44",X"83",X"04",X"89",
		X"73",X"73",X"73",X"73",X"77",X"04",X"3F",X"73",X"04",X"D9",X"F9",X"D5",X"04",X"DD",X"11",X"39",
		X"39",X"04",X"D9",X"F9",X"D5",X"04",X"DD",X"11",X"71",X"75",X"04",X"3D",X"71",X"71",X"71",X"75",
		X"39",X"04",X"D9",X"F9",X"D5",X"04",X"3F",X"73",X"73",X"77",X"04",X"3F",X"73",X"73",X"BB",X"39",
		X"39",X"04",X"D9",X"F9",X"D5",X"42",X"DD",X"39",X"F9",X"D5",X"04",X"3D",X"71",X"71",X"71",X"71",
		X"0C",X"08",X"02",X"02",X"02",X"02",X"06",X"06",X"06",X"06",X"0E",X"0A",X"06",X"06",X"08",X"08",
		X"02",X"02",X"02",X"02",X"02",X"06",X"02",X"02",X"08",X"4E",X"06",X"0C",X"08",X"02",X"02",X"02",
		X"02",X"02",X"02",X"06",X"08",X"0E",X"84",X"06",X"02",X"02",X"84",X"02",X"02",X"02",X"08",X"06",
		X"02",X"02",X"84",X"02",X"02",X"02",X"08",X"0E",X"02",X"02",X"02",X"02",X"02",X"02",X"48",X"02",
		X"0C",X"20",X"53",X"1B",X"3B",X"22",X"8C",X"8D",X"BB",X"12",X"42",X"22",X"8A",X"14",X"42",X"24",
		X"FD",X"FF",X"60",X"4E",X"1E",X"26",X"FC",X"26",X"26",X"C0",X"79",X"53",X"EC",X"00",X"A4",X"00",
		X"22",X"C5",X"14",X"EC",X"EF",X"2F",X"82",X"CA",X"7B",X"14",X"26",X"9D",X"08",X"BE",X"42",X"AC",
		X"AC",X"02",X"7B",X"14",X"26",X"9D",X"08",X"BE",X"FD",X"E7",X"20",X"D1",X"53",X"8B",X"8D",X"9D",
		X"83",X"76",X"72",X"3C",X"B5",X"02",X"B8",X"BC",X"FF",X"B3",X"06",X"B5",X"06",X"B7",X"44",X"B9",
		X"B0",X"3C",X"B0",X"1C",X"90",X"0D",X"81",X"B0",X"B0",X"12",X"90",X"03",X"81",X"B9",X"00",X"2D",
		X"03",X"B8",X"B2",X"76",X"72",X"2D",X"FF",X"B3",X"38",X"3A",X"41",X"3E",X"41",X"32",X"36",X"38",
		X"87",X"81",X"83",X"81",X"83",X"B0",X"45",X"70",X"B9",X"04",X"3A",X"81",X"70",X"B0",X"70",X"3E",
		X"02",X"02",X"02",X"06",X"08",X"0E",X"8A",X"08",X"02",X"02",X"48",X"06",X"02",X"02",X"02",X"06",
		X"48",X"06",X"06",X"06",X"08",X"02",X"02",X"02",X"02",X"08",X"06",X"08",X"4E",X"44",X"06",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"46",X"0C",X"06",X"08",
		X"08",X"0A",X"06",X"46",X"06",X"06",X"06",X"08",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"04",X"DD",X"39",X"04",X"D9",X"F9",X"F9",X"F9",X"95",X"99",X"F9",X"D5",X"42",X"D9",X"F9",X"F9",
		X"F9",X"F9",X"D5",X"40",X"D9",X"F9",X"D5",X"04",X"95",X"95",X"77",X"04",X"DD",X"39",X"04",X"3F",
		X"71",X"71",X"75",X"04",X"D9",X"F9",X"D5",X"04",X"39",X"42",X"DD",X"B7",X"73",X"73",X"77",X"04",
		X"75",X"04",X"3D",X"71",X"B9",X"B5",X"71",X"75",X"0A",X"D9",X"F9",X"D5",X"04",X"3D",X"71",X"75",
		X"5B",X"EB",X"89",X"FB",X"22",X"00",X"00",X"FB",X"53",X"E6",X"45",X"2E",X"4B",X"C0",X"81",X"79",
		X"44",X"1E",X"E4",X"4C",X"5C",X"E1",X"13",X"15",X"4D",X"42",X"83",X"F3",X"87",X"E4",X"86",X"5C",
		X"89",X"9F",X"33",X"0F",X"5E",X"0C",X"00",X"42",X"B5",X"9D",X"89",X"1D",X"4A",X"C0",X"3F",X"00",
		X"06",X"06",X"06",X"06",X"22",X"C8",X"8B",X"5B",X"26",X"1C",X"26",X"C4",X"04",X"86",X"EC",X"06",
		X"0E",X"FD",X"80",X"EC",X"02",X"15",X"33",X"28",X"5E",X"0C",X"00",X"22",X"6D",X"8B",X"42",X"FC",
		X"2B",X"8B",X"1D",X"8A",X"C0",X"75",X"CA",X"CA",X"0E",X"0E",X"0E",X"C0",X"C0",X"C0",X"C0",X"CA",
		X"B5",X"A8",X"2A",X"22",X"DF",X"8B",X"5B",X"EB",X"A8",X"2A",X"9F",X"57",X"BD",X"C0",X"BB",X"EA",
		X"8D",X"FD",X"46",X"59",X"BD",X"8B",X"FD",X"0C",X"5B",X"14",X"8D",X"33",X"13",X"E4",X"01",X"90",
		X"97",X"7D",X"04",X"DD",X"39",X"04",X"3D",X"71",X"F9",X"D5",X"04",X"DD",X"B7",X"73",X"73",X"73",
		X"F9",X"D5",X"04",X"3F",X"77",X"04",X"3F",X"73",X"F9",X"D5",X"04",X"DD",X"39",X"42",X"B1",X"F9",
		X"F9",X"D5",X"04",X"DD",X"39",X"04",X"3D",X"71",X"F9",X"D5",X"04",X"3D",X"71",X"71",X"71",X"75",
		X"00",X"00",X"00",X"00",X"34",X"02",X"04",X"02",X"02",X"08",X"0E",X"4E",X"0C",X"08",X"0E",X"02",
		X"4E",X"06",X"0C",X"08",X"08",X"4E",X"06",X"0C",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"06",
		X"0E",X"0A",X"06",X"06",X"08",X"02",X"02",X"02",X"02",X"08",X"0E",X"02",X"02",X"02",X"0E",X"02",
		X"0C",X"08",X"02",X"04",X"02",X"02",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7D",X"38",X"10",X"F8",X"10",X"09",X"16",
		X"8F",X"99",X"E6",X"B4",X"8F",X"8D",X"8F",X"8D",X"04",X"B7",X"44",X"B9",X"00",X"12",X"16",X"1A",
		X"41",X"47",X"74",X"76",X"B2",X"74",X"76",X"B2",X"B5",X"06",X"B7",X"44",X"B9",X"04",X"90",X"B0",
		X"76",X"70",X"74",X"70",X"3C",X"74",X"70",X"3C",X"B5",X"04",X"B7",X"44",X"B9",X"00",X"72",X"76",
		X"3C",X"38",X"32",X"72",X"76",X"72",X"0D",X"32",X"BC",X"A0",X"90",X"AA",X"BC",X"A0",X"90",X"98",
		X"3C",X"81",X"36",X"81",X"0D",X"81",X"0B",X"81",X"00",X"5E",X"FD",X"00",X"60",X"46",X"82",X"04",
		X"A1",X"E4",X"42",X"5C",X"22",X"B4",X"5C",X"2D",X"0A",X"EC",X"FF",X"A4",X"44",X"58",X"22",X"0B",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"16",X"5E",X"5A",X"90",X"9A",X"98",X"1A",X"94",
		X"12",X"98",X"52",X"5E",X"5C",X"20",X"20",X"20",X"32",X"76",X"32",X"7A",X"BA",X"B4",X"32",X"22",
		X"05",X"47",X"B6",X"4D",X"14",X"83",X"E8",X"89",X"EC",X"00",X"A4",X"4A",X"58",X"17",X"00",X"80",
		X"06",X"FD",X"0C",X"A0",X"C0",X"FA",X"87",X"1D",X"4A",X"58",X"B3",X"1D",X"04",X"A4",X"48",X"58",
		X"C2",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",
		X"00",X"00",X"00",X"FF",X"FD",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"95",X"77",X"04",X"3F",X"95",X"95",X"95",X"95",X"77",X"04",X"3D",X"71",X"71",X"71",X"75",X"04",
		X"11",X"11",X"11",X"39",X"04",X"D9",X"F9",X"D5",X"71",X"75",X"04",X"3D",X"71",X"71",X"71",X"75",
		X"11",X"11",X"11",X"39",X"04",X"D9",X"F9",X"D5",X"BB",X"39",X"04",X"DD",X"B7",X"73",X"73",X"77",
		X"73",X"73",X"73",X"77",X"04",X"D9",X"F9",X"D5",X"39",X"04",X"DD",X"39",X"40",X"D9",X"F9",X"F5",
		X"75",X"04",X"D9",X"F9",X"D5",X"04",X"DD",X"39",X"39",X"04",X"DD",X"39",X"48",X"DD",X"39",X"04",
		X"39",X"0A",X"DD",X"39",X"04",X"DD",X"B5",X"71",X"71",X"71",X"B9",X"39",X"04",X"D9",X"F9",X"D5",
		X"75",X"04",X"3F",X"77",X"04",X"3F",X"73",X"73",X"73",X"73",X"73",X"77",X"04",X"D9",X"F9",X"D5",
		X"39",X"40",X"D9",X"F9",X"F5",X"71",X"71",X"75",X"71",X"71",X"75",X"04",X"3D",X"71",X"71",X"75",
		X"39",X"0A",X"D9",X"F9",X"D5",X"04",X"DD",X"B5",X"5D",X"F9",X"F9",X"F9",X"D5",X"04",X"DD",X"11",
		X"75",X"04",X"D9",X"00",X"00",X"00",X"00",X"3C",X"02",X"46",X"02",X"02",X"0E",X"0C",X"06",X"06",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"06",X"0C",X"0E",X"06",X"06",X"06",X"0E",X"06",
		X"02",X"02",X"02",X"02",X"02",X"02",X"06",X"02",X"0C",X"06",X"0E",X"06",X"4A",X"0C",X"06",X"08",
		X"DD",X"39",X"04",X"D9",X"F9",X"D5",X"04",X"DD",X"F9",X"D5",X"0A",X"DD",X"39",X"0A",X"DD",X"39",
		X"3D",X"71",X"71",X"71",X"B9",X"39",X"04",X"5D",X"B9",X"39",X"04",X"3D",X"71",X"71",X"B9",X"39",
		X"02",X"02",X"04",X"02",X"08",X"06",X"86",X"0C",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"80",X"06",X"0C",X"08",X"06",X"80",X"06",X"0C",X"48",X"06",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"86",X"02",X"02",X"02",X"04",X"02",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E2",X"10",X"20",X"10",X"E6",X"36",X"10",X"F8",
		X"42",X"8E",X"42",X"4C",X"31",X"31",X"31",X"62",X"47",X"86",X"89",X"48",X"70",X"47",X"24",X"89",
		X"C8",X"58",X"48",X"01",X"65",X"65",X"EF",X"65",X"9A",X"75",X"FF",X"9E",X"9A",X"BB",X"9E",X"FF",
		X"02",X"02",X"02",X"06",X"0E",X"0C",X"06",X"06",X"06",X"02",X"02",X"02",X"46",X"02",X"02",X"B9",
		X"3A",X"10",X"F6",X"10",X"0B",X"16",X"C7",X"16",X"20",X"20",X"DD",X"31",X"24",X"20",X"20",X"20",
		X"98",X"4D",X"86",X"19",X"48",X"D2",X"4D",X"CC",X"4D",X"CA",X"88",X"48",X"04",X"65",X"65",X"01",
		X"0A",X"75",X"FF",X"9E",X"9A",X"BB",X"FF",X"9E",X"6F",X"65",X"04",X"0F",X"4D",X"84",X"00",X"00",
		X"BB",X"39",X"04",X"3F",X"73",X"73",X"BB",X"39",X"F9",X"D5",X"04",X"DD",X"39",X"42",X"DD",X"39",
		X"39",X"04",X"DD",X"39",X"04",X"D9",X"F9",X"D5",X"71",X"75",X"04",X"3F",X"77",X"04",X"3D",X"75",
		X"77",X"04",X"3F",X"77",X"04",X"D9",X"F9",X"D5",X"BB",X"39",X"0A",X"DD",X"39",X"4C",X"D9",X"F9",
		X"3D",X"71",X"71",X"B9",X"39",X"04",X"3D",X"71",X"71",X"71",X"B9",X"F9",X"D5",X"04",X"3F",X"77",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"02",X"00",
		X"02",X"00",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",
		X"FF",X"10",X"F9",X"91",X"95",X"95",X"95",X"95",X"F9",X"F9",X"F9",X"D5",X"04",X"D9",X"F9",X"F9",
		X"95",X"99",X"F9",X"D5",X"0A",X"D9",X"F9",X"D5",X"D5",X"04",X"D9",X"F9",X"F9",X"F9",X"D5",X"40",
		X"DD",X"39",X"04",X"DD",X"39",X"04",X"3D",X"71",X"71",X"71",X"71",X"75",X"04",X"D9",X"F9",X"F7",
		X"3F",X"77",X"04",X"3F",X"77",X"04",X"3F",X"73",X"B7",X"73",X"73",X"77",X"04",X"D9",X"F9",X"D5",
		X"DD",X"39",X"0A",X"D9",X"F9",X"D5",X"04",X"3D",X"04",X"79",X"97",X"97",X"97",X"7D",X"04",X"DD",
		X"3D",X"75",X"04",X"D9",X"F9",X"D5",X"04",X"DD",X"04",X"D9",X"F9",X"F9",X"F9",X"D5",X"04",X"3F",
		X"75",X"04",X"D9",X"F9",X"F7",X"73",X"73",X"77",X"73",X"73",X"77",X"04",X"3F",X"73",X"BB",X"39",
		X"39",X"04",X"D9",X"F9",X"D5",X"84",X"DD",X"39",X"F9",X"D5",X"04",X"3D",X"75",X"04",X"3D",X"71",
		X"97",X"7D",X"04",X"3F",X"77",X"04",X"3F",X"77",X"F9",X"D5",X"04",X"DD",X"39",X"04",X"3F",X"73",
		X"F9",X"D5",X"40",X"DD",X"39",X"04",X"3F",X"77",X"DD",X"39",X"04",X"B1",X"F9",X"F9",X"F9",X"D5",
		X"02",X"02",X"02",X"06",X"08",X"06",X"80",X"06",X"06",X"06",X"08",X"06",X"02",X"02",X"02",X"02",
		X"0E",X"8A",X"08",X"06",X"02",X"02",X"02",X"02",X"02",X"02",X"06",X"06",X"08",X"06",X"80",X"06",
		X"02",X"4A",X"06",X"02",X"02",X"02",X"06",X"0E",X"06",X"0E",X"06",X"06",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"0E",X"06",X"06",X"02",X"06",X"0E",X"06",X"0C",X"0E",X"0C",X"06",
		X"06",X"0C",X"08",X"02",X"02",X"02",X"08",X"48",X"06",X"08",X"4E",X"06",X"06",X"08",X"06",X"08",
		X"02",X"4E",X"02",X"02",X"02",X"06",X"08",X"06",X"02",X"02",X"4E",X"02",X"02",X"02",X"06",X"08",
		X"4E",X"06",X"06",X"08",X"02",X"02",X"02",X"08",X"0E",X"08",X"48",X"06",X"0C",X"0E",X"08",X"48",
		X"02",X"02",X"48",X"06",X"02",X"02",X"02",X"02",X"06",X"80",X"06",X"0C",X"08",X"06",X"02",X"02",
		X"FF",X"65",X"89",X"47",X"88",X"00",X"00",X"C3",X"00",X"2D",X"47",X"CA",X"9A",X"10",X"9A",X"9A",
		X"01",X"65",X"04",X"01",X"65",X"65",X"9A",X"00",X"D5",X"04",X"DD",X"D1",X"95",X"95",X"95",X"95",
		X"95",X"99",X"F9",X"F9",X"F9",X"F9",X"D5",X"04",X"D5",X"04",X"DD",X"39",X"40",X"DD",X"39",X"0A",
		X"39",X"0A",X"D9",X"F9",X"D5",X"04",X"DD",X"39",X"39",X"04",X"3D",X"75",X"04",X"3F",X"95",X"95",
		X"00",X"00",X"CB",X"4D",X"68",X"00",X"00",X"9A",X"21",X"75",X"FF",X"FF",X"65",X"64",X"21",X"04",
		X"64",X"00",X"98",X"0A",X"00",X"00",X"9A",X"FB",X"95",X"9D",X"39",X"04",X"3F",X"95",X"95",X"95",
		X"D1",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"39",X"40",X"D9",X"F9",X"D5",X"04",X"3D",X"71",
		X"71",X"75",X"04",X"3D",X"71",X"71",X"71",X"75",X"75",X"04",X"D9",X"F9",X"D5",X"04",X"DD",X"B7",
		X"3F",X"73",X"73",X"73",X"77",X"04",X"DD",X"B7",X"73",X"73",X"BB",X"F9",X"D5",X"0A",X"DD",X"11",
		X"D9",X"F9",X"F5",X"71",X"71",X"75",X"04",X"DD",X"97",X"97",X"7D",X"04",X"DD",X"39",X"04",X"3D",
		X"D9",X"F9",X"F7",X"73",X"73",X"77",X"04",X"3F",X"F9",X"F9",X"D5",X"04",X"3F",X"77",X"04",X"DD",
		X"D9",X"F9",X"D5",X"42",X"DD",X"39",X"04",X"B1",X"DD",X"39",X"04",X"D9",X"F9",X"D5",X"04",X"3D",
		X"F5",X"FF",X"9A",X"9A",X"02",X"01",X"65",X"04",X"BB",X"7B",X"D6",X"95",X"5A",X"F8",X"85",X"1D",
		X"06",X"FD",X"0C",X"A0",X"80",X"EC",X"02",X"A4",X"9D",X"04",X"17",X"A5",X"C2",X"B3",X"17",X"5B",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"02",
		X"FF",X"00",X"00",X"FF",X"FD",X"00",X"00",X"00",X"FF",X"00",X"00",X"02",X"FF",X"02",X"FF",X"00",
		X"95",X"95",X"77",X"04",X"3F",X"95",X"95",X"95",X"D9",X"F9",X"D5",X"04",X"DD",X"39",X"8A",X"DD",
		X"04",X"DD",X"39",X"04",X"3D",X"71",X"71",X"71",X"04",X"3D",X"75",X"04",X"3D",X"75",X"04",X"DD",
		X"04",X"3F",X"77",X"04",X"3F",X"73",X"73",X"73",X"04",X"DD",X"39",X"04",X"DD",X"39",X"04",X"3F",
		X"42",X"DD",X"39",X"04",X"DD",X"39",X"0A",X"DD",X"71",X"71",X"75",X"04",X"3D",X"71",X"75",X"04",
		X"04",X"DD",X"B7",X"73",X"73",X"77",X"04",X"DD",X"D9",X"F9",X"D5",X"04",X"DD",X"39",X"04",X"DD",
		X"71",X"71",X"75",X"04",X"3D",X"75",X"04",X"3D",X"04",X"3F",X"77",X"04",X"DD",X"39",X"04",X"3D",
		X"73",X"73",X"77",X"04",X"DD",X"39",X"04",X"3F",X"0A",X"DD",X"39",X"04",X"DD",X"39",X"48",X"DD",
		X"04",X"DD",X"39",X"04",X"DD",X"B5",X"71",X"71",X"04",X"DD",X"B5",X"71",X"71",X"75",X"04",X"3D",
		X"71",X"71",X"71",X"75",X"04",X"DD",X"39",X"04",X"11",X"11",X"39",X"04",X"DD",X"B5",X"71",X"71",
		X"02",X"02",X"02",X"02",X"02",X"06",X"02",X"02",X"44",X"06",X"0E",X"0C",X"06",X"06",X"02",X"02",
		X"06",X"0E",X"06",X"02",X"02",X"02",X"06",X"0E",X"0C",X"0E",X"06",X"06",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"0E",X"06",X"4A",X"02",X"02",X"02",X"02",X"02",X"02",X"4A",X"06",
		X"39",X"0C",X"DD",X"39",X"04",X"B1",X"F9",X"F9",X"04",X"D9",X"F9",X"D5",X"04",X"DD",X"39",X"04",
		X"F9",X"F9",X"F9",X"D5",X"04",X"3D",X"71",X"71",X"04",X"D9",X"00",X"34",X"04",X"02",X"86",X"02",
		X"08",X"06",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"0C",X"08",X"06",
		X"08",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"0E",X"08",X"48",X"06",X"0C",X"0E",X"08",X"48",
		X"02",X"0C",X"08",X"06",X"86",X"0C",X"08",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"31",X"CA",X"24",X"CA",X"10",X"07",X"16",X"C9",X"16",X"52",X"42",X"8E",
		X"42",X"8E",X"42",X"8E",X"42",X"00",X"00",X"36",X"B9",X"B2",X"47",X"2E",X"58",X"B9",X"F6",X"47",
		X"01",X"44",X"98",X"9A",X"9A",X"9A",X"FF",X"DE",X"8A",X"10",X"9A",X"75",X"6F",X"04",X"75",X"FF",
		X"44",X"06",X"40",X"02",X"02",X"02",X"02",X"02",X"CA",X"24",X"CA",X"E2",X"10",X"20",X"10",X"E6",
		X"14",X"8C",X"44",X"8C",X"44",X"8C",X"44",X"20",X"20",X"8C",X"44",X"8C",X"44",X"8C",X"00",X"00",
		X"19",X"B9",X"32",X"4D",X"2C",X"88",X"B9",X"76",X"64",X"04",X"10",X"9A",X"FE",X"9A",X"8A",X"90",
		X"FE",X"9A",X"0A",X"75",X"FF",X"FF",X"FF",X"75",X"49",X"4D",X"CA",X"00",X"00",X"89",X"4D",X"22",
		X"0A",X"DD",X"39",X"04",X"DD",X"39",X"04",X"D9",X"0A",X"DD",X"39",X"04",X"3D",X"71",X"71",X"B9",
		X"04",X"DD",X"39",X"04",X"3D",X"71",X"71",X"71",X"04",X"3F",X"77",X"04",X"3F",X"73",X"73",X"73",
		X"04",X"DD",X"39",X"04",X"3F",X"73",X"73",X"73",X"D5",X"04",X"DD",X"39",X"0C",X"DD",X"39",X"04",
		X"71",X"71",X"75",X"04",X"3D",X"71",X"71",X"71",X"04",X"3D",X"71",X"75",X"04",X"3F",X"77",X"04",
		X"00",X"00",X"02",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"02",X"02",X"02",
		X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",
		X"99",X"F9",X"D5",X"04",X"D9",X"F9",X"F9",X"F9",X"F9",X"91",X"95",X"95",X"95",X"95",X"95",X"95",
		X"04",X"D9",X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",X"D9",X"F9",X"D5",X"04",X"3D",X"75",X"04",X"3F",
		X"71",X"B9",X"39",X"04",X"DD",X"39",X"04",X"3D",X"73",X"73",X"77",X"04",X"DD",X"11",X"39",X"04",
		X"73",X"BB",X"39",X"04",X"3F",X"77",X"04",X"DD",X"0A",X"DD",X"11",X"39",X"46",X"DD",X"39",X"0A",
		X"75",X"04",X"DD",X"11",X"39",X"04",X"3D",X"75",X"39",X"04",X"3D",X"75",X"04",X"DD",X"39",X"04",
		X"39",X"04",X"3F",X"73",X"77",X"04",X"DD",X"39",X"77",X"04",X"DD",X"39",X"04",X"3F",X"77",X"04",
		X"04",X"3F",X"77",X"04",X"3F",X"73",X"73",X"73",X"04",X"DD",X"B7",X"73",X"73",X"77",X"04",X"DD",
		X"04",X"DD",X"39",X"0A",X"DD",X"39",X"04",X"D9",X"71",X"71",X"71",X"75",X"04",X"79",X"97",X"97",
		X"04",X"3D",X"75",X"04",X"DD",X"39",X"04",X"D9",X"73",X"73",X"BB",X"39",X"04",X"D9",X"F9",X"F9",
		X"04",X"D9",X"F9",X"D5",X"04",X"DD",X"39",X"0C",X"04",X"3D",X"71",X"71",X"71",X"75",X"04",X"DD",
		X"06",X"06",X"08",X"06",X"80",X"02",X"02",X"02",X"84",X"02",X"02",X"02",X"08",X"0E",X"8A",X"08",
		X"84",X"02",X"02",X"02",X"08",X"06",X"80",X"02",X"06",X"06",X"08",X"02",X"02",X"02",X"02",X"02",
		X"06",X"4A",X"0C",X"06",X"0E",X"06",X"4A",X"0C",X"02",X"02",X"02",X"02",X"02",X"02",X"06",X"02",
		X"06",X"0E",X"06",X"0C",X"0E",X"06",X"02",X"02",X"06",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"06",X"02",X"02",X"02",X"08",X"4E",X"06",X"06",X"08",X"06",X"02",X"02",X"02",
		X"C2",X"08",X"06",X"C2",X"08",X"06",X"02",X"02",X"06",X"08",X"4E",X"06",X"06",X"08",X"06",X"08",
		X"48",X"02",X"02",X"02",X"06",X"02",X"02",X"02",X"06",X"0C",X"08",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"08",X"06",X"80",X"06",X"0C",X"08",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"47",X"8E",X"00",X"00",X"CF",X"47",X"C4",X"00",X"EF",X"65",X"01",X"65",X"65",X"EF",X"65",X"65",
		X"00",X"00",X"9A",X"9A",X"FB",X"65",X"10",X"F9",X"95",X"95",X"95",X"9D",X"D1",X"95",X"95",X"95",
		X"DD",X"D1",X"95",X"95",X"95",X"95",X"99",X"F9",X"D9",X"F9",X"F9",X"F9",X"F9",X"D5",X"04",X"DD",
		X"04",X"3D",X"71",X"71",X"71",X"75",X"04",X"DD",X"95",X"95",X"77",X"04",X"3F",X"77",X"04",X"3D",
		X"FE",X"9A",X"9B",X"FF",X"65",X"EF",X"65",X"64",X"00",X"00",X"21",X"65",X"04",X"9A",X"8A",X"21",
		X"10",X"F9",X"91",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"9D",
		X"99",X"F9",X"D5",X"0E",X"DD",X"39",X"4A",X"DD",X"71",X"75",X"04",X"DD",X"39",X"04",X"3D",X"71",
		X"04",X"3F",X"77",X"04",X"3D",X"75",X"04",X"3D",X"73",X"77",X"04",X"3F",X"77",X"04",X"3F",X"73",
		X"73",X"73",X"77",X"04",X"DD",X"B7",X"73",X"73",X"39",X"46",X"DD",X"39",X"0A",X"DD",X"39",X"0A",
		X"11",X"39",X"04",X"3D",X"75",X"04",X"79",X"97",X"75",X"04",X"DD",X"39",X"04",X"3D",X"75",X"04",
		X"73",X"77",X"04",X"DD",X"39",X"04",X"D9",X"F9",X"39",X"04",X"3F",X"77",X"04",X"DD",X"39",X"04",
		X"F9",X"F9",X"F9",X"D5",X"0A",X"DD",X"39",X"0A",X"71",X"71",X"71",X"71",X"75",X"04",X"DD",X"39",
		X"22",X"00",X"00",X"02",X"00",X"80",X"A4",X"11",X"FD",X"04",X"95",X"42",X"A0",X"28",X"80",X"7D",
		X"FD",X"A0",X"15",X"06",X"A0",X"2C",X"00",X"68",X"A0",X"2A",X"F8",X"3D",X"B1",X"A4",X"0E",X"90",
		X"EB",X"A0",X"A2",X"98",X"A2",X"0C",X"FF",X"33",X"1D",X"A6",X"5E",X"68",X"FA",X"3D",X"4E",X"15",
		X"5E",X"FA",X"2F",X"15",X"5A",X"A0",X"28",X"8A",X"93",X"50",X"A4",X"11",X"90",X"F2",X"27",X"5E",
		X"12",X"1B",X"3B",X"0C",X"28",X"5B",X"DC",X"68",X"82",X"FD",X"58",X"64",X"7C",X"A2",X"A0",X"44",
		X"B4",X"A2",X"FA",X"A4",X"08",X"14",X"F8",X"A4",X"90",X"A1",X"3D",X"02",X"20",X"82",X"13",X"F2",
		X"4E",X"4E",X"5E",X"7B",X"16",X"0B",X"12",X"A4",X"BD",X"17",X"46",X"26",X"00",X"58",X"4E",X"08",
		X"00",X"10",X"B1",X"08",X"00",X"18",X"4E",X"08",X"12",X"9C",X"12",X"16",X"22",X"0C",X"90",X"EC",
		X"0A",X"40",X"0E",X"E1",X"46",X"39",X"48",X"FD",X"74",X"9B",X"74",X"AD",X"7A",X"7A",X"D7",X"7A",
		X"28",X"24",X"83",X"85",X"28",X"85",X"28",X"68",X"48",X"FD",X"FF",X"FF",X"FF",X"E4",X"00",X"5E",
		X"EC",X"02",X"A4",X"69",X"14",X"EC",X"8C",X"A4",X"00",X"5E",X"FD",X"02",X"55",X"C9",X"A8",X"7F",
		X"8C",X"A4",X"69",X"1C",X"4C",X"48",X"17",X"C9",X"A8",X"7F",X"C8",X"8A",X"EC",X"06",X"A4",X"69",
		X"5B",X"9C",X"AA",X"C6",X"84",X"5B",X"12",X"AC",X"F0",X"9F",X"3B",X"E8",X"5E",X"22",X"EC",X"5E",
		X"2C",X"AA",X"4C",X"00",X"C0",X"7F",X"33",X"B2",X"5C",X"5E",X"DF",X"33",X"77",X"B4",X"66",X"E4",
		X"08",X"EC",X"11",X"67",X"DE",X"B6",X"22",X"8E",X"20",X"34",X"CC",X"08",X"C0",X"DC",X"5E",X"57",
		X"B5",X"70",X"AA",X"BD",X"B1",X"48",X"C0",X"04",X"9B",X"26",X"9C",X"26",X"DC",X"C0",X"86",X"77",
		X"DE",X"9B",X"0C",X"66",X"5B",X"DC",X"68",X"0C",X"F3",X"A4",X"C2",X"FC",X"A4",X"64",X"14",X"26",
		X"4E",X"3D",X"06",X"1D",X"A2",X"FD",X"A8",X"20",X"DC",X"68",X"E4",X"10",X"90",X"0E",X"3D",X"02",
		X"90",X"3D",X"80",X"55",X"41",X"A2",X"6F",X"A4",X"6A",X"20",X"F9",X"A2",X"35",X"E4",X"0C",X"06",
		X"E8",X"BE",X"26",X"B4",X"26",X"80",X"F1",X"E6",X"80",X"F1",X"E6",X"E6",X"CA",X"15",X"D6",X"A4",
		X"FF",X"02",X"00",X"00",X"02",X"FF",X"00",X"00",X"64",X"9A",X"64",X"9A",X"9A",X"9A",X"9A",X"9A",
		X"2A",X"2A",X"2A",X"24",X"24",X"24",X"24",X"02",X"42",X"80",X"4C",X"70",X"80",X"B0",X"8E",X"88",
		X"9A",X"9A",X"64",X"9A",X"64",X"94",X"54",X"2B",X"83",X"02",X"02",X"02",X"02",X"00",X"00",X"00",
		X"00",X"00",X"00",X"9A",X"64",X"9A",X"64",X"9A",X"64",X"9A",X"64",X"94",X"54",X"2B",X"89",X"50",
		X"69",X"14",X"82",X"02",X"00",X"C0",X"6B",X"26",X"27",X"E4",X"04",X"5C",X"2F",X"20",X"40",X"EC",
		X"B1",X"03",X"0C",X"00",X"42",X"82",X"04",X"5E",X"00",X"5E",X"A4",X"29",X"5A",X"22",X"CE",X"5E",
		X"53",X"F0",X"FD",X"0C",X"20",X"08",X"22",X"1D",X"F0",X"FD",X"02",X"60",X"08",X"0C",X"00",X"C0",
		X"60",X"40",X"0C",X"04",X"FD",X"08",X"60",X"04",X"BE",X"55",X"3C",X"20",X"EC",X"02",X"04",X"53",
		X"E2",X"55",X"E2",X"2B",X"EA",X"22",X"EC",X"1D",X"EA",X"A0",X"EC",X"99",X"07",X"50",X"52",X"1E",
		X"4F",X"6E",X"01",X"E6",X"01",X"16",X"94",X"1A",X"6E",X"01",X"E6",X"01",X"1C",X"94",X"1A",X"1A",
		X"01",X"49",X"04",X"90",X"58",X"12",X"D2",X"1A",X"80",X"80",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",
		X"1A",X"94",X"10",X"98",X"9E",X"5E",X"6E",X"0B",X"10",X"10",X"5E",X"9C",X"1A",X"94",X"6E",X"03",
		X"5E",X"68",X"FA",X"3D",X"4E",X"15",X"BA",X"A0",X"2F",X"15",X"BA",X"A0",X"28",X"8A",X"15",X"B4",
		X"1E",X"80",X"29",X"B3",X"93",X"FD",X"18",X"15",X"0C",X"02",X"17",X"EB",X"A0",X"F6",X"3D",X"02",
		X"D3",X"22",X"00",X"58",X"0C",X"08",X"A4",X"11",X"BB",X"22",X"00",X"10",X"0C",X"08",X"A4",X"11",
		X"80",X"B9",X"0C",X"08",X"A4",X"11",X"90",X"EC",X"D3",X"80",X"40",X"0C",X"26",X"5B",X"DC",X"68",
		X"90",X"9D",X"08",X"97",X"00",X"A2",X"11",X"5E",X"A4",X"02",X"5C",X"A4",X"00",X"90",X"F7",X"E4",
		X"EC",X"04",X"A4",X"C9",X"5C",X"E4",X"10",X"90",X"A4",X"C9",X"5C",X"F0",X"A3",X"3D",X"02",X"60",
		X"3D",X"04",X"60",X"0A",X"EC",X"08",X"A4",X"E9",X"80",X"A4",X"E9",X"5C",X"F0",X"A3",X"3D",X"40",
		X"01",X"90",X"3D",X"06",X"1D",X"2A",X"1E",X"5B",X"4E",X"3D",X"06",X"FD",X"06",X"20",X"40",X"0C",
		X"17",X"C9",X"A8",X"4C",X"28",X"17",X"C9",X"A8",X"C9",X"A8",X"4C",X"50",X"17",X"C9",X"A8",X"4C",
		X"59",X"82",X"AC",X"0C",X"0C",X"DB",X"22",X"48",X"FD",X"B1",X"55",X"DD",X"A8",X"FD",X"B3",X"55",
		X"B7",X"55",X"BE",X"AA",X"FD",X"BB",X"55",X"0E",X"55",X"B7",X"AA",X"FD",X"F1",X"55",X"FB",X"AA",
		X"02",X"9F",X"5E",X"22",X"6C",X"5E",X"DF",X"F2",X"DF",X"F8",X"03",X"84",X"33",X"3B",X"EC",X"04",
		X"82",X"EC",X"5E",X"9B",X"26",X"DC",X"26",X"9C",X"66",X"B6",X"82",X"06",X"00",X"C0",X"CA",X"26",
		X"04",X"00",X"C0",X"80",X"22",X"8E",X"5E",X"F0",X"CC",X"02",X"C0",X"00",X"DB",X"7C",X"00",X"DB",
		X"02",X"DB",X"66",X"DB",X"66",X"80",X"02",X"53",X"AC",X"02",X"22",X"20",X"5E",X"FC",X"26",X"2D",
		X"82",X"00",X"00",X"60",X"5F",X"E4",X"04",X"5C",X"17",X"4D",X"0A",X"F0",X"7F",X"C8",X"A0",X"1E",
		X"40",X"5B",X"7B",X"A4",X"80",X"F7",X"A4",X"11",X"E4",X"10",X"90",X"3D",X"30",X"15",X"56",X"26",
		X"10",X"90",X"3D",X"80",X"15",X"56",X"26",X"CC",X"A4",X"E4",X"00",X"90",X"27",X"20",X"B9",X"5B",
		X"7D",X"FF",X"20",X"B7",X"80",X"3B",X"57",X"06",X"10",X"0C",X"08",X"EC",X"10",X"BE",X"68",X"20",
		X"11",X"90",X"E4",X"10",X"90",X"3D",X"80",X"55",X"22",X"00",X"60",X"66",X"F8",X"AB",X"20",X"F7",
		X"04",X"A8",X"40",X"D1",X"42",X"A9",X"4E",X"D0",X"9A",X"9B",X"74",X"9B",X"74",X"65",X"74",X"9A",
		X"9A",X"85",X"28",X"85",X"28",X"24",X"24",X"24",X"48",X"99",X"4A",X"09",X"84",X"A1",X"86",X"9B",
		X"D4",X"6B",X"AB",X"9B",X"74",X"9B",X"74",X"65",X"28",X"24",X"83",X"29",X"02",X"98",X"0C",X"F1",
		X"FF",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"9D",X"D4",X"6B",X"AB",X"2A",X"2A",X"2A",
		X"40",X"5A",X"3D",X"4E",X"57",X"EE",X"57",X"EE",X"EC",X"AC",X"A4",X"44",X"58",X"53",X"06",X"08",
		X"02",X"08",X"02",X"02",X"02",X"86",X"AE",X"26",X"AE",X"F4",X"AE",X"0D",X"AE",X"CB",X"AE",X"A3",
		X"EA",X"37",X"EA",X"0D",X"EA",X"04",X"EC",X"58",X"EA",X"BC",X"EA",X"B5",X"EA",X"02",X"00",X"04",
		X"E0",X"D1",X"E0",X"35",X"E0",X"79",X"E0",X"BD",X"E2",X"64",X"E2",X"D0",X"E2",X"12",X"E2",X"82",
		X"D2",X"D6",X"6E",X"43",X"6E",X"81",X"7B",X"04",X"94",X"98",X"10",X"14",X"9A",X"98",X"98",X"5E",
		X"10",X"90",X"58",X"12",X"D2",X"1A",X"94",X"10",X"01",X"6F",X"04",X"A2",X"10",X"5E",X"94",X"10",
		X"96",X"6E",X"0F",X"00",X"6E",X"00",X"01",X"00",X"90",X"9A",X"16",X"56",X"5A",X"12",X"5C",X"10",
		X"A0",X"10",X"DA",X"DC",X"DE",X"6E",X"4D",X"6E",X"66",X"68",X"6A",X"6C",X"10",X"A2",X"E2",X"E0",
		X"90",X"F2",X"0D",X"5E",X"FA",X"1D",X"04",X"7E",X"F2",X"2F",X"20",X"8A",X"A4",X"0E",X"90",X"F8",
		X"FA",X"FD",X"04",X"D5",X"06",X"A0",X"17",X"14",X"4E",X"4E",X"4E",X"4E",X"DE",X"0C",X"00",X"17",
		X"93",X"50",X"A4",X"11",X"90",X"F2",X"27",X"BE",X"5A",X"A0",X"F2",X"0F",X"0F",X"03",X"1D",X"A2",
		X"15",X"54",X"A0",X"E6",X"E6",X"E6",X"E6",X"33",X"FC",X"27",X"E3",X"15",X"AB",X"A0",X"1D",X"A6",
		X"33",X"F8",X"FD",X"10",X"64",X"78",X"A2",X"E0",X"FD",X"18",X"64",X"B0",X"A2",X"E0",X"06",X"64",
		X"38",X"14",X"E4",X"00",X"90",X"1E",X"E4",X"10",X"3D",X"4E",X"1E",X"F2",X"3D",X"B1",X"4E",X"4E",
		X"11",X"90",X"E4",X"10",X"90",X"3D",X"80",X"60",X"00",X"58",X"B1",X"08",X"00",X"10",X"4E",X"08",
		X"00",X"18",X"B1",X"08",X"5E",X"10",X"12",X"9E",X"02",X"BE",X"6A",X"20",X"F9",X"6F",X"A4",X"06",
		X"FF",X"FF",X"FF",X"9B",X"74",X"9B",X"74",X"9B",X"7A",X"7A",X"7A",X"9D",X"D4",X"6B",X"AB",X"50",
		X"02",X"D9",X"0A",X"40",X"0E",X"E1",X"46",X"39",X"FD",X"02",X"55",X"C9",X"A8",X"7F",X"C8",X"A4",
		X"69",X"1C",X"4C",X"00",X"17",X"C9",X"A8",X"E4",X"C8",X"8E",X"EC",X"04",X"A4",X"69",X"14",X"EC",
		X"A8",X"E4",X"00",X"5E",X"FD",X"02",X"55",X"C9",X"14",X"EC",X"8C",X"A4",X"69",X"1C",X"4C",X"C0",
		X"DF",X"FA",X"03",X"C6",X"84",X"22",X"4E",X"5E",X"DF",X"F2",X"57",X"6E",X"9F",X"FD",X"FF",X"15",
		X"DE",X"33",X"EC",X"06",X"9F",X"9E",X"9B",X"22",X"42",X"5C",X"5E",X"E4",X"B4",X"5C",X"23",X"60",
		X"5E",X"F0",X"9F",X"EA",X"BE",X"82",X"00",X"00",X"62",X"57",X"62",X"57",X"62",X"57",X"62",X"2F",
		X"3D",X"4E",X"53",X"77",X"5B",X"12",X"AC",X"77",X"22",X"4E",X"5E",X"F0",X"9F",X"AC",X"00",X"77",
		X"6C",X"5B",X"DC",X"68",X"93",X"8C",X"00",X"22",X"FC",X"A4",X"54",X"14",X"E4",X"01",X"90",X"4E",
		X"02",X"E8",X"A4",X"69",X"12",X"0C",X"62",X"5B",X"1D",X"68",X"1E",X"5B",X"DC",X"68",X"E4",X"10",
		X"00",X"90",X"B7",X"22",X"0E",X"90",X"6F",X"BE",X"D3",X"33",X"93",X"A4",X"11",X"90",X"13",X"EC",
		X"E6",X"13",X"B2",X"26",X"EC",X"EE",X"BE",X"26",X"B3",X"D3",X"80",X"D9",X"A2",X"11",X"5E",X"0C",
		X"FF",X"02",X"00",X"00",X"02",X"FF",X"00",X"9A",X"64",X"9A",X"64",X"94",X"54",X"2B",X"89",X"2A",
		X"02",X"02",X"02",X"D0",X"04",X"40",X"0E",X"30",X"C2",X"94",X"54",X"2B",X"89",X"65",X"64",X"9A",
		X"89",X"85",X"28",X"2A",X"52",X"50",X"28",X"24",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"9A",X"9A",X"9A",X"65",X"64",X"9A",X"9A",X"9A",X"28",X"24",X"83",X"22",X"18",X"18",X"40",X"D0",
		X"FC",X"A4",X"E9",X"5C",X"82",X"04",X"00",X"C0",X"04",X"A4",X"59",X"5C",X"A4",X"D9",X"5C",X"22",
		X"02",X"48",X"00",X"7B",X"A1",X"EC",X"02",X"A4",X"EC",X"00",X"A4",X"2B",X"5A",X"0C",X"88",X"5F",
		X"5A",X"53",X"22",X"FD",X"58",X"53",X"0A",X"1B",X"82",X"E4",X"86",X"5C",X"0C",X"02",X"FD",X"02",
		X"0C",X"06",X"DF",X"13",X"17",X"B4",X"6A",X"57",X"22",X"00",X"00",X"24",X"95",X"5A",X"53",X"E4",
		X"EA",X"10",X"EC",X"8B",X"EA",X"82",X"EC",X"A9",X"50",X"10",X"96",X"16",X"5E",X"94",X"1A",X"6E",
		X"18",X"52",X"98",X"10",X"10",X"10",X"6E",X"4F",X"10",X"90",X"58",X"12",X"D2",X"6E",X"4F",X"6E",
		X"94",X"10",X"5E",X"5C",X"1A",X"6E",X"0B",X"6E",X"80",X"80",X"49",X"04",X"90",X"58",X"12",X"D2",
		X"6E",X"01",X"85",X"04",X"1E",X"12",X"5A",X"1A",X"6E",X"01",X"94",X"04",X"94",X"1A",X"12",X"18",
		X"F2",X"0F",X"0F",X"03",X"1D",X"A2",X"5E",X"FA",X"A0",X"E6",X"E6",X"E6",X"E6",X"F0",X"9D",X"80",
		X"1A",X"A0",X"F6",X"7D",X"B1",X"15",X"1A",X"A0",X"7D",X"02",X"DE",X"0C",X"00",X"A2",X"11",X"5E",
		X"90",X"AC",X"00",X"68",X"20",X"F7",X"28",X"80",X"90",X"EC",X"10",X"BE",X"68",X"20",X"F9",X"28",
		X"4E",X"BE",X"68",X"20",X"F9",X"28",X"80",X"B9",X"17",X"B8",X"A2",X"F6",X"1D",X"A0",X"A4",X"09",
		X"A4",X"11",X"90",X"6F",X"A4",X"00",X"5C",X"E8",X"00",X"90",X"6E",X"1E",X"3D",X"31",X"60",X"0A",
		X"6E",X"5E",X"3D",X"30",X"60",X"0A",X"EC",X"02",X"0A",X"EC",X"40",X"A4",X"E9",X"5C",X"F0",X"A3",
		X"5C",X"F0",X"A3",X"3D",X"08",X"60",X"0A",X"EC",X"60",X"0A",X"EC",X"20",X"A4",X"E9",X"5C",X"E4",
		X"DC",X"68",X"E4",X"01",X"90",X"4E",X"4E",X"4E",X"64",X"5B",X"DC",X"68",X"17",X"C8",X"A4",X"0E",
		X"4C",X"A0",X"17",X"C9",X"A8",X"4C",X"E8",X"17",X"98",X"17",X"C9",X"A8",X"E4",X"00",X"5E",X"2F",
		X"5E",X"DB",X"7C",X"00",X"DB",X"3C",X"02",X"FC",X"76",X"AA",X"FD",X"B5",X"55",X"8F",X"AA",X"FD",
		X"AC",X"FD",X"BD",X"55",X"29",X"AA",X"FD",X"BF",X"FD",X"FF",X"55",X"57",X"AA",X"BC",X"3B",X"EC",
		X"09",X"5B",X"9C",X"AA",X"84",X"5B",X"12",X"AC",X"9F",X"5E",X"22",X"6C",X"5E",X"DF",X"F2",X"0B",
		X"C0",X"00",X"33",X"9B",X"DF",X"77",X"93",X"B4",X"5C",X"22",X"8E",X"5E",X"F0",X"9F",X"B2",X"82",
		X"9F",X"EA",X"BE",X"82",X"00",X"00",X"20",X"08",X"3C",X"02",X"C2",X"DB",X"BA",X"00",X"DB",X"B8",
		X"17",X"63",X"A8",X"22",X"CE",X"5E",X"F0",X"9F",X"26",X"2D",X"26",X"2D",X"26",X"2D",X"26",X"2D",
		X"2F",X"55",X"8B",X"22",X"6F",X"A4",X"00",X"5E",X"82",X"02",X"00",X"C0",X"AF",X"EC",X"10",X"A4",
		X"90",X"E4",X"10",X"90",X"3D",X"80",X"60",X"BD",X"0C",X"40",X"5B",X"7B",X"A4",X"80",X"F7",X"E4",
		X"02",X"0C",X"08",X"A4",X"11",X"90",X"5B",X"7B",X"7B",X"A4",X"A4",X"11",X"90",X"E4",X"00",X"90",
		X"F6",X"FD",X"80",X"D5",X"63",X"A4",X"22",X"00",X"F9",X"28",X"80",X"BF",X"5B",X"B9",X"E4",X"A4",
		X"DF",X"A4",X"17",X"56",X"26",X"A4",X"11",X"90",X"53",X"A0",X"A2",X"AA",X"A2",X"A0",X"A4",X"00",
		X"82",X"40",X"8C",X"A8",X"8E",X"9A",X"9A",X"9A",X"9B",X"9A",X"9A",X"9A",X"9A",X"65",X"64",X"9A",
		X"24",X"29",X"02",X"98",X"0C",X"F1",X"0E",X"61",X"74",X"9B",X"74",X"9D",X"D4",X"6B",X"AB",X"9D",
		X"74",X"9A",X"9B",X"85",X"28",X"2A",X"52",X"50",X"0E",X"61",X"48",X"99",X"4A",X"FD",X"FF",X"FF",
		X"7A",X"AD",X"7A",X"7A",X"D7",X"7A",X"7A",X"7A",X"2A",X"85",X"28",X"85",X"28",X"68",X"02",X"D9",
		X"6E",X"CC",X"C8",X"07",X"FD",X"C0",X"20",X"04",X"02",X"04",X"02",X"02",X"02",X"02",X"48",X"02",
		X"AE",X"A4",X"AE",X"12",X"AE",X"D4",X"AE",X"74",X"AE",X"22",X"EA",X"00",X"EA",X"FB",X"AE",X"3E",
		X"E0",X"D4",X"E0",X"E8",X"EA",X"9E",X"EA",X"97",X"00",X"06",X"00",X"E9",X"E0",X"19",X"E0",X"5D",
		X"E0",X"00",X"E2",X"44",X"E2",X"C4",X"E2",X"7E",X"EC",X"0D",X"E2",X"8F",X"E2",X"A1",X"E2",X"EB",
		X"90",X"9A",X"96",X"50",X"10",X"96",X"98",X"12",X"5C",X"6E",X"0F",X"6E",X"01",X"6F",X"04",X"A2",
		X"5E",X"5C",X"58",X"D2",X"10",X"6E",X"0F",X"6E",X"A4",X"10",X"90",X"58",X"12",X"D2",X"1A",X"94",
		X"8D",X"06",X"14",X"5E",X"5C",X"9A",X"96",X"10",X"1C",X"5E",X"94",X"10",X"10",X"10",X"A0",X"A0",
		X"01",X"E5",X"04",X"D8",X"10",X"60",X"62",X"64",X"A0",X"6E",X"07",X"6E",X"01",X"3A",X"06",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"2C",X"12",X"5C",X"2E",X"10",X"6E",X"0F",X"6E",X"01",
		X"2C",X"6E",X"03",X"6E",X"01",X"1A",X"02",X"2C",X"6E",X"01",X"50",X"02",X"2C",X"90",X"52",X"5C",
		X"02",X"2C",X"5A",X"52",X"16",X"56",X"D2",X"2C",X"A2",X"A0",X"10",X"DA",X"DC",X"DE",X"6E",X"CF",
		X"10",X"DA",X"DC",X"DE",X"6E",X"CF",X"6E",X"01",X"6C",X"6E",X"07",X"6E",X"01",X"1B",X"04",X"10",
		X"A8",X"01",X"43",X"45",X"4B",X"4D",X"6E",X"43",X"94",X"D2",X"10",X"10",X"5E",X"56",X"6E",X"4F",
		X"10",X"10",X"10",X"94",X"10",X"5A",X"6E",X"4F",X"52",X"5C",X"10",X"10",X"A2",X"10",X"16",X"94",
		X"01",X"40",X"06",X"A4",X"10",X"16",X"5E",X"52",X"18",X"52",X"98",X"10",X"6E",X"4F",X"6E",X"01",
		X"10",X"10",X"A4",X"10",X"16",X"94",X"1A",X"18",X"06",X"1C",X"94",X"1A",X"1A",X"10",X"10",X"90",
		X"87",X"8D",X"41",X"8D",X"87",X"8D",X"41",X"8D",X"BE",X"F0",X"F0",X"BA",X"B6",X"70",X"83",X"8B",
		X"8B",X"85",X"87",X"49",X"45",X"41",X"0D",X"81",X"81",X"8D",X"83",X"41",X"03",X"FF",X"1E",X"A0",
		X"BE",X"20",X"5C",X"80",X"5A",X"80",X"58",X"80",X"3C",X"A0",X"3E",X"10",X"B0",X"B1",X"F7",X"E6",
		X"41",X"78",X"B2",X"B4",X"B6",X"B6",X"B2",X"87",X"F4",X"F0",X"BC",X"BA",X"8D",X"78",X"83",X"21",
		X"8D",X"06",X"10",X"12",X"18",X"18",X"52",X"98",X"10",X"12",X"98",X"10",X"10",X"10",X"A0",X"A0",
		X"01",X"D4",X"04",X"10",X"10",X"10",X"10",X"10",X"02",X"02",X"6E",X"01",X"90",X"10",X"10",X"10",
		X"5A",X"52",X"18",X"9E",X"12",X"D2",X"10",X"5A",X"10",X"6E",X"03",X"6E",X"01",X"6E",X"01",X"1B",
		X"1E",X"10",X"10",X"6E",X"03",X"6E",X"01",X"7C",X"56",X"D2",X"6E",X"03",X"6E",X"01",X"51",X"04",
		X"EC",X"02",X"A4",X"88",X"5C",X"53",X"0F",X"6E",X"1E",X"9A",X"94",X"1A",X"E6",X"E6",X"6E",X"0B",
		X"58",X"52",X"96",X"98",X"E6",X"E6",X"E6",X"E6",X"98",X"5E",X"14",X"5E",X"56",X"1A",X"E6",X"E6",
		X"16",X"94",X"D2",X"14",X"12",X"14",X"D2",X"E6",X"02",X"06",X"02",X"02",X"02",X"06",X"04",X"04",
		X"08",X"0C",X"04",X"04",X"04",X"04",X"08",X"04",X"02",X"02",X"02",X"02",X"04",X"08",X"08",X"08",
		X"0B",X"7E",X"95",X"F5",X"E4",X"28",X"C0",X"B5",X"21",X"88",X"29",X"8E",X"61",X"8C",X"69",X"8C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B6",X"20",X"00",X"48",X"00",X"44",X"CE",X"00",
		X"D2",X"02",X"0C",X"40",X"00",X"00",X"04",X"00",X"D2",X"04",X"0C",X"44",X"00",X"00",X"04",X"00",
		X"D2",X"08",X"0C",X"48",X"00",X"0C",X"04",X"00",X"AC",X"0E",X"0F",X"7E",X"00",X"00",X"08",X"00",
		X"6E",X"01",X"76",X"04",X"96",X"98",X"12",X"94",X"01",X"48",X"06",X"5A",X"96",X"10",X"90",X"12",
		X"01",X"76",X"04",X"10",X"10",X"10",X"10",X"10",X"76",X"04",X"12",X"16",X"98",X"10",X"52",X"52",
		X"76",X"04",X"98",X"50",X"1A",X"D2",X"10",X"5A",X"06",X"5E",X"98",X"98",X"5E",X"5A",X"1A",X"5C",
		X"80",X"19",X"91",X"EC",X"E4",X"04",X"5C",X"3F",X"EB",X"EC",X"C9",X"EC",X"07",X"A8",X"25",X"EC",
		X"DB",X"7C",X"A0",X"DB",X"3C",X"A2",X"AC",X"03",X"DB",X"7C",X"90",X"DB",X"3C",X"92",X"AC",X"09",
		X"FF",X"4A",X"DB",X"42",X"DB",X"7C",X"00",X"DB",X"06",X"AC",X"41",X"DB",X"7C",X"80",X"DB",X"3C",
		X"AC",X"41",X"DB",X"7C",X"20",X"DB",X"3C",X"22",X"47",X"DB",X"7C",X"A0",X"DB",X"3C",X"A2",X"AA",
		X"DB",X"7C",X"10",X"DB",X"3C",X"12",X"AA",X"DB",X"7C",X"90",X"DB",X"3C",X"92",X"AA",X"DB",X"7C",
		X"E6",X"E6",X"6E",X"03",X"6E",X"01",X"1B",X"04",X"E6",X"E6",X"E6",X"E6",X"6E",X"03",X"6E",X"01",
		X"14",X"9A",X"96",X"1A",X"E6",X"E6",X"6E",X"07",X"90",X"E6",X"E6",X"E6",X"E6",X"E6",X"E6",X"E6",
		X"6E",X"03",X"6E",X"81",X"7C",X"04",X"96",X"9A",X"5A",X"12",X"5C",X"6E",X"43",X"6E",X"01",X"5A",
		X"00",X"00",X"6C",X"01",X"0D",X"47",X"4B",X"4D",X"10",X"10",X"6E",X"89",X"6E",X"81",X"A4",X"01",
		X"10",X"10",X"6E",X"4F",X"6E",X"01",X"44",X"06",X"5E",X"5C",X"1A",X"6E",X"4F",X"6E",X"01",X"44",
		X"4F",X"6E",X"01",X"48",X"06",X"90",X"9A",X"16",X"4C",X"06",X"98",X"12",X"14",X"58",X"1A",X"10",
		X"90",X"94",X"52",X"1E",X"50",X"98",X"6E",X"4F",X"4F",X"6E",X"01",X"76",X"02",X"2C",X"12",X"5E",
		X"EA",X"5E",X"22",X"00",X"5A",X"9F",X"77",X"F2",X"84",X"53",X"64",X"D5",X"14",X"D5",X"D4",X"D5",
		X"BA",X"B2",X"BA",X"B2",X"70",X"70",X"3A",X"3C",X"78",X"B2",X"BA",X"B6",X"76",X"78",X"B6",X"BC",
		X"B2",X"B6",X"B8",X"BA",X"74",X"76",X"78",X"B6",X"B2",X"BA",X"B2",X"70",X"50",X"10",X"70",X"3E",
		X"BA",X"B6",X"B2",X"B2",X"B6",X"8B",X"BA",X"B6",X"BC",X"74",X"78",X"83",X"81",X"83",X"FF",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"10",X"6E",X"07",X"6E",X"01",X"7C",X"04",X"10",X"6E",X"07",X"6E",X"01",X"7C",X"04",X"5A",
		X"5C",X"6E",X"43",X"6E",X"01",X"7C",X"04",X"10",X"6E",X"0B",X"6E",X"01",X"EA",X"04",X"10",X"10",
		X"A2",X"10",X"6E",X"03",X"6E",X"01",X"7C",X"04",X"0F",X"6E",X"01",X"76",X"04",X"54",X"9A",X"5C",
		X"4F",X"6E",X"01",X"76",X"04",X"9E",X"52",X"98",X"6E",X"01",X"76",X"04",X"98",X"50",X"1A",X"10",
		X"02",X"02",X"06",X"02",X"02",X"02",X"08",X"02",X"02",X"78",X"0A",X"02",X"02",X"02",X"C0",X"08",
		X"06",X"08",X"8C",X"08",X"06",X"02",X"02",X"02",X"02",X"04",X"08",X"04",X"08",X"4C",X"04",X"08",
		X"04",X"08",X"04",X"02",X"02",X"02",X"02",X"04",X"02",X"04",X"02",X"44",X"02",X"02",X"02",X"02",
		X"08",X"00",X"04",X"10",X"02",X"EC",X"EA",X"80",X"02",X"EC",X"EA",X"80",X"22",X"25",X"10",X"82",
		X"C8",X"B0",X"47",X"40",X"00",X"02",X"0C",X"00",X"9C",X"48",X"FF",X"49",X"00",X"04",X"40",X"00",
		X"AC",X"E0",X"FD",X"84",X"F1",X"08",X"4E",X"F9",X"02",X"04",X"08",X"40",X"80",X"20",X"10",X"01",
		X"05",X"45",X"85",X"C5",X"27",X"6B",X"E1",X"17",X"DD",X"E8",X"DF",X"E8",X"B3",X"06",X"B5",X"06",
		X"F2",X"F2",X"F0",X"8F",X"BC",X"BA",X"B8",X"B6",X"83",X"8B",X"41",X"8B",X"83",X"8B",X"41",X"8B",
		X"85",X"A8",X"17",X"EC",X"AF",X"EC",X"8F",X"A8",X"A4",X"02",X"5E",X"17",X"4D",X"0A",X"5B",X"14",
		X"4D",X"0A",X"7F",X"C8",X"A0",X"7F",X"C8",X"4E",X"0A",X"7F",X"C8",X"A2",X"17",X"4D",X"0A",X"7F",
		X"17",X"4D",X"0A",X"7F",X"C8",X"80",X"17",X"4D",X"E4",X"02",X"5E",X"E8",X"3D",X"4E",X"A4",X"02",
		X"03",X"EE",X"57",X"1E",X"60",X"A6",X"DB",X"42",X"DB",X"7C",X"80",X"DB",X"3C",X"82",X"AC",X"0F",
		X"14",X"A1",X"14",X"81",X"14",X"B0",X"14",X"90",X"12",X"A1",X"12",X"81",X"12",X"B0",X"12",X"90",
		X"10",X"A1",X"10",X"6F",X"10",X"6D",X"10",X"6B",X"10",X"53",X"10",X"73",X"10",X"42",X"12",X"62",
		X"12",X"53",X"12",X"73",X"12",X"42",X"14",X"62",X"14",X"53",X"14",X"55",X"14",X"57",X"14",X"59",
		X"14",X"53",X"14",X"55",X"14",X"57",X"14",X"59",X"14",X"14",X"5F",X"14",X"91",X"14",X"00",X"5E",
		X"5A",X"96",X"10",X"90",X"12",X"16",X"E6",X"5A",X"02",X"2C",X"12",X"56",X"12",X"14",X"1A",X"52",
		X"5A",X"12",X"16",X"56",X"D2",X"2C",X"6E",X"03",X"56",X"D2",X"2C",X"6E",X"07",X"6E",X"01",X"50",
		X"6E",X"07",X"6E",X"01",X"BC",X"04",X"80",X"10",X"6E",X"01",X"F0",X"04",X"88",X"10",X"AA",X"A0",
		X"DA",X"04",X"60",X"62",X"64",X"66",X"68",X"6A",X"5E",X"52",X"56",X"12",X"56",X"1A",X"E6",X"E6",
		X"6E",X"81",X"08",X"06",X"5A",X"1A",X"5A",X"5E",X"6E",X"01",X"08",X"06",X"14",X"12",X"18",X"10",
		X"6E",X"01",X"40",X"06",X"A2",X"10",X"16",X"5E",X"1A",X"18",X"52",X"98",X"10",X"6E",X"4F",X"6E",
		X"5C",X"96",X"10",X"A2",X"10",X"16",X"94",X"1A",X"40",X"06",X"A2",X"10",X"16",X"5E",X"52",X"5C",
		X"52",X"98",X"96",X"6E",X"4F",X"6E",X"01",X"40",X"58",X"12",X"D2",X"10",X"10",X"10",X"10",X"10",
		X"87",X"8D",X"41",X"8D",X"AD",X"A7",X"BA",X"BC",X"41",X"8B",X"83",X"8B",X"41",X"8B",X"0D",X"8D",
		X"81",X"8D",X"8B",X"81",X"81",X"0D",X"81",X"8D",X"56",X"80",X"58",X"80",X"5A",X"80",X"5C",X"80",
		X"54",X"80",X"1E",X"80",X"1C",X"80",X"3A",X"A0",X"B3",X"00",X"B5",X"04",X"B7",X"44",X"B9",X"00",
		X"78",X"B6",X"BA",X"BC",X"BC",X"BA",X"8D",X"F8",X"41",X"BA",X"BC",X"BE",X"F0",X"B2",X"B6",X"B8",
		X"52",X"5E",X"5C",X"12",X"58",X"10",X"10",X"10",X"A0",X"10",X"DA",X"DC",X"DE",X"6E",X"8B",X"6E",
		X"10",X"10",X"6E",X"0E",X"0E",X"0E",X"02",X"02",X"6E",X"0F",X"6E",X"01",X"D6",X"04",X"D8",X"10",
		X"1C",X"1E",X"10",X"16",X"5E",X"10",X"10",X"10",X"04",X"E6",X"5A",X"12",X"18",X"10",X"18",X"5E",
		X"04",X"10",X"10",X"10",X"14",X"58",X"52",X"5C",X"E6",X"56",X"52",X"58",X"58",X"1A",X"94",X"10",
		X"01",X"57",X"04",X"10",X"56",X"52",X"5A",X"12",X"6E",X"01",X"57",X"04",X"10",X"96",X"98",X"D2",
		X"6E",X"0B",X"6E",X"01",X"5D",X"04",X"10",X"5E",X"E6",X"6E",X"0F",X"6E",X"01",X"5D",X"04",X"10",
		X"E6",X"E6",X"E6",X"6E",X"0F",X"6E",X"01",X"02",X"04",X"02",X"02",X"02",X"02",X"04",X"08",X"08",
		X"08",X"08",X"08",X"0C",X"04",X"04",X"04",X"04",X"0C",X"04",X"04",X"04",X"04",X"0C",X"08",X"0A",
		X"81",X"88",X"89",X"4E",X"C1",X"8A",X"C9",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C9",X"8C",X"C9",X"8C",X"C9",X"8C",X"B4",X"20",X"F7",X"0F",X"00",X"04",X"4E",X"00",
		X"D2",X"02",X"0C",X"42",X"00",X"00",X"04",X"00",X"D2",X"06",X"0C",X"46",X"00",X"00",X"04",X"00",
		X"28",X"00",X"0C",X"40",X"04",X"00",X"44",X"00",X"B0",X"08",X"00",X"00",X"00",X"00",X"40",X"00",
		X"94",X"52",X"5C",X"1E",X"10",X"6E",X"4F",X"6E",X"16",X"E6",X"5A",X"1A",X"5C",X"6E",X"4F",X"6E",
		X"10",X"10",X"10",X"10",X"6E",X"0B",X"6E",X"01",X"52",X"2C",X"10",X"10",X"6E",X"0F",X"6E",X"01",
		X"1A",X"1A",X"98",X"6E",X"4F",X"6E",X"01",X"48",X"6E",X"4F",X"6E",X"01",X"E4",X"04",X"5C",X"FD",
		X"DE",X"08",X"8D",X"EC",X"47",X"EC",X"48",X"00",X"41",X"A8",X"67",X"EC",X"4B",X"A8",X"A3",X"EC",
		X"DB",X"7C",X"10",X"DB",X"3C",X"12",X"AC",X"03",X"53",X"4A",X"6F",X"E3",X"F5",X"22",X"EE",X"0C",
		X"3C",X"02",X"AA",X"DB",X"7C",X"04",X"DB",X"3C",X"82",X"AA",X"DB",X"7C",X"84",X"DB",X"3C",X"86",
		X"AA",X"DB",X"7C",X"24",X"DB",X"3C",X"26",X"AC",X"DB",X"7C",X"A4",X"DB",X"3C",X"A6",X"AC",X"05",
		X"7C",X"14",X"DB",X"3C",X"16",X"AC",X"05",X"DB",X"94",X"DB",X"3C",X"96",X"AC",X"07",X"53",X"91",
		X"10",X"9A",X"94",X"16",X"50",X"52",X"5C",X"E6",X"51",X"04",X"10",X"5A",X"12",X"16",X"50",X"52",
		X"6E",X"01",X"51",X"04",X"10",X"94",X"5E",X"5A",X"6E",X"07",X"6E",X"01",X"2A",X"01",X"03",X"0B",
		X"90",X"1A",X"94",X"10",X"90",X"12",X"16",X"E6",X"12",X"5C",X"6E",X"43",X"6E",X"01",X"6E",X"81",
		X"6E",X"4F",X"6E",X"81",X"A0",X"01",X"10",X"10",X"43",X"45",X"4B",X"4D",X"6E",X"43",X"6E",X"81",
		X"14",X"5E",X"5C",X"9A",X"96",X"10",X"10",X"5C",X"06",X"14",X"5E",X"5C",X"9A",X"96",X"10",X"6E",
		X"56",X"5A",X"12",X"5C",X"6E",X"4F",X"6E",X"01",X"10",X"6E",X"4F",X"6E",X"01",X"4C",X"06",X"9A",
		X"6E",X"01",X"44",X"04",X"A0",X"A0",X"A0",X"6E",X"96",X"9A",X"56",X"1A",X"2C",X"6E",X"0B",X"6E",
		X"22",X"B5",X"E2",X"9F",X"84",X"26",X"86",X"FC",X"B4",X"D5",X"7F",X"0A",X"02",X"7F",X"80",X"88",
		X"3E",X"61",X"67",X"69",X"49",X"0D",X"BC",X"BA",X"F4",X"F0",X"F0",X"BC",X"B6",X"78",X"65",X"61",
		X"BA",X"BC",X"BE",X"F0",X"B2",X"B6",X"B8",X"BA",X"70",X"65",X"63",X"65",X"74",X"30",X"45",X"BC",
		X"B2",X"70",X"70",X"32",X"36",X"74",X"61",X"78",X"2C",X"0F",X"B0",X"B1",X"CB",X"E8",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"10",X"10",X"90",X"52",X"5C",X"56",X"D2",X"96",X"10",X"90",X"12",X"16",X"E6",X"5A",X"12",
		X"10",X"10",X"52",X"5C",X"56",X"D2",X"10",X"10",X"A2",X"E2",X"E0",X"A0",X"E4",X"A2",X"E2",X"E0",
		X"10",X"10",X"10",X"10",X"96",X"9A",X"1A",X"6E",X"52",X"5E",X"94",X"10",X"10",X"10",X"10",X"6E",
		X"50",X"10",X"10",X"10",X"10",X"10",X"6E",X"4F",X"16",X"50",X"12",X"96",X"1A",X"10",X"6E",X"4F",
		X"02",X"02",X"06",X"02",X"02",X"08",X"02",X"02",X"08",X"C0",X"0A",X"02",X"02",X"02",X"8E",X"04",
		X"BC",X"02",X"02",X"02",X"02",X"06",X"02",X"02",X"04",X"08",X"04",X"08",X"46",X"02",X"02",X"02",
		X"04",X"04",X"4C",X"04",X"08",X"04",X"08",X"04",X"06",X"02",X"02",X"02",X"06",X"02",X"02",X"06",
		X"10",X"10",X"4C",X"EA",X"EC",X"80",X"15",X"16",X"5E",X"E4",X"AC",X"88",X"C4",X"2F",X"51",X"86",
		X"C8",X"B0",X"47",X"40",X"00",X"02",X"0C",X"00",X"9C",X"00",X"04",X"44",X"0E",X"06",X"48",X"00",
		X"24",X"02",X"02",X"0C",X"00",X"02",X"0E",X"00",X"00",X"9E",X"D8",X"32",X"3E",X"7A",X"B8",X"F6",
		X"99",X"E6",X"B7",X"E6",X"D0",X"E8",X"8B",X"E8",X"B7",X"44",X"B9",X"04",X"81",X"F8",X"F6",X"F4",
		X"B6",X"B4",X"83",X"61",X"41",X"30",X"54",X"58",X"83",X"8B",X"41",X"8B",X"8B",X"C1",X"89",X"8F",
		X"53",X"EC",X"53",X"7F",X"C8",X"48",X"EC",X"30",X"8D",X"17",X"4D",X"0A",X"7F",X"C8",X"4A",X"17",
		X"17",X"4D",X"0A",X"7F",X"C8",X"6E",X"17",X"4D",X"C8",X"A6",X"17",X"4D",X"0A",X"7F",X"C8",X"4C",
		X"0A",X"6F",X"A4",X"88",X"5C",X"17",X"F8",X"0A",X"5E",X"5E",X"57",X"03",X"0C",X"00",X"DB",X"22",
		X"DB",X"7C",X"00",X"DB",X"3C",X"02",X"AC",X"0F",X"DB",X"7C",X"20",X"DB",X"3C",X"22",X"AC",X"45",
		X"14",X"A0",X"14",X"80",X"14",X"B1",X"12",X"91",X"12",X"A0",X"12",X"80",X"12",X"B1",X"10",X"91",
		X"10",X"69",X"10",X"67",X"10",X"65",X"10",X"63",X"12",X"52",X"12",X"72",X"12",X"43",X"12",X"63",
		X"14",X"52",X"14",X"72",X"14",X"43",X"14",X"63",X"14",X"5B",X"14",X"5D",X"14",X"5F",X"14",X"91",
		X"14",X"5B",X"14",X"5D",X"14",X"5F",X"14",X"91",X"53",X"00",X"00",X"A0",X"4B",X"00",X"BA",X"B6");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
