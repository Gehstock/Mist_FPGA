library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity col2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(7 downto 0);
	data : out std_logic_vector(3 downto 0)
);
end entity;

architecture prom of col2 is
	type rom is array(0 to  255) of std_logic_vector(3 downto 0);
	signal rom_data: rom := (
		"1111","1100","0000","1111","1111","1011","1111","0000","1111","1010","1111","1101","1111","1100","1111","0011",
		"1111","0011","1011","1111","1111","0000","1101","0011","1111","1111","1100","0000","1111","1111","1010","0000",
		"1111","1111","1010","0011","1111","0000","0011","0101","1111","1101","0000","0101","1111","1100","0011","1010",
		"1111","0000","0000","1100","1111","1111","1011","0011","1111","1110","1010","1100","1111","1011","1111","1111",
		"1111","1100","0000","1111","1111","1011","1111","0000","1111","1010","1111","1101","1111","0011","1010","0000",
		"1111","0011","1010","0000","1111","0011","1010","0000","1111","0011","1010","0000","1111","1111","1010","0000",
		"1111","1111","1010","0011","1111","0000","0011","0101","1111","1101","0000","0101","1111","1100","0011","1010",
		"1111","0000","0000","1100","1111","1111","1011","0011","1111","1110","1010","1100","1111","1011","1111","1111",
		"1111","1100","0000","1111","1111","1011","1111","0000","1111","1010","1111","1101","1111","1010","1111","0000",
		"1111","1010","1111","0000","1111","1010","1111","0000","1111","1010","1111","0000","1111","1111","1010","0000",
		"1111","1111","1010","0011","1111","0000","0011","0101","1111","1101","0000","0101","1111","1100","0011","1010",
		"1111","0000","0000","1100","1111","1111","1011","0011","1111","1110","1010","1100","1111","1011","1111","1111",
		"1111","1100","0000","1111","1111","1011","1111","0000","1111","1010","1111","1101","1111","1100","0000","1011",
		"1111","1100","0000","1011","1111","1100","0000","1011","1111","1100","0000","1011","1111","1111","1010","0000",
		"1111","1111","1010","0011","1111","0000","0011","0101","1111","1101","0000","0101","1111","1100","0011","1010",
		"1111","0000","0000","1100","1111","1111","1011","0011","1111","1110","1010","1100","1111","1011","1111","1111");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
