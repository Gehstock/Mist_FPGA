library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity twotiger_sp_bits_4 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of twotiger_sp_bits_4 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0F",X"EE",X"00",X"00",
		X"0E",X"EF",X"0E",X"00",X"0E",X"EF",X"EF",X"00",X"0E",X"EF",X"EE",X"00",X"EE",X"5E",X"5E",X"00",
		X"5F",X"55",X"55",X"00",X"5E",X"55",X"55",X"00",X"5E",X"55",X"FF",X"00",X"6F",X"FF",X"EE",X"00",
		X"EE",X"EE",X"00",X"00",X"0E",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",
		X"0E",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"0E",X"00",X"00",X"0E",X"EF",X"00",X"00",
		X"0F",X"FF",X"00",X"00",X"0E",X"FF",X"00",X"00",X"EE",X"FF",X"00",X"00",X"5E",X"55",X"0E",X"00",
		X"5E",X"55",X"EF",X"00",X"E6",X"55",X"FF",X"00",X"0E",X"FF",X"5E",X"00",X"0F",X"EE",X"55",X"00",
		X"0E",X"E0",X"55",X"00",X"00",X"E0",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"E5",X"00",
		X"0E",X"00",X"E5",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"0E",X"00",X"00",X"55",X"EE",X"00",X"00",
		X"55",X"EF",X"00",X"00",X"E5",X"FF",X"00",X"00",X"EF",X"EF",X"00",X"00",X"EE",X"5E",X"E0",X"00",
		X"0E",X"55",X"5E",X"00",X"00",X"55",X"55",X"00",X"00",X"EE",X"55",X"00",X"00",X"FE",X"55",X"00",
		X"0F",X"FF",X"65",X"00",X"00",X"FF",X"FE",X"00",X"00",X"FF",X"EE",X"00",X"00",X"FF",X"E5",X"00",
		X"00",X"FE",X"E5",X"00",X"00",X"E0",X"E5",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"0E",X"EE",X"00",X"00",
		X"E5",X"FF",X"00",X"00",X"55",X"FF",X"00",X"00",X"55",X"5F",X"0E",X"00",X"E6",X"55",X"EE",X"00",
		X"0E",X"55",X"EF",X"00",X"0F",X"55",X"FF",X"00",X"0E",X"FE",X"FF",X"00",X"0E",X"EE",X"EE",X"00",
		X"F0",X"FF",X"55",X"00",X"00",X"FF",X"55",X"00",X"00",X"FE",X"55",X"00",X"00",X"E0",X"55",X"00",
		X"00",X"00",X"E5",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"EE",X"E0",X"00",X"00",X"E5",X"5E",X"00",X"00",X"55",X"55",X"00",X"00",
		X"E5",X"5F",X"00",X"00",X"E6",X"5F",X"00",X"00",X"0E",X"5E",X"00",X"00",X"00",X"55",X"EE",X"00",
		X"00",X"55",X"FF",X"00",X"0E",X"55",X"FF",X"00",X"F0",X"EE",X"FF",X"00",X"00",X"FE",X"EF",X"00",
		X"00",X"F6",X"55",X"00",X"00",X"FE",X"55",X"00",X"00",X"E0",X"55",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"00",X"00",X"00",X"5E",X"E0",X"00",X"00",X"55",X"5E",X"00",X"00",X"E5",X"5F",X"00",X"00",
		X"E5",X"5F",X"00",X"00",X"0E",X"5E",X"00",X"00",X"0E",X"5E",X"00",X"00",X"00",X"55",X"0E",X"00",
		X"00",X"55",X"EF",X"00",X"0F",X"55",X"EF",X"00",X"0F",X"E1",X"FF",X"00",X"00",X"FE",X"FF",X"00",
		X"00",X"FE",X"EF",X"00",X"00",X"FF",X"5E",X"00",X"00",X"FF",X"55",X"00",X"00",X"FE",X"55",X"00",
		X"00",X"EE",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0E",X"EE",X"E0",X"00",X"0E",X"5E",X"E0",X"00",X"0E",X"55",X"E0",X"00",
		X"00",X"5E",X"E0",X"00",X"00",X"EF",X"00",X"00",X"00",X"EF",X"00",X"00",X"00",X"5E",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"E5",X"EE",X"00",X"00",X"F1",X"EE",X"00",X"00",X"FE",X"FF",X"00",
		X"00",X"FE",X"EF",X"00",X"00",X"FF",X"5E",X"00",X"00",X"FF",X"55",X"00",X"00",X"FF",X"55",X"00",
		X"00",X"EE",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",
		X"EE",X"00",X"00",X"00",X"E5",X"E0",X"00",X"00",X"E6",X"5E",X"E0",X"00",X"EE",X"55",X"E0",X"00",
		X"0E",X"5E",X"E0",X"00",X"00",X"5E",X"E0",X"00",X"00",X"EF",X"00",X"00",X"0E",X"5E",X"00",X"00",
		X"0E",X"55",X"00",X"00",X"F0",X"55",X"EE",X"00",X"00",X"EE",X"FF",X"00",X"00",X"EF",X"FF",X"00",
		X"00",X"EE",X"FF",X"00",X"00",X"FF",X"EF",X"00",X"00",X"FF",X"5E",X"00",X"00",X"FE",X"55",X"00",
		X"00",X"E0",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"5E",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",
		X"0E",X"EE",X"00",X"00",X"0E",X"55",X"00",X"00",X"00",X"55",X"E0",X"00",X"00",X"E5",X"FE",X"00",
		X"00",X"55",X"FE",X"00",X"00",X"5E",X"FE",X"00",X"0F",X"5E",X"E0",X"00",X"00",X"5E",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E1",X"0E",X"00",X"00",X"EF",X"EF",X"00",
		X"00",X"FE",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"EE",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"E5",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"5E",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"E0",X"00",X"00",X"0E",X"00",X"00",X"00",
		X"0E",X"EE",X"00",X"00",X"0E",X"55",X"00",X"00",X"00",X"55",X"E0",X"00",X"00",X"E5",X"FE",X"00",
		X"00",X"55",X"FE",X"00",X"0F",X"5E",X"FE",X"00",X"00",X"5E",X"FE",X"00",X"00",X"55",X"E0",X"00",
		X"00",X"5E",X"00",X"00",X"00",X"FE",X"00",X"00",X"00",X"E1",X"00",X"00",X"00",X"EF",X"E0",X"00",
		X"00",X"EE",X"FE",X"00",X"00",X"FE",X"FF",X"00",X"00",X"EE",X"FF",X"00",X"00",X"00",X"FE",X"00",
		X"00",X"00",X"FE",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"5E",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"E5",X"E0",X"00",X"00",X"5E",X"FE",X"00",
		X"00",X"55",X"FE",X"00",X"0E",X"55",X"FE",X"00",X"00",X"5E",X"FE",X"00",X"00",X"5E",X"E0",X"00",
		X"00",X"55",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"FE",X"00",X"00",X"00",X"E1",X"00",X"00",
		X"00",X"FE",X"E0",X"00",X"00",X"EE",X"FE",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"FE",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"FE",X"00",X"00",X"00",X"E0",X"00",X"00",
		X"00",X"5E",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"5E",X"EE",X"00",X"00",X"55",X"FE",X"00",
		X"00",X"55",X"FF",X"00",X"00",X"55",X"FF",X"00",X"00",X"55",X"FE",X"00",X"00",X"55",X"E0",X"00",
		X"00",X"55",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E1",X"00",X"00",X"00",X"E1",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"EE",X"E0",X"00",X"00",X"E0",X"FE",X"00",X"00",X"00",X"FE",X"00",
		X"00",X"00",X"FE",X"00",X"00",X"0E",X"E0",X"00",X"00",X"0E",X"5E",X"00",X"00",X"0E",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"5E",X"00",X"00",X"00",X"E5",X"00",X"00",X"0F",X"5E",X"00",X"00",X"0F",X"5E",X"E0",X"00",
		X"00",X"55",X"FE",X"00",X"00",X"55",X"FE",X"00",X"00",X"5E",X"FF",X"00",X"00",X"5E",X"FE",X"00",
		X"00",X"5E",X"EE",X"00",X"00",X"E5",X"E0",X"00",X"00",X"1E",X"00",X"00",X"00",X"1E",X"00",X"00",
		X"00",X"EF",X"00",X"00",X"00",X"E6",X"00",X"00",X"00",X"0E",X"E0",X"00",X"00",X"00",X"FE",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"E5",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"5F",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"55",X"EE",X"00",X"00",X"55",X"FE",X"00",X"00",X"5E",X"FF",X"00",
		X"00",X"55",X"FF",X"00",X"00",X"E5",X"FE",X"00",X"00",X"1E",X"E0",X"00",X"00",X"1E",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E6",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"55",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"5E",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"EF",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"EE",X"00",X"00",X"55",X"FF",X"00",
		X"00",X"55",X"FF",X"00",X"00",X"E5",X"FF",X"00",X"00",X"E5",X"FE",X"00",X"00",X"E5",X"E0",X"00",
		X"00",X"55",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"E5",X"00",X"00",
		X"00",X"E6",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"55",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"E5",X"00",X"00",
		X"00",X"F5",X"00",X"00",X"00",X"65",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"E2",X"00",X"00",
		X"00",X"65",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"65",X"00",X"00",X"00",X"F5",X"00",X"00",
		X"00",X"65",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"65",X"00",X"00",X"00",X"E5",X"00",X"00",
		X"00",X"FE",X"00",X"00",X"00",X"1E",X"00",X"00",X"00",X"1E",X"00",X"00",X"00",X"FE",X"00",X"00",
		X"00",X"E5",X"00",X"00",X"00",X"65",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"E5",X"00",X"00",
		X"00",X"E5",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"EE",X"EE",X"00",X"00",X"99",X"99",X"00",X"EE",X"99",X"99",X"00",X"BB",X"EE",X"99",X"00",
		X"BB",X"BB",X"99",X"00",X"EB",X"BB",X"EE",X"E0",X"EB",X"EE",X"BB",X"E0",X"EB",X"99",X"BB",X"00",
		X"BB",X"99",X"BB",X"00",X"EE",X"99",X"BE",X"00",X"00",X"EE",X"EE",X"00",X"00",X"99",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9E",X"00",X"00",
		X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"EE",X"EE",X"00",X"00",X"BB",X"AA",X"00",X"EE",X"BB",X"AA",X"00",X"AA",X"BB",X"EE",X"00",
		X"AA",X"BB",X"BB",X"00",X"EE",X"EE",X"BB",X"E0",X"BB",X"BB",X"BB",X"E0",X"BB",X"BB",X"BB",X"E0",
		X"BE",X"BB",X"BB",X"E0",X"EF",X"EE",X"BB",X"00",X"0E",X"1E",X"BB",X"00",X"00",X"BB",X"EE",X"00",
		X"00",X"1E",X"00",X"00",X"00",X"BE",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9E",X"00",X"00",
		X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E1",X"00",X"00",X"00",X"3F",X"00",X"00",
		X"00",X"3F",X"00",X"00",X"00",X"1F",X"00",X"00",X"00",X"E3",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"2E",X"00",X"00",X"00",X"22",X"00",X"00",
		X"03",X"22",X"F0",X"00",X"EE",X"EF",X"00",X"00",X"3E",X"EF",X"30",X"00",X"EE",X"EE",X"00",X"00",
		X"EE",X"EE",X"EE",X"00",X"EE",X"EE",X"EE",X"00",X"EE",X"EE",X"F2",X"00",X"2E",X"EE",X"EE",X"00",
		X"2E",X"33",X"E2",X"00",X"EE",X"F1",X"EE",X"E0",X"EE",X"FF",X"E2",X"E0",X"EE",X"3F",X"E2",X"00",
		X"2E",X"11",X"E2",X"00",X"E1",X"11",X"2E",X"00",X"E1",X"13",X"EE",X"00",X"EE",X"13",X"00",X"00",
		X"E1",X"EE",X"EE",X"00",X"E1",X"FE",X"3E",X"00",X"E1",X"FE",X"1E",X"00",X"11",X"EE",X"1E",X"00",
		X"1E",X"E2",X"EE",X"00",X"EE",X"22",X"03",X"00",X"00",X"22",X"00",X"00",X"00",X"2E",X"00",X"00",
		X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"1E",X"00",X"00",X"03",X"22",X"00",X"00",
		X"03",X"22",X"11",X"00",X"EE",X"EF",X"11",X"00",X"3E",X"EF",X"11",X"00",X"E1",X"EE",X"10",X"00",
		X"11",X"EE",X"1E",X"00",X"1E",X"EE",X"13",X"00",X"EE",X"EE",X"12",X"00",X"3E",X"EE",X"3E",X"00",
		X"13",X"EE",X"13",X"00",X"11",X"EE",X"1E",X"E0",X"EE",X"EE",X"13",X"E0",X"1E",X"EE",X"11",X"00",
		X"2E",X"EE",X"E1",X"00",X"1E",X"EE",X"2E",X"00",X"EE",X"EE",X"EE",X"00",X"EE",X"EE",X"33",X"00",
		X"3E",X"EE",X"13",X"00",X"EE",X"EE",X"33",X"00",X"EE",X"EE",X"EE",X"00",X"EE",X"EE",X"EE",X"00",
		X"EE",X"E2",X"EE",X"00",X"EE",X"22",X"03",X"00",X"10",X"22",X"00",X"00",X"11",X"2E",X"00",X"00",
		X"31",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"2B",X"EA",X"00",X"00",X"2B",X"AE",X"00",X"00",X"00",X"AA",X"00",X"00",X"A2",X"AA",X"00",X"00",
		X"AA",X"AA",X"EE",X"00",X"EE",X"A1",X"AA",X"00",X"EE",X"33",X"3A",X"00",X"0E",X"A3",X"BA",X"00",
		X"0E",X"A3",X"EA",X"00",X"0E",X"AA",X"EE",X"00",X"0E",X"AA",X"EE",X"00",X"0E",X"AA",X"3E",X"00",
		X"0E",X"AA",X"EE",X"00",X"EE",X"A3",X"BB",X"00",X"EE",X"A3",X"9B",X"00",X"0E",X"39",X"99",X"00",
		X"EE",X"99",X"99",X"00",X"EB",X"99",X"EE",X"00",X"EB",X"99",X"00",X"00",X"E9",X"EE",X"00",X"00",
		X"E9",X"00",X"00",X"00",X"EE",X"00",X"E0",X"00",X"00",X"00",X"3E",X"00",X"00",X"00",X"3E",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"AE",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"EA",X"00",X"00",X"00",X"EA",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"AE",X"00",X"00",X"00",X"A1",X"00",X"00",X"00",X"AE",X"00",X"00",
		X"00",X"2E",X"00",X"00",X"00",X"E2",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AE",X"00",X"00",
		X"00",X"AE",X"00",X"00",X"0A",X"0A",X"00",X"00",X"AA",X"0A",X"00",X"00",X"AE",X"EE",X"00",X"00",
		X"E0",X"0E",X"00",X"00",X"0E",X"AA",X"00",X"00",X"0E",X"EA",X"00",X"00",X"AE",X"EA",X"00",X"00",
		X"AE",X"EE",X"00",X"00",X"EE",X"EE",X"00",X"00",X"AE",X"AA",X"00",X"00",X"A1",X"AE",X"00",X"00",
		X"EA",X"AA",X"00",X"00",X"2A",X"EE",X"00",X"00",X"EE",X"AE",X"00",X"00",X"3E",X"AA",X"00",X"00",
		X"EE",X"AA",X"00",X"00",X"E2",X"E3",X"00",X"00",X"2A",X"AE",X"00",X"00",X"AE",X"E1",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",
		X"EE",X"EE",X"EE",X"00",X"EE",X"EE",X"77",X"00",X"AE",X"EE",X"77",X"00",X"AA",X"55",X"AA",X"00",
		X"AA",X"5E",X"EE",X"00",X"EE",X"EE",X"77",X"00",X"BB",X"EE",X"BB",X"00",X"BB",X"BE",X"EE",X"00",
		X"EB",X"BB",X"EE",X"00",X"EE",X"9B",X"99",X"E0",X"0E",X"B9",X"9B",X"E0",X"00",X"B9",X"2B",X"E0",
		X"00",X"FE",X"E0",X"20",X"00",X"00",X"F0",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"01",X"FF",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"F1",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"01",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"00",X"9E",X"00",X"00",X"EE",X"99",X"00",X"00",X"99",X"AA",X"00",X"00",X"99",X"1A",X"00",
		X"00",X"22",X"12",X"00",X"EE",X"EE",X"EE",X"00",X"E1",X"E2",X"EE",X"00",X"EE",X"1E",X"EE",X"00",
		X"0E",X"11",X"1E",X"00",X"00",X"31",X"11",X"00",X"0E",X"33",X"E1",X"00",X"E2",X"13",X"E1",X"00",
		X"2E",X"13",X"EE",X"00",X"2F",X"11",X"EE",X"E0",X"2E",X"11",X"EE",X"E0",X"22",X"11",X"EE",X"00",
		X"EE",X"11",X"EE",X"00",X"00",X"1E",X"1E",X"00",X"0F",X"E1",X"33",X"00",X"0E",X"11",X"E1",X"00",
		X"0E",X"E1",X"EE",X"00",X"0E",X"EE",X"EE",X"00",X"0E",X"2E",X"EE",X"00",X"3E",X"E2",X"EE",X"00",
		X"00",X"EE",X"EE",X"00",X"00",X"22",X"E0",X"00",X"00",X"22",X"E0",X"00",X"00",X"E2",X"E0",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"E0",X"21",X"00",X"11",X"2E",X"01",X"00",X"1A",X"99",X"11",X"00",X"1A",X"11",X"11",X"00",
		X"11",X"11",X"11",X"00",X"11",X"11",X"1E",X"00",X"3E",X"E1",X"EE",X"00",X"E1",X"EE",X"EE",X"00",
		X"3E",X"11",X"EE",X"00",X"11",X"EE",X"EE",X"00",X"11",X"EE",X"33",X"00",X"E1",X"EE",X"11",X"00",
		X"E1",X"EE",X"11",X"01",X"EE",X"EE",X"EE",X"10",X"EE",X"11",X"EE",X"00",X"3E",X"E1",X"EE",X"00",
		X"1E",X"E1",X"11",X"00",X"11",X"1E",X"EE",X"10",X"00",X"EE",X"E3",X"10",X"EE",X"1E",X"E3",X"10",
		X"E1",X"EE",X"E3",X"30",X"E1",X"EE",X"E3",X"00",X"31",X"EE",X"EE",X"00",X"13",X"31",X"EE",X"00",
		X"11",X"1E",X"11",X"00",X"12",X"11",X"11",X"00",X"11",X"11",X"EE",X"00",X"11",X"11",X"E0",X"00",
		X"EE",X"11",X"E1",X"00",X"EE",X"1E",X"03",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"02",X"00",X"6F",X"00",
		X"02",X"20",X"02",X"00",X"00",X"F0",X"F0",X"00",X"00",X"F0",X"20",X"00",X"62",X"F0",X"02",X"00",
		X"F0",X"FF",X"02",X"00",X"02",X"2F",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"26",X"00",X"00",
		X"00",X"26",X"00",X"20",X"60",X"26",X"00",X"20",X"FF",X"22",X"02",X"00",X"F2",X"22",X"22",X"00",
		X"22",X"22",X"22",X"00",X"02",X"22",X"20",X"00",X"02",X"22",X"00",X"00",X"00",X"22",X"00",X"20",
		X"00",X"22",X"00",X"20",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",
		X"00",X"60",X"00",X"00",X"00",X"26",X"00",X"00",X"00",X"02",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"00",X"00",X"62",X"02",X"00",X"00",X"00",X"62",X"60",X"00",X"00",X"66",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"66",X"02",X"00",X"60",X"22",X"00",X"00",X"20",X"62",X"60",X"00",
		X"00",X"62",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"66",X"00",X"00",
		X"00",X"62",X"02",X"00",X"62",X"62",X"60",X"20",X"20",X"26",X"60",X"00",X"00",X"26",X"22",X"60",
		X"00",X"22",X"22",X"60",X"00",X"22",X"20",X"60",X"00",X"22",X"20",X"00",X"00",X"22",X"20",X"00",
		X"00",X"70",X"20",X"00",X"00",X"72",X"20",X"00",X"00",X"72",X"20",X"00",X"00",X"22",X"20",X"00",
		X"00",X"22",X"20",X"00",X"00",X"22",X"20",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"88",X"00",X"00",X"00",X"86",X"00",X"00",X"00",X"64",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"4C",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"4E",X"00",X"00",X"00",X"9E",X"00",
		X"00",X"00",X"9E",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"9E",X"00",
		X"00",X"00",X"9E",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"9E",X"00",
		X"00",X"00",X"9E",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"EE",X"00",X"00",X"E7",X"F7",X"00",
		X"00",X"F7",X"F7",X"00",X"77",X"00",X"77",X"00",X"00",X"00",X"F0",X"00",X"FF",X"FF",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"E0",X"00",X"00",X"E6",X"FE",X"00",X"00",X"06",X"FF",X"00",X"00",X"00",X"EF",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"0E",X"AE",X"00",X"00",X"EE",X"FF",X"00",X"00",X"6E",X"FF",X"EE",X"00",
		X"66",X"FE",X"FF",X"E0",X"66",X"FE",X"66",X"FE",X"AA",X"FF",X"6B",X"FF",X"FF",X"FF",X"BF",X"BE",
		X"FF",X"FF",X"BB",X"E0",X"FF",X"EE",X"BB",X"00",X"FF",X"EE",X"EE",X"00",X"EE",X"EE",X"E0",X"00",
		X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",
		X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"EE",X"00",X"00",X"0E",X"9E",X"00",X"00",
		X"0E",X"9E",X"00",X"00",X"0E",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",
		X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"BE",X"00",X"00",X"00",X"EB",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"EE",X"E0",X"00",X"00",X"BB",X"EE",X"00",X"00",X"EB",X"BB",X"00",
		X"00",X"0E",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"77",X"00",X"77",X"F7",X"F7",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"0E",X"AA",X"00",X"00",X"EB",X"EE",X"00",X"00",X"0E",X"EF",X"00",
		X"00",X"00",X"CC",X"00",X"E7",X"7F",X"CC",X"F7",X"70",X"07",X"EE",X"07",X"00",X"00",X"77",X"00",
		X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"00",X"CC",X"00",X"E0",X"00",X"EC",X"00",X"E0",X"00",X"EC",X"EE",
		X"E0",X"00",X"CC",X"CC",X"EE",X"00",X"CC",X"EE",X"BE",X"00",X"EE",X"E0",X"BE",X"07",X"BB",X"E0",
		X"BB",X"07",X"BB",X"CC",X"EE",X"7F",X"EE",X"77",X"70",X"07",X"77",X"07",X"10",X"10",X"07",X"06",
		X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"2E",X"00",X"00",
		X"00",X"2E",X"00",X"00",X"00",X"2E",X"00",X"00",X"00",X"2E",X"00",X"00",X"00",X"2E",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"22",X"EE",X"00",X"00",X"22",X"E2",X"00",X"EE",X"EE",X"22",X"00",
		X"22",X"22",X"22",X"00",X"22",X"22",X"EE",X"00",X"22",X"EE",X"EE",X"00",X"22",X"22",X"E2",X"00",
		X"EE",X"22",X"EE",X"00",X"00",X"22",X"0E",X"00",X"00",X"EE",X"00",X"00",X"00",X"22",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"2E",X"00",X"00",X"00",X"2E",X"00",X"00",X"00",X"2E",X"00",X"00",
		X"00",X"2E",X"00",X"00",X"00",X"2E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"2E",X"00",X"00",X"00",X"66",X"00",X"00",
		X"02",X"62",X"50",X"00",X"26",X"E5",X"00",X"00",X"66",X"E5",X"60",X"00",X"EE",X"EE",X"00",X"00",
		X"EE",X"22",X"EE",X"00",X"EE",X"26",X"EE",X"00",X"EE",X"66",X"52",X"00",X"2E",X"22",X"EE",X"00",
		X"2E",X"2E",X"E2",X"00",X"EE",X"EE",X"EE",X"E0",X"EE",X"EE",X"E2",X"E0",X"EE",X"EE",X"E2",X"00",
		X"2E",X"EE",X"E2",X"00",X"E2",X"E2",X"2E",X"00",X"E2",X"22",X"EE",X"00",X"EE",X"22",X"00",X"00",
		X"E6",X"66",X"EE",X"00",X"E6",X"5E",X"2E",X"00",X"E6",X"5E",X"7E",X"00",X"22",X"EE",X"6E",X"00",
		X"2E",X"E6",X"EE",X"00",X"EE",X"22",X"06",X"00",X"00",X"22",X"00",X"00",X"00",X"2E",X"00",X"00",
		X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0F",X"EE",X"00",X"00",
		X"0E",X"ED",X"0E",X"00",X"0E",X"ED",X"ED",X"00",X"0E",X"ED",X"EE",X"00",X"EE",X"CE",X"CE",X"00",
		X"CF",X"CC",X"CC",X"00",X"CE",X"CC",X"CC",X"00",X"CE",X"CC",X"BB",X"00",X"BB",X"BB",X"EE",X"00",
		X"EE",X"EE",X"00",X"00",X"0E",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",
		X"0E",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"0E",X"00",X"00",X"0E",X"ED",X"00",X"00",
		X"0F",X"DD",X"00",X"00",X"0E",X"DD",X"00",X"00",X"EE",X"DD",X"00",X"00",X"CE",X"CC",X"0E",X"00",
		X"CE",X"CC",X"ED",X"00",X"EB",X"CC",X"DD",X"00",X"0E",X"BB",X"CD",X"00",X"0F",X"EE",X"CC",X"00",
		X"0E",X"E0",X"CC",X"00",X"00",X"E0",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"EC",X"00",
		X"0E",X"00",X"EC",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"0E",X"00",X"00",X"CC",X"EE",X"00",X"00",
		X"CC",X"ED",X"00",X"00",X"EC",X"DD",X"00",X"00",X"EB",X"ED",X"00",X"00",X"EE",X"CE",X"E0",X"00",
		X"0E",X"CC",X"CE",X"00",X"00",X"CC",X"CC",X"00",X"00",X"EE",X"CC",X"00",X"00",X"DE",X"CC",X"00",
		X"0F",X"DD",X"CC",X"00",X"00",X"DD",X"BE",X"00",X"00",X"DD",X"EE",X"00",X"00",X"DD",X"EC",X"00",
		X"00",X"DE",X"EC",X"00",X"00",X"E0",X"EC",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"0E",X"EE",X"00",X"00",
		X"EC",X"DD",X"00",X"00",X"CC",X"DD",X"00",X"00",X"CC",X"CD",X"0E",X"00",X"EB",X"CC",X"EE",X"00",
		X"0E",X"CC",X"ED",X"00",X"0F",X"CC",X"DD",X"00",X"0E",X"BE",X"DD",X"00",X"0E",X"EE",X"EE",X"00",
		X"F0",X"DD",X"CC",X"00",X"00",X"DD",X"CC",X"00",X"00",X"DE",X"CC",X"00",X"00",X"E0",X"CC",X"00",
		X"00",X"00",X"EC",X"00",X"00",X"00",X"EC",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"EE",X"E0",X"00",X"00",X"EC",X"CE",X"00",X"00",X"CC",X"CC",X"00",X"00",
		X"EC",X"CD",X"00",X"00",X"EB",X"CD",X"00",X"00",X"0E",X"CE",X"00",X"00",X"00",X"CC",X"EE",X"00",
		X"00",X"CC",X"DD",X"00",X"0E",X"CC",X"DD",X"00",X"F0",X"EE",X"DD",X"00",X"00",X"DE",X"ED",X"00",
		X"00",X"DB",X"CC",X"00",X"00",X"DE",X"CC",X"00",X"00",X"E0",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"00",X"00",X"00",X"CE",X"E0",X"00",X"00",X"CC",X"CE",X"00",X"00",X"EC",X"CD",X"00",X"00",
		X"EC",X"CD",X"00",X"00",X"0E",X"CE",X"00",X"00",X"0E",X"CE",X"00",X"00",X"00",X"CC",X"0E",X"00",
		X"00",X"CC",X"ED",X"00",X"0F",X"CC",X"ED",X"00",X"0F",X"E2",X"DD",X"00",X"00",X"DE",X"DD",X"00",
		X"00",X"DE",X"ED",X"00",X"00",X"DD",X"CE",X"00",X"00",X"DD",X"CC",X"00",X"00",X"DE",X"CC",X"00",
		X"00",X"EE",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0E",X"EE",X"E0",X"00",X"0E",X"CE",X"E0",X"00",X"0E",X"CC",X"E0",X"00",
		X"00",X"CE",X"E0",X"00",X"00",X"CD",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"CE",X"00",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"EC",X"EE",X"00",X"00",X"D2",X"EE",X"00",X"00",X"DE",X"DD",X"00",
		X"00",X"DE",X"ED",X"00",X"00",X"DD",X"CE",X"00",X"00",X"DD",X"CC",X"00",X"00",X"DD",X"CC",X"00",
		X"00",X"EE",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",
		X"EE",X"00",X"00",X"00",X"EC",X"E0",X"00",X"00",X"EB",X"CE",X"E0",X"00",X"EE",X"CC",X"E0",X"00",
		X"0E",X"CE",X"E0",X"00",X"00",X"CE",X"E0",X"00",X"00",X"ED",X"00",X"00",X"0E",X"CE",X"00",X"00",
		X"0E",X"CC",X"00",X"00",X"F0",X"CC",X"EE",X"00",X"00",X"EE",X"DD",X"00",X"00",X"EB",X"DD",X"00",
		X"00",X"EE",X"DD",X"00",X"00",X"DD",X"ED",X"00",X"00",X"DD",X"CE",X"00",X"00",X"DE",X"CC",X"00",
		X"00",X"E0",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CE",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",
		X"0E",X"EE",X"00",X"00",X"0E",X"CC",X"00",X"00",X"00",X"CC",X"E0",X"00",X"00",X"EC",X"DE",X"00",
		X"00",X"CC",X"DE",X"00",X"00",X"CE",X"DE",X"00",X"0F",X"CE",X"E0",X"00",X"00",X"CE",X"00",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"EC",X"00",X"00",X"00",X"E2",X"0E",X"00",X"00",X"EF",X"ED",X"00",
		X"00",X"DE",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"EE",X"DD",X"00",X"00",X"00",X"DD",X"00",
		X"00",X"00",X"EC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CE",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"E0",X"00",X"00",X"0E",X"00",X"00",X"00",
		X"0E",X"EE",X"00",X"00",X"0E",X"CC",X"00",X"00",X"00",X"CC",X"E0",X"00",X"00",X"EC",X"DE",X"00",
		X"00",X"CC",X"DE",X"00",X"0F",X"CE",X"DE",X"00",X"00",X"CE",X"DE",X"00",X"00",X"CC",X"E0",X"00",
		X"00",X"CE",X"00",X"00",X"00",X"BE",X"00",X"00",X"00",X"E2",X"00",X"00",X"00",X"EF",X"E0",X"00",
		X"00",X"EE",X"DE",X"00",X"00",X"DE",X"DD",X"00",X"00",X"EE",X"DD",X"00",X"00",X"00",X"DD",X"00",
		X"00",X"00",X"DE",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CE",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"EC",X"E0",X"00",X"00",X"CE",X"DE",X"00",
		X"00",X"CC",X"DE",X"00",X"0E",X"CC",X"DE",X"00",X"00",X"CE",X"DE",X"00",X"00",X"CE",X"E0",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"EC",X"00",X"00",X"00",X"BE",X"00",X"00",X"00",X"E2",X"00",X"00",
		X"00",X"DE",X"E0",X"00",X"00",X"EE",X"DE",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",
		X"00",X"00",X"DE",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"FE",X"00",X"00",X"00",X"E0",X"00",X"00",
		X"00",X"CE",X"00",X"00",X"00",X"EC",X"00",X"00",X"00",X"CE",X"EE",X"00",X"00",X"CC",X"DE",X"00",
		X"00",X"CC",X"DD",X"00",X"00",X"CC",X"DD",X"00",X"00",X"CC",X"DE",X"00",X"00",X"CC",X"E0",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E2",X"00",X"00",X"00",X"E2",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"EE",X"E0",X"00",X"00",X"E0",X"DE",X"00",X"00",X"00",X"DE",X"00",
		X"00",X"00",X"DE",X"00",X"00",X"0E",X"E0",X"00",X"00",X"0E",X"CE",X"00",X"00",X"0E",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"CE",X"00",X"00",X"00",X"EC",X"00",X"00",X"0F",X"CE",X"00",X"00",X"0F",X"CE",X"E0",X"00",
		X"00",X"CC",X"DE",X"00",X"00",X"CC",X"DE",X"00",X"00",X"CE",X"DD",X"00",X"00",X"CE",X"DE",X"00",
		X"00",X"CE",X"EE",X"00",X"00",X"EC",X"E0",X"00",X"00",X"2E",X"00",X"00",X"00",X"2E",X"00",X"00",
		X"00",X"EB",X"00",X"00",X"00",X"EB",X"00",X"00",X"00",X"0E",X"E0",X"00",X"00",X"00",X"DE",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"EC",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"CF",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"CC",X"EE",X"00",X"00",X"CC",X"DE",X"00",X"00",X"CE",X"DD",X"00",
		X"00",X"CC",X"DD",X"00",X"00",X"EC",X"DE",X"00",X"00",X"2E",X"E0",X"00",X"00",X"2E",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EB",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"EC",X"00",X"00",X"00",X"CC",X"00",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"CE",X"00",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"EF",X"00",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"EE",X"00",X"00",X"CC",X"DD",X"00",
		X"00",X"CC",X"DD",X"00",X"00",X"EC",X"DD",X"00",X"00",X"EC",X"DE",X"00",X"00",X"EC",X"E0",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"EC",X"00",X"00",X"00",X"BC",X"00",X"00",X"00",X"EC",X"00",X"00",
		X"00",X"EB",X"00",X"00",X"00",X"EC",X"00",X"00",X"00",X"EC",X"00",X"00",X"00",X"CC",X"00",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"EC",X"00",X"00",
		X"00",X"BC",X"00",X"00",X"00",X"BC",X"00",X"00",X"00",X"BC",X"00",X"00",X"00",X"E2",X"00",X"00",
		X"00",X"BC",X"00",X"00",X"00",X"BC",X"00",X"00",X"00",X"BC",X"00",X"00",X"00",X"BC",X"00",X"00",
		X"00",X"BC",X"00",X"00",X"00",X"BC",X"00",X"00",X"00",X"BC",X"00",X"00",X"00",X"EC",X"00",X"00",
		X"00",X"FE",X"00",X"00",X"00",X"2E",X"00",X"00",X"00",X"2E",X"00",X"00",X"00",X"FE",X"00",X"00",
		X"00",X"EC",X"00",X"00",X"00",X"BC",X"00",X"00",X"00",X"BC",X"00",X"00",X"00",X"EC",X"00",X"00",
		X"00",X"EC",X"00",X"00",X"00",X"EC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"E2",X"EE",X"00",X"EE",X"22",X"2E",X"00",X"E3",X"22",X"22",X"00",X"EE",X"22",X"22",X"00",
		X"0E",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"0E",X"22",X"2E",X"E0",X"0E",X"23",X"22",X"E0",
		X"0E",X"2E",X"22",X"00",X"EE",X"2E",X"22",X"00",X"E2",X"EE",X"22",X"00",X"33",X"EE",X"22",X"00",
		X"EE",X"22",X"22",X"00",X"EE",X"22",X"22",X"EE",X"E2",X"22",X"22",X"3E",X"E2",X"22",X"22",X"3E",
		X"EE",X"22",X"22",X"EE",X"0E",X"22",X"32",X"00",X"0E",X"22",X"32",X"00",X"0E",X"22",X"EE",X"00",
		X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"0E",X"22",X"22",X"00",X"70",X"07",X"77",X"00",
		X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"EF",X"00",X"00",
		X"00",X"FF",X"E0",X"00",X"00",X"FF",X"FE",X"00",X"00",X"FF",X"5F",X"00",X"00",X"FF",X"FF",X"00",
		X"00",X"FF",X"F5",X"00",X"00",X"E5",X"55",X"00",X"00",X"0E",X"55",X"00",X"00",X"0E",X"55",X"00",
		X"00",X"0E",X"55",X"00",X"00",X"0E",X"55",X"00",X"00",X"60",X"5E",X"00",X"00",X"00",X"5E",X"00",
		X"E0",X"00",X"EF",X"00",X"E4",X"00",X"FF",X"00",X"E5",X"E0",X"EF",X"00",X"E5",X"E0",X"0E",X"00",
		X"5E",X"E0",X"00",X"00",X"55",X"E0",X"00",X"00",X"E5",X"E0",X"00",X"00",X"0E",X"EE",X"00",X"00",
		X"E5",X"E4",X"60",X"00",X"55",X"5E",X"00",X"00",X"55",X"5E",X"00",X"00",X"55",X"5E",X"00",X"00",
		X"E5",X"E0",X"00",X"00",X"E5",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"EF",X"00",X"00",
		X"00",X"FF",X"E0",X"00",X"00",X"FF",X"FE",X"00",X"00",X"FF",X"CF",X"00",X"00",X"FF",X"FF",X"00",
		X"00",X"FF",X"FC",X"00",X"00",X"EC",X"CC",X"00",X"00",X"0E",X"CC",X"00",X"00",X"0E",X"CC",X"00",
		X"00",X"0E",X"CC",X"00",X"00",X"0E",X"CC",X"00",X"00",X"60",X"CE",X"00",X"00",X"00",X"CE",X"00",
		X"E0",X"00",X"EF",X"00",X"E4",X"00",X"FF",X"00",X"EC",X"E0",X"EF",X"00",X"EC",X"E0",X"0E",X"00",
		X"CE",X"E0",X"00",X"00",X"CB",X"E0",X"00",X"00",X"EC",X"E0",X"00",X"00",X"0E",X"EE",X"00",X"00",
		X"EC",X"E4",X"60",X"00",X"CC",X"CE",X"00",X"00",X"CC",X"CE",X"00",X"00",X"CC",X"CE",X"00",X"00",
		X"EC",X"E0",X"00",X"00",X"EC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"00",X"00",
		X"55",X"55",X"E0",X"00",X"55",X"55",X"5E",X"00",X"5B",X"BB",X"BB",X"00",X"5B",X"BB",X"BB",X"00",
		X"5B",X"BB",X"BB",X"00",X"E5",X"BB",X"BB",X"00",X"E5",X"BB",X"BB",X"00",X"E5",X"BB",X"BB",X"00",
		X"E5",X"BB",X"BB",X"00",X"E5",X"BB",X"BB",X"70",X"E5",X"BB",X"BB",X"07",X"75",X"BB",X"BB",X"00",
		X"E0",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"0F",X"00",X"0F",X"30",X"30",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"30",
		X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"30",
		X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"30",
		X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"30",
		X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"F0",X"03",X"03",X"00",X"00",X"F0",X"F0",X"00",
		X"00",X"30",X"00",X"00",X"03",X"22",X"00",X"00",X"21",X"00",X"00",X"00",X"20",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"5E",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"E0",X"00",X"00",
		X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"BE",X"00",X"00",X"10",X"BE",X"00",X"00",
		X"11",X"BE",X"00",X"00",X"31",X"BE",X"00",X"00",X"13",X"EF",X"00",X"00",X"31",X"5F",X"00",X"00",
		X"E1",X"5E",X"00",X"00",X"66",X"E5",X"00",X"00",X"66",X"E5",X"00",X"00",X"E6",X"E5",X"00",X"00",
		X"0E",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"EF",X"00",X"00",X"00",X"E5",X"00",X"00",
		X"00",X"30",X"00",X"00",X"03",X"22",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"CE",X"00",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CE",X"00",X"00",X"00",X"E0",X"00",X"00",
		X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"BE",X"00",X"00",X"00",X"BE",X"00",X"00",
		X"00",X"BE",X"00",X"00",X"30",X"BE",X"00",X"00",X"13",X"EF",X"00",X"00",X"33",X"CF",X"00",X"00",
		X"E3",X"CE",X"00",X"00",X"DD",X"EC",X"00",X"00",X"DD",X"EC",X"00",X"00",X"ED",X"EC",X"00",X"00",
		X"0E",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"EF",X"00",X"00",X"00",X"EC",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
