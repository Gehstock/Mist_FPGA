library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity bg1_rom is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of bg1_rom is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"0F",X"1E",X"3C",X"78",X"F0",X"E1",X"C3",X"87",X"F0",X"E1",X"C3",X"87",X"0F",X"1E",X"3C",X"78",
		X"0F",X"1E",X"3C",X"78",X"F0",X"E1",X"C3",X"87",X"38",X"6C",X"C6",X"83",X"83",X"C6",X"6C",X"38",
		X"C7",X"93",X"39",X"7C",X"7C",X"39",X"93",X"C7",X"38",X"6C",X"C6",X"83",X"83",X"C6",X"6C",X"38",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"3C",X"78",X"F0",X"F0",X"F0",X"78",X"3C",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C0",X"C0",X"C0",X"CC",X"CC",X"0C",X"0C",X"0C",
		X"3F",X"3F",X"3F",X"33",X"33",X"F3",X"F3",X"F3",X"C0",X"C0",X"C0",X"CC",X"CC",X"0C",X"0C",X"0C",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"F8",X"88",X"F8",X"00",X"F8",X"88",X"F8",
		X"00",X"48",X"F8",X"08",X"00",X"F8",X"88",X"F8",X"00",X"48",X"F8",X"08",X"00",X"E8",X"A8",X"B8",
		X"00",X"B8",X"A8",X"E8",X"00",X"F8",X"88",X"F8",X"00",X"B8",X"A8",X"E8",X"00",X"E8",X"A8",X"B8",
		X"00",X"88",X"A8",X"F8",X"00",X"F8",X"88",X"F8",X"00",X"88",X"A8",X"F8",X"00",X"E8",X"A8",X"B8",
		X"00",X"F0",X"10",X"F8",X"00",X"F8",X"88",X"F8",X"00",X"F0",X"10",X"F8",X"00",X"E8",X"A8",X"B8",
		X"00",X"E8",X"A8",X"B8",X"00",X"F8",X"88",X"F8",X"00",X"F8",X"A8",X"B8",X"00",X"F8",X"88",X"F8",
		X"00",X"80",X"80",X"F8",X"00",X"F8",X"88",X"F8",X"00",X"F8",X"A8",X"F8",X"00",X"F8",X"88",X"F8",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"F7",X"F7",X"F7",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F3",X"F3",X"F3",X"F1",X"E1",X"E1",X"E1",X"C1",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C3",X"C3",X"C3",X"C3",X"C3",X"C3",X"C3",X"C1",
		X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"7F",X"3F",X"E0",X"F0",X"F8",X"FC",X"FC",X"FC",X"FC",X"FE",
		X"3F",X"3F",X"3F",X"1F",X"1F",X"1F",X"1F",X"8F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"CF",X"C7",X"E7",X"E3",X"E3",X"F3",X"F3",X"F1",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"C0",X"E0",
		X"3C",X"FE",X"7F",X"7F",X"3F",X"3F",X"3F",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"1E",X"1E",X"1F",X"0F",X"0F",X"06",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FE",X"FC",X"FC",X"FC",X"FE",X"64",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"80",X"C0",X"40",X"00",X"00",X"00",X"FE",X"FF",X"FF",X"F7",X"F0",X"E0",X"F8",X"FE",
		X"00",X"00",X"C0",X"F0",X"E0",X"E0",X"E0",X"C0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FC",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"3F",X"3F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"E7",X"C2",X"82",X"80",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"E0",X"C0",X"C0",X"80",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"0F",X"1F",X"3F",X"3F",X"3F",X"7F",X"7F",
		X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"5F",X"5F",
		X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"F1",X"F8",X"FC",X"FC",
		X"7F",X"FF",X"FF",X"7F",X"27",X"23",X"01",X"01",X"80",X"8F",X"38",X"F0",X"F0",X"F0",X"F8",X"F8",
		X"6F",X"6F",X"EF",X"EF",X"EF",X"EF",X"EF",X"CF",X"00",X"00",X"00",X"00",X"00",X"81",X"E3",X"FF",
		X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"03",X"0F",X"01",X"00",X"00",X"00",X"01",X"63",
		X"F0",X"F0",X"C0",X"00",X"00",X"00",X"00",X"00",X"8F",X"0F",X"0F",X"07",X"02",X"00",X"00",X"00",
		X"FF",X"F8",X"F0",X"F0",X"E0",X"C0",X"80",X"80",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"0F",X"01",X"00",X"01",X"07",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"73",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"E0",X"F8",X"FC",X"FE",
		X"00",X"00",X"01",X"83",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"03",X"07",X"07",X"0F",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"07",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FC",X"F8",X"F0",X"E0",X"E0",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"83",X"31",X"F0",X"90",X"10",X"00",X"00",X"FF",X"FF",X"FE",X"F8",X"F3",X"EE",X"EC",X"CC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",
		X"87",X"00",X"00",X"00",X"06",X"0C",X"08",X"18",X"FF",X"FF",X"FF",X"FE",X"FE",X"FC",X"FC",X"F8",
		X"03",X"13",X"30",X"E0",X"E0",X"C0",X"80",X"00",X"18",X"1C",X"1E",X"0F",X"0F",X"07",X"03",X"00",
		X"F8",X"F8",X"F0",X"F0",X"F0",X"E0",X"E0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"F0",X"F0",
		X"00",X"00",X"00",X"0F",X"3F",X"7F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"80",X"C0",X"FF",X"FF",
		X"F8",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"00",X"FF",X"FF",X"FF",X"FF",X"7F",X"03",X"00",X"F0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"87",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FE",X"F8",X"E3",X"CF",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"FF",X"FF",X"FF",X"7F",
		X"FF",X"0F",X"E0",X"FE",X"7F",X"1F",X"03",X"00",X"FF",X"EF",X"E7",X"E1",X"E0",X"F0",X"F8",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F1",X"E7",X"CF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"F8",X"F8",
		X"3F",X"9F",X"CF",X"07",X"13",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"FB",X"FF",
		X"FF",X"CF",X"1F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FD",X"F9",X"F7",X"FC",X"F1",X"C7",X"7F",X"3F",
		X"0F",X"E0",X"FF",X"FF",X"3F",X"03",X"C0",X"F0",X"30",X"9F",X"C7",X"F0",X"FC",X"FE",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"FC",X"F8",X"F8",X"E0",X"80",X"00",X"63",X"C9",X"C9",X"88",X"8C",X"86",X"86",X"86",
		X"F0",X"E0",X"C1",X"81",X"83",X"83",X"87",X"8F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"7C",X"70",X"F8",X"F0",X"F8",X"FC",X"FE",
		X"86",X"83",X"83",X"81",X"C1",X"C0",X"E1",X"F0",X"CF",X"EF",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"F0",X"F0",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FE",X"FC",X"FC",X"FC",X"78",X"30",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"1E",X"00",X"7F",X"FF",X"23",X"01",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"1F",X"C7",X"F3",X"F9",X"7D",X"7D",
		X"7D",X"7D",X"FD",X"FD",X"F9",X"F9",X"F9",X"F1",X"E1",X"03",X"03",X"03",X"02",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"80",X"01",X"01",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FE",X"F8",X"F0",X"E0",X"E0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"00",X"00",X"00",X"00",X"C0",X"C3",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"07",X"0F",X"1F",X"1F",X"1F",X"1F",X"0F",X"0F",
		X"0F",X"1F",X"BF",X"BF",X"BF",X"BF",X"BF",X"80",X"80",X"B8",X"B8",X"B8",X"B8",X"B8",X"38",X"38",
		X"78",X"F8",X"F8",X"F8",X"F8",X"F8",X"78",X"38",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"F0",X"D8",X"CC",X"FE",X"FE",X"F2",X"00",X"00",X"03",X"03",X"03",X"01",X"00",X"00",
		X"F6",X"FC",X"FC",X"C8",X"D8",X"F0",X"00",X"00",X"00",X"01",X"03",X"03",X"03",X"03",X"00",X"00",
		X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"02",X"08",X"00",X"00",X"08",
		X"88",X"20",X"00",X"48",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"1C",X"00",X"00",X"00",X"00",X"04",X"0E",X"1F",X"1F",
		X"3C",X"48",X"C4",X"3E",X"0E",X"04",X"00",X"00",X"1F",X"1F",X"0E",X"04",X"00",X"00",X"00",X"00",
		X"00",X"00",X"40",X"E0",X"F0",X"F2",X"F6",X"BE",X"00",X"00",X"00",X"00",X"03",X"07",X"07",X"03",
		X"3E",X"36",X"72",X"F0",X"E0",X"40",X"00",X"00",X"03",X"06",X"04",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"40",X"60",X"70",X"38",X"38",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"38",X"38",X"38",X"70",X"60",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"D8",X"4C",X"66",X"26",X"32",X"32",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"32",X"32",X"26",X"66",X"4C",X"D8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"22",X"22",X"EE",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"0E",
		X"00",X"22",X"22",X"EE",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"0E",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FA",X"FA",X"FA",X"FA",X"7A",X"00",X"00",X"00",X"07",X"03",X"01",X"00",X"1A",
		X"3A",X"9A",X"40",X"A0",X"D0",X"00",X"00",X"00",X"1D",X"1E",X"1F",X"1F",X"1F",X"00",X"00",X"00",
		X"00",X"3C",X"20",X"1C",X"20",X"1C",X"00",X"BC",X"00",X"44",X"6C",X"68",X"6E",X"6C",X"68",X"6E",
		X"00",X"FC",X"00",X"FC",X"18",X"24",X"24",X"00",X"6E",X"68",X"6E",X"6C",X"68",X"6C",X"44",X"00",
		X"00",X"00",X"F8",X"1C",X"0C",X"0E",X"1E",X"FE",X"00",X"00",X"03",X"07",X"0E",X"1E",X"1F",X"1F",
		X"7E",X"3E",X"3E",X"3C",X"70",X"E0",X"00",X"00",X"1C",X"18",X"18",X"08",X"0C",X"07",X"00",X"00",
		X"00",X"00",X"00",X"60",X"B0",X"D8",X"D8",X"D8",X"00",X"00",X"00",X"07",X"0F",X"1F",X"1F",X"19",
		X"D8",X"D8",X"D8",X"B0",X"60",X"00",X"00",X"00",X"19",X"1F",X"1F",X"0F",X"07",X"00",X"00",X"00",
		X"00",X"00",X"00",X"E0",X"F1",X"F9",X"FF",X"F9",X"00",X"00",X"00",X"07",X"07",X"07",X"07",X"07",
		X"F1",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"1F",X"1E",X"0C",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"60",X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"60",X"60",X"60",X"00",X"00",X"00",X"00",X"00",X"E7",X"E7",X"00",
		X"00",X"00",X"00",X"00",X"00",X"79",X"79",X"00",X"00",X"00",X"00",X"00",X"00",X"9E",X"9E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"06",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"06",
		X"00",X"00",X"00",X"00",X"00",X"07",X"07",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"60",
		X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"00",X"00",X"60",X"60",X"60",X"60",X"60",X"60",X"60",
		X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"06",X"06",X"06",X"06",X"06",X"06",X"06",
		X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"00",X"60",X"60",X"60",X"00",X"00",X"60",X"60",X"60",
		X"00",X"60",X"60",X"60",X"60",X"00",X"00",X"60",X"60",X"00",X"00",X"60",X"60",X"60",X"60",X"00",
		X"06",X"06",X"06",X"00",X"00",X"06",X"06",X"06",X"06",X"00",X"00",X"06",X"06",X"06",X"06",X"00",
		X"00",X"06",X"06",X"06",X"06",X"00",X"00",X"06",X"60",X"80",X"80",X"00",X"00",X"00",X"00",X"00",
		X"60",X"60",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"E7",X"E7",X"00",X"00",X"00",X"00",X"00",X"00",X"9E",X"9E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"79",X"79",X"00",X"00",X"00",X"00",X"00",X"06",X"01",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"06",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"F0",X"F8",X"3C",X"1E",X"07",
		X"00",X"00",X"00",X"00",X"00",X"03",X"0F",X"3F",X"80",X"C0",X"60",X"30",X"08",X"04",X"F0",X"FF",
		X"03",X"01",X"00",X"00",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"F0",X"C0",X"00",
		X"FF",X"F0",X"04",X"08",X"30",X"60",X"C0",X"80",X"FF",X"FF",X"FF",X"F0",X"00",X"00",X"01",X"03",
		X"00",X"C0",X"F0",X"FC",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"1E",X"3C",X"F8",X"F0",X"E0",X"C0",X"80",X"3F",X"0F",X"03",X"00",X"00",X"00",X"00",X"00",
		X"01",X"03",X"07",X"0F",X"1F",X"3C",X"70",X"C0",X"00",X"C0",X"F0",X"FC",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"3F",X"0F",X"03",X"03",X"0F",X"3F",X"FF",X"FF",X"7F",X"3F",X"1F",X"0F",X"07",X"03",X"01",
		X"01",X"03",X"07",X"0F",X"1F",X"3F",X"7F",X"FF",X"FF",X"3F",X"0F",X"03",X"03",X"0F",X"3F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FC",X"F0",X"C0",X"00",X"C0",X"70",X"3C",X"1F",X"0F",X"07",X"03",X"01",
		X"00",X"00",X"00",X"00",X"1C",X"3C",X"7F",X"FF",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"E0",
		X"00",X"00",X"00",X"00",X"03",X"0F",X"0F",X"07",X"00",X"00",X"00",X"00",X"6C",X"FE",X"FC",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"FD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"1F",X"1E",X"7F",X"FF",X"FF",X"FF",X"7E",X"3C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"7C",X"7F",X"7F",X"7E",X"70",X"38",X"18",X"C6",X"0F",X"0F",X"8F",X"E6",X"F0",X"38",X"18",
		X"03",X"80",X"C0",X"FF",X"FF",X"78",X"18",X"78",X"FF",X"7F",X"FF",X"FF",X"7E",X"7C",X"F0",X"FC",
		X"FC",X"FC",X"F8",X"F1",X"E0",X"00",X"00",X"00",X"CF",X"CF",X"C7",X"C3",X"81",X"00",X"00",X"00",
		X"3F",X"3F",X"3F",X"3F",X"1F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F8",X"FC",X"FC",
		X"00",X"00",X"60",X"E0",X"80",X"01",X"33",X"FB",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"18",X"18",X"18",X"38",X"F0",X"E0",X"80",
		X"D8",X"88",X"D8",X"78",X"18",X"78",X"FF",X"FF",X"FE",X"FF",X"FE",X"FC",X"F0",X"7C",X"3E",X"0F",
		X"00",X"00",X"80",X"C0",X"E0",X"E0",X"F0",X"F0",X"00",X"1E",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"03",X"FC",X"70",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"EE",X"CC",X"00",X"00",X"00",X"00",X"1F",X"1F",X"3F",X"3F",X"1F",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"E0",X"C0",X"C0",X"80",X"00",X"1F",X"1F",X"1F",X"83",X"8F",X"DF",X"DF",X"90",
		X"F0",X"F0",X"E7",X"EF",X"DF",X"81",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"1E",X"00",
		X"03",X"03",X"01",X"01",X"00",X"38",X"7C",X"7E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"20",X"60",X"E0",X"E0",X"E0",X"E0",X"00",X"00",X"00",X"78",X"FC",X"FE",X"FE",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"F8",X"F8",
		X"FE",X"FE",X"FE",X"FC",X"78",X"00",X"00",X"01",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"60",X"20",X"00",X"40",X"FC",X"FC",X"F8",X"C0",X"FE",X"7C",X"38",X"00",X"10",X"1F",X"1F",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"F8",X"F8",X"F8",X"70",X"0E",X"07",X"21",X"E1",
		X"E1",X"F1",X"F8",X"F8",X"F8",X"78",X"30",X"00",X"01",X"03",X"01",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"E0",X"60",X"00",X"00",X"00",X"00",X"00",X"3F",X"3F",X"3F",X"1B",X"00",X"00",X"00",X"00",
		X"F0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"7E",X"00",X"00",X"00",X"00",
		X"1F",X"3F",X"3F",X"3F",X"3E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"38",X"78",X"F8",X"F8",X"F8",X"F8",X"F8",X"78",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"FC",
		X"00",X"00",X"00",X"00",X"78",X"FC",X"FC",X"1F",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",
		X"38",X"38",X"B8",X"B8",X"B8",X"B8",X"B8",X"80",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"0F",X"1F",X"3F",X"FF",X"FF",X"DF",X"0F",X"0E",X"0C",X"0C",X"0E",X"07",X"07",X"03",X"00",
		X"80",X"BF",X"BF",X"BF",X"BF",X"BF",X"1F",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",
		X"0F",X"DF",X"FF",X"FF",X"3F",X"1F",X"0F",X"0F",X"00",X"03",X"07",X"07",X"0E",X"0C",X"0C",X"0E",
		X"0F",X"0F",X"1F",X"1F",X"1F",X"1F",X"0F",X"07",X"FC",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"FE",X"FC",X"78",X"00",X"00",X"00",X"00",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"E3",
		X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"61",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"F8",X"F8",X"FE",X"FF",X"FF",X"FF",X"7F",X"CF",X"DD",X"F8",X"F8",X"FD",X"7F",X"7F",X"CF",
		X"E7",X"EF",X"FF",X"FF",X"FC",X"F8",X"F8",X"FC",X"01",X"07",X"0F",X"1F",X"3F",X"7F",X"FF",X"FF",
		X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"E7",X"C3",X"CE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FC",X"FC",X"3F",X"1F",X"1F",X"1F",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"7C",X"7E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"F9",X"FC",X"EC",X"60",
		X"1F",X"FF",X"FF",X"FF",X"FF",X"7E",X"00",X"00",X"7F",X"3F",X"1F",X"07",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"60",X"70",X"38",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"07",X"FF",X"FF",X"7F",X"1F",X"0F",X"0F",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"02",X"02",X"01",X"00",X"03",
		X"3F",X"FF",X"3F",X"0F",X"1F",X"3F",X"7F",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"F8",
		X"80",X"80",X"00",X"00",X"00",X"80",X"E0",X"FB",X"0F",X"38",X"61",X"42",X"C2",X"C1",X"81",X"00",
		X"DC",X"18",X"30",X"60",X"80",X"00",X"00",X"00",X"F1",X"C3",X"00",X"00",X"00",X"00",X"00",X"00",
		X"79",X"3D",X"1D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"F0",X"FC",X"7E",X"3E",X"0F",X"07",X"83",X"00",X"00",X"06",X"0C",X"00",X"00",X"03",X"07",
		X"00",X"00",X"00",X"00",X"F0",X"F8",X"FC",X"FC",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",
		X"00",X"18",X"3C",X"3C",X"18",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"07",X"07",X"47",X"E7",
		X"47",X"E3",X"40",X"00",X"18",X"18",X"00",X"80",X"FC",X"FC",X"FC",X"F6",X"F2",X"03",X"81",X"C1",
		X"03",X"03",X"03",X"01",X"80",X"C0",X"C7",X"9F",X"00",X"18",X"18",X"00",X"01",X"33",X"33",X"01",
		X"43",X"03",X"03",X"03",X"01",X"01",X"00",X"00",X"86",X"CF",X"4F",X"66",X"20",X"20",X"00",X"00",
		X"F0",X"F2",X"E7",X"F2",X"F8",X"B8",X"90",X"D3",X"7F",X"FF",X"FF",X"FF",X"FF",X"F7",X"E3",X"80",
		X"00",X"00",X"30",X"39",X"39",X"11",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"00",X"00",X"C0",X"C0",X"C0",X"80",X"D7",X"D7",X"43",X"00",X"01",X"07",X"3F",X"32",
		X"E3",X"F7",X"7C",X"18",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F8",X"F8",X"F8",X"FC",X"FC",X"FE",X"7E",X"CF",X"DD",X"F8",X"F8",X"FD",X"7F",X"7F",X"CF",
		X"3F",X"7F",X"FF",X"FF",X"F7",X"F0",X"E0",X"C0",X"CE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"F8",X"F8",X"C0",X"E0",X"E0",X"00",X"80",X"FF",X"FF",X"BF",X"3F",X"1F",X"0F",X"07",X"03",
		X"00",X"C0",X"F0",X"FC",X"FC",X"00",X"00",X"80",X"0E",X"1F",X"1F",X"03",X"31",X"60",X"03",X"07",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"F0",X"10",X"10",X"10",X"10",
		X"00",X"00",X"00",X"FF",X"10",X"10",X"10",X"10",X"00",X"00",X"00",X"1F",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"F0",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"FF",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"1F",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"F0",X"00",X"00",X"00",X"00",
		X"10",X"10",X"10",X"FF",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"1F",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
