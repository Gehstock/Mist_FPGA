library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ps01 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ps01 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"C3",X"C6",X"05",X"00",X"00",X"F5",X"C5",X"D5",X"E5",X"C3",X"A7",X"51",X"00",
		X"F5",X"C5",X"D5",X"E5",X"C3",X"40",X"00",X"00",X"C3",X"6E",X"0A",X"E5",X"FF",X"11",X"05",X"09",
		X"3A",X"03",X"23",X"67",X"C9",X"0C",X"49",X"01",X"C3",X"D8",X"02",X"AB",X"07",X"21",X"F0",X"20",
		X"C3",X"D6",X"04",X"2A",X"21",X"20",X"01",X"04",X"C3",X"2F",X"0B",X"06",X"57",X"00",X"00",X"43",
		X"21",X"00",X"23",X"35",X"23",X"34",X"CD",X"1B",X"04",X"DB",X"01",X"0F",X"DA",X"90",X"00",X"3A",
		X"09",X"23",X"A7",X"CA",X"6B",X"00",X"3A",X"0A",X"23",X"FE",X"18",X"D2",X"67",X"00",X"C6",X"01",
		X"27",X"32",X"0A",X"23",X"CD",X"8F",X"04",X"AF",X"32",X"09",X"23",X"3A",X"08",X"23",X"A7",X"CA",
		X"87",X"00",X"3A",X"0D",X"23",X"A7",X"C2",X"64",X"09",X"3A",X"0A",X"23",X"A7",X"C2",X"95",X"00",
		X"3A",X"0B",X"23",X"A7",X"C2",X"64",X"09",X"CD",X"A9",X"16",X"E1",X"D1",X"C1",X"F1",X"FB",X"C9",
		X"3E",X"01",X"C3",X"68",X"00",X"3A",X"4C",X"20",X"A7",X"C2",X"87",X"00",X"3E",X"01",X"32",X"4C",
		X"20",X"AF",X"32",X"0B",X"23",X"31",X"FF",X"23",X"FB",X"CD",X"D9",X"01",X"CD",X"A0",X"04",X"21",
		X"16",X"30",X"11",X"79",X"42",X"0E",X"04",X"CD",X"E6",X"02",X"D3",X"05",X"3A",X"0A",X"23",X"3D",
		X"D3",X"05",X"21",X"12",X"28",X"0E",X"14",X"C2",X"B9",X"01",X"11",X"12",X"05",X"CD",X"E6",X"02",
		X"DB",X"01",X"E6",X"04",X"CA",X"BC",X"00",X"06",X"99",X"AF",X"32",X"0C",X"23",X"3A",X"0A",X"23",
		X"80",X"27",X"32",X"0A",X"23",X"CD",X"8F",X"04",X"21",X"0D",X"23",X"34",X"21",X"00",X"00",X"22",
		X"18",X"23",X"22",X"1C",X"23",X"CD",X"15",X"02",X"CD",X"20",X"02",X"CD",X"2B",X"02",X"CD",X"A0",
		X"04",X"CD",X"6E",X"01",X"06",X"20",X"CD",X"2E",X"09",X"21",X"01",X"01",X"22",X"04",X"23",X"DB",
		X"02",X"07",X"DC",X"B1",X"4B",X"21",X"03",X"23",X"36",X"22",X"E5",X"CD",X"CB",X"07",X"E1",X"36",
		X"21",X"CD",X"CB",X"07",X"CD",X"7F",X"01",X"CD",X"DE",X"01",X"CD",X"92",X"0A",X"CD",X"86",X"08",
		X"CD",X"0C",X"15",X"CD",X"D4",X"01",X"21",X"37",X"20",X"AF",X"BE",X"C2",X"3B",X"14",X"E7",X"2E",
		X"4D",X"7E",X"FE",X"0A",X"CA",X"57",X"01",X"FE",X"0B",X"D2",X"33",X"15",X"CD",X"8C",X"01",X"CD",
		X"73",X"08",X"D3",X"05",X"C3",X"36",X"01",X"2E",X"49",X"AF",X"BE",X"C2",X"4C",X"01",X"34",X"2E",
		X"00",X"36",X"00",X"2E",X"13",X"36",X"00",X"21",X"E3",X"20",X"34",X"C3",X"4C",X"01",X"DB",X"02",
		X"E6",X"03",X"21",X"4F",X"21",X"F5",X"86",X"77",X"F1",X"21",X"4F",X"22",X"86",X"77",X"C9",X"3A",
		X"0C",X"23",X"A7",X"C0",X"21",X"01",X"2E",X"06",X"28",X"C3",X"CB",X"03",X"CD",X"AF",X"01",X"7E",
		X"A7",X"C8",X"06",X"50",X"CD",X"9F",X"03",X"B8",X"D8",X"CD",X"E4",X"08",X"34",X"CD",X"DE",X"01",
		X"CD",X"AF",X"01",X"36",X"00",X"21",X"4A",X"20",X"34",X"11",X"49",X"4E",X"C3",X"41",X"4E",X"21",
		X"04",X"23",X"3A",X"03",X"23",X"0F",X"D8",X"23",X"C9",X"11",X"FD",X"04",X"CD",X"E6",X"02",X"DB",
		X"01",X"0F",X"0F",X"DA",X"CD",X"01",X"0F",X"DA",X"D7",X"00",X"C3",X"BC",X"00",X"3E",X"01",X"06",
		X"98",X"C3",X"DA",X"00",X"3E",X"01",X"C3",X"DA",X"01",X"AF",X"32",X"08",X"23",X"C9",X"CD",X"E4",
		X"08",X"7E",X"3D",X"C8",X"4F",X"21",X"03",X"34",X"11",X"B7",X"42",X"C5",X"06",X"10",X"CD",X"DB",
		X"03",X"C1",X"0D",X"C2",X"E8",X"01",X"C9",X"C3",X"00",X"57",X"23",X"11",X"15",X"23",X"1A",X"BE",
		X"1B",X"2B",X"1A",X"CA",X"0A",X"02",X"D0",X"C3",X"0C",X"02",X"BE",X"D0",X"7E",X"12",X"13",X"23",
		X"7E",X"12",X"C3",X"9A",X"04",X"06",X"00",X"11",X"00",X"40",X"21",X"00",X"20",X"C3",X"BB",X"04",
		X"06",X"50",X"21",X"00",X"21",X"11",X"00",X"41",X"C3",X"BB",X"04",X"06",X"50",X"21",X"00",X"22",
		X"C3",X"25",X"02",X"7E",X"3D",X"21",X"03",X"34",X"CA",X"41",X"02",X"24",X"24",X"3D",X"C2",X"3B",
		X"02",X"06",X"10",X"CD",X"CB",X"03",X"C3",X"6E",X"03",X"21",X"07",X"28",X"11",X"54",X"02",X"0E",
		X"13",X"C3",X"54",X"03",X"06",X"00",X"0C",X"04",X"1B",X"0E",X"15",X"04",X"11",X"1B",X"0F",X"0B",
		X"00",X"18",X"04",X"11",X"26",X"1B",X"27",X"3A",X"03",X"23",X"0F",X"DA",X"77",X"02",X"06",X"20",
		X"21",X"07",X"23",X"70",X"C3",X"C6",X"02",X"06",X"00",X"C3",X"70",X"02",X"CD",X"F7",X"01",X"CD",
		X"15",X"02",X"CD",X"5A",X"15",X"CD",X"5F",X"15",X"21",X"03",X"23",X"11",X"53",X"41",X"06",X"05",
		X"CD",X"BB",X"04",X"21",X"00",X"00",X"22",X"0C",X"23",X"CD",X"F0",X"04",X"CD",X"77",X"02",X"CD",
		X"A0",X"04",X"21",X"13",X"2D",X"11",X"54",X"02",X"0E",X"0A",X"CD",X"54",X"03",X"CD",X"6E",X"03",
		X"C3",X"E0",X"05",X"CD",X"48",X"03",X"23",X"11",X"15",X"23",X"1A",X"BE",X"1B",X"2B",X"1A",X"CA",
		X"0A",X"02",X"D0",X"C3",X"0C",X"02",X"F3",X"78",X"D3",X"06",X"06",X"0A",X"0E",X"00",X"0D",X"C2",
		X"CE",X"02",X"05",X"C2",X"CC",X"02",X"FB",X"C9",X"4E",X"23",X"46",X"23",X"79",X"86",X"77",X"23",
		X"78",X"86",X"77",X"C9",X"0E",X"02",X"1A",X"D5",X"CD",X"F2",X"02",X"D1",X"13",X"0D",X"C2",X"E6",
		X"02",X"C9",X"CD",X"3F",X"05",X"06",X"05",X"D3",X"05",X"CD",X"DB",X"03",X"C5",X"AF",X"77",X"01",
		X"20",X"00",X"09",X"77",X"09",X"77",X"09",X"C1",X"C9",X"CD",X"48",X"03",X"3A",X"11",X"23",X"A7",
		X"C8",X"AF",X"32",X"11",X"23",X"E5",X"2A",X"12",X"23",X"EB",X"E1",X"7E",X"83",X"27",X"77",X"5F",
		X"23",X"7E",X"8A",X"27",X"77",X"57",X"23",X"7E",X"23",X"66",X"6F",X"7A",X"CD",X"30",X"03",X"7B",
		X"D5",X"F5",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"CD",X"43",X"03",X"F1",X"E6",X"0F",X"CD",X"43",
		X"03",X"D1",X"C9",X"C6",X"1C",X"C3",X"F2",X"02",X"3A",X"03",X"23",X"0F",X"21",X"18",X"23",X"D8",
		X"21",X"1C",X"23",X"C9",X"D5",X"1A",X"CD",X"F2",X"02",X"D1",X"3E",X"07",X"32",X"00",X"23",X"3A",
		X"00",X"23",X"3D",X"D3",X"05",X"C2",X"5F",X"03",X"13",X"0D",X"C2",X"54",X"03",X"C9",X"3E",X"40",
		X"C3",X"78",X"03",X"3E",X"80",X"C3",X"78",X"03",X"32",X"00",X"23",X"3A",X"00",X"23",X"A7",X"D3",
		X"05",X"C2",X"7B",X"03",X"C9",X"3E",X"20",X"C3",X"78",X"03",X"3E",X"05",X"C3",X"78",X"03",X"E5",
		X"D5",X"11",X"00",X"04",X"19",X"3E",X"1C",X"CD",X"F2",X"02",X"D1",X"E1",X"C3",X"2B",X"03",X"CD",
		X"48",X"03",X"7E",X"23",X"66",X"6F",X"29",X"29",X"29",X"29",X"7C",X"C9",X"F7",X"C5",X"E5",X"1A",
		X"D3",X"03",X"DB",X"03",X"AE",X"77",X"23",X"13",X"AF",X"D3",X"03",X"DB",X"03",X"AE",X"77",X"E1",
		X"01",X"20",X"00",X"09",X"C1",X"05",X"C2",X"AD",X"03",X"C9",X"F7",X"C5",X"E5",X"AF",X"77",X"E1",
		X"01",X"20",X"00",X"09",X"C1",X"05",X"C2",X"CB",X"03",X"C9",X"F7",X"C5",X"1A",X"77",X"13",X"01",
		X"20",X"00",X"09",X"C1",X"05",X"C2",X"DB",X"03",X"C9",X"F7",X"C5",X"E5",X"1A",X"D3",X"03",X"DB",
		X"03",X"77",X"23",X"13",X"AF",X"D3",X"03",X"DB",X"03",X"77",X"E1",X"01",X"20",X"00",X"09",X"C1",
		X"05",X"C2",X"EA",X"03",X"C9",X"3A",X"0D",X"23",X"A7",X"C8",X"DB",X"02",X"E6",X"04",X"DB",X"01",
		X"C8",X"3A",X"03",X"23",X"0F",X"DB",X"00",X"D0",X"DB",X"01",X"C9",X"DB",X"00",X"E6",X"04",X"C8",
		X"3A",X"4B",X"20",X"A7",X"C0",X"06",X"04",X"CD",X"56",X"09",X"31",X"FF",X"23",X"06",X"04",X"C5",
		X"CD",X"F0",X"04",X"C1",X"05",X"C2",X"2F",X"04",X"3E",X"01",X"32",X"4B",X"20",X"CD",X"D9",X"01",
		X"FB",X"11",X"80",X"41",X"21",X"16",X"30",X"0E",X"04",X"CD",X"54",X"03",X"CD",X"6E",X"03",X"C3",
		X"C6",X"05",X"0E",X"08",X"11",X"27",X"05",X"21",X"03",X"25",X"CD",X"E6",X"02",X"0E",X"08",X"21",
		X"02",X"25",X"CD",X"E6",X"02",X"0E",X"08",X"21",X"01",X"25",X"C3",X"E6",X"02",X"21",X"18",X"23",
		X"C3",X"79",X"04",X"21",X"1C",X"23",X"C3",X"79",X"04",X"5E",X"23",X"56",X"23",X"7E",X"23",X"66",
		X"6F",X"C3",X"8F",X"03",X"0E",X"07",X"21",X"01",X"35",X"11",X"7D",X"42",X"C3",X"E6",X"02",X"3A",
		X"0A",X"23",X"21",X"01",X"3C",X"C3",X"30",X"03",X"00",X"00",X"21",X"14",X"23",X"C3",X"79",X"04",
		X"CD",X"F0",X"04",X"CD",X"61",X"0A",X"CD",X"52",X"04",X"CD",X"6D",X"04",X"CD",X"73",X"04",X"CD",
		X"9A",X"04",X"CD",X"84",X"04",X"CD",X"8F",X"04",X"C3",X"E9",X"0A",X"1A",X"77",X"23",X"13",X"05",
		X"C2",X"BB",X"04",X"C9",X"E5",X"23",X"23",X"5E",X"23",X"56",X"23",X"4E",X"23",X"46",X"E1",X"D5",
		X"5E",X"23",X"56",X"EB",X"D1",X"C9",X"7D",X"E6",X"07",X"D3",X"00",X"C5",X"06",X"03",X"7C",X"1F",
		X"67",X"7D",X"1F",X"6F",X"05",X"C2",X"DE",X"04",X"7C",X"E6",X"3F",X"F6",X"20",X"67",X"C1",X"C9",
		X"21",X"00",X"24",X"36",X"00",X"23",X"7C",X"FE",X"40",X"C2",X"F3",X"04",X"C9",X"1D",X"1B",X"0E",
		X"11",X"1B",X"1E",X"0F",X"0B",X"00",X"18",X"04",X"11",X"12",X"1B",X"01",X"14",X"13",X"13",X"0E",
		X"0D",X"1B",X"0E",X"0D",X"0B",X"18",X"1B",X"1D",X"0F",X"0B",X"00",X"18",X"04",X"11",X"1B",X"1B",
		X"01",X"14",X"13",X"13",X"0E",X"0D",X"1B",X"07",X"08",X"2B",X"12",X"02",X"0E",X"11",X"04",X"0F",
		X"0B",X"00",X"18",X"04",X"11",X"2B",X"1D",X"0F",X"0B",X"00",X"18",X"04",X"11",X"2B",X"1E",X"11",
		X"84",X"41",X"A7",X"C8",X"E5",X"21",X"00",X"00",X"C5",X"01",X"05",X"00",X"09",X"3D",X"C2",X"49",
		X"05",X"19",X"EB",X"C1",X"E1",X"C9",X"F7",X"C5",X"E5",X"1A",X"D3",X"03",X"DB",X"03",X"2F",X"A6",
		X"77",X"23",X"13",X"1A",X"D3",X"03",X"DB",X"03",X"2F",X"A6",X"77",X"23",X"13",X"AF",X"D3",X"03",
		X"DB",X"03",X"2F",X"A6",X"77",X"E1",X"01",X"20",X"00",X"09",X"C1",X"05",X"C2",X"57",X"05",X"C9",
		X"21",X"04",X"20",X"CD",X"C4",X"04",X"F7",X"C5",X"E5",X"1A",X"D3",X"03",X"DB",X"03",X"AE",X"77",
		X"23",X"13",X"0D",X"C2",X"89",X"05",X"AF",X"D3",X"03",X"DB",X"03",X"AE",X"77",X"E1",X"01",X"20",
		X"00",X"09",X"C1",X"05",X"C2",X"87",X"05",X"C9",X"C5",X"E5",X"1A",X"77",X"23",X"13",X"0D",X"C2",
		X"AA",X"05",X"E1",X"01",X"20",X"00",X"09",X"C1",X"05",X"C2",X"A8",X"05",X"C9",X"21",X"4A",X"20",
		X"AF",X"BE",X"C2",X"0E",X"4E",X"C9",X"31",X"FF",X"23",X"CD",X"15",X"02",X"21",X"00",X"23",X"11",
		X"50",X"41",X"06",X"30",X"CD",X"BB",X"04",X"CD",X"20",X"02",X"CD",X"2B",X"02",X"CD",X"A7",X"50",
		X"AF",X"D3",X"04",X"D3",X"06",X"CD",X"D4",X"01",X"FB",X"CD",X"A0",X"04",X"CD",X"6E",X"03",X"CD",
		X"A8",X"06",X"CD",X"00",X"50",X"CD",X"F7",X"06",X"CD",X"A0",X"04",X"01",X"51",X"45",X"CD",X"64",
		X"0A",X"21",X"1A",X"27",X"11",X"7F",X"45",X"0E",X"15",X"CD",X"E6",X"02",X"21",X"18",X"29",X"0E",
		X"11",X"CD",X"E6",X"02",X"21",X"15",X"29",X"11",X"1A",X"46",X"01",X"02",X"10",X"CD",X"A8",X"05",
		X"21",X"13",X"29",X"E5",X"11",X"FE",X"42",X"06",X"12",X"CD",X"DB",X"03",X"E1",X"2E",X"11",X"E5",
		X"11",X"4F",X"44",X"06",X"11",X"CD",X"DB",X"03",X"E1",X"2E",X"0E",X"E5",X"11",X"E7",X"42",X"06",
		X"0B",X"CD",X"DB",X"03",X"E1",X"2E",X"0C",X"E5",X"11",X"DB",X"42",X"06",X"0C",X"CD",X"DB",X"03",
		X"E1",X"2E",X"0A",X"E5",X"11",X"10",X"43",X"06",X"03",X"CD",X"DB",X"03",X"E1",X"2E",X"08",X"11",
		X"E1",X"44",X"06",X"03",X"CD",X"DB",X"03",X"CD",X"6E",X"03",X"11",X"A5",X"45",X"1A",X"FE",X"FF",
		X"CA",X"84",X"06",X"1A",X"6F",X"13",X"1A",X"67",X"13",X"0E",X"0A",X"CD",X"E6",X"02",X"CD",X"85",
		X"03",X"C3",X"6D",X"06",X"06",X"0C",X"11",X"1A",X"46",X"C5",X"21",X"15",X"29",X"01",X"02",X"10",
		X"CD",X"A8",X"05",X"3E",X"08",X"CD",X"78",X"03",X"C1",X"05",X"C2",X"89",X"06",X"CD",X"6E",X"03",
		X"CD",X"7A",X"4C",X"D3",X"05",X"C3",X"E9",X"05",X"21",X"08",X"C6",X"11",X"01",X"30",X"3E",X"03",
		X"DF",X"21",X"08",X"26",X"11",X"73",X"44",X"06",X"08",X"CD",X"DB",X"03",X"24",X"0E",X"16",X"C3",
		X"E6",X"02",X"21",X"14",X"2C",X"11",X"67",X"44",X"0E",X"0C",X"CD",X"54",X"03",X"06",X"08",X"AF",
		X"C5",X"21",X"14",X"CC",X"11",X"01",X"18",X"F5",X"DF",X"CD",X"8A",X"03",X"F1",X"3C",X"FE",X"08",
		X"C2",X"D1",X"06",X"C1",X"05",X"C2",X"CF",X"06",X"3E",X"06",X"21",X"14",X"CC",X"11",X"01",X"18",
		X"DF",X"CD",X"6E",X"03",X"C3",X"F0",X"04",X"CD",X"D9",X"01",X"CD",X"15",X"02",X"CD",X"5A",X"15",
		X"CD",X"5F",X"15",X"CD",X"A0",X"04",X"CD",X"92",X"0A",X"DB",X"02",X"E6",X"10",X"CA",X"15",X"07",
		X"06",X"20",X"CD",X"33",X"09",X"21",X"0B",X"23",X"34",X"CD",X"CB",X"07",X"CD",X"D4",X"01",X"21",
		X"37",X"20",X"AF",X"BE",X"C2",X"2C",X"07",X"D3",X"05",X"C3",X"1F",X"07",X"36",X"00",X"21",X"0B",
		X"23",X"36",X"00",X"CD",X"51",X"07",X"CD",X"15",X"02",X"CD",X"5A",X"15",X"CD",X"5F",X"15",X"DB",
		X"02",X"E6",X"10",X"CA",X"4B",X"07",X"06",X"DF",X"CD",X"3D",X"09",X"CD",X"F0",X"04",X"C3",X"D4",
		X"01",X"CD",X"48",X"16",X"06",X"08",X"CD",X"2E",X"09",X"2A",X"04",X"20",X"E5",X"01",X"02",X"18",
		X"CD",X"0F",X"09",X"E1",X"E5",X"FF",X"11",X"03",X"07",X"AF",X"DF",X"E1",X"11",X"B1",X"44",X"01",
		X"02",X"18",X"CD",X"AB",X"07",X"3E",X"40",X"CD",X"78",X"03",X"06",X"F7",X"CD",X"3D",X"09",X"06",
		X"08",X"AF",X"C5",X"2A",X"04",X"20",X"F5",X"FF",X"F1",X"11",X"03",X"07",X"F5",X"DF",X"3E",X"01",
		X"CD",X"78",X"03",X"F1",X"3C",X"FE",X"08",X"C2",X"83",X"07",X"C1",X"05",X"C2",X"81",X"07",X"2A",
		X"04",X"20",X"FF",X"AF",X"11",X"03",X"07",X"DF",X"C3",X"6E",X"03",X"F7",X"C5",X"E5",X"1A",X"D3",
		X"03",X"DB",X"03",X"77",X"23",X"13",X"0D",X"C2",X"AE",X"07",X"AF",X"D3",X"03",X"DB",X"03",X"77",
		X"E1",X"01",X"20",X"00",X"09",X"C1",X"05",X"C2",X"AC",X"07",X"C9",X"06",X"01",X"21",X"00",X"20",
		X"70",X"2E",X"4F",X"70",X"2E",X"72",X"70",X"2E",X"84",X"70",X"2E",X"7B",X"70",X"2E",X"8D",X"70",
		X"CD",X"42",X"0B",X"70",X"2E",X"13",X"70",X"2E",X"39",X"70",X"2E",X"4E",X"7E",X"FE",X"07",X"D2",
		X"65",X"08",X"FE",X"06",X"CA",X"58",X"08",X"FE",X"05",X"CA",X"58",X"08",X"FE",X"04",X"CA",X"45");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
