library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity gamate_bios_bit is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of gamate_bios_bit is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"4C",X"01",X"F3",X"4C",X"E0",X"F2",X"4C",X"EB",X"F2",X"4C",X"F6",X"F2",X"4C",X"90",X"F5",X"4C",
		X"67",X"FB",X"4C",X"1D",X"F3",X"4C",X"C7",X"F5",X"4C",X"AE",X"F3",X"4C",X"F7",X"F4",X"4C",X"7B",
		X"F4",X"4C",X"4A",X"F5",X"4C",X"1A",X"F6",X"4C",X"2F",X"F6",X"4C",X"18",X"FF",X"4C",X"21",X"FF",
		X"4C",X"79",X"FB",X"4C",X"5A",X"FF",X"4C",X"A9",X"FB",X"A9",X"00",X"85",X"16",X"85",X"17",X"85",
		X"15",X"A5",X"16",X"8D",X"02",X"50",X"A5",X"17",X"8D",X"03",X"50",X"20",X"90",X"F5",X"A9",X"B8",
		X"85",X"00",X"85",X"02",X"A9",X"F1",X"85",X"01",X"85",X"03",X"A9",X"58",X"85",X"1C",X"A9",X"10",
		X"85",X"1D",X"A2",X"20",X"A0",X"90",X"20",X"C7",X"F5",X"A0",X"00",X"20",X"EB",X"F2",X"8C",X"03",
		X"50",X"C8",X"C0",X"60",X"90",X"F5",X"20",X"F6",X"F2",X"A9",X"06",X"85",X"21",X"A9",X"10",X"85",
		X"00",X"85",X"02",X"A9",X"F1",X"85",X"01",X"85",X"03",X"A9",X"38",X"85",X"1C",X"A9",X"18",X"85",
		X"1D",X"A2",X"30",X"A0",X"A4",X"20",X"C7",X"F5",X"A9",X"68",X"85",X"00",X"85",X"02",X"A9",X"F2",
		X"85",X"01",X"85",X"03",X"A9",X"08",X"85",X"1C",X"A9",X"08",X"85",X"1D",X"A2",X"68",X"A0",X"B4",
		X"20",X"C7",X"F5",X"A9",X"70",X"85",X"00",X"85",X"02",X"A9",X"F2",X"85",X"01",X"85",X"03",X"A9",
		X"50",X"85",X"1C",X"A9",X"08",X"85",X"1D",X"A2",X"28",X"A0",X"BE",X"20",X"C7",X"F5",X"C6",X"21",
		X"F0",X"2B",X"20",X"F6",X"F2",X"A9",X"58",X"85",X"1C",X"A9",X"28",X"85",X"1D",X"A2",X"20",X"A0",
		X"A4",X"A9",X"00",X"20",X"18",X"FF",X"A9",X"58",X"85",X"1C",X"A9",X"28",X"85",X"1D",X"A2",X"20",
		X"A0",X"A4",X"A9",X"00",X"20",X"21",X"FF",X"20",X"F6",X"F2",X"4C",X"7D",X"F0",X"A0",X"06",X"20",
		X"F6",X"F2",X"88",X"10",X"FA",X"A9",X"01",X"85",X"0C",X"A9",X"FF",X"85",X"0A",X"4C",X"20",X"60",
		X"00",X"7F",X"7F",X"7F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"7F",X"7F",X"7F",X"00",X"FF",X"80",X"FF",X"80",X"87",X"80",X"83",
		X"80",X"87",X"80",X"FF",X"80",X"FF",X"80",X"87",X"80",X"83",X"80",X"87",X"80",X"FF",X"80",X"FF",
		X"00",X"81",X"01",X"E1",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"C0",X"00",X"F0",X"00",X"F8",
		X"00",X"F8",X"00",X"F8",X"00",X"F3",X"03",X"C3",X"00",X"FF",X"F8",X"FF",X"78",X"7F",X"78",X"7F",
		X"78",X"7F",X"78",X"7F",X"78",X"7F",X"78",X"7F",X"78",X"7F",X"78",X"7F",X"78",X"FF",X"F8",X"FF",
		X"00",X"E7",X"07",X"E7",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",
		X"00",X"80",X"00",X"80",X"00",X"F0",X"00",X"F0",X"00",X"FF",X"FC",X"FF",X"3C",X"3F",X"3C",X"3F",
		X"3C",X"3F",X"3C",X"3F",X"3C",X"3F",X"3C",X"3F",X"3C",X"3F",X"3C",X"3F",X"3C",X"3F",X"3C",X"3F",
		X"00",X"FF",X"00",X"FF",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",
		X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"00",X"00",X"07",X"1C",X"38",X"70",X"70",
		X"E0",X"E0",X"E0",X"E0",X"70",X"70",X"3E",X"1F",X"00",X"00",X"00",X"E8",X"38",X"18",X"08",X"00",
		X"00",X"00",X"7C",X"38",X"38",X"38",X"F9",X"BB",X"00",X"00",X"00",X"03",X"03",X"07",X"0D",X"09",
		X"19",X"30",X"3F",X"60",X"C0",X"C0",X"80",X"C1",X"00",X"00",X"00",X"01",X"00",X"80",X"81",X"81",
		X"C1",X"C1",X"C1",X"C3",X"C2",X"E2",X"E2",X"F7",X"00",X"00",X"00",X"C0",X"E0",X"E0",X"E0",X"60",
		X"61",X"71",X"33",X"34",X"34",X"3C",X"18",X"18",X"00",X"00",X"00",X"38",X"70",X"70",X"F0",X"B0",
		X"B0",X"30",X"70",X"70",X"61",X"61",X"E3",X"F7",X"00",X"00",X"00",X"06",X"06",X"0F",X"1B",X"13",
		X"33",X"61",X"7F",X"C1",X"81",X"81",X"01",X"83",X"00",X"00",X"00",X"1F",X"31",X"63",X"03",X"03",
		X"83",X"83",X"87",X"87",X"86",X"C6",X"C6",X"EF",X"00",X"00",X"00",X"FB",X"99",X"89",X"81",X"01",
		X"01",X"01",X"03",X"03",X"03",X"03",X"03",X"07",X"00",X"00",X"00",X"FF",X"C3",X"C0",X"84",X"84",
		X"8C",X"F8",X"88",X"00",X"03",X"06",X"06",X"FE",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",
		X"00",X"00",X"00",X"F1",X"5B",X"5F",X"55",X"51",X"3C",X"42",X"B9",X"A5",X"B9",X"A5",X"42",X"3C",
		X"00",X"38",X"44",X"BA",X"A2",X"BA",X"44",X"38",X"00",X"00",X"F8",X"CC",X"F8",X"CC",X"CC",X"F8",
		X"00",X"00",X"78",X"30",X"30",X"30",X"30",X"78",X"00",X"00",X"FC",X"30",X"30",X"30",X"30",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"78",X"CC",X"C0",X"C0",X"CC",X"78",
		X"00",X"00",X"78",X"CC",X"CC",X"CC",X"CC",X"78",X"00",X"00",X"F8",X"CC",X"CC",X"F8",X"D0",X"CC",
		X"00",X"00",X"F8",X"CC",X"CC",X"F8",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"30",
		X"00",X"38",X"44",X"BA",X"A2",X"BA",X"44",X"38",X"3F",X"19",X"19",X"1F",X"19",X"19",X"19",X"3F",
		X"3E",X"9C",X"9C",X"1C",X"9C",X"9C",X"9C",X"3E",X"FE",X"38",X"38",X"38",X"38",X"38",X"38",X"38",
		X"A5",X"0B",X"C9",X"08",X"90",X"FA",X"A9",X"00",X"85",X"0B",X"60",X"A5",X"0B",X"C9",X"05",X"90",
		X"FA",X"A9",X"00",X"85",X"0B",X"60",X"A5",X"0B",X"C9",X"18",X"90",X"FA",X"A9",X"00",X"85",X"0B",
		X"60",X"A9",X"C0",X"85",X"00",X"85",X"02",X"A9",X"F2",X"85",X"01",X"85",X"03",X"A9",X"20",X"85",
		X"1C",X"A9",X"08",X"85",X"1D",X"A2",X"40",X"A0",X"8C",X"20",X"C7",X"F5",X"60",X"8A",X"4A",X"4A",
		X"4A",X"09",X"80",X"85",X"18",X"84",X"19",X"A0",X"00",X"B1",X"00",X"85",X"1B",X"C8",X"B1",X"00",
		X"20",X"3A",X"F3",X"E6",X"18",X"C6",X"1B",X"D0",X"F4",X"60",X"85",X"1A",X"98",X"48",X"A9",X"40",
		X"05",X"15",X"8D",X"01",X"50",X"A5",X"18",X"8D",X"04",X"50",X"A5",X"19",X"8D",X"05",X"50",X"A5",
		X"1A",X"C9",X"61",X"B0",X"41",X"C9",X"41",X"B0",X"25",X"A2",X"00",X"C9",X"20",X"F0",X"0E",X"B0",
		X"05",X"A2",X"00",X"4C",X"6D",X"F3",X"38",X"E9",X"2F",X"0A",X"0A",X"0A",X"AA",X"86",X"1A",X"A0",
		X"07",X"BD",X"29",X"60",X"8D",X"07",X"50",X"E8",X"88",X"10",X"F6",X"4C",X"AB",X"F3",X"38",X"E9",
		X"41",X"0A",X"0A",X"0A",X"AA",X"86",X"1A",X"A0",X"07",X"BD",X"81",X"60",X"8D",X"07",X"50",X"E8",
		X"88",X"10",X"F6",X"4C",X"AB",X"F3",X"38",X"E9",X"61",X"0A",X"0A",X"0A",X"AA",X"86",X"1A",X"A0",
		X"07",X"BD",X"51",X"61",X"8D",X"07",X"50",X"E8",X"88",X"10",X"F6",X"68",X"A8",X"60",X"A5",X"00",
		X"48",X"A5",X"01",X"48",X"A9",X"40",X"05",X"15",X"8D",X"01",X"50",X"A0",X"00",X"B1",X"00",X"C9",
		X"FE",X"D0",X"03",X"4C",X"F2",X"F3",X"85",X"19",X"A9",X"00",X"85",X"18",X"20",X"75",X"F4",X"B1",
		X"00",X"C9",X"FF",X"F0",X"17",X"85",X"1A",X"20",X"75",X"F4",X"B1",X"00",X"85",X"1B",X"A5",X"06",
		X"85",X"02",X"A5",X"07",X"85",X"03",X"20",X"30",X"F4",X"4C",X"CC",X"F3",X"20",X"75",X"F4",X"4C",
		X"BD",X"F3",X"68",X"85",X"01",X"68",X"85",X"00",X"A0",X"00",X"B1",X"00",X"C9",X"FE",X"D0",X"03",
		X"4C",X"2F",X"F4",X"85",X"19",X"A9",X"80",X"85",X"18",X"20",X"75",X"F4",X"B1",X"00",X"C9",X"FF",
		X"F0",X"17",X"85",X"1A",X"20",X"75",X"F4",X"B1",X"00",X"85",X"1B",X"A5",X"08",X"85",X"02",X"A5",
		X"09",X"85",X"03",X"20",X"30",X"F4",X"4C",X"09",X"F4",X"20",X"75",X"F4",X"4C",X"FA",X"F3",X"60",
		X"48",X"98",X"48",X"A5",X"1A",X"D0",X"0A",X"A5",X"18",X"18",X"65",X"1B",X"85",X"18",X"4C",X"71",
		X"F4",X"C9",X"20",X"90",X"07",X"E6",X"03",X"38",X"E9",X"20",X"B0",X"F5",X"0A",X"0A",X"0A",X"85",
		X"1A",X"A5",X"18",X"8D",X"04",X"50",X"A5",X"19",X"0A",X"0A",X"0A",X"8D",X"05",X"50",X"A4",X"1A",
		X"A2",X"07",X"B1",X"02",X"8D",X"07",X"50",X"C8",X"CA",X"10",X"F7",X"E6",X"18",X"C6",X"1B",X"D0",
		X"E0",X"68",X"A8",X"68",X"60",X"C8",X"D0",X"02",X"E6",X"01",X"60",X"A5",X"00",X"48",X"A5",X"01",
		X"48",X"A9",X"40",X"05",X"15",X"8D",X"01",X"50",X"A0",X"00",X"B1",X"00",X"C9",X"FE",X"D0",X"03",
		X"4C",X"BC",X"F4",X"85",X"19",X"A9",X"00",X"85",X"18",X"20",X"75",X"F4",X"B1",X"00",X"C9",X"FF",
		X"F0",X"14",X"85",X"1A",X"A9",X"01",X"85",X"1B",X"A5",X"06",X"85",X"02",X"A5",X"07",X"85",X"03",
		X"20",X"30",X"F4",X"4C",X"99",X"F4",X"20",X"75",X"F4",X"4C",X"8A",X"F4",X"68",X"85",X"01",X"68",
		X"85",X"00",X"A0",X"00",X"B1",X"00",X"C9",X"FE",X"D0",X"03",X"4C",X"F6",X"F4",X"85",X"19",X"A9",
		X"80",X"85",X"18",X"20",X"75",X"F4",X"B1",X"00",X"C9",X"FF",X"F0",X"14",X"85",X"1A",X"A9",X"01",
		X"85",X"1B",X"A5",X"08",X"85",X"02",X"A5",X"09",X"85",X"03",X"20",X"30",X"F4",X"4C",X"D3",X"F4",
		X"20",X"75",X"F4",X"4C",X"C4",X"F4",X"60",X"A9",X"00",X"05",X"15",X"8D",X"01",X"50",X"A0",X"E6",
		X"8C",X"05",X"50",X"A9",X"00",X"A2",X"20",X"8D",X"04",X"50",X"8D",X"07",X"50",X"CA",X"D0",X"FA",
		X"C8",X"C0",X"FF",X"D0",X"EB",X"A0",X"00",X"B1",X"00",X"C9",X"FE",X"F0",X"2C",X"18",X"69",X"E6",
		X"8D",X"05",X"50",X"A9",X"00",X"8D",X"04",X"50",X"20",X"75",X"F4",X"B1",X"00",X"C9",X"FF",X"F0",
		X"13",X"85",X"1A",X"20",X"75",X"F4",X"B1",X"00",X"AA",X"A5",X"1A",X"8D",X"07",X"50",X"CA",X"D0",
		X"FA",X"4C",X"28",X"F5",X"20",X"75",X"F4",X"D0",X"CE",X"60",X"A9",X"00",X"05",X"15",X"8D",X"01",
		X"50",X"A0",X"E6",X"8C",X"05",X"50",X"A9",X"00",X"A2",X"20",X"8D",X"04",X"50",X"8D",X"07",X"50",
		X"CA",X"D0",X"FA",X"C8",X"C0",X"FF",X"D0",X"EB",X"A0",X"00",X"B1",X"00",X"C9",X"FE",X"F0",X"1F",
		X"18",X"69",X"E6",X"8D",X"05",X"50",X"A9",X"00",X"8D",X"04",X"50",X"20",X"75",X"F4",X"B1",X"00",
		X"C9",X"FF",X"F0",X"06",X"8D",X"07",X"50",X"4C",X"7B",X"F5",X"20",X"75",X"F4",X"D0",X"DB",X"60",
		X"A9",X"80",X"05",X"15",X"8D",X"01",X"50",X"A9",X"00",X"85",X"1E",X"20",X"AD",X"F5",X"A9",X"80",
		X"85",X"1E",X"20",X"AD",X"F5",X"A9",X"40",X"05",X"15",X"8D",X"01",X"50",X"60",X"A0",X"00",X"A5",
		X"1E",X"8D",X"04",X"50",X"8C",X"05",X"50",X"A2",X"20",X"A9",X"00",X"8D",X"07",X"50",X"CA",X"D0",
		X"FA",X"C8",X"C0",X"C8",X"D0",X"E9",X"60",X"86",X"18",X"84",X"19",X"46",X"18",X"46",X"18",X"46",
		X"18",X"A5",X"18",X"48",X"A9",X"40",X"05",X"15",X"8D",X"01",X"50",X"46",X"1C",X"46",X"1C",X"46",
		X"1C",X"20",X"F5",X"F5",X"A5",X"02",X"85",X"00",X"A5",X"03",X"85",X"01",X"68",X"09",X"80",X"85",
		X"18",X"20",X"F5",X"F5",X"60",X"A5",X"1C",X"85",X"1E",X"A0",X"00",X"A5",X"18",X"8D",X"04",X"50",
		X"A5",X"19",X"8D",X"05",X"50",X"A5",X"1D",X"85",X"1F",X"B1",X"00",X"8D",X"07",X"50",X"C8",X"C6",
		X"1F",X"D0",X"F6",X"E6",X"18",X"C6",X"1E",X"D0",X"E2",X"60",X"A2",X"10",X"A0",X"00",X"A9",X"FF",
		X"99",X"23",X"00",X"99",X"28",X"00",X"98",X"18",X"69",X"08",X"A8",X"CA",X"D0",X"F0",X"60",X"48",
		X"98",X"48",X"8A",X"48",X"A2",X"08",X"A0",X"00",X"B9",X"28",X"00",X"C9",X"FF",X"F0",X"19",X"B9",
		X"26",X"00",X"4A",X"4A",X"4A",X"85",X"18",X"85",X"1E",X"B9",X"27",X"00",X"29",X"F8",X"85",X"19",
		X"4A",X"4A",X"4A",X"85",X"1F",X"20",X"C4",X"F6",X"98",X"18",X"69",X"08",X"A8",X"CA",X"D0",X"D8",
		X"A2",X"08",X"A0",X"00",X"B9",X"68",X"00",X"C9",X"FF",X"F0",X"19",X"B9",X"66",X"00",X"4A",X"4A",
		X"4A",X"85",X"18",X"85",X"1E",X"B9",X"67",X"00",X"29",X"F8",X"85",X"19",X"4A",X"4A",X"4A",X"85",
		X"1F",X"20",X"9D",X"F9",X"98",X"18",X"69",X"08",X"A8",X"CA",X"D0",X"D8",X"A2",X"08",X"A0",X"00",
		X"8A",X"48",X"A2",X"00",X"B9",X"21",X"00",X"9D",X"00",X"03",X"C8",X"E8",X"E0",X"08",X"D0",X"F4",
		X"68",X"AA",X"AD",X"02",X"03",X"C9",X"FF",X"F0",X"0F",X"20",X"88",X"F7",X"20",X"ED",X"F7",X"20",
		X"A1",X"F8",X"20",X"CE",X"F8",X"20",X"FA",X"F8",X"CA",X"D0",X"D5",X"20",X"63",X"F9",X"68",X"AA",
		X"68",X"A8",X"68",X"60",X"98",X"48",X"8A",X"48",X"A9",X"40",X"05",X"15",X"8D",X"01",X"50",X"A5",
		X"1F",X"18",X"69",X"E6",X"85",X"1F",X"A0",X"00",X"A9",X"03",X"85",X"1B",X"A6",X"1E",X"A5",X"1F",
		X"85",X"1D",X"8D",X"05",X"50",X"8E",X"04",X"50",X"AD",X"06",X"50",X"99",X"08",X"03",X"E6",X"1D",
		X"A5",X"1D",X"8D",X"05",X"50",X"8E",X"04",X"50",X"AD",X"06",X"50",X"99",X"09",X"03",X"E6",X"1D",
		X"A5",X"1D",X"8D",X"05",X"50",X"8E",X"04",X"50",X"AD",X"06",X"50",X"99",X"0A",X"03",X"C8",X"C8",
		X"C8",X"E8",X"C6",X"1B",X"D0",X"C8",X"A0",X"00",X"A9",X"03",X"85",X"1C",X"A6",X"18",X"A9",X"03",
		X"85",X"1D",X"8E",X"04",X"50",X"A5",X"19",X"8D",X"05",X"50",X"B9",X"08",X"03",X"20",X"4B",X"F7",
		X"C8",X"C6",X"1D",X"D0",X"F5",X"E8",X"C6",X"1C",X"D0",X"E4",X"A5",X"18",X"C9",X"80",X"B0",X"06",
		X"09",X"80",X"85",X"18",X"D0",X"D0",X"68",X"AA",X"68",X"A8",X"60",X"85",X"1A",X"8A",X"48",X"98",
		X"48",X"A5",X"06",X"85",X"02",X"A5",X"07",X"85",X"03",X"A6",X"18",X"E0",X"80",X"90",X"08",X"A5",
		X"08",X"85",X"02",X"A5",X"09",X"85",X"03",X"A5",X"1A",X"C9",X"20",X"90",X"07",X"E6",X"03",X"38",
		X"E9",X"20",X"B0",X"F5",X"0A",X"0A",X"0A",X"A8",X"A2",X"08",X"B1",X"02",X"8D",X"07",X"50",X"C8",
		X"CA",X"D0",X"F7",X"68",X"A8",X"68",X"AA",X"60",X"48",X"8A",X"48",X"98",X"48",X"A9",X"40",X"05",
		X"15",X"8D",X"01",X"50",X"AD",X"00",X"03",X"4A",X"4A",X"4A",X"85",X"18",X"AD",X"01",X"03",X"85",
		X"19",X"A9",X"08",X"85",X"00",X"A9",X"03",X"85",X"01",X"A6",X"18",X"A0",X"00",X"A5",X"19",X"85",
		X"1B",X"A5",X"1B",X"8D",X"05",X"50",X"8E",X"04",X"50",X"AD",X"06",X"50",X"91",X"00",X"E6",X"1B",
		X"C8",X"C0",X"30",X"F0",X"0C",X"C0",X"20",X"F0",X"04",X"C0",X"10",X"D0",X"E4",X"E8",X"4C",X"AD",
		X"F7",X"A5",X"18",X"AA",X"C9",X"80",X"B0",X"0F",X"A9",X"38",X"85",X"00",X"A9",X"03",X"85",X"01",
		X"8A",X"09",X"80",X"85",X"18",X"D0",X"C2",X"68",X"A8",X"68",X"AA",X"68",X"60",X"48",X"8A",X"48",
		X"98",X"48",X"A9",X"40",X"05",X"15",X"8D",X"01",X"50",X"A9",X"68",X"85",X"00",X"A9",X"03",X"85",
		X"01",X"A9",X"00",X"85",X"1B",X"AD",X"02",X"03",X"A8",X"20",X"4E",X"F8",X"20",X"95",X"F8",X"98",
		X"18",X"69",X"02",X"20",X"4E",X"F8",X"20",X"95",X"F8",X"98",X"18",X"69",X"01",X"20",X"4E",X"F8",
		X"20",X"95",X"F8",X"98",X"18",X"69",X"03",X"20",X"4E",X"F8",X"A5",X"1B",X"D0",X"0D",X"E6",X"1B",
		X"A9",X"98",X"85",X"00",X"A9",X"03",X"85",X"01",X"4C",X"05",X"F8",X"A0",X"0F",X"A9",X"00",X"99",
		X"88",X"03",X"99",X"B8",X"03",X"88",X"10",X"F7",X"68",X"A8",X"68",X"AA",X"68",X"60",X"85",X"1A",
		X"8A",X"48",X"98",X"48",X"A5",X"06",X"85",X"02",X"A5",X"07",X"85",X"03",X"A5",X"1B",X"F0",X"08",
		X"A5",X"08",X"85",X"02",X"A5",X"09",X"85",X"03",X"A5",X"1A",X"C9",X"20",X"90",X"07",X"E6",X"03",
		X"38",X"E9",X"20",X"B0",X"F5",X"0A",X"0A",X"0A",X"A8",X"A5",X"00",X"48",X"A2",X"08",X"86",X"1C",
		X"A2",X"00",X"B1",X"02",X"81",X"00",X"C8",X"E6",X"00",X"C6",X"1C",X"D0",X"F5",X"68",X"85",X"00",
		X"68",X"A8",X"68",X"AA",X"60",X"A5",X"00",X"18",X"69",X"08",X"85",X"00",X"90",X"02",X"E6",X"01",
		X"60",X"48",X"8A",X"48",X"98",X"48",X"AD",X"00",X"03",X"29",X"07",X"F0",X"1B",X"A8",X"A2",X"0F",
		X"5E",X"68",X"03",X"7E",X"78",X"03",X"7E",X"88",X"03",X"5E",X"98",X"03",X"7E",X"A8",X"03",X"7E",
		X"B8",X"03",X"CA",X"10",X"EB",X"88",X"D0",X"E6",X"68",X"A8",X"68",X"AA",X"68",X"60",X"48",X"8A",
		X"48",X"98",X"48",X"A2",X"2F",X"BD",X"68",X"03",X"1D",X"98",X"03",X"49",X"FF",X"A8",X"3D",X"08",
		X"03",X"1D",X"68",X"03",X"9D",X"68",X"03",X"98",X"3D",X"38",X"03",X"1D",X"98",X"03",X"9D",X"98",
		X"03",X"CA",X"10",X"E1",X"68",X"A8",X"68",X"AA",X"68",X"60",X"48",X"8A",X"48",X"98",X"48",X"A9",
		X"40",X"05",X"15",X"8D",X"01",X"50",X"AD",X"00",X"03",X"4A",X"4A",X"4A",X"85",X"18",X"AA",X"AD",
		X"01",X"03",X"85",X"19",X"A0",X"00",X"A5",X"19",X"8D",X"05",X"50",X"8E",X"04",X"50",X"B9",X"68",
		X"03",X"8D",X"07",X"50",X"C8",X"C0",X"30",X"F0",X"0C",X"C0",X"20",X"F0",X"04",X"C0",X"10",X"D0",
		X"ED",X"E8",X"4C",X"16",X"F9",X"A5",X"18",X"09",X"80",X"85",X"18",X"AA",X"A0",X"00",X"A5",X"19",
		X"8D",X"05",X"50",X"8E",X"04",X"50",X"B9",X"98",X"03",X"8D",X"07",X"50",X"C8",X"C0",X"30",X"F0",
		X"0C",X"C0",X"20",X"F0",X"04",X"C0",X"10",X"D0",X"ED",X"E8",X"4C",X"3E",X"F9",X"68",X"A8",X"68",
		X"AA",X"68",X"60",X"48",X"98",X"48",X"8A",X"48",X"A2",X"08",X"A0",X"00",X"8A",X"48",X"A2",X"00",
		X"B9",X"61",X"00",X"9D",X"00",X"03",X"C8",X"E8",X"E0",X"08",X"D0",X"F4",X"68",X"AA",X"AD",X"02",
		X"03",X"C9",X"FF",X"F0",X"0F",X"20",X"13",X"FA",X"20",X"74",X"FA",X"20",X"B3",X"FA",X"20",X"DA",
		X"FA",X"20",X"06",X"FB",X"CA",X"D0",X"D5",X"68",X"AA",X"68",X"A8",X"68",X"60",X"98",X"48",X"8A",
		X"48",X"A9",X"40",X"05",X"15",X"8D",X"01",X"50",X"A5",X"1F",X"18",X"69",X"E6",X"85",X"1F",X"A0",
		X"00",X"A9",X"02",X"85",X"1B",X"A6",X"1E",X"A5",X"1F",X"85",X"1D",X"8D",X"05",X"50",X"8E",X"04",
		X"50",X"AD",X"06",X"50",X"99",X"08",X"03",X"E6",X"1D",X"A5",X"1D",X"8D",X"05",X"50",X"8E",X"04",
		X"50",X"AD",X"06",X"50",X"99",X"09",X"03",X"C8",X"C8",X"E8",X"C6",X"1B",X"D0",X"D9",X"A0",X"00",
		X"A9",X"02",X"85",X"1C",X"A6",X"18",X"A9",X"02",X"85",X"1D",X"8E",X"04",X"50",X"A5",X"19",X"8D",
		X"05",X"50",X"B9",X"08",X"03",X"20",X"4B",X"F7",X"C8",X"C6",X"1D",X"D0",X"F5",X"E8",X"C6",X"1C",
		X"D0",X"E4",X"A5",X"18",X"C9",X"80",X"B0",X"06",X"09",X"80",X"85",X"18",X"D0",X"D0",X"68",X"AA",
		X"68",X"A8",X"60",X"48",X"8A",X"48",X"98",X"48",X"A9",X"40",X"05",X"15",X"8D",X"01",X"50",X"AD",
		X"00",X"03",X"4A",X"4A",X"4A",X"85",X"18",X"AD",X"01",X"03",X"85",X"19",X"A9",X"08",X"85",X"00",
		X"A9",X"03",X"85",X"01",X"A6",X"18",X"A0",X"00",X"A5",X"19",X"85",X"1B",X"A5",X"1B",X"8D",X"05",
		X"50",X"8E",X"04",X"50",X"AD",X"06",X"50",X"91",X"00",X"E6",X"1B",X"C8",X"C0",X"10",X"F0",X"08",
		X"C0",X"08",X"D0",X"E8",X"E8",X"4C",X"38",X"FA",X"A5",X"18",X"AA",X"C9",X"80",X"B0",X"0F",X"A9",
		X"38",X"85",X"00",X"A9",X"03",X"85",X"01",X"8A",X"09",X"80",X"85",X"18",X"D0",X"C6",X"68",X"A8",
		X"68",X"AA",X"68",X"60",X"48",X"8A",X"48",X"98",X"48",X"A9",X"68",X"85",X"00",X"A9",X"03",X"85",
		X"01",X"A9",X"00",X"85",X"1B",X"AD",X"02",X"03",X"A8",X"20",X"4E",X"F8",X"20",X"95",X"F8",X"A5",
		X"1B",X"D0",X"0D",X"E6",X"1B",X"A9",X"98",X"85",X"00",X"A9",X"03",X"85",X"01",X"4C",X"85",X"FA",
		X"A0",X"07",X"A9",X"00",X"99",X"70",X"03",X"99",X"A0",X"03",X"88",X"10",X"F7",X"68",X"A8",X"68",
		X"AA",X"68",X"60",X"48",X"8A",X"48",X"98",X"48",X"AD",X"00",X"03",X"29",X"07",X"F0",X"15",X"A8",
		X"A2",X"07",X"5E",X"68",X"03",X"7E",X"70",X"03",X"5E",X"98",X"03",X"7E",X"A0",X"03",X"CA",X"10",
		X"F1",X"88",X"D0",X"EC",X"68",X"A8",X"68",X"AA",X"68",X"60",X"48",X"8A",X"48",X"98",X"48",X"A2",
		X"0F",X"BD",X"68",X"03",X"1D",X"98",X"03",X"49",X"FF",X"A8",X"3D",X"08",X"03",X"1D",X"68",X"03",
		X"9D",X"68",X"03",X"98",X"3D",X"38",X"03",X"1D",X"98",X"03",X"9D",X"98",X"03",X"CA",X"10",X"E1",
		X"68",X"A8",X"68",X"AA",X"68",X"60",X"48",X"8A",X"48",X"98",X"48",X"A9",X"40",X"05",X"15",X"8D",
		X"01",X"50",X"AD",X"00",X"03",X"4A",X"4A",X"4A",X"85",X"18",X"AA",X"AD",X"01",X"03",X"85",X"19",
		X"A0",X"00",X"A5",X"19",X"8D",X"05",X"50",X"8E",X"04",X"50",X"B9",X"68",X"03",X"8D",X"07",X"50",
		X"C8",X"C0",X"10",X"F0",X"08",X"C0",X"08",X"D0",X"F1",X"E8",X"4C",X"22",X"FB",X"A5",X"18",X"09",
		X"80",X"85",X"18",X"AA",X"A0",X"00",X"A5",X"19",X"8D",X"05",X"50",X"8E",X"04",X"50",X"B9",X"98",
		X"03",X"8D",X"07",X"50",X"C8",X"C0",X"10",X"F0",X"08",X"C0",X"08",X"D0",X"F1",X"E8",X"4C",X"46",
		X"FB",X"68",X"A8",X"68",X"AA",X"68",X"60",X"A9",X"19",X"85",X"1D",X"A9",X"FF",X"85",X"1C",X"A2",
		X"00",X"A0",X"E6",X"A9",X"00",X"20",X"18",X"FF",X"60",X"98",X"48",X"8A",X"48",X"A5",X"12",X"05",
		X"13",X"D0",X"06",X"A9",X"FF",X"85",X"12",X"85",X"13",X"A5",X"13",X"29",X"04",X"0A",X"0A",X"0A",
		X"0A",X"0A",X"85",X"14",X"A5",X"12",X"29",X"10",X"0A",X"0A",X"0A",X"45",X"14",X"0A",X"26",X"12",
		X"26",X"13",X"68",X"AA",X"68",X"A8",X"A5",X"12",X"60",X"20",X"90",X"F5",X"A9",X"00",X"8D",X"02",
		X"50",X"8D",X"03",X"50",X"8D",X"E0",X"00",X"8D",X"E1",X"00",X"8D",X"E2",X"00",X"8D",X"E5",X"00",
		X"8D",X"E6",X"00",X"A9",X"70",X"8D",X"E3",X"00",X"A9",X"80",X"8D",X"E7",X"00",X"20",X"EB",X"FB",
		X"AD",X"E1",X"00",X"AE",X"E0",X"00",X"A0",X"00",X"20",X"5A",X"FF",X"A9",X"A1",X"85",X"00",X"A9",
		X"00",X"85",X"01",X"A2",X"10",X"A0",X"10",X"20",X"1D",X"F3",X"60",X"A0",X"00",X"B1",X"E2",X"18",
		X"6D",X"E0",X"00",X"8D",X"E0",X"00",X"AD",X"E1",X"00",X"69",X"00",X"8D",X"E1",X"00",X"C8",X"D0",
		X"EC",X"EE",X"E3",X"00",X"AD",X"E3",X"00",X"CD",X"E7",X"00",X"D0",X"E1",X"60",X"78",X"A9",X"00",
		X"85",X"0C",X"A2",X"FF",X"9A",X"58",X"D8",X"A9",X"00",X"85",X"0B",X"A9",X"FF",X"85",X"12",X"85",
		X"13",X"20",X"79",X"FB",X"A5",X"0B",X"F0",X"F9",X"4C",X"2E",X"FC",X"4C",X"39",X"F0",X"A9",X"00",
		X"85",X"0C",X"A9",X"20",X"8D",X"00",X"59",X"AD",X"00",X"5A",X"29",X"01",X"F0",X"2D",X"AD",X"00",
		X"5A",X"29",X"02",X"F0",X"0F",X"20",X"BF",X"FD",X"58",X"A2",X"FF",X"9A",X"A9",X"00",X"8D",X"00",
		X"59",X"4C",X"39",X"F0",X"A2",X"00",X"BD",X"65",X"FC",X"9D",X"00",X"02",X"E8",X"E0",X"10",X"D0",
		X"F5",X"78",X"4C",X"00",X"02",X"AD",X"00",X"58",X"6C",X"FC",X"FF",X"A9",X"55",X"8D",X"00",X"44",
		X"A5",X"0B",X"69",X"3C",X"C5",X"0B",X"D0",X"FC",X"A9",X"AA",X"8D",X"00",X"44",X"78",X"4C",X"00",
		X"FD",X"A9",X"00",X"85",X"0C",X"20",X"5E",X"FD",X"20",X"96",X"FD",X"58",X"A5",X"0B",X"69",X"32",
		X"C5",X"0B",X"D0",X"FC",X"A9",X"00",X"8D",X"00",X"59",X"A9",X"00",X"8D",X"00",X"44",X"4C",X"99",
		X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C3",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"A2",X"00",X"A9",X"55",X"8D",X"00",X"02",X"95",X"00",X"E8",X"D0",X"FB",X"B5",X"00",X"CD",X"00",
		X"02",X"D0",X"48",X"49",X"FF",X"95",X"00",X"E8",X"D0",X"F2",X"AD",X"00",X"02",X"49",X"FF",X"8D",
		X"00",X"02",X"C9",X"55",X"D0",X"E6",X"A9",X"00",X"85",X"E2",X"A9",X"01",X"85",X"E3",X"A0",X"00",
		X"A9",X"55",X"85",X"E4",X"91",X"E2",X"C8",X"D0",X"FB",X"B1",X"E2",X"C5",X"E4",X"D0",X"1C",X"49",
		X"FF",X"91",X"E2",X"C8",X"D0",X"F3",X"A5",X"E4",X"49",X"FF",X"85",X"E4",X"C9",X"55",X"D0",X"E9",
		X"E6",X"E3",X"A5",X"E3",X"C9",X"04",X"D0",X"D8",X"4C",X"81",X"FC",X"4C",X"00",X"FF",X"A9",X"55",
		X"85",X"E4",X"A9",X"00",X"85",X"E8",X"85",X"0A",X"A5",X"E4",X"8D",X"00",X"44",X"AD",X"00",X"4C",
		X"AD",X"00",X"4C",X"AD",X"00",X"4C",X"AD",X"00",X"4C",X"AD",X"00",X"4C",X"AD",X"00",X"4C",X"AD",
		X"00",X"4C",X"AD",X"00",X"4C",X"A5",X"E8",X"F0",X"FC",X"A5",X"0A",X"C5",X"E4",X"D0",X"CC",X"49",
		X"FF",X"C9",X"55",X"D0",X"CB",X"60",X"A9",X"00",X"85",X"E0",X"85",X"E1",X"85",X"E7",X"85",X"E2",
		X"A9",X"E2",X"85",X"E5",X"A9",X"58",X"85",X"E6",X"A9",X"F0",X"85",X"E3",X"20",X"3F",X"FE",X"60",
		X"42",X"49",X"54",X"20",X"43",X"4F",X"52",X"50",X"4F",X"52",X"41",X"54",X"49",X"4F",X"4E",X"78",
		X"D8",X"A2",X"00",X"BD",X"B0",X"FD",X"85",X"04",X"A0",X"09",X"06",X"04",X"2A",X"2A",X"2A",X"8D",
		X"00",X"60",X"88",X"D0",X"F5",X"E8",X"E0",X"0F",X"D0",X"E9",X"A2",X"00",X"AD",X"00",X"60",X"4A",
		X"4A",X"26",X"04",X"E8",X"E0",X"08",X"D0",X"F4",X"A5",X"04",X"C9",X"47",X"D0",X"07",X"20",X"F8",
		X"FD",X"20",X"21",X"FE",X"60",X"4C",X"0D",X"FF",X"A2",X"00",X"BD",X"05",X"60",X"DD",X"08",X"FE",
		X"D0",X"F3",X"E8",X"E0",X"19",X"D0",X"F3",X"60",X"43",X"4F",X"50",X"59",X"52",X"49",X"47",X"48",
		X"54",X"20",X"42",X"49",X"54",X"20",X"43",X"4F",X"52",X"50",X"4F",X"52",X"41",X"54",X"49",X"4F",
		X"4E",X"A9",X"70",X"85",X"E3",X"A9",X"00",X"85",X"E2",X"85",X"E0",X"85",X"E1",X"AD",X"00",X"60",
		X"85",X"E5",X"AD",X"01",X"60",X"85",X"E6",X"A9",X"80",X"85",X"E7",X"20",X"3F",X"FE",X"60",X"A0",
		X"00",X"B1",X"E2",X"18",X"65",X"E0",X"85",X"E0",X"A5",X"E1",X"69",X"00",X"85",X"E1",X"C8",X"D0",
		X"F0",X"E6",X"E3",X"A5",X"E3",X"C5",X"E7",X"D0",X"E8",X"A5",X"E5",X"C5",X"E0",X"D0",X"07",X"A5",
		X"E6",X"C5",X"E1",X"D0",X"01",X"60",X"4C",X"F5",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"A9",X"00",X"8D",X"00",X"59",X"A9",X"FF",X"8D",X"00",X"44",X"4C",X"05",X"FF",X"A9",X"00",X"8D",
		X"00",X"59",X"B9",X"00",X"60",X"4C",X"12",X"FF",X"48",X"A9",X"00",X"85",X"A8",X"68",X"4C",X"27",
		X"FF",X"48",X"A9",X"80",X"85",X"A8",X"68",X"85",X"1A",X"84",X"19",X"8A",X"4A",X"4A",X"4A",X"05",
		X"A8",X"85",X"18",X"A9",X"40",X"05",X"15",X"8D",X"01",X"50",X"A5",X"1C",X"4A",X"4A",X"4A",X"AA",
		X"A5",X"19",X"8D",X"05",X"50",X"A5",X"18",X"8D",X"04",X"50",X"A5",X"1A",X"A4",X"1D",X"8D",X"07",
		X"50",X"88",X"D0",X"FA",X"E6",X"18",X"CA",X"D0",X"E7",X"60",X"48",X"29",X"0F",X"09",X"30",X"85",
		X"A3",X"68",X"4A",X"4A",X"4A",X"4A",X"29",X"0F",X"09",X"30",X"85",X"A2",X"8A",X"29",X"0F",X"09",
		X"30",X"85",X"A5",X"8A",X"4A",X"4A",X"4A",X"4A",X"29",X"0F",X"09",X"30",X"85",X"A4",X"C0",X"FF",
		X"D0",X"09",X"A0",X"20",X"84",X"A6",X"84",X"A7",X"4C",X"9D",X"FF",X"98",X"29",X"0F",X"09",X"30",
		X"85",X"A7",X"98",X"4A",X"4A",X"4A",X"4A",X"29",X"0F",X"09",X"30",X"85",X"A6",X"A0",X"00",X"B9",
		X"A2",X"00",X"C9",X"30",X"D0",X"0A",X"A9",X"20",X"99",X"A2",X"00",X"C8",X"C0",X"05",X"90",X"EF",
		X"A9",X"06",X"85",X"A1",X"60",X"78",X"08",X"48",X"98",X"48",X"E6",X"0B",X"A0",X"03",X"18",X"B9",
		X"0E",X"00",X"69",X"01",X"99",X"0E",X"00",X"90",X"03",X"88",X"10",X"F2",X"A5",X"0C",X"F0",X"03",
		X"20",X"26",X"60",X"68",X"A8",X"68",X"28",X"58",X"40",X"08",X"48",X"AD",X"00",X"48",X"85",X"0A",
		X"A9",X"FF",X"85",X"E8",X"A5",X"0C",X"F0",X"03",X"20",X"23",X"60",X"68",X"28",X"40",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"D9",X"FF",X"0D",X"FC",X"B5",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
