library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity GFX1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of GFX1 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"CC",X"EE",X"11",X"11",X"33",X"EE",X"CC",X"00",X"11",X"33",X"66",X"44",X"44",X"33",X"11",X"00",
		X"11",X"11",X"FF",X"FF",X"11",X"11",X"00",X"00",X"00",X"00",X"77",X"77",X"22",X"00",X"00",X"00",
		X"11",X"99",X"DD",X"DD",X"FF",X"77",X"33",X"00",X"33",X"77",X"55",X"44",X"44",X"66",X"22",X"00",
		X"66",X"FF",X"99",X"99",X"99",X"33",X"22",X"00",X"44",X"66",X"77",X"55",X"44",X"44",X"00",X"00",
		X"44",X"FF",X"FF",X"44",X"44",X"CC",X"CC",X"00",X"00",X"77",X"77",X"66",X"33",X"11",X"00",X"00",
		X"EE",X"FF",X"11",X"11",X"11",X"33",X"22",X"00",X"00",X"55",X"55",X"55",X"55",X"77",X"77",X"00",
		X"66",X"FF",X"99",X"99",X"99",X"FF",X"EE",X"00",X"00",X"44",X"44",X"44",X"66",X"33",X"11",X"00",
		X"00",X"00",X"88",X"FF",X"77",X"00",X"00",X"00",X"66",X"77",X"55",X"44",X"44",X"66",X"66",X"00",
		X"66",X"77",X"DD",X"DD",X"99",X"99",X"66",X"00",X"00",X"33",X"44",X"44",X"55",X"77",X"33",X"00",
		X"CC",X"EE",X"BB",X"99",X"99",X"99",X"00",X"00",X"33",X"77",X"44",X"44",X"44",X"77",X"33",X"00",
		X"FF",X"FF",X"44",X"44",X"44",X"FF",X"FF",X"00",X"11",X"33",X"66",X"44",X"66",X"33",X"11",X"00",
		X"66",X"FF",X"99",X"99",X"99",X"FF",X"FF",X"00",X"33",X"77",X"44",X"44",X"44",X"77",X"77",X"00",
		X"22",X"33",X"11",X"11",X"33",X"EE",X"CC",X"00",X"22",X"66",X"44",X"44",X"66",X"33",X"11",X"00",
		X"CC",X"EE",X"33",X"11",X"11",X"FF",X"FF",X"00",X"11",X"33",X"66",X"44",X"44",X"77",X"77",X"00",
		X"11",X"99",X"99",X"99",X"FF",X"FF",X"00",X"00",X"44",X"44",X"44",X"44",X"77",X"77",X"00",X"00",
		X"00",X"88",X"88",X"88",X"88",X"FF",X"FF",X"00",X"44",X"44",X"44",X"44",X"44",X"77",X"77",X"00",
		X"00",X"00",X"08",X"0C",X"0E",X"0C",X"08",X"00",X"00",X"07",X"0F",X"0F",X"07",X"0F",X"0F",X"07",
		X"22",X"66",X"44",X"55",X"77",X"55",X"CC",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"11",X"11",X"11",X"33",X"22",X"22",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"22",X"22",X"22",X"33",X"11",X"11",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",
		X"88",X"88",X"CC",X"55",X"77",X"55",X"44",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FB",X"F7",X"DD",X"88",X"00",X"00",X"00",X"00",X"F3",X"F3",X"70",X"30",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"88",X"D9",X"FB",X"00",X"00",X"00",X"00",X"00",X"00",X"41",X"C3",
		X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"00",X"00",X"70",X"03",X"03",X"03",X"CF",X"1F",
		X"88",X"08",X"08",X"08",X"08",X"C0",X"00",X"00",X"FF",X"EF",X"01",X"01",X"10",X"00",X"00",X"00",
		X"CC",X"22",X"22",X"22",X"22",X"EE",X"22",X"00",X"44",X"55",X"55",X"77",X"00",X"77",X"22",X"00",
		X"CC",X"22",X"22",X"CC",X"CC",X"22",X"22",X"CC",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C1",X"EF",X"2E",X"EF",X"C1",X"00",X"00",X"77",X"17",X"DB",X"FF",X"DB",X"17",X"77",X"00",
		X"F0",X"F0",X"70",X"70",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"E4",X"C8",X"C0",X"80",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F3",X"F0",X"E0",X"00",X"00",
		X"00",X"00",X"00",X"80",X"C0",X"C0",X"E0",X"E0",X"00",X"00",X"E0",X"FC",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"30",X"71",X"72",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"DD",X"00",X"EE",X"DD",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"DD",X"00",X"EE",X"DD",X"00",X"00",
		X"22",X"22",X"33",X"00",X"22",X"22",X"22",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"88",X"88",X"00",X"88",X"88",X"88",X"88",X"44",X"44",X"DD",X"00",X"77",X"44",X"44",X"DD",
		X"00",X"00",X"44",X"88",X"EE",X"88",X"44",X"00",X"00",X"00",X"11",X"00",X"33",X"00",X"11",X"00",
		X"00",X"88",X"88",X"88",X"88",X"88",X"00",X"00",X"00",X"22",X"22",X"22",X"22",X"22",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"CC",X"22",X"22",X"66",X"CC",X"88",X"00",X"33",X"77",X"CC",X"88",X"88",X"77",X"33",X"00",
		X"22",X"22",X"EE",X"EE",X"22",X"22",X"00",X"00",X"00",X"00",X"FF",X"FF",X"44",X"00",X"00",X"00",
		X"22",X"22",X"AA",X"AA",X"EE",X"EE",X"66",X"00",X"66",X"FF",X"BB",X"99",X"99",X"CC",X"44",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"66",X"44",X"00",X"88",X"DD",X"FF",X"BB",X"99",X"88",X"00",X"00",
		X"88",X"EE",X"EE",X"88",X"88",X"88",X"88",X"00",X"00",X"FF",X"FF",X"CC",X"66",X"33",X"11",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"66",X"44",X"00",X"11",X"BB",X"AA",X"AA",X"AA",X"EE",X"EE",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"EE",X"CC",X"00",X"00",X"99",X"99",X"99",X"DD",X"77",X"33",X"00",
		X"00",X"00",X"00",X"EE",X"EE",X"00",X"00",X"00",X"CC",X"EE",X"BB",X"99",X"88",X"CC",X"CC",X"00",
		X"CC",X"EE",X"AA",X"AA",X"22",X"22",X"CC",X"00",X"00",X"66",X"99",X"99",X"BB",X"FF",X"66",X"00",
		X"88",X"CC",X"66",X"22",X"22",X"22",X"00",X"00",X"77",X"FF",X"99",X"99",X"99",X"FF",X"66",X"00",
		X"00",X"00",X"00",X"00",X"88",X"44",X"22",X"00",X"88",X"44",X"22",X"11",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"FF",
		X"00",X"00",X"88",X"DD",X"00",X"00",X"00",X"00",X"66",X"99",X"99",X"88",X"88",X"CC",X"66",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"EE",X"88",X"88",X"88",X"EE",X"EE",X"00",X"33",X"77",X"CC",X"88",X"CC",X"77",X"33",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"EE",X"EE",X"00",X"66",X"FF",X"99",X"99",X"99",X"FF",X"FF",X"00",
		X"44",X"66",X"22",X"22",X"66",X"CC",X"88",X"00",X"44",X"CC",X"88",X"88",X"CC",X"77",X"33",X"00",
		X"88",X"CC",X"66",X"22",X"22",X"EE",X"EE",X"00",X"33",X"77",X"CC",X"88",X"88",X"FF",X"FF",X"00",
		X"22",X"22",X"22",X"22",X"EE",X"EE",X"00",X"00",X"88",X"99",X"99",X"99",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"00",X"88",X"99",X"99",X"99",X"99",X"FF",X"FF",X"00",
		X"EE",X"EE",X"22",X"22",X"66",X"CC",X"88",X"00",X"99",X"99",X"99",X"88",X"CC",X"77",X"33",X"00",
		X"EE",X"EE",X"00",X"00",X"00",X"EE",X"EE",X"00",X"FF",X"FF",X"11",X"11",X"11",X"FF",X"FF",X"00",
		X"22",X"22",X"EE",X"EE",X"22",X"22",X"00",X"00",X"88",X"88",X"FF",X"FF",X"88",X"88",X"00",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"66",X"44",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"22",X"66",X"EE",X"CC",X"88",X"EE",X"EE",X"00",X"88",X"CC",X"66",X"33",X"11",X"FF",X"FF",X"00",
		X"22",X"22",X"22",X"22",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"EE",X"EE",X"00",X"88",X"00",X"EE",X"EE",X"00",X"FF",X"FF",X"77",X"33",X"77",X"FF",X"FF",X"00",
		X"EE",X"EE",X"CC",X"88",X"00",X"EE",X"EE",X"00",X"FF",X"FF",X"11",X"33",X"77",X"FF",X"FF",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"EE",X"CC",X"00",X"77",X"FF",X"88",X"88",X"88",X"FF",X"77",X"00",
		X"00",X"88",X"88",X"88",X"88",X"EE",X"EE",X"00",X"77",X"FF",X"88",X"88",X"88",X"FF",X"FF",X"00",
		X"AA",X"CC",X"EE",X"AA",X"22",X"EE",X"CC",X"00",X"77",X"FF",X"88",X"88",X"88",X"FF",X"77",X"00",
		X"22",X"66",X"EE",X"CC",X"88",X"EE",X"EE",X"00",X"77",X"FF",X"99",X"88",X"88",X"FF",X"FF",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"66",X"44",X"00",X"00",X"55",X"DD",X"99",X"99",X"FF",X"66",X"00",
		X"00",X"00",X"EE",X"EE",X"00",X"00",X"00",X"00",X"88",X"88",X"FF",X"FF",X"88",X"88",X"00",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"EE",X"CC",X"00",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"00",
		X"00",X"88",X"CC",X"EE",X"CC",X"88",X"00",X"00",X"FF",X"FF",X"11",X"00",X"11",X"FF",X"FF",X"00",
		X"EE",X"EE",X"CC",X"88",X"CC",X"EE",X"EE",X"00",X"FF",X"FF",X"11",X"33",X"11",X"FF",X"FF",X"00",
		X"66",X"EE",X"CC",X"88",X"CC",X"EE",X"66",X"00",X"CC",X"EE",X"77",X"33",X"77",X"EE",X"CC",X"00",
		X"00",X"00",X"EE",X"EE",X"00",X"00",X"00",X"00",X"EE",X"FF",X"11",X"11",X"FF",X"EE",X"00",X"00",
		X"22",X"22",X"22",X"AA",X"EE",X"EE",X"66",X"00",X"CC",X"EE",X"FF",X"BB",X"99",X"88",X"88",X"00",
		X"00",X"00",X"00",X"00",X"88",X"22",X"00",X"00",X"00",X"CC",X"EE",X"FF",X"33",X"00",X"00",X"00",
		X"F1",X"F3",X"F7",X"EE",X"FC",X"FF",X"FF",X"00",X"00",X"10",X"30",X"70",X"71",X"73",X"33",X"00",
		X"F0",X"F0",X"FF",X"FF",X"00",X"10",X"30",X"70",X"70",X"70",X"73",X"33",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"C0",X"EE",X"EE",X"00",X"CC",X"88",X"00",X"F0",X"F0",X"FF",X"FF",X"00",
		X"80",X"C0",X"EE",X"EE",X"CC",X"88",X"00",X"00",X"F0",X"F0",X"FF",X"FF",X"71",X"F3",X"F7",X"EE",
		X"00",X"00",X"00",X"F0",X"F0",X"FF",X"FF",X"00",X"00",X"00",X"00",X"70",X"70",X"73",X"33",X"00",
		X"F0",X"F0",X"FF",X"FF",X"00",X"00",X"00",X"00",X"70",X"70",X"73",X"33",X"00",X"00",X"00",X"00",
		X"66",X"E6",X"E6",X"EE",X"CC",X"88",X"00",X"00",X"00",X"00",X"10",X"F0",X"F1",X"FF",X"FF",X"00",
		X"00",X"00",X"80",X"C8",X"EC",X"EE",X"66",X"66",X"E0",X"F0",X"FF",X"FF",X"11",X"00",X"00",X"00",
		X"F1",X"F3",X"F7",X"FE",X"FC",X"FF",X"FF",X"00",X"00",X"10",X"30",X"70",X"71",X"73",X"33",X"00",
		X"F0",X"F0",X"FF",X"FF",X"CC",X"EE",X"77",X"73",X"70",X"70",X"73",X"33",X"11",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"C0",X"EE",X"EE",X"00",X"88",X"88",X"00",X"F0",X"F0",X"FF",X"FF",X"00",
		X"80",X"C0",X"EE",X"EE",X"00",X"00",X"00",X"00",X"F0",X"F0",X"FF",X"FF",X"00",X"00",X"00",X"88",
		X"30",X"30",X"30",X"F0",X"F0",X"FF",X"FF",X"00",X"73",X"73",X"73",X"73",X"73",X"73",X"33",X"00",
		X"00",X"C0",X"C0",X"EE",X"FF",X"BB",X"11",X"10",X"00",X"10",X"30",X"70",X"71",X"73",X"73",X"73",
		X"E6",X"E6",X"E6",X"E6",X"E6",X"EE",X"EE",X"00",X"DC",X"DC",X"DC",X"FC",X"FC",X"FF",X"FF",X"00",
		X"00",X"00",X"00",X"88",X"CC",X"EE",X"E6",X"E6",X"00",X"E0",X"F0",X"F3",X"F7",X"FE",X"DC",X"DC",
		X"30",X"30",X"30",X"F0",X"F0",X"FF",X"FF",X"00",X"73",X"73",X"73",X"73",X"73",X"73",X"33",X"00",
		X"00",X"00",X"30",X"30",X"30",X"30",X"30",X"30",X"00",X"60",X"60",X"73",X"73",X"73",X"73",X"73",
		X"E6",X"E6",X"E6",X"E6",X"E6",X"EE",X"EE",X"00",X"DC",X"DC",X"DC",X"FC",X"FC",X"FF",X"FF",X"00",
		X"00",X"80",X"C0",X"E6",X"E6",X"E6",X"E6",X"E6",X"00",X"10",X"10",X"90",X"DC",X"DC",X"DC",X"DC",
		X"71",X"71",X"71",X"F1",X"F1",X"FF",X"FF",X"00",X"73",X"73",X"73",X"73",X"73",X"73",X"33",X"00",
		X"80",X"C0",X"EE",X"FF",X"BB",X"31",X"31",X"31",X"10",X"30",X"70",X"71",X"73",X"73",X"73",X"73",
		X"00",X"00",X"00",X"80",X"C0",X"EE",X"EE",X"00",X"88",X"88",X"88",X"F8",X"F8",X"FF",X"FF",X"00",
		X"00",X"C0",X"E2",X"E6",X"EE",X"CC",X"88",X"00",X"00",X"00",X"10",X"F0",X"F8",X"FF",X"FF",X"88",
		X"00",X"00",X"00",X"F8",X"FC",X"FF",X"77",X"00",X"73",X"73",X"73",X"33",X"11",X"00",X"00",X"00",
		X"00",X"C0",X"E6",X"EE",X"CC",X"88",X"00",X"00",X"00",X"10",X"30",X"70",X"71",X"73",X"73",X"73",
		X"E6",X"E6",X"E6",X"EE",X"CC",X"88",X"00",X"00",X"10",X"10",X"30",X"F0",X"F1",X"FF",X"FF",X"00",
		X"00",X"00",X"00",X"88",X"CC",X"EE",X"E6",X"E6",X"00",X"00",X"33",X"33",X"11",X"10",X"10",X"10",
		X"00",X"00",X"88",X"FC",X"FE",X"77",X"33",X"00",X"73",X"73",X"33",X"11",X"00",X"00",X"00",X"00",
		X"70",X"F0",X"F3",X"F7",X"EE",X"CC",X"88",X"00",X"00",X"00",X"10",X"30",X"70",X"71",X"73",X"73",
		X"00",X"00",X"00",X"C0",X"C0",X"EE",X"EE",X"00",X"F3",X"F3",X"F3",X"F3",X"F3",X"FF",X"FF",X"00",
		X"80",X"C0",X"EE",X"EE",X"00",X"00",X"00",X"00",X"F0",X"F0",X"FF",X"FF",X"F3",X"F3",X"F3",X"F3",
		X"30",X"30",X"30",X"F1",X"FB",X"FF",X"EE",X"00",X"73",X"73",X"73",X"73",X"33",X"11",X"00",X"00",
		X"00",X"00",X"10",X"B8",X"B8",X"30",X"30",X"30",X"00",X"20",X"70",X"71",X"73",X"73",X"73",X"73",
		X"E6",X"E6",X"E6",X"E6",X"E6",X"EE",X"CC",X"00",X"DC",X"DC",X"DC",X"FC",X"B8",X"10",X"00",X"00",
		X"00",X"00",X"00",X"88",X"CC",X"EE",X"E6",X"E6",X"00",X"E0",X"F0",X"F3",X"F7",X"FE",X"DC",X"DC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"22",X"44",X"FF",X"44",X"22",X"00",
		X"E0",X"78",X"78",X"96",X"1E",X"1E",X"FF",X"FF",X"FC",X"CE",X"CE",X"CE",X"DE",X"EF",X"77",X"33",
		X"F3",X"3C",X"3C",X"3C",X"B7",X"7F",X"EE",X"CC",X"70",X"E1",X"E1",X"96",X"87",X"87",X"FF",X"FF",
		X"00",X"AA",X"AA",X"AA",X"AA",X"CC",X"00",X"00",X"00",X"11",X"22",X"22",X"22",X"11",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"11",X"22",X"22",X"11",X"33",X"00",X"00",
		X"71",X"71",X"71",X"F1",X"F1",X"FF",X"FF",X"00",X"00",X"00",X"00",X"70",X"70",X"73",X"33",X"00",
		X"F0",X"F0",X"FF",X"FF",X"71",X"71",X"71",X"71",X"70",X"70",X"73",X"33",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"C0",X"EE",X"EE",X"00",X"88",X"88",X"88",X"F8",X"F8",X"FF",X"FF",X"00",
		X"80",X"C0",X"EE",X"EE",X"00",X"00",X"00",X"00",X"F0",X"F0",X"FF",X"FF",X"88",X"88",X"88",X"88",
		X"D3",X"87",X"97",X"0F",X"2F",X"07",X"00",X"00",X"33",X"10",X"10",X"10",X"00",X"00",X"00",X"00",
		X"0C",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"4F",X"1F",X"0F",X"4F",X"0E",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"00",X"00",X"00",X"08",X"0E",X"8E",X"1F",X"0F",
		X"00",X"00",X"00",X"07",X"4F",X"0F",X"A7",X"87",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",
		X"EF",X"47",X"07",X"07",X"03",X"01",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"0C",X"0C",X"08",X"08",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0E",X"00",X"00",
		X"00",X"00",X"00",X"08",X"08",X"0C",X"0C",X"0C",X"00",X"00",X"0E",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"00",X"00",X"01",X"03",X"87",X"87",X"87",X"47",X"00",X"00",X"00",X"10",X"10",X"30",X"30",X"10",
		X"0F",X"0B",X"0C",X"0F",X"01",X"00",X"00",X"00",X"02",X"01",X"01",X"00",X"00",X"00",X"00",X"00",
		X"68",X"68",X"68",X"68",X"68",X"0C",X"00",X"00",X"0F",X"0F",X"07",X"0C",X"0F",X"03",X"00",X"00",
		X"00",X"00",X"0C",X"68",X"68",X"68",X"6E",X"6E",X"00",X"00",X"03",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"01",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"02",
		X"87",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"10",X"00",X"01",X"01",X"01",X"00",X"00",X"00",
		X"08",X"0C",X"0C",X"08",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"0C",X"0C",X"0C",X"00",X"00",X"0C",X"0F",X"CF",X"2F",X"0F",X"0F",
		X"00",X"00",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"20",
		X"D2",X"63",X"52",X"30",X"00",X"00",X"00",X"00",X"02",X"02",X"04",X"00",X"00",X"00",X"00",X"00",
		X"68",X"84",X"C0",X"80",X"00",X"00",X"00",X"00",X"F5",X"E1",X"5A",X"BE",X"E0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"48",X"84",X"C2",X"E0",X"00",X"00",X"E0",X"B4",X"7C",X"E1",X"5B",X"A5",
		X"00",X"00",X"00",X"30",X"52",X"61",X"F1",X"BC",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"03",
		X"0F",X"0F",X"0D",X"0F",X"0F",X"1E",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"24",X"2C",X"68",X"48",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"48",X"68",X"24",X"2C",
		X"00",X"F0",X"1E",X"0F",X"0D",X"0F",X"0F",X"0D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"F1",X"E0",X"E0",X"00",X"00",X"00",X"00",X"20",X"20",X"10",X"10",X"00",X"00",X"00",X"00",
		X"22",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"DD",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"F1",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"20",
		X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"23",X"33",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"2E",X"EE",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"EE",X"EE",
		X"00",X"00",X"00",X"00",X"11",X"33",X"33",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FD",X"FE",X"FF",X"77",X"33",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"CC",X"CC",X"4C",X"CC",X"00",X"00",X"00",X"FF",X"F7",X"FF",X"F9",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"CC",X"CC",X"CC",X"CC",X"C4",X"00",X"00",X"00",X"FF",X"FF",X"F7",X"FB",X"F9",
		X"00",X"00",X"00",X"33",X"77",X"FE",X"FD",X"FD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",
		X"22",X"66",X"00",X"11",X"08",X"01",X"01",X"01",X"77",X"00",X"04",X"08",X"00",X"01",X"02",X"04",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"00",X"00",X"00",X"33",X"00",X"00",X"33",X"77",X"00",X"00",X"00",
		X"00",X"00",X"00",X"CC",X"48",X"48",X"CC",X"CC",X"00",X"00",X"00",X"FF",X"23",X"FF",X"11",X"71",
		X"00",X"00",X"00",X"55",X"CC",X"C4",X"C9",X"00",X"00",X"00",X"00",X"00",X"11",X"32",X"75",X"75",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"FF",X"F0",X"F0",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"E6",X"E6",X"E6",X"E6",X"00",X"00",X"00",X"00",X"E6",X"E6",X"E6",X"E6",
		X"00",X"00",X"00",X"00",X"E6",X"E6",X"E6",X"E6",X"00",X"00",X"00",X"00",X"E6",X"E6",X"E6",X"E6",
		X"00",X"0E",X"4A",X"6A",X"6A",X"4A",X"0E",X"00",X"00",X"07",X"25",X"65",X"65",X"25",X"07",X"00",
		X"00",X"99",X"CC",X"EE",X"E6",X"E6",X"E6",X"E6",X"00",X"FF",X"FF",X"F0",X"F0",X"FC",X"FE",X"F6",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"FF",X"F0",X"F0",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"F0",X"F0",X"FF",X"FF",X"FF",
		X"00",X"FF",X"FF",X"F0",X"F0",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"F0",X"F0",X"FF",X"FF",X"00",
		X"E6",X"E6",X"E6",X"E6",X"E6",X"E6",X"E6",X"E6",X"76",X"76",X"76",X"76",X"76",X"76",X"76",X"76",
		X"E6",X"E6",X"E6",X"E6",X"E6",X"E6",X"E6",X"E6",X"76",X"76",X"76",X"76",X"76",X"76",X"76",X"E6",
		X"00",X"FF",X"FF",X"F0",X"F0",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"F0",X"F0",X"FF",X"FF",X"00",
		X"E6",X"E6",X"E6",X"E6",X"EE",X"CC",X"88",X"00",X"76",X"FE",X"FC",X"F0",X"F0",X"FF",X"FF",X"00",
		X"00",X"FF",X"FF",X"F0",X"F0",X"F3",X"F7",X"F6",X"00",X"11",X"33",X"77",X"76",X"76",X"76",X"76",
		X"E6",X"E6",X"E6",X"E6",X"EE",X"CC",X"88",X"00",X"76",X"FE",X"FC",X"F0",X"F0",X"FF",X"FF",X"00",
		X"00",X"FF",X"FF",X"F0",X"F0",X"F3",X"F7",X"F6",X"00",X"11",X"33",X"77",X"76",X"76",X"76",X"76",
		X"00",X"FF",X"FF",X"F0",X"F0",X"F3",X"F7",X"F6",X"00",X"11",X"33",X"77",X"76",X"76",X"76",X"76",
		X"00",X"88",X"CC",X"EE",X"E6",X"E6",X"E6",X"E6",X"00",X"FF",X"FF",X"F0",X"F0",X"FC",X"FE",X"76",
		X"E6",X"E6",X"E6",X"E6",X"EE",X"CC",X"88",X"00",X"76",X"FE",X"FC",X"F0",X"F0",X"FF",X"FF",X"00",
		X"E6",X"F7",X"F3",X"F0",X"F0",X"FF",X"FF",X"00",X"76",X"76",X"76",X"76",X"77",X"33",X"11",X"00",
		X"E6",X"F7",X"F3",X"F0",X"F0",X"FF",X"FF",X"00",X"76",X"76",X"76",X"76",X"77",X"33",X"11",X"00",
		X"00",X"88",X"CC",X"EE",X"E6",X"E6",X"E6",X"E6",X"00",X"FF",X"FF",X"F0",X"F0",X"FC",X"FE",X"F6",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"E2",X"E2",X"F1",X"F1",X"F1",X"F1",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F1",X"F1",X"F1",X"F1",X"E2",X"E2",X"CC",X"00",
		X"00",X"33",X"74",X"74",X"F8",X"F8",X"F8",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"F8",X"F8",X"F8",X"74",X"74",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",
		X"00",X"00",X"00",X"00",X"33",X"74",X"F8",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"F8",X"74",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"FF",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"FF",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"E2",X"F1",X"F1",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F1",X"F1",X"E2",X"CC",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"F8",X"F8",X"F9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F9",X"F8",X"F8",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"F1",X"F1",X"F9",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F9",X"F1",X"F1",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"88",X"F7",X"F0",X"F0",X"F0",X"F1",X"F1",X"F1",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F7",X"88",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F1",X"F1",X"F1",
		X"F8",X"F8",X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"11",X"FE",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",X"F0",X"F0",X"F0",X"FE",X"11",X"00",X"00",X"00",
		X"24",X"2C",X"2C",X"24",X"24",X"2C",X"2C",X"24",X"C2",X"C3",X"C3",X"C2",X"C2",X"C3",X"C3",X"C2",
		X"24",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"C2",X"C3",X"C3",X"C3",X"C3",X"C2",X"C2",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"0C",X"22",X"C0",X"C2",X"C2",X"C3",X"C3",X"C3",X"C3",X"C2",
		X"00",X"00",X"00",X"00",X"08",X"0C",X"0C",X"0C",X"0E",X"0E",X"0A",X"0F",X"0F",X"0E",X"0B",X"0F",
		X"0C",X"04",X"0C",X"08",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0D",X"0F",X"0F",X"0E",X"0A",X"0E",
		X"0C",X"0C",X"0C",X"04",X"0C",X"0C",X"0C",X"04",X"0F",X"0F",X"0D",X"0F",X"0F",X"0E",X"0B",X"0F",
		X"3C",X"34",X"3C",X"F0",X"0C",X"0C",X"04",X"0C",X"69",X"69",X"69",X"F0",X"0F",X"0E",X"0B",X"0F",
		X"0C",X"04",X"0C",X"04",X"F0",X"3C",X"3C",X"3C",X"0F",X"0F",X"0D",X"0F",X"F0",X"68",X"69",X"69",
		X"20",X"20",X"20",X"F0",X"00",X"00",X"00",X"00",X"30",X"30",X"30",X"F0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"F0",X"20",X"20",X"20",X"00",X"00",X"00",X"00",X"F0",X"30",X"30",X"30",
		X"80",X"00",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"10",X"00",X"00",X"00",X"11",X"70",X"F0",
		X"97",X"09",X"09",X"96",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"70",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"30",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"F7",X"FF",X"F9",X"F1",X"F3",X"F3",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"10",X"00",X"00",X"00",X"11",X"30",X"30",
		X"97",X"83",X"03",X"96",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"30",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"33",X"41",X"C3",
		X"00",X"00",X"00",X"00",X"00",X"88",X"D9",X"FB",X"00",X"00",X"70",X"03",X"03",X"03",X"CF",X"1F",
		X"88",X"08",X"08",X"08",X"08",X"C0",X"00",X"00",X"F3",X"F3",X"70",X"30",X"00",X"00",X"00",X"00",
		X"FB",X"F7",X"DD",X"88",X"00",X"00",X"00",X"00",X"FF",X"EF",X"01",X"01",X"10",X"00",X"00",X"00",
		X"03",X"03",X"07",X"8F",X"8F",X"8E",X"88",X"88",X"00",X"10",X"32",X"47",X"47",X"67",X"32",X"12",
		X"33",X"B6",X"97",X"1F",X"1F",X"3F",X"B7",X"97",X"CC",X"E6",X"F7",X"F3",X"F9",X"FC",X"FC",X"FD",
		X"88",X"8E",X"8F",X"8F",X"07",X"03",X"03",X"00",X"03",X"47",X"67",X"77",X"33",X"11",X"00",X"00",
		X"1F",X"1F",X"3F",X"FE",X"FF",X"FF",X"33",X"00",X"F9",X"F3",X"F7",X"F7",X"FF",X"EE",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"03",X"0F",X"0F",X"03",X"00",X"12",X"16",X"8F",X"8F",X"CF",X"56",X"16",
		X"FF",X"F4",X"B6",X"3E",X"3F",X"7F",X"F7",X"B7",X"00",X"CC",X"EE",X"F7",X"F3",X"FB",X"F9",X"FB",
		X"03",X"0F",X"0F",X"03",X"00",X"00",X"00",X"00",X"07",X"8F",X"CF",X"FF",X"77",X"33",X"00",X"00",
		X"3F",X"3E",X"7E",X"FC",X"FF",X"FF",X"00",X"00",X"F3",X"F7",X"FF",X"FF",X"EE",X"CC",X"00",X"00",
		X"00",X"00",X"00",X"07",X"87",X"87",X"87",X"00",X"00",X"88",X"88",X"98",X"9A",X"8B",X"47",X"67",
		X"00",X"00",X"00",X"95",X"97",X"1F",X"1F",X"3F",X"00",X"00",X"EE",X"FF",X"F3",X"F9",X"FD",X"FD",
		X"87",X"87",X"87",X"07",X"00",X"00",X"00",X"00",X"FE",X"56",X"47",X"8B",X"89",X"88",X"88",X"00",
		X"B7",X"97",X"1F",X"1F",X"1D",X"00",X"00",X"00",X"FD",X"F9",X"F3",X"FF",X"FF",X"EE",X"00",X"00",
		X"00",X"00",X"03",X"43",X"CB",X"CB",X"8B",X"88",X"00",X"00",X"44",X"88",X"89",X"45",X"23",X"33",
		X"00",X"00",X"00",X"C2",X"C3",X"0F",X"0F",X"1F",X"00",X"00",X"77",X"FF",X"F9",X"FC",X"FE",X"FE",
		X"88",X"88",X"8B",X"CB",X"CB",X"43",X"03",X"00",X"77",X"23",X"23",X"45",X"88",X"88",X"44",X"00",
		X"D3",X"C3",X"0F",X"0F",X"1F",X"00",X"00",X"00",X"FE",X"FE",X"FC",X"F9",X"FF",X"FF",X"77",X"00",
		X"00",X"00",X"00",X"00",X"10",X"1E",X"DE",X"89",X"00",X"00",X"00",X"00",X"73",X"C2",X"C3",X"F3",
		X"00",X"00",X"00",X"00",X"88",X"D9",X"FB",X"FB",X"00",X"00",X"00",X"00",X"00",X"EF",X"1F",X"1F",
		X"1E",X"1E",X"00",X"00",X"00",X"00",X"00",X"00",X"F1",X"F0",X"70",X"00",X"00",X"00",X"00",X"00",
		X"F7",X"DD",X"88",X"00",X"00",X"00",X"00",X"00",X"EF",X"CF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"33",X"41",X"C3",
		X"00",X"00",X"00",X"00",X"00",X"88",X"D9",X"FB",X"00",X"00",X"70",X"03",X"03",X"03",X"CF",X"1F",
		X"88",X"08",X"08",X"08",X"08",X"C0",X"00",X"00",X"F3",X"F3",X"70",X"30",X"00",X"00",X"00",X"00",
		X"FB",X"F7",X"DD",X"88",X"00",X"00",X"00",X"00",X"FF",X"EF",X"01",X"01",X"10",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"77",X"22",X"00",
		X"00",X"00",X"00",X"00",X"30",X"2D",X"0F",X"06",X"00",X"00",X"00",X"00",X"00",X"0C",X"0C",X"0E",
		X"00",X"10",X"3C",X"3C",X"00",X"00",X"00",X"00",X"00",X"31",X"76",X"9B",X"97",X"F3",X"70",X"30",
		X"07",X"47",X"FF",X"F7",X"89",X"C0",X"C0",X"80",X"8E",X"EE",X"EF",X"0B",X"1B",X"CF",X"77",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"AC",X"AC",X"00",X"00",X"00",X"00",X"33",X"11",X"10",X"30",
		X"00",X"00",X"00",X"00",X"0F",X"E7",X"F3",X"F3",X"00",X"00",X"00",X"00",X"08",X"0C",X"77",X"FF",
		X"88",X"8F",X"8F",X"6E",X"4E",X"00",X"00",X"00",X"30",X"30",X"10",X"00",X"00",X"00",X"00",X"00",
		X"F3",X"F3",X"F3",X"E6",X"00",X"00",X"00",X"00",X"FF",X"FF",X"77",X"07",X"03",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"2C",X"2C",X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"70",X"70",
		X"00",X"00",X"00",X"01",X"CD",X"E6",X"F7",X"F7",X"00",X"00",X"00",X"0C",X"0C",X"EF",X"EF",X"EE",
		X"1E",X"1E",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"30",X"10",X"00",X"00",X"00",X"00",X"00",
		X"F7",X"E6",X"CD",X"01",X"00",X"00",X"00",X"00",X"EF",X"EF",X"0C",X"0C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"EE",X"CC",X"1E",X"1E",X"00",X"00",X"00",X"00",X"00",X"31",X"70",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"89",X"DD",X"FF",X"00",X"00",X"00",X"00",X"0F",X"0F",X"EF",X"EF",
		X"00",X"4C",X"4C",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"70",X"31",X"67",X"00",X"00",X"00",
		X"FF",X"FF",X"DD",X"8F",X"0E",X"00",X"00",X"00",X"EE",X"EF",X"EF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"EE",X"11",X"11",X"33",X"EE",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"66",X"44",X"44",X"33",X"11",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"11",X"FF",X"FF",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"77",X"22",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"99",X"DD",X"DD",X"FF",X"77",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"77",X"55",X"44",X"44",X"66",X"22",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"FF",X"99",X"99",X"99",X"33",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"66",X"77",X"55",X"44",X"44",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"FF",X"FF",X"44",X"44",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"77",X"66",X"33",X"11",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"FF",X"11",X"11",X"11",X"33",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"77",X"77",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"FF",X"99",X"99",X"99",X"FF",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"44",X"44",X"66",X"33",X"11",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"88",X"FF",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"77",X"55",X"44",X"44",X"66",X"66",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"77",X"DD",X"DD",X"99",X"99",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"44",X"44",X"55",X"77",X"33",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"EE",X"BB",X"99",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"77",X"44",X"44",X"44",X"77",X"33",X"00",
		X"00",X"CC",X"22",X"22",X"CC",X"00",X"CC",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"88",X"88",X"77",X"00",X"77",X"88",
		X"22",X"CC",X"00",X"CC",X"66",X"22",X"66",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"11",X"33",X"22",X"33",X"11",X"88",X"77",X"00",X"DD",X"22",X"22",X"22",X"88",
		X"00",X"CC",X"22",X"22",X"CC",X"00",X"CC",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"88",X"88",X"77",X"00",X"77",X"88",
		X"22",X"CC",X"00",X"88",X"EE",X"88",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"88",X"77",X"00",X"00",X"FF",X"88",X"44",X"33",
		X"00",X"CC",X"22",X"22",X"CC",X"00",X"CC",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"88",X"88",X"77",X"00",X"77",X"88",
		X"22",X"CC",X"00",X"CC",X"66",X"22",X"22",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"11",X"11",X"11",X"11",X"11",X"88",X"77",X"00",X"33",X"22",X"22",X"22",X"EE",
		X"00",X"CC",X"22",X"22",X"CC",X"00",X"CC",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"88",X"88",X"77",X"00",X"77",X"88",
		X"22",X"CC",X"00",X"CC",X"66",X"22",X"22",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"11",X"11",X"11",X"11",X"00",X"88",X"77",X"00",X"33",X"22",X"22",X"AA",X"FF",
		X"00",X"00",X"00",X"10",X"20",X"D8",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"30",X"70",X"70",X"43",X"06",X"86",X"C3",X"E0",X"C0",X"80",X"C0",X"73",X"77",X"55",X"EE",
		X"CC",X"CC",X"D8",X"20",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C3",X"86",X"06",X"43",X"70",X"70",X"30",X"10",X"EE",X"55",X"77",X"73",X"C0",X"80",X"C0",X"E0",
		X"00",X"00",X"00",X"20",X"40",X"A0",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",
		X"00",X"00",X"30",X"70",X"96",X"03",X"03",X"97",X"00",X"00",X"F0",X"C0",X"E6",X"FF",X"BB",X"DD",
		X"88",X"88",X"A0",X"40",X"20",X"00",X"00",X"00",X"10",X"10",X"10",X"00",X"00",X"00",X"00",X"00",
		X"97",X"03",X"03",X"96",X"70",X"30",X"00",X"00",X"DD",X"BB",X"FF",X"E6",X"C0",X"F0",X"00",X"00",
		X"80",X"00",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"10",X"00",X"00",X"00",X"11",X"70",X"F0",
		X"97",X"09",X"09",X"96",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"70",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"30",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"F7",X"FF",X"F9",X"F1",X"F3",X"F3",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"10",X"00",X"00",X"00",X"11",X"30",X"30",
		X"97",X"83",X"03",X"96",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"30",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"CC",X"6E",X"6E",X"EE",X"EE",X"EE",X"EE",X"00",X"00",X"10",X"10",X"10",X"00",X"00",X"00",
		X"00",X"00",X"87",X"87",X"80",X"00",X"61",X"61",X"00",X"11",X"0F",X"0F",X"33",X"33",X"0F",X"0F",
		X"EE",X"CC",X"E6",X"FB",X"FC",X"FC",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"11",X"30",X"77",X"44",X"44",X"30",X"10",
		X"80",X"08",X"C4",X"E6",X"6E",X"6E",X"6E",X"6E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"03",X"70",X"30",X"23",X"23",X"23",X"23",
		X"EE",X"CC",X"E6",X"FB",X"FC",X"FC",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"11",X"30",X"77",X"47",X"47",X"30",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"30",X"30",
		X"00",X"00",X"00",X"00",X"00",X"F0",X"30",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"30",X"30",X"30",X"F0",X"00",X"00",X"00",
		X"20",X"20",X"20",X"20",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"C0",X"EE",X"EE",X"CC",X"88",X"00",X"00",X"70",X"70",X"73",X"33",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"FF",X"FF",X"00",X"10",X"30",X"70",X"F0",X"F0",X"FF",X"FF",X"71",X"F3",X"F7",X"EE",
		X"00",X"00",X"00",X"80",X"C0",X"EE",X"EE",X"00",X"00",X"10",X"30",X"70",X"71",X"73",X"33",X"00",
		X"F1",X"F3",X"F7",X"EE",X"FC",X"FF",X"FF",X"00",X"CC",X"88",X"00",X"F0",X"F0",X"FF",X"FF",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"88",X"88",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"77",X"77",X"77",X"FF",X"FF",X"FF",
		X"00",X"88",X"88",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"77",X"77",X"77",X"66",
		X"00",X"00",X"88",X"88",X"CC",X"CC",X"CC",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"33",X"33",X"77",X"77",X"FF",
		X"00",X"88",X"CC",X"CC",X"CC",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"77",X"77",X"33",X"33",X"33",X"11",
		X"00",X"00",X"CC",X"EE",X"EE",X"EE",X"EE",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"33",X"77",
		X"88",X"CC",X"EE",X"EE",X"EE",X"EE",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"77",X"33",X"33",X"11",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"44",X"EE",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"77",
		X"CC",X"EE",X"EE",X"EE",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"77",X"33",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",
		X"CC",X"EE",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"33",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"22",X"44",X"11",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"11",X"00",X"00",X"00",X"11",X"99",X"44",X"00",X"00",
		X"00",X"22",X"11",X"88",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"22",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"22",X"22",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
