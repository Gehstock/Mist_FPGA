library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity guzzler_tile_bit1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of guzzler_tile_bit1 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"00",X"07",X"00",X"07",X"00",X"07",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"8E",X"00",X"07",X"00",X"07",X"00",X"07",X"00",
		X"00",X"02",X"03",X"03",X"03",X"03",X"03",X"01",X"00",X"02",X"03",X"03",X"03",X"03",X"03",X"01",
		X"00",X"02",X"03",X"03",X"03",X"03",X"03",X"01",X"00",X"02",X"03",X"03",X"03",X"03",X"03",X"01",
		X"04",X"06",X"03",X"01",X"0E",X"01",X"03",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"06",X"03",X"01",X"0E",X"01",X"03",X"02",
		X"1F",X"3E",X"E7",X"F8",X"08",X"E4",X"1F",X"FF",X"E0",X"78",X"FC",X"1E",X"6E",X"6F",X"0B",X"F9",
		X"F8",X"38",X"7C",X"03",X"1C",X"F0",X"E0",X"3F",X"19",X"69",X"6B",X"0A",X"FE",X"1C",X"38",X"F0",
		X"1F",X"3E",X"E0",X"F0",X"03",X"EC",X"18",X"F8",X"F0",X"38",X"0C",X"FE",X"0E",X"6F",X"6B",X"19",
		X"FF",X"3F",X"74",X"08",X"18",X"F7",X"E0",X"3F",X"F9",X"09",X"6B",X"6A",X"16",X"FC",X"78",X"E0",
		X"FF",X"73",X"D8",X"86",X"03",X"FF",X"3F",X"FF",X"F0",X"F8",X"38",X"1E",X"C7",X"F3",X"FB",X"FB",
		X"FF",X"63",X"07",X"18",X"FC",X"98",X"3F",X"0F",X"F3",X"E3",X"E7",X"C7",X"0E",X"1C",X"F8",X"F0",
		X"00",X"07",X"1E",X"0F",X"FC",X"39",X"0E",X"3F",X"1C",X"C6",X"F3",X"37",X"1C",X"06",X"18",X"C7",
		X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"71",X"3C",X"70",X"06",X"FC",X"1F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"70",X"30",X"08",X"00",X"02",X"00",
		X"81",X"81",X"81",X"81",X"81",X"81",X"FF",X"FF",X"FF",X"FF",X"81",X"81",X"81",X"81",X"81",X"81",
		X"00",X"00",X"06",X"0F",X"3F",X"95",X"70",X"38",X"0D",X"F7",X"1E",X"70",X"39",X"E7",X"03",X"1B",
		X"1C",X"3F",X"0D",X"03",X"00",X"07",X"01",X"00",X"CF",X"81",X"FB",X"A1",X"70",X"F8",X"BF",X"73",
		X"06",X"0F",X"69",X"78",X"5C",X"4C",X"CE",X"E6",X"88",X"DC",X"D4",X"52",X"71",X"31",X"31",X"19",
		X"E7",X"43",X"13",X"37",X"1B",X"19",X"58",X"30",X"19",X"0D",X"8E",X"86",X"84",X"44",X"64",X"38",
		X"30",X"78",X"48",X"4D",X"40",X"60",X"20",X"00",X"00",X"08",X"04",X"04",X"08",X"10",X"10",X"08",
		X"00",X"00",X"00",X"00",X"06",X"06",X"00",X"00",X"00",X"08",X"08",X"08",X"08",X"08",X"00",X"00",
		X"1C",X"3E",X"61",X"41",X"43",X"3E",X"1C",X"00",X"01",X"01",X"7F",X"7F",X"21",X"01",X"00",X"00",
		X"31",X"79",X"59",X"4D",X"4F",X"67",X"23",X"00",X"46",X"6F",X"79",X"59",X"49",X"43",X"02",X"00",
		X"04",X"7F",X"7F",X"64",X"34",X"1C",X"0C",X"00",X"0E",X"5F",X"51",X"51",X"51",X"77",X"76",X"00",
		X"06",X"0F",X"49",X"49",X"69",X"3F",X"1E",X"00",X"60",X"70",X"58",X"4F",X"47",X"40",X"40",X"00",
		X"36",X"4F",X"4D",X"5D",X"59",X"79",X"36",X"00",X"3C",X"7E",X"4B",X"49",X"49",X"78",X"30",X"00",
		X"38",X"44",X"42",X"21",X"42",X"44",X"38",X"00",X"0D",X"26",X"77",X"59",X"4D",X"57",X"22",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3C",X"5A",X"99",X"BD",X"BD",X"99",X"42",X"3C",X"1F",X"3F",X"64",X"44",X"64",X"3F",X"1F",X"00",
		X"36",X"7F",X"49",X"49",X"49",X"7F",X"7F",X"00",X"22",X"63",X"41",X"41",X"63",X"3E",X"1C",X"00",
		X"1C",X"3E",X"63",X"41",X"41",X"7F",X"7F",X"00",X"41",X"49",X"49",X"49",X"49",X"7F",X"7F",X"00",
		X"40",X"48",X"48",X"48",X"48",X"7F",X"7F",X"00",X"4F",X"4F",X"49",X"49",X"63",X"3E",X"1C",X"00",
		X"7F",X"7F",X"08",X"08",X"08",X"7F",X"7F",X"00",X"00",X"41",X"7F",X"7F",X"41",X"00",X"00",X"00",
		X"7E",X"7F",X"01",X"01",X"01",X"03",X"02",X"00",X"41",X"63",X"37",X"1E",X"0C",X"7F",X"7F",X"00",
		X"01",X"01",X"01",X"01",X"01",X"7F",X"7F",X"00",X"7F",X"7F",X"38",X"1C",X"38",X"7F",X"7F",X"00",
		X"7F",X"7F",X"0E",X"1C",X"38",X"7F",X"7F",X"00",X"3E",X"7F",X"41",X"41",X"41",X"7F",X"3E",X"00",
		X"30",X"78",X"48",X"48",X"48",X"7F",X"7F",X"00",X"3D",X"7F",X"46",X"45",X"41",X"7F",X"3E",X"00",
		X"39",X"7B",X"4E",X"44",X"44",X"7F",X"7F",X"00",X"26",X"6F",X"4D",X"59",X"59",X"7B",X"32",X"00",
		X"40",X"40",X"7F",X"7F",X"40",X"40",X"00",X"00",X"7E",X"7F",X"03",X"03",X"03",X"7F",X"7E",X"00",
		X"78",X"7C",X"06",X"03",X"06",X"7C",X"78",X"00",X"7C",X"7F",X"06",X"1C",X"06",X"7F",X"7C",X"00",
		X"63",X"77",X"3E",X"1C",X"3E",X"77",X"63",X"00",X"60",X"78",X"0F",X"0F",X"78",X"60",X"00",X"00",
		X"61",X"71",X"79",X"5D",X"4F",X"47",X"43",X"00",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",
		X"00",X"00",X"01",X"03",X"03",X"07",X"0D",X"08",X"00",X"00",X"80",X"E0",X"30",X"30",X"50",X"70",
		X"0C",X"0E",X"0F",X"05",X"06",X"03",X"00",X"00",X"30",X"10",X"80",X"60",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"05",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"02",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"0E",X"09",X"1A",X"15",X"00",X"07",X"18",X"33",X"2C",X"6B",X"54",X"55",
		X"15",X"1A",X"09",X"0E",X"03",X"00",X"00",X"00",X"55",X"54",X"6B",X"2C",X"33",X"1C",X"07",X"00",
		X"00",X"00",X"03",X"04",X"03",X"00",X"03",X"04",X"00",X"00",X"E0",X"10",X"E0",X"00",X"E0",X"10",
		X"03",X"00",X"00",X"04",X"04",X"07",X"00",X"00",X"E0",X"00",X"60",X"90",X"90",X"A0",X"00",X"00",
		X"00",X"00",X"03",X"04",X"03",X"00",X"03",X"04",X"00",X"00",X"C0",X"20",X"C0",X"00",X"C0",X"20",
		X"03",X"00",X"02",X"05",X"05",X"02",X"00",X"00",X"C0",X"00",X"C0",X"20",X"20",X"C0",X"00",X"00",
		X"03",X"04",X"03",X"00",X"03",X"04",X"03",X"00",X"C0",X"20",X"C0",X"00",X"C0",X"20",X"C0",X"00",
		X"03",X"04",X"03",X"00",X"00",X"07",X"02",X"00",X"C0",X"20",X"C0",X"00",X"20",X"E0",X"20",X"00",
		X"03",X"04",X"03",X"00",X"03",X"04",X"03",X"00",X"C0",X"20",X"C0",X"00",X"C0",X"20",X"C0",X"00",
		X"03",X"04",X"03",X"00",X"03",X"04",X"04",X"02",X"C0",X"20",X"C0",X"00",X"20",X"A0",X"A0",X"60",
		X"03",X"04",X"03",X"00",X"03",X"04",X"03",X"00",X"C0",X"20",X"C0",X"00",X"C0",X"20",X"C0",X"00",
		X"03",X"04",X"03",X"00",X"06",X"05",X"05",X"04",X"C0",X"20",X"C0",X"00",X"C0",X"20",X"20",X"40",
		X"03",X"04",X"03",X"00",X"03",X"04",X"03",X"00",X"C0",X"20",X"C0",X"00",X"C0",X"20",X"C0",X"00",
		X"03",X"04",X"03",X"00",X"00",X"07",X"04",X"03",X"C0",X"20",X"C0",X"00",X"40",X"E0",X"40",X"C0",
		X"03",X"04",X"03",X"00",X"03",X"04",X"03",X"00",X"C0",X"20",X"C0",X"00",X"C0",X"20",X"C0",X"00",
		X"03",X"04",X"03",X"00",X"00",X"05",X"05",X"07",X"C0",X"20",X"C0",X"00",X"C0",X"20",X"20",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3B",X"3E",X"1F",X"0F",X"0F",X"0D",X"1D",X"1F",X"00",X"60",X"C0",X"80",X"C0",X"C0",X"80",X"80",
		X"41",X"8F",X"9F",X"BF",X"FF",X"FF",X"7F",X"7F",X"20",X"38",X"3C",X"3E",X"1A",X"18",X"0C",X"08",
		X"7F",X"31",X"61",X"61",X"BF",X"81",X"40",X"20",X"02",X"06",X"07",X"03",X"02",X"02",X"04",X"00",
		X"00",X"06",X"0F",X"0F",X"1E",X"17",X"00",X"01",X"20",X"38",X"7C",X"FE",X"BE",X"33",X"3A",X"18",
		X"03",X"01",X"09",X"01",X"06",X"02",X"00",X"00",X"98",X"D8",X"9C",X"0D",X"0E",X"2E",X"2C",X"18",
		X"00",X"01",X"03",X"07",X"07",X"0E",X"0E",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"FF",X"E7",X"81",X"3C",X"66",X"C3",X"99",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",
		X"81",X"AF",X"AF",X"EF",X"EB",X"EB",X"CB",X"CB",X"81",X"FD",X"FD",X"FF",X"87",X"87",X"83",X"83",
		X"CB",X"C3",X"C3",X"E7",X"FF",X"BD",X"BD",X"81",X"83",X"83",X"87",X"87",X"FF",X"FD",X"FD",X"81",
		X"81",X"C3",X"C3",X"E3",X"E3",X"F3",X"F3",X"DB",X"81",X"83",X"83",X"83",X"83",X"83",X"83",X"83",
		X"DB",X"CF",X"CF",X"C7",X"C7",X"C3",X"C3",X"81",X"83",X"83",X"83",X"83",X"FF",X"FF",X"FF",X"81",
		X"81",X"C3",X"C3",X"C3",X"C3",X"D3",X"D3",X"D3",X"81",X"B3",X"B3",X"FB",X"FB",X"CF",X"CF",X"CF",
		X"D3",X"D3",X"D3",X"D3",X"FF",X"FF",X"FF",X"81",X"C9",X"C9",X"C9",X"C9",X"FF",X"FF",X"FF",X"81",
		X"50",X"D1",X"D3",X"F7",X"F7",X"7E",X"7E",X"3C",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"50",X"D0",X"D0",X"F0",X"F0",X"70",X"70",X"30",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"00",X"01",X"03",X"06",X"04",X"0C",X"08",X"00",X"7E",X"C7",X"05",X"05",X"05",X"05",X"05",X"05",
		X"00",X"81",X"C3",X"66",X"64",X"7C",X"58",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"00",X"80",X"C0",X"60",X"60",X"70",X"50",X"50",X"50",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"50",
		X"05",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"04",X"04",X"06",X"06",X"06",X"07",X"06",X"06",X"04",X"38",X"20",X"30",X"18",X"0C",X"04",
		X"08",X"64",X"C8",X"90",X"C0",X"60",X"30",X"10",X"20",X"40",X"40",X"20",X"20",X"40",X"40",X"40",
		X"1E",X"21",X"1E",X"00",X"1E",X"21",X"1E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1E",X"21",X"1E",X"00",X"06",X"29",X"29",X"3A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1C",X"39",X"73",X"7F",X"7F",X"3F",X"1F",X"0F",X"00",X"80",X"00",X"70",X"E0",X"C0",X"80",X"80",
		X"0D",X"0D",X"0D",X"0D",X"18",X"18",X"1D",X"1F",X"C0",X"C0",X"E0",X"E0",X"E0",X"C0",X"C0",X"C0",
		X"5F",X"DE",X"FE",X"FE",X"FC",X"FC",X"F8",X"F8",X"FF",X"81",X"81",X"81",X"81",X"81",X"81",X"FF",
		X"3C",X"3F",X"3F",X"3F",X"37",X"21",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"54",X"54",X"54",X"52",X"52",X"52",X"51",X"52",X"52",X"54",X"78",X"60",X"70",X"58",X"5C",X"54",
		X"58",X"74",X"D8",X"90",X"C0",X"60",X"70",X"50",X"60",X"40",X"40",X"60",X"60",X"40",X"40",X"40",
		X"00",X"00",X"1E",X"21",X"1E",X"00",X"1E",X"21",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1E",X"00",X"19",X"25",X"25",X"13",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"1E",X"21",X"1E",X"00",X"1E",X"21",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1E",X"00",X"06",X"29",X"29",X"3A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"1E",X"21",X"1E",X"00",X"1E",X"21",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1E",X"00",X"16",X"29",X"29",X"16",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1E",X"21",X"1E",X"00",X"1E",X"21",X"1E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1E",X"21",X"1E",X"00",X"01",X"3F",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1E",X"21",X"1E",X"00",X"1E",X"21",X"1E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1E",X"21",X"1E",X"00",X"19",X"25",X"25",X"13",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1E",X"21",X"1E",X"00",X"1E",X"21",X"1E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1E",X"21",X"1E",X"00",X"36",X"29",X"29",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1E",X"21",X"1E",X"00",X"1E",X"21",X"1E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1E",X"21",X"1E",X"00",X"02",X"3F",X"22",X"1E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"04",X"3E",X"1F",X"78",X"3C",X"00",X"7F",X"FF",X"71",X"C0",X"E3",X"00",X"F3",
		X"F8",X"70",X"9F",X"79",X"07",X"00",X"00",X"00",X"1F",X"C0",X"80",X"F8",X"9F",X"3F",X"07",X"00",
		X"04",X"FC",X"FC",X"FE",X"FE",X"FE",X"FF",X"06",X"06",X"FC",X"F8",X"E0",X"F0",X"F8",X"FC",X"04",
		X"08",X"FC",X"F8",X"90",X"C0",X"E0",X"E0",X"10",X"20",X"C0",X"C0",X"E0",X"E0",X"C0",X"C0",X"40",
		X"54",X"FC",X"FC",X"FE",X"FE",X"FE",X"FF",X"52",X"52",X"FC",X"F8",X"E0",X"F0",X"F8",X"FC",X"54",
		X"58",X"FC",X"F8",X"90",X"C0",X"E0",X"F0",X"50",X"60",X"C0",X"C0",X"E0",X"E0",X"C0",X"C0",X"40",
		X"00",X"00",X"00",X"30",X"38",X"3C",X"3C",X"3E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3C",X"3C",X"38",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"30",X"78",X"70",X"3B",X"7B",X"7B",X"FB",X"00",X"00",X"00",X"00",X"F8",X"FC",X"FC",X"FC",
		X"FB",X"7B",X"3B",X"70",X"70",X"30",X"00",X"00",X"FC",X"FC",X"F8",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"07",X"1F",X"38",X"27",X"1F",X"38",X"00",X"C0",X"E0",X"F8",X"1C",X"E4",X"F8",X"1C",
		X"27",X"1F",X"3F",X"30",X"07",X"0F",X"07",X"00",X"E4",X"F8",X"FC",X"0C",X"E0",X"B0",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C3",X"00",X"00",X"00",X"00",X"70",X"0C",X"03",X"01",
		X"C7",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"18",X"0F",X"1C",X"06",X"38",X"5C",X"3F",X"8C",X"F8",X"80",X"0F",X"3F",X"1F",X"FF",
		X"70",X"E3",X"EF",X"39",X"67",X"4E",X"00",X"00",X"3F",X"0F",X"99",X"03",X"FA",X"20",X"FF",X"39",
		X"00",X"00",X"03",X"04",X"03",X"00",X"03",X"04",X"00",X"00",X"C0",X"20",X"C0",X"00",X"C0",X"20",
		X"03",X"00",X"03",X"04",X"04",X"02",X"00",X"00",X"C0",X"00",X"20",X"A0",X"A0",X"60",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"81",X"43",X"41",X"01",X"03",X"03",X"00",X"00",X"40",X"C0",X"C0",X"C6",X"86",X"06",X"06",X"02",
		X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"80",X"00",X"0C",X"0C",X"0C",X"1C",X"18",X"18",X"00",
		X"20",X"40",X"80",X"81",X"03",X"03",X"00",X"00",X"00",X"20",X"F0",X"F8",X"A0",X"06",X"06",X"06",
		X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"20",X"06",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"40",X"80",X"81",X"03",X"03",X"00",X"00",X"00",X"00",X"0C",X"CC",X"EC",X"6C",X"E4",X"60",
		X"00",X"00",X"00",X"00",X"00",X"40",X"20",X"18",X"46",X"06",X"06",X"06",X"02",X"00",X"00",X"00",
		X"41",X"83",X"83",X"80",X"80",X"00",X"00",X"00",X"F0",X"F0",X"28",X"18",X"18",X"18",X"18",X"00",
		X"00",X"00",X"00",X"81",X"80",X"83",X"83",X"41",X"00",X"06",X"C6",X"C6",X"C6",X"C2",X"C0",X"80",
		X"11",X"23",X"43",X"80",X"81",X"00",X"00",X"00",X"80",X"C0",X"C2",X"C6",X"C6",X"C6",X"06",X"00",
		X"00",X"00",X"00",X"80",X"80",X"43",X"23",X"11",X"00",X"18",X"18",X"18",X"18",X"28",X"F0",X"F0",
		X"81",X"43",X"41",X"01",X"03",X"03",X"00",X"00",X"40",X"E0",X"F0",X"FE",X"FE",X"FE",X"FE",X"F2",
		X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"80",X"30",X"1C",X"1C",X"3C",X"1C",X"18",X"18",X"00",
		X"20",X"40",X"80",X"81",X"03",X"03",X"00",X"00",X"00",X"E0",X"F0",X"F8",X"F0",X"FE",X"FE",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"20",X"3E",X"12",X"10",X"30",X"00",X"20",X"00",X"00",
		X"20",X"40",X"80",X"81",X"03",X"03",X"00",X"00",X"00",X"E0",X"FC",X"FC",X"FC",X"FC",X"F4",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"40",X"20",X"18",X"7E",X"1E",X"1E",X"3E",X"12",X"20",X"00",X"00",
		X"22",X"43",X"87",X"83",X"03",X"03",X"00",X"00",X"BE",X"FC",X"F8",X"F8",X"F8",X"F8",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"40",X"40",X"5F",X"DF",X"38",X"1E",X"1E",X"3E",X"1E",X"2A",X"E8",X"E8",
		X"41",X"83",X"83",X"80",X"80",X"00",X"00",X"00",X"F0",X"F0",X"F8",X"78",X"78",X"38",X"38",X"70",
		X"00",X"00",X"00",X"81",X"80",X"83",X"83",X"41",X"70",X"3E",X"FE",X"FE",X"FE",X"F2",X"E0",X"80",
		X"21",X"43",X"83",X"80",X"80",X"80",X"80",X"C0",X"F0",X"F0",X"F2",X"7E",X"7E",X"3E",X"3E",X"70",
		X"C0",X"80",X"80",X"80",X"80",X"83",X"43",X"21",X"70",X"3E",X"3E",X"7E",X"7E",X"72",X"F0",X"F0",
		X"11",X"23",X"43",X"80",X"81",X"00",X"00",X"00",X"80",X"E0",X"F2",X"FE",X"FE",X"FE",X"3E",X"70",
		X"00",X"00",X"00",X"80",X"80",X"43",X"23",X"11",X"70",X"38",X"38",X"78",X"78",X"78",X"F0",X"F0",
		X"11",X"23",X"43",X"80",X"80",X"00",X"00",X"00",X"F0",X"F0",X"F3",X"7E",X"7F",X"3F",X"3F",X"7F",
		X"00",X"00",X"00",X"80",X"80",X"43",X"23",X"11",X"7F",X"3F",X"3F",X"7F",X"7E",X"73",X"F0",X"F0",
		X"81",X"47",X"47",X"07",X"07",X"07",X"07",X"07",X"40",X"E0",X"F0",X"FE",X"FE",X"FE",X"FE",X"F2",
		X"07",X"01",X"01",X"01",X"01",X"41",X"40",X"80",X"70",X"7C",X"7C",X"7C",X"7C",X"58",X"18",X"00",
		X"20",X"47",X"87",X"87",X"07",X"07",X"07",X"07",X"00",X"E0",X"F0",X"F8",X"F0",X"FE",X"FE",X"FE",
		X"07",X"01",X"01",X"01",X"01",X"41",X"40",X"20",X"3E",X"32",X"30",X"30",X"30",X"20",X"00",X"00",
		X"20",X"47",X"87",X"87",X"07",X"07",X"07",X"07",X"00",X"E0",X"FC",X"FC",X"FC",X"FC",X"F4",X"F0",
		X"07",X"01",X"01",X"01",X"01",X"41",X"20",X"18",X"7E",X"3E",X"3E",X"3E",X"32",X"20",X"00",X"00",
		X"22",X"47",X"87",X"87",X"07",X"07",X"07",X"07",X"BE",X"FC",X"FC",X"FC",X"F8",X"F8",X"F0",X"F0",
		X"07",X"01",X"01",X"01",X"41",X"41",X"51",X"DF",X"F8",X"FE",X"FE",X"FE",X"FE",X"EA",X"E8",X"E8",
		X"41",X"87",X"87",X"87",X"81",X"01",X"01",X"01",X"F0",X"F0",X"F8",X"F8",X"78",X"78",X"78",X"70",
		X"01",X"01",X"01",X"81",X"87",X"87",X"87",X"41",X"70",X"7E",X"FE",X"FE",X"FE",X"F2",X"E0",X"80",
		X"41",X"87",X"87",X"87",X"81",X"81",X"81",X"C1",X"F0",X"F0",X"FA",X"FE",X"3E",X"3E",X"3E",X"38",
		X"C1",X"81",X"81",X"81",X"87",X"87",X"87",X"41",X"38",X"3E",X"3E",X"3E",X"FE",X"FA",X"F0",X"F0",
		X"11",X"27",X"47",X"87",X"81",X"01",X"01",X"01",X"80",X"E0",X"F2",X"FE",X"FE",X"BE",X"3E",X"38",
		X"01",X"01",X"01",X"81",X"87",X"47",X"27",X"11",X"38",X"3C",X"3C",X"3C",X"FC",X"F4",X"F0",X"F0",
		X"11",X"27",X"47",X"87",X"81",X"01",X"01",X"01",X"F0",X"F0",X"FB",X"FE",X"3F",X"3F",X"3F",X"3F",
		X"01",X"01",X"01",X"81",X"87",X"47",X"27",X"11",X"3F",X"3F",X"3F",X"3F",X"FE",X"FB",X"F0",X"F0",
		X"81",X"4F",X"5F",X"3F",X"7F",X"7F",X"7F",X"7F",X"40",X"E0",X"F0",X"FE",X"FE",X"FE",X"FE",X"F2",
		X"7F",X"31",X"61",X"61",X"31",X"41",X"40",X"80",X"70",X"7C",X"7C",X"7C",X"7C",X"58",X"18",X"00",
		X"20",X"4F",X"9F",X"BF",X"7F",X"7F",X"7F",X"7F",X"00",X"E0",X"F0",X"F8",X"F0",X"FE",X"FE",X"FE",
		X"7F",X"31",X"61",X"61",X"31",X"41",X"40",X"20",X"3E",X"32",X"30",X"30",X"30",X"20",X"00",X"00",
		X"20",X"4F",X"9F",X"BF",X"7F",X"7F",X"7F",X"7F",X"00",X"E0",X"FC",X"FC",X"FC",X"FC",X"F4",X"F0",
		X"7F",X"31",X"61",X"61",X"31",X"41",X"20",X"18",X"7E",X"3E",X"3E",X"3E",X"32",X"20",X"00",X"00",
		X"22",X"4F",X"9F",X"BF",X"7F",X"7F",X"7F",X"7F",X"BE",X"FC",X"FC",X"FC",X"F8",X"F8",X"F0",X"F0",
		X"7F",X"31",X"61",X"61",X"71",X"41",X"51",X"DF",X"F8",X"FE",X"FE",X"FE",X"FE",X"EA",X"E8",X"E8",
		X"41",X"87",X"9F",X"BF",X"B9",X"71",X"71",X"39",X"F0",X"F0",X"F8",X"F8",X"78",X"78",X"78",X"70",
		X"39",X"71",X"71",X"B9",X"BF",X"9F",X"87",X"41",X"70",X"7E",X"FE",X"FE",X"FE",X"F2",X"E0",X"80",
		X"21",X"CF",X"9F",X"BF",X"B1",X"E1",X"E1",X"FF",X"F0",X"F0",X"FA",X"FE",X"3E",X"3E",X"3E",X"38",
		X"FF",X"E1",X"E1",X"B1",X"BF",X"9F",X"CF",X"21",X"38",X"3E",X"3E",X"3E",X"FE",X"FA",X"F0",X"F0",
		X"11",X"27",X"5F",X"BF",X"B1",X"61",X"61",X"31",X"80",X"E0",X"F2",X"FE",X"FE",X"BE",X"3E",X"38",
		X"31",X"61",X"61",X"B1",X"BF",X"5F",X"27",X"11",X"38",X"3C",X"3C",X"3C",X"FC",X"F4",X"F0",X"F0",
		X"11",X"2F",X"5F",X"BF",X"B1",X"61",X"61",X"3F",X"F0",X"F0",X"FB",X"FE",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"61",X"61",X"B1",X"BF",X"5F",X"2F",X"11",X"3F",X"3F",X"3F",X"3F",X"FE",X"FB",X"F0",X"F0",
		X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"E8",X"E8",X"E8",X"E8",X"E8",X"E8",X"E8",X"E8",
		X"5F",X"5F",X"7F",X"7F",X"77",X"23",X"00",X"00",X"E8",X"E8",X"F8",X"F8",X"B8",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"5C",X"7F",X"7F",X"77",X"23",X"00",X"00",X"40",X"E8",X"F8",X"F8",X"B8",X"10",X"00",X"00",
		X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"E8",X"E8",X"E8",X"E8",X"E8",X"E8",X"E8",X"E8",
		X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"E8",X"E8",X"E8",X"E8",X"E8",X"E8",X"E8",X"E8",
		X"00",X"00",X"00",X"00",X"5F",X"5F",X"5F",X"5F",X"00",X"00",X"00",X"00",X"E8",X"E8",X"E8",X"E8",
		X"5F",X"5F",X"7F",X"7F",X"77",X"23",X"00",X"00",X"E8",X"E8",X"F8",X"F8",X"B8",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"5F",X"5F",X"7F",X"7F",X"77",X"23",X"00",X"00",X"E8",X"E8",X"F8",X"F8",X"B8",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"5C",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"40",X"E8",X"E8",X"E8",X"E8",X"E8",X"E8",X"E8",
		X"00",X"1F",X"3C",X"1F",X"0F",X"1F",X"3F",X"3F",X"00",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"1F",X"0F",X"1F",X"3C",X"1F",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"1E",X"3C",X"1E",X"0F",X"1E",X"3C",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1E",X"0F",X"1E",X"3C",X"1E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"00",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"1F",X"3C",X"1F",X"0F",X"1F",X"3F",X"3F",X"00",X"F0",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"1F",X"0F",X"1F",X"3C",X"1F",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"00",X"F0",X"00",X"00",X"00",
		X"00",X"1F",X"3C",X"1F",X"0F",X"1F",X"3F",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"0F",X"1F",X"3C",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FE",X"00",X"FE",X"FF",X"FE",X"FC",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FF",X"FE",X"00",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"1E",X"1C",X"18",X"0F",X"00",X"00",X"00",X"1C",X"3C",X"38",X"10",X"0F",X"18",X"1C",X"0E",
		X"0C",X"0E",X"06",X"03",X"0F",X"06",X"0E",X"0C",X"04",X"06",X"03",X"01",X"0E",X"01",X"03",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"3E",X"3E",X"7E",
		X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7E",X"7E",X"7E",X"7A",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"BA",
		X"E0",X"E0",X"E0",X"00",X"00",X"00",X"00",X"00",X"DA",X"EA",X"DA",X"BA",X"DA",X"EA",X"70",X"00",
		X"00",X"01",X"00",X"01",X"7F",X"7F",X"1E",X"3C",X"00",X"F0",X"70",X"F8",X"FC",X"FC",X"7E",X"BE",
		X"7C",X"1E",X"7E",X"CF",X"1F",X"3F",X"03",X"07",X"3E",X"5E",X"1E",X"3E",X"FE",X"F6",X"C4",X"00",
		X"0F",X"39",X"7F",X"7C",X"FF",X"F8",X"F1",X"FF",X"C0",X"F0",X"F8",X"FC",X"FC",X"FE",X"FE",X"FE",
		X"FF",X"FF",X"7F",X"3F",X"3B",X"73",X"06",X"00",X"FE",X"FE",X"FE",X"FC",X"FC",X"78",X"70",X"E0",
		X"0F",X"38",X"7F",X"79",X"FF",X"F8",X"FC",X"FF",X"C0",X"F0",X"D8",X"CC",X"CE",X"DE",X"7E",X"FE",
		X"FF",X"FF",X"7F",X"7F",X"3F",X"1B",X"13",X"02",X"FE",X"FE",X"FC",X"FC",X"F8",X"60",X"40",X"00",
		X"07",X"1C",X"3F",X"7E",X"7F",X"FC",X"F1",X"FF",X"E0",X"F8",X"EC",X"64",X"E6",X"E6",X"CE",X"9E",
		X"FF",X"FF",X"FF",X"7F",X"7F",X"3D",X"1C",X"0E",X"FE",X"FE",X"FC",X"F8",X"B8",X"9C",X"C0",X"00",
		X"08",X"0D",X"0F",X"2F",X"26",X"3F",X"BF",X"9F",X"00",X"F8",X"FC",X"FE",X"32",X"1B",X"B9",X"C9",
		X"FF",X"FF",X"7F",X"7E",X"3F",X"0F",X"03",X"00",X"C9",X"B9",X"1B",X"32",X"FE",X"FC",X"F8",X"00",
		X"00",X"03",X"0F",X"3F",X"7E",X"7F",X"FF",X"FF",X"00",X"F8",X"FC",X"FE",X"7E",X"3F",X"FF",X"DF",
		X"9F",X"BF",X"3F",X"26",X"2F",X"0F",X"0D",X"08",X"DF",X"FF",X"3F",X"7E",X"FE",X"FC",X"F8",X"00",
		X"01",X"00",X"03",X"1C",X"3F",X"79",X"E3",X"FF",X"C0",X"C2",X"C6",X"E6",X"FE",X"FC",X"F8",X"F8",
		X"FF",X"BF",X"3F",X"7F",X"5F",X"10",X"00",X"00",X"FA",X"FE",X"FC",X"EC",X"C8",X"00",X"00",X"00",
		X"00",X"00",X"03",X"1C",X"3F",X"38",X"71",X"77",X"00",X"04",X"C4",X"EC",X"FC",X"FC",X"F8",X"FA",
		X"FF",X"DF",X"9F",X"3F",X"67",X"4C",X"08",X"00",X"FA",X"FE",X"FE",X"FC",X"E0",X"00",X"00",X"00",
		X"00",X"00",X"04",X"1F",X"38",X"71",X"F7",X"FF",X"00",X"04",X"E4",X"EC",X"FC",X"FC",X"F8",X"F8",
		X"9F",X"3F",X"7F",X"4F",X"0B",X"01",X"00",X"00",X"FA",X"FA",X"FE",X"FE",X"E6",X"82",X"C0",X"00",
		X"00",X"00",X"00",X"03",X"0F",X"04",X"3E",X"9F",X"18",X"38",X"70",X"F2",X"FE",X"7E",X"3E",X"FC",
		X"FF",X"FF",X"7E",X"7C",X"3F",X"0F",X"00",X"00",X"3C",X"FF",X"3F",X"7F",X"F9",X"F1",X"70",X"00",
		X"00",X"00",X"0F",X"1F",X"3C",X"7E",X"3F",X"FF",X"00",X"70",X"F1",X"F9",X"7F",X"3F",X"FF",X"3C",
		X"7F",X"3E",X"7C",X"0F",X"03",X"00",X"00",X"00",X"FC",X"3E",X"7E",X"FE",X"F2",X"70",X"38",X"18",
		X"66",X"8E",X"88",X"40",X"40",X"28",X"10",X"10",X"30",X"38",X"1C",X"0E",X"1E",X"1C",X"00",X"00",
		X"10",X"10",X"28",X"40",X"40",X"88",X"8E",X"66",X"00",X"00",X"1C",X"1E",X"0E",X"1C",X"38",X"30",
		X"00",X"01",X"62",X"72",X"32",X"B1",X"18",X"00",X"B8",X"3C",X"0E",X"06",X"02",X"02",X"00",X"00",
		X"00",X"00",X"51",X"12",X"32",X"3A",X"19",X"00",X"00",X"00",X"02",X"02",X"06",X"0E",X"3C",X"B8",
		X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"00",X"70",X"88",X"34",X"34",X"04",X"88",X"70",X"88",
		X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"34",X"34",X"04",X"88",X"70",X"00",X"00",X"00",
		X"0F",X"04",X"02",X"01",X"01",X"00",X"00",X"00",X"80",X"60",X"10",X"38",X"68",X"F8",X"84",X"F8",
		X"01",X"01",X"02",X"04",X"0F",X"00",X"00",X"00",X"E8",X"38",X"10",X"60",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F8",
		X"3F",X"0F",X"07",X"03",X"00",X"00",X"00",X"00",X"FE",X"FE",X"FE",X"FC",X"F8",X"00",X"00",X"00",
		X"00",X"1C",X"3E",X"70",X"63",X"65",X"2C",X"0C",X"00",X"38",X"7C",X"0E",X"C6",X"E6",X"74",X"10",
		X"0C",X"2C",X"65",X"63",X"70",X"3E",X"1C",X"00",X"10",X"74",X"E6",X"C6",X"0E",X"7C",X"38",X"00",
		X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"60",X"60",X"70",X"30",X"3C",X"1F",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",
		X"00",X"07",X"1F",X"3C",X"30",X"70",X"60",X"60",X"1E",X"3F",X"7F",X"FF",X"FF",X"FF",X"7F",X"1E",
		X"1E",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
