library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity travusa_cpu is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of travusa_cpu is
	type rom is array(0 to  28671) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"F3",X"31",X"80",X"E9",X"ED",X"56",X"3A",X"07",X"71",X"CB",X"47",X"C2",X"E0",X"62",X"C3",X"3C",
		X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"08",X"D9",X"CD",X"EB",X"00",X"CD",X"70",X"00",
		X"D9",X"08",X"FB",X"ED",X"4D",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F5",X"C5",X"D5",X"E5",X"E1",X"D1",X"C1",X"F1",X"ED",X"45",
		X"C3",X"40",X"5E",X"35",X"C0",X"3E",X"02",X"77",X"3A",X"00",X"D0",X"E6",X"08",X"28",X"46",X"3A",
		X"1C",X"E6",X"FE",X"00",X"C8",X"3E",X"00",X"32",X"1C",X"E6",X"21",X"19",X"E6",X"35",X"C0",X"3A",
		X"18",X"E6",X"6F",X"26",X"00",X"11",X"CB",X"00",X"19",X"7E",X"32",X"19",X"E6",X"11",X"10",X"00",
		X"19",X"3A",X"07",X"E2",X"86",X"32",X"07",X"E2",X"C6",X"F6",X"30",X"05",X"3E",X"09",X"32",X"07",
		X"E2",X"3E",X"05",X"CD",X"75",X"22",X"3A",X"F4",X"83",X"FE",X"43",X"C0",X"3A",X"07",X"E2",X"C6",
		X"30",X"32",X"FC",X"83",X"C9",X"3E",X"01",X"32",X"1C",X"E6",X"C9",X"01",X"02",X"03",X"01",X"01",
		X"01",X"01",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"03",
		X"04",X"05",X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"21",X"00",X"E0",X"11",X"20",
		X"C8",X"01",X"60",X"00",X"ED",X"B0",X"1E",X"A0",X"01",X"60",X"00",X"ED",X"B0",X"11",X"20",X"C9",
		X"01",X"60",X"00",X"ED",X"B0",X"1E",X"A0",X"01",X"60",X"00",X"ED",X"B0",X"0E",X"1C",X"7E",X"ED",
		X"79",X"23",X"7E",X"E6",X"7F",X"01",X"40",X"00",X"CB",X"3F",X"30",X"01",X"04",X"20",X"F9",X"7E",
		X"CB",X"07",X"E6",X"01",X"A8",X"5F",X"ED",X"A3",X"3A",X"00",X"88",X"0E",X"80",X"ED",X"A3",X"0E",
		X"60",X"ED",X"A3",X"0E",X"A0",X"ED",X"A3",X"7E",X"2F",X"D3",X"C0",X"C9",X"06",X"20",X"C5",X"21",
		X"00",X"C9",X"06",X"00",X"36",X"00",X"23",X"10",X"FB",X"C1",X"10",X"F2",X"3E",X"01",X"32",X"19",
		X"E6",X"32",X"1B",X"E6",X"3A",X"04",X"D0",X"2F",X"E6",X"0F",X"32",X"18",X"E6",X"6F",X"26",X"00",
		X"11",X"F4",X"5E",X"19",X"7E",X"32",X"19",X"E6",X"3A",X"04",X"D0",X"2F",X"E6",X"F0",X"CB",X"3F",
		X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"32",X"1A",X"E6",X"6F",X"26",X"00",X"19",X"7E",X"00",X"00",
		X"00",X"3E",X"00",X"32",X"07",X"E2",X"3E",X"00",X"32",X"1C",X"E6",X"32",X"1D",X"E6",X"FB",X"21",
		X"00",X"E2",X"11",X"01",X"E2",X"01",X"00",X"02",X"36",X"00",X"ED",X"B0",X"CD",X"61",X"38",X"CD",
		X"F4",X"0D",X"21",X"60",X"E2",X"11",X"61",X"E2",X"36",X"20",X"01",X"12",X"00",X"ED",X"B0",X"3E",
		X"30",X"32",X"65",X"E2",X"32",X"6B",X"E2",X"21",X"FA",X"0D",X"11",X"6C",X"E2",X"01",X"06",X"00",
		X"ED",X"B0",X"21",X"00",X"80",X"11",X"01",X"80",X"01",X"FF",X"07",X"3E",X"20",X"77",X"ED",X"B0",
		X"3A",X"03",X"D0",X"2F",X"E6",X"03",X"C6",X"01",X"32",X"9A",X"E3",X"3A",X"03",X"D0",X"2F",X"E6",
		X"04",X"CB",X"3F",X"CB",X"3F",X"32",X"10",X"E6",X"3A",X"03",X"D0",X"CB",X"3F",X"CB",X"3F",X"CB",
		X"3F",X"CB",X"3F",X"CB",X"3F",X"2F",X"E6",X"07",X"32",X"9B",X"E3",X"CD",X"64",X"3E",X"3E",X"00",
		X"32",X"07",X"E2",X"3E",X"00",X"32",X"2D",X"E3",X"32",X"EB",X"E2",X"CD",X"75",X"3D",X"F5",X"CD",
		X"83",X"0D",X"F1",X"32",X"19",X"E3",X"FE",X"01",X"CA",X"A7",X"03",X"C3",X"1E",X"02",X"3E",X"00",
		X"32",X"41",X"E2",X"32",X"42",X"E2",X"32",X"43",X"E2",X"32",X"13",X"E2",X"3E",X"10",X"32",X"06",
		X"E2",X"3E",X"01",X"32",X"00",X"E2",X"3A",X"9A",X"E3",X"32",X"03",X"E2",X"21",X"57",X"09",X"11",
		X"60",X"E2",X"01",X"06",X"00",X"ED",X"B0",X"21",X"57",X"09",X"11",X"66",X"E2",X"01",X"06",X"00",
		X"ED",X"B0",X"3E",X"00",X"32",X"18",X"E3",X"32",X"01",X"E2",X"CD",X"2B",X"03",X"CD",X"88",X"03",
		X"3E",X"01",X"32",X"00",X"E2",X"CD",X"34",X"04",X"CD",X"2B",X"03",X"3E",X"00",X"32",X"41",X"E2",
		X"32",X"42",X"E2",X"32",X"43",X"E2",X"CD",X"69",X"03",X"3A",X"10",X"E6",X"FE",X"00",X"28",X"05",
		X"3E",X"01",X"32",X"01",X"D0",X"3E",X"02",X"32",X"00",X"E2",X"CD",X"34",X"04",X"CD",X"69",X"03",
		X"3E",X"00",X"32",X"01",X"D0",X"32",X"41",X"E2",X"32",X"42",X"E2",X"32",X"43",X"E2",X"3A",X"23",
		X"E6",X"FE",X"FF",X"28",X"0E",X"CD",X"4A",X"03",X"3E",X"01",X"32",X"00",X"E2",X"CD",X"E7",X"02",
		X"CD",X"2B",X"03",X"3A",X"33",X"E6",X"FE",X"FF",X"28",X"22",X"CD",X"69",X"03",X"3A",X"10",X"E6",
		X"FE",X"00",X"28",X"05",X"3E",X"01",X"32",X"01",X"D0",X"3E",X"02",X"32",X"00",X"E2",X"CD",X"E7",
		X"02",X"3E",X"00",X"32",X"01",X"D0",X"CD",X"88",X"03",X"C3",X"9E",X"02",X"3A",X"23",X"E6",X"FE",
		X"FF",X"C2",X"9E",X"02",X"C3",X"03",X"02",X"CD",X"A0",X"38",X"3E",X"00",X"32",X"13",X"E2",X"32",
		X"41",X"E2",X"32",X"42",X"E2",X"32",X"43",X"E2",X"32",X"31",X"E3",X"32",X"01",X"E2",X"21",X"03",
		X"E2",X"35",X"7E",X"FE",X"FF",X"C0",X"CD",X"B1",X"06",X"3A",X"03",X"D0",X"E6",X"10",X"C4",X"26",
		X"43",X"3A",X"03",X"D0",X"E6",X"10",X"C0",X"CD",X"98",X"3E",X"F5",X"3E",X"00",X"32",X"EB",X"E2",
		X"F1",X"FE",X"00",X"C8",X"3A",X"9A",X"E3",X"32",X"03",X"E2",X"C9",X"3A",X"18",X"E3",X"32",X"20",
		X"E6",X"3A",X"06",X"E2",X"32",X"22",X"E6",X"3A",X"03",X"E2",X"32",X"23",X"E6",X"3A",X"04",X"E2",
		X"32",X"24",X"E6",X"3A",X"2D",X"E3",X"32",X"25",X"E6",X"C9",X"3A",X"20",X"E6",X"32",X"18",X"E3",
		X"3A",X"22",X"E6",X"32",X"06",X"E2",X"3A",X"23",X"E6",X"32",X"03",X"E2",X"3A",X"24",X"E6",X"32",
		X"04",X"E2",X"3A",X"25",X"E6",X"32",X"2D",X"E3",X"C9",X"3A",X"30",X"E6",X"32",X"18",X"E3",X"3A",
		X"32",X"E6",X"32",X"06",X"E2",X"3A",X"33",X"E6",X"32",X"03",X"E2",X"3A",X"34",X"E6",X"32",X"04",
		X"E2",X"3A",X"35",X"E6",X"32",X"2D",X"E3",X"C9",X"3A",X"18",X"E3",X"32",X"30",X"E6",X"3A",X"06",
		X"E2",X"32",X"32",X"E6",X"3A",X"03",X"E2",X"32",X"33",X"E6",X"3A",X"04",X"E2",X"32",X"34",X"E6",
		X"3A",X"2D",X"E3",X"32",X"35",X"E6",X"C9",X"3E",X"00",X"32",X"41",X"E2",X"32",X"42",X"E2",X"32",
		X"43",X"E2",X"32",X"13",X"E2",X"3E",X"10",X"32",X"06",X"E2",X"3E",X"01",X"32",X"00",X"E2",X"3A",
		X"9A",X"E3",X"32",X"03",X"E2",X"21",X"57",X"09",X"11",X"60",X"E2",X"01",X"06",X"00",X"ED",X"B0",
		X"21",X"57",X"09",X"11",X"66",X"E2",X"01",X"06",X"00",X"ED",X"B0",X"3E",X"00",X"32",X"18",X"E3",
		X"32",X"01",X"E2",X"CD",X"D4",X"38",X"3E",X"00",X"32",X"13",X"E2",X"32",X"41",X"E2",X"32",X"42",
		X"E2",X"32",X"43",X"E2",X"32",X"31",X"E3",X"32",X"01",X"E2",X"21",X"03",X"E2",X"35",X"7E",X"FE",
		X"FF",X"20",X"2B",X"CD",X"B1",X"06",X"3A",X"03",X"D0",X"E6",X"10",X"C4",X"26",X"43",X"3A",X"03",
		X"D0",X"E6",X"10",X"C2",X"03",X"02",X"CD",X"98",X"3E",X"F5",X"3E",X"00",X"32",X"EB",X"E2",X"F1",
		X"FE",X"00",X"CA",X"03",X"02",X"3A",X"9A",X"E3",X"32",X"03",X"E2",X"C3",X"2E",X"04",X"CD",X"44",
		X"04",X"C3",X"E6",X"03",X"CD",X"83",X"0D",X"3E",X"00",X"32",X"30",X"E3",X"3E",X"00",X"32",X"83",
		X"E3",X"32",X"84",X"E3",X"3E",X"00",X"32",X"1E",X"E3",X"32",X"1F",X"E3",X"32",X"30",X"E3",X"32",
		X"04",X"E2",X"32",X"05",X"E2",X"3E",X"01",X"32",X"4F",X"E2",X"CD",X"E0",X"3F",X"CD",X"D8",X"34",
		X"CD",X"81",X"34",X"CD",X"1D",X"0B",X"CD",X"C6",X"37",X"3E",X"F0",X"32",X"8B",X"E3",X"3E",X"20",
		X"32",X"8C",X"E3",X"3E",X"02",X"32",X"E5",X"E2",X"32",X"E6",X"E2",X"3E",X"00",X"32",X"87",X"E3",
		X"32",X"1F",X"E3",X"32",X"83",X"E3",X"32",X"84",X"E3",X"CD",X"CA",X"07",X"CD",X"24",X"0C",X"FE",
		X"00",X"20",X"06",X"CD",X"9C",X"04",X"C3",X"5A",X"04",X"3E",X"FF",X"C9",X"01",X"00",X"00",X"11",
		X"00",X"00",X"3E",X"00",X"F5",X"CD",X"64",X"1C",X"F1",X"3C",X"FE",X"18",X"20",X"F6",X"21",X"1E",
		X"E3",X"34",X"21",X"35",X"09",X"CD",X"FB",X"3F",X"3A",X"2D",X"E3",X"C6",X"31",X"32",X"2E",X"82",
		X"3E",X"02",X"11",X"00",X"00",X"1D",X"20",X"FD",X"15",X"20",X"FA",X"3D",X"20",X"F7",X"3A",X"1E",
		X"E3",X"CB",X"27",X"47",X"21",X"F3",X"81",X"CD",X"84",X"33",X"11",X"00",X"08",X"1D",X"20",X"FD",
		X"15",X"20",X"FA",X"10",X"F2",X"11",X"00",X"00",X"1D",X"20",X"FD",X"15",X"20",X"FA",X"3A",X"2D",
		X"E3",X"3C",X"4F",X"57",X"21",X"33",X"82",X"3A",X"1E",X"E3",X"CB",X"27",X"47",X"3E",X"0A",X"CD",
		X"A0",X"33",X"CD",X"84",X"33",X"1E",X"00",X"1D",X"20",X"FD",X"0D",X"20",X"F0",X"4A",X"10",X"ED",
		X"06",X"04",X"11",X"00",X"00",X"1D",X"20",X"FD",X"15",X"20",X"FA",X"10",X"F8",X"21",X"18",X"E3",
		X"34",X"C9",X"3A",X"4E",X"E2",X"FE",X"01",X"C2",X"2D",X"05",X"3E",X"00",X"C9",X"3A",X"10",X"E2",
		X"47",X"3A",X"11",X"E2",X"4F",X"CD",X"7C",X"3A",X"7D",X"3C",X"3C",X"3C",X"E6",X"0F",X"47",X"7D",
		X"E6",X"E0",X"B0",X"6F",X"11",X"20",X"00",X"19",X"7E",X"FE",X"19",X"CA",X"26",X"06",X"3A",X"10",
		X"E2",X"D6",X"08",X"32",X"52",X"E2",X"C6",X"18",X"32",X"54",X"E2",X"3A",X"11",X"E2",X"D6",X"08",
		X"32",X"53",X"E2",X"C6",X"10",X"32",X"55",X"E2",X"DD",X"21",X"84",X"E0",X"06",X"09",X"DD",X"7E",
		X"02",X"FE",X"00",X"C2",X"A4",X"05",X"DD",X"23",X"DD",X"23",X"DD",X"23",X"DD",X"23",X"04",X"78",
		X"FE",X"18",X"C2",X"8E",X"05",X"DD",X"21",X"E4",X"E0",X"06",X"30",X"C3",X"6E",X"05",X"FE",X"34",
		X"C2",X"9C",X"05",X"DD",X"21",X"44",X"E1",X"06",X"40",X"C3",X"6E",X"05",X"FE",X"44",X"C2",X"6E",
		X"05",X"3E",X"00",X"C9",X"DD",X"7E",X"02",X"FE",X"7D",X"CA",X"76",X"05",X"FE",X"7E",X"CA",X"76",
		X"05",X"FE",X"75",X"CA",X"76",X"05",X"FE",X"76",X"CA",X"76",X"05",X"FE",X"77",X"CA",X"76",X"05",
		X"FE",X"78",X"CA",X"76",X"05",X"E6",X"FC",X"FE",X"68",X"CA",X"76",X"05",X"FE",X"6C",X"CA",X"76",
		X"05",X"FE",X"28",X"CA",X"76",X"05",X"FE",X"30",X"CA",X"76",X"05",X"C5",X"DD",X"46",X"03",X"DD",
		X"4E",X"00",X"CD",X"21",X"29",X"C1",X"7A",X"FE",X"00",X"C2",X"76",X"05",X"3E",X"07",X"CD",X"75",
		X"22",X"3E",X"00",X"32",X"1E",X"E3",X"32",X"31",X"E3",X"78",X"E6",X"1F",X"FE",X"04",X"D2",X"03",
		X"06",X"C6",X"09",X"DD",X"46",X"03",X"DD",X"4E",X"00",X"16",X"03",X"1E",X"28",X"C5",X"D5",X"F5",
		X"11",X"00",X"00",X"1D",X"C2",X"13",X"06",X"15",X"C2",X"13",X"06",X"3E",X"07",X"CD",X"75",X"22",
		X"F1",X"D1",X"C1",X"CD",X"64",X"1C",X"3A",X"10",X"E2",X"47",X"3A",X"11",X"E2",X"4F",X"11",X"30",
		X"03",X"3E",X"01",X"CD",X"64",X"1C",X"C5",X"78",X"C6",X"10",X"47",X"3E",X"00",X"CD",X"64",X"1C",
		X"C1",X"2E",X"30",X"C5",X"01",X"00",X"40",X"0D",X"C2",X"47",X"06",X"10",X"FA",X"3E",X"07",X"CD",
		X"75",X"22",X"C1",X"16",X"03",X"2C",X"7D",X"FE",X"34",X"CA",X"75",X"06",X"5D",X"3E",X"01",X"CD",
		X"64",X"1C",X"C5",X"78",X"C6",X"10",X"47",X"3E",X"00",X"CD",X"64",X"1C",X"3E",X"02",X"CD",X"64",
		X"1C",X"C1",X"C3",X"43",X"06",X"11",X"00",X"00",X"01",X"00",X"00",X"2E",X"00",X"7D",X"CD",X"64",
		X"1C",X"2C",X"7D",X"FE",X"18",X"C2",X"7D",X"06",X"3E",X"FF",X"C9",X"45",X"58",X"54",X"45",X"4E",
		X"44",X"45",X"44",X"20",X"50",X"4C",X"41",X"59",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"47",X"41",X"4D",X"45",X"20",X"4F",X"56",X"45",X"52",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"3A",X"80",X"E1",X"F5",X"3E",X"00",X"32",X"80",X"E1",X"21",X"9E",X"06",X"11",X"89",X"81",
		X"01",X"0F",X"00",X"ED",X"B0",X"3E",X"30",X"32",X"EC",X"E2",X"3A",X"EC",X"E2",X"E6",X"02",X"C6",
		X"02",X"21",X"89",X"85",X"11",X"8A",X"85",X"01",X"0F",X"00",X"77",X"ED",X"B0",X"01",X"00",X"10",
		X"0D",X"20",X"FD",X"10",X"FB",X"21",X"EC",X"E2",X"35",X"20",X"DF",X"F1",X"32",X"80",X"E1",X"C9",
		X"3A",X"80",X"E1",X"F5",X"3E",X"00",X"32",X"80",X"E1",X"21",X"8B",X"06",X"11",X"89",X"81",X"01",
		X"0F",X"00",X"ED",X"B0",X"3E",X"20",X"32",X"EC",X"E2",X"3A",X"EC",X"E2",X"E6",X"02",X"C6",X"02",
		X"21",X"89",X"85",X"11",X"8A",X"85",X"01",X"0F",X"00",X"77",X"ED",X"B0",X"01",X"00",X"20",X"0D",
		X"20",X"FD",X"10",X"FB",X"21",X"EC",X"E2",X"35",X"20",X"DF",X"21",X"89",X"81",X"11",X"8A",X"81",
		X"36",X"00",X"01",X"0F",X"00",X"ED",X"B0",X"3E",X"01",X"32",X"EB",X"E2",X"F1",X"32",X"80",X"E1",
		X"CD",X"B7",X"0A",X"CD",X"1E",X"0D",X"C9",X"3E",X"01",X"32",X"19",X"E3",X"32",X"00",X"E2",X"3E",
		X"00",X"32",X"03",X"E2",X"32",X"18",X"E3",X"CD",X"83",X"0D",X"3E",X"00",X"32",X"30",X"E3",X"3E",
		X"00",X"32",X"83",X"E3",X"32",X"84",X"E3",X"3E",X"00",X"32",X"1E",X"E3",X"32",X"1F",X"E3",X"32",
		X"30",X"E3",X"32",X"04",X"E2",X"32",X"05",X"E2",X"3E",X"01",X"32",X"4F",X"E2",X"CD",X"E0",X"3F",
		X"CD",X"46",X"1C",X"E6",X"07",X"32",X"18",X"E3",X"CD",X"83",X"0D",X"CD",X"D8",X"34",X"CD",X"81",
		X"34",X"CD",X"1D",X"0B",X"CD",X"C6",X"37",X"3E",X"F0",X"32",X"8B",X"E3",X"3E",X"20",X"32",X"8C",
		X"E3",X"3E",X"02",X"32",X"E5",X"E2",X"32",X"E6",X"E2",X"3E",X"00",X"32",X"87",X"E3",X"32",X"1F",
		X"E3",X"32",X"83",X"E3",X"32",X"84",X"E3",X"3E",X"01",X"32",X"01",X"E2",X"3E",X"01",X"32",X"41",
		X"E2",X"CD",X"24",X"0C",X"3E",X"00",X"32",X"01",X"E2",X"C9",X"3A",X"90",X"E3",X"47",X"3A",X"18",
		X"E3",X"E6",X"0F",X"80",X"6F",X"26",X"00",X"CB",X"25",X"CB",X"14",X"CB",X"25",X"CB",X"14",X"CB",
		X"25",X"CB",X"14",X"11",X"05",X"08",X"19",X"7E",X"32",X"00",X"E6",X"23",X"7E",X"32",X"01",X"E6",
		X"23",X"7E",X"32",X"02",X"E6",X"23",X"7E",X"32",X"2F",X"E3",X"23",X"7E",X"32",X"E5",X"E2",X"23",
		X"7E",X"32",X"E6",X"E2",X"C9",X"08",X"04",X"04",X"01",X"03",X"03",X"00",X"00",X"08",X"03",X"03",
		X"01",X"03",X"03",X"00",X"00",X"07",X"03",X"02",X"00",X"03",X"03",X"00",X"00",X"07",X"03",X"02",
		X"00",X"02",X"02",X"00",X"00",X"06",X"02",X"02",X"00",X"02",X"02",X"00",X"00",X"06",X"02",X"02",
		X"00",X"02",X"02",X"00",X"00",X"05",X"02",X"02",X"00",X"01",X"01",X"00",X"00",X"05",X"02",X"02",
		X"00",X"01",X"01",X"00",X"00",X"04",X"02",X"02",X"00",X"01",X"01",X"00",X"00",X"04",X"02",X"02",
		X"00",X"02",X"02",X"00",X"00",X"04",X"01",X"02",X"00",X"01",X"01",X"00",X"00",X"04",X"01",X"01",
		X"00",X"01",X"01",X"00",X"00",X"04",X"01",X"01",X"00",X"01",X"01",X"00",X"00",X"04",X"01",X"01",
		X"00",X"01",X"01",X"00",X"00",X"05",X"01",X"02",X"00",X"01",X"01",X"00",X"00",X"05",X"01",X"02",
		X"00",X"01",X"01",X"00",X"00",X"05",X"01",X"02",X"00",X"01",X"01",X"00",X"00",X"05",X"01",X"02",
		X"00",X"01",X"01",X"00",X"00",X"05",X"01",X"02",X"00",X"01",X"01",X"00",X"00",X"05",X"01",X"02",
		X"00",X"01",X"01",X"00",X"00",X"05",X"01",X"02",X"00",X"01",X"01",X"00",X"00",X"05",X"01",X"02",
		X"00",X"01",X"01",X"00",X"00",X"05",X"01",X"02",X"00",X"01",X"01",X"00",X"00",X"05",X"01",X"02",
		X"00",X"01",X"01",X"00",X"00",X"05",X"01",X"02",X"00",X"01",X"01",X"00",X"00",X"05",X"01",X"02",
		X"00",X"01",X"01",X"00",X"00",X"05",X"01",X"02",X"00",X"01",X"01",X"00",X"00",X"05",X"01",X"02",
		X"00",X"01",X"01",X"00",X"00",X"05",X"01",X"02",X"00",X"01",X"01",X"00",X"00",X"05",X"01",X"02",
		X"00",X"01",X"01",X"00",X"00",X"05",X"01",X"02",X"00",X"01",X"01",X"00",X"00",X"05",X"01",X"02",
		X"00",X"01",X"01",X"00",X"00",X"05",X"01",X"02",X"00",X"01",X"01",X"00",X"00",X"05",X"01",X"02",
		X"00",X"01",X"01",X"00",X"00",X"05",X"01",X"02",X"00",X"01",X"01",X"00",X"00",X"05",X"01",X"02",
		X"00",X"01",X"01",X"00",X"00",X"05",X"01",X"02",X"00",X"01",X"01",X"00",X"00",X"05",X"01",X"02",
		X"00",X"01",X"01",X"00",X"00",X"05",X"81",X"EB",X"42",X"4F",X"4E",X"55",X"53",X"20",X"20",X"20",
		X"30",X"30",X"30",X"20",X"20",X"FD",X"82",X"2B",X"20",X"20",X"20",X"31",X"58",X"20",X"20",X"20",
		X"30",X"30",X"30",X"20",X"20",X"FF",X"FF",X"20",X"20",X"20",X"20",X"30",X"30",X"20",X"20",X"20",
		X"CD",X"47",X"0A",X"3A",X"78",X"E2",X"D6",X"04",X"E6",X"1F",X"32",X"78",X"E2",X"3A",X"83",X"E3",
		X"D6",X"28",X"32",X"83",X"E3",X"3A",X"84",X"E3",X"DE",X"00",X"32",X"84",X"E3",X"20",X"0D",X"3E",
		X"00",X"32",X"83",X"E3",X"32",X"84",X"E3",X"3E",X"02",X"32",X"78",X"E2",X"3E",X"00",X"32",X"41",
		X"E2",X"32",X"42",X"E2",X"32",X"43",X"E2",X"32",X"46",X"E2",X"32",X"4A",X"E2",X"32",X"04",X"E2",
		X"32",X"05",X"E2",X"32",X"00",X"E3",X"32",X"10",X"E3",X"3E",X"FF",X"32",X"85",X"E1",X"3E",X"40",
		X"32",X"84",X"E1",X"3E",X"48",X"32",X"83",X"E1",X"3E",X"01",X"32",X"79",X"E2",X"32",X"7A",X"E2",
		X"32",X"7B",X"E2",X"32",X"7C",X"E2",X"32",X"7D",X"E2",X"32",X"80",X"E1",X"32",X"81",X"E1",X"32",
		X"82",X"E1",X"3A",X"18",X"E3",X"E6",X"0F",X"6F",X"26",X"00",X"06",X"05",X"CB",X"25",X"CB",X"14",
		X"10",X"FA",X"11",X"00",X"4E",X"19",X"11",X"80",X"EB",X"01",X"20",X"00",X"ED",X"B0",X"3E",X"00",
		X"32",X"78",X"E2",X"CD",X"23",X"19",X"CD",X"6D",X"19",X"21",X"3C",X"0A",X"11",X"AB",X"81",X"01",
		X"08",X"00",X"ED",X"B0",X"11",X"AB",X"85",X"21",X"AA",X"85",X"36",X"0C",X"01",X"0A",X"00",X"ED",
		X"B0",X"3A",X"19",X"E3",X"FE",X"01",X"28",X"20",X"21",X"78",X"0D",X"11",X"6A",X"81",X"01",X"08",
		X"00",X"ED",X"B0",X"21",X"6A",X"85",X"11",X"6B",X"85",X"36",X"0C",X"01",X"0A",X"00",X"ED",X"B0",
		X"3A",X"00",X"E2",X"C6",X"30",X"32",X"71",X"81",X"CD",X"1E",X"0D",X"C9",X"52",X"45",X"41",X"44",
		X"59",X"21",X"20",X"20",X"20",X"20",X"20",X"3E",X"88",X"32",X"1D",X"E3",X"3E",X"01",X"32",X"12",
		X"E2",X"3E",X"00",X"32",X"14",X"E2",X"3E",X"01",X"32",X"15",X"E2",X"3E",X"00",X"32",X"16",X"E2",
		X"32",X"17",X"E2",X"32",X"18",X"E2",X"32",X"1A",X"E2",X"32",X"1B",X"E2",X"32",X"26",X"E2",X"32",
		X"27",X"E2",X"32",X"28",X"E2",X"32",X"2A",X"E2",X"32",X"2B",X"E2",X"21",X"80",X"E2",X"11",X"81",
		X"E2",X"36",X"00",X"01",X"4F",X"00",X"ED",X"B0",X"3E",X"01",X"32",X"3C",X"E2",X"32",X"3D",X"E2",
		X"32",X"3E",X"E2",X"32",X"3F",X"E2",X"32",X"D1",X"E2",X"32",X"D2",X"E2",X"32",X"D3",X"E2",X"32",
		X"04",X"E3",X"32",X"1E",X"E2",X"32",X"2E",X"E2",X"3E",X"50",X"32",X"40",X"E2",X"3E",X"00",X"32",
		X"01",X"E2",X"3E",X"00",X"32",X"78",X"E2",X"3E",X"00",X"32",X"E0",X"E2",X"32",X"90",X"E3",X"32",
		X"91",X"E3",X"32",X"46",X"E2",X"32",X"4A",X"E2",X"32",X"4E",X"E2",X"32",X"A0",X"E3",X"32",X"B0",
		X"E3",X"32",X"C0",X"E3",X"32",X"D0",X"E3",X"32",X"E8",X"E3",X"32",X"80",X"E2",X"32",X"88",X"E2",
		X"32",X"90",X"E2",X"32",X"98",X"E2",X"32",X"A0",X"E2",X"32",X"A8",X"E2",X"32",X"B0",X"E2",X"32",
		X"B8",X"E2",X"32",X"C0",X"E2",X"32",X"C8",X"E2",X"32",X"10",X"E3",X"32",X"20",X"E3",X"32",X"87",
		X"E3",X"32",X"8A",X"E3",X"32",X"E0",X"E3",X"32",X"E1",X"E3",X"32",X"E2",X"E3",X"32",X"E3",X"E3",
		X"32",X"E4",X"E3",X"32",X"E5",X"E3",X"32",X"E6",X"E3",X"32",X"E7",X"E3",X"C9",X"3E",X"FF",X"32",
		X"85",X"E1",X"3E",X"40",X"32",X"84",X"E1",X"3E",X"48",X"32",X"83",X"E1",X"3E",X"01",X"32",X"79",
		X"E2",X"32",X"7A",X"E2",X"32",X"7B",X"E2",X"32",X"7C",X"E2",X"32",X"7D",X"E2",X"32",X"80",X"E1",
		X"32",X"81",X"E1",X"32",X"82",X"E1",X"3E",X"03",X"32",X"78",X"E2",X"3A",X"18",X"E3",X"E6",X"0F",
		X"6F",X"26",X"00",X"06",X"05",X"CB",X"25",X"CB",X"14",X"10",X"FA",X"11",X"00",X"4E",X"19",X"11",
		X"80",X"EB",X"01",X"20",X"00",X"ED",X"B0",X"3E",X"00",X"32",X"78",X"E2",X"CD",X"23",X"19",X"CD",
		X"6D",X"19",X"21",X"62",X"0D",X"11",X"AB",X"81",X"01",X"08",X"00",X"ED",X"B0",X"11",X"AB",X"85",
		X"21",X"AA",X"85",X"36",X"07",X"01",X"0A",X"00",X"ED",X"B0",X"11",X"EC",X"85",X"21",X"EB",X"85",
		X"36",X"07",X"01",X"0A",X"00",X"ED",X"B0",X"21",X"6D",X"0D",X"11",X"EB",X"81",X"01",X"08",X"00",
		X"ED",X"B0",X"3A",X"18",X"E3",X"CB",X"3F",X"CB",X"3F",X"E6",X"0F",X"C6",X"31",X"32",X"B1",X"81",
		X"3A",X"18",X"E3",X"E6",X"03",X"C6",X"31",X"32",X"F1",X"81",X"3A",X"19",X"E3",X"FE",X"01",X"28",
		X"20",X"21",X"78",X"0D",X"11",X"6A",X"81",X"01",X"08",X"00",X"ED",X"B0",X"21",X"6A",X"85",X"11",
		X"6B",X"85",X"36",X"07",X"01",X"0A",X"00",X"ED",X"B0",X"3A",X"00",X"E2",X"C6",X"30",X"32",X"71",
		X"81",X"3A",X"41",X"E2",X"47",X"3A",X"42",X"E2",X"4F",X"3A",X"43",X"E2",X"C5",X"F5",X"CD",X"47",
		X"0A",X"F1",X"32",X"43",X"E2",X"C1",X"78",X"32",X"41",X"E2",X"79",X"FE",X"01",X"20",X"0A",X"3E",
		X"02",X"32",X"42",X"E2",X"3E",X"0F",X"32",X"00",X"E3",X"CD",X"1E",X"0D",X"3A",X"00",X"E3",X"FE",
		X"00",X"C8",X"3A",X"10",X"E2",X"32",X"01",X"E3",X"3A",X"11",X"E2",X"32",X"02",X"E3",X"3E",X"34",
		X"32",X"03",X"E3",X"C9",X"3E",X"10",X"CD",X"75",X"22",X"CD",X"CA",X"07",X"CD",X"B7",X"2E",X"3E",
		X"EA",X"32",X"D0",X"E2",X"CD",X"68",X"18",X"CD",X"DD",X"1D",X"CD",X"0E",X"1E",X"CD",X"57",X"1E",
		X"CD",X"4F",X"1F",X"CD",X"55",X"20",X"CD",X"89",X"22",X"CD",X"62",X"25",X"CD",X"02",X"27",X"CD",
		X"02",X"27",X"CD",X"3B",X"28",X"CD",X"00",X"2D",X"CD",X"A5",X"2D",X"CD",X"A5",X"2D",X"CD",X"21",
		X"39",X"CD",X"B0",X"39",X"CD",X"C3",X"3A",X"CD",X"04",X"3B",X"CD",X"A5",X"3B",X"CD",X"EC",X"3B",
		X"CD",X"55",X"20",X"CD",X"22",X"3C",X"CD",X"22",X"3C",X"CD",X"3B",X"32",X"CD",X"47",X"17",X"CD",
		X"03",X"18",X"CD",X"5E",X"2D",X"CD",X"1A",X"10",X"CD",X"9D",X"11",X"CD",X"9D",X"11",X"CD",X"95",
		X"0F",X"CD",X"95",X"37",X"CD",X"74",X"21",X"CD",X"CB",X"21",X"CD",X"5C",X"37",X"CD",X"E7",X"36",
		X"CD",X"20",X"37",X"3E",X"01",X"CD",X"01",X"1B",X"CD",X"15",X"17",X"CD",X"33",X"3D",X"CD",X"55",
		X"20",X"CD",X"A5",X"3B",X"01",X"00",X"02",X"0D",X"20",X"FD",X"10",X"FB",X"3A",X"84",X"E3",X"FE",
		X"01",X"20",X"12",X"3A",X"83",X"E3",X"FE",X"40",X"20",X"03",X"3E",X"00",X"C9",X"FE",X"30",X"20",
		X"03",X"C3",X"D5",X"0C",X"00",X"3A",X"01",X"E2",X"FE",X"00",X"28",X"06",X"3A",X"07",X"E2",X"FE",
		X"00",X"C0",X"CD",X"22",X"05",X"FE",X"FF",X"CA",X"F0",X"0C",X"CD",X"56",X"3D",X"C3",X"2C",X"0C",
		X"3A",X"01",X"E2",X"FE",X"00",X"28",X"02",X"E1",X"C9",X"3A",X"03",X"E2",X"FE",X"00",X"20",X"16",
		X"3A",X"06",X"E2",X"E6",X"F0",X"FE",X"00",X"28",X"0D",X"3A",X"EB",X"E2",X"FE",X"01",X"28",X"06",
		X"CD",X"F0",X"06",X"C3",X"2C",X"0C",X"3E",X"11",X"CD",X"75",X"22",X"3E",X"FF",X"C9",X"3E",X"03",
		X"01",X"00",X"00",X"0D",X"20",X"FD",X"05",X"20",X"FA",X"3D",X"20",X"F7",X"3E",X"00",X"32",X"D0",
		X"E2",X"CD",X"B1",X"1C",X"3E",X"06",X"32",X"14",X"E2",X"CD",X"CD",X"1C",X"01",X"00",X"08",X"0D",
		X"20",X"FD",X"10",X"FB",X"3A",X"14",X"E2",X"EE",X"01",X"32",X"14",X"E2",X"3A",X"10",X"E2",X"3C",
		X"32",X"10",X"E2",X"FE",X"80",X"20",X"E2",X"21",X"6A",X"81",X"06",X"00",X"36",X"20",X"23",X"10",
		X"FB",X"C9",X"53",X"54",X"41",X"47",X"45",X"20",X"20",X"20",X"20",X"20",X"20",X"53",X"43",X"45",
		X"4E",X"45",X"20",X"20",X"20",X"20",X"20",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"20",X"20",
		X"20",X"20",X"20",X"3E",X"01",X"32",X"12",X"E2",X"3E",X"00",X"32",X"14",X"E2",X"3E",X"01",X"32",
		X"15",X"E2",X"3E",X"00",X"32",X"16",X"E2",X"32",X"17",X"E2",X"32",X"18",X"E2",X"32",X"1A",X"E2",
		X"32",X"1B",X"E2",X"32",X"26",X"E2",X"32",X"27",X"E2",X"32",X"28",X"E2",X"32",X"2A",X"E2",X"32",
		X"2B",X"E2",X"21",X"80",X"E2",X"11",X"81",X"E2",X"36",X"00",X"01",X"4F",X"00",X"ED",X"B0",X"3E",
		X"01",X"32",X"3C",X"E2",X"32",X"3D",X"E2",X"32",X"3E",X"E2",X"32",X"3F",X"E2",X"32",X"D1",X"E2",
		X"32",X"D2",X"E2",X"32",X"D3",X"E2",X"32",X"04",X"E3",X"32",X"1E",X"E2",X"32",X"2E",X"E2",X"3E",
		X"50",X"32",X"40",X"E2",X"3E",X"00",X"32",X"01",X"E2",X"3E",X"00",X"32",X"78",X"E2",X"3E",X"88",
		X"32",X"1D",X"E3",X"C9",X"3E",X"00",X"32",X"13",X"E2",X"C9",X"35",X"30",X"30",X"30",X"30",X"30",
		X"30",X"3A",X"18",X"E3",X"E6",X"0F",X"6F",X"26",X"00",X"06",X"06",X"CB",X"25",X"CB",X"14",X"10",
		X"FA",X"3A",X"83",X"E3",X"FE",X"D0",X"20",X"00",X"E5",X"3A",X"83",X"E3",X"E6",X"0F",X"FE",X"00",
		X"20",X"19",X"06",X"F0",X"0E",X"C0",X"CD",X"7C",X"3A",X"26",X"81",X"7D",X"E6",X"1F",X"C6",X"40",
		X"6F",X"3E",X"1A",X"77",X"11",X"00",X"04",X"19",X"3E",X"16",X"77",X"E1",X"11",X"52",X"45",X"19",
		X"3A",X"84",X"E3",X"FE",X"00",X"C0",X"3A",X"83",X"E3",X"4F",X"7E",X"FE",X"FF",X"C8",X"B9",X"28",
		X"05",X"23",X"23",X"23",X"18",X"F4",X"23",X"7E",X"FE",X"00",X"20",X"09",X"23",X"7E",X"32",X"85",
		X"E3",X"23",X"C3",X"4A",X"0E",X"FE",X"01",X"20",X"09",X"23",X"7E",X"32",X"80",X"E3",X"23",X"C3",
		X"4A",X"0E",X"FE",X"02",X"20",X"09",X"23",X"7E",X"32",X"81",X"E3",X"23",X"C3",X"4A",X"0E",X"FE",
		X"03",X"20",X"09",X"23",X"7E",X"32",X"82",X"E3",X"23",X"C3",X"4A",X"0E",X"FE",X"04",X"20",X"3D",
		X"23",X"23",X"E5",X"C5",X"3E",X"00",X"32",X"8E",X"E3",X"3A",X"20",X"E3",X"FE",X"00",X"20",X"28",
		X"3E",X"01",X"32",X"20",X"E3",X"3E",X"00",X"32",X"21",X"E3",X"3E",X"04",X"32",X"22",X"E3",X"CD",
		X"46",X"1C",X"E6",X"0C",X"C6",X"50",X"32",X"24",X"E3",X"3E",X"00",X"32",X"25",X"E3",X"CD",X"46",
		X"1C",X"E6",X"03",X"C6",X"02",X"32",X"26",X"E3",X"C1",X"E1",X"C3",X"4A",X"0E",X"FE",X"05",X"20",
		X"09",X"23",X"7E",X"32",X"1D",X"E3",X"23",X"C3",X"4A",X"0E",X"FE",X"06",X"20",X"1C",X"23",X"7E",
		X"32",X"2B",X"E3",X"23",X"3E",X"01",X"32",X"87",X"E3",X"32",X"88",X"E3",X"32",X"89",X"E3",X"3E",
		X"00",X"32",X"8A",X"E3",X"32",X"8D",X"E3",X"C3",X"4A",X"0E",X"FE",X"07",X"20",X"1C",X"23",X"7E",
		X"32",X"2B",X"E3",X"23",X"3E",X"01",X"32",X"87",X"E3",X"32",X"88",X"E3",X"32",X"89",X"E3",X"32",
		X"8D",X"E3",X"3E",X"00",X"32",X"8A",X"E3",X"C3",X"4A",X"0E",X"FE",X"08",X"20",X"3C",X"23",X"E5",
		X"C5",X"3E",X"01",X"32",X"8E",X"E3",X"3A",X"20",X"E3",X"FE",X"00",X"20",X"28",X"3E",X"01",X"32",
		X"20",X"E3",X"3E",X"00",X"32",X"21",X"E3",X"3E",X"04",X"32",X"22",X"E3",X"CD",X"46",X"1C",X"E6",
		X"0C",X"3E",X"50",X"32",X"24",X"E3",X"3E",X"00",X"32",X"25",X"E3",X"CD",X"46",X"1C",X"E6",X"03",
		X"C6",X"02",X"32",X"26",X"E3",X"C1",X"E1",X"C3",X"4A",X"0E",X"FE",X"09",X"20",X"0A",X"23",X"E5",
		X"CD",X"05",X"32",X"E1",X"23",X"C3",X"4A",X"0E",X"FE",X"0A",X"20",X"0A",X"23",X"3E",X"01",X"32",
		X"2F",X"E3",X"23",X"C3",X"4A",X"0E",X"FE",X"0B",X"20",X"0A",X"23",X"3E",X"00",X"32",X"2F",X"E3",
		X"23",X"C3",X"4A",X"0E",X"FE",X"0D",X"20",X"09",X"23",X"7E",X"32",X"2E",X"E3",X"23",X"C3",X"4A",
		X"0E",X"23",X"C3",X"4A",X"0E",X"DD",X"21",X"A0",X"E3",X"3E",X"09",X"32",X"86",X"E3",X"DD",X"7E",
		X"00",X"FE",X"00",X"CA",X"CB",X"0F",X"DD",X"46",X"01",X"DD",X"4E",X"02",X"DD",X"56",X"03",X"DD",
		X"5E",X"04",X"3A",X"86",X"E3",X"CD",X"64",X"1C",X"DD",X"46",X"05",X"DD",X"4E",X"06",X"DD",X"56",
		X"07",X"DD",X"5E",X"08",X"3A",X"86",X"E3",X"3C",X"CD",X"64",X"1C",X"11",X"10",X"00",X"DD",X"19",
		X"3A",X"86",X"E3",X"3C",X"3C",X"32",X"86",X"E3",X"FE",X"0D",X"20",X"0C",X"3A",X"8D",X"E3",X"FE",
		X"00",X"28",X"0A",X"3E",X"11",X"32",X"86",X"E3",X"FE",X"15",X"C2",X"9E",X"0F",X"3A",X"E0",X"E3",
		X"FE",X"00",X"C8",X"DD",X"21",X"E0",X"E3",X"DD",X"46",X"00",X"DD",X"4E",X"01",X"DD",X"56",X"02",
		X"DD",X"5E",X"03",X"3E",X"15",X"CD",X"64",X"1C",X"DD",X"46",X"04",X"DD",X"4E",X"05",X"DD",X"56",
		X"06",X"DD",X"5E",X"07",X"3E",X"16",X"CD",X"64",X"1C",X"C9",X"3A",X"1F",X"E3",X"FE",X"00",X"C0",
		X"21",X"88",X"E3",X"35",X"C0",X"CD",X"46",X"1C",X"E6",X"1F",X"C6",X"02",X"77",X"3A",X"87",X"E3",
		X"FE",X"00",X"C8",X"FE",X"02",X"CA",X"69",X"10",X"3A",X"30",X"E2",X"FE",X"00",X"C0",X"3A",X"34",
		X"E2",X"FE",X"00",X"C0",X"3A",X"38",X"E2",X"FE",X"00",X"C0",X"3A",X"8D",X"E3",X"FE",X"00",X"28",
		X"13",X"DD",X"21",X"80",X"E2",X"06",X"04",X"DD",X"7E",X"00",X"FE",X"00",X"C0",X"11",X"08",X"00",
		X"DD",X"19",X"10",X"F3",X"3E",X"02",X"32",X"87",X"E3",X"DD",X"21",X"A0",X"E3",X"DD",X"7E",X"00",
		X"FE",X"00",X"CA",X"8D",X"10",X"11",X"10",X"00",X"DD",X"19",X"DD",X"E5",X"D1",X"0E",X"E0",X"3A",
		X"8D",X"E3",X"FE",X"00",X"20",X"02",X"0E",X"C0",X"7B",X"B9",X"20",X"E1",X"C9",X"3E",X"03",X"DD",
		X"77",X"0D",X"CD",X"46",X"1C",X"E6",X"01",X"20",X"0A",X"3A",X"11",X"E2",X"C6",X"A0",X"38",X"03",
		X"C3",X"17",X"11",X"3E",X"00",X"DD",X"77",X"0F",X"CD",X"46",X"1C",X"E6",X"03",X"FE",X"00",X"CA",
		X"5C",X"11",X"FE",X"02",X"CA",X"9A",X"11",X"FE",X"01",X"CA",X"17",X"11",X"3E",X"F6",X"DD",X"77",
		X"01",X"DD",X"77",X"05",X"3E",X"50",X"DD",X"77",X"02",X"3E",X"40",X"DD",X"77",X"06",X"3E",X"60",
		X"DD",X"77",X"04",X"3E",X"61",X"DD",X"77",X"08",X"3E",X"00",X"DD",X"77",X"09",X"CD",X"46",X"1C",
		X"E6",X"0F",X"C6",X"08",X"DD",X"77",X"0A",X"3E",X"01",X"DD",X"77",X"0B",X"3E",X"01",X"DD",X"77",
		X"00",X"3E",X"08",X"DD",X"77",X"03",X"DD",X"77",X"07",X"CD",X"46",X"1C",X"E6",X"01",X"C0",X"3A",
		X"8B",X"E3",X"FE",X"00",X"C8",X"3D",X"32",X"8B",X"E3",X"3E",X"09",X"DD",X"77",X"03",X"DD",X"77",
		X"07",X"3E",X"05",X"DD",X"77",X"0D",X"C9",X"3E",X"08",X"DD",X"77",X"01",X"D6",X"0F",X"DD",X"77",
		X"05",X"3A",X"11",X"E2",X"D6",X"10",X"F5",X"CD",X"46",X"1C",X"E6",X"1F",X"47",X"F1",X"80",X"DD",
		X"77",X"02",X"DD",X"77",X"06",X"3E",X"70",X"DD",X"77",X"04",X"3E",X"77",X"DD",X"77",X"08",X"3E",
		X"40",X"DD",X"77",X"09",X"3E",X"01",X"DD",X"77",X"0B",X"3E",X"02",X"DD",X"77",X"00",X"3E",X"00",
		X"DD",X"77",X"0C",X"3E",X"48",X"DD",X"77",X"03",X"DD",X"77",X"07",X"C9",X"3E",X"F0",X"DD",X"77",
		X"01",X"3E",X"00",X"DD",X"77",X"05",X"CD",X"46",X"1C",X"E6",X"7F",X"C6",X"30",X"DD",X"77",X"02",
		X"DD",X"77",X"06",X"3E",X"70",X"DD",X"77",X"04",X"3E",X"77",X"DD",X"77",X"08",X"3E",X"00",X"DD",
		X"77",X"09",X"3E",X"01",X"DD",X"77",X"0B",X"3E",X"02",X"DD",X"77",X"00",X"3E",X"08",X"DD",X"77",
		X"03",X"DD",X"77",X"07",X"3E",X"00",X"DD",X"77",X"0C",X"C9",X"C3",X"BC",X"10",X"21",X"89",X"E3",
		X"35",X"C0",X"3A",X"00",X"E6",X"32",X"89",X"E3",X"DD",X"21",X"A0",X"E3",X"DD",X"7E",X"00",X"FE",
		X"00",X"C2",X"CC",X"11",X"11",X"10",X"00",X"DD",X"19",X"DD",X"E5",X"D1",X"0E",X"E0",X"3A",X"8D",
		X"E3",X"FE",X"00",X"20",X"02",X"0E",X"C0",X"7B",X"B9",X"20",X"E1",X"C9",X"DD",X"7E",X"03",X"E6",
		X"0F",X"47",X"DD",X"7E",X"09",X"B0",X"DD",X"77",X"03",X"DD",X"7E",X"07",X"E6",X"0F",X"47",X"DD",
		X"7E",X"09",X"B0",X"DD",X"77",X"07",X"DD",X"7E",X"00",X"FE",X"01",X"CA",X"BF",X"12",X"FE",X"02",
		X"CA",X"FB",X"13",X"FE",X"03",X"CA",X"5C",X"13",X"FE",X"04",X"CA",X"05",X"12",X"FE",X"05",X"CA",
		X"21",X"12",X"C3",X"B4",X"11",X"DD",X"35",X"0B",X"C2",X"B4",X"11",X"3E",X"02",X"DD",X"77",X"0B",
		X"DD",X"34",X"04",X"DD",X"34",X"08",X"DD",X"7E",X"04",X"FE",X"34",X"C2",X"B4",X"11",X"C3",X"F3",
		X"12",X"DD",X"7E",X"0F",X"FE",X"00",X"28",X"36",X"DD",X"35",X"01",X"DD",X"35",X"01",X"DD",X"35",
		X"01",X"DD",X"34",X"05",X"DD",X"34",X"05",X"DD",X"34",X"05",X"DD",X"35",X"01",X"DD",X"35",X"01",
		X"DD",X"34",X"05",X"DD",X"34",X"05",X"DD",X"35",X"0F",X"DD",X"7E",X"0F",X"E6",X"7F",X"FE",X"00",
		X"C2",X"B4",X"11",X"3E",X"00",X"DD",X"77",X"0F",X"CD",X"B5",X"29",X"C3",X"B4",X"11",X"DD",X"35",
		X"0B",X"C2",X"B4",X"11",X"3E",X"02",X"DD",X"77",X"0B",X"3A",X"E3",X"E3",X"C6",X"02",X"32",X"E3",
		X"E3",X"3A",X"E7",X"E3",X"C6",X"02",X"32",X"E7",X"E3",X"FE",X"71",X"20",X"26",X"3E",X"00",X"32",
		X"E0",X"E3",X"32",X"E4",X"E3",X"32",X"8A",X"E3",X"01",X"00",X"00",X"11",X"00",X"00",X"3E",X"15",
		X"CD",X"64",X"1C",X"3E",X"16",X"CD",X"64",X"1C",X"CD",X"EB",X"29",X"3E",X"03",X"DD",X"77",X"0B",
		X"C3",X"B4",X"11",X"FE",X"6D",X"20",X"10",X"3A",X"E0",X"E3",X"C6",X"10",X"32",X"E0",X"E3",X"3A",
		X"E4",X"E3",X"C6",X"10",X"32",X"E4",X"E3",X"3E",X"03",X"DD",X"77",X"0B",X"C3",X"B4",X"11",X"DD",
		X"7E",X"0F",X"FE",X"00",X"C2",X"D8",X"15",X"DD",X"7E",X"09",X"FE",X"00",X"28",X"14",X"DD",X"7E",
		X"01",X"3C",X"3C",X"DD",X"77",X"01",X"DD",X"77",X"05",X"E6",X"FC",X"FE",X"FC",X"28",X"14",X"C3",
		X"F9",X"12",X"DD",X"7E",X"01",X"3D",X"3D",X"DD",X"77",X"01",X"DD",X"77",X"05",X"E6",X"FC",X"FE",
		X"FC",X"20",X"06",X"CD",X"DC",X"16",X"C3",X"B4",X"11",X"DD",X"35",X"0B",X"20",X"17",X"3E",X"02",
		X"DD",X"77",X"0B",X"DD",X"7E",X"04",X"3C",X"3C",X"FE",X"68",X"20",X"02",X"3E",X"60",X"DD",X"77",
		X"04",X"3C",X"DD",X"77",X"08",X"DD",X"35",X"0A",X"C2",X"B4",X"11",X"DD",X"7E",X"09",X"FE",X"00",
		X"C2",X"47",X"13",X"CD",X"46",X"1C",X"E6",X"01",X"CA",X"47",X"13",X"3E",X"79",X"DD",X"77",X"04",
		X"3E",X"7A",X"DD",X"77",X"08",X"3E",X"03",X"DD",X"77",X"00",X"CD",X"46",X"1C",X"E6",X"0F",X"C6",
		X"01",X"DD",X"77",X"0B",X"C3",X"B4",X"11",X"DD",X"7E",X"09",X"EE",X"40",X"DD",X"77",X"09",X"CD",
		X"46",X"1C",X"E6",X"0F",X"C6",X"08",X"DD",X"77",X"0A",X"C3",X"B4",X"11",X"DD",X"34",X"02",X"DD",
		X"34",X"02",X"DD",X"34",X"06",X"DD",X"34",X"06",X"DD",X"35",X"0B",X"C2",X"B4",X"11",X"CD",X"46",
		X"1C",X"E6",X"07",X"C6",X"02",X"DD",X"77",X"0B",X"DD",X"7E",X"04",X"FE",X"79",X"20",X"1C",X"3E",
		X"7B",X"DD",X"77",X"04",X"3C",X"DD",X"77",X"08",X"DD",X"7E",X"02",X"C6",X"06",X"DD",X"77",X"02",
		X"DD",X"7E",X"06",X"C6",X"06",X"DD",X"77",X"06",X"C3",X"D6",X"13",X"FE",X"7B",X"20",X"1A",X"3E",
		X"72",X"DD",X"77",X"04",X"3E",X"75",X"DD",X"77",X"08",X"DD",X"7E",X"02",X"D6",X"0C",X"DD",X"77",
		X"02",X"D6",X"10",X"DD",X"77",X"06",X"C3",X"D6",X"13",X"3E",X"70",X"DD",X"77",X"04",X"3E",X"77",
		X"DD",X"77",X"08",X"DD",X"7E",X"01",X"C6",X"10",X"DD",X"77",X"05",X"DD",X"7E",X"02",X"DD",X"77",
		X"06",X"3E",X"02",X"DD",X"77",X"00",X"C3",X"B4",X"11",X"3A",X"11",X"E2",X"DD",X"BE",X"02",X"38",
		X"0D",X"DD",X"34",X"02",X"DD",X"34",X"06",X"DD",X"34",X"02",X"DD",X"34",X"06",X"C9",X"DD",X"35",
		X"02",X"DD",X"35",X"06",X"DD",X"35",X"02",X"DD",X"35",X"06",X"C9",X"DD",X"7E",X"0F",X"FE",X"00",
		X"C2",X"3B",X"16",X"DD",X"7E",X"0C",X"FE",X"00",X"C2",X"0B",X"15",X"DD",X"7E",X"03",X"E6",X"0F",
		X"FE",X"09",X"CC",X"D9",X"13",X"DD",X"7E",X"0E",X"FE",X"00",X"28",X"18",X"3A",X"11",X"E2",X"DD",
		X"BE",X"02",X"38",X"08",X"DD",X"34",X"02",X"DD",X"34",X"06",X"18",X"32",X"DD",X"35",X"02",X"DD",
		X"35",X"06",X"18",X"2A",X"DD",X"E5",X"D1",X"7B",X"FE",X"B0",X"28",X"04",X"FE",X"A0",X"20",X"1E",
		X"DD",X"7E",X"00",X"FE",X"02",X"20",X"17",X"DD",X"7E",X"09",X"FE",X"00",X"20",X"10",X"DD",X"7E",
		X"01",X"C6",X"B0",X"DA",X"5E",X"14",X"3E",X"01",X"DD",X"77",X"0C",X"DD",X"77",X"0E",X"DD",X"7E",
		X"03",X"E6",X"0F",X"FE",X"09",X"20",X"3C",X"DD",X"7E",X"0C",X"FE",X"00",X"20",X"35",X"CD",X"46",
		X"1C",X"E6",X"07",X"FE",X"03",X"20",X"2C",X"DD",X"7E",X"09",X"FE",X"00",X"20",X"12",X"DD",X"7E",
		X"01",X"C6",X"B8",X"DA",X"A3",X"14",X"3E",X"01",X"DD",X"77",X"0C",X"DD",X"77",X"0E",X"18",X"13",
		X"3A",X"10",X"E2",X"C6",X"20",X"DD",X"BE",X"01",X"D2",X"A3",X"14",X"3E",X"01",X"DD",X"77",X"0C",
		X"DD",X"77",X"0E",X"DD",X"7E",X"02",X"D6",X"04",X"DD",X"77",X"06",X"DD",X"7E",X"02",X"E6",X"FC",
		X"47",X"3A",X"11",X"E2",X"E6",X"FC",X"B8",X"28",X"10",X"38",X"07",X"3E",X"71",X"DD",X"77",X"04",
		X"18",X"0C",X"3E",X"73",X"DD",X"77",X"04",X"18",X"05",X"3E",X"70",X"DD",X"77",X"04",X"DD",X"7E",
		X"09",X"FE",X"00",X"CA",X"F2",X"14",X"DD",X"7E",X"01",X"3C",X"3C",X"3C",X"3C",X"DD",X"77",X"01",
		X"D6",X"10",X"DD",X"77",X"05",X"DD",X"7E",X"01",X"E6",X"FC",X"FE",X"FC",X"C2",X"0B",X"15",X"C3",
		X"F3",X"12",X"DD",X"7E",X"01",X"3D",X"3D",X"3D",X"3D",X"DD",X"77",X"01",X"C6",X"10",X"DD",X"77",
		X"05",X"DD",X"7E",X"01",X"E6",X"FC",X"FE",X"FC",X"CA",X"F3",X"12",X"DD",X"35",X"0B",X"C2",X"B4",
		X"11",X"DD",X"7E",X"0C",X"FE",X"00",X"C2",X"2E",X"15",X"DD",X"7E",X"08",X"3C",X"FE",X"79",X"20",
		X"02",X"3E",X"77",X"DD",X"77",X"08",X"3E",X"04",X"DD",X"77",X"0B",X"C3",X"B4",X"11",X"DD",X"34",
		X"0C",X"DD",X"7E",X"0C",X"FE",X"02",X"20",X"20",X"3E",X"72",X"DD",X"77",X"04",X"3E",X"75",X"DD",
		X"77",X"08",X"DD",X"7E",X"01",X"DD",X"77",X"05",X"DD",X"7E",X"02",X"D6",X"10",X"DD",X"77",X"06",
		X"3E",X"04",X"DD",X"77",X"0B",X"C3",X"B4",X"11",X"FE",X"03",X"20",X"12",X"3E",X"74",X"DD",X"77",
		X"04",X"3E",X"76",X"DD",X"77",X"08",X"3E",X"04",X"DD",X"77",X"0B",X"C3",X"B4",X"11",X"FE",X"04",
		X"20",X"28",X"3E",X"72",X"DD",X"77",X"04",X"3E",X"75",X"DD",X"77",X"08",X"3E",X"04",X"DD",X"77",
		X"0B",X"DD",X"7E",X"09",X"EE",X"40",X"DD",X"77",X"09",X"DD",X"7E",X"03",X"E6",X"0F",X"DD",X"B6",
		X"09",X"DD",X"77",X"03",X"DD",X"77",X"07",X"C3",X"B4",X"11",X"3E",X"70",X"DD",X"77",X"04",X"3E",
		X"77",X"DD",X"77",X"08",X"3E",X"00",X"DD",X"77",X"0C",X"3E",X"01",X"DD",X"77",X"0B",X"DD",X"7E",
		X"09",X"FE",X"00",X"C2",X"C7",X"15",X"DD",X"7E",X"01",X"C6",X"10",X"DD",X"77",X"05",X"DD",X"7E",
		X"02",X"DD",X"77",X"06",X"C3",X"B4",X"11",X"DD",X"7E",X"01",X"D6",X"10",X"DD",X"77",X"05",X"DD",
		X"7E",X"02",X"DD",X"77",X"06",X"C3",X"B4",X"11",X"DD",X"35",X"0B",X"C2",X"B4",X"11",X"3E",X"02",
		X"DD",X"77",X"0B",X"DD",X"35",X"0F",X"DD",X"7E",X"0F",X"FE",X"80",X"C2",X"B4",X"11",X"3E",X"00",
		X"DD",X"77",X"0F",X"DD",X"7E",X"04",X"FE",X"79",X"20",X"0C",X"3E",X"60",X"DD",X"77",X"04",X"3C",
		X"DD",X"77",X"08",X"C3",X"B4",X"11",X"FE",X"7B",X"20",X"11",X"3E",X"79",X"DD",X"77",X"04",X"3C",
		X"DD",X"77",X"08",X"3E",X"82",X"DD",X"77",X"0F",X"C3",X"B4",X"11",X"FE",X"72",X"20",X"19",X"3E",
		X"7B",X"DD",X"77",X"04",X"3C",X"DD",X"77",X"08",X"DD",X"7E",X"02",X"C6",X"10",X"DD",X"77",X"02",
		X"3E",X"82",X"DD",X"77",X"0F",X"C3",X"B4",X"11",X"C3",X"B4",X"11",X"DD",X"7E",X"09",X"FE",X"00",
		X"CA",X"5F",X"16",X"DD",X"7E",X"01",X"3C",X"3C",X"3C",X"3C",X"DD",X"77",X"01",X"D6",X"10",X"DD",
		X"77",X"05",X"DD",X"7E",X"01",X"E6",X"FC",X"FE",X"FC",X"C2",X"78",X"16",X"C3",X"F3",X"12",X"DD",
		X"7E",X"01",X"3D",X"3D",X"3D",X"3D",X"DD",X"77",X"01",X"C6",X"10",X"DD",X"77",X"05",X"DD",X"7E",
		X"01",X"E6",X"FC",X"FE",X"FC",X"CA",X"F3",X"12",X"DD",X"35",X"0B",X"C2",X"B4",X"11",X"3E",X"02",
		X"DD",X"77",X"0B",X"DD",X"7E",X"0F",X"E6",X"10",X"C2",X"AF",X"16",X"DD",X"7E",X"02",X"C6",X"02",
		X"DD",X"77",X"02",X"DD",X"7E",X"06",X"C6",X"02",X"DD",X"77",X"06",X"DD",X"7E",X"02",X"C6",X"50",
		X"D2",X"A9",X"16",X"CD",X"B5",X"29",X"C3",X"B4",X"11",X"DD",X"35",X"0F",X"C3",X"B4",X"11",X"DD",
		X"34",X"02",X"DD",X"34",X"02",X"DD",X"34",X"06",X"DD",X"34",X"06",X"DD",X"7E",X"02",X"C6",X"E0",
		X"DA",X"C9",X"16",X"CD",X"B5",X"29",X"C3",X"B4",X"11",X"DD",X"35",X"0F",X"DD",X"7E",X"0F",X"FE",
		X"10",X"C2",X"B4",X"11",X"3E",X"00",X"DD",X"77",X"0F",X"C3",X"B4",X"11",X"DD",X"E5",X"D1",X"7B",
		X"D6",X"A0",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"6F",X"26",X"00",X"11",X"11",X"17",
		X"19",X"06",X"0F",X"3E",X"00",X"DD",X"E5",X"DD",X"77",X"00",X"DD",X"23",X"10",X"F9",X"DD",X"E1",
		X"7E",X"F5",X"01",X"00",X"00",X"11",X"00",X"00",X"CD",X"64",X"1C",X"F1",X"3C",X"CD",X"64",X"1C",
		X"C9",X"09",X"0B",X"11",X"13",X"DD",X"21",X"A0",X"E3",X"06",X"04",X"DD",X"7E",X"00",X"FE",X"00",
		X"28",X"1D",X"FE",X"05",X"28",X"19",X"DD",X"7E",X"09",X"FE",X"00",X"20",X"12",X"DD",X"35",X"01",
		X"DD",X"35",X"05",X"DD",X"7E",X"01",X"C5",X"E6",X"FC",X"FE",X"FC",X"CC",X"DC",X"16",X"C1",X"11",
		X"10",X"00",X"DD",X"19",X"10",X"D5",X"C9",X"3A",X"2F",X"E3",X"FE",X"01",X"C8",X"3A",X"E0",X"E2",
		X"FE",X"00",X"C0",X"3A",X"87",X"E3",X"FE",X"02",X"C0",X"21",X"E7",X"E2",X"35",X"C0",X"3A",X"E5",
		X"E2",X"77",X"DD",X"21",X"A0",X"E3",X"DD",X"7E",X"00",X"FE",X"02",X"20",X"30",X"DD",X"7E",X"02",
		X"E6",X"C0",X"47",X"3A",X"11",X"E2",X"E6",X"C0",X"B8",X"20",X"22",X"DD",X"7E",X"09",X"FE",X"00",
		X"20",X"0E",X"DD",X"7E",X"01",X"47",X"3A",X"10",X"E2",X"B8",X"D2",X"9D",X"17",X"C3",X"B1",X"17",
		X"DD",X"7E",X"01",X"47",X"3A",X"10",X"E2",X"B8",X"38",X"03",X"C3",X"B1",X"17",X"11",X"10",X"00",
		X"DD",X"19",X"DD",X"E5",X"D1",X"7B",X"FE",X"C0",X"C2",X"66",X"17",X"3E",X"04",X"32",X"E7",X"E2",
		X"C9",X"DD",X"7E",X"09",X"FE",X"00",X"28",X"15",X"DD",X"7E",X"01",X"C6",X"08",X"32",X"E2",X"E2",
		X"3E",X"43",X"32",X"E4",X"E2",X"3E",X"01",X"32",X"E1",X"E2",X"C3",X"DF",X"17",X"DD",X"7E",X"01",
		X"D6",X"08",X"32",X"E2",X"E2",X"3E",X"03",X"32",X"E4",X"E2",X"3E",X"00",X"32",X"E1",X"E2",X"DD",
		X"7E",X"02",X"32",X"E3",X"E2",X"3E",X"04",X"32",X"E8",X"E2",X"3E",X"01",X"32",X"E0",X"E2",X"3A",
		X"E2",X"E2",X"47",X"3A",X"E3",X"E2",X"4F",X"3A",X"E4",X"E2",X"57",X"1E",X"4C",X"3E",X"10",X"CD",
		X"64",X"1C",X"C9",X"DD",X"21",X"E0",X"E2",X"DD",X"7E",X"00",X"FE",X"00",X"C8",X"DD",X"35",X"08",
		X"C0",X"DD",X"7E",X"06",X"DD",X"77",X"08",X"DD",X"7E",X"01",X"FE",X"00",X"20",X"25",X"DD",X"35",
		X"02",X"DD",X"35",X"02",X"DD",X"35",X"02",X"DD",X"35",X"02",X"DD",X"7E",X"02",X"E6",X"FC",X"FE",
		X"FC",X"20",X"25",X"3E",X"00",X"DD",X"77",X"00",X"01",X"00",X"00",X"11",X"00",X"00",X"3E",X"10",
		X"C3",X"64",X"1C",X"DD",X"34",X"02",X"DD",X"34",X"02",X"DD",X"34",X"02",X"DD",X"34",X"02",X"DD",
		X"7E",X"02",X"E6",X"FC",X"FE",X"FC",X"28",X"DB",X"DD",X"46",X"02",X"DD",X"4E",X"03",X"DD",X"56",
		X"04",X"1E",X"4D",X"3E",X"10",X"C3",X"64",X"1C",X"DD",X"E5",X"E5",X"C5",X"21",X"08",X"E2",X"01",
		X"00",X"06",X"71",X"23",X"10",X"FC",X"3E",X"00",X"32",X"11",X"E6",X"32",X"12",X"E6",X"3A",X"00",
		X"D0",X"CB",X"3F",X"38",X"05",X"3E",X"01",X"32",X"11",X"E6",X"CB",X"3F",X"38",X"05",X"3E",X"01",
		X"32",X"12",X"E6",X"3A",X"01",X"E2",X"FE",X"00",X"C2",X"EE",X"18",X"3A",X"00",X"E2",X"FE",X"01",
		X"28",X"12",X"3A",X"03",X"D0",X"E6",X"04",X"EE",X"04",X"28",X"09",X"DD",X"21",X"08",X"E2",X"3A",
		X"02",X"D0",X"18",X"07",X"DD",X"21",X"08",X"E2",X"3A",X"01",X"D0",X"CB",X"3F",X"38",X"03",X"DD",
		X"34",X"05",X"CB",X"3F",X"38",X"03",X"DD",X"34",X"04",X"CB",X"3F",X"38",X"03",X"DD",X"34",X"03",
		X"CB",X"3F",X"38",X"03",X"DD",X"34",X"02",X"CB",X"3F",X"38",X"03",X"DD",X"34",X"01",X"CB",X"3F",
		X"CB",X"3F",X"CB",X"3F",X"38",X"03",X"DD",X"34",X"00",X"C1",X"E1",X"DD",X"E1",X"C9",X"21",X"9F",
		X"E3",X"7E",X"E6",X"01",X"32",X"08",X"E2",X"3A",X"9E",X"E3",X"FE",X"00",X"20",X"07",X"3E",X"01",
		X"32",X"0A",X"E2",X"18",X"09",X"FE",X"01",X"20",X"05",X"3E",X"01",X"32",X"0B",X"E2",X"35",X"20",
		X"0D",X"CD",X"46",X"1C",X"E6",X"0F",X"C6",X"02",X"77",X"2B",X"7E",X"EE",X"01",X"77",X"C1",X"E1",
		X"DD",X"E1",X"C9",X"3A",X"78",X"E2",X"3D",X"3D",X"E6",X"1F",X"F6",X"80",X"6F",X"26",X"EB",X"06",
		X"08",X"11",X"00",X"EC",X"7E",X"CD",X"46",X"19",X"23",X"7D",X"E6",X"1F",X"F6",X"80",X"6F",X"7B",
		X"C6",X"08",X"5F",X"10",X"EF",X"C9",X"E5",X"D5",X"C5",X"67",X"2E",X"00",X"CB",X"3C",X"CB",X"1D",
		X"CB",X"3C",X"CB",X"1D",X"01",X"00",X"50",X"09",X"06",X"08",X"C5",X"01",X"08",X"00",X"ED",X"B0",
		X"01",X"38",X"00",X"EB",X"09",X"EB",X"C1",X"10",X"F1",X"C1",X"D1",X"E1",X"C9",X"21",X"06",X"1C",
		X"11",X"00",X"81",X"01",X"40",X"00",X"ED",X"B0",X"21",X"00",X"85",X"06",X"40",X"36",X"A0",X"23",
		X"10",X"FB",X"26",X"EC",X"3A",X"79",X"E2",X"6F",X"11",X"00",X"83",X"06",X"08",X"E5",X"D5",X"C5",
		X"01",X"20",X"00",X"ED",X"B0",X"C1",X"D1",X"E1",X"C5",X"EB",X"01",X"20",X"00",X"09",X"EB",X"01",
		X"40",X"00",X"09",X"C1",X"10",X"E7",X"26",X"EE",X"3A",X"79",X"E2",X"6F",X"21",X"00",X"83",X"11",
		X"00",X"87",X"06",X"00",X"7E",X"CD",X"80",X"1A",X"12",X"23",X"13",X"10",X"01",X"C9",X"C3",X"B4",
		X"19",X"E5",X"D5",X"C5",X"47",X"3A",X"7C",X"E2",X"80",X"4F",X"E6",X"01",X"32",X"7C",X"E2",X"79",
		X"CB",X"3F",X"4F",X"3A",X"81",X"E1",X"81",X"32",X"81",X"E1",X"3A",X"7D",X"E2",X"80",X"4F",X"E6",
		X"03",X"32",X"7D",X"E2",X"79",X"CB",X"3F",X"CB",X"3F",X"4F",X"3A",X"82",X"E1",X"81",X"32",X"82",
		X"E1",X"3A",X"7B",X"E2",X"80",X"47",X"E6",X"07",X"32",X"7B",X"E2",X"78",X"CB",X"3F",X"CB",X"3F",
		X"CB",X"3F",X"20",X"0F",X"3A",X"7A",X"E2",X"47",X"3A",X"7B",X"E2",X"80",X"32",X"80",X"E1",X"C1",
		X"D1",X"E1",X"C9",X"47",X"CB",X"20",X"CB",X"20",X"CB",X"20",X"3A",X"7A",X"E2",X"80",X"32",X"7A",
		X"E2",X"3A",X"79",X"E2",X"3D",X"32",X"79",X"E2",X"FE",X"FF",X"20",X"12",X"3A",X"78",X"E2",X"3D",
		X"3D",X"E6",X"7F",X"32",X"78",X"E2",X"3E",X"0F",X"32",X"79",X"E2",X"CD",X"23",X"19",X"3A",X"7A",
		X"E2",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"6F",X"3E",X"1F",X"95",X"3C",X"E6",X"1F",X"6F",X"26",
		X"83",X"3A",X"79",X"E2",X"5F",X"16",X"EC",X"E5",X"06",X"08",X"1A",X"77",X"C5",X"01",X"20",X"00",
		X"09",X"EB",X"01",X"40",X"00",X"09",X"EB",X"C1",X"10",X"F0",X"E1",X"E5",X"D5",X"11",X"40",X"FE",
		X"19",X"11",X"20",X"00",X"06",X"0E",X"36",X"00",X"19",X"10",X"FB",X"D1",X"E1",X"C3",X"04",X"1A",
		X"0E",X"A7",X"FE",X"8D",X"CA",X"FF",X"1A",X"FE",X"91",X"CA",X"FF",X"1A",X"0D",X"FE",X"8E",X"CA",
		X"FF",X"1A",X"FE",X"90",X"CA",X"FF",X"1A",X"0E",X"A5",X"FE",X"8F",X"28",X"62",X"0E",X"A4",X"FE",
		X"70",X"28",X"5C",X"FE",X"76",X"28",X"58",X"FE",X"77",X"28",X"54",X"0D",X"FE",X"6E",X"28",X"4F",
		X"FE",X"6F",X"28",X"4B",X"FE",X"74",X"28",X"47",X"FE",X"75",X"28",X"43",X"0D",X"FE",X"8D",X"28",
		X"3E",X"FE",X"6D",X"28",X"3A",X"FE",X"73",X"28",X"36",X"FE",X"90",X"28",X"32",X"0D",X"FE",X"6C",
		X"28",X"2D",X"FE",X"68",X"28",X"29",X"FE",X"72",X"28",X"25",X"FE",X"6C",X"28",X"21",X"FE",X"69",
		X"28",X"1D",X"FE",X"6A",X"28",X"19",X"FE",X"6B",X"28",X"15",X"FE",X"71",X"28",X"11",X"FE",X"78",
		X"28",X"0D",X"FE",X"79",X"28",X"09",X"FE",X"8E",X"28",X"05",X"FE",X"91",X"28",X"01",X"0D",X"79",
		X"C9",X"E5",X"D5",X"C5",X"47",X"3A",X"7C",X"E2",X"80",X"4F",X"E6",X"01",X"32",X"7C",X"E2",X"79",
		X"CB",X"3F",X"4F",X"3A",X"81",X"E1",X"91",X"32",X"81",X"E1",X"3A",X"7D",X"E2",X"80",X"4F",X"E6",
		X"03",X"32",X"7D",X"E2",X"79",X"CB",X"3F",X"CB",X"3F",X"4F",X"3A",X"82",X"E1",X"91",X"32",X"82",
		X"E1",X"3A",X"7B",X"E2",X"2F",X"E6",X"07",X"80",X"47",X"E6",X"07",X"2F",X"E6",X"07",X"32",X"7B",
		X"E2",X"78",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"20",X"0F",X"3A",X"7A",X"E2",X"47",X"3A",X"7B",
		X"E2",X"80",X"32",X"80",X"E1",X"C1",X"D1",X"E1",X"C9",X"47",X"CB",X"20",X"CB",X"20",X"CB",X"20",
		X"3A",X"7A",X"E2",X"90",X"32",X"7A",X"E2",X"CD",X"01",X"0E",X"21",X"83",X"E3",X"34",X"20",X"02",
		X"23",X"34",X"3A",X"79",X"E2",X"3C",X"32",X"79",X"E2",X"FE",X"20",X"20",X"12",X"3A",X"78",X"E2",
		X"3C",X"3C",X"E6",X"7F",X"32",X"78",X"E2",X"3E",X"10",X"32",X"79",X"E2",X"CD",X"23",X"19",X"3A",
		X"7A",X"E2",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"6F",X"3E",X"1F",X"95",X"3D",X"E6",X"1F",X"6F",
		X"26",X"83",X"3A",X"79",X"E2",X"C6",X"1E",X"5F",X"16",X"EC",X"E5",X"06",X"08",X"1A",X"77",X"C5",
		X"01",X"20",X"00",X"09",X"EB",X"01",X"40",X"00",X"09",X"EB",X"C1",X"10",X"F0",X"E1",X"E5",X"D5",
		X"11",X"40",X"FE",X"19",X"EB",X"21",X"00",X"04",X"19",X"EB",X"7E",X"FE",X"1A",X"20",X"05",X"3E",
		X"00",X"32",X"2C",X"E3",X"06",X"0E",X"36",X"00",X"3E",X"00",X"12",X"C5",X"D5",X"01",X"20",X"00",
		X"09",X"EB",X"E1",X"09",X"EB",X"C1",X"10",X"EE",X"D1",X"E1",X"11",X"00",X"04",X"EB",X"19",X"06",
		X"08",X"1A",X"CD",X"80",X"1A",X"77",X"C5",X"01",X"20",X"00",X"09",X"E5",X"EB",X"09",X"EB",X"E1",
		X"C1",X"10",X"EE",X"C3",X"4A",X"1B",X"3D",X"3E",X"3D",X"3E",X"3D",X"3E",X"3D",X"3E",X"3D",X"3E",
		X"3D",X"3E",X"3D",X"3E",X"3D",X"3E",X"3D",X"3E",X"3D",X"3E",X"3D",X"3E",X"3D",X"3E",X"3D",X"3E",
		X"3D",X"3E",X"3D",X"3E",X"3D",X"3E",X"3F",X"40",X"3F",X"40",X"3F",X"40",X"3F",X"40",X"3F",X"40",
		X"3F",X"40",X"3F",X"40",X"3F",X"40",X"3F",X"40",X"3F",X"40",X"3F",X"40",X"3F",X"40",X"3F",X"40",
		X"3F",X"40",X"3F",X"40",X"3F",X"40",X"E5",X"D5",X"C5",X"3A",X"0E",X"E2",X"6F",X"26",X"20",X"7E",
		X"47",X"3A",X"0F",X"E2",X"80",X"32",X"0F",X"E2",X"2C",X"7D",X"32",X"0E",X"E2",X"3A",X"0F",X"E2",
		X"C1",X"D1",X"E1",X"C9",X"DD",X"E5",X"E5",X"D5",X"C5",X"6F",X"CB",X"25",X"CB",X"25",X"26",X"E0",
		X"C5",X"01",X"60",X"00",X"09",X"C1",X"E5",X"DD",X"E1",X"DD",X"71",X"00",X"DD",X"70",X"03",X"DD",
		X"72",X"01",X"DD",X"73",X"02",X"C5",X"01",X"60",X"00",X"DD",X"09",X"C1",X"DD",X"71",X"00",X"DD",
		X"70",X"03",X"DD",X"72",X"01",X"DD",X"73",X"02",X"C5",X"01",X"60",X"00",X"DD",X"09",X"C1",X"DD",
		X"71",X"00",X"DD",X"70",X"03",X"DD",X"72",X"01",X"DD",X"73",X"02",X"C1",X"D1",X"E1",X"DD",X"E1",
		X"C9",X"3E",X"10",X"32",X"10",X"E2",X"3E",X"60",X"32",X"11",X"E2",X"3E",X"01",X"32",X"12",X"E2",
		X"3E",X"00",X"32",X"14",X"E2",X"3E",X"01",X"32",X"15",X"E2",X"C3",X"CD",X"1C",X"3E",X"01",X"32",
		X"12",X"E2",X"3A",X"4E",X"E2",X"FE",X"00",X"28",X"0D",X"21",X"4F",X"E2",X"35",X"20",X"03",X"3E",
		X"04",X"77",X"7E",X"32",X"12",X"E2",X"3A",X"10",X"E2",X"47",X"3A",X"11",X"E2",X"4F",X"3A",X"12",
		X"E2",X"57",X"1E",X"01",X"3E",X"00",X"CD",X"64",X"1C",X"1E",X"02",X"3A",X"13",X"E2",X"FE",X"00",
		X"28",X"06",X"1E",X"03",X"FE",X"01",X"28",X"00",X"3A",X"12",X"E2",X"57",X"3A",X"10",X"E2",X"C6",
		X"10",X"47",X"3A",X"11",X"E2",X"4F",X"3E",X"01",X"CD",X"64",X"1C",X"3A",X"10",X"E2",X"D6",X"07",
		X"47",X"3A",X"11",X"E2",X"4F",X"16",X"01",X"3A",X"14",X"E2",X"FE",X"00",X"20",X"03",X"3A",X"1F",
		X"E2",X"5F",X"3E",X"02",X"CD",X"64",X"1C",X"3A",X"43",X"E2",X"FE",X"01",X"CA",X"C1",X"1D",X"3A",
		X"16",X"E2",X"FE",X"00",X"28",X"16",X"3A",X"1B",X"E2",X"47",X"3A",X"1C",X"E2",X"4F",X"3A",X"1A",
		X"E2",X"5F",X"16",X"01",X"3E",X"03",X"CD",X"64",X"1C",X"C3",X"80",X"1D",X"3A",X"10",X"E2",X"C6",
		X"20",X"47",X"3A",X"11",X"E2",X"4F",X"3A",X"18",X"E2",X"C6",X"0A",X"5F",X"16",X"01",X"3A",X"17",
		X"E2",X"FE",X"00",X"20",X"06",X"01",X"00",X"00",X"11",X"00",X"00",X"3E",X"03",X"CD",X"64",X"1C",
		X"3A",X"26",X"E2",X"FE",X"00",X"28",X"16",X"3A",X"2B",X"E2",X"47",X"3A",X"2C",X"E2",X"4F",X"3A",
		X"2A",X"E2",X"5F",X"16",X"01",X"3E",X"04",X"CD",X"64",X"1C",X"C3",X"C1",X"1D",X"3A",X"10",X"E2",
		X"C6",X"20",X"47",X"3A",X"11",X"E2",X"4F",X"3A",X"28",X"E2",X"C6",X"0A",X"5F",X"16",X"01",X"3A",
		X"27",X"E2",X"FE",X"00",X"20",X"06",X"01",X"00",X"00",X"11",X"00",X"00",X"3E",X"04",X"CD",X"64",
		X"1C",X"3A",X"42",X"E2",X"FE",X"00",X"CA",X"DC",X"1D",X"3A",X"01",X"E3",X"47",X"3A",X"02",X"E3",
		X"4F",X"16",X"01",X"3A",X"03",X"E3",X"5F",X"3E",X"07",X"CD",X"64",X"1C",X"C9",X"3A",X"0B",X"E2",
		X"FE",X"00",X"28",X"10",X"3A",X"11",X"E2",X"3D",X"3D",X"E6",X"FE",X"FE",X"10",X"20",X"02",X"3E",
		X"12",X"32",X"11",X"E2",X"3A",X"0A",X"E2",X"FE",X"00",X"28",X"10",X"3A",X"11",X"E2",X"3C",X"3C",
		X"E6",X"FE",X"FE",X"B0",X"20",X"02",X"3E",X"AE",X"32",X"11",X"E2",X"C3",X"CD",X"1C",X"3A",X"0C",
		X"E2",X"FE",X"00",X"28",X"18",X"3E",X"00",X"32",X"14",X"E2",X"3A",X"10",X"E2",X"3D",X"3D",X"E6",
		X"FE",X"FE",X"20",X"20",X"02",X"3E",X"22",X"32",X"10",X"E2",X"C3",X"CD",X"1C",X"3A",X"0D",X"E2",
		X"FE",X"00",X"20",X"04",X"32",X"14",X"E2",X"C9",X"3A",X"14",X"E2",X"FE",X"00",X"20",X"05",X"3E",
		X"06",X"32",X"14",X"E2",X"3A",X"10",X"E2",X"3C",X"3C",X"E6",X"FE",X"FE",X"B2",X"20",X"02",X"3E",
		X"B0",X"32",X"10",X"E2",X"C3",X"CD",X"1C",X"3A",X"10",X"E2",X"C6",X"18",X"47",X"3A",X"11",X"E2",
		X"4F",X"CD",X"7C",X"3A",X"11",X"C1",X"FF",X"19",X"7E",X"E6",X"FC",X"FE",X"14",X"CA",X"9E",X"1E",
		X"23",X"7E",X"E6",X"FC",X"FE",X"14",X"CA",X"9E",X"1E",X"23",X"7E",X"E6",X"FC",X"FE",X"14",X"28",
		X"1D",X"11",X"1E",X"00",X"19",X"7E",X"E6",X"FC",X"FE",X"14",X"CA",X"9E",X"1E",X"23",X"7E",X"E6",
		X"FC",X"FE",X"14",X"28",X"09",X"23",X"7E",X"E6",X"FC",X"FE",X"14",X"C2",X"0A",X"1F",X"11",X"00",
		X"04",X"19",X"7E",X"CB",X"27",X"DA",X"0A",X"1F",X"11",X"00",X"FC",X"19",X"7E",X"E6",X"03",X"CB",
		X"27",X"5F",X"16",X"00",X"E5",X"21",X"15",X"21",X"19",X"56",X"23",X"5E",X"E1",X"19",X"E5",X"FD",
		X"E1",X"DD",X"21",X"90",X"E3",X"DD",X"7E",X"02",X"FD",X"77",X"00",X"DD",X"7E",X"03",X"FD",X"77",
		X"01",X"DD",X"7E",X"04",X"FD",X"77",X"20",X"DD",X"7E",X"05",X"FD",X"77",X"21",X"11",X"00",X"04",
		X"FD",X"19",X"DD",X"7E",X"06",X"FD",X"77",X"00",X"DD",X"7E",X"07",X"FD",X"77",X"01",X"DD",X"7E",
		X"08",X"FD",X"77",X"20",X"DD",X"7E",X"09",X"FD",X"77",X"21",X"CD",X"A5",X"3C",X"3E",X"96",X"CD",
		X"A0",X"33",X"3E",X"04",X"CD",X"75",X"22",X"C3",X"0D",X"1F",X"CD",X"1D",X"21",X"3A",X"1A",X"E2",
		X"EE",X"01",X"32",X"1A",X"E2",X"3A",X"2A",X"E2",X"EE",X"01",X"32",X"2A",X"E2",X"21",X"15",X"E2",
		X"35",X"20",X"23",X"3E",X"04",X"77",X"3A",X"1F",X"E2",X"06",X"08",X"FE",X"08",X"20",X"02",X"06",
		X"09",X"78",X"32",X"1F",X"E2",X"3A",X"14",X"E2",X"FE",X"00",X"28",X"0A",X"3C",X"FE",X"08",X"20",
		X"02",X"3E",X"06",X"32",X"14",X"E2",X"3E",X"01",X"32",X"12",X"E2",X"CD",X"CD",X"1C",X"C9",X"3A",
		X"17",X"E2",X"FE",X"00",X"28",X"05",X"32",X"05",X"E2",X"18",X"06",X"3A",X"27",X"E2",X"32",X"05",
		X"E2",X"CD",X"5C",X"37",X"3A",X"43",X"E2",X"FE",X"00",X"C0",X"3A",X"16",X"E2",X"FE",X"00",X"C2",
		X"E9",X"1F",X"3A",X"26",X"E2",X"FE",X"00",X"20",X"08",X"3A",X"27",X"E2",X"FE",X"00",X"C2",X"E9",
		X"1F",X"3A",X"08",X"E2",X"FE",X"00",X"20",X"41",X"3A",X"17",X"E2",X"FE",X"00",X"CA",X"E9",X"1F",
		X"3E",X"01",X"CD",X"75",X"22",X"3A",X"17",X"E2",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",
		X"CB",X"3F",X"CB",X"3F",X"CB",X"27",X"C6",X"0E",X"32",X"1A",X"E2",X"3E",X"06",X"32",X"1D",X"E2",
		X"3E",X"00",X"32",X"18",X"E2",X"3E",X"01",X"32",X"16",X"E2",X"3A",X"10",X"E2",X"C6",X"10",X"32",
		X"1B",X"E2",X"3A",X"11",X"E2",X"32",X"1C",X"E2",X"C9",X"3A",X"17",X"E2",X"C6",X"08",X"D2",X"D3",
		X"1F",X"3E",X"FF",X"32",X"17",X"E2",X"21",X"1E",X"E2",X"35",X"20",X"0C",X"3E",X"04",X"77",X"3A",
		X"18",X"E2",X"3C",X"E6",X"03",X"32",X"18",X"E2",X"C9",X"3A",X"26",X"E2",X"FE",X"00",X"C0",X"3A",
		X"08",X"E2",X"FE",X"00",X"20",X"3F",X"3A",X"27",X"E2",X"FE",X"00",X"C8",X"3E",X"01",X"CD",X"75",
		X"22",X"3A",X"27",X"E2",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",
		X"CB",X"27",X"C6",X"0E",X"32",X"2A",X"E2",X"3E",X"06",X"32",X"2D",X"E2",X"3E",X"00",X"32",X"28",
		X"E2",X"3E",X"01",X"32",X"26",X"E2",X"3A",X"10",X"E2",X"C6",X"10",X"32",X"2B",X"E2",X"3A",X"11",
		X"E2",X"32",X"2C",X"E2",X"C9",X"3A",X"27",X"E2",X"C6",X"08",X"D2",X"3F",X"20",X"3E",X"FF",X"32",
		X"27",X"E2",X"21",X"2E",X"E2",X"35",X"20",X"0C",X"3E",X"04",X"77",X"3A",X"28",X"E2",X"3C",X"E6",
		X"03",X"32",X"28",X"E2",X"C9",X"CD",X"7F",X"20",X"3A",X"16",X"E2",X"FE",X"00",X"C8",X"3A",X"1B",
		X"E2",X"47",X"3A",X"1D",X"E2",X"80",X"32",X"1B",X"E2",X"FE",X"F8",X"DA",X"7C",X"20",X"3E",X"00",
		X"32",X"16",X"E2",X"32",X"17",X"E2",X"32",X"18",X"E2",X"C3",X"CD",X"1C",X"C3",X"CD",X"1C",X"3A",
		X"26",X"E2",X"FE",X"00",X"C8",X"3A",X"2B",X"E2",X"47",X"3A",X"2D",X"E2",X"80",X"32",X"2B",X"E2",
		X"FE",X"F8",X"DA",X"A0",X"20",X"3E",X"00",X"32",X"26",X"E2",X"32",X"27",X"E2",X"32",X"28",X"E2",
		X"C9",X"3A",X"16",X"E2",X"FE",X"00",X"20",X"03",X"3E",X"FF",X"C9",X"3A",X"6E",X"E0",X"D6",X"0E",
		X"CB",X"3F",X"6F",X"26",X"00",X"11",X"D3",X"20",X"CB",X"25",X"CB",X"25",X"19",X"46",X"23",X"4E",
		X"23",X"56",X"23",X"5E",X"3A",X"6C",X"E0",X"67",X"78",X"84",X"47",X"3A",X"6F",X"E0",X"6F",X"79",
		X"85",X"4F",X"C9",X"F8",X"F4",X"18",X"20",X"F8",X"F4",X"18",X"20",X"F4",X"F4",X"20",X"20",X"F0",
		X"F4",X"28",X"28",X"3A",X"26",X"E2",X"FE",X"00",X"20",X"03",X"3E",X"FF",X"C9",X"3A",X"72",X"E0",
		X"D6",X"0E",X"CB",X"3F",X"6F",X"26",X"00",X"11",X"D3",X"20",X"CB",X"25",X"CB",X"25",X"19",X"46",
		X"23",X"4E",X"23",X"56",X"23",X"5E",X"3A",X"70",X"E0",X"67",X"78",X"84",X"47",X"3A",X"73",X"E0",
		X"6F",X"79",X"85",X"4F",X"C9",X"00",X"00",X"FF",X"FF",X"FF",X"E0",X"FF",X"DF",X"3A",X"10",X"E2",
		X"C6",X"18",X"47",X"3A",X"11",X"E2",X"4F",X"CD",X"7C",X"3A",X"7E",X"FE",X"18",X"28",X"08",X"11",
		X"20",X"00",X"19",X"7E",X"FE",X"18",X"C0",X"3E",X"09",X"CD",X"75",X"22",X"E5",X"11",X"00",X"04",
		X"19",X"7E",X"E1",X"CB",X"27",X"D8",X"3E",X"00",X"77",X"11",X"00",X"04",X"19",X"77",X"21",X"06",
		X"E2",X"7E",X"C6",X"0C",X"77",X"C6",X"40",X"30",X"16",X"3A",X"03",X"E2",X"3C",X"E6",X"0F",X"32",
		X"03",X"E2",X"3E",X"10",X"77",X"F5",X"CD",X"C6",X"37",X"3E",X"06",X"CD",X"75",X"22",X"F1",X"C6",
		X"40",X"38",X"E6",X"C9",X"21",X"10",X"E2",X"46",X"23",X"4E",X"CD",X"7C",X"3A",X"23",X"23",X"11",
		X"E0",X"FF",X"19",X"7E",X"FE",X"1A",X"28",X"10",X"11",X"20",X"00",X"19",X"7E",X"FE",X"1A",X"28",
		X"07",X"19",X"7E",X"FE",X"1A",X"28",X"01",X"C9",X"11",X"00",X"04",X"E5",X"19",X"7E",X"E1",X"CB",
		X"27",X"D8",X"3E",X"00",X"77",X"3E",X"01",X"32",X"13",X"E2",X"3A",X"2C",X"E3",X"3C",X"E6",X"0F",
		X"32",X"2C",X"E3",X"FE",X"0A",X"20",X"05",X"3E",X"09",X"32",X"2C",X"E3",X"3E",X"64",X"CD",X"A0",
		X"33",X"21",X"1E",X"E3",X"34",X"3E",X"02",X"CD",X"75",X"22",X"C9",X"3A",X"13",X"E2",X"FE",X"00",
		X"C8",X"21",X"10",X"E2",X"46",X"23",X"4E",X"CD",X"7C",X"3A",X"7E",X"FE",X"6C",X"28",X"0B",X"FE",
		X"72",X"28",X"07",X"FE",X"68",X"28",X"03",X"FE",X"69",X"C0",X"3E",X"00",X"32",X"13",X"E2",X"21",
		X"00",X"83",X"06",X"1F",X"7E",X"FE",X"03",X"28",X"06",X"23",X"10",X"F8",X"C3",X"13",X"22",X"3E",
		X"2B",X"23",X"77",X"2B",X"3A",X"2C",X"E3",X"C6",X"21",X"77",X"3E",X"28",X"11",X"00",X"04",X"19",
		X"77",X"23",X"77",X"3A",X"2C",X"E3",X"6F",X"26",X"00",X"11",X"65",X"22",X"19",X"06",X"0A",X"7E",
		X"CD",X"A0",X"33",X"10",X"FA",X"3A",X"2C",X"E3",X"FE",X"09",X"20",X"29",X"21",X"1A",X"36",X"11",
		X"B3",X"84",X"01",X"0A",X"00",X"ED",X"B0",X"01",X"08",X"00",X"3A",X"2D",X"E3",X"FE",X"03",X"28",
		X"01",X"3C",X"32",X"2D",X"E3",X"47",X"CB",X"27",X"80",X"6F",X"26",X"00",X"11",X"B3",X"84",X"19",
		X"3E",X"12",X"77",X"23",X"77",X"3E",X"00",X"32",X"2C",X"E3",X"21",X"1E",X"E3",X"34",X"3E",X"03",
		X"CD",X"75",X"22",X"C9",X"C9",X"05",X"0A",X"0F",X"14",X"19",X"1E",X"23",X"28",X"2D",X"32",X"32",
		X"32",X"32",X"32",X"32",X"32",X"F5",X"3A",X"01",X"E2",X"FE",X"00",X"28",X"02",X"F1",X"C9",X"F1",
		X"32",X"00",X"D0",X"F6",X"80",X"32",X"00",X"D0",X"C9",X"3A",X"87",X"E3",X"FE",X"00",X"C0",X"21",
		X"50",X"E2",X"35",X"C0",X"3A",X"40",X"E2",X"77",X"21",X"51",X"E2",X"34",X"7E",X"E6",X"07",X"77",
		X"5F",X"16",X"00",X"CB",X"23",X"CB",X"23",X"CB",X"23",X"CB",X"23",X"CB",X"12",X"3A",X"2E",X"E3",
		X"47",X"0E",X"00",X"CB",X"38",X"CB",X"19",X"21",X"E2",X"22",X"19",X"09",X"06",X"03",X"56",X"23",
		X"5E",X"23",X"D5",X"DD",X"E1",X"DD",X"7E",X"00",X"FE",X"00",X"C0",X"7E",X"DD",X"77",X"01",X"23",
		X"7E",X"DD",X"77",X"03",X"3E",X"01",X"DD",X"77",X"00",X"3E",X"00",X"DD",X"77",X"02",X"23",X"10",
		X"DD",X"C9",X"E2",X"30",X"00",X"18",X"E2",X"34",X"00",X"18",X"E2",X"38",X"00",X"18",X"00",X"00",
		X"00",X"00",X"E2",X"30",X"00",X"18",X"E2",X"34",X"00",X"18",X"E2",X"38",X"00",X"18",X"00",X"00",
		X"00",X"00",X"E2",X"30",X"00",X"18",X"E2",X"34",X"00",X"18",X"E2",X"38",X"00",X"18",X"00",X"00",
		X"00",X"00",X"E2",X"30",X"01",X"18",X"E2",X"34",X"01",X"18",X"E2",X"38",X"01",X"18",X"00",X"00",
		X"00",X"00",X"E2",X"30",X"01",X"18",X"E2",X"34",X"03",X"18",X"E2",X"38",X"02",X"18",X"00",X"00",
		X"00",X"00",X"E2",X"30",X"03",X"18",X"E2",X"34",X"03",X"18",X"E2",X"38",X"01",X"18",X"00",X"00",
		X"00",X"00",X"E2",X"30",X"00",X"18",X"E2",X"34",X"00",X"18",X"E2",X"38",X"00",X"18",X"00",X"00",
		X"00",X"00",X"E2",X"30",X"00",X"18",X"E2",X"34",X"00",X"18",X"E2",X"38",X"00",X"18",X"00",X"00",
		X"00",X"00",X"E2",X"30",X"00",X"20",X"E2",X"34",X"00",X"20",X"E2",X"38",X"00",X"20",X"00",X"00",
		X"00",X"00",X"E2",X"30",X"00",X"20",X"E2",X"34",X"00",X"18",X"E2",X"38",X"00",X"20",X"00",X"00",
		X"00",X"00",X"E2",X"30",X"00",X"18",X"E2",X"34",X"00",X"18",X"E2",X"38",X"00",X"18",X"00",X"00",
		X"00",X"00",X"E2",X"30",X"01",X"20",X"E2",X"34",X"01",X"18",X"E2",X"38",X"01",X"20",X"00",X"00",
		X"00",X"00",X"E2",X"30",X"01",X"18",X"E2",X"34",X"03",X"18",X"E2",X"38",X"02",X"18",X"00",X"00",
		X"00",X"00",X"E2",X"30",X"03",X"20",X"E2",X"34",X"03",X"20",X"E2",X"38",X"01",X"20",X"00",X"00",
		X"00",X"00",X"E2",X"30",X"00",X"18",X"E2",X"34",X"00",X"18",X"E2",X"38",X"00",X"20",X"00",X"00",
		X"00",X"00",X"E2",X"30",X"00",X"18",X"E2",X"34",X"00",X"18",X"E2",X"38",X"00",X"18",X"00",X"00",
		X"00",X"00",X"E2",X"30",X"00",X"24",X"E2",X"34",X"00",X"18",X"E2",X"38",X"00",X"24",X"00",X"00",
		X"00",X"00",X"E2",X"30",X"00",X"24",X"E2",X"34",X"00",X"24",X"E2",X"38",X"00",X"24",X"00",X"00",
		X"00",X"00",X"E2",X"30",X"00",X"18",X"E2",X"34",X"00",X"20",X"E2",X"38",X"00",X"24",X"00",X"00",
		X"00",X"00",X"E2",X"30",X"01",X"24",X"E2",X"34",X"01",X"18",X"E2",X"38",X"01",X"24",X"00",X"00",
		X"00",X"00",X"E2",X"30",X"01",X"18",X"E2",X"34",X"03",X"1C",X"E2",X"38",X"02",X"24",X"00",X"00",
		X"00",X"00",X"E2",X"30",X"03",X"24",X"E2",X"34",X"03",X"24",X"E2",X"38",X"01",X"24",X"00",X"00",
		X"00",X"00",X"E2",X"30",X"00",X"18",X"E2",X"34",X"00",X"24",X"E2",X"38",X"00",X"24",X"00",X"00",
		X"00",X"00",X"E2",X"30",X"00",X"24",X"E2",X"34",X"00",X"18",X"E2",X"38",X"00",X"24",X"00",X"00",
		X"00",X"00",X"E2",X"30",X"00",X"1C",X"E2",X"34",X"00",X"1C",X"E2",X"38",X"00",X"1C",X"00",X"00",
		X"00",X"00",X"E2",X"30",X"00",X"1C",X"E2",X"34",X"00",X"1C",X"E2",X"38",X"00",X"1C",X"00",X"00",
		X"00",X"00",X"E2",X"30",X"00",X"24",X"E2",X"34",X"00",X"24",X"E2",X"38",X"00",X"24",X"00",X"00",
		X"00",X"00",X"E2",X"30",X"01",X"24",X"E2",X"34",X"01",X"18",X"E2",X"38",X"01",X"1C",X"00",X"00",
		X"00",X"00",X"E2",X"30",X"01",X"1C",X"E2",X"34",X"03",X"1C",X"E2",X"38",X"02",X"1C",X"00",X"00",
		X"00",X"00",X"E2",X"30",X"03",X"24",X"E2",X"34",X"03",X"24",X"E2",X"38",X"01",X"24",X"00",X"00",
		X"00",X"00",X"E2",X"30",X"00",X"18",X"E2",X"34",X"00",X"18",X"E2",X"38",X"00",X"18",X"00",X"00",
		X"00",X"00",X"E2",X"30",X"00",X"18",X"E2",X"34",X"00",X"18",X"E2",X"38",X"00",X"18",X"00",X"00",
		X"00",X"00",X"E2",X"30",X"00",X"18",X"E2",X"34",X"00",X"18",X"E2",X"38",X"00",X"18",X"00",X"00",
		X"00",X"00",X"E2",X"30",X"00",X"1C",X"E2",X"34",X"00",X"1C",X"E2",X"38",X"00",X"1C",X"00",X"00",
		X"00",X"00",X"E2",X"30",X"00",X"24",X"E2",X"34",X"00",X"24",X"E2",X"38",X"00",X"24",X"00",X"00",
		X"00",X"00",X"E2",X"30",X"01",X"24",X"E2",X"34",X"01",X"18",X"E2",X"38",X"01",X"1C",X"00",X"00",
		X"00",X"00",X"E2",X"30",X"01",X"18",X"E2",X"34",X"03",X"18",X"E2",X"38",X"02",X"18",X"00",X"00",
		X"00",X"00",X"E2",X"30",X"03",X"24",X"E2",X"34",X"03",X"24",X"E2",X"38",X"01",X"24",X"00",X"00",
		X"00",X"00",X"E2",X"30",X"00",X"18",X"E2",X"34",X"00",X"18",X"E2",X"38",X"00",X"18",X"00",X"00",
		X"00",X"00",X"E2",X"30",X"00",X"18",X"E2",X"34",X"00",X"18",X"E2",X"38",X"00",X"18",X"00",X"00",
		X"00",X"00",X"21",X"3C",X"E2",X"35",X"C0",X"CD",X"46",X"1C",X"E6",X"1F",X"C6",X"10",X"77",X"DD",
		X"21",X"30",X"E2",X"FD",X"21",X"E4",X"E0",X"0E",X"00",X"06",X"90",X"CD",X"9D",X"25",X"DD",X"21",
		X"34",X"E2",X"FD",X"21",X"84",X"E0",X"06",X"50",X"0E",X"04",X"CD",X"9D",X"25",X"DD",X"21",X"38",
		X"E2",X"FD",X"21",X"44",X"E1",X"06",X"10",X"0E",X"04",X"C3",X"9D",X"25",X"C9",X"DD",X"7E",X"00",
		X"FE",X"01",X"C0",X"DD",X"7E",X"02",X"FE",X"04",X"C8",X"DD",X"7E",X"01",X"FE",X"03",X"CA",X"BB",
		X"25",X"FE",X"02",X"CA",X"BB",X"25",X"FE",X"01",X"CA",X"54",X"26",X"C5",X"DD",X"5E",X"02",X"16",
		X"00",X"CB",X"23",X"CB",X"23",X"FD",X"19",X"78",X"C6",X"10",X"47",X"CD",X"46",X"1C",X"E6",X"1F",
		X"4F",X"78",X"91",X"47",X"FD",X"70",X"00",X"3E",X"F6",X"FD",X"77",X"03",X"DD",X"7E",X"03",X"FD",
		X"77",X"02",X"3E",X"04",X"FD",X"77",X"01",X"51",X"CB",X"3A",X"CB",X"3A",X"CB",X"3A",X"E5",X"5A",
		X"16",X"00",X"21",X"0F",X"26",X"19",X"7E",X"E1",X"C1",X"06",X"00",X"21",X"F0",X"E3",X"09",X"77",
		X"DD",X"34",X"02",X"DD",X"7E",X"02",X"FE",X"04",X"C0",X"3E",X"02",X"DD",X"77",X"00",X"C9",X"10",
		X"18",X"08",X"00",X"DD",X"5E",X"02",X"16",X"00",X"CB",X"23",X"CB",X"23",X"FD",X"19",X"78",X"D6",
		X"0A",X"FD",X"77",X"00",X"3E",X"F6",X"FD",X"77",X"03",X"FD",X"77",X"07",X"DD",X"7E",X"03",X"FD",
		X"77",X"02",X"FD",X"77",X"06",X"3E",X"04",X"FD",X"77",X"01",X"FD",X"77",X"05",X"78",X"C6",X"0A",
		X"FD",X"77",X"04",X"DD",X"7E",X"02",X"3C",X"3C",X"DD",X"77",X"02",X"FE",X"04",X"C0",X"3E",X"02",
		X"DD",X"77",X"00",X"C9",X"DD",X"5E",X"02",X"16",X"00",X"CB",X"23",X"CB",X"23",X"FD",X"19",X"DD",
		X"7E",X"02",X"FE",X"01",X"20",X"2E",X"78",X"D6",X"0A",X"FD",X"77",X"00",X"78",X"C6",X"0A",X"FD",
		X"77",X"04",X"3E",X"F6",X"FD",X"77",X"03",X"FD",X"77",X"07",X"3E",X"04",X"FD",X"77",X"01",X"FD",
		X"77",X"05",X"DD",X"7E",X"03",X"FD",X"77",X"02",X"FD",X"77",X"06",X"DD",X"7E",X"02",X"C6",X"02",
		X"DD",X"77",X"02",X"C9",X"FD",X"70",X"00",X"DD",X"7E",X"03",X"FD",X"77",X"02",X"3E",X"04",X"FD",
		X"77",X"01",X"3E",X"F6",X"FD",X"77",X"03",X"DD",X"7E",X"02",X"3C",X"DD",X"77",X"02",X"FE",X"04",
		X"C0",X"3E",X"02",X"DD",X"77",X"00",X"C9",X"78",X"D6",X"20",X"FD",X"77",X"00",X"C6",X"10",X"FD",
		X"77",X"04",X"C6",X"10",X"FD",X"77",X"08",X"C6",X"10",X"FD",X"77",X"0C",X"DD",X"7E",X"03",X"FD",
		X"77",X"02",X"FD",X"77",X"06",X"FD",X"77",X"0A",X"FD",X"77",X"0E",X"3E",X"F6",X"FD",X"77",X"03",
		X"FD",X"77",X"07",X"FD",X"77",X"0B",X"FD",X"77",X"0F",X"3E",X"04",X"FD",X"77",X"01",X"FD",X"77",
		X"05",X"FD",X"77",X"09",X"FD",X"77",X"0D",X"3E",X"04",X"DD",X"77",X"02",X"3E",X"02",X"DD",X"77",
		X"00",X"C9",X"21",X"57",X"E2",X"35",X"C0",X"3A",X"01",X"E6",X"77",X"21",X"3E",X"E2",X"35",X"20",
		X"0A",X"3E",X"02",X"77",X"3E",X"00",X"32",X"3F",X"E2",X"18",X"05",X"3E",X"01",X"32",X"3F",X"E2",
		X"21",X"FD",X"E3",X"35",X"20",X"09",X"3E",X"03",X"77",X"3E",X"00",X"2B",X"77",X"18",X"04",X"3E",
		X"01",X"2B",X"77",X"DD",X"21",X"30",X"E2",X"FD",X"21",X"E4",X"E0",X"CD",X"51",X"27",X"DD",X"21",
		X"34",X"E2",X"FD",X"21",X"84",X"E0",X"CD",X"51",X"27",X"DD",X"21",X"38",X"E2",X"FD",X"21",X"44",
		X"E1",X"DD",X"7E",X"00",X"FE",X"00",X"C8",X"DD",X"46",X"02",X"78",X"FE",X"00",X"C8",X"06",X"00",
		X"FD",X"E5",X"3A",X"FC",X"E3",X"FE",X"00",X"20",X"35",X"DD",X"7E",X"01",X"FE",X"01",X"28",X"2E",
		X"FD",X"7E",X"02",X"E6",X"FC",X"FE",X"28",X"28",X"25",X"FD",X"7E",X"00",X"FE",X"00",X"28",X"1E",
		X"DD",X"E5",X"E1",X"7D",X"D6",X"30",X"80",X"C6",X"F0",X"6F",X"26",X"E3",X"34",X"7E",X"E6",X"1F",
		X"6F",X"26",X"00",X"11",X"E3",X"30",X"19",X"7E",X"FD",X"86",X"00",X"FD",X"77",X"00",X"3A",X"3F",
		X"E2",X"FE",X"00",X"20",X"27",X"FD",X"7E",X"02",X"FE",X"2B",X"20",X"10",X"3E",X"00",X"FD",X"77",
		X"00",X"FD",X"77",X"01",X"FD",X"77",X"02",X"FD",X"77",X"03",X"18",X"10",X"FD",X"7E",X"02",X"E6",
		X"FC",X"4F",X"FD",X"7E",X"02",X"3C",X"E6",X"03",X"81",X"FD",X"77",X"02",X"FD",X"7E",X"02",X"E6",
		X"F8",X"FE",X"28",X"20",X"12",X"FD",X"34",X"03",X"FD",X"34",X"03",X"FD",X"34",X"03",X"FD",X"7E",
		X"03",X"E6",X"F8",X"28",X"10",X"18",X"1E",X"FD",X"7E",X"03",X"D6",X"02",X"E6",X"FE",X"FD",X"77",
		X"03",X"FE",X"F8",X"20",X"10",X"3E",X"00",X"FD",X"77",X"01",X"FD",X"77",X"02",X"FD",X"77",X"00",
		X"3E",X"FA",X"FD",X"77",X"03",X"FD",X"23",X"FD",X"23",X"FD",X"23",X"FD",X"23",X"04",X"78",X"DD",
		X"BE",X"02",X"C2",X"62",X"27",X"FD",X"E1",X"DD",X"7E",X"00",X"FE",X"02",X"C0",X"FD",X"7E",X"00",
		X"FE",X"00",X"C0",X"FD",X"7E",X"04",X"FE",X"00",X"C0",X"FD",X"7E",X"08",X"FE",X"00",X"C0",X"FD",
		X"7E",X"0C",X"FE",X"00",X"C0",X"3E",X"00",X"DD",X"77",X"00",X"C9",X"CD",X"A1",X"20",X"FE",X"FF",
		X"28",X"1A",X"78",X"32",X"52",X"E2",X"79",X"32",X"53",X"E2",X"78",X"82",X"32",X"54",X"E2",X"79",
		X"83",X"32",X"55",X"E2",X"3E",X"01",X"32",X"56",X"E2",X"CD",X"CB",X"2A",X"CD",X"E3",X"20",X"FE",
		X"FF",X"28",X"1A",X"78",X"32",X"52",X"E2",X"79",X"32",X"53",X"E2",X"78",X"82",X"32",X"54",X"E2",
		X"79",X"83",X"32",X"55",X"E2",X"3E",X"02",X"32",X"56",X"E2",X"CD",X"CB",X"2A",X"3A",X"44",X"E2",
		X"D6",X"10",X"32",X"53",X"E2",X"C6",X"20",X"32",X"55",X"E2",X"3A",X"45",X"E2",X"D6",X"18",X"32",
		X"52",X"E2",X"C6",X"20",X"32",X"54",X"E2",X"3E",X"03",X"32",X"56",X"E2",X"3A",X"46",X"E2",X"FE",
		X"01",X"CC",X"CB",X"2A",X"3A",X"48",X"E2",X"D6",X"10",X"32",X"53",X"E2",X"C6",X"20",X"32",X"55",
		X"E2",X"3A",X"49",X"E2",X"D6",X"18",X"32",X"52",X"E2",X"C6",X"20",X"32",X"54",X"E2",X"3E",X"04",
		X"32",X"56",X"E2",X"3A",X"4A",X"E2",X"FE",X"01",X"CC",X"CB",X"2A",X"3A",X"07",X"E3",X"FE",X"00",
		X"28",X"22",X"3A",X"08",X"E3",X"D6",X"08",X"32",X"53",X"E2",X"C6",X"10",X"32",X"55",X"E2",X"3A",
		X"09",X"E3",X"D6",X"08",X"32",X"52",X"E2",X"C6",X"10",X"32",X"54",X"E2",X"3E",X"05",X"32",X"56",
		X"E2",X"CD",X"CB",X"2A",X"3A",X"10",X"E3",X"FE",X"00",X"28",X"25",X"3A",X"11",X"E3",X"D6",X"08",
		X"32",X"53",X"E2",X"C6",X"10",X"32",X"55",X"E2",X"3A",X"12",X"E3",X"C6",X"08",X"32",X"54",X"E2",
		X"3A",X"16",X"E3",X"D6",X"10",X"32",X"52",X"E2",X"3E",X"06",X"32",X"56",X"E2",X"CD",X"CB",X"2A",
		X"C9",X"16",X"FF",X"3A",X"52",X"E2",X"B8",X"D0",X"3A",X"54",X"E2",X"B8",X"D8",X"3A",X"53",X"E2",
		X"B9",X"D0",X"3A",X"55",X"E2",X"B9",X"D8",X"16",X"00",X"C9",X"DD",X"21",X"80",X"E2",X"DD",X"7E",
		X"00",X"FE",X"00",X"28",X"18",X"DD",X"7E",X"03",X"E6",X"FC",X"FE",X"30",X"28",X"0F",X"DD",X"46",
		X"01",X"DD",X"4E",X"04",X"CD",X"21",X"29",X"7A",X"FE",X"00",X"CC",X"30",X"2B",X"11",X"08",X"00",
		X"DD",X"19",X"DD",X"E5",X"D1",X"7B",X"FE",X"D0",X"20",X"D4",X"C9",X"DD",X"21",X"A0",X"E3",X"DD",
		X"7E",X"00",X"FE",X"00",X"20",X"0E",X"11",X"10",X"00",X"DD",X"19",X"DD",X"E5",X"D1",X"7B",X"FE",
		X"E0",X"20",X"EC",X"C9",X"FE",X"04",X"28",X"EE",X"FE",X"05",X"28",X"EA",X"FE",X"01",X"CA",X"06",
		X"2A",X"DD",X"46",X"02",X"DD",X"4E",X"01",X"CD",X"21",X"29",X"7A",X"FE",X"00",X"20",X"D7",X"3A",
		X"56",X"E2",X"FE",X"03",X"CA",X"03",X"31",X"FE",X"04",X"CA",X"4D",X"31",X"CD",X"7A",X"2A",X"7A",
		X"FE",X"00",X"C2",X"76",X"29",X"DD",X"7E",X"03",X"06",X"4B",X"FE",X"09",X"20",X"02",X"06",X"64",
		X"78",X"CD",X"A0",X"33",X"3E",X"07",X"CD",X"75",X"22",X"3E",X"02",X"DD",X"77",X"0B",X"3E",X"04",
		X"DD",X"77",X"00",X"3E",X"30",X"DD",X"77",X"04",X"DD",X"77",X"08",X"3E",X"03",X"DD",X"77",X"03",
		X"DD",X"77",X"07",X"3E",X"04",X"DD",X"77",X"00",X"C3",X"76",X"29",X"3E",X"04",X"DD",X"77",X"00",
		X"3E",X"30",X"DD",X"77",X"04",X"DD",X"77",X"08",X"3E",X"03",X"DD",X"77",X"03",X"DD",X"77",X"07",
		X"3E",X"04",X"DD",X"77",X"00",X"C9",X"DD",X"46",X"02",X"DD",X"4E",X"01",X"CD",X"21",X"29",X"7A",
		X"FE",X"00",X"C2",X"76",X"29",X"3A",X"56",X"E2",X"FE",X"04",X"CA",X"97",X"31",X"CD",X"7A",X"2A",
		X"7A",X"FE",X"00",X"C2",X"76",X"29",X"3E",X"96",X"CD",X"A0",X"33",X"3A",X"8A",X"E3",X"FE",X"01",
		X"CA",X"B5",X"29",X"3E",X"00",X"DD",X"77",X"09",X"DD",X"77",X"0F",X"3E",X"7D",X"DD",X"77",X"04",
		X"3E",X"7E",X"DD",X"77",X"08",X"3E",X"05",X"DD",X"77",X"00",X"DD",X"7E",X"01",X"32",X"E0",X"E3",
		X"C6",X"10",X"32",X"E4",X"E3",X"DD",X"7E",X"02",X"D6",X"08",X"32",X"E1",X"E3",X"32",X"E5",X"E3",
		X"3E",X"03",X"32",X"E2",X"E3",X"32",X"E6",X"E3",X"3E",X"68",X"32",X"E3",X"E3",X"3E",X"69",X"32",
		X"E7",X"E3",X"3E",X"01",X"32",X"8A",X"E3",X"C3",X"76",X"29",X"CD",X"83",X"2A",X"D5",X"CD",X"92",
		X"2C",X"D1",X"C9",X"3A",X"56",X"E2",X"FE",X"01",X"28",X"13",X"FE",X"02",X"28",X"0F",X"FE",X"03",
		X"28",X"1F",X"FE",X"04",X"28",X"1B",X"FE",X"05",X"20",X"20",X"C3",X"B1",X"2A",X"3A",X"17",X"E2",
		X"47",X"3A",X"56",X"E2",X"FE",X"01",X"28",X"04",X"3A",X"27",X"E2",X"47",X"78",X"E6",X"80",X"20",
		X"09",X"16",X"01",X"DD",X"35",X"0D",X"C0",X"16",X"00",X"C9",X"DD",X"7E",X"0D",X"D6",X"04",X"DD",
		X"77",X"0D",X"F2",X"C8",X"2A",X"16",X"00",X"C9",X"16",X"01",X"C9",X"3A",X"E8",X"E3",X"FE",X"01",
		X"CC",X"5C",X"33",X"3A",X"87",X"E3",X"FE",X"02",X"20",X"0C",X"CD",X"6B",X"29",X"3A",X"8D",X"E3",
		X"FE",X"00",X"CA",X"3A",X"29",X"C9",X"DD",X"21",X"E4",X"E0",X"DD",X"7E",X"02",X"FE",X"00",X"28",
		X"18",X"DD",X"7E",X"02",X"E6",X"FC",X"FE",X"28",X"28",X"0F",X"DD",X"46",X"00",X"DD",X"4E",X"03",
		X"CD",X"21",X"29",X"7A",X"FE",X"00",X"CC",X"7A",X"2C",X"DD",X"23",X"DD",X"23",X"DD",X"23",X"DD",
		X"23",X"DD",X"E5",X"E1",X"7D",X"FE",X"F4",X"20",X"06",X"DD",X"21",X"84",X"E0",X"18",X"CB",X"FE",
		X"94",X"20",X"06",X"DD",X"21",X"44",X"E1",X"18",X"C1",X"FE",X"54",X"20",X"BD",X"C3",X"3A",X"29",
		X"DD",X"7E",X"00",X"FE",X"20",X"C8",X"3E",X"30",X"DD",X"77",X"03",X"DD",X"E5",X"3E",X"05",X"CD",
		X"A0",X"33",X"3E",X"07",X"CD",X"75",X"22",X"DD",X"E1",X"DD",X"7E",X"00",X"FE",X"02",X"28",X"0D",
		X"FE",X"03",X"28",X"09",X"FE",X"04",X"28",X"05",X"FE",X"05",X"C2",X"92",X"2C",X"3A",X"25",X"E3",
		X"3C",X"32",X"25",X"E3",X"FE",X"04",X"C2",X"92",X"2C",X"3A",X"8E",X"E3",X"FE",X"01",X"CA",X"2C",
		X"2C",X"3A",X"90",X"E3",X"6F",X"3A",X"91",X"E3",X"67",X"7E",X"E6",X"FC",X"FE",X"80",X"CA",X"92",
		X"2C",X"3A",X"7A",X"E2",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"6F",X"3E",X"1F",X"95",X"3D",X"6F",
		X"26",X"80",X"DD",X"7E",X"01",X"2F",X"E6",X"F8",X"5F",X"16",X"00",X"CB",X"23",X"CB",X"12",X"CB",
		X"23",X"CB",X"12",X"19",X"DD",X"7E",X"04",X"C6",X"0C",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"85",
		X"2D",X"E6",X"1F",X"47",X"7D",X"E6",X"E0",X"B0",X"6F",X"E6",X"1F",X"FE",X"1F",X"20",X"01",X"2B",
		X"DD",X"E5",X"FD",X"E5",X"E5",X"FD",X"E1",X"DD",X"21",X"90",X"E3",X"DD",X"75",X"00",X"DD",X"74",
		X"01",X"FD",X"7E",X"00",X"DD",X"77",X"02",X"FD",X"7E",X"01",X"DD",X"77",X"03",X"FD",X"7E",X"20",
		X"DD",X"77",X"04",X"FD",X"7E",X"21",X"DD",X"77",X"05",X"3E",X"14",X"FD",X"77",X"00",X"3C",X"FD",
		X"77",X"01",X"3C",X"FD",X"77",X"20",X"3C",X"FD",X"77",X"21",X"11",X"00",X"04",X"FD",X"19",X"FD",
		X"7E",X"00",X"DD",X"77",X"06",X"FD",X"7E",X"01",X"DD",X"77",X"07",X"FD",X"7E",X"20",X"DD",X"77",
		X"08",X"FD",X"7E",X"21",X"DD",X"77",X"09",X"3E",X"18",X"FD",X"77",X"00",X"FD",X"77",X"01",X"FD",
		X"77",X"20",X"FD",X"77",X"21",X"FD",X"E1",X"DD",X"E1",X"C3",X"92",X"2C",X"3A",X"7A",X"E2",X"CB",
		X"3F",X"CB",X"3F",X"CB",X"3F",X"6F",X"3E",X"1F",X"95",X"3D",X"6F",X"26",X"80",X"DD",X"7E",X"01",
		X"2F",X"E6",X"F8",X"5F",X"16",X"00",X"CB",X"23",X"CB",X"12",X"CB",X"23",X"CB",X"12",X"19",X"DD",
		X"7E",X"04",X"C6",X"0C",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"85",X"E6",X"1F",X"47",X"7D",X"E6",
		X"E0",X"B0",X"6F",X"7E",X"FE",X"20",X"28",X"05",X"FE",X"00",X"C2",X"92",X"2C",X"3E",X"18",X"77",
		X"11",X"00",X"04",X"19",X"3E",X"1B",X"77",X"C3",X"92",X"2C",X"3E",X"07",X"CD",X"75",X"22",X"3E",
		X"28",X"DD",X"77",X"02",X"3E",X"03",X"DD",X"77",X"01",X"DD",X"E5",X"3E",X"01",X"CD",X"A0",X"33",
		X"DD",X"E1",X"3A",X"56",X"E2",X"FE",X"01",X"20",X"0F",X"3A",X"17",X"E2",X"E6",X"80",X"C0",X"3E",
		X"00",X"32",X"16",X"E2",X"32",X"17",X"E2",X"C9",X"FE",X"02",X"20",X"0F",X"3A",X"27",X"E2",X"E6",
		X"80",X"C0",X"3E",X"00",X"32",X"16",X"E2",X"32",X"17",X"E2",X"C9",X"FE",X"03",X"20",X"11",X"3E",
		X"00",X"32",X"44",X"E2",X"32",X"45",X"E2",X"32",X"46",X"E2",X"32",X"47",X"E2",X"C3",X"5B",X"39",
		X"FE",X"04",X"20",X"11",X"3E",X"00",X"32",X"48",X"E2",X"32",X"49",X"E2",X"32",X"4A",X"E2",X"32",
		X"4B",X"E2",X"C3",X"5B",X"39",X"FE",X"05",X"20",X"16",X"3E",X"00",X"32",X"07",X"E3",X"32",X"08",
		X"E3",X"32",X"09",X"E3",X"01",X"00",X"00",X"11",X"00",X"00",X"3E",X"08",X"C3",X"64",X"1C",X"C9",
		X"3A",X"1F",X"E3",X"FE",X"00",X"C0",X"3A",X"8D",X"E3",X"FE",X"00",X"28",X"06",X"3A",X"87",X"E3",
		X"FE",X"00",X"C0",X"21",X"D1",X"E2",X"35",X"C0",X"CD",X"46",X"1C",X"E6",X"0F",X"C6",X"10",X"77",
		X"3A",X"D0",X"E2",X"FE",X"00",X"C8",X"CD",X"9C",X"2E",X"FE",X"FF",X"C8",X"3A",X"D0",X"E2",X"3D",
		X"32",X"D0",X"E2",X"3E",X"01",X"DD",X"77",X"00",X"3E",X"F6",X"DD",X"77",X"04",X"3E",X"03",X"DD",
		X"77",X"02",X"3E",X"2C",X"DD",X"77",X"03",X"CD",X"46",X"1C",X"E6",X"7F",X"47",X"CD",X"46",X"1C",
		X"E6",X"1F",X"80",X"C6",X"20",X"DD",X"77",X"01",X"3E",X"01",X"DD",X"77",X"05",X"C9",X"FD",X"21",
		X"94",X"E0",X"CD",X"70",X"2D",X"FD",X"21",X"F4",X"E0",X"CD",X"70",X"2D",X"FD",X"21",X"54",X"E1",
		X"DD",X"21",X"80",X"E2",X"06",X"0A",X"11",X"08",X"00",X"DD",X"7E",X"00",X"FE",X"00",X"28",X"18",
		X"DD",X"7E",X"01",X"FD",X"77",X"00",X"DD",X"7E",X"02",X"FD",X"77",X"01",X"DD",X"7E",X"03",X"FD",
		X"77",X"02",X"DD",X"7E",X"04",X"FD",X"77",X"03",X"DD",X"19",X"FD",X"23",X"FD",X"23",X"FD",X"23",
		X"FD",X"23",X"10",X"D5",X"C9",X"21",X"D2",X"E2",X"35",X"C0",X"3A",X"02",X"E6",X"77",X"21",X"D3",
		X"E2",X"35",X"21",X"8F",X"E3",X"35",X"7E",X"3E",X"01",X"32",X"28",X"E3",X"DD",X"21",X"80",X"E2",
		X"DD",X"7E",X"00",X"FE",X"01",X"CA",X"0C",X"2E",X"FE",X"02",X"28",X"0E",X"FE",X"03",X"28",X"0A",
		X"FE",X"04",X"28",X"06",X"FE",X"05",X"28",X"02",X"18",X"13",X"DD",X"7E",X"03",X"FE",X"00",X"28",
		X"14",X"DD",X"7E",X"02",X"FE",X"00",X"28",X"0D",X"CD",X"5C",X"2F",X"18",X"08",X"FE",X"20",X"20",
		X"03",X"C3",X"F5",X"2D",X"00",X"11",X"08",X"00",X"DD",X"19",X"DD",X"E5",X"D1",X"7B",X"FE",X"D0",
		X"20",X"BE",X"3A",X"D3",X"E2",X"FE",X"00",X"C0",X"3E",X"04",X"77",X"C9",X"DD",X"35",X"05",X"20",
		X"44",X"DD",X"7E",X"03",X"FE",X"33",X"20",X"2B",X"3E",X"00",X"DD",X"77",X"00",X"DD",X"77",X"01",
		X"DD",X"77",X"02",X"DD",X"77",X"03",X"DD",X"77",X"04",X"DD",X"E5",X"E1",X"7D",X"D6",X"80",X"CB",
		X"3F",X"CB",X"3F",X"CB",X"3F",X"C6",X"0D",X"01",X"00",X"00",X"11",X"00",X"00",X"CD",X"64",X"1C",
		X"C3",X"F5",X"2D",X"E6",X"FC",X"47",X"DD",X"7E",X"03",X"3C",X"E6",X"03",X"80",X"DD",X"77",X"03",
		X"3E",X"02",X"DD",X"77",X"05",X"DD",X"7E",X"03",X"E6",X"FC",X"FE",X"30",X"20",X"03",X"C3",X"F5",
		X"2D",X"DD",X"7E",X"04",X"3D",X"3D",X"E6",X"FE",X"FE",X"F8",X"CA",X"18",X"2E",X"DD",X"77",X"04",
		X"3A",X"D3",X"E2",X"E6",X"01",X"FE",X"00",X"20",X"20",X"3A",X"11",X"E2",X"DD",X"BE",X"01",X"28",
		X"18",X"38",X"0B",X"3A",X"80",X"E3",X"DD",X"86",X"01",X"DD",X"77",X"01",X"18",X"0B",X"3A",X"80",
		X"E3",X"47",X"DD",X"7E",X"01",X"90",X"DD",X"77",X"01",X"C3",X"F5",X"2D",X"DD",X"21",X"80",X"E2",
		X"11",X"08",X"00",X"DD",X"7E",X"00",X"FE",X"00",X"C8",X"DD",X"19",X"DD",X"E5",X"E1",X"3A",X"1D",
		X"E3",X"BD",X"20",X"EF",X"3E",X"FF",X"C9",X"3A",X"8D",X"E3",X"FE",X"00",X"28",X"06",X"3A",X"87",
		X"E3",X"FE",X"00",X"C0",X"21",X"22",X"E3",X"35",X"C0",X"3A",X"A0",X"E2",X"FE",X"00",X"20",X"2A",
		X"3A",X"A8",X"E2",X"FE",X"00",X"20",X"23",X"3A",X"B0",X"E2",X"FE",X"00",X"20",X"1C",X"3A",X"B8",
		X"E2",X"FE",X"00",X"20",X"15",X"3A",X"20",X"E3",X"FE",X"02",X"20",X"0E",X"3E",X"00",X"32",X"20",
		X"E3",X"32",X"23",X"E3",X"32",X"21",X"E3",X"32",X"25",X"E3",X"3E",X"0C",X"77",X"3A",X"20",X"E3",
		X"FE",X"01",X"C0",X"3A",X"21",X"E3",X"6F",X"26",X"00",X"CB",X"25",X"CB",X"25",X"CB",X"25",X"11",
		X"A0",X"E2",X"19",X"E5",X"DD",X"E1",X"3A",X"26",X"E3",X"DD",X"77",X"00",X"3E",X"A0",X"DD",X"77",
		X"01",X"3E",X"F6",X"DD",X"77",X"04",X"06",X"03",X"3A",X"8E",X"E3",X"FE",X"00",X"28",X"02",X"06",
		X"01",X"DD",X"70",X"02",X"3A",X"24",X"E3",X"DD",X"77",X"03",X"3E",X"03",X"DD",X"77",X"05",X"3E",
		X"00",X"DD",X"77",X"06",X"3E",X"08",X"DD",X"77",X"07",X"3A",X"21",X"E3",X"3C",X"FE",X"04",X"20",
		X"07",X"3E",X"02",X"32",X"20",X"E3",X"3E",X"00",X"32",X"21",X"E3",X"C9",X"DD",X"7E",X"00",X"FE",
		X"00",X"20",X"18",X"3E",X"00",X"DD",X"77",X"01",X"DD",X"77",X"02",X"DD",X"77",X"03",X"DD",X"77",
		X"04",X"DD",X"77",X"05",X"DD",X"77",X"06",X"DD",X"77",X"07",X"C9",X"DD",X"35",X"04",X"DD",X"7E",
		X"03",X"E6",X"FC",X"FE",X"30",X"CA",X"12",X"30",X"DD",X"7E",X"05",X"FE",X"00",X"20",X"0C",X"DD",
		X"34",X"01",X"DD",X"34",X"01",X"DD",X"34",X"01",X"C3",X"12",X"30",X"FE",X"01",X"20",X"53",X"DD",
		X"34",X"04",X"DD",X"34",X"04",X"DD",X"34",X"04",X"DD",X"7E",X"02",X"E6",X"1F",X"F6",X"40",X"DD",
		X"77",X"02",X"DD",X"7E",X"04",X"E6",X"FC",X"FE",X"F8",X"20",X"57",X"3E",X"01",X"32",X"23",X"E3",
		X"3E",X"00",X"DD",X"77",X"00",X"DD",X"77",X"01",X"DD",X"77",X"02",X"DD",X"77",X"03",X"DD",X"77",
		X"04",X"DD",X"77",X"05",X"DD",X"77",X"06",X"DD",X"77",X"07",X"DD",X"E5",X"E1",X"7D",X"D6",X"80",
		X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"C6",X"0D",X"01",X"00",X"00",X"11",X"00",X"00",X"CD",X"64",
		X"1C",X"C9",X"FE",X"02",X"20",X"0B",X"DD",X"35",X"01",X"DD",X"35",X"01",X"DD",X"35",X"01",X"18",
		X"11",X"DD",X"35",X"04",X"DD",X"35",X"04",X"DD",X"35",X"04",X"DD",X"7E",X"02",X"E6",X"1F",X"DD",
		X"77",X"02",X"3A",X"28",X"E3",X"FE",X"01",X"C2",X"33",X"30",X"DD",X"7E",X"03",X"3C",X"FE",X"34",
		X"CA",X"BB",X"2F",X"DD",X"7E",X"03",X"E6",X"FC",X"47",X"DD",X"7E",X"03",X"3C",X"E6",X"03",X"80",
		X"DD",X"77",X"03",X"DD",X"35",X"07",X"C0",X"DD",X"34",X"06",X"DD",X"7E",X"00",X"D6",X"02",X"5F",
		X"16",X"00",X"CB",X"23",X"CB",X"23",X"CB",X"23",X"CB",X"23",X"CB",X"23",X"DD",X"7E",X"06",X"CB",
		X"27",X"6F",X"26",X"00",X"19",X"11",X"63",X"30",X"19",X"7E",X"DD",X"77",X"05",X"23",X"7E",X"DD",
		X"77",X"07",X"C9",X"00",X"00",X"02",X"20",X"03",X"10",X"00",X"20",X"01",X"44",X"01",X"44",X"01",
		X"44",X"01",X"44",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"04",X"03",X"04",X"00",X"02",X"01",X"02",X"02",X"20",X"03",
		X"30",X"01",X"F0",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"03",X"20",X"02",X"20",X"01",X"10",X"00",X"18",X"01",X"00",X"01",
		X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"30",X"03",X"08",X"00",X"30",X"03",X"08",X"02",X"30",X"01",
		X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"02",X"02",X"02",X"01",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"00",X"FF",
		X"00",X"00",X"00",X"3E",X"0A",X"CD",X"A0",X"33",X"CD",X"92",X"2C",X"3E",X"08",X"CD",X"75",X"22",
		X"DD",X"7E",X"02",X"C6",X"08",X"DD",X"77",X"02",X"DD",X"7E",X"06",X"C6",X"08",X"DD",X"77",X"06",
		X"DD",X"7E",X"0F",X"FE",X"00",X"28",X"08",X"3E",X"02",X"DD",X"77",X"0F",X"C3",X"76",X"29",X"3E",
		X"02",X"DD",X"77",X"0F",X"DD",X"7E",X"04",X"06",X"71",X"FE",X"73",X"28",X"09",X"FE",X"71",X"28",
		X"05",X"FE",X"70",X"28",X"01",X"47",X"78",X"DD",X"77",X"04",X"C3",X"76",X"29",X"3E",X"0A",X"CD",
		X"A0",X"33",X"CD",X"92",X"2C",X"3E",X"08",X"CD",X"75",X"22",X"DD",X"7E",X"02",X"D6",X"08",X"DD",
		X"77",X"02",X"DD",X"7E",X"06",X"D6",X"08",X"DD",X"77",X"06",X"DD",X"7E",X"0F",X"FE",X"00",X"28",
		X"08",X"3E",X"12",X"DD",X"77",X"0F",X"C3",X"76",X"29",X"3E",X"12",X"DD",X"77",X"0F",X"DD",X"7E",
		X"04",X"06",X"73",X"FE",X"73",X"28",X"09",X"FE",X"71",X"28",X"05",X"FE",X"70",X"28",X"01",X"47",
		X"78",X"DD",X"77",X"04",X"C3",X"76",X"29",X"3E",X"32",X"CD",X"A0",X"33",X"CD",X"92",X"2C",X"DD",
		X"7E",X"0F",X"FE",X"00",X"20",X"12",X"3E",X"84",X"DD",X"77",X"0F",X"3E",X"79",X"DD",X"77",X"04",
		X"3E",X"7A",X"DD",X"77",X"08",X"C3",X"76",X"29",X"3E",X"88",X"DD",X"77",X"0F",X"DD",X"7E",X"04",
		X"01",X"7C",X"7B",X"FE",X"79",X"28",X"35",X"01",X"00",X"72",X"FE",X"7B",X"20",X"0B",X"DD",X"7E",
		X"06",X"DD",X"77",X"02",X"DD",X"7E",X"04",X"18",X"23",X"3E",X"64",X"CD",X"A0",X"33",X"3E",X"05",
		X"DD",X"77",X"00",X"3E",X"49",X"DD",X"77",X"04",X"3C",X"DD",X"77",X"08",X"3E",X"03",X"DD",X"77",
		X"03",X"DD",X"77",X"07",X"3E",X"88",X"DD",X"77",X"0F",X"C3",X"76",X"29",X"DD",X"70",X"04",X"DD",
		X"71",X"08",X"C3",X"76",X"29",X"3A",X"E8",X"E3",X"FE",X"00",X"C0",X"3E",X"01",X"32",X"E8",X"E3",
		X"CD",X"46",X"1C",X"E6",X"01",X"32",X"E9",X"E3",X"CD",X"46",X"1C",X"E6",X"1F",X"06",X"50",X"80",
		X"32",X"EB",X"E3",X"3E",X"F6",X"32",X"EA",X"E3",X"3E",X"4B",X"32",X"EC",X"E3",X"CD",X"46",X"1C",
		X"E6",X"0F",X"47",X"3A",X"8C",X"E3",X"80",X"32",X"ED",X"E3",X"C9",X"DD",X"21",X"E8",X"E3",X"3A",
		X"E8",X"E3",X"FE",X"00",X"C8",X"FE",X"02",X"20",X"24",X"DD",X"35",X"05",X"C0",X"3E",X"01",X"DD",
		X"77",X"05",X"DD",X"7E",X"04",X"3C",X"FE",X"34",X"28",X"23",X"DD",X"77",X"04",X"DD",X"46",X"02",
		X"DD",X"4E",X"03",X"16",X"03",X"DD",X"5E",X"04",X"3E",X"17",X"C3",X"64",X"1C",X"DD",X"21",X"E8",
		X"E3",X"DD",X"35",X"02",X"DD",X"7E",X"02",X"E6",X"FC",X"FE",X"FC",X"20",X"1C",X"3E",X"00",X"DD",
		X"77",X"00",X"DD",X"77",X"01",X"DD",X"77",X"02",X"DD",X"77",X"03",X"32",X"E8",X"E3",X"01",X"00",
		X"00",X"11",X"00",X"00",X"3E",X"17",X"C3",X"64",X"1C",X"DD",X"35",X"06",X"DD",X"7E",X"06",X"E6",
		X"01",X"CA",X"F9",X"32",X"CD",X"46",X"1C",X"E6",X"1F",X"FE",X"10",X"20",X"08",X"DD",X"7E",X"01",
		X"EE",X"01",X"DD",X"77",X"01",X"DD",X"7E",X"01",X"FE",X"00",X"20",X"20",X"DD",X"34",X"03",X"DD",
		X"34",X"03",X"DD",X"34",X"03",X"DD",X"34",X"03",X"DD",X"7E",X"03",X"C6",X"58",X"30",X"2A",X"3E",
		X"A8",X"DD",X"77",X"03",X"3E",X"01",X"DD",X"77",X"01",X"C3",X"F9",X"32",X"DD",X"35",X"03",X"DD",
		X"35",X"03",X"DD",X"35",X"03",X"DD",X"35",X"03",X"DD",X"7E",X"03",X"C6",X"B0",X"38",X"0A",X"3E",
		X"50",X"DD",X"77",X"03",X"3E",X"00",X"DD",X"77",X"01",X"DD",X"46",X"02",X"DD",X"4E",X"03",X"16",
		X"03",X"DD",X"5E",X"04",X"3E",X"17",X"CD",X"64",X"1C",X"DD",X"35",X"05",X"C0",X"CD",X"46",X"1C",
		X"E6",X"1F",X"47",X"3A",X"8C",X"E3",X"80",X"DD",X"77",X"05",X"3A",X"7A",X"E2",X"CB",X"3F",X"CB",
		X"3F",X"CB",X"3F",X"6F",X"3E",X"1F",X"95",X"3D",X"6F",X"26",X"80",X"DD",X"7E",X"03",X"2F",X"E6",
		X"F8",X"5F",X"16",X"00",X"CB",X"23",X"CB",X"12",X"CB",X"23",X"CB",X"12",X"19",X"DD",X"7E",X"02",
		X"C6",X"0C",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"85",X"E6",X"1F",X"47",X"7D",X"E6",X"E0",X"B0",
		X"6F",X"3E",X"19",X"77",X"11",X"00",X"04",X"19",X"3E",X"19",X"77",X"C9",X"DD",X"21",X"E8",X"E3",
		X"DD",X"46",X"03",X"DD",X"4E",X"02",X"CD",X"21",X"29",X"7A",X"FE",X"00",X"C0",X"3E",X"02",X"DD",
		X"77",X"00",X"3E",X"30",X"DD",X"77",X"04",X"3E",X"02",X"DD",X"77",X"05",X"3E",X"64",X"CD",X"A0",
		X"33",X"C3",X"92",X"2C",X"3E",X"0B",X"CD",X"75",X"22",X"3E",X"01",X"E5",X"D5",X"C5",X"DD",X"E5",
		X"FD",X"E5",X"E5",X"DD",X"E1",X"CD",X"CE",X"33",X"FD",X"E1",X"DD",X"E1",X"C1",X"D1",X"E1",X"C9",
		X"E5",X"D5",X"C5",X"DD",X"E5",X"FD",X"E5",X"47",X"3A",X"01",X"E2",X"FE",X"00",X"20",X"17",X"3A",
		X"00",X"E2",X"DD",X"21",X"64",X"E2",X"FE",X"01",X"28",X"04",X"DD",X"21",X"6A",X"E2",X"CD",X"CE",
		X"33",X"10",X"FB",X"CD",X"5F",X"34",X"FD",X"E1",X"DD",X"E1",X"C1",X"D1",X"E1",X"C9",X"DD",X"E5",
		X"C5",X"06",X"05",X"DD",X"7E",X"00",X"FE",X"20",X"20",X"02",X"3E",X"30",X"3C",X"FE",X"3A",X"28",
		X"07",X"DD",X"77",X"00",X"C1",X"DD",X"E1",X"C9",X"3E",X"30",X"DD",X"77",X"00",X"DD",X"2B",X"10",
		X"E2",X"3A",X"03",X"E2",X"C6",X"02",X"32",X"03",X"E2",X"C5",X"CD",X"C6",X"37",X"06",X"10",X"C5",
		X"3E",X"06",X"CD",X"75",X"22",X"01",X"00",X"80",X"0D",X"20",X"FD",X"10",X"FB",X"C1",X"10",X"EF",
		X"3A",X"18",X"E3",X"D6",X"02",X"E6",X"1F",X"32",X"18",X"E3",X"C1",X"C1",X"DD",X"E1",X"C9",X"E5",
		X"D5",X"C5",X"DD",X"E5",X"E1",X"11",X"52",X"34",X"3A",X"02",X"E2",X"FE",X"00",X"28",X"03",X"11",
		X"58",X"34",X"2B",X"2B",X"2B",X"06",X"04",X"1A",X"BE",X"28",X"04",X"C1",X"D1",X"E1",X"C9",X"13",
		X"23",X"10",X"F4",X"3A",X"03",X"E2",X"FE",X"04",X"28",X"04",X"3C",X"32",X"03",X"E2",X"C1",X"D1",
		X"E1",X"C9",X"35",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"21",
		X"60",X"E2",X"11",X"22",X"80",X"01",X"06",X"00",X"ED",X"B0",X"21",X"66",X"E2",X"11",X"37",X"80",
		X"01",X"06",X"00",X"ED",X"B0",X"21",X"6C",X"E2",X"11",X"2D",X"80",X"01",X"06",X"00",X"ED",X"B0",
		X"C9",X"21",X"00",X"84",X"06",X"20",X"36",X"03",X"23",X"10",X"FB",X"21",X"0A",X"84",X"06",X"0A",
		X"36",X"0D",X"23",X"10",X"FB",X"21",X"20",X"84",X"06",X"1F",X"36",X"06",X"23",X"10",X"FB",X"21",
		X"2A",X"84",X"06",X"0A",X"36",X"08",X"23",X"10",X"FB",X"21",X"B7",X"34",X"11",X"01",X"80",X"01",
		X"1F",X"00",X"ED",X"B0",X"C3",X"5F",X"34",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"31",X"20",
		X"20",X"20",X"48",X"49",X"20",X"53",X"43",X"4F",X"52",X"45",X"20",X"20",X"20",X"50",X"4C",X"41",
		X"59",X"45",X"52",X"32",X"20",X"20",X"20",X"20",X"21",X"40",X"80",X"06",X"C0",X"36",X"00",X"23",
		X"10",X"FB",X"21",X"40",X"84",X"06",X"C0",X"36",X"14",X"23",X"10",X"FB",X"21",X"67",X"36",X"11",
		X"42",X"80",X"01",X"10",X"00",X"ED",X"B0",X"11",X"42",X"84",X"01",X"10",X"00",X"ED",X"B0",X"21",
		X"87",X"36",X"11",X"62",X"80",X"01",X"10",X"00",X"ED",X"B0",X"11",X"62",X"84",X"01",X"10",X"00",
		X"ED",X"B0",X"21",X"A7",X"36",X"11",X"A2",X"80",X"01",X"10",X"00",X"ED",X"B0",X"11",X"A2",X"84",
		X"01",X"10",X"00",X"ED",X"B0",X"21",X"C7",X"36",X"11",X"C2",X"80",X"01",X"10",X"00",X"ED",X"B0",
		X"11",X"C2",X"84",X"01",X"10",X"00",X"ED",X"B0",X"21",X"47",X"36",X"11",X"00",X"E0",X"01",X"14",
		X"00",X"ED",X"B0",X"21",X"FC",X"35",X"11",X"B3",X"80",X"01",X"0B",X"00",X"ED",X"B0",X"21",X"0B",
		X"36",X"11",X"B3",X"84",X"01",X"0B",X"00",X"ED",X"B0",X"21",X"35",X"36",X"11",X"87",X"80",X"01",
		X"08",X"00",X"ED",X"B0",X"21",X"3E",X"36",X"11",X"E7",X"80",X"01",X"08",X"00",X"ED",X"B0",X"21",
		X"87",X"84",X"11",X"88",X"84",X"01",X"08",X"00",X"36",X"13",X"ED",X"B0",X"21",X"E7",X"84",X"11",
		X"E8",X"84",X"01",X"08",X"00",X"36",X"13",X"ED",X"B0",X"01",X"01",X"02",X"ED",X"43",X"52",X"80",
		X"01",X"03",X"04",X"ED",X"43",X"72",X"80",X"01",X"05",X"06",X"ED",X"43",X"5D",X"80",X"01",X"07",
		X"08",X"ED",X"43",X"7D",X"80",X"01",X"1B",X"1B",X"ED",X"43",X"52",X"84",X"ED",X"43",X"72",X"84",
		X"ED",X"43",X"5D",X"84",X"ED",X"43",X"7D",X"84",X"21",X"54",X"84",X"11",X"55",X"84",X"01",X"08",
		X"00",X"36",X"1D",X"ED",X"B0",X"21",X"74",X"84",X"11",X"75",X"84",X"01",X"08",X"00",X"36",X"1D",
		X"ED",X"B0",X"21",X"29",X"36",X"11",X"98",X"80",X"01",X"03",X"00",X"ED",X"B0",X"21",X"2E",X"36",
		X"11",X"98",X"84",X"01",X"03",X"00",X"ED",X"B0",X"CD",X"E7",X"36",X"CD",X"5C",X"37",X"CD",X"20",
		X"37",X"CD",X"C6",X"37",X"21",X"2D",X"E3",X"35",X"CD",X"2C",X"22",X"C9",X"31",X"58",X"20",X"32",
		X"58",X"20",X"33",X"58",X"20",X"34",X"58",X"20",X"20",X"20",X"20",X"12",X"12",X"14",X"11",X"11",
		X"14",X"11",X"11",X"14",X"11",X"11",X"14",X"14",X"14",X"14",X"11",X"11",X"14",X"11",X"11",X"14",
		X"11",X"11",X"14",X"11",X"11",X"14",X"14",X"14",X"14",X"50",X"4F",X"57",X"20",X"20",X"13",X"13",
		X"13",X"13",X"13",X"13",X"13",X"4C",X"41",X"53",X"45",X"52",X"20",X"20",X"20",X"20",X"53",X"48",
		X"49",X"45",X"4C",X"44",X"20",X"20",X"20",X"C0",X"00",X"34",X"9C",X"C0",X"00",X"34",X"AC",X"C0",
		X"00",X"34",X"BC",X"C0",X"00",X"34",X"CC",X"C0",X"00",X"34",X"DC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"05",X"06",X"1B",X"1B",X"15",X"15",X"15",X"15",X"15",X"15",X"15",
		X"15",X"15",X"15",X"15",X"15",X"1B",X"1B",X"03",X"04",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"07",X"08",X"1B",X"1B",X"15",X"15",X"15",X"15",X"15",X"15",X"15",
		X"15",X"15",X"15",X"15",X"15",X"1B",X"1B",X"01",X"02",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"05",X"06",X"1B",X"1B",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",
		X"1C",X"1C",X"1C",X"1C",X"1C",X"1B",X"1B",X"03",X"04",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"07",X"08",X"1B",X"1B",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",
		X"1C",X"1C",X"1C",X"1C",X"1C",X"1B",X"1B",X"3A",X"05",X"E2",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",
		X"CB",X"3F",X"6F",X"26",X"00",X"11",X"49",X"37",X"19",X"7E",X"E6",X"0F",X"47",X"21",X"44",X"80",
		X"11",X"64",X"80",X"78",X"FE",X"00",X"28",X"0A",X"3E",X"10",X"77",X"3E",X"11",X"12",X"23",X"13",
		X"10",X"F1",X"7D",X"FE",X"50",X"C8",X"3E",X"12",X"77",X"3E",X"13",X"12",X"23",X"13",X"18",X"F2",
		X"3A",X"04",X"E2",X"E6",X"0F",X"47",X"21",X"54",X"80",X"11",X"74",X"80",X"78",X"FE",X"00",X"28",
		X"0A",X"3E",X"10",X"77",X"3E",X"11",X"12",X"23",X"13",X"10",X"F1",X"7D",X"FE",X"5D",X"C8",X"3E",
		X"12",X"77",X"3E",X"13",X"12",X"23",X"13",X"18",X"F2",X"00",X"01",X"02",X"03",X"04",X"05",X"06",
		X"07",X"08",X"09",X"0A",X"0B",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"3A",X"06",X"E2",X"CB",
		X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"E6",X"0F",X"6F",X"26",X"00",X"11",X"49",X"37",X"19",
		X"7E",X"47",X"21",X"A4",X"80",X"11",X"C4",X"80",X"78",X"FE",X"00",X"28",X"0A",X"3E",X"10",X"77",
		X"3E",X"11",X"12",X"23",X"13",X"10",X"F1",X"7D",X"FE",X"B0",X"C8",X"3E",X"12",X"77",X"3E",X"13",
		X"12",X"23",X"13",X"18",X"F2",X"21",X"7F",X"E2",X"35",X"C0",X"3E",X"08",X"77",X"21",X"7E",X"E2",
		X"35",X"7E",X"E6",X"07",X"6F",X"26",X"00",X"11",X"BA",X"37",X"19",X"4E",X"21",X"00",X"87",X"06",
		X"00",X"7E",X"E6",X"8F",X"B1",X"77",X"23",X"10",X"F8",X"C9",X"20",X"30",X"40",X"50",X"50",X"40",
		X"30",X"20",X"20",X"20",X"20",X"20",X"21",X"01",X"E0",X"11",X"04",X"00",X"3A",X"03",X"E2",X"47",
		X"78",X"FE",X"00",X"28",X"05",X"36",X"01",X"19",X"10",X"F6",X"7D",X"FE",X"15",X"D8",X"36",X"00",
		X"19",X"18",X"F7",X"CD",X"0C",X"39",X"C9",X"79",X"5E",X"1C",X"CB",X"22",X"19",X"ED",X"78",X"F5",
		X"D1",X"19",X"0E",X"E2",X"ED",X"79",X"C9",X"21",X"C3",X"00",X"60",X"F0",X"ED",X"79",X"CD",X"0C",
		X"39",X"3E",X"41",X"ED",X"79",X"CD",X"0C",X"39",X"ED",X"78",X"47",X"CD",X"0C",X"39",X"CD",X"E3",
		X"37",X"0E",X"E1",X"3E",X"F1",X"ED",X"79",X"CD",X"0C",X"39",X"3E",X"24",X"ED",X"79",X"CD",X"0C",
		X"39",X"ED",X"78",X"4F",X"CD",X"0C",X"39",X"C5",X"C9",X"00",X"00",X"21",X"C3",X"26",X"43",X"F2",
		X"ED",X"79",X"CD",X"0C",X"39",X"3E",X"47",X"ED",X"79",X"CD",X"0C",X"39",X"ED",X"78",X"47",X"CD",
		X"0C",X"39",X"CD",X"E3",X"37",X"0E",X"E1",X"3E",X"F3",X"ED",X"79",X"CD",X"0C",X"39",X"3E",X"2E",
		X"ED",X"79",X"CD",X"0C",X"39",X"ED",X"78",X"4F",X"CD",X"0C",X"39",X"C5",X"C9",X"00",X"00",X"00",
		X"21",X"C9",X"26",X"43",X"F0",X"ED",X"79",X"CD",X"0C",X"39",X"3E",X"01",X"ED",X"79",X"CD",X"0C",
		X"39",X"ED",X"78",X"47",X"FE",X"00",X"C8",X"31",X"00",X"20",X"C3",X"66",X"00",X"CD",X"0C",X"39",
		X"CD",X"E3",X"37",X"0E",X"E1",X"3E",X"F5",X"ED",X"79",X"CD",X"0C",X"39",X"3E",X"FF",X"ED",X"79",
		X"CD",X"0C",X"39",X"ED",X"78",X"4F",X"CD",X"0C",X"39",X"C5",X"C9",X"00",X"00",X"00",X"00",X"21",
		X"C3",X"44",X"04",X"F6",X"ED",X"79",X"CD",X"0C",X"39",X"3E",X"44",X"ED",X"79",X"CD",X"0C",X"39",
		X"ED",X"78",X"47",X"CD",X"0C",X"39",X"CD",X"E3",X"37",X"0E",X"E1",X"3E",X"F7",X"ED",X"79",X"CD",
		X"0C",X"39",X"3E",X"C4",X"ED",X"79",X"CD",X"0C",X"39",X"ED",X"78",X"4F",X"CD",X"0C",X"39",X"C5",
		X"C9",X"00",X"00",X"21",X"C3",X"34",X"04",X"F8",X"ED",X"79",X"CD",X"0C",X"39",X"3E",X"AE",X"ED",
		X"79",X"CD",X"0C",X"39",X"ED",X"78",X"47",X"CD",X"0C",X"39",X"CD",X"E3",X"37",X"0E",X"E1",X"3E",
		X"F9",X"ED",X"79",X"CD",X"0C",X"39",X"3E",X"61",X"ED",X"79",X"CD",X"0C",X"39",X"ED",X"78",X"4F",
		X"CD",X"0C",X"39",X"C5",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C9",X"3A",X"08",X"E2",X"FE",X"00",X"C8",X"3A",X"41",X"E2",X"FE",X"00",X"C8",X"3A",X"46",X"E2",
		X"FE",X"00",X"C0",X"3A",X"4A",X"E2",X"FE",X"00",X"C0",X"3E",X"01",X"32",X"46",X"E2",X"32",X"4A",
		X"E2",X"3A",X"10",X"E2",X"32",X"44",X"E2",X"32",X"48",X"E2",X"3A",X"11",X"E2",X"32",X"45",X"E2",
		X"32",X"49",X"E2",X"3E",X"0C",X"32",X"47",X"E2",X"32",X"4B",X"E2",X"3A",X"46",X"E2",X"FE",X"00",
		X"20",X"0E",X"01",X"00",X"00",X"11",X"00",X"00",X"3E",X"05",X"CD",X"64",X"1C",X"C3",X"87",X"39",
		X"1E",X"39",X"FE",X"01",X"28",X"02",X"1E",X"3D",X"16",X"02",X"3A",X"44",X"E2",X"47",X"3A",X"45",
		X"E2",X"4F",X"3E",X"05",X"CD",X"64",X"1C",X"3A",X"4A",X"E2",X"FE",X"00",X"20",X"0B",X"01",X"00",
		X"00",X"11",X"00",X"00",X"3E",X"06",X"C3",X"64",X"1C",X"1E",X"3A",X"FE",X"01",X"28",X"02",X"1E",
		X"3E",X"16",X"02",X"3A",X"48",X"E2",X"47",X"3A",X"49",X"E2",X"4F",X"3E",X"06",X"C3",X"64",X"1C",
		X"3A",X"46",X"E2",X"47",X"3A",X"4A",X"E2",X"80",X"FE",X"00",X"C8",X"CD",X"20",X"3A",X"CD",X"C4",
		X"39",X"C3",X"5B",X"39",X"DD",X"21",X"44",X"E2",X"DD",X"7E",X"02",X"FE",X"00",X"C8",X"FE",X"02",
		X"20",X"06",X"DD",X"35",X"03",X"C0",X"18",X"19",X"3A",X"10",X"E2",X"DD",X"77",X"00",X"DD",X"34",
		X"01",X"DD",X"34",X"01",X"DD",X"34",X"01",X"DD",X"34",X"01",X"DD",X"7E",X"01",X"FE",X"B0",X"38",
		X"0F",X"3E",X"00",X"DD",X"77",X"00",X"DD",X"77",X"01",X"DD",X"77",X"02",X"DD",X"77",X"03",X"C9",
		X"DD",X"35",X"03",X"28",X"EC",X"DD",X"46",X"00",X"DD",X"4E",X"01",X"CD",X"7C",X"3A",X"FE",X"20",
		X"C8",X"FE",X"00",X"C8",X"C9",X"3E",X"02",X"DD",X"77",X"02",X"3E",X"04",X"DD",X"77",X"03",X"C9",
		X"DD",X"21",X"48",X"E2",X"DD",X"7E",X"02",X"FE",X"00",X"C8",X"FE",X"02",X"20",X"06",X"DD",X"35",
		X"03",X"C0",X"18",X"19",X"3A",X"10",X"E2",X"DD",X"77",X"00",X"DD",X"35",X"01",X"DD",X"35",X"01",
		X"DD",X"35",X"01",X"DD",X"35",X"01",X"DD",X"7E",X"01",X"E6",X"F0",X"20",X"0F",X"3E",X"00",X"DD",
		X"77",X"00",X"DD",X"77",X"01",X"DD",X"77",X"02",X"DD",X"77",X"03",X"C9",X"DD",X"35",X"03",X"28",
		X"EC",X"DD",X"46",X"00",X"DD",X"4E",X"01",X"CD",X"7C",X"3A",X"FE",X"20",X"C8",X"FE",X"00",X"C8",
		X"C9",X"3E",X"02",X"DD",X"77",X"02",X"3E",X"04",X"DD",X"77",X"03",X"C9",X"79",X"2F",X"4F",X"CB",
		X"38",X"CB",X"38",X"CB",X"38",X"CB",X"39",X"CB",X"39",X"CB",X"39",X"69",X"26",X"00",X"58",X"16",
		X"00",X"06",X"05",X"CB",X"25",X"CB",X"14",X"10",X"FA",X"19",X"11",X"00",X"80",X"19",X"E5",X"C1",
		X"3A",X"7A",X"E2",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"6F",X"3E",X"1F",X"95",X"3D",X"E6",X"1F",
		X"6F",X"79",X"E6",X"1F",X"85",X"E6",X"1F",X"6F",X"79",X"E6",X"E0",X"85",X"4F",X"C5",X"E1",X"4F",
		X"7D",X"7E",X"C9",X"3A",X"42",X"E2",X"FE",X"02",X"C0",X"DD",X"21",X"00",X"E3",X"DD",X"35",X"00",
		X"20",X"0B",X"3E",X"01",X"32",X"42",X"E2",X"3E",X"34",X"DD",X"77",X"03",X"C9",X"DD",X"6E",X"00",
		X"CB",X"3D",X"26",X"00",X"11",X"F5",X"3A",X"19",X"DD",X"7E",X"01",X"96",X"DD",X"77",X"01",X"3E",
		X"38",X"DD",X"77",X"03",X"C9",X"01",X"01",X"02",X"02",X"02",X"03",X"03",X"04",X"04",X"05",X"06",
		X"07",X"08",X"08",X"08",X"3A",X"42",X"E2",X"FE",X"01",X"C0",X"DD",X"21",X"00",X"E3",X"DD",X"35",
		X"04",X"C0",X"3E",X"01",X"DD",X"77",X"04",X"DD",X"7E",X"03",X"06",X"34",X"FE",X"34",X"20",X"02",
		X"06",X"35",X"DD",X"70",X"03",X"3A",X"10",X"E2",X"D6",X"40",X"30",X"02",X"3E",X"60",X"C6",X"28",
		X"DD",X"77",X"05",X"3A",X"11",X"E2",X"C6",X"10",X"FE",X"B0",X"38",X"02",X"3E",X"B0",X"DD",X"77",
		X"06",X"3A",X"10",X"E2",X"47",X"3A",X"11",X"E2",X"C6",X"10",X"4F",X"CD",X"7C",X"3A",X"FE",X"20",
		X"28",X"0A",X"FE",X"00",X"28",X"06",X"3A",X"11",X"E2",X"DD",X"77",X"06",X"DD",X"7E",X"01",X"DD",
		X"BE",X"05",X"28",X"0A",X"30",X"05",X"DD",X"34",X"01",X"18",X"03",X"DD",X"35",X"01",X"DD",X"7E",
		X"02",X"DD",X"BE",X"06",X"28",X"0A",X"30",X"05",X"DD",X"34",X"02",X"18",X"03",X"DD",X"35",X"02",
		X"DD",X"7E",X"07",X"FE",X"00",X"C0",X"3A",X"08",X"E2",X"FE",X"00",X"C8",X"3E",X"01",X"DD",X"77",
		X"07",X"DD",X"7E",X"01",X"C6",X"08",X"DD",X"77",X"08",X"DD",X"7E",X"02",X"DD",X"77",X"09",X"3E",
		X"36",X"DD",X"77",X"0A",X"C9",X"3A",X"07",X"E3",X"FE",X"00",X"C8",X"3A",X"08",X"E3",X"3C",X"3C",
		X"3C",X"3C",X"E6",X"FC",X"FE",X"FC",X"20",X"19",X"3E",X"00",X"32",X"07",X"E3",X"32",X"08",X"E3",
		X"32",X"09",X"E3",X"32",X"0A",X"E3",X"01",X"00",X"00",X"11",X"00",X"00",X"3E",X"08",X"C3",X"64",
		X"1C",X"32",X"08",X"E3",X"3A",X"0A",X"E3",X"EE",X"01",X"32",X"0A",X"E3",X"5F",X"16",X"03",X"3A",
		X"08",X"E3",X"47",X"3A",X"09",X"E3",X"4F",X"3E",X"08",X"C3",X"64",X"1C",X"3A",X"43",X"E2",X"FE",
		X"01",X"C0",X"3A",X"10",X"E3",X"FE",X"00",X"C0",X"3A",X"08",X"E2",X"FE",X"00",X"C8",X"3E",X"01",
		X"32",X"10",X"E3",X"3A",X"10",X"E2",X"C6",X"10",X"32",X"11",X"E3",X"32",X"15",X"E3",X"3A",X"11",
		X"E2",X"32",X"12",X"E3",X"32",X"16",X"E3",X"3E",X"3B",X"32",X"13",X"E3",X"3E",X"10",X"32",X"14",
		X"E3",X"C9",X"3A",X"10",X"E3",X"FE",X"00",X"C8",X"DD",X"21",X"10",X"E3",X"DD",X"7E",X"04",X"FE",
		X"00",X"28",X"20",X"DD",X"35",X"04",X"DD",X"7E",X"02",X"3C",X"DD",X"77",X"02",X"FE",X"B0",X"38",
		X"05",X"3E",X"B0",X"DD",X"77",X"02",X"DD",X"7E",X"06",X"3D",X"FE",X"18",X"30",X"02",X"3E",X"18",
		X"DD",X"77",X"06",X"DD",X"34",X"01",X"DD",X"34",X"01",X"DD",X"34",X"01",X"DD",X"34",X"05",X"DD",
		X"34",X"05",X"DD",X"34",X"05",X"DD",X"7E",X"01",X"E6",X"FC",X"FE",X"FC",X"20",X"16",X"01",X"00",
		X"00",X"11",X"00",X"00",X"3E",X"03",X"CD",X"64",X"1C",X"3E",X"04",X"CD",X"64",X"1C",X"3E",X"00",
		X"32",X"10",X"E3",X"C9",X"DD",X"46",X"01",X"DD",X"4E",X"02",X"16",X"03",X"DD",X"5E",X"03",X"3E",
		X"03",X"CD",X"64",X"1C",X"DD",X"46",X"05",X"DD",X"4E",X"06",X"16",X"03",X"DD",X"5E",X"03",X"3E",
		X"04",X"CD",X"64",X"1C",X"C9",X"3E",X"C8",X"CD",X"A0",X"33",X"06",X"04",X"3A",X"41",X"E2",X"FE",
		X"00",X"28",X"0B",X"06",X"02",X"3A",X"42",X"E2",X"FE",X"00",X"28",X"02",X"06",X"01",X"21",X"30",
		X"E3",X"7E",X"80",X"77",X"32",X"04",X"E2",X"FE",X"08",X"C2",X"20",X"37",X"3E",X"15",X"CD",X"75",
		X"22",X"3E",X"00",X"77",X"32",X"04",X"E2",X"3A",X"31",X"E3",X"5F",X"16",X"00",X"21",X"25",X"3D",
		X"19",X"7E",X"21",X"31",X"E3",X"34",X"7E",X"FE",X"04",X"20",X"03",X"3E",X"03",X"77",X"FE",X"01",
		X"CA",X"1F",X"3D",X"FE",X"02",X"CA",X"03",X"3D",X"3E",X"01",X"32",X"43",X"E2",X"3E",X"00",X"32",
		X"10",X"E3",X"C9",X"3E",X"02",X"32",X"42",X"E2",X"3A",X"10",X"E2",X"32",X"01",X"E3",X"3A",X"11",
		X"E2",X"32",X"02",X"E3",X"3E",X"0F",X"32",X"00",X"E3",X"3E",X"38",X"32",X"03",X"E3",X"C9",X"3E",
		X"01",X"32",X"41",X"E2",X"C9",X"02",X"03",X"04",X"05",X"06",X"07",X"08",X"09",X"0A",X"0B",X"0C",
		X"0D",X"0E",X"0F",X"3E",X"00",X"32",X"4E",X"E2",X"3A",X"09",X"E2",X"FE",X"00",X"C8",X"3A",X"06",
		X"E2",X"FE",X"00",X"C8",X"3E",X"01",X"32",X"4E",X"E2",X"21",X"EA",X"E2",X"35",X"C0",X"3E",X"04",
		X"77",X"21",X"06",X"E2",X"35",X"C9",X"3A",X"EB",X"E2",X"FE",X"00",X"C8",X"21",X"EA",X"E2",X"35",
		X"C0",X"3E",X"10",X"77",X"21",X"06",X"E2",X"35",X"7E",X"FE",X"00",X"28",X"03",X"FE",X"FF",X"C0",
		X"E1",X"3E",X"FF",X"C9",X"C9",X"3A",X"07",X"E2",X"FE",X"00",X"C2",X"B1",X"3D",X"CD",X"F8",X"37",
		X"CD",X"22",X"3E",X"3A",X"07",X"E2",X"FE",X"00",X"C2",X"B1",X"3D",X"CD",X"A5",X"3F",X"CD",X"22",
		X"3E",X"3A",X"07",X"E2",X"FE",X"00",X"C2",X"B1",X"3D",X"3E",X"01",X"32",X"01",X"E2",X"CD",X"46",
		X"1C",X"E6",X"0F",X"32",X"18",X"E3",X"CD",X"47",X"07",X"3E",X"00",X"32",X"01",X"E2",X"C3",X"7D",
		X"3D",X"CD",X"5E",X"3F",X"CD",X"07",X"43",X"3A",X"07",X"E2",X"FE",X"01",X"20",X"2C",X"CD",X"68",
		X"3F",X"CD",X"76",X"3F",X"CD",X"3B",X"3E",X"FE",X"FF",X"20",X"0B",X"3A",X"07",X"E2",X"FE",X"01",
		X"C2",X"EA",X"3D",X"C3",X"C1",X"3D",X"FE",X"02",X"CA",X"C1",X"3D",X"3A",X"07",X"E2",X"FE",X"00",
		X"CA",X"B1",X"3D",X"3D",X"32",X"07",X"E2",X"3E",X"01",X"C9",X"CD",X"6F",X"3F",X"CD",X"76",X"3F",
		X"CD",X"3B",X"3E",X"FE",X"FF",X"28",X"F6",X"FE",X"02",X"CA",X"0D",X"3E",X"3A",X"07",X"E2",X"FE",
		X"00",X"CA",X"ED",X"3D",X"3D",X"E6",X"0F",X"32",X"07",X"E2",X"3E",X"01",X"C9",X"3A",X"07",X"E2",
		X"FE",X"00",X"CA",X"B1",X"3D",X"3D",X"FE",X"00",X"CA",X"05",X"3E",X"3D",X"32",X"07",X"E2",X"3E",
		X"02",X"C9",X"3E",X"00",X"32",X"01",X"E2",X"16",X"80",X"01",X"00",X"30",X"0D",X"20",X"FD",X"10",
		X"FB",X"3A",X"07",X"E2",X"FE",X"00",X"C0",X"15",X"20",X"EF",X"C9",X"16",X"10",X"D5",X"CD",X"68",
		X"18",X"D1",X"3A",X"11",X"E6",X"FE",X"00",X"28",X"03",X"3E",X"01",X"C9",X"3A",X"12",X"E6",X"FE",
		X"00",X"28",X"03",X"3E",X"02",X"C9",X"01",X"00",X"02",X"0D",X"20",X"FD",X"10",X"FB",X"15",X"20",
		X"DC",X"3E",X"FF",X"C9",X"21",X"4E",X"41",X"11",X"10",X"E4",X"01",X"E0",X"00",X"ED",X"B0",X"C9",
		X"21",X"40",X"80",X"11",X"41",X"80",X"01",X"BF",X"03",X"36",X"00",X"ED",X"B0",X"21",X"40",X"84",
		X"11",X"41",X"84",X"01",X"BF",X"03",X"36",X"00",X"ED",X"B0",X"21",X"00",X"E0",X"11",X"01",X"E0",
		X"01",X"85",X"01",X"36",X"00",X"ED",X"B0",X"C9",X"3E",X"08",X"32",X"2B",X"E3",X"CD",X"70",X"3E",
		X"CD",X"2C",X"38",X"3E",X"13",X"CD",X"75",X"22",X"CD",X"70",X"3E",X"21",X"C6",X"42",X"CD",X"FB",
		X"3F",X"21",X"F5",X"42",X"CD",X"FB",X"3F",X"CD",X"07",X"43",X"3E",X"01",X"32",X"29",X"E3",X"3E",
		X"39",X"32",X"2A",X"E3",X"CD",X"68",X"18",X"3A",X"08",X"E2",X"FE",X"00",X"20",X"F6",X"CD",X"68",
		X"18",X"3A",X"0C",X"E2",X"FE",X"00",X"C4",X"22",X"3F",X"3A",X"0D",X"E2",X"FE",X"00",X"C4",X"22",
		X"3F",X"3A",X"08",X"E2",X"FE",X"00",X"28",X"03",X"C3",X"41",X"3F",X"01",X"00",X"40",X"0D",X"20",
		X"FD",X"10",X"FB",X"21",X"2B",X"E3",X"35",X"20",X"D5",X"3E",X"0A",X"77",X"2B",X"35",X"7E",X"FE",
		X"2F",X"28",X"06",X"32",X"4F",X"82",X"C3",X"EB",X"3E",X"3E",X"00",X"C9",X"11",X"60",X"E2",X"3A",
		X"00",X"E2",X"FE",X"01",X"28",X"03",X"11",X"66",X"E2",X"21",X"57",X"09",X"01",X"06",X"00",X"ED",
		X"B0",X"C9",X"3A",X"29",X"E3",X"FE",X"01",X"28",X"0C",X"21",X"F5",X"42",X"CD",X"FB",X"3F",X"3E",
		X"01",X"32",X"29",X"E3",X"C9",X"21",X"FE",X"42",X"CD",X"FB",X"3F",X"3E",X"00",X"32",X"29",X"E3",
		X"C9",X"3A",X"29",X"E3",X"FE",X"00",X"CA",X"5B",X"3F",X"3A",X"07",X"E2",X"FE",X"00",X"CA",X"CE",
		X"3E",X"3D",X"32",X"07",X"E2",X"CD",X"0C",X"3F",X"3E",X"01",X"C9",X"3E",X"00",X"C9",X"CD",X"70",
		X"3E",X"21",X"FE",X"41",X"CD",X"FB",X"3F",X"C9",X"21",X"85",X"42",X"CD",X"FB",X"3F",X"C9",X"21",
		X"A6",X"42",X"CD",X"FB",X"3F",X"C9",X"21",X"C1",X"86",X"11",X"C2",X"86",X"3A",X"C8",X"86",X"06",
		X"0C",X"FE",X"01",X"28",X"18",X"06",X"07",X"FE",X"04",X"28",X"12",X"06",X"01",X"FE",X"07",X"28",
		X"0C",X"06",X"05",X"FE",X"0C",X"28",X"06",X"06",X"04",X"FE",X"05",X"28",X"00",X"78",X"06",X"1F",
		X"77",X"23",X"10",X"FC",X"C9",X"CD",X"70",X"3E",X"21",X"CD",X"40",X"CD",X"FB",X"3F",X"CD",X"B5",
		X"3F",X"CD",X"07",X"43",X"C9",X"21",X"10",X"E4",X"11",X"A8",X"81",X"06",X"0A",X"C5",X"E5",X"D5",
		X"21",X"00",X"04",X"19",X"EB",X"21",X"EE",X"41",X"01",X"0F",X"00",X"ED",X"B0",X"D1",X"E1",X"01",
		X"10",X"00",X"ED",X"B0",X"E5",X"EB",X"11",X"10",X"00",X"19",X"EB",X"E1",X"C1",X"10",X"DE",X"C9",
		X"21",X"00",X"E0",X"11",X"01",X"E0",X"01",X"90",X"01",X"36",X"00",X"ED",X"B0",X"21",X"00",X"80",
		X"11",X"01",X"80",X"01",X"FF",X"07",X"36",X"00",X"ED",X"B0",X"C9",X"4E",X"23",X"56",X"23",X"5E",
		X"23",X"7E",X"FE",X"FF",X"C8",X"FE",X"FE",X"20",X"05",X"23",X"4E",X"23",X"18",X"F3",X"FE",X"FD",
		X"20",X"07",X"23",X"56",X"23",X"5E",X"23",X"18",X"E8",X"12",X"E5",X"21",X"00",X"04",X"19",X"71",
		X"E1",X"13",X"23",X"C3",X"01",X"40",X"CD",X"E0",X"3F",X"CD",X"81",X"34",X"21",X"36",X"40",X"CD",
		X"FB",X"3F",X"CD",X"07",X"43",X"C9",X"03",X"81",X"8A",X"50",X"52",X"4F",X"47",X"52",X"41",X"4D",
		X"4D",X"45",X"44",X"20",X"42",X"59",X"FD",X"82",X"0A",X"FE",X"06",X"4B",X"59",X"4C",X"45",X"20",
		X"48",X"4F",X"44",X"47",X"45",X"54",X"54",X"53",X"FD",X"82",X"4A",X"54",X"4F",X"4E",X"59",X"20",
		X"20",X"57",X"49",X"4E",X"44",X"53",X"4F",X"52",X"FD",X"82",X"CB",X"FE",X"01",X"49",X"4E",X"53",
		X"45",X"52",X"54",X"20",X"43",X"4F",X"49",X"4E",X"FD",X"83",X"4D",X"FE",X"0B",X"43",X"20",X"31",
		X"39",X"38",X"38",X"FD",X"83",X"87",X"FE",X"0A",X"56",X"49",X"53",X"49",X"4F",X"4E",X"20",X"45",
		X"4C",X"45",X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",X"53",X"FE",X"10",X"FD",X"80",X"C7",X"80",
		X"81",X"82",X"83",X"84",X"85",X"86",X"87",X"80",X"81",X"00",X"00",X"88",X"89",X"8A",X"8B",X"8C",
		X"8D",X"FE",X"1A",X"FD",X"80",X"E7",X"8E",X"8F",X"90",X"91",X"92",X"93",X"94",X"95",X"8E",X"8F",
		X"00",X"00",X"96",X"97",X"98",X"99",X"9A",X"9B",X"FF",X"FF",X"FF",X"FF",X"FF",X"10",X"80",X"C7",
		X"80",X"81",X"82",X"83",X"84",X"85",X"86",X"87",X"80",X"81",X"00",X"00",X"88",X"89",X"8A",X"8B",
		X"8C",X"8D",X"FE",X"1A",X"FD",X"80",X"E7",X"8E",X"8F",X"90",X"91",X"92",X"93",X"94",X"95",X"8E",
		X"8F",X"00",X"00",X"96",X"97",X"98",X"99",X"9A",X"9B",X"FE",X"02",X"FD",X"81",X"2D",X"54",X"4F",
		X"50",X"20",X"54",X"45",X"4E",X"FD",X"81",X"4E",X"41",X"4C",X"49",X"45",X"4E",X"FD",X"81",X"6D",
		X"4B",X"49",X"43",X"4B",X"45",X"52",X"53",X"FE",X"01",X"FD",X"83",X"0B",X"49",X"4E",X"53",X"45",
		X"52",X"54",X"20",X"43",X"4F",X"49",X"4E",X"FD",X"83",X"4D",X"FE",X"0B",X"43",X"20",X"31",X"39",
		X"38",X"38",X"FD",X"83",X"87",X"FE",X"0A",X"56",X"49",X"53",X"49",X"4F",X"4E",X"20",X"45",X"4C",
		X"45",X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",X"53",X"FF",X"FF",X"FF",X"FF",X"FF",X"20",X"31",
		X"2E",X"20",X"35",X"30",X"30",X"30",X"30",X"30",X"20",X"20",X"4B",X"2E",X"48",X"20",X"20",X"32",
		X"2E",X"20",X"34",X"30",X"30",X"30",X"30",X"30",X"20",X"20",X"54",X"2E",X"57",X"20",X"20",X"33",
		X"2E",X"20",X"33",X"30",X"30",X"30",X"30",X"30",X"20",X"20",X"42",X"47",X"4A",X"20",X"20",X"34",
		X"2E",X"20",X"32",X"30",X"30",X"30",X"30",X"30",X"20",X"20",X"42",X"4F",X"42",X"20",X"20",X"35",
		X"2E",X"20",X"31",X"30",X"30",X"30",X"30",X"30",X"20",X"20",X"52",X"4F",X"4E",X"20",X"20",X"36",
		X"2E",X"20",X"20",X"35",X"30",X"30",X"30",X"30",X"20",X"20",X"2E",X"2E",X"2E",X"20",X"20",X"37",
		X"2E",X"20",X"20",X"34",X"30",X"30",X"30",X"30",X"20",X"20",X"50",X"43",X"51",X"20",X"20",X"38",
		X"2E",X"20",X"20",X"33",X"30",X"30",X"30",X"30",X"20",X"20",X"41",X"2E",X"50",X"20",X"20",X"39",
		X"2E",X"20",X"20",X"31",X"30",X"30",X"30",X"30",X"20",X"20",X"50",X"48",X"4C",X"20",X"31",X"30",
		X"2E",X"20",X"20",X"20",X"35",X"30",X"30",X"30",X"20",X"20",X"49",X"56",X"4E",X"20",X"06",X"06",
		X"06",X"06",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"09",X"09",X"09",X"09",X"03",X"81",
		X"8A",X"50",X"52",X"4F",X"47",X"52",X"41",X"4D",X"4D",X"45",X"44",X"20",X"42",X"59",X"FD",X"82",
		X"0A",X"FE",X"06",X"4B",X"59",X"4C",X"45",X"20",X"48",X"4F",X"44",X"47",X"45",X"54",X"54",X"53",
		X"FD",X"82",X"4A",X"54",X"4F",X"4E",X"59",X"20",X"20",X"57",X"49",X"4E",X"44",X"53",X"4F",X"52",
		X"FD",X"83",X"4D",X"FE",X"0B",X"43",X"20",X"31",X"39",X"38",X"38",X"FD",X"83",X"87",X"FE",X"0A",
		X"56",X"49",X"53",X"49",X"4F",X"4E",X"20",X"45",X"4C",X"45",X"43",X"54",X"52",X"4F",X"4E",X"49",
		X"43",X"53",X"FE",X"10",X"FD",X"80",X"C7",X"80",X"81",X"82",X"83",X"84",X"85",X"86",X"87",X"80",
		X"81",X"00",X"00",X"88",X"89",X"8A",X"8B",X"8C",X"8D",X"FE",X"1A",X"FD",X"80",X"E7",X"8E",X"8F",
		X"90",X"91",X"92",X"93",X"94",X"95",X"8E",X"8F",X"00",X"00",X"96",X"97",X"98",X"99",X"9A",X"9B",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"82",X"C2",X"50",X"52",X"45",X"53",X"53",X"20",X"4F",X"4E",
		X"45",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"20",X"42",X"55",X"54",X"54",X"4F",X"4E",X"20",
		X"4F",X"4E",X"4C",X"59",X"FF",X"FF",X"01",X"82",X"C2",X"20",X"20",X"50",X"52",X"45",X"53",X"53",
		X"20",X"4F",X"4E",X"45",X"20",X"4F",X"52",X"20",X"54",X"57",X"4F",X"20",X"50",X"4C",X"41",X"59",
		X"45",X"52",X"53",X"20",X"20",X"FF",X"05",X"80",X"E9",X"43",X"4F",X"4E",X"54",X"49",X"4E",X"55",
		X"45",X"20",X"50",X"4C",X"41",X"59",X"FE",X"0C",X"FD",X"81",X"4E",X"59",X"45",X"53",X"FE",X"01",
		X"FD",X"81",X"CB",X"50",X"52",X"45",X"53",X"53",X"20",X"46",X"49",X"52",X"45",X"FE",X"06",X"FD",
		X"82",X"4F",X"39",X"FF",X"FF",X"0C",X"81",X"4E",X"59",X"45",X"53",X"20",X"FF",X"FF",X"0C",X"81",
		X"4E",X"4E",X"4F",X"20",X"20",X"FF",X"FF",X"21",X"37",X"45",X"11",X"F4",X"83",X"01",X"0A",X"00",
		X"ED",X"B0",X"21",X"43",X"45",X"11",X"F4",X"87",X"01",X"0A",X"00",X"ED",X"B0",X"3A",X"07",X"E2",
		X"C6",X"30",X"32",X"FC",X"83",X"C9",X"DD",X"21",X"60",X"E2",X"3A",X"00",X"E2",X"FE",X"01",X"28",
		X"04",X"DD",X"21",X"66",X"E2",X"3E",X"00",X"32",X"ED",X"E2",X"FD",X"21",X"14",X"E4",X"DD",X"E5",
		X"FD",X"E5",X"06",X"05",X"DD",X"7E",X"00",X"FD",X"BE",X"00",X"28",X"0B",X"FE",X"00",X"28",X"07",
		X"FD",X"BE",X"00",X"30",X"1B",X"18",X"06",X"DD",X"23",X"FD",X"23",X"10",X"E7",X"FD",X"E1",X"DD",
		X"E1",X"11",X"10",X"00",X"FD",X"19",X"21",X"ED",X"E2",X"34",X"7E",X"FE",X"0A",X"20",X"CF",X"C9",
		X"3E",X"12",X"CD",X"75",X"22",X"FD",X"E1",X"DD",X"E1",X"FD",X"E5",X"E1",X"7D",X"FE",X"14",X"20",
		X"0B",X"DD",X"E5",X"E1",X"11",X"6C",X"E2",X"01",X"06",X"00",X"ED",X"B0",X"3A",X"ED",X"E2",X"CB",
		X"27",X"CB",X"27",X"CB",X"27",X"6F",X"26",X"00",X"11",X"CD",X"44",X"19",X"56",X"23",X"5E",X"23",
		X"46",X"23",X"4E",X"D5",X"23",X"56",X"23",X"5E",X"EB",X"D1",X"E5",X"21",X"10",X"00",X"19",X"EB",
		X"E5",X"09",X"EB",X"09",X"EB",X"ED",X"B8",X"E1",X"11",X"0B",X"00",X"19",X"FD",X"22",X"ED",X"E2",
		X"FD",X"E5",X"D1",X"DD",X"E5",X"E1",X"01",X"06",X"00",X"ED",X"B0",X"EB",X"23",X"23",X"DD",X"E1",
		X"E5",X"FD",X"E1",X"3E",X"31",X"E5",X"D5",X"21",X"11",X"E4",X"11",X"10",X"00",X"06",X"09",X"3E",
		X"31",X"77",X"E5",X"F5",X"23",X"36",X"2E",X"23",X"36",X"00",X"F1",X"E1",X"3C",X"19",X"10",X"F1",
		X"2B",X"36",X"31",X"23",X"36",X"30",X"D1",X"E1",X"CD",X"70",X"3E",X"CD",X"B5",X"3F",X"21",X"25",
		X"45",X"CD",X"FB",X"3F",X"DD",X"E5",X"D1",X"21",X"00",X"04",X"19",X"EB",X"D5",X"E1",X"2B",X"36",
		X"0C",X"01",X"18",X"00",X"ED",X"B0",X"11",X"0C",X"00",X"DD",X"19",X"3E",X"41",X"DD",X"77",X"00",
		X"DD",X"77",X"01",X"DD",X"77",X"02",X"FD",X"77",X"00",X"FD",X"77",X"01",X"FD",X"77",X"02",X"3E",
		X"03",X"32",X"ED",X"E2",X"CD",X"68",X"18",X"3A",X"0D",X"E2",X"FE",X"00",X"28",X"15",X"DD",X"34",
		X"00",X"DD",X"7E",X"00",X"FE",X"5F",X"20",X"02",X"3E",X"41",X"DD",X"77",X"00",X"FD",X"77",X"00",
		X"C3",X"85",X"44",X"3A",X"0C",X"E2",X"FE",X"00",X"28",X"15",X"DD",X"35",X"00",X"DD",X"7E",X"00",
		X"FE",X"40",X"20",X"02",X"3E",X"5E",X"DD",X"77",X"00",X"FD",X"77",X"00",X"C3",X"85",X"44",X"3A",
		X"08",X"E2",X"FE",X"00",X"CA",X"34",X"44",X"DD",X"23",X"FD",X"23",X"21",X"ED",X"E2",X"35",X"C2",
		X"9B",X"44",X"C3",X"B4",X"44",X"DD",X"E5",X"E1",X"11",X"00",X"04",X"19",X"7E",X"EE",X"08",X"77",
		X"01",X"00",X"40",X"0D",X"20",X"FD",X"10",X"FB",X"C3",X"34",X"44",X"DD",X"E5",X"E1",X"11",X"00",
		X"04",X"19",X"7E",X"EE",X"08",X"77",X"01",X"00",X"80",X"0D",X"20",X"FD",X"10",X"FB",X"01",X"00",
		X"40",X"C3",X"93",X"44",X"CD",X"B5",X"3F",X"3E",X"04",X"01",X"00",X"00",X"0D",X"20",X"FD",X"10",
		X"FB",X"3D",X"20",X"F8",X"CD",X"81",X"34",X"3E",X"11",X"CD",X"75",X"22",X"C9",X"E4",X"10",X"00",
		X"E0",X"81",X"A8",X"00",X"00",X"E4",X"20",X"00",X"D0",X"81",X"C8",X"00",X"00",X"E4",X"30",X"00",
		X"C0",X"81",X"E8",X"00",X"00",X"E4",X"40",X"00",X"B0",X"82",X"08",X"00",X"00",X"E4",X"50",X"00",
		X"A0",X"82",X"28",X"00",X"00",X"E4",X"60",X"00",X"90",X"82",X"48",X"00",X"00",X"E4",X"70",X"00",
		X"80",X"82",X"68",X"00",X"00",X"E4",X"80",X"00",X"70",X"82",X"88",X"00",X"00",X"E4",X"90",X"00",
		X"60",X"82",X"A8",X"00",X"00",X"E4",X"A0",X"00",X"50",X"82",X"C8",X"00",X"00",X"E4",X"B0",X"00",
		X"40",X"82",X"E8",X"00",X"00",X"0C",X"83",X"09",X"45",X"4E",X"54",X"45",X"52",X"20",X"49",X"4E",
		X"20",X"4E",X"41",X"4D",X"45",X"FF",X"FF",X"43",X"52",X"45",X"44",X"49",X"54",X"53",X"20",X"20",
		X"20",X"20",X"20",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",
		X"04",X"04",X"C0",X"05",X"88",X"1F",X"01",X"01",X"1E",X"02",X"04",X"1D",X"03",X"04",X"E0",X"05",
		X"98",X"22",X"04",X"01",X"40",X"04",X"01",X"80",X"04",X"01",X"B0",X"04",X"01",X"60",X"08",X"01",
		X"98",X"08",X"01",X"D1",X"08",X"01",X"77",X"09",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"20",X"05",X"98",X"1F",X"01",X"01",X"1E",X"02",X"04",X"1D",X"03",X"04",X"40",X"05",
		X"98",X"10",X"04",X"01",X"55",X"04",X"01",X"82",X"04",X"01",X"B6",X"04",X"01",X"E2",X"04",X"01",
		X"31",X"08",X"01",X"68",X"08",X"01",X"98",X"08",X"01",X"C8",X"08",X"01",X"FE",X"08",X"01",X"E0",
		X"06",X"05",X"01",X"0D",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"20",X"05",X"98",X"1F",X"01",X"01",X"1E",X"02",X"04",X"1D",X"03",X"04",X"40",X"05",
		X"98",X"10",X"04",X"01",X"55",X"04",X"01",X"82",X"04",X"01",X"B6",X"04",X"01",X"E2",X"04",X"01",
		X"31",X"08",X"01",X"68",X"08",X"01",X"98",X"08",X"01",X"C8",X"08",X"01",X"F2",X"07",X"01",X"08",
		X"06",X"05",X"01",X"0D",X"04",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"C0",X"05",X"88",X"1F",X"01",X"01",X"1E",X"02",X"04",X"1D",X"03",X"04",X"E0",X"05",
		X"98",X"22",X"04",X"01",X"40",X"04",X"01",X"80",X"04",X"01",X"B0",X"04",X"01",X"60",X"08",X"01",
		X"98",X"08",X"01",X"D1",X"08",X"01",X"33",X"08",X"04",X"09",X"06",X"01",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"20",X"05",X"98",X"1F",X"01",X"01",X"1E",X"02",X"04",X"1D",X"03",X"04",X"40",X"05",
		X"98",X"10",X"04",X"01",X"55",X"04",X"01",X"82",X"04",X"01",X"B6",X"04",X"01",X"E2",X"04",X"01",
		X"31",X"08",X"01",X"68",X"08",X"01",X"98",X"08",X"01",X"C8",X"08",X"01",X"FE",X"08",X"01",X"E0",
		X"07",X"05",X"01",X"0D",X"01",X"55",X"06",X"22",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"20",X"05",X"98",X"1F",X"01",X"01",X"1E",X"02",X"04",X"1D",X"03",X"04",X"40",X"05",
		X"98",X"10",X"04",X"01",X"55",X"04",X"01",X"82",X"04",X"01",X"B6",X"04",X"01",X"E2",X"04",X"01",
		X"31",X"08",X"01",X"68",X"08",X"01",X"98",X"08",X"01",X"C8",X"08",X"01",X"FE",X"08",X"01",X"44",
		X"07",X"05",X"01",X"0D",X"04",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"C0",X"05",X"88",X"1F",X"01",X"01",X"1E",X"02",X"04",X"1D",X"03",X"04",X"E0",X"05",
		X"98",X"22",X"04",X"01",X"40",X"04",X"01",X"80",X"04",X"01",X"B0",X"04",X"01",X"60",X"08",X"01",
		X"98",X"08",X"01",X"D1",X"08",X"01",X"77",X"09",X"00",X"57",X"07",X"02",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"20",X"05",X"98",X"1F",X"01",X"01",X"1E",X"02",X"04",X"1D",X"03",X"04",X"40",X"05",
		X"98",X"10",X"04",X"01",X"55",X"04",X"01",X"82",X"04",X"01",X"B6",X"04",X"01",X"E2",X"04",X"01",
		X"31",X"08",X"01",X"68",X"08",X"01",X"98",X"08",X"01",X"C8",X"08",X"01",X"FE",X"08",X"01",X"E0",
		X"06",X"05",X"01",X"0D",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"20",X"05",X"98",X"1F",X"01",X"01",X"1E",X"02",X"04",X"1D",X"03",X"04",X"40",X"05",
		X"98",X"10",X"04",X"01",X"55",X"04",X"01",X"82",X"04",X"01",X"B6",X"04",X"01",X"E2",X"04",X"01",
		X"31",X"08",X"01",X"68",X"08",X"01",X"98",X"08",X"01",X"C8",X"08",X"01",X"F2",X"07",X"01",X"08",
		X"06",X"05",X"01",X"0D",X"04",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"C0",X"05",X"88",X"1F",X"01",X"01",X"1E",X"02",X"04",X"1D",X"03",X"04",X"E0",X"05",
		X"98",X"22",X"04",X"01",X"40",X"04",X"01",X"80",X"04",X"01",X"B0",X"04",X"01",X"60",X"08",X"01",
		X"98",X"08",X"01",X"D1",X"08",X"01",X"33",X"08",X"04",X"09",X"06",X"01",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"20",X"05",X"98",X"1F",X"01",X"01",X"1E",X"02",X"04",X"1D",X"03",X"04",X"40",X"05",
		X"98",X"10",X"04",X"01",X"55",X"04",X"01",X"82",X"04",X"01",X"B6",X"04",X"01",X"E2",X"04",X"01",
		X"31",X"08",X"01",X"68",X"08",X"01",X"98",X"08",X"01",X"C8",X"08",X"01",X"FE",X"08",X"01",X"E0",
		X"07",X"05",X"01",X"0D",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"20",X"05",X"98",X"1F",X"01",X"01",X"1E",X"02",X"04",X"1D",X"03",X"04",X"40",X"05",
		X"98",X"10",X"04",X"01",X"55",X"04",X"01",X"82",X"04",X"01",X"B6",X"04",X"01",X"E2",X"04",X"01",
		X"31",X"08",X"01",X"68",X"08",X"01",X"98",X"08",X"01",X"C8",X"08",X"01",X"FE",X"08",X"01",X"44",
		X"06",X"05",X"01",X"0D",X"04",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"C0",X"05",X"88",X"1F",X"01",X"01",X"1E",X"02",X"04",X"1D",X"03",X"04",X"E0",X"05",
		X"98",X"22",X"04",X"01",X"40",X"04",X"01",X"80",X"04",X"01",X"B0",X"04",X"01",X"60",X"08",X"01",
		X"98",X"08",X"01",X"D1",X"08",X"01",X"77",X"09",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"20",X"05",X"98",X"1F",X"01",X"01",X"1E",X"02",X"04",X"1D",X"03",X"04",X"40",X"05",
		X"98",X"10",X"04",X"01",X"55",X"04",X"01",X"82",X"04",X"01",X"B6",X"04",X"01",X"E2",X"04",X"01",
		X"31",X"08",X"01",X"68",X"08",X"01",X"98",X"08",X"01",X"C8",X"08",X"01",X"FE",X"08",X"01",X"E0",
		X"06",X"05",X"01",X"0D",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"20",X"05",X"98",X"1F",X"01",X"01",X"1E",X"02",X"04",X"1D",X"03",X"04",X"40",X"05",
		X"98",X"10",X"04",X"01",X"55",X"04",X"01",X"82",X"04",X"01",X"B6",X"04",X"01",X"E2",X"04",X"01",
		X"31",X"08",X"01",X"68",X"08",X"01",X"98",X"08",X"01",X"C8",X"08",X"01",X"F2",X"07",X"01",X"08",
		X"06",X"05",X"01",X"0D",X"04",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"C0",X"05",X"88",X"1F",X"01",X"01",X"1E",X"02",X"04",X"1D",X"03",X"04",X"E0",X"05",
		X"98",X"22",X"04",X"01",X"40",X"04",X"01",X"80",X"04",X"01",X"B0",X"04",X"01",X"60",X"08",X"01",
		X"98",X"08",X"01",X"D1",X"08",X"01",X"33",X"08",X"04",X"09",X"06",X"01",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"20",X"05",X"98",X"1F",X"01",X"01",X"1E",X"02",X"04",X"1D",X"03",X"04",X"40",X"05",
		X"98",X"10",X"04",X"01",X"55",X"04",X"01",X"82",X"04",X"01",X"B6",X"04",X"01",X"E2",X"04",X"01",
		X"31",X"08",X"01",X"68",X"08",X"01",X"98",X"08",X"01",X"C8",X"08",X"01",X"FE",X"08",X"01",X"E0",
		X"07",X"05",X"01",X"0D",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"20",X"05",X"98",X"1F",X"01",X"01",X"1E",X"02",X"04",X"1D",X"03",X"04",X"40",X"05",
		X"98",X"10",X"04",X"01",X"55",X"04",X"01",X"82",X"04",X"01",X"B6",X"04",X"01",X"E2",X"04",X"01",
		X"31",X"08",X"01",X"68",X"08",X"01",X"98",X"08",X"01",X"C8",X"08",X"01",X"FE",X"08",X"01",X"44",
		X"06",X"05",X"01",X"0D",X"04",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"C0",X"05",X"88",X"1F",X"01",X"01",X"1E",X"02",X"04",X"1D",X"03",X"04",X"E0",X"05",
		X"98",X"22",X"04",X"01",X"40",X"04",X"01",X"80",X"04",X"01",X"B0",X"04",X"01",X"60",X"08",X"01",
		X"98",X"08",X"01",X"D1",X"08",X"01",X"77",X"09",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"20",X"05",X"98",X"1F",X"01",X"01",X"1E",X"02",X"04",X"1D",X"03",X"04",X"40",X"05",
		X"98",X"10",X"04",X"01",X"55",X"04",X"01",X"82",X"04",X"01",X"B6",X"04",X"01",X"E2",X"04",X"01",
		X"31",X"08",X"01",X"68",X"08",X"01",X"98",X"08",X"01",X"C8",X"08",X"01",X"FE",X"08",X"01",X"E0",
		X"06",X"05",X"01",X"0D",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"20",X"05",X"98",X"1F",X"01",X"01",X"1E",X"02",X"04",X"1D",X"03",X"04",X"40",X"05",
		X"98",X"10",X"04",X"01",X"55",X"04",X"01",X"82",X"04",X"01",X"B6",X"04",X"01",X"E2",X"04",X"01",
		X"31",X"08",X"01",X"68",X"08",X"01",X"98",X"08",X"01",X"C8",X"08",X"01",X"F2",X"07",X"01",X"08",
		X"06",X"05",X"01",X"0D",X"04",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"C0",X"05",X"88",X"1F",X"01",X"01",X"1E",X"02",X"04",X"1D",X"03",X"04",X"E0",X"05",
		X"98",X"22",X"04",X"01",X"40",X"04",X"01",X"80",X"04",X"01",X"B0",X"04",X"01",X"60",X"08",X"01",
		X"98",X"08",X"01",X"D1",X"08",X"01",X"33",X"08",X"04",X"09",X"06",X"01",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"20",X"05",X"98",X"1F",X"01",X"01",X"1E",X"02",X"04",X"1D",X"03",X"04",X"40",X"05",
		X"98",X"10",X"04",X"01",X"55",X"04",X"01",X"82",X"04",X"01",X"B6",X"04",X"01",X"E2",X"04",X"01",
		X"31",X"08",X"01",X"68",X"08",X"01",X"98",X"08",X"01",X"C8",X"08",X"01",X"FE",X"08",X"01",X"E0",
		X"07",X"05",X"01",X"0D",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"20",X"05",X"98",X"1F",X"01",X"01",X"1E",X"02",X"04",X"1D",X"03",X"04",X"40",X"05",
		X"98",X"10",X"04",X"01",X"55",X"04",X"01",X"82",X"04",X"01",X"B6",X"04",X"01",X"E2",X"04",X"01",
		X"31",X"08",X"01",X"68",X"08",X"01",X"98",X"08",X"01",X"C8",X"08",X"01",X"FE",X"08",X"01",X"44",
		X"06",X"05",X"01",X"0D",X"04",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"20",X"05",X"98",X"1F",X"01",X"01",X"1E",X"02",X"04",X"1D",X"03",X"04",X"40",X"05",
		X"98",X"10",X"04",X"01",X"55",X"04",X"01",X"82",X"04",X"01",X"B6",X"04",X"01",X"E2",X"04",X"01",
		X"31",X"08",X"01",X"68",X"08",X"01",X"98",X"08",X"01",X"C8",X"08",X"01",X"FE",X"08",X"01",X"E0",
		X"06",X"05",X"01",X"0D",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"20",X"05",X"98",X"1F",X"01",X"01",X"1E",X"02",X"04",X"1D",X"03",X"04",X"40",X"05",
		X"98",X"10",X"04",X"01",X"55",X"04",X"01",X"82",X"04",X"01",X"B6",X"04",X"01",X"E2",X"04",X"01",
		X"31",X"08",X"01",X"68",X"08",X"01",X"98",X"08",X"01",X"C8",X"08",X"01",X"F2",X"07",X"01",X"08",
		X"06",X"05",X"01",X"0D",X"04",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"C0",X"05",X"88",X"1F",X"01",X"01",X"1E",X"02",X"04",X"1D",X"03",X"04",X"E0",X"05",
		X"98",X"22",X"04",X"01",X"40",X"04",X"01",X"80",X"04",X"01",X"B0",X"04",X"01",X"60",X"08",X"01",
		X"98",X"08",X"01",X"D1",X"08",X"01",X"33",X"08",X"04",X"09",X"06",X"01",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"20",X"05",X"98",X"1F",X"01",X"01",X"1E",X"02",X"04",X"1D",X"03",X"04",X"40",X"05",
		X"98",X"10",X"04",X"01",X"55",X"04",X"01",X"82",X"04",X"01",X"B6",X"04",X"01",X"E2",X"04",X"01",
		X"31",X"08",X"01",X"68",X"08",X"01",X"98",X"08",X"01",X"C8",X"08",X"01",X"FE",X"08",X"01",X"E0",
		X"07",X"05",X"01",X"0D",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"20",X"05",X"98",X"1F",X"01",X"01",X"1E",X"02",X"04",X"1D",X"03",X"04",X"40",X"05",
		X"98",X"10",X"04",X"01",X"55",X"04",X"01",X"82",X"04",X"01",X"B6",X"04",X"01",X"E2",X"04",X"01",
		X"31",X"08",X"01",X"68",X"08",X"01",X"98",X"08",X"01",X"C8",X"08",X"01",X"FE",X"08",X"01",X"44",
		X"06",X"05",X"01",X"0D",X"04",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"C0",X"05",X"88",X"1F",X"01",X"01",X"1E",X"02",X"04",X"1D",X"03",X"04",X"E0",X"05",
		X"98",X"22",X"04",X"01",X"40",X"04",X"01",X"80",X"04",X"01",X"B0",X"04",X"01",X"60",X"08",X"01",
		X"98",X"08",X"01",X"D1",X"08",X"01",X"77",X"09",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"20",X"05",X"98",X"1F",X"01",X"01",X"1E",X"02",X"04",X"1D",X"03",X"04",X"40",X"05",
		X"98",X"10",X"04",X"01",X"55",X"04",X"01",X"82",X"04",X"01",X"B6",X"04",X"01",X"E2",X"04",X"01",
		X"31",X"08",X"01",X"68",X"08",X"01",X"98",X"08",X"01",X"C8",X"08",X"01",X"FE",X"08",X"01",X"E0",
		X"06",X"05",X"01",X"0D",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"05",X"14",X"0F",X"04",X"02",X"03",X"12",X"06",X"07",X"37",X"38",X"00",X"11",X"02",X"03",X"00",
		X"04",X"37",X"38",X"0A",X"0F",X"02",X"03",X"06",X"07",X"37",X"38",X"08",X"09",X"08",X"37",X"38",
		X"34",X"24",X"24",X"26",X"24",X"24",X"26",X"24",X"37",X"38",X"24",X"14",X"24",X"24",X"2F",X"24",
		X"37",X"38",X"00",X"00",X"24",X"24",X"26",X"24",X"37",X"38",X"25",X"26",X"25",X"2F",X"37",X"38",
		X"2A",X"2A",X"2B",X"29",X"18",X"19",X"18",X"37",X"38",X"18",X"10",X"00",X"18",X"1A",X"18",X"19",
		X"37",X"38",X"29",X"04",X"02",X"03",X"18",X"37",X"38",X"18",X"1A",X"32",X"18",X"1A",X"37",X"38",
		X"33",X"28",X"28",X"36",X"28",X"28",X"35",X"37",X"38",X"32",X"28",X"28",X"34",X"28",X"0A",X"37",
		X"38",X"11",X"28",X"28",X"36",X"28",X"16",X"37",X"38",X"15",X"28",X"28",X"28",X"00",X"37",X"38",
		X"0C",X"1B",X"1B",X"1C",X"1B",X"1B",X"0D",X"37",X"38",X"0C",X"1B",X"1D",X"1B",X"0D",X"37",X"38",
		X"0C",X"1B",X"1C",X"1C",X"1E",X"1B",X"0D",X"37",X"38",X"0C",X"1B",X"1C",X"1E",X"1C",X"37",X"38",
		X"1C",X"1F",X"20",X"1F",X"30",X"31",X"37",X"38",X"20",X"1F",X"1C",X"1F",X"1F",X"36",X"37",X"38",
		X"1F",X"1F",X"34",X"1F",X"17",X"1F",X"37",X"38",X"2B",X"2C",X"1A",X"1F",X"30",X"31",X"37",X"38",
		X"22",X"21",X"21",X"34",X"21",X"21",X"21",X"22",X"21",X"22",X"36",X"21",X"22",X"34",X"37",X"38",
		X"1E",X"1A",X"0C",X"0D",X"13",X"14",X"15",X"16",X"18",X"1A",X"1C",X"1C",X"1C",X"1B",X"37",X"38",
		X"33",X"36",X"33",X"33",X"36",X"35",X"34",X"33",X"35",X"33",X"33",X"34",X"36",X"33",X"37",X"38",
		X"33",X"35",X"36",X"33",X"33",X"34",X"33",X"33",X"33",X"05",X"36",X"33",X"35",X"33",X"37",X"38",
		X"05",X"14",X"0F",X"04",X"02",X"03",X"12",X"06",X"07",X"37",X"38",X"00",X"11",X"02",X"03",X"00",
		X"04",X"37",X"38",X"0A",X"0F",X"02",X"03",X"06",X"07",X"37",X"38",X"08",X"09",X"08",X"37",X"38",
		X"34",X"24",X"24",X"26",X"24",X"24",X"26",X"24",X"37",X"38",X"24",X"14",X"24",X"24",X"2F",X"24",
		X"37",X"38",X"00",X"00",X"24",X"24",X"26",X"24",X"37",X"38",X"25",X"26",X"25",X"2F",X"37",X"38",
		X"2A",X"2A",X"2B",X"29",X"18",X"19",X"18",X"37",X"38",X"18",X"10",X"00",X"18",X"1A",X"18",X"19",
		X"37",X"38",X"29",X"04",X"02",X"03",X"18",X"37",X"38",X"18",X"1A",X"32",X"18",X"1A",X"37",X"38",
		X"33",X"28",X"28",X"36",X"28",X"28",X"35",X"37",X"38",X"32",X"28",X"28",X"34",X"28",X"0A",X"37",
		X"38",X"11",X"28",X"28",X"36",X"28",X"16",X"37",X"38",X"15",X"28",X"28",X"28",X"00",X"37",X"38",
		X"0C",X"1B",X"1B",X"1C",X"1B",X"1B",X"0D",X"37",X"38",X"0C",X"1B",X"1D",X"1B",X"0D",X"37",X"38",
		X"0C",X"1B",X"1C",X"1C",X"1E",X"1B",X"0D",X"37",X"38",X"0C",X"1B",X"1C",X"1E",X"1C",X"37",X"38",
		X"1C",X"1F",X"20",X"1F",X"30",X"31",X"37",X"38",X"20",X"1F",X"1C",X"1F",X"1F",X"36",X"37",X"38",
		X"1F",X"1F",X"34",X"1F",X"17",X"1F",X"37",X"38",X"2B",X"2C",X"1A",X"1F",X"30",X"31",X"37",X"38",
		X"22",X"21",X"21",X"34",X"21",X"21",X"21",X"22",X"21",X"22",X"36",X"21",X"22",X"34",X"37",X"38",
		X"1E",X"1A",X"0C",X"0D",X"13",X"14",X"15",X"16",X"18",X"1A",X"1C",X"1C",X"1C",X"1B",X"37",X"38",
		X"33",X"36",X"33",X"33",X"36",X"35",X"34",X"33",X"35",X"33",X"33",X"34",X"36",X"33",X"37",X"38",
		X"33",X"35",X"36",X"33",X"33",X"34",X"33",X"33",X"33",X"05",X"36",X"33",X"35",X"33",X"37",X"38",
		X"3D",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"3E",X"7D",X"54",X"55",X"1B",X"60",X"61",X"62",X"7E",
		X"7D",X"56",X"57",X"1F",X"63",X"7A",X"64",X"7E",X"7D",X"1C",X"3A",X"1C",X"65",X"66",X"67",X"7E",
		X"7D",X"1C",X"1C",X"54",X"55",X"7A",X"20",X"3A",X"7D",X"20",X"24",X"56",X"57",X"7A",X"1C",X"7E",
		X"7D",X"23",X"1B",X"1B",X"1B",X"1B",X"3A",X"7E",X"3F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"40",
		X"3D",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"3E",X"7D",X"1D",X"1B",X"1B",X"1B",X"1B",X"1B",X"3A",
		X"7D",X"41",X"42",X"7A",X"7A",X"7A",X"7A",X"7E",X"3A",X"43",X"44",X"7A",X"1D",X"1B",X"1B",X"3A",
		X"7D",X"1C",X"36",X"59",X"31",X"59",X"5A",X"7E",X"7D",X"23",X"31",X"7A",X"4F",X"7A",X"5C",X"7E",
		X"7D",X"7A",X"5D",X"5E",X"34",X"5E",X"5F",X"7E",X"3F",X"7F",X"7F",X"7F",X"3A",X"7F",X"7F",X"40",
		X"3D",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"3E",X"3A",X"1B",X"1B",X"1B",X"3D",X"7C",X"7C",X"7C",
		X"7D",X"60",X"61",X"62",X"7D",X"00",X"01",X"02",X"3A",X"63",X"57",X"64",X"7D",X"03",X"03",X"00",
		X"7D",X"65",X"66",X"67",X"3F",X"7F",X"7F",X"7F",X"7D",X"1C",X"7A",X"7A",X"54",X"55",X"1C",X"7E",
		X"7D",X"23",X"1B",X"1B",X"56",X"57",X"25",X"7E",X"3F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"40",
		X"3D",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"3E",X"3E",X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",X"3A",
		X"7A",X"7C",X"7C",X"7C",X"7C",X"7C",X"42",X"7E",X"1B",X"1B",X"1E",X"1F",X"54",X"55",X"7E",X"7E",
		X"7F",X"7A",X"1C",X"1C",X"56",X"57",X"7E",X"7E",X"7D",X"7D",X"1C",X"23",X"1B",X"25",X"7E",X"3A",
		X"7D",X"3F",X"3A",X"7F",X"7F",X"7F",X"44",X"7E",X"3F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"40",
		X"3D",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"3E",X"7D",X"3D",X"7C",X"7C",X"7C",X"3E",X"1D",X"3A",
		X"7D",X"7D",X"26",X"27",X"28",X"7E",X"1C",X"7E",X"7D",X"7D",X"2B",X"2C",X"2D",X"7E",X"1C",X"7E",
		X"7D",X"3F",X"7F",X"7F",X"7F",X"40",X"25",X"7E",X"3A",X"1B",X"1B",X"1B",X"1B",X"54",X"55",X"7E",
		X"7D",X"1D",X"1B",X"1B",X"1B",X"56",X"57",X"7E",X"3F",X"3A",X"7F",X"7F",X"7F",X"7F",X"7F",X"40",
		X"3D",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"3E",X"3A",X"1B",X"1F",X"7A",X"54",X"55",X"1D",X"3A",
		X"7D",X"06",X"07",X"08",X"56",X"57",X"1C",X"7E",X"7D",X"0B",X"0C",X"0D",X"23",X"1B",X"25",X"7E",
		X"7D",X"0E",X"0F",X"0F",X"0F",X"0F",X"10",X"7E",X"7D",X"11",X"4F",X"7A",X"7A",X"4F",X"12",X"3A",
		X"7D",X"13",X"14",X"14",X"14",X"14",X"15",X"7E",X"3F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"40",
		X"3D",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"3E",X"3A",X"06",X"07",X"07",X"07",X"08",X"7A",X"7E",
		X"7D",X"09",X"7A",X"7A",X"7A",X"4C",X"4D",X"4D",X"7D",X"0B",X"0C",X"0C",X"0C",X"0D",X"1C",X"7E",
		X"7D",X"20",X"1B",X"1B",X"54",X"55",X"1C",X"06",X"3A",X"26",X"27",X"28",X"56",X"57",X"20",X"09",
		X"7D",X"2B",X"2C",X"2D",X"24",X"1B",X"25",X"09",X"3F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"09",
		X"3D",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"3E",X"7D",X"06",X"07",X"08",X"1D",X"1B",X"1B",X"3A",
		X"4D",X"4E",X"7A",X"0A",X"1C",X"50",X"51",X"7E",X"7D",X"0B",X"0C",X"0D",X"24",X"52",X"53",X"7E",
		X"07",X"07",X"08",X"24",X"1B",X"1B",X"1E",X"3A",X"4F",X"4F",X"0A",X"7A",X"54",X"55",X"1C",X"7E",
		X"4F",X"4F",X"0A",X"7A",X"56",X"57",X"25",X"7E",X"4F",X"4F",X"0A",X"7F",X"7F",X"7F",X"7F",X"40",
		X"3D",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"3E",X"7D",X"1D",X"1B",X"1B",X"1B",X"1B",X"1E",X"3A",
		X"7D",X"23",X"54",X"55",X"58",X"59",X"37",X"7E",X"7D",X"7A",X"56",X"57",X"5B",X"7A",X"5C",X"7E",
		X"3A",X"1B",X"1B",X"22",X"5B",X"7A",X"5C",X"7E",X"7D",X"7A",X"54",X"55",X"5B",X"7A",X"5C",X"7E",
		X"7D",X"7A",X"56",X"57",X"5D",X"5E",X"5F",X"3A",X"3F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"40",
		X"3D",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"3E",X"3A",X"1E",X"1B",X"41",X"45",X"42",X"7A",X"7E",
		X"7D",X"1C",X"7A",X"43",X"48",X"44",X"7A",X"7E",X"7D",X"20",X"54",X"55",X"7A",X"1C",X"7A",X"7E",
		X"7D",X"1C",X"56",X"57",X"1B",X"24",X"1B",X"3A",X"7D",X"1C",X"7A",X"7A",X"7A",X"7A",X"7A",X"7E",
		X"3A",X"24",X"1B",X"1B",X"1F",X"7A",X"7A",X"7E",X"3F",X"7F",X"7F",X"7F",X"3A",X"7F",X"7F",X"40",
		X"3D",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"3E",X"7D",X"41",X"42",X"7A",X"41",X"45",X"42",X"7E",
		X"7D",X"43",X"44",X"1F",X"46",X"88",X"47",X"7E",X"7D",X"1C",X"3A",X"1C",X"43",X"48",X"44",X"7E",
		X"7D",X"1C",X"1C",X"54",X"55",X"7A",X"20",X"3A",X"7D",X"20",X"3A",X"56",X"57",X"7A",X"1C",X"7E",
		X"7D",X"23",X"1B",X"1B",X"1B",X"1B",X"3A",X"7E",X"3F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"40",
		X"3D",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"3E",X"7D",X"1D",X"1B",X"54",X"89",X"89",X"1B",X"3A",
		X"7D",X"41",X"42",X"8C",X"88",X"8A",X"7A",X"7E",X"3A",X"43",X"44",X"56",X"8B",X"57",X"1B",X"3A",
		X"7D",X"1C",X"36",X"59",X"31",X"59",X"5A",X"7E",X"7D",X"23",X"31",X"7A",X"7A",X"7A",X"5C",X"7E",
		X"7D",X"7A",X"5D",X"5E",X"34",X"5E",X"5F",X"7E",X"3F",X"7F",X"7F",X"7F",X"3A",X"7F",X"7F",X"40",
		X"3D",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"3E",X"3A",X"1E",X"1E",X"1E",X"1E",X"1E",X"1E",X"3A",
		X"7D",X"20",X"21",X"21",X"21",X"21",X"21",X"3A",X"3A",X"21",X"21",X"21",X"21",X"21",X"21",X"3A",
		X"7D",X"20",X"21",X"21",X"21",X"21",X"21",X"3A",X"7D",X"20",X"21",X"21",X"21",X"21",X"21",X"3A",
		X"7D",X"23",X"24",X"24",X"24",X"24",X"24",X"3A",X"3F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"40",
		X"3D",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"3E",X"3A",X"1E",X"1E",X"1E",X"1E",X"1E",X"1E",X"3A",
		X"3A",X"21",X"21",X"21",X"21",X"21",X"22",X"7E",X"3A",X"21",X"21",X"21",X"21",X"21",X"22",X"7E",
		X"3A",X"21",X"21",X"21",X"21",X"21",X"22",X"7E",X"3A",X"21",X"21",X"21",X"21",X"21",X"21",X"3A",
		X"3A",X"24",X"24",X"24",X"24",X"24",X"25",X"7E",X"3F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"40",
		X"3D",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"3E",X"7D",X"3D",X"7C",X"7C",X"7C",X"3E",X"1D",X"3A",
		X"7D",X"7D",X"50",X"89",X"51",X"7E",X"1C",X"7E",X"7D",X"7D",X"52",X"8B",X"53",X"7E",X"1C",X"7E",
		X"7D",X"3F",X"7F",X"7F",X"7A",X"7E",X"22",X"7E",X"3A",X"1B",X"1E",X"1B",X"7D",X"7E",X"1C",X"7E",
		X"7D",X"1D",X"24",X"1B",X"3F",X"40",X"25",X"7E",X"3F",X"3A",X"7F",X"7F",X"7F",X"7F",X"7F",X"40",
		X"3D",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"3E",X"3A",X"00",X"01",X"01",X"01",X"02",X"1D",X"3A",
		X"7D",X"03",X"03",X"03",X"03",X"00",X"1C",X"7E",X"7D",X"7A",X"1D",X"1B",X"24",X"1B",X"25",X"7E",
		X"7D",X"0E",X"0F",X"0F",X"0F",X"0F",X"10",X"7E",X"7D",X"11",X"7A",X"7A",X"7A",X"7A",X"12",X"3A",
		X"7D",X"13",X"14",X"14",X"14",X"14",X"15",X"7E",X"3F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"40",
		X"3D",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"3E",X"3A",X"00",X"00",X"08",X"3A",X"3A",X"3A",X"3A",
		X"7D",X"09",X"7A",X"0A",X"3A",X"3A",X"3A",X"3A",X"7D",X"0B",X"0C",X"0D",X"7A",X"7A",X"1C",X"7E",
		X"7D",X"20",X"1B",X"1B",X"54",X"55",X"1C",X"7E",X"3A",X"1E",X"1E",X"1E",X"8C",X"8A",X"20",X"3A",
		X"7D",X"23",X"24",X"25",X"56",X"57",X"25",X"7E",X"3F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"40",
		X"3D",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"3E",X"7D",X"4F",X"1B",X"1B",X"1B",X"3A",X"1E",X"3A",
		X"7D",X"7A",X"7A",X"7A",X"7A",X"7A",X"1C",X"7E",X"7D",X"7A",X"7A",X"3A",X"1B",X"1B",X"25",X"7E",
		X"7D",X"7A",X"3A",X"24",X"1B",X"1B",X"1E",X"3A",X"7D",X"7A",X"7A",X"50",X"51",X"7A",X"1C",X"7E",
		X"7D",X"7A",X"7A",X"52",X"53",X"1B",X"25",X"7E",X"3F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"40",
		X"3D",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"3E",X"3A",X"1B",X"1B",X"1E",X"1B",X"3A",X"3A",X"7E",
		X"7D",X"7A",X"54",X"55",X"58",X"59",X"37",X"7E",X"7D",X"7A",X"56",X"57",X"5B",X"88",X"5C",X"7E",
		X"3A",X"1B",X"1B",X"22",X"5B",X"88",X"5C",X"7E",X"7D",X"7A",X"54",X"55",X"5B",X"88",X"5C",X"7E",
		X"7D",X"7A",X"56",X"57",X"5D",X"5E",X"5F",X"3A",X"3F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"40",
		X"3D",X"7C",X"7C",X"7C",X"06",X"07",X"07",X"08",X"3A",X"1F",X"7A",X"7A",X"09",X"7A",X"7A",X"0A",
		X"7D",X"1C",X"7A",X"7A",X"0B",X"0C",X"0C",X"0D",X"7D",X"20",X"54",X"55",X"7A",X"1C",X"7A",X"7E",
		X"7D",X"1C",X"56",X"57",X"1B",X"24",X"1B",X"3A",X"7D",X"1C",X"7A",X"7A",X"7A",X"7A",X"7A",X"7E",
		X"3A",X"24",X"1B",X"1B",X"1F",X"7A",X"7A",X"7E",X"3F",X"7F",X"7F",X"7F",X"3A",X"7F",X"7F",X"40",
		X"60",X"61",X"61",X"61",X"61",X"61",X"61",X"62",X"63",X"50",X"51",X"7A",X"7A",X"7A",X"7A",X"64",
		X"63",X"52",X"53",X"1F",X"1D",X"3A",X"7A",X"64",X"63",X"7A",X"7A",X"36",X"37",X"7A",X"7A",X"64",
		X"63",X"7A",X"7A",X"38",X"39",X"7A",X"7A",X"64",X"63",X"3A",X"1B",X"22",X"23",X"50",X"51",X"64",
		X"63",X"7A",X"7A",X"23",X"1B",X"52",X"53",X"64",X"65",X"66",X"66",X"66",X"66",X"66",X"66",X"67",
		X"41",X"45",X"82",X"61",X"61",X"61",X"80",X"45",X"3A",X"1B",X"31",X"3A",X"3A",X"3A",X"5C",X"21",
		X"46",X"7A",X"5B",X"3A",X"70",X"3A",X"5C",X"21",X"46",X"7A",X"5B",X"3A",X"76",X"3A",X"16",X"4D",
		X"46",X"7A",X"5B",X"3A",X"77",X"3A",X"5C",X"21",X"3A",X"1B",X"31",X"3A",X"3A",X"3A",X"5C",X"21",
		X"46",X"7A",X"5D",X"5E",X"5E",X"5E",X"5F",X"21",X"43",X"48",X"48",X"48",X"48",X"21",X"21",X"21",
		X"21",X"21",X"21",X"21",X"45",X"45",X"45",X"42",X"21",X"58",X"59",X"59",X"59",X"5A",X"7A",X"47",
		X"21",X"5B",X"0E",X"0F",X"10",X"5C",X"7A",X"47",X"4D",X"17",X"13",X"14",X"15",X"5C",X"1D",X"3A",
		X"21",X"5D",X"5E",X"5E",X"5E",X"5F",X"1C",X"47",X"21",X"21",X"21",X"21",X"21",X"7A",X"1C",X"47",
		X"21",X"20",X"7A",X"1D",X"1B",X"1B",X"25",X"47",X"21",X"48",X"48",X"48",X"48",X"48",X"48",X"44",
		X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"04",X"03",X"3A",
		X"3A",X"3A",X"3A",X"3A",X"3A",X"05",X"04",X"3A",X"3A",X"3A",X"3A",X"04",X"03",X"3A",X"3A",X"3A",
		X"3A",X"3A",X"3A",X"05",X"04",X"3A",X"3A",X"3A",X"3A",X"04",X"03",X"3A",X"3A",X"3A",X"3A",X"3A",
		X"3A",X"05",X"04",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",
		X"41",X"42",X"41",X"42",X"41",X"42",X"41",X"42",X"43",X"44",X"43",X"44",X"43",X"44",X"43",X"44",
		X"41",X"42",X"41",X"42",X"41",X"42",X"41",X"42",X"43",X"44",X"43",X"44",X"43",X"44",X"43",X"44",
		X"41",X"42",X"41",X"42",X"41",X"42",X"41",X"42",X"43",X"44",X"43",X"44",X"43",X"44",X"43",X"44",
		X"41",X"42",X"41",X"42",X"41",X"42",X"41",X"42",X"43",X"44",X"43",X"44",X"43",X"44",X"43",X"44",
		X"41",X"42",X"41",X"42",X"41",X"42",X"41",X"42",X"43",X"44",X"43",X"44",X"43",X"44",X"43",X"44",
		X"41",X"42",X"41",X"42",X"50",X"51",X"41",X"42",X"43",X"44",X"43",X"44",X"52",X"53",X"43",X"44",
		X"41",X"42",X"41",X"42",X"41",X"42",X"41",X"42",X"43",X"44",X"43",X"44",X"43",X"44",X"43",X"44",
		X"41",X"42",X"50",X"51",X"41",X"42",X"41",X"42",X"43",X"44",X"52",X"53",X"43",X"44",X"43",X"44",
		X"41",X"42",X"3A",X"3A",X"41",X"42",X"41",X"42",X"43",X"44",X"3A",X"3A",X"43",X"44",X"43",X"44",
		X"41",X"42",X"41",X"42",X"41",X"42",X"41",X"42",X"43",X"44",X"43",X"44",X"43",X"44",X"43",X"44",
		X"41",X"42",X"41",X"42",X"3A",X"3A",X"41",X"42",X"43",X"44",X"43",X"44",X"3A",X"3A",X"43",X"44",
		X"3A",X"3A",X"41",X"42",X"41",X"42",X"41",X"42",X"3A",X"3A",X"43",X"44",X"43",X"44",X"43",X"44",
		X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",
		X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",
		X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",
		X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",
		X"54",X"55",X"54",X"55",X"54",X"55",X"3A",X"3A",X"56",X"57",X"56",X"57",X"56",X"57",X"3A",X"3A",
		X"3A",X"3A",X"54",X"55",X"54",X"55",X"54",X"55",X"3A",X"3A",X"56",X"57",X"56",X"57",X"56",X"57",
		X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",
		X"54",X"55",X"54",X"55",X"3A",X"3A",X"54",X"55",X"56",X"57",X"56",X"57",X"3A",X"3A",X"56",X"57",
		X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",
		X"54",X"55",X"00",X"02",X"54",X"55",X"54",X"55",X"56",X"57",X"03",X"00",X"56",X"57",X"56",X"57",
		X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",
		X"54",X"55",X"54",X"55",X"00",X"02",X"54",X"55",X"56",X"57",X"56",X"57",X"03",X"00",X"56",X"57",
		X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",
		X"54",X"55",X"1E",X"1B",X"54",X"55",X"54",X"55",X"56",X"57",X"23",X"1F",X"56",X"57",X"56",X"57",
		X"54",X"55",X"7A",X"20",X"1E",X"1B",X"54",X"55",X"56",X"57",X"1D",X"25",X"3A",X"7A",X"56",X"57",
		X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"56",X"57",X"56",X"57",X"56",X"57",X"56",X"57",
		X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",
		X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",
		X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",
		X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",
		X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"1D",X"1F",X"3A",X"3A",X"3A",X"3A",X"3A",
		X"3A",X"23",X"7A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"1D",X"1F",X"3A",X"3A",X"3A",
		X"3A",X"3A",X"3A",X"23",X"25",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"7A",X"1F",X"3A",
		X"3A",X"3A",X"3A",X"3A",X"3A",X"23",X"25",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",
		X"60",X"62",X"03",X"03",X"60",X"62",X"03",X"03",X"65",X"67",X"60",X"62",X"65",X"67",X"60",X"62",
		X"60",X"62",X"65",X"67",X"60",X"62",X"65",X"67",X"65",X"67",X"60",X"62",X"65",X"67",X"60",X"62",
		X"60",X"62",X"65",X"67",X"60",X"62",X"65",X"67",X"65",X"67",X"60",X"62",X"65",X"67",X"60",X"62",
		X"60",X"62",X"65",X"67",X"60",X"62",X"65",X"67",X"65",X"67",X"60",X"62",X"65",X"67",X"60",X"62",
		X"60",X"62",X"60",X"62",X"60",X"62",X"60",X"62",X"65",X"67",X"65",X"67",X"65",X"67",X"65",X"67",
		X"60",X"62",X"1D",X"1F",X"1D",X"1F",X"60",X"62",X"65",X"67",X"23",X"1D",X"1F",X"25",X"65",X"67",
		X"60",X"62",X"1D",X"23",X"25",X"1F",X"60",X"62",X"65",X"67",X"23",X"25",X"23",X"25",X"65",X"67",
		X"60",X"62",X"60",X"62",X"60",X"62",X"60",X"62",X"65",X"67",X"65",X"67",X"65",X"67",X"65",X"67",
		X"1D",X"1F",X"1D",X"1F",X"1D",X"1F",X"3D",X"3E",X"23",X"25",X"23",X"25",X"23",X"25",X"3F",X"40",
		X"1D",X"1F",X"3D",X"3E",X"1D",X"1F",X"1D",X"1F",X"23",X"25",X"3F",X"40",X"23",X"25",X"23",X"25",
		X"1D",X"1F",X"1D",X"1F",X"1D",X"1F",X"1D",X"1F",X"23",X"25",X"23",X"25",X"23",X"25",X"23",X"25",
		X"1D",X"1F",X"1D",X"1F",X"3D",X"3E",X"1D",X"1F",X"23",X"25",X"23",X"25",X"3F",X"40",X"23",X"25",
		X"3D",X"3E",X"3D",X"3E",X"3D",X"3E",X"3D",X"3E",X"3F",X"40",X"3F",X"40",X"3F",X"40",X"3F",X"40",
		X"3D",X"3E",X"3D",X"3E",X"3D",X"3E",X"3D",X"3E",X"3F",X"40",X"3F",X"40",X"3F",X"40",X"3F",X"40",
		X"3D",X"3E",X"3D",X"3E",X"3D",X"3E",X"3D",X"3E",X"3F",X"40",X"3F",X"40",X"3F",X"40",X"3F",X"40",
		X"3D",X"3E",X"3D",X"3E",X"3D",X"3E",X"3D",X"3E",X"3F",X"40",X"3F",X"40",X"3F",X"40",X"3F",X"40",
		X"3D",X"3E",X"3D",X"3E",X"3D",X"3E",X"3D",X"3E",X"3D",X"3E",X"3F",X"40",X"3D",X"3E",X"3F",X"40",
		X"3F",X"40",X"3D",X"3E",X"3F",X"40",X"3D",X"3E",X"3D",X"3E",X"3F",X"40",X"3D",X"3E",X"3F",X"40",
		X"3F",X"40",X"3D",X"3E",X"3F",X"40",X"3D",X"3E",X"3D",X"3E",X"3F",X"40",X"3D",X"3E",X"3F",X"40",
		X"3F",X"40",X"3D",X"3E",X"3F",X"40",X"3D",X"3E",X"3D",X"3E",X"3F",X"40",X"3D",X"3E",X"3F",X"40",
		X"3D",X"3E",X"3D",X"3E",X"3D",X"3E",X"3D",X"3E",X"3D",X"3E",X"3F",X"40",X"3D",X"3E",X"3F",X"40",
		X"3F",X"40",X"50",X"51",X"3F",X"40",X"3D",X"3E",X"3D",X"3E",X"52",X"53",X"3D",X"3E",X"3F",X"40",
		X"3F",X"40",X"3D",X"3E",X"3F",X"40",X"3D",X"3E",X"3D",X"3E",X"3F",X"40",X"3D",X"3E",X"3F",X"40",
		X"3F",X"40",X"3D",X"3E",X"3F",X"40",X"50",X"51",X"3D",X"3E",X"3F",X"40",X"3D",X"3E",X"52",X"53",
		X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",
		X"00",X"02",X"4F",X"4F",X"00",X"02",X"00",X"02",X"03",X"00",X"4F",X"4F",X"03",X"00",X"03",X"00",
		X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",
		X"00",X"02",X"00",X"02",X"4F",X"4F",X"00",X"02",X"03",X"00",X"03",X"00",X"4F",X"4F",X"03",X"00",
		X"2E",X"30",X"2E",X"30",X"2E",X"30",X"2E",X"30",X"33",X"35",X"33",X"35",X"33",X"35",X"33",X"35",
		X"30",X"2E",X"30",X"2E",X"30",X"2E",X"30",X"2E",X"35",X"33",X"35",X"33",X"35",X"33",X"35",X"33",
		X"2E",X"30",X"2E",X"30",X"2E",X"30",X"2E",X"30",X"33",X"35",X"33",X"35",X"33",X"35",X"33",X"35",
		X"30",X"2E",X"30",X"2E",X"30",X"2E",X"30",X"2E",X"35",X"33",X"35",X"33",X"35",X"33",X"35",X"33",
		X"41",X"42",X"41",X"42",X"41",X"42",X"41",X"42",X"43",X"44",X"46",X"47",X"43",X"44",X"46",X"47",
		X"41",X"42",X"43",X"44",X"41",X"42",X"43",X"44",X"43",X"44",X"41",X"42",X"43",X"44",X"41",X"42",
		X"41",X"42",X"43",X"44",X"41",X"42",X"43",X"44",X"43",X"44",X"41",X"42",X"43",X"44",X"41",X"42",
		X"41",X"42",X"43",X"44",X"41",X"42",X"43",X"44",X"43",X"44",X"41",X"42",X"43",X"44",X"41",X"42",
		X"41",X"42",X"41",X"42",X"41",X"42",X"41",X"42",X"46",X"47",X"43",X"44",X"46",X"47",X"43",X"44",
		X"43",X"44",X"41",X"42",X"43",X"44",X"41",X"42",X"41",X"42",X"46",X"47",X"41",X"42",X"46",X"47",
		X"46",X"47",X"43",X"44",X"46",X"47",X"43",X"44",X"43",X"44",X"41",X"42",X"43",X"44",X"41",X"42",
		X"41",X"42",X"46",X"47",X"41",X"42",X"46",X"47",X"46",X"47",X"43",X"44",X"46",X"47",X"43",X"44",
		X"41",X"42",X"41",X"42",X"41",X"42",X"41",X"42",X"43",X"44",X"46",X"47",X"43",X"44",X"46",X"47",
		X"41",X"42",X"43",X"44",X"50",X"51",X"43",X"44",X"43",X"44",X"41",X"42",X"52",X"53",X"41",X"42",
		X"50",X"51",X"43",X"44",X"41",X"42",X"43",X"44",X"52",X"53",X"41",X"42",X"43",X"44",X"41",X"42",
		X"41",X"42",X"43",X"44",X"41",X"42",X"43",X"44",X"43",X"44",X"41",X"42",X"43",X"44",X"50",X"51",
		X"41",X"42",X"41",X"42",X"41",X"42",X"41",X"42",X"46",X"47",X"43",X"44",X"46",X"47",X"43",X"44",
		X"43",X"44",X"41",X"42",X"43",X"44",X"41",X"42",X"41",X"42",X"46",X"47",X"54",X"55",X"46",X"47",
		X"46",X"47",X"43",X"44",X"46",X"47",X"43",X"44",X"43",X"44",X"41",X"42",X"56",X"57",X"41",X"42",
		X"54",X"55",X"46",X"47",X"41",X"42",X"46",X"47",X"46",X"47",X"43",X"44",X"46",X"47",X"43",X"44",
		X"3D",X"3E",X"3D",X"3E",X"3D",X"3E",X"3D",X"3E",X"7D",X"7E",X"3D",X"3E",X"7D",X"7E",X"7D",X"7E",
		X"3F",X"40",X"7D",X"7E",X"3D",X"3E",X"3F",X"40",X"3D",X"3E",X"3F",X"40",X"7D",X"7E",X"3D",X"3E",
		X"7D",X"7E",X"3D",X"3E",X"3F",X"40",X"7D",X"7E",X"3F",X"40",X"7D",X"7E",X"3D",X"3E",X"3F",X"40",
		X"3D",X"3E",X"3F",X"40",X"7D",X"7E",X"3D",X"3E",X"7D",X"7E",X"3D",X"3E",X"3F",X"40",X"7D",X"7E",
		X"3D",X"3E",X"3D",X"3E",X"3D",X"3E",X"3D",X"3E",X"54",X"55",X"7D",X"7E",X"7D",X"7E",X"3D",X"3E",
		X"7D",X"7E",X"3D",X"3E",X"3F",X"40",X"7D",X"7E",X"56",X"57",X"7D",X"7E",X"3D",X"3E",X"3F",X"40",
		X"3D",X"3E",X"3F",X"40",X"7D",X"7E",X"3D",X"3E",X"7D",X"7E",X"3D",X"3E",X"3F",X"40",X"7D",X"7E",
		X"3F",X"40",X"7D",X"7E",X"54",X"55",X"3F",X"40",X"3D",X"3E",X"3F",X"40",X"7D",X"7E",X"3D",X"3E",
		X"3D",X"3E",X"3D",X"3E",X"3D",X"3E",X"3D",X"3E",X"7D",X"7E",X"7D",X"7E",X"3D",X"3E",X"3F",X"40",
		X"3D",X"3E",X"3F",X"40",X"7D",X"7E",X"3D",X"3E",X"7D",X"7E",X"54",X"55",X"3F",X"40",X"7D",X"7E",
		X"3F",X"40",X"7D",X"7E",X"3D",X"3E",X"3F",X"40",X"3D",X"3E",X"56",X"57",X"7D",X"7E",X"3D",X"3E",
		X"7D",X"7E",X"3D",X"3E",X"3F",X"40",X"7D",X"7E",X"3F",X"40",X"7D",X"7E",X"3D",X"3E",X"3F",X"40",
		X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"1D",X"1B",X"60",X"61",X"62",X"3A",X"3A",
		X"3A",X"70",X"3A",X"63",X"7A",X"64",X"3A",X"41",X"3A",X"76",X"3A",X"65",X"66",X"67",X"3A",X"43",
		X"3A",X"76",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"77",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",
		X"3A",X"23",X"1B",X"1B",X"1B",X"1B",X"1F",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"1C",X"3A",
		X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",
		X"42",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"44",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",
		X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"41",X"42",X"3A",X"3A",
		X"3A",X"3A",X"3A",X"3A",X"43",X"44",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",
		X"26",X"27",X"27",X"27",X"27",X"27",X"27",X"28",X"29",X"41",X"42",X"41",X"42",X"41",X"42",X"2A",
		X"29",X"43",X"44",X"43",X"44",X"43",X"44",X"2A",X"29",X"41",X"42",X"54",X"55",X"41",X"42",X"2A",
		X"29",X"43",X"44",X"56",X"57",X"43",X"44",X"2A",X"29",X"41",X"42",X"41",X"42",X"41",X"42",X"2A",
		X"29",X"43",X"44",X"43",X"44",X"43",X"44",X"2A",X"2B",X"2C",X"2C",X"2C",X"2C",X"2C",X"2C",X"2D",
		X"26",X"27",X"27",X"27",X"27",X"27",X"27",X"28",X"29",X"3D",X"3E",X"3D",X"3E",X"3D",X"3E",X"2A",
		X"29",X"3F",X"40",X"3F",X"40",X"3F",X"40",X"2A",X"29",X"3D",X"3E",X"3D",X"3E",X"3D",X"3E",X"2A",
		X"29",X"3F",X"40",X"3F",X"40",X"3F",X"40",X"2A",X"29",X"3D",X"3E",X"3D",X"3E",X"3D",X"3E",X"2A",
		X"29",X"3F",X"40",X"3F",X"40",X"3F",X"40",X"2A",X"2B",X"2C",X"2C",X"2C",X"2C",X"2C",X"2C",X"2D",
		X"26",X"27",X"27",X"27",X"27",X"27",X"27",X"28",X"29",X"3D",X"3E",X"3D",X"3E",X"3D",X"3E",X"2A",
		X"29",X"3F",X"40",X"3F",X"40",X"3F",X"40",X"2A",X"29",X"3D",X"3E",X"54",X"55",X"3D",X"3E",X"2A",
		X"29",X"3F",X"40",X"56",X"57",X"3F",X"40",X"2A",X"29",X"3D",X"3E",X"3D",X"3E",X"54",X"55",X"2A",
		X"29",X"3F",X"40",X"3F",X"40",X"56",X"57",X"2A",X"2B",X"2C",X"2C",X"2C",X"2C",X"2C",X"2C",X"2D",
		X"26",X"27",X"27",X"27",X"27",X"27",X"27",X"28",X"29",X"3D",X"3E",X"3D",X"3E",X"54",X"55",X"2A",
		X"29",X"3F",X"40",X"3F",X"40",X"56",X"57",X"2A",X"29",X"3D",X"3E",X"7A",X"7A",X"3F",X"40",X"2A",
		X"29",X"3F",X"40",X"7A",X"7A",X"3D",X"3E",X"2A",X"29",X"7A",X"7A",X"3D",X"3E",X"54",X"55",X"2A",
		X"29",X"7A",X"7A",X"3F",X"40",X"56",X"57",X"2A",X"2B",X"2C",X"2C",X"2C",X"2C",X"2C",X"2C",X"2D",
		X"26",X"27",X"27",X"27",X"27",X"27",X"27",X"28",X"29",X"3D",X"3E",X"7A",X"7A",X"3D",X"3E",X"2A",
		X"29",X"3F",X"40",X"7A",X"7A",X"3F",X"40",X"2A",X"29",X"7A",X"7A",X"54",X"55",X"3D",X"3E",X"2A",
		X"29",X"7A",X"7A",X"56",X"57",X"3F",X"40",X"2A",X"29",X"3D",X"3E",X"3D",X"3E",X"3D",X"3E",X"2A",
		X"29",X"3F",X"40",X"3F",X"40",X"3F",X"40",X"2A",X"2B",X"2C",X"2C",X"2C",X"2C",X"2C",X"2C",X"2D",
		X"3D",X"7C",X"7C",X"7C",X"3E",X"8E",X"03",X"03",X"7D",X"7A",X"7A",X"7A",X"7E",X"90",X"8E",X"03",
		X"7D",X"7A",X"7A",X"7A",X"7E",X"90",X"6B",X"6C",X"7D",X"7A",X"7A",X"7A",X"7E",X"71",X"72",X"72",
		X"7D",X"7A",X"7A",X"7A",X"6E",X"68",X"68",X"78",X"7D",X"7A",X"7A",X"74",X"79",X"79",X"79",X"79",
		X"7D",X"7A",X"74",X"79",X"79",X"79",X"79",X"79",X"7D",X"7A",X"4F",X"8F",X"4F",X"8F",X"4F",X"8F",
		X"03",X"03",X"8D",X"3D",X"7C",X"7C",X"7C",X"3E",X"03",X"8D",X"91",X"7D",X"7A",X"7A",X"7A",X"7E",
		X"6C",X"6D",X"91",X"7D",X"7A",X"7A",X"7A",X"7E",X"72",X"72",X"73",X"7D",X"7A",X"7A",X"7A",X"7E",
		X"68",X"78",X"78",X"6F",X"7A",X"7A",X"7A",X"7E",X"79",X"79",X"79",X"79",X"75",X"7A",X"7A",X"7E",
		X"79",X"79",X"79",X"79",X"79",X"75",X"7A",X"7E",X"4F",X"8F",X"4F",X"8F",X"4F",X"8F",X"7A",X"7E",
		X"21",X"1E",X"E6",X"35",X"7E",X"FE",X"FF",X"00",X"3E",X"01",X"77",X"CD",X"A1",X"5E",X"3A",X"00",
		X"D0",X"E6",X"08",X"28",X"46",X"3A",X"1C",X"E6",X"FE",X"00",X"C8",X"3E",X"00",X"32",X"1C",X"E6",
		X"21",X"19",X"E6",X"35",X"C0",X"3A",X"18",X"E6",X"6F",X"26",X"00",X"11",X"F4",X"5E",X"19",X"7E",
		X"32",X"19",X"E6",X"11",X"10",X"00",X"19",X"3A",X"07",X"E2",X"86",X"32",X"07",X"E2",X"C6",X"F6",
		X"30",X"05",X"3E",X"09",X"32",X"07",X"E2",X"3E",X"05",X"CD",X"34",X"5F",X"3A",X"F4",X"83",X"FE",
		X"43",X"C0",X"3A",X"07",X"E2",X"C6",X"30",X"32",X"FC",X"83",X"C9",X"3E",X"01",X"32",X"1C",X"E6",
		X"C9",X"3A",X"00",X"D0",X"E6",X"04",X"28",X"46",X"3A",X"1D",X"E6",X"FE",X"00",X"C8",X"3E",X"00",
		X"32",X"1D",X"E6",X"21",X"1B",X"E6",X"35",X"C0",X"3A",X"1A",X"E6",X"6F",X"26",X"00",X"11",X"14",
		X"5F",X"19",X"7E",X"32",X"1B",X"E6",X"11",X"10",X"00",X"19",X"3A",X"07",X"E2",X"86",X"32",X"07",
		X"E2",X"C6",X"F6",X"30",X"05",X"3E",X"09",X"32",X"07",X"E2",X"3E",X"05",X"CD",X"34",X"5F",X"3A",
		X"F4",X"83",X"FE",X"43",X"C0",X"3A",X"07",X"E2",X"C6",X"30",X"32",X"FC",X"83",X"C9",X"3E",X"01",
		X"32",X"1D",X"E6",X"C9",X"01",X"01",X"02",X"03",X"04",X"02",X"02",X"02",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"00",X"01",X"02",X"03",X"04",X"05",X"06",X"07",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"F5",X"3A",X"01",X"E2",X"FE",X"00",X"28",X"02",X"F1",X"C9",X"F1",X"F5",
		X"32",X"00",X"D0",X"F6",X"80",X"32",X"00",X"D0",X"F1",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"CD",X"26",X"40",X"CD",X"22",X"3E",X"CD",X"70",X"3E",X"21",X"19",X"60",X"CD",X"FB",X"3F",X"CD",
		X"07",X"43",X"CD",X"22",X"3E",X"CD",X"22",X"3E",X"C9",X"01",X"80",X"81",X"57",X"45",X"41",X"50",
		X"4F",X"4E",X"53",X"FE",X"06",X"FD",X"80",X"C7",X"32",X"20",X"50",X"4F",X"57",X"53",X"20",X"47",
		X"49",X"56",X"45",X"53",X"20",X"53",X"49",X"44",X"45",X"20",X"41",X"52",X"4D",X"53",X"FD",X"80",
		X"E2",X"50",X"4C",X"55",X"53",X"20",X"34",X"20",X"50",X"4F",X"57",X"53",X"20",X"47",X"49",X"56",
		X"45",X"53",X"20",X"53",X"4C",X"41",X"56",X"45",X"20",X"53",X"48",X"49",X"50",X"FD",X"81",X"02",
		X"50",X"4C",X"55",X"53",X"20",X"38",X"20",X"50",X"4F",X"57",X"53",X"20",X"47",X"49",X"56",X"45",
		X"53",X"20",X"57",X"41",X"56",X"45",X"20",X"47",X"55",X"4E",X"FE",X"01",X"FD",X"81",X"41",X"50",
		X"4F",X"57",X"45",X"52",X"20",X"4F",X"52",X"42",X"53",X"20",X"FE",X"16",X"1A",X"FE",X"06",X"FD",
		X"81",X"87",X"50",X"49",X"43",X"4B",X"20",X"55",X"50",X"20",X"31",X"30",X"20",X"49",X"4E",X"20",
		X"41",X"20",X"52",X"4F",X"57",X"20",X"41",X"4E",X"44",X"FD",X"81",X"A2",X"50",X"4C",X"41",X"43",
		X"45",X"20",X"4F",X"4E",X"20",X"44",X"52",X"4F",X"50",X"20",X"5A",X"4F",X"4E",X"45",X"20",X"46",
		X"4F",X"52",X"20",X"32",X"58",X"20",X"33",X"58",X"FD",X"81",X"C2",X"41",X"4E",X"44",X"20",X"34",
		X"58",X"20",X"42",X"4F",X"4E",X"55",X"53",X"20",X"4D",X"49",X"53",X"53",X"20",X"41",X"4E",X"59",
		X"20",X"42",X"45",X"46",X"4F",X"52",X"45",X"FD",X"81",X"E2",X"44",X"52",X"4F",X"50",X"20",X"5A",
		X"4F",X"4E",X"45",X"20",X"41",X"4E",X"44",X"20",X"4E",X"4F",X"20",X"42",X"4F",X"4E",X"55",X"53",
		X"FE",X"01",X"FD",X"82",X"21",X"53",X"48",X"49",X"45",X"4C",X"44",X"53",X"20",X"FE",X"06",X"18",
		X"FE",X"06",X"FD",X"82",X"67",X"50",X"49",X"43",X"4B",X"20",X"55",X"50",X"20",X"53",X"48",X"49",
		X"45",X"4C",X"44",X"53",X"20",X"54",X"4F",X"20",X"46",X"49",X"4C",X"4C",X"FD",X"82",X"82",X"53",
		X"48",X"49",X"45",X"4C",X"44",X"20",X"47",X"55",X"41",X"47",X"45",X"FD",X"82",X"C7",X"46",X"49",
		X"4C",X"4C",X"20",X"53",X"48",X"49",X"45",X"4C",X"44",X"20",X"47",X"55",X"41",X"47",X"45",X"20",
		X"46",X"4F",X"52",X"FD",X"82",X"E2",X"45",X"58",X"54",X"52",X"41",X"20",X"53",X"48",X"49",X"50",
		X"FD",X"83",X"27",X"48",X"4F",X"4C",X"44",X"20",X"42",X"4F",X"4D",X"42",X"20",X"42",X"55",X"54",
		X"54",X"4F",X"4E",X"20",X"44",X"4F",X"57",X"4E",X"FD",X"83",X"42",X"46",X"4F",X"52",X"20",X"53",
		X"48",X"49",X"45",X"4C",X"44",X"20",X"55",X"4E",X"54",X"49",X"4C",X"20",X"47",X"55",X"41",X"47",
		X"45",X"20",X"45",X"4D",X"50",X"54",X"59",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"31",X"F7",X"39",X"6F",X"ED",X"79",X"AC",X"CB",X"08",X"ED",X"5A",X"E5",X"26",X"62",X"BA",X"3E",
		X"F8",X"D1",X"12",X"E6",X"E7",X"6F",X"A8",X"77",X"E9",X"33",X"1F",X"1F",X"C9",X"FE",X"35",X"CA",
		X"00",X"31",X"10",X"FC",X"CD",X"F5",X"C7",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
