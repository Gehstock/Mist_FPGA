library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity rom5t32 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of rom5t32 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"77",X"5E",X"00",X"FF",X"75",X"00",X"FF",X"36",X"80",X"FF",X"77",X"80",X"FF",X"5F",X"00",X"80",
		X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"14",X"36",X"00",X"FF",X"14",X"00",
		X"16",X"C2",X"32",X"3D",X"22",X"42",X"6F",X"C3",X"31",X"CA",X"3A",X"42",X"22",X"42",X"CA",X"A7",
		X"DD",X"32",X"C3",X"20",X"17",X"6F",X"FF",X"FF",X"3E",X"17",X"32",X"05",X"22",X"42",X"06",X"3E",
		X"26",X"1D",X"CA",X"A7",X"42",X"55",X"43",X"3A",X"43",X"3A",X"A7",X"22",X"F2",X"CA",X"3A",X"45",
		X"33",X"FE",X"65",X"DA",X"3E",X"42",X"32",X"01",X"3D",X"22",X"43",X"32",X"3A",X"22",X"20",X"D4",
		X"00",X"22",X"00",X"00",X"D3",X"2A",X"3E",X"20",X"22",X"49",X"7B",X"C3",X"AF",X"42",X"49",X"32",
		X"86",X"C3",X"2A",X"42",X"20",X"D3",X"26",X"7C",X"94",X"3D",X"D6",X"85",X"6F",X"01",X"3D",X"26",
		X"3E",X"22",X"32",X"00",X"22",X"46",X"3A",X"C9",X"94",X"25",X"D6",X"85",X"6F",X"02",X"44",X"22",
		X"A7",X"42",X"B2",X"CA",X"AF",X"42",X"48",X"32",X"20",X"E2",X"3A",X"A7",X"22",X"48",X"AA",X"CA",
		X"C9",X"42",X"CA",X"A7",X"42",X"A1",X"32",X"AF",X"3A",X"22",X"22",X"45",X"33",X"FE",X"BB",X"D2",
		X"42",X"BB",X"3A",X"C9",X"22",X"47",X"CA",X"A7",X"22",X"48",X"45",X"3A",X"FE",X"22",X"DA",X"33",
		X"32",X"01",X"22",X"47",X"49",X"3A",X"A7",X"22",X"42",X"C7",X"32",X"3D",X"22",X"47",X"3E",X"C9",
		X"17",X"D2",X"CD",X"43",X"42",X"E9",X"58",X"CD",X"78",X"C2",X"3A",X"47",X"22",X"45",X"26",X"FE",
		X"2A",X"47",X"22",X"44",X"43",X"06",X"46",X"3A",X"3E",X"1D",X"32",X"A0",X"22",X"43",X"F2",X"C3",
		X"57",X"0A",X"FF",X"C9",X"FF",X"FF",X"FF",X"FF",X"E6",X"22",X"87",X"03",X"0A",X"4F",X"03",X"5F",
		X"44",X"2A",X"06",X"22",X"C3",X"47",X"42",X"EE",X"45",X"05",X"44",X"4F",X"44",X"AC",X"44",X"00",
		X"42",X"E9",X"58",X"CD",X"3A",X"1D",X"22",X"46",X"49",X"3A",X"A7",X"22",X"8E",X"C2",X"CD",X"47",
		X"22",X"44",X"D6",X"7D",X"6F",X"40",X"DE",X"7C",X"32",X"3C",X"22",X"46",X"03",X"E6",X"2A",X"F5",
		X"2A",X"43",X"22",X"44",X"C6",X"7D",X"6F",X"1F",X"67",X"00",X"44",X"22",X"F1",X"22",X"47",X"C2",
		X"42",X"E9",X"AA",X"CD",X"C9",X"1D",X"40",X"CD",X"CE",X"7C",X"67",X"00",X"44",X"22",X"CD",X"22",
		X"40",X"A9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CD",X"42",X"46",X"D6",X"28",X"CD",X"C3",X"0A",
		X"20",X"AB",X"01",X"FE",X"7A",X"DA",X"3E",X"43",X"E2",X"3A",X"A7",X"20",X"74",X"CA",X"3A",X"43",
		X"43",X"6A",X"0C",X"3E",X"07",X"36",X"C0",X"C3",X"C3",X"46",X"43",X"7C",X"A7",X"3A",X"C3",X"20",
		X"0F",X"07",X"00",X"FF",X"07",X"00",X"FF",X"07",X"80",X"19",X"0F",X"C0",X"FF",X"1F",X"80",X"00",
		X"FF",X"07",X"00",X"00",X"07",X"07",X"00",X"FF",X"00",X"00",X"07",X"07",X"00",X"FF",X"07",X"00",
		X"00",X"FF",X"02",X"00",X"FF",X"07",X"00",X"00",X"07",X"00",X"FF",X"07",X"00",X"00",X"07",X"07",
		X"00",X"00",X"02",X"02",X"00",X"FF",X"02",X"00",X"02",X"02",X"00",X"FF",X"02",X"00",X"FF",X"02",
		X"00",X"00",X"04",X"0E",X"00",X"FF",X"04",X"00",X"FF",X"02",X"00",X"00",X"02",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"08",X"FF",X"FF",X"00",X"C0",X"FF",X"00",X"00",X"FF",X"1C",X"00",X"FF",X"08",
		X"FF",X"10",X"00",X"00",X"00",X"10",X"FF",X"FF",X"38",X"EF",X"00",X"07",X"00",X"FF",X"38",X"00",
		X"00",X"00",X"01",X"00",X"FF",X"00",X"FF",X"FF",X"00",X"00",X"00",X"80",X"01",X"03",X"00",X"FF",
		X"20",X"3E",X"0F",X"C3",X"3E",X"40",X"D3",X"00",X"E2",X"32",X"3E",X"20",X"D3",X"20",X"C9",X"01",
		X"40",X"FE",X"14",X"C2",X"DF",X"40",X"C3",X"C9",X"21",X"07",X"24",X"00",X"00",X"36",X"7C",X"23",
		X"E2",X"3A",X"A7",X"20",X"35",X"CA",X"F1",X"40",X"0C",X"92",X"FF",X"FF",X"FF",X"FF",X"F5",X"FF",
		X"3B",X"3B",X"C9",X"F1",X"10",X"3E",X"27",X"C3",X"20",X"F6",X"36",X"C3",X"F1",X"40",X"07",X"D3",
		X"C3",X"20",X"40",X"27",X"04",X"21",X"11",X"3E",X"97",X"40",X"27",X"C3",X"97",X"40",X"EA",X"32",
		X"CD",X"D5",X"09",X"F1",X"11",X"00",X"FD",X"E0",X"40",X"90",X"00",X"06",X"02",X"0E",X"C5",X"E5",
		X"C2",X"D5",X"40",X"59",X"C1",X"D1",X"04",X"E1",X"7C",X"19",X"C1",X"D1",X"FE",X"90",X"C5",X"2C",
		X"13",X"13",X"DF",X"D5",X"59",X"C3",X"DF",X"40",X"FE",X"78",X"CA",X"0B",X"40",X"7F",X"C5",X"E5",
		X"20",X"C3",X"FF",X"4E",X"FF",X"FF",X"EA",X"3B",X"DF",X"DF",X"DF",X"DF",X"DF",X"DF",X"DF",X"DF",
		X"26",X"02",X"26",X"26",X"26",X"06",X"26",X"00",X"26",X"19",X"26",X"08",X"26",X"0B",X"26",X"04",
		X"CA",X"43",X"17",X"EA",X"28",X"CD",X"C2",X"0A",X"26",X"0C",X"26",X"04",X"26",X"12",X"4E",X"C3",
		X"17",X"EA",X"3C",X"A7",X"32",X"27",X"20",X"AD",X"40",X"AC",X"AD",X"3A",X"FE",X"20",X"CA",X"99",
		X"F3",X"08",X"45",X"C3",X"3E",X"08",X"D3",X"00",X"E2",X"CD",X"C3",X"09",X"17",X"EA",X"53",X"D2",
		X"41",X"76",X"E2",X"3A",X"A7",X"20",X"E8",X"CA",X"D3",X"01",X"D3",X"06",X"D3",X"07",X"C3",X"04",
		X"03",X"DB",X"E3",X"C3",X"3A",X"40",X"20",X"E2",X"DB",X"40",X"07",X"00",X"C3",X"07",X"15",X"F9",
		X"DB",X"C9",X"E6",X"03",X"C9",X"10",X"23",X"23",X"CA",X"A7",X"40",X"F9",X"00",X"DB",X"10",X"E6",
		X"CD",X"C5",X"0B",X"D3",X"0A",X"C1",X"C5",X"0B",X"23",X"E5",X"2E",X"66",X"C1",X"1D",X"0B",X"0A",
		X"D3",X"C3",X"67",X"0B",X"3A",X"F5",X"20",X"E2",X"D3",X"CD",X"C1",X"0B",X"0B",X"0A",X"C1",X"C5",
		X"00",X"CE",X"32",X"27",X"20",X"AB",X"F1",X"C9",X"CA",X"A7",X"41",X"2F",X"3A",X"F1",X"20",X"AB",
		X"C9",X"20",X"1B",X"2B",X"DA",X"B8",X"41",X"5A",X"A7",X"3A",X"CE",X"20",X"27",X"00",X"A7",X"32",
		X"FF",X"FF",X"1B",X"2B",X"DA",X"B8",X"41",X"6A",X"33",X"C8",X"C3",X"33",X"05",X"03",X"FF",X"FF",
		X"FF",X"FF",X"A5",X"11",X"21",X"20",X"20",X"A1",X"33",X"C8",X"C3",X"33",X"05",X"18",X"FF",X"FF",
		X"FF",X"FF",X"A9",X"11",X"21",X"20",X"20",X"A1",X"03",X"06",X"C3",X"EF",X"05",X"03",X"FF",X"FF",
		X"E2",X"32",X"C3",X"20",X"00",X"B6",X"FF",X"FF",X"03",X"06",X"C3",X"EF",X"05",X"18",X"00",X"3E",
		X"FF",X"05",X"70",X"E8",X"07",X"05",X"50",X"FF",X"78",X"78",X"07",X"05",X"78",X"FF",X"07",X"F8",
		X"40",X"FF",X"01",X"00",X"FF",X"00",X"F0",X"FF",X"07",X"60",X"FF",X"03",X"40",X"60",X"01",X"03",
		X"F0",X"FF",X"0B",X"A0",X"FF",X"0E",X"C0",X"E0",X"0E",X"F0",X"FF",X"0A",X"D0",X"F0",X"0B",X"0E",
		X"00",X"80",X"00",X"02",X"FF",X"FF",X"20",X"E0",X"06",X"0E",X"C0",X"FF",X"06",X"80",X"FF",X"02",
		X"C0",X"E0",X"16",X"17",X"C0",X"FF",X"1B",X"80",X"1D",X"1D",X"E0",X"FF",X"1B",X"E0",X"FF",X"17",
		X"05",X"00",X"FF",X"00",X"C0",X"FF",X"3B",X"C0",X"FF",X"0B",X"00",X"80",X"05",X"0B",X"00",X"FF",
		X"2F",X"80",X"FF",X"2B",X"00",X"80",X"1B",X"3B",X"FF",X"3B",X"C0",X"40",X"2F",X"3A",X"C0",X"FF",
		X"00",X"0A",X"FF",X"FF",X"80",X"80",X"77",X"77",X"00",X"FF",X"1B",X"00",X"FF",X"0A",X"00",X"00",
		X"43",X"DE",X"43",X"D3",X"43",X"C8",X"43",X"81",X"43",X"F0",X"45",X"91",X"45",X"7F",X"45",X"64",
		X"E0",X"FF",X"EC",X"00",X"E1",X"1E",X"00",X"E7",X"80",X"C0",X"FB",X"7F",X"C3",X"C1",X"03",X"01",
		X"0E",X"00",X"F0",X"FF",X"E6",X"00",X"3B",X"10",X"FF",X"07",X"00",X"E0",X"00",X"EA",X"7E",X"71",
		X"3C",X"13",X"08",X"00",X"F0",X"FF",X"E0",X"00",X"00",X"3C",X"FF",X"1C",X"00",X"D0",X"38",X"BF",
		X"27",X"03",X"E0",X"FF",X"EE",X"00",X"01",X"C0",X"03",X"70",X"FF",X"7E",X"00",X"F0",X"E0",X"EA",
		X"C0",X"FF",X"FD",X"00",X"00",X"00",X"FF",X"07",X"FF",X"03",X"00",X"E0",X"80",X"BF",X"03",X"01",
		X"1E",X"00",X"00",X"00",X"FF",X"1C",X"00",X"00",X"00",X"80",X"00",X"7F",X"0E",X"00",X"00",X"FF",
		X"FE",X"5F",X"F0",X"70",X"38",X"FF",X"7B",X"80",X"00",X"00",X"08",X"00",X"FF",X"FF",X"E0",X"F0",
		X"80",X"7A",X"9F",X"1C",X"03",X"00",X"BC",X"FF",X"38",X"C7",X"00",X"F9",X"FF",X"01",X"00",X"B8",
		X"00",X"F4",X"0E",X"EF",X"0F",X"04",X"02",X"00",X"F9",X"00",X"0E",X"04",X"00",X"0F",X"FF",X"07",
		X"00",X"BC",X"F8",X"FA",X"09",X"00",X"B8",X"FF",X"3C",X"FF",X"F8",X"00",X"00",X"9C",X"FF",X"1F",
		X"70",X"FF",X"3F",X"00",X"00",X"C0",X"FF",X"01",X"7B",X"00",X"FF",X"F0",X"00",X"F8",X"E0",X"6F",
		X"07",X"00",X"00",X"00",X"FF",X"07",X"00",X"00",X"00",X"E0",X"80",X"1F",X"03",X"00",X"80",X"FF",
		X"A7",X"22",X"E2",X"CA",X"3D",X"46",X"4A",X"32",X"00",X"00",X"02",X"00",X"FF",X"FF",X"4A",X"3A",
		X"4B",X"3A",X"FE",X"22",X"DA",X"02",X"46",X"F9",X"C9",X"22",X"43",X"3A",X"32",X"22",X"22",X"4A",
		X"3E",X"C9",X"C3",X"08",X"46",X"F2",X"FF",X"FF",X"1F",X"00",X"4B",X"32",X"CD",X"22",X"40",X"27",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"47",X"10",X"46",X"10",X"46",X"76",X"45",X"9E",
		X"80",X"FF",X"B3",X"00",X"87",X"78",X"03",X"9C",X"00",X"00",X"EE",X"FD",X"0F",X"05",X"0F",X"07",
		X"39",X"01",X"C0",X"FF",X"9B",X"00",X"EF",X"40",X"FF",X"1F",X"00",X"80",X"00",X"AB",X"F8",X"C7",
		X"F0",X"4E",X"20",X"00",X"C0",X"FF",X"83",X"00",X"00",X"F0",X"FF",X"70",X"00",X"C0",X"E0",X"FE",
		X"80",X"AB",X"9F",X"0F",X"80",X"FF",X"BB",X"00",X"0F",X"C0",X"00",X"F9",X"FF",X"01",X"00",X"C0",
		X"0E",X"06",X"00",X"FF",X"F7",X"00",X"03",X"00",X"07",X"00",X"FF",X"0F",X"00",X"80",X"00",X"FE",
		X"00",X"FF",X"78",X"00",X"00",X"00",X"FF",X"70",X"FF",X"1C",X"00",X"00",X"00",X"FE",X"38",X"01",
		X"45",X"3A",X"FE",X"22",X"DA",X"3D",X"47",X"8E",X"00",X"00",X"00",X"00",X"20",X"00",X"FF",X"FF",
		X"43",X"32",X"C3",X"22",X"47",X"F8",X"08",X"CD",X"08",X"CD",X"CD",X"43",X"1D",X"58",X"A0",X"3E",
		X"46",X"32",X"E6",X"22",X"F5",X"03",X"44",X"2A",X"CD",X"43",X"1D",X"58",X"46",X"3A",X"3C",X"22",
		X"22",X"67",X"22",X"44",X"C2",X"F1",X"47",X"BE",X"7D",X"22",X"40",X"C6",X"7C",X"6F",X"00",X"CE",
		X"00",X"DE",X"22",X"67",X"22",X"44",X"08",X"CD",X"44",X"2A",X"7D",X"22",X"01",X"D6",X"7C",X"6F",
		X"A7",X"22",X"D2",X"CA",X"3E",X"47",X"32",X"A0",X"CD",X"43",X"1D",X"AA",X"F5",X"C9",X"43",X"3A",
		X"43",X"4A",X"48",X"4F",X"52",X"48",X"49",X"4E",X"22",X"43",X"C3",X"F1",X"01",X"45",X"FF",X"FF",
		X"41",X"48",X"4D",X"42",X"50",X"55",X"45",X"52",X"53",X"20",X"20",X"4C",X"53",X"41",X"54",X"54",
		X"D3",X"AF",X"C3",X"01",X"42",X"7B",X"FF",X"FF",X"52",X"59",X"D3",X"AF",X"C3",X"01",X"42",X"6C",
		X"E0",X"FC",X"E7",X"1F",X"FF",X"1C",X"DC",X"00",X"F8",X"E0",X"3F",X"73",X"3C",X"7E",X"00",X"FF",
		X"C3",X"5E",X"83",X"3D",X"00",X"07",X"FF",X"00",X"1D",X"C1",X"0E",X"C3",X"00",X"01",X"80",X"FF",
		X"7E",X"FE",X"02",X"3F",X"FF",X"01",X"DE",X"00",X"1E",X"00",X"BC",X"E7",X"03",X"07",X"00",X"FF",
		X"9C",X"00",X"1D",X"70",X"00",X"FF",X"E0",X"F8",X"3C",X"3C",X"00",X"FF",X"38",X"5C",X"FF",X"3D",
		X"00",X"FF",X"80",X"C0",X"FF",X"03",X"00",X"FF",X"FF",X"1F",X"F0",X"00",X"0F",X"C0",X"00",X"01",
		X"C0",X"00",X"7F",X"00",X"C1",X"7E",X"01",X"0E",X"3E",X"80",X"E7",X"F7",X"07",X"C3",X"FF",X"03",
		X"FF",X"00",X"E0",X"00",X"D5",X"38",X"73",X"3C",X"00",X"FF",X"10",X"C0",X"3C",X"DD",X"1C",X"E1",
		X"FF",X"3B",X"E0",X"00",X"7F",X"E0",X"13",X"27",X"00",X"08",X"00",X"FF",X"70",X"E0",X"7E",X"C1",
		X"C0",X"00",X"D5",X"80",X"03",X"03",X"00",X"FF",X"00",X"FF",X"C0",X"E0",X"03",X"CD",X"FF",X"03",
		X"7F",X"00",X"01",X"0E",X"00",X"FF",X"00",X"00",X"00",X"C0",X"07",X"D9",X"FF",X"01",X"80",X"00",
		X"00",X"08",X"FF",X"FF",X"E0",X"80",X"FD",X"CF",X"1C",X"EF",X"FF",X"00",X"00",X"00",X"3C",X"00",
		X"9F",X"5F",X"03",X"70",X"FF",X"00",X"70",X"00",X"F0",X"F9",X"00",X"01",X"00",X"FF",X"80",X"F0",
		X"0E",X"78",X"0F",X"F5",X"02",X"1C",X"FF",X"00",X"77",X"04",X"38",X"0F",X"00",X"07",X"00",X"FF",
		X"F8",X"F8",X"09",X"DF",X"FF",X"04",X"78",X"00",X"78",X"00",X"F0",X"9C",X"0E",X"1F",X"00",X"FF",
		X"70",X"00",X"76",X"C0",X"00",X"01",X"00",X"FF",X"F3",X"F0",X"00",X"FF",X"E0",X"70",X"FF",X"F5",
		X"3B",X"00",X"00",X"07",X"00",X"FF",X"00",X"00",X"80",X"E0",X"03",X"5F",X"FF",X"00",X"C0",X"00",
		X"9C",X"DE",X"1F",X"0F",X"FF",X"0F",X"00",X"00",X"02",X"0F",X"FF",X"00",X"00",X"FF",X"F8",X"00",
		X"40",X"00",X"F0",X"77",X"70",X"87",X"FF",X"03",X"FD",X"00",X"07",X"F8",X"07",X"39",X"00",X"FF",
		X"00",X"FF",X"C0",X"80",X"F9",X"07",X"01",X"EF",X"80",X"00",X"57",X"E0",X"CF",X"F0",X"01",X"20",
		X"00",X"FF",X"00",X"80",X"0F",X"37",X"FF",X"0F",X"FF",X"00",X"80",X"00",X"FE",X"80",X"4D",X"9F",
		X"00",X"00",X"1C",X"67",X"FF",X"07",X"00",X"00",X"00",X"00",X"57",X"00",X"0F",X"0E",X"00",X"FF",
		X"70",X"BC",X"FF",X"03",X"00",X"00",X"F0",X"00",X"FE",X"00",X"05",X"38",X"00",X"FF",X"00",X"00",
		X"1F",X"F7",X"00",X"07",X"C0",X"FF",X"DF",X"00",X"00",X"20",X"FF",X"FF",X"C0",X"7F",X"DF",X"DF",
		X"00",X"FF",X"20",X"00",X"FF",X"00",X"00",X"FF",X"1F",X"F8",X"FF",X"00",X"00",X"00",X"20",X"F8",
		X"40",X"E0",X"00",X"FF",X"40",X"00",X"FF",X"00",X"BF",X"00",X"1F",X"E0",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"FF",X"FF",X"F8",X"FC",X"00",X"FF",X"C0",X"00",X"01",X"80",X"FF",X"00",
		X"0E",X"71",X"FF",X"7E",X"00",X"AE",X"E0",X"1E",X"3F",X"17",X"3C",X"1C",X"CE",X"FF",X"1E",X"E0",
		X"00",X"C3",X"FF",X"01",X"80",X"FD",X"C3",X"3F",X"E7",X"07",X"6F",X"FF",X"BE",X"00",X"03",X"C1",
		X"FF",X"07",X"00",X"AF",X"7E",X"3E",X"02",X"00",X"83",X"01",X"0F",X"FF",X"3E",X"00",X"00",X"E7",
		X"38",X"1F",X"FC",X"FF",X"0F",X"00",X"FF",X"70",X"EE",X"FF",X"1E",X"00",X"FF",X"3C",X"00",X"FE",
		X"00",X"C0",X"FF",X"01",X"00",X"00",X"80",X"00",X"00",X"F8",X"E0",X"07",X"E0",X"FF",X"01",X"00",
		X"FF",X"42",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"21",X"3E",X"01",X"D3",X"8F",X"C3");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
