library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity dderby_bg_bits_1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of dderby_bg_bits_1 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"50",X"85",X"54",X"85",X"56",X"95",X"56",X"15",X"56",X"55",X"52",X"55",X"58",X"55",X"48",
		X"00",X"55",X"00",X"05",X"00",X"15",X"00",X"55",X"05",X"55",X"05",X"55",X"01",X"54",X"02",X"52",
		X"55",X"20",X"54",X"80",X"52",X"00",X"48",X"00",X"60",X"00",X"20",X"00",X"80",X"00",X"00",X"00",
		X"00",X"A8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"FF",X"FF",
		X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"FF",X"FF",
		X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"FF",X"FF",
		X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"FF",X"FF",
		X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"FF",X"FF",
		X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"FF",X"FF",
		X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"FF",X"FF",
		X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"FF",X"FF",
		X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"15",X"54",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"15",X"54",
		X"00",X"00",X"00",X"00",X"15",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"15",X"54",
		X"00",X"00",X"00",X"00",X"15",X"54",X"00",X"14",X"15",X"54",X"14",X"00",X"14",X"00",X"15",X"54",
		X"00",X"00",X"00",X"00",X"15",X"54",X"00",X"14",X"15",X"54",X"00",X"14",X"00",X"14",X"15",X"54",
		X"00",X"00",X"00",X"00",X"00",X"14",X"14",X"14",X"14",X"14",X"15",X"54",X"00",X"14",X"00",X"14",
		X"00",X"00",X"00",X"00",X"15",X"54",X"10",X"00",X"15",X"54",X"00",X"14",X"00",X"14",X"15",X"54",
		X"00",X"00",X"00",X"00",X"15",X"54",X"14",X"00",X"14",X"00",X"15",X"54",X"14",X"14",X"15",X"54",
		X"00",X"00",X"00",X"00",X"05",X"54",X"04",X"14",X"00",X"14",X"00",X"14",X"00",X"14",X"00",X"14",
		X"00",X"00",X"00",X"00",X"15",X"54",X"14",X"14",X"15",X"54",X"14",X"14",X"14",X"14",X"15",X"54",
		X"00",X"00",X"00",X"00",X"15",X"54",X"14",X"14",X"14",X"14",X"15",X"54",X"00",X"14",X"15",X"54",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"15",X"54",X"14",X"14",X"14",X"14",X"15",X"54",X"14",X"14",X"14",X"14",
		X"00",X"00",X"00",X"00",X"15",X"50",X"15",X"50",X"14",X"10",X"15",X"54",X"14",X"14",X"15",X"54",
		X"00",X"00",X"00",X"00",X"15",X"54",X"14",X"00",X"14",X"00",X"14",X"00",X"14",X"00",X"15",X"54",
		X"00",X"00",X"00",X"00",X"15",X"50",X"14",X"54",X"14",X"14",X"14",X"14",X"14",X"54",X"15",X"50",
		X"00",X"00",X"00",X"00",X"15",X"54",X"14",X"00",X"15",X"50",X"14",X"00",X"14",X"00",X"15",X"54",
		X"00",X"00",X"00",X"00",X"15",X"50",X"14",X"00",X"14",X"00",X"15",X"40",X"14",X"00",X"14",X"00",
		X"00",X"00",X"00",X"00",X"15",X"54",X"14",X"00",X"14",X"00",X"14",X"14",X"14",X"14",X"15",X"54",
		X"00",X"00",X"00",X"00",X"14",X"14",X"14",X"14",X"14",X"14",X"15",X"54",X"14",X"14",X"14",X"14",
		X"00",X"00",X"00",X"00",X"15",X"54",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"15",X"54",
		X"00",X"00",X"00",X"00",X"01",X"55",X"00",X"14",X"00",X"14",X"14",X"14",X"14",X"14",X"15",X"54",
		X"00",X"00",X"00",X"00",X"14",X"54",X"15",X"40",X"15",X"00",X"15",X"40",X"14",X"50",X"14",X"14",
		X"00",X"00",X"00",X"00",X"14",X"00",X"14",X"00",X"14",X"00",X"14",X"00",X"14",X"14",X"15",X"54",
		X"00",X"00",X"00",X"00",X"15",X"54",X"14",X"44",X"14",X"44",X"14",X"44",X"14",X"44",X"14",X"44",
		X"00",X"00",X"00",X"00",X"14",X"14",X"15",X"14",X"15",X"54",X"14",X"54",X"14",X"54",X"14",X"14",
		X"00",X"00",X"00",X"00",X"15",X"54",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"15",X"54",
		X"00",X"00",X"00",X"00",X"15",X"54",X"14",X"14",X"14",X"14",X"15",X"54",X"14",X"00",X"14",X"00",
		X"00",X"00",X"00",X"00",X"15",X"54",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"54",X"15",X"54",
		X"00",X"00",X"00",X"00",X"15",X"54",X"14",X"14",X"15",X"54",X"14",X"50",X"14",X"14",X"14",X"14",
		X"00",X"00",X"00",X"00",X"15",X"50",X"10",X"00",X"15",X"50",X"00",X"50",X"00",X"50",X"15",X"50",
		X"00",X"00",X"00",X"00",X"15",X"54",X"11",X"44",X"01",X"40",X"01",X"40",X"01",X"40",X"05",X"50",
		X"00",X"00",X"00",X"00",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"15",X"54",
		X"00",X"00",X"00",X"00",X"15",X"14",X"05",X"10",X"05",X"10",X"05",X"50",X"01",X"40",X"01",X"40",
		X"00",X"00",X"00",X"00",X"14",X"44",X"14",X"44",X"14",X"44",X"14",X"44",X"14",X"44",X"15",X"54",
		X"00",X"00",X"00",X"00",X"15",X"14",X"05",X"10",X"01",X"40",X"04",X"50",X"10",X"10",X"10",X"14",
		X"00",X"00",X"00",X"00",X"14",X"14",X"05",X"10",X"05",X"40",X"01",X"40",X"01",X"40",X"01",X"40",
		X"00",X"00",X"00",X"00",X"15",X"54",X"00",X"50",X"01",X"40",X"05",X"00",X"14",X"00",X"15",X"54",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"DF",X"AB",X"FD",X"AA",X"DD",X"6B",X"DF",X"AA",X"FD",X"AB",X"DD",X"6A",X"DF",X"AB",X"FD",X"AA",
		X"99",X"A5",X"55",X"55",X"55",X"96",X"59",X"65",X"55",X"55",X"3F",X"FF",X"99",X"66",X"55",X"55",
		X"95",X"56",X"69",X"66",X"55",X"95",X"55",X"56",X"05",X"55",X"56",X"9A",X"12",X"55",X"51",X"56",
		X"55",X"55",X"96",X"59",X"55",X"55",X"55",X"95",X"55",X"55",X"A9",X"59",X"95",X"55",X"55",X"65",
		X"56",X"59",X"55",X"55",X"95",X"55",X"51",X"65",X"55",X"51",X"FF",X"FD",X"59",X"65",X"55",X"55",
		X"59",X"65",X"59",X"55",X"59",X"64",X"55",X"95",X"55",X"55",X"3F",X"FF",X"91",X"49",X"55",X"55",
		X"10",X"44",X"96",X"65",X"99",X"65",X"59",X"65",X"59",X"65",X"6A",X"A9",X"95",X"55",X"95",X"95",
		X"90",X"21",X"95",X"65",X"95",X"69",X"66",X"59",X"66",X"55",X"A6",X"65",X"95",X"55",X"95",X"65",
		X"00",X"64",X"95",X"65",X"95",X"A5",X"99",X"96",X"59",X"96",X"69",X"56",X"65",X"95",X"65",X"95",
		X"94",X"09",X"59",X"19",X"5A",X"59",X"5A",X"65",X"55",X"65",X"3F",X"FF",X"99",X"66",X"55",X"55",
		X"CC",X"DF",X"F0",X"1F",X"CC",X"DF",X"F0",X"1F",X"CC",X"DF",X"F0",X"1F",X"CC",X"DF",X"F0",X"1F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",X"FF",X"F5",X"FF",X"FF",X"FF",X"E6",X"F7",X"DD",X"FB",
		X"FF",X"F5",X"FF",X"FD",X"FF",X"F5",X"FF",X"D5",X"FF",X"55",X"F7",X"55",X"FF",X"55",X"FF",X"D5",
		X"55",X"55",X"55",X"5B",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"FF",X"55",X"57",X"55",X"5F",X"55",X"FF",X"55",X"D9",X"57",X"F7",X"57",X"FF",X"7D",X"FF",
		X"DB",X"FF",X"D7",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"5F",X"57",X"57",X"75",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"D5",X"57",X"FD",X"DF",X"FF",X"FF",
		X"FF",X"D5",X"7F",X"FD",X"FF",X"D5",X"FF",X"5D",X"FF",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FE",X"FE",X"7F",X"FF",X"FF",X"EF",X"FF",X"FB",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"7F",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"E7",X"FF",X"D7",X"FF",X"FF",X"FF",X"FF",X"FB",X"FF",X"D7",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"E7",X"FF",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"F9",X"FD",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"5F",X"FF",X"7F",X"FF",X"F7",X"FF",X"5F",X"FF",
		X"FF",X"75",X"7D",X"57",X"55",X"5F",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"7F",X"FD",X"5D",X"75",X"D7",X"55",X"D5",X"55",X"55",X"55",X"D5",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"D5",X"FF",X"F5",
		X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"CC",X"DF",X"F0",X"1F",X"CC",X"DD",X"F0",X"1F",X"CC",X"DE",X"F0",X"1F",X"CC",X"DF",X"F0",X"1F",
		X"FD",X"AB",X"DD",X"6A",X"DF",X"AB",X"FD",X"AA",X"DD",X"6B",X"DF",X"AA",X"FD",X"AB",X"DD",X"6A",
		X"DD",X"6A",X"DF",X"AB",X"FD",X"AB",X"DD",X"6A",X"DF",X"AB",X"FD",X"AA",X"DD",X"6B",X"DF",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"B3",X"33",X"CC",X"CC",X"F3",X"00",X"CC",X"CC",X"F0",X"35",X"CC",X"DF",X"F0",X"1F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"FF",X"FF",
		X"00",X"00",X"95",X"55",X"95",X"55",X"95",X"55",X"95",X"55",X"95",X"55",X"95",X"55",X"FF",X"FF",
		X"00",X"00",X"A5",X"55",X"A5",X"55",X"A5",X"55",X"A5",X"55",X"A5",X"55",X"A5",X"55",X"FF",X"FF",
		X"00",X"00",X"A9",X"55",X"A9",X"55",X"A9",X"55",X"A9",X"55",X"A9",X"55",X"A9",X"55",X"FF",X"FF",
		X"00",X"00",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"FF",X"FF",
		X"00",X"00",X"AA",X"95",X"AA",X"95",X"AA",X"95",X"AA",X"95",X"AA",X"95",X"AA",X"95",X"FF",X"FF",
		X"00",X"00",X"AA",X"A5",X"AA",X"A5",X"AA",X"A5",X"AA",X"A5",X"AA",X"A5",X"AA",X"A5",X"FF",X"FF",
		X"00",X"00",X"AA",X"A9",X"AA",X"A9",X"AA",X"A9",X"AA",X"A9",X"AA",X"A9",X"AA",X"A9",X"FF",X"FF",
		X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"2A",X"A8",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"2A",X"A8",
		X"00",X"00",X"00",X"00",X"2A",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"2A",X"A8",
		X"00",X"00",X"00",X"00",X"2A",X"A8",X"00",X"28",X"2A",X"A8",X"28",X"00",X"28",X"00",X"2A",X"A8",
		X"00",X"00",X"00",X"00",X"2A",X"A8",X"00",X"28",X"2A",X"A8",X"00",X"28",X"00",X"28",X"2A",X"A8",
		X"00",X"00",X"00",X"00",X"00",X"28",X"28",X"28",X"28",X"28",X"2A",X"A8",X"00",X"28",X"00",X"28",
		X"00",X"00",X"00",X"00",X"2A",X"A8",X"20",X"00",X"2A",X"A8",X"00",X"28",X"00",X"28",X"2A",X"A8",
		X"00",X"00",X"00",X"00",X"2A",X"A8",X"28",X"00",X"28",X"00",X"2A",X"A8",X"28",X"28",X"2A",X"A8",
		X"00",X"00",X"00",X"00",X"0A",X"A8",X"08",X"28",X"00",X"28",X"00",X"28",X"00",X"28",X"00",X"28",
		X"00",X"00",X"00",X"00",X"2A",X"A8",X"28",X"28",X"2A",X"A8",X"28",X"28",X"28",X"28",X"2A",X"A8",
		X"00",X"00",X"00",X"00",X"2A",X"A8",X"28",X"28",X"28",X"28",X"2A",X"A8",X"00",X"28",X"2A",X"A8",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"2A",X"A8",X"28",X"28",X"28",X"28",X"2A",X"A8",X"28",X"28",X"28",X"28",
		X"00",X"00",X"00",X"00",X"2A",X"A0",X"2A",X"A0",X"28",X"20",X"2A",X"A8",X"28",X"28",X"2A",X"A8",
		X"00",X"00",X"00",X"00",X"2A",X"A8",X"28",X"00",X"28",X"00",X"28",X"00",X"28",X"00",X"2A",X"A8",
		X"00",X"00",X"00",X"00",X"2A",X"A0",X"28",X"A8",X"28",X"28",X"28",X"28",X"28",X"A8",X"2A",X"A0",
		X"00",X"00",X"00",X"00",X"2A",X"A8",X"28",X"00",X"2A",X"A0",X"28",X"00",X"28",X"00",X"2A",X"A8",
		X"00",X"00",X"00",X"00",X"2A",X"A0",X"28",X"00",X"28",X"00",X"2A",X"80",X"28",X"00",X"28",X"00",
		X"00",X"00",X"00",X"00",X"2A",X"A8",X"28",X"00",X"28",X"00",X"28",X"28",X"28",X"28",X"2A",X"A8",
		X"00",X"00",X"00",X"00",X"28",X"28",X"28",X"28",X"28",X"28",X"2A",X"A8",X"28",X"28",X"28",X"28",
		X"00",X"00",X"00",X"00",X"2A",X"A8",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"2A",X"A8",
		X"00",X"00",X"00",X"00",X"02",X"AA",X"00",X"28",X"00",X"28",X"28",X"28",X"28",X"28",X"2A",X"A8",
		X"00",X"00",X"00",X"00",X"28",X"A8",X"2A",X"80",X"2A",X"00",X"2A",X"80",X"28",X"A0",X"28",X"28",
		X"00",X"00",X"00",X"00",X"28",X"00",X"28",X"00",X"28",X"00",X"28",X"00",X"28",X"28",X"2A",X"A8",
		X"00",X"00",X"00",X"00",X"2A",X"A8",X"28",X"88",X"28",X"88",X"28",X"88",X"28",X"88",X"28",X"88",
		X"00",X"00",X"00",X"00",X"28",X"28",X"2A",X"28",X"2A",X"A8",X"28",X"A8",X"28",X"A8",X"28",X"28",
		X"00",X"00",X"00",X"00",X"2A",X"A8",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"2A",X"A8",
		X"00",X"00",X"00",X"00",X"2A",X"A8",X"28",X"28",X"28",X"28",X"2A",X"A8",X"28",X"00",X"28",X"00",
		X"00",X"00",X"00",X"00",X"2A",X"A8",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"A8",X"2A",X"A8",
		X"00",X"00",X"00",X"00",X"2A",X"A8",X"28",X"28",X"2A",X"A8",X"28",X"A0",X"28",X"28",X"28",X"28",
		X"00",X"00",X"00",X"00",X"2A",X"A0",X"20",X"00",X"2A",X"A0",X"00",X"A0",X"00",X"A0",X"2A",X"A0",
		X"00",X"00",X"00",X"00",X"2A",X"A8",X"22",X"88",X"02",X"80",X"02",X"80",X"02",X"80",X"0A",X"A0",
		X"00",X"00",X"00",X"00",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"2A",X"A8",
		X"00",X"00",X"00",X"00",X"2A",X"28",X"0A",X"20",X"0A",X"20",X"0A",X"A0",X"02",X"80",X"02",X"80",
		X"00",X"00",X"00",X"00",X"28",X"88",X"28",X"88",X"28",X"88",X"28",X"88",X"28",X"88",X"2A",X"A8",
		X"00",X"00",X"00",X"00",X"2A",X"28",X"0A",X"20",X"02",X"80",X"08",X"A0",X"20",X"20",X"20",X"28",
		X"00",X"00",X"00",X"00",X"28",X"28",X"0A",X"20",X"0A",X"80",X"02",X"80",X"02",X"80",X"02",X"80",
		X"00",X"00",X"00",X"00",X"2A",X"A8",X"00",X"A0",X"02",X"80",X"0A",X"00",X"28",X"00",X"2A",X"A8",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"33",X"33",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"55",X"55",X"FF",X"FF",X"FD",X"FD",
		X"FF",X"FF",X"33",X"33",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"55",X"55",X"FF",X"FF",X"E7",X"9F",
		X"FF",X"FF",X"33",X"33",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"55",X"55",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"30",X"C3",X"FF",X"FF",X"5D",X"75",X"61",X"86",X"AA",X"AA",X"AA",X"AA",X"EE",X"EE",
		X"FF",X"FF",X"C3",X"0C",X"FF",X"FF",X"75",X"D7",X"86",X"18",X"AA",X"AA",X"AA",X"AA",X"EE",X"EE",
		X"FF",X"FF",X"5C",X"75",X"FF",X"FF",X"D7",X"5D",X"18",X"61",X"AA",X"AA",X"AA",X"AA",X"EE",X"EE",
		X"FF",X"FF",X"30",X"C3",X"FF",X"FF",X"1C",X"71",X"61",X"86",X"AA",X"AA",X"AA",X"AA",X"EE",X"EE",
		X"02",X"FF",X"0F",X"4C",X"39",X"3F",X"B5",X"E7",X"D7",X"44",X"D2",X"6A",X"DD",X"AA",X"FD",X"AA",
		X"15",X"46",X"0A",X"15",X"5F",X"45",X"55",X"55",X"15",X"5F",X"15",X"55",X"1F",X"55",X"15",X"55",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"C1",X"A1",X"06",X"A8",X"06",X"A4",X"C5",X"15",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"00",
		X"A9",X"55",X"A5",X"3D",X"55",X"15",X"55",X"55",X"55",X"55",X"55",X"F5",X"55",X"55",X"55",X"55",
		X"54",X"01",X"55",X"E5",X"15",X"A9",X"55",X"25",X"7D",X"55",X"55",X"55",X"55",X"5F",X"55",X"55",
		X"AA",X"54",X"A5",X"57",X"55",X"57",X"55",X"57",X"5F",X"56",X"55",X"56",X"55",X"56",X"40",X"54",
		X"00",X"00",X"00",X"00",X"00",X"00",X"39",X"00",X"AA",X"4C",X"41",X"50",X"00",X"50",X"6D",X"5E",
		X"00",X"00",X"00",X"00",X"00",X"01",X"40",X"41",X"40",X"11",X"5B",X"55",X"6A",X"55",X"59",X"05",
		X"00",X"00",X"00",X"00",X"00",X"41",X"6D",X"00",X"69",X"7D",X"06",X"69",X"01",X"65",X"E5",X"55",
		X"AA",X"22",X"AA",X"88",X"8A",X"A2",X"A2",X"A8",X"88",X"AA",X"A2",X"28",X"88",X"A0",X"A2",X"20",
		X"22",X"2A",X"88",X"AA",X"22",X"A2",X"8A",X"8A",X"AA",X"22",X"28",X"8A",X"0A",X"22",X"08",X"8A",
		X"02",X"22",X"02",X"8A",X"00",X"A2",X"20",X"2A",X"80",X"22",X"20",X"0A",X"80",X"02",X"AA",X"AA",
		X"88",X"80",X"A2",X"80",X"8A",X"00",X"A8",X"00",X"88",X"00",X"A0",X"00",X"80",X"00",X"AA",X"AA",
		X"55",X"55",X"15",X"55",X"15",X"55",X"15",X"55",X"05",X"55",X"01",X"55",X"01",X"55",X"00",X"55",
		X"55",X"55",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"50",X"55",X"40",X"55",X"40",X"55",X"00",
		X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"85",X"00",X"15",X"00",X"55",X"01",X"55",
		X"55",X"40",X"55",X"50",X"55",X"50",X"55",X"54",X"05",X"56",X"41",X"56",X"61",X"56",X"25",X"56",
		X"85",X"56",X"15",X"52",X"D5",X"48",X"55",X"20",X"54",X"80",X"52",X"00",X"48",X"00",X"A0",X"00",
		X"05",X"54",X"05",X"52",X"15",X"49",X"55",X"43",X"55",X"55",X"54",X"55",X"02",X"55",X"00",X"AA",
		X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"02",X"00",X"0D",X"00",X"05",X"00",X"55",X"00",X"D5",
		X"55",X"55",X"55",X"55",X"55",X"54",X"55",X"56",X"55",X"02",X"54",X"A8",X"55",X"50",X"55",X"58",
		X"00",X"95",X"03",X"55",X"01",X"54",X"01",X"55",X"01",X"55",X"03",X"55",X"00",X"55",X"00",X"2A",
		X"55",X"78",X"00",X"20",X"2A",X"80",X"54",X"00",X"56",X"00",X"52",X"00",X"48",X"00",X"A0",X"00",
		X"00",X"55",X"01",X"55",X"01",X"55",X"05",X"54",X"05",X"54",X"05",X"56",X"01",X"52",X"02",X"A8",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"05",X"00",X"05",X"00",X"15",X"00",X"15",X"00",X"55",
		X"15",X"00",X"55",X"40",X"55",X"61",X"55",X"65",X"55",X"15",X"55",X"55",X"55",X"55",X"55",X"55",
		X"15",X"51",X"15",X"51",X"15",X"41",X"15",X"45",X"95",X"95",X"0A",X"15",X"00",X"01",X"00",X"02",
		X"54",X"80",X"54",X"80",X"56",X"00",X"52",X"00",X"52",X"00",X"58",X"00",X"58",X"00",X"A0",X"00",
		X"15",X"80",X"55",X"40",X"55",X"60",X"55",X"60",X"55",X"60",X"55",X"20",X"55",X"20",X"55",X"80",
		X"55",X"00",X"55",X"50",X"55",X"54",X"55",X"56",X"55",X"56",X"45",X"56",X"25",X"56",X"95",X"56",
		X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"05",X"00",X"15",X"00",X"55",X"01",X"55",X"05",X"54",
		X"05",X"54",X"05",X"51",X"05",X"55",X"05",X"55",X"01",X"55",X"00",X"55",X"00",X"25",X"00",X"0A",
		X"95",X"52",X"55",X"58",X"55",X"48",X"55",X"20",X"54",X"80",X"52",X"00",X"68",X"00",X"A0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"05",X"00",X"05",X"00",X"15",
		X"00",X"55",X"00",X"55",X"01",X"55",X"01",X"55",X"01",X"55",X"00",X"55",X"00",X"15",X"00",X"0A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"05",X"00",X"15",X"40",X"55",X"40",X"55",X"60",X"55",X"60",X"55",X"20",X"54",X"80",X"56",X"00",
		X"52",X"00",X"48",X"00",X"40",X"00",X"55",X"00",X"55",X"80",X"55",X"80",X"5A",X"00",X"A0",X"00",
		X"01",X"40",X"05",X"50",X"15",X"54",X"15",X"54",X"55",X"58",X"55",X"58",X"55",X"60",X"55",X"60",
		X"55",X"80",X"55",X"80",X"54",X"80",X"56",X"00",X"52",X"00",X"58",X"00",X"48",X"00",X"A0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",
		X"00",X"05",X"00",X"05",X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"05",X"00",X"00",
		X"55",X"54",X"55",X"55",X"55",X"56",X"55",X"56",X"55",X"42",X"55",X"48",X"55",X"60",X"55",X"20",
		X"00",X"15",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"0A",X"00",X"05",X"00",X"01",
		X"00",X"05",X"00",X"15",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"15",X"00",X"05",X"00",X"0A",
		X"55",X"80",X"54",X"80",X"56",X"00",X"52",X"00",X"58",X"00",X"48",X"00",X"20",X"00",X"80",X"00",
		X"00",X"05",X"00",X"15",X"00",X"15",X"00",X"55",X"00",X"55",X"01",X"55",X"01",X"55",X"05",X"55",
		X"00",X"50",X"81",X"54",X"61",X"55",X"65",X"55",X"45",X"56",X"45",X"56",X"55",X"58",X"55",X"48",
		X"05",X"55",X"15",X"51",X"15",X"51",X"55",X"51",X"55",X"41",X"15",X"41",X"05",X"49",X"0A",X"A0",
		X"55",X"60",X"55",X"20",X"55",X"80",X"55",X"80",X"54",X"80",X"54",X"80",X"54",X"80",X"AA",X"00",
		X"00",X"15",X"00",X"55",X"00",X"55",X"00",X"55",X"01",X"55",X"01",X"55",X"01",X"55",X"05",X"55",
		X"55",X"40",X"55",X"50",X"55",X"54",X"55",X"55",X"41",X"55",X"25",X"55",X"95",X"54",X"55",X"52",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"05",X"55",X"05",X"55",X"15",X"55",X"15",X"55",X"55",X"51",X"55",X"41",X"15",X"48",X"0A",X"A0",
		X"55",X"48",X"51",X"A0",X"52",X"00",X"54",X"00",X"55",X"00",X"55",X"60",X"55",X"60",X"15",X"80",
		X"00",X"01",X"00",X"15",X"00",X"55",X"00",X"55",X"80",X"55",X"80",X"25",X"80",X"15",X"00",X"55",
		X"2A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"40",X"55",X"50",X"55",X"54",X"55",X"54",X"55",X"56",X"51",X"56",X"49",X"56",X"55",X"52",
		X"00",X"55",X"01",X"55",X"01",X"55",X"01",X"55",X"01",X"56",X"01",X"55",X"01",X"55",X"00",X"55",
		X"55",X"48",X"15",X"60",X"95",X"60",X"55",X"60",X"55",X"60",X"55",X"60",X"55",X"80",X"56",X"00",
		X"01",X"55",X"02",X"55",X"01",X"54",X"05",X"55",X"05",X"55",X"15",X"55",X"05",X"55",X"09",X"15",
		X"00",X"2A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"0F",X"00",X"0D",
		X"00",X"0A",X"00",X"95",X"02",X"95",X"09",X"56",X"D5",X"59",X"55",X"63",X"F1",X"7F",X"01",X"FF",
		X"80",X"00",X"70",X"01",X"55",X"55",X"AF",X"44",X"6A",X"D4",X"DA",X"B5",X"F9",X"AA",X"FA",X"66",
		X"00",X"00",X"40",X"03",X"D0",X"32",X"F4",X"D9",X"37",X"36",X"68",X"0F",X"AF",X"FF",X"95",X"59",
		X"00",X"0C",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"57",X"FF",X"57",X"17",X"5C",X"65",X"3D",X"99",X"30",X"45",X"35",X"39",X"35",X"F5",X"35",X"F5",
		X"FA",X"99",X"C9",X"55",X"E9",X"5A",X"E5",X"6A",X"D9",X"5A",X"D6",X"55",X"F5",X"95",X"FF",X"69",
		X"5A",X"A6",X"AA",X"95",X"AA",X"67",X"A9",X"97",X"AA",X"5F",X"6A",X"5E",X"56",X"7A",X"59",X"6A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",
		X"34",X"F4",X"35",X"17",X"35",X"57",X"35",X"53",X"0D",X"0F",X"03",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"C3",X"FF",X"00",X"3F",X"00",X"0F",X"0F",X"0F",X"00",X"03",
		X"95",X"6A",X"EA",X"AA",X"FF",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",
		X"00",X"C0",X"00",X"00",X"03",X"30",X"00",X"FF",X"00",X"0F",X"C0",X"00",X"C0",X"03",X"3C",X"00",
		X"00",X"00",X"00",X"04",X"00",X"00",X"30",X"00",X"3C",X"F0",X"3C",X"00",X"0C",X"31",X"FC",X"00",
		X"FC",X"F0",X"31",X"55",X"00",X"55",X"05",X"55",X"01",X"54",X"35",X"41",X"71",X"01",X"05",X"46",
		X"00",X"00",X"2A",X"00",X"79",X"80",X"AE",X"60",X"AF",X"CF",X"FF",X"FB",X"FE",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FC",X"BB",X"BB",X"AA",X"BF",X"AA",X"AB",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"BF",X"00",X"EE",X"00",
		X"00",X"C0",X"0C",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"30",
		X"AA",X"AA",X"BE",X"A7",X"FA",X"9F",X"EA",X"7F",X"A9",X"FF",X"A8",X"FC",X"A7",X"F6",X"93",X"DA",
		X"72",X"AA",X"FF",X"EA",X"FF",X"FA",X"FF",X"FA",X"FF",X"FA",X"0F",X"FA",X"A3",X"FF",X"A8",X"F5",
		X"FE",X"00",X"EF",X"80",X"FE",X"20",X"BE",X"B8",X"A7",X"BC",X"E4",X"38",X"E9",X"6E",X"CA",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"03",X"00",X"3F",X"03",X"FC",X"40",X"0F",X"90",X"0F",
		X"9F",X"29",X"7F",X"A1",X"3D",X"B7",X"FD",X"9F",X"FD",X"7C",X"FD",X"71",X"FD",X"63",X"FD",X"64",
		X"98",X"36",X"5A",X"36",X"D6",X"FD",X"F6",X"1D",X"F6",X"7F",X"F6",X"DF",X"76",X"7F",X"55",X"FF",
		X"72",X"BF",X"9C",X"AF",X"A7",X"2B",X"A9",X"CA",X"6A",X"72",X"DA",X"9C",X"F6",X"A7",X"FD",X"A9",
		X"EC",X"3F",X"FB",X"00",X"FE",X"C0",X"FF",X"F3",X"BB",X"BF",X"AA",X"23",X"2B",X"2F",X"CE",X"00",
		X"1D",X"59",X"5C",X"56",X"5F",X"55",X"57",X"15",X"57",X"D1",X"41",X"FF",X"00",X"65",X"00",X"15",
		X"55",X"7F",X"94",X"FF",X"50",X"FF",X"47",X"CC",X"1F",X"15",X"FC",X"5A",X"55",X"56",X"95",X"95",
		X"FF",X"6A",X"FF",X"DA",X"0F",X"F5",X"3C",X"FD",X"3C",X"FF",X"FC",X"FF",X"3F",X"FC",X"BF",X"FC",
		X"73",X"2C",X"9C",X"F0",X"A7",X"00",X"57",X"C0",X"FF",X"C0",X"3D",X"00",X"F1",X"00",X"01",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"00",X"3C",X"00",X"00",X"00",X"00",X"30",X"30",X"00",X"03",X"0C",X"00",
		X"00",X"C0",X"00",X"31",X"00",X"30",X"3C",X"30",X"00",X"30",X"00",X"C0",X"C0",X"00",X"03",X"00",
		X"00",X"55",X"05",X"55",X"01",X"5D",X"04",X"40",X"01",X"50",X"00",X"54",X"00",X"40",X"43",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"00",X"30",X"03",X"F3",X"00",X"0F",X"03",X"CC",X"C0",X"F3",X"0F",X"00",X"00",X"C0",
		X"FC",X"00",X"0F",X"00",X"C0",X"00",X"CC",X"00",X"3F",X"00",X"00",X"00",X"03",X"00",X"30",X"00",
		X"03",X"14",X"00",X"05",X"00",X"55",X"01",X"45",X"04",X"05",X"00",X"54",X"04",X"15",X"00",X"15",
		X"C0",X"00",X"00",X"00",X"00",X"C0",X"C0",X"00",X"00",X"03",X"00",X"0F",X"00",X"3F",X"00",X"00",
		X"00",X"3F",X"00",X"F3",X"00",X"0F",X"00",X"30",X"00",X"30",X"33",X"C0",X"FF",X"FC",X"FC",X"0F",
		X"00",X"00",X"C3",X"00",X"3C",X"30",X"00",X"C0",X"F0",X"0F",X"C0",X"3C",X"03",X"03",X"FF",X"FF",
		X"00",X"05",X"00",X"44",X"C0",X"05",X"3C",X"03",X"00",X"0C",X"C0",X"3F",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"30",X"00",X"0F",X"FF",X"00",X"F3",X"C0",X"FF",
		X"00",X"CF",X"FF",X"FF",X"00",X"0F",X"03",X"FF",X"0C",X"FF",X"F0",X"F0",X"FF",X"C0",X"FF",X"F0",
		X"FF",X"FC",X"0F",X"FF",X"FF",X"FC",X"FF",X"F3",X"FF",X"FF",X"40",X"44",X"CF",X"F0",X"03",X"C0",
		X"3F",X"3C",X"30",X"00",X"C3",X"04",X"00",X"04",X"00",X"00",X"40",X"FF",X"3F",X"05",X"55",X"55",
		X"45",X"5C",X"16",X"51",X"65",X"01",X"55",X"81",X"55",X"00",X"05",X"05",X"05",X"55",X"05",X"55",
		X"55",X"61",X"55",X"A2",X"59",X"14",X"6A",X"45",X"59",X"98",X"69",X"59",X"5A",X"46",X"5A",X"A6",
		X"83",X"FD",X"9F",X"C3",X"99",X"44",X"AA",X"98",X"A5",X"53",X"A4",X"C0",X"99",X"54",X"75",X"95",
		X"15",X"40",X"15",X"40",X"54",X"00",X"D5",X"40",X"55",X"40",X"55",X"00",X"55",X"40",X"55",X"50",
		X"55",X"59",X"55",X"66",X"55",X"69",X"55",X"65",X"55",X"55",X"55",X"55",X"15",X"05",X"58",X"4C",
		X"9A",X"9A",X"69",X"EA",X"AA",X"AA",X"AB",X"AB",X"6A",X"AB",X"66",X"BA",X"5A",X"AE",X"46",X"AA",
		X"00",X"8D",X"31",X"45",X"06",X"16",X"56",X"6D",X"99",X"6A",X"E9",X"AD",X"AE",X"A9",X"A9",X"A9",
		X"55",X"40",X"55",X"40",X"55",X"40",X"95",X"40",X"55",X"00",X"95",X"13",X"65",X"00",X"95",X"03",
		X"5C",X"44",X"71",X"55",X"D5",X"53",X"13",X"3F",X"F0",X"3C",X"FF",X"0C",X"FF",X"00",X"FF",X"00",
		X"41",X"AB",X"A1",X"1A",X"04",X"41",X"F3",X"0F",X"CC",X"CF",X"FF",X"FF",X"CC",X"34",X"54",X"5A",
		X"AA",X"05",X"A6",X"31",X"80",X"3C",X"FF",X"F0",X"C0",X"33",X"00",X"0F",X"15",X"55",X"59",X"55",
		X"51",X"03",X"55",X"03",X"30",X"0C",X"CF",X"3F",X"FC",X"C0",X"0F",X"FF",X"53",X"FF",X"40",X"0F",
		X"00",X"55",X"15",X"55",X"55",X"55",X"55",X"55",X"14",X"50",X"FC",X"05",X"55",X"55",X"55",X"55",
		X"69",X"9A",X"A6",X"AA",X"56",X"95",X"95",X"0C",X"3C",X"FF",X"44",X"05",X"55",X"54",X"55",X"00",
		X"55",X"54",X"A5",X"55",X"55",X"50",X"30",X"FC",X"FF",X"FF",X"00",X"00",X"40",X"00",X"10",X"00",
		X"03",X"FF",X"0C",X"F3",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"3F",X"00",X"F3",X"F0");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
