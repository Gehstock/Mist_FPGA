`define BUILD_DATE "190831"
`define BUILD_TIME "162534"
