library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity guzzler_prog2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of guzzler_prog2 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"21",X"71",X"85",X"CB",X"C6",X"21",X"80",X"83",X"06",X"80",X"AF",X"77",X"23",X"10",X"FC",X"21",
		X"4B",X"E0",X"CD",X"7B",X"5C",X"3E",X"23",X"06",X"02",X"FF",X"3A",X"80",X"83",X"FE",X"01",X"20",
		X"F4",X"3E",X"23",X"06",X"3C",X"FF",X"21",X"75",X"E0",X"22",X"1C",X"80",X"21",X"20",X"84",X"22",
		X"29",X"80",X"21",X"55",X"E0",X"CD",X"7B",X"5C",X"3E",X"23",X"06",X"02",X"FF",X"3A",X"80",X"83",
		X"FE",X"02",X"20",X"F4",X"21",X"65",X"E0",X"CD",X"73",X"5C",X"C9",X"03",X"9F",X"E0",X"04",X"BA",
		X"E0",X"05",X"D5",X"E0",X"FF",X"03",X"09",X"E2",X"04",X"25",X"E4",X"05",X"39",X"E4",X"06",X"00",
		X"E6",X"07",X"60",X"3D",X"FF",X"11",X"12",X"13",X"14",X"15",X"16",X"17",X"18",X"19",X"1A",X"1B",
		X"1C",X"1D",X"1E",X"1F",X"FF",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"93",X"E0",X"96",X"E0",X"00",
		X"00",X"00",X"00",X"01",X"12",X"91",X"02",X"81",X"D4",X"92",X"80",X"00",X"90",X"FF",X"FF",X"31",
		X"20",X"87",X"DD",X"21",X"98",X"83",X"21",X"4E",X"80",X"22",X"A5",X"83",X"DD",X"36",X"01",X"01",
		X"DD",X"36",X"0C",X"03",X"DD",X"36",X"0B",X"7E",X"18",X"34",X"31",X"00",X"87",X"DD",X"21",X"B0",
		X"83",X"21",X"55",X"80",X"22",X"BD",X"83",X"DD",X"36",X"01",X"02",X"DD",X"36",X"0C",X"02",X"DD",
		X"36",X"0B",X"9E",X"18",X"19",X"31",X"E0",X"86",X"DD",X"21",X"C8",X"83",X"21",X"5C",X"80",X"22",
		X"D5",X"83",X"DD",X"36",X"01",X"04",X"DD",X"36",X"0C",X"01",X"DD",X"36",X"0B",X"BE",X"DD",X"36",
		X"09",X"01",X"DD",X"7E",X"0C",X"06",X"01",X"CD",X"7C",X"36",X"DD",X"75",X"05",X"DD",X"74",X"06",
		X"DD",X"5E",X"0D",X"DD",X"56",X"0E",X"D5",X"13",X"13",X"13",X"ED",X"A0",X"7E",X"DD",X"77",X"02",
		X"23",X"DD",X"75",X"03",X"DD",X"74",X"04",X"EB",X"36",X"10",X"23",X"36",X"40",X"DD",X"36",X"0A",
		X"40",X"23",X"DD",X"7E",X"0B",X"77",X"E1",X"36",X"00",X"3E",X"23",X"06",X"3C",X"FF",X"DD",X"CB",
		X"00",X"7E",X"C2",X"93",X"E1",X"DD",X"CB",X"00",X"76",X"C2",X"EF",X"E1",X"DD",X"7E",X"0A",X"FE",
		X"90",X"38",X"48",X"DD",X"CB",X"01",X"46",X"20",X"13",X"3A",X"81",X"83",X"DD",X"CB",X"01",X"4E",
		X"28",X"06",X"FE",X"01",X"28",X"06",X"18",X"36",X"FE",X"02",X"38",X"32",X"CD",X"3E",X"E3",X"DD",
		X"6E",X"0D",X"DD",X"66",X"0E",X"E5",X"23",X"23",X"23",X"77",X"23",X"23",X"34",X"E1",X"36",X"00",
		X"DD",X"E5",X"E1",X"11",X"09",X"00",X"19",X"01",X"04",X"00",X"11",X"69",X"83",X"ED",X"B0",X"3E",
		X"01",X"01",X"A0",X"36",X"FF",X"DD",X"CB",X"00",X"FE",X"18",X"6B",X"CD",X"5B",X"E3",X"CD",X"08",
		X"E3",X"18",X"63",X"3A",X"73",X"80",X"CB",X"7F",X"20",X"5C",X"DD",X"6E",X"0D",X"DD",X"66",X"0E",
		X"E5",X"11",X"06",X"00",X"19",X"E1",X"36",X"00",X"DD",X"CB",X"01",X"56",X"20",X"0E",X"DD",X"CB",
		X"00",X"BE",X"DD",X"CB",X"00",X"F6",X"21",X"81",X"83",X"34",X"18",X"3A",X"3E",X"23",X"06",X"3C",
		X"FF",X"FD",X"21",X"80",X"80",X"11",X"0B",X"00",X"FD",X"CB",X"01",X"7E",X"28",X"0E",X"FD",X"CB",
		X"02",X"46",X"28",X"08",X"FD",X"36",X"00",X"40",X"FD",X"CB",X"01",X"BE",X"FD",X"19",X"FD",X"7E",
		X"00",X"FE",X"FF",X"20",X"E3",X"21",X"81",X"83",X"36",X"03",X"2B",X"36",X"01",X"18",X"0F",X"3A",
		X"81",X"83",X"FE",X"03",X"28",X"08",X"3E",X"23",X"06",X"02",X"FF",X"C3",X"2E",X"E1",X"DD",X"6E",
		X"0D",X"DD",X"66",X"0E",X"36",X"40",X"3E",X"60",X"FF",X"31",X"20",X"87",X"DD",X"21",X"98",X"83",
		X"DD",X"E5",X"E1",X"AF",X"06",X"18",X"77",X"23",X"10",X"FC",X"3E",X"23",X"06",X"10",X"FF",X"DD",
		X"36",X"09",X"01",X"DD",X"36",X"0A",X"00",X"DD",X"36",X"0B",X"A0",X"DD",X"36",X"0C",X"04",X"21",
		X"4E",X"80",X"22",X"A5",X"83",X"3E",X"04",X"06",X"01",X"CD",X"7C",X"36",X"22",X"9D",X"83",X"11",
		X"51",X"80",X"ED",X"A0",X"7E",X"DD",X"77",X"02",X"23",X"22",X"9B",X"83",X"EB",X"36",X"10",X"23",
		X"36",X"00",X"23",X"36",X"A0",X"AF",X"32",X"4E",X"80",X"DD",X"CB",X"00",X"7E",X"28",X"34",X"3A",
		X"73",X"80",X"CB",X"7F",X"C2",X"EE",X"E2",X"DD",X"CB",X"00",X"BE",X"DD",X"34",X"0C",X"DD",X"7E",
		X"0C",X"DD",X"46",X"09",X"CD",X"7C",X"36",X"22",X"9D",X"83",X"11",X"51",X"80",X"ED",X"A0",X"7E",
		X"DD",X"77",X"02",X"23",X"22",X"9B",X"83",X"AF",X"32",X"4E",X"80",X"DD",X"7E",X"07",X"FE",X"03",
		X"CA",X"F6",X"E2",X"CD",X"5B",X"E3",X"CD",X"08",X"E3",X"DD",X"CB",X"00",X"76",X"20",X"0F",X"CD",
		X"C3",X"E3",X"B7",X"28",X"09",X"DD",X"CB",X"00",X"F6",X"3E",X"02",X"CD",X"DC",X"34",X"DD",X"46",
		X"0A",X"DD",X"4E",X"07",X"78",X"FE",X"50",X"38",X"35",X"79",X"B7",X"28",X"0F",X"78",X"FE",X"70",
		X"38",X"2C",X"79",X"FE",X"01",X"28",X"05",X"78",X"FE",X"A0",X"38",X"22",X"CD",X"3E",X"E3",X"32",
		X"51",X"80",X"AF",X"32",X"4E",X"80",X"11",X"69",X"83",X"21",X"A1",X"83",X"01",X"04",X"00",X"ED",
		X"B0",X"3E",X"01",X"01",X"AA",X"36",X"FF",X"DD",X"CB",X"00",X"FE",X"DD",X"34",X"07",X"3E",X"23",
		X"06",X"02",X"FF",X"C3",X"59",X"E2",X"3E",X"23",X"06",X"3C",X"FF",X"3E",X"40",X"32",X"4E",X"80",
		X"3E",X"02",X"32",X"80",X"83",X"3E",X"60",X"FF",X"DD",X"7E",X"02",X"B7",X"28",X"04",X"DD",X"35",
		X"02",X"C9",X"DD",X"6E",X"03",X"DD",X"66",X"04",X"7E",X"FE",X"FF",X"20",X"06",X"DD",X"6E",X"05",
		X"DD",X"66",X"06",X"DD",X"5E",X"0D",X"DD",X"56",X"0E",X"D5",X"13",X"13",X"13",X"ED",X"A0",X"7E",
		X"DD",X"77",X"02",X"23",X"DD",X"75",X"03",X"DD",X"74",X"04",X"E1",X"36",X"00",X"C9",X"21",X"2E",
		X"7A",X"11",X"04",X"00",X"DD",X"7E",X"0C",X"3D",X"28",X"03",X"19",X"18",X"FA",X"DD",X"7E",X"09",
		X"CB",X"3F",X"FE",X"04",X"20",X"01",X"3D",X"5F",X"19",X"7E",X"C9",X"DD",X"7E",X"08",X"B7",X"28",
		X"04",X"DD",X"35",X"08",X"C9",X"DD",X"6E",X"0D",X"DD",X"66",X"0E",X"E5",X"DD",X"7E",X"09",X"11",
		X"05",X"00",X"E6",X"03",X"20",X"01",X"13",X"19",X"DD",X"7E",X"09",X"CB",X"47",X"28",X"09",X"7E",
		X"C6",X"02",X"77",X"DD",X"77",X"0A",X"18",X"21",X"CB",X"4F",X"28",X"09",X"7E",X"D6",X"02",X"77",
		X"DD",X"77",X"0A",X"18",X"14",X"CB",X"57",X"28",X"09",X"7E",X"D6",X"02",X"77",X"DD",X"77",X"0B",
		X"18",X"07",X"7E",X"C6",X"02",X"77",X"DD",X"77",X"0B",X"E1",X"36",X"00",X"DD",X"7E",X"0C",X"FE",
		X"04",X"30",X"0A",X"DD",X"CB",X"00",X"6E",X"20",X"04",X"3E",X"02",X"18",X"02",X"3E",X"01",X"DD",
		X"77",X"08",X"C9",X"DD",X"6E",X"0D",X"DD",X"66",X"0E",X"23",X"23",X"23",X"11",X"54",X"85",X"AF",
		X"12",X"13",X"01",X"04",X"00",X"ED",X"B0",X"3E",X"01",X"12",X"21",X"80",X"80",X"E5",X"23",X"CB",
		X"7E",X"28",X"1C",X"23",X"23",X"23",X"23",X"11",X"5A",X"85",X"ED",X"A0",X"ED",X"A0",X"23",X"23",
		X"ED",X"A0",X"ED",X"A0",X"3E",X"01",X"21",X"54",X"85",X"CD",X"30",X"55",X"B7",X"20",X"0D",X"E1",
		X"11",X"0B",X"00",X"19",X"7E",X"FE",X"FF",X"20",X"D4",X"AF",X"18",X"18",X"E1",X"E5",X"23",X"4E",
		X"79",X"E6",X"7F",X"06",X"00",X"E6",X"03",X"20",X"08",X"06",X"02",X"CB",X"61",X"20",X"02",X"06",
		X"01",X"E1",X"3E",X"01",X"C9",X"31",X"00",X"87",X"DD",X"21",X"E0",X"83",X"21",X"55",X"80",X"22",
		X"E7",X"83",X"3E",X"23",X"06",X"08",X"FF",X"18",X"16",X"31",X"E0",X"86",X"DD",X"21",X"F0",X"83",
		X"21",X"5C",X"80",X"22",X"F7",X"83",X"DD",X"36",X"00",X"01",X"3E",X"23",X"06",X"C0",X"FF",X"DD",
		X"CB",X"00",X"7E",X"20",X"03",X"CD",X"7D",X"E4",X"DD",X"6E",X"07",X"DD",X"66",X"08",X"23",X"23",
		X"CB",X"7E",X"28",X"06",X"CD",X"29",X"E5",X"3E",X"60",X"FF",X"DD",X"CB",X"00",X"76",X"20",X"03",
		X"CD",X"99",X"E5",X"CD",X"63",X"E5",X"3E",X"23",X"06",X"03",X"FF",X"18",X"D2",X"DD",X"CB",X"00",
		X"76",X"20",X"5B",X"21",X"21",X"84",X"CB",X"76",X"20",X"04",X"CB",X"66",X"28",X"07",X"3E",X"23",
		X"06",X"01",X"FF",X"18",X"EE",X"CB",X"F6",X"23",X"36",X"40",X"DD",X"6E",X"07",X"DD",X"66",X"08",
		X"E5",X"23",X"36",X"84",X"23",X"36",X"00",X"23",X"EB",X"21",X"81",X"7A",X"DD",X"CB",X"00",X"46",
		X"28",X"03",X"21",X"86",X"7A",X"DD",X"75",X"04",X"DD",X"74",X"05",X"ED",X"A0",X"7E",X"DD",X"77",
		X"01",X"23",X"DD",X"75",X"02",X"DD",X"74",X"03",X"EB",X"36",X"12",X"23",X"36",X"B0",X"23",X"36",
		X"A0",X"E1",X"36",X"00",X"DD",X"36",X"09",X"20",X"DD",X"CB",X"00",X"F6",X"18",X"4A",X"DD",X"7E",
		X"09",X"B7",X"28",X"05",X"DD",X"35",X"09",X"18",X"3F",X"DD",X"CB",X"00",X"B6",X"DD",X"CB",X"00",
		X"FE",X"21",X"58",X"7A",X"DD",X"CB",X"00",X"46",X"28",X"03",X"21",X"70",X"7A",X"DD",X"75",X"04",
		X"DD",X"74",X"05",X"DD",X"5E",X"07",X"DD",X"56",X"08",X"D5",X"13",X"13",X"13",X"ED",X"A0",X"7E",
		X"DD",X"77",X"01",X"23",X"DD",X"75",X"02",X"DD",X"74",X"03",X"EB",X"36",X"12",X"DD",X"CB",X"00",
		X"46",X"28",X"02",X"36",X"16",X"E1",X"36",X"00",X"C9",X"DD",X"6E",X"07",X"DD",X"66",X"08",X"E5",
		X"23",X"23",X"23",X"36",X"3D",X"23",X"36",X"10",X"E1",X"36",X"00",X"E5",X"AF",X"32",X"2D",X"80",
		X"3E",X"23",X"06",X"40",X"FF",X"E1",X"E5",X"23",X"23",X"23",X"36",X"3F",X"23",X"36",X"0E",X"E1",
		X"36",X"00",X"3E",X"23",X"06",X"40",X"FF",X"DD",X"6E",X"07",X"DD",X"66",X"08",X"36",X"40",X"23",
		X"CB",X"BE",X"C9",X"DD",X"7E",X"01",X"B7",X"28",X"04",X"DD",X"35",X"01",X"C9",X"DD",X"6E",X"02",
		X"DD",X"66",X"03",X"7E",X"FE",X"FF",X"20",X"06",X"DD",X"6E",X"04",X"DD",X"66",X"05",X"DD",X"5E",
		X"07",X"DD",X"56",X"08",X"D5",X"13",X"13",X"13",X"ED",X"A0",X"7E",X"DD",X"77",X"01",X"23",X"DD",
		X"75",X"02",X"DD",X"74",X"03",X"E1",X"36",X"00",X"C9",X"DD",X"6E",X"07",X"DD",X"66",X"08",X"E5",
		X"11",X"05",X"00",X"19",X"7E",X"DD",X"CB",X"00",X"46",X"20",X"04",X"D6",X"02",X"18",X"02",X"D6",
		X"03",X"77",X"E1",X"36",X"00",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"31",X"A0",X"87",X"FD",X"2A",X"29",X"80",X"FD",X"23",X"DD",X"21",X"42",X"84",X"01",X"01",X"00",
		X"18",X"3F",X"31",X"80",X"87",X"FD",X"2A",X"29",X"80",X"01",X"05",X"00",X"FD",X"09",X"DD",X"21",
		X"4C",X"84",X"01",X"03",X"00",X"18",X"2A",X"31",X"60",X"87",X"FD",X"2A",X"29",X"80",X"01",X"09",
		X"00",X"FD",X"09",X"DD",X"21",X"56",X"84",X"01",X"05",X"00",X"18",X"15",X"31",X"40",X"87",X"FD",
		X"2A",X"29",X"80",X"01",X"0D",X"00",X"FD",X"09",X"DD",X"21",X"60",X"84",X"01",X"07",X"00",X"18",
		X"00",X"CD",X"1A",X"E8",X"3E",X"23",X"06",X"02",X"FF",X"DD",X"6E",X"04",X"DD",X"66",X"05",X"23",
		X"23",X"CB",X"7E",X"CA",X"15",X"E7",X"FD",X"CB",X"00",X"FE",X"FD",X"CB",X"00",X"DE",X"3E",X"36",
		X"CD",X"CA",X"1B",X"21",X"42",X"79",X"CD",X"68",X"E8",X"E1",X"DD",X"46",X"01",X"3E",X"23",X"FF",
		X"E1",X"01",X"05",X"00",X"09",X"3E",X"FF",X"BE",X"20",X"EC",X"3E",X"23",X"06",X"01",X"FF",X"3A",
		X"70",X"85",X"CB",X"4F",X"28",X"09",X"3A",X"24",X"85",X"CB",X"7F",X"20",X"06",X"18",X"EB",X"CB",
		X"67",X"20",X"E7",X"DD",X"6E",X"04",X"DD",X"66",X"05",X"23",X"23",X"CB",X"6E",X"28",X"4C",X"3A",
		X"71",X"85",X"CB",X"47",X"28",X"05",X"21",X"CC",X"E8",X"18",X"1E",X"11",X"A8",X"E8",X"DD",X"6E",
		X"04",X"DD",X"66",X"05",X"23",X"23",X"CB",X"76",X"EB",X"28",X"03",X"21",X"B0",X"E8",X"3A",X"71",
		X"85",X"CB",X"7F",X"20",X"04",X"23",X"23",X"23",X"23",X"11",X"54",X"85",X"01",X"04",X"00",X"ED",
		X"B0",X"3E",X"01",X"21",X"54",X"85",X"01",X"00",X"08",X"DD",X"5E",X"04",X"DD",X"56",X"05",X"CD",
		X"80",X"53",X"FD",X"CB",X"00",X"DE",X"3E",X"23",X"06",X"40",X"FF",X"FD",X"CB",X"00",X"9E",X"DD",
		X"6E",X"04",X"DD",X"66",X"05",X"36",X"40",X"23",X"CB",X"BE",X"FD",X"36",X"02",X"00",X"FD",X"36",
		X"03",X"00",X"3E",X"60",X"FF",X"3A",X"71",X"85",X"CB",X"47",X"20",X"55",X"2A",X"29",X"80",X"7E",
		X"FE",X"01",X"20",X"4D",X"21",X"71",X"85",X"CB",X"6E",X"20",X"0B",X"3A",X"00",X"C0",X"FE",X"04",
		X"38",X"3F",X"CB",X"EE",X"18",X"3B",X"21",X"DA",X"E8",X"06",X"05",X"0E",X"00",X"5E",X"23",X"56",
		X"23",X"1A",X"B7",X"20",X"01",X"0C",X"10",X"F5",X"79",X"FE",X"02",X"38",X"24",X"06",X"07",X"21",
		X"8C",X"82",X"11",X"08",X"00",X"7E",X"FE",X"00",X"28",X"04",X"19",X"04",X"18",X"F7",X"78",X"01",
		X"83",X"44",X"FF",X"21",X"00",X"C7",X"01",X"40",X"00",X"16",X"00",X"CD",X"82",X"5A",X"3E",X"60",
		X"FF",X"FD",X"CB",X"00",X"76",X"28",X"6C",X"FD",X"35",X"01",X"28",X"36",X"FD",X"CB",X"00",X"6E",
		X"20",X"14",X"3E",X"37",X"CD",X"CA",X"1B",X"FD",X"CB",X"00",X"EE",X"21",X"DC",X"78",X"CD",X"68",
		X"E8",X"E1",X"E1",X"C3",X"54",X"E6",X"DD",X"35",X"01",X"C2",X"54",X"E6",X"DD",X"6E",X"02",X"DD",
		X"66",X"03",X"3E",X"FF",X"BE",X"20",X"03",X"21",X"DC",X"78",X"CD",X"68",X"E8",X"E1",X"E1",X"C3",
		X"54",X"E6",X"FD",X"CB",X"00",X"AE",X"FD",X"CB",X"00",X"B6",X"2A",X"29",X"80",X"23",X"06",X"04",
		X"11",X"04",X"00",X"CB",X"7E",X"20",X"04",X"CB",X"76",X"20",X"08",X"19",X"10",X"F5",X"3E",X"57",
		X"CD",X"CA",X"1B",X"FD",X"CB",X"00",X"E6",X"DD",X"36",X"06",X"10",X"21",X"80",X"78",X"CD",X"68",
		X"E8",X"E1",X"E1",X"FD",X"CB",X"00",X"66",X"28",X"0F",X"DD",X"7E",X"06",X"B7",X"28",X"05",X"DD",
		X"35",X"06",X"18",X"04",X"FD",X"CB",X"00",X"A6",X"DD",X"35",X"01",X"C2",X"54",X"E6",X"DD",X"6E",
		X"02",X"DD",X"66",X"03",X"3E",X"FF",X"BE",X"20",X"09",X"21",X"80",X"78",X"DD",X"75",X"02",X"DD",
		X"74",X"03",X"CD",X"68",X"E8",X"E1",X"E1",X"C3",X"54",X"E6",X"2A",X"1C",X"80",X"11",X"16",X"00",
		X"19",X"5E",X"23",X"56",X"EB",X"09",X"5E",X"23",X"56",X"FD",X"73",X"02",X"FD",X"72",X"03",X"21",
		X"80",X"78",X"23",X"23",X"23",X"23",X"7E",X"DD",X"77",X"01",X"23",X"DD",X"75",X"02",X"DD",X"74",
		X"03",X"11",X"54",X"85",X"21",X"80",X"78",X"01",X"04",X"00",X"ED",X"B0",X"FD",X"7E",X"02",X"12",
		X"13",X"FD",X"7E",X"03",X"12",X"3E",X"00",X"06",X"08",X"0E",X"00",X"21",X"54",X"85",X"CD",X"80",
		X"53",X"DD",X"75",X"04",X"DD",X"74",X"05",X"C9",X"5D",X"54",X"E3",X"E5",X"EB",X"11",X"54",X"85",
		X"01",X"04",X"00",X"ED",X"B0",X"7E",X"DD",X"77",X"01",X"23",X"DD",X"75",X"02",X"DD",X"74",X"03",
		X"E3",X"E5",X"3E",X"01",X"01",X"00",X"08",X"DD",X"5E",X"04",X"DD",X"56",X"05",X"21",X"54",X"85",
		X"CD",X"80",X"53",X"C9",X"02",X"04",X"00",X"00",X"C4",X"C5",X"00",X"00",X"C6",X"C7",X"02",X"04",
		X"00",X"00",X"CC",X"CD",X"00",X"00",X"CE",X"CF",X"94",X"E8",X"00",X"0A",X"B8",X"E8",X"00",X"0A",
		X"9E",X"E8",X"00",X"0A",X"C2",X"E8",X"00",X"0A",X"02",X"04",X"00",X"00",X"68",X"69",X"00",X"00",
		X"6A",X"6B",X"02",X"04",X"00",X"00",X"70",X"71",X"00",X"00",X"72",X"73",X"D0",X"E8",X"00",X"0E",
		X"02",X"04",X"00",X"00",X"C4",X"C5",X"00",X"00",X"C6",X"C7",X"80",X"83",X"A0",X"83",X"C0",X"83",
		X"E0",X"83",X"00",X"84",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"6C",X"78",X"00",X"72",X"78",X"08",X"96",X"78",X"01",X"A8",X"84",X"08",X"B6",X"90",X"04",
		X"C0",X"96",X"08",X"C0",X"90",X"98",X"C0",X"9C",X"88",X"C0",X"9C",X"80",X"C0",X"9C",X"00",X"C0",
		X"9C",X"01",X"C0",X"B3",X"00",X"CC",X"C0",X"04",X"CE",X"C0",X"00",X"D8",X"B0",X"90",X"D8",X"A9",
		X"80",X"D8",X"A9",X"00",X"D8",X"A9",X"08",X"D8",X"A9",X"00",X"D8",X"C8",X"02",X"D8",X"CA",X"00",
		X"90",X"D8",X"01",X"8D",X"D8",X"91",X"92",X"D8",X"81",X"92",X"D8",X"00",X"B3",X"D8",X"02",X"B8",
		X"D8",X"00",X"5E",X"D8",X"01",X"5C",X"D8",X"91",X"6E",X"D8",X"81",X"6E",X"D8",X"00",X"80",X"D8",
		X"02",X"82",X"D8",X"00",X"5A",X"D8",X"04",X"58",X"D8",X"94",X"48",X"A8",X"84",X"48",X"A8",X"00",
		X"48",X"A5",X"08",X"48",X"A2",X"02",X"48",X"B2",X"91",X"33",X"C0",X"81",X"33",X"C0",X"04",X"53",
		X"C0",X"01",X"60",X"B2",X"04",X"72",X"A8",X"00",X"78",X"8C",X"08",X"78",X"8A",X"00",X"78",X"9E",
		X"04",X"78",X"A0",X"00",X"78",X"50",X"02",X"78",X"4A",X"01",X"6E",X"48",X"08",X"B8",X"48",X"98",
		X"C0",X"4A",X"88",X"C0",X"4A",X"80",X"C0",X"4A",X"04",X"C0",X"4A",X"02",X"C0",X"38",X"00",X"B3",
		X"30",X"04",X"B0",X"30",X"00",X"A8",X"21",X"02",X"A8",X"1E",X"08",X"93",X"18",X"04",X"78",X"2B",
		X"02",X"78",X"18",X"00",X"39",X"18",X"08",X"36",X"18",X"98",X"30",X"22",X"88",X"30",X"22",X"80",
		X"30",X"22",X"04",X"30",X"22",X"02",X"30",X"18",X"08",X"1E",X"18",X"00",X"18",X"62",X"04",X"18",
		X"65",X"94",X"18",X"5F",X"84",X"18",X"5F",X"00",X"18",X"5F",X"08",X"18",X"5F",X"01",X"18",X"9B",
		X"91",X"1A",X"A8",X"81",X"1A",X"A8",X"00",X"86",X"18",X"08",X"84",X"18",X"00",X"78",X"28",X"04",
		X"78",X"2C",X"00",X"78",X"1F",X"02",X"78",X"1C",X"00",X"65",X"18",X"08",X"3B",X"18",X"98",X"30",
		X"27",X"88",X"30",X"27",X"80",X"30",X"27",X"00",X"30",X"27",X"00",X"B3",X"30",X"04",X"AC",X"30",
		X"02",X"A8",X"20",X"00",X"86",X"18",X"08",X"84",X"18",X"04",X"78",X"2C",X"02",X"78",X"1C",X"00",
		X"41",X"18",X"08",X"3E",X"18",X"00",X"30",X"23",X"04",X"30",X"27",X"08",X"30",X"18",X"00",X"30",
		X"25",X"01",X"30",X"27",X"00",X"4A",X"30",X"02",X"4D",X"30",X"00",X"30",X"30",X"01",X"30",X"30",
		X"91",X"36",X"30",X"81",X"36",X"30",X"02",X"5B",X"30",X"92",X"50",X"30",X"82",X"50",X"30",X"01",
		X"33",X"C0",X"04",X"50",X"C0",X"01",X"60",X"B0",X"91",X"76",X"A8",X"81",X"76",X"A8",X"80",X"76",
		X"A8",X"00",X"C0",X"4D",X"02",X"C0",X"5D",X"00",X"B0",X"60",X"08",X"AD",X"60",X"00",X"A8",X"6D",
		X"02",X"A8",X"6F",X"00",X"8B",X"78",X"08",X"88",X"78",X"98",X"78",X"7E",X"88",X"78",X"7E",X"00",
		X"78",X"92",X"04",X"78",X"95",X"00",X"78",X"7B",X"02",X"78",X"78",X"00",X"5E",X"78",X"90",X"4B",
		X"78",X"80",X"4B",X"78",X"00",X"48",X"78",X"04",X"35",X"78",X"00",X"30",X"66",X"01",X"30",X"63",
		X"04",X"55",X"60",X"01",X"60",X"4B",X"08",X"75",X"48",X"00",X"78",X"60",X"04",X"78",X"A5",X"94",
		X"78",X"86",X"84",X"78",X"86",X"00",X"78",X"83",X"08",X"78",X"80",X"00",X"78",X"97",X"01",X"78",
		X"9A",X"04",X"8B",X"A8",X"00",X"90",X"96",X"01",X"90",X"94",X"08",X"B3",X"90",X"00",X"C0",X"B8",
		X"01",X"C0",X"BA",X"08",X"D6",X"C0",X"00",X"D8",X"D8",X"02",X"D8",X"D8",X"00",X"BB",X"D8",X"01",
		X"B8",X"D8",X"00",X"C8",X"D8",X"02",X"CB",X"D8",X"92",X"C4",X"D8",X"82",X"C4",X"00",X"00",X"00",
		X"08",X"76",X"78",X"01",X"78",X"88",X"08",X"86",X"90",X"98",X"90",X"96",X"88",X"90",X"96",X"00",
		X"90",X"96",X"02",X"90",X"A8",X"92",X"7C",X"A8",X"82",X"7C",X"A8",X"80",X"7C",X"A8",X"00",X"74",
		X"A8",X"04",X"56",X"A8",X"00",X"48",X"95",X"01",X"48",X"92",X"04",X"6D",X"90",X"94",X"78",X"71",
		X"84",X"78",X"71",X"00",X"78",X"6A",X"01",X"78",X"68",X"91",X"78",X"63",X"81",X"78",X"60",X"04",
		X"A2",X"60",X"02",X"A8",X"4A",X"01",X"4A",X"48",X"91",X"54",X"48",X"81",X"54",X"48",X"80",X"54",
		X"48",X"94",X"78",X"6B",X"84",X"78",X"6B",X"00",X"78",X"55",X"02",X"78",X"52",X"08",X"4E",X"48",
		X"01",X"48",X"5B",X"91",X"58",X"60",X"81",X"58",X"60",X"91",X"84",X"60",X"81",X"84",X"60",X"02",
		X"64",X"D8",X"00",X"51",X"D8",X"04",X"1A",X"D8",X"00",X"18",X"C6",X"01",X"18",X"89",X"00",X"27",
		X"78",X"90",X"58",X"78",X"80",X"58",X"78",X"00",X"58",X"78",X"04",X"70",X"78",X"02",X"78",X"65",
		X"92",X"76",X"60",X"82",X"76",X"60",X"00",X"76",X"60",X"04",X"54",X"60",X"08",X"48",X"4C",X"00",
		X"48",X"59",X"01",X"48",X"5C",X"00",X"5B",X"60",X"90",X"72",X"60",X"80",X"72",X"60",X"04",X"43",
		X"78",X"00",X"30",X"5B",X"01",X"30",X"41",X"00",X"50",X"30",X"08",X"6D",X"30",X"01",X"78",X"40",
		X"08",X"8D",X"48",X"98",X"90",X"4D",X"88",X"90",X"4D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"76",X"78",X"08",X"89",X"78",X"00",X"90",X"88",X"02",X"90",X"8A",X"00",X"6E",X"90",X"01",
		X"62",X"90",X"91",X"72",X"90",X"81",X"72",X"90",X"04",X"72",X"90",X"01",X"78",X"7C",X"00",X"8B",
		X"78",X"08",X"B8",X"78",X"00",X"C0",X"87",X"90",X"C0",X"9A",X"80",X"C0",X"9A",X"04",X"C0",X"9A",
		X"00",X"C0",X"65",X"02",X"C0",X"63",X"00",X"AD",X"60",X"04",X"AA",X"60",X"01",X"A8",X"50",X"91",
		X"AE",X"48",X"81",X"AE",X"48",X"00",X"AE",X"48",X"02",X"AE",X"48",X"08",X"97",X"48",X"04",X"90",
		X"5B",X"02",X"90",X"4B",X"00",X"76",X"48",X"90",X"4C",X"48",X"80",X"4C",X"48",X"00",X"4C",X"48",
		X"08",X"1F",X"48",X"00",X"18",X"52",X"90",X"18",X"5F",X"80",X"18",X"5F",X"00",X"18",X"5F",X"01",
		X"18",X"5F",X"08",X"2B",X"60",X"00",X"30",X"77",X"90",X"30",X"8F",X"80",X"30",X"8F",X"00",X"80",
		X"60",X"08",X"7D",X"60",X"00",X"78",X"72",X"04",X"78",X"75",X"01",X"78",X"55",X"00",X"85",X"48",
		X"90",X"8B",X"48",X"80",X"8B",X"48",X"00",X"8B",X"48",X"90",X"B0",X"48",X"80",X"B0",X"48",X"00",
		X"B0",X"48",X"08",X"CD",X"48",X"00",X"D8",X"5D",X"02",X"D8",X"5F",X"00",X"C2",X"60",X"04",X"71",
		X"60",X"00",X"60",X"50",X"02",X"60",X"4D",X"90",X"4C",X"48",X"80",X"4C",X"48",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C3",X"AB",X"F0",X"CD",X"12",X"F0",X"21",X"08",X"C1",X"11",X"80",X"98",X"01",X"20",X"00",X"ED",
		X"B0",X"C9",X"DD",X"21",X"28",X"C1",X"DD",X"CB",X"00",X"7E",X"C8",X"DD",X"CB",X"00",X"76",X"28",
		X"11",X"21",X"00",X"88",X"36",X"00",X"2C",X"20",X"FB",X"21",X"FD",X"98",X"36",X"00",X"2C",X"20",
		X"FB",X"C9",X"11",X"2C",X"C1",X"DD",X"7E",X"00",X"E6",X"0F",X"21",X"F0",X"88",X"B7",X"28",X"19",
		X"CB",X"3F",X"30",X"11",X"F5",X"1A",X"D5",X"E5",X"11",X"F0",X"FF",X"06",X"04",X"77",X"3C",X"19",
		X"10",X"FB",X"E1",X"D1",X"F1",X"13",X"23",X"18",X"E4",X"DD",X"7E",X"00",X"E6",X"F0",X"DD",X"77",
		X"00",X"DD",X"7E",X"02",X"DD",X"CB",X"01",X"6E",X"28",X"02",X"D6",X"60",X"5F",X"DD",X"7E",X"03",
		X"DD",X"CB",X"01",X"66",X"28",X"02",X"D6",X"60",X"57",X"DD",X"4E",X"01",X"3A",X"00",X"B8",X"CB",
		X"67",X"20",X"11",X"3A",X"00",X"80",X"CB",X"6F",X"28",X"0A",X"3E",X"10",X"A9",X"4F",X"7A",X"C6",
		X"08",X"57",X"18",X"04",X"3E",X"88",X"92",X"57",X"79",X"32",X"FD",X"98",X"7B",X"32",X"FE",X"98",
		X"7A",X"32",X"FF",X"98",X"C9",X"5E",X"23",X"56",X"23",X"EB",X"C9",X"ED",X"73",X"08",X"C2",X"31",
		X"80",X"C2",X"3E",X"23",X"06",X"2D",X"FF",X"21",X"30",X"C1",X"06",X"B4",X"36",X"00",X"23",X"10",
		X"FB",X"21",X"00",X"C1",X"06",X"30",X"36",X"00",X"23",X"10",X"FB",X"FD",X"21",X"00",X"C1",X"21",
		X"24",X"C0",X"CB",X"C6",X"21",X"63",X"90",X"01",X"1A",X"1A",X"11",X"06",X"00",X"C5",X"36",X"00",
		X"2C",X"10",X"FB",X"C1",X"19",X"0D",X"20",X"F5",X"3A",X"00",X"80",X"CB",X"6F",X"20",X"05",X"3A",
		X"D4",X"85",X"18",X"03",X"3A",X"D5",X"85",X"3D",X"FD",X"77",X"00",X"3D",X"FE",X"1F",X"38",X"02",
		X"3E",X"1E",X"F5",X"5F",X"16",X"00",X"21",X"45",X"F2",X"19",X"7E",X"FD",X"77",X"01",X"F1",X"6F",
		X"26",X"00",X"29",X"29",X"11",X"68",X"F2",X"19",X"FD",X"75",X"02",X"FD",X"74",X"03",X"3E",X"23",
		X"06",X"10",X"FF",X"DD",X"21",X"1C",X"F2",X"CD",X"8A",X"5A",X"3E",X"23",X"06",X"10",X"FF",X"21",
		X"A9",X"91",X"DD",X"21",X"13",X"C0",X"16",X"9C",X"1E",X"07",X"06",X"05",X"0E",X"00",X"CD",X"B9",
		X"5B",X"3A",X"71",X"85",X"CB",X"7F",X"28",X"39",X"3E",X"23",X"06",X"10",X"FF",X"DD",X"21",X"29",
		X"F2",X"CD",X"8A",X"5A",X"11",X"00",X"C2",X"21",X"13",X"C0",X"01",X"05",X"00",X"ED",X"B0",X"21",
		X"04",X"C2",X"11",X"17",X"C0",X"06",X"05",X"CD",X"75",X"5B",X"3E",X"23",X"06",X"10",X"FF",X"21",
		X"A9",X"91",X"DD",X"21",X"13",X"C0",X"16",X"9C",X"1E",X"07",X"06",X"05",X"0E",X"00",X"CD",X"B9",
		X"5B",X"3E",X"23",X"06",X"10",X"FF",X"CD",X"E1",X"F2",X"3E",X"23",X"06",X"20",X"FF",X"DD",X"21",
		X"33",X"F2",X"CD",X"8A",X"5A",X"FD",X"7E",X"00",X"3C",X"06",X"00",X"FE",X"0A",X"38",X"05",X"04",
		X"D6",X"0A",X"18",X"F7",X"4F",X"21",X"56",X"95",X"78",X"B7",X"28",X"10",X"F5",X"C5",X"3E",X"23",
		X"06",X"02",X"FF",X"C1",X"F1",X"C6",X"30",X"77",X"CB",X"DC",X"36",X"07",X"21",X"36",X"95",X"C5",
		X"3E",X"23",X"06",X"02",X"FF",X"C1",X"79",X"C6",X"30",X"77",X"CB",X"DC",X"36",X"07",X"3E",X"23",
		X"06",X"1E",X"FF",X"3A",X"00",X"B0",X"E6",X"03",X"FE",X"03",X"20",X"31",X"3A",X"00",X"B8",X"E6",
		X"0C",X"FE",X"0C",X"20",X"28",X"21",X"20",X"80",X"11",X"D4",X"85",X"3A",X"00",X"80",X"CB",X"6F",
		X"28",X"02",X"13",X"23",X"3A",X"00",X"B8",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",
		X"3F",X"CB",X"3F",X"3C",X"86",X"77",X"EB",X"34",X"FD",X"34",X"00",X"18",X"88",X"3E",X"23",X"06",
		X"1E",X"FF",X"21",X"24",X"C0",X"CB",X"86",X"ED",X"7B",X"08",X"C2",X"C9",X"04",X"05",X"C9",X"92",
		X"9C",X"00",X"00",X"42",X"4F",X"4E",X"55",X"53",X"00",X"00",X"02",X"09",X"92",X"9C",X"00",X"01",
		X"58",X"32",X"00",X"02",X"0A",X"D6",X"92",X"9C",X"00",X"07",X"4E",X"45",X"58",X"54",X"20",X"52",
		X"4F",X"55",X"4E",X"44",X"00",X"01",X"01",X"01",X"17",X"17",X"17",X"02",X"02",X"02",X"18",X"18",
		X"18",X"15",X"15",X"15",X"19",X"19",X"19",X"03",X"03",X"03",X"1A",X"1A",X"1A",X"04",X"04",X"04",
		X"1B",X"1B",X"1B",X"16",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"01",X"05",X"00",X"00",X"01",X"05",X"00",X"00",X"01",X"05",X"00",X"00",X"02",X"00",
		X"00",X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"02",X"05",X"00",X"00",X"02",X"05",
		X"00",X"00",X"02",X"05",X"00",X"00",X"03",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"03",X"00",
		X"00",X"00",X"03",X"05",X"00",X"00",X"03",X"05",X"00",X"00",X"03",X"05",X"00",X"00",X"04",X"00",
		X"00",X"00",X"04",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"04",X"05",X"00",X"00",X"04",X"05",
		X"00",X"00",X"04",X"05",X"00",X"00",X"05",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",X"00",
		X"00",X"00",X"05",X"05",X"00",X"00",X"05",X"05",X"00",X"00",X"05",X"05",X"00",X"00",X"06",X"00",
		X"00",X"CD",X"33",X"F5",X"DD",X"21",X"30",X"C1",X"11",X"14",X"00",X"06",X"09",X"FD",X"CB",X"06",
		X"46",X"28",X"0A",X"CD",X"75",X"F3",X"3E",X"23",X"06",X"01",X"FF",X"18",X"11",X"DD",X"CB",X"00",
		X"46",X"28",X"07",X"C5",X"D5",X"CD",X"D0",X"F3",X"D1",X"C1",X"DD",X"19",X"10",X"DF",X"3E",X"23",
		X"06",X"01",X"FF",X"FD",X"35",X"04",X"C2",X"E4",X"F2",X"FD",X"7E",X"07",X"FD",X"77",X"04",X"FD",
		X"35",X"05",X"20",X"04",X"FD",X"36",X"05",X"03",X"FD",X"7E",X"05",X"C6",X"06",X"21",X"FF",X"9D",
		X"11",X"E0",X"FF",X"06",X"08",X"77",X"2B",X"77",X"23",X"19",X"10",X"F9",X"FD",X"6E",X"02",X"FD",
		X"66",X"03",X"11",X"17",X"C0",X"06",X"05",X"CD",X"8B",X"5B",X"21",X"A9",X"91",X"DD",X"21",X"13",
		X"C0",X"16",X"9C",X"1E",X"07",X"06",X"05",X"0E",X"00",X"CD",X"B9",X"5B",X"FD",X"7E",X"01",X"CD",
		X"5C",X"57",X"21",X"13",X"C0",X"06",X"05",X"AF",X"B6",X"23",X"10",X"FC",X"C2",X"E4",X"F2",X"3E",
		X"00",X"32",X"00",X"A8",X"C9",X"21",X"A5",X"90",X"01",X"16",X"16",X"C5",X"E5",X"7E",X"B7",X"28",
		X"38",X"FE",X"FF",X"20",X"04",X"3E",X"04",X"18",X"1E",X"FE",X"04",X"38",X"1A",X"D6",X"A8",X"38",
		X"28",X"FE",X"03",X"30",X"24",X"5F",X"16",X"00",X"E5",X"21",X"CD",X"F3",X"19",X"CD",X"C6",X"F3",
		X"BE",X"E1",X"30",X"15",X"34",X"18",X"12",X"3D",X"5F",X"16",X"00",X"E5",X"21",X"C9",X"F3",X"19",
		X"CD",X"C6",X"F3",X"BE",X"E1",X"30",X"02",X"36",X"A8",X"23",X"10",X"C1",X"E1",X"C1",X"11",X"20",
		X"00",X"19",X"0D",X"20",X"B6",X"C9",X"ED",X"5F",X"C9",X"40",X"10",X"02",X"01",X"08",X"08",X"08",
		X"CD",X"0F",X"F4",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"2B",X"DD",X"75",X"02",X"DD",X"74",X"03",
		X"7D",X"B4",X"CC",X"38",X"F4",X"DD",X"6E",X"04",X"DD",X"66",X"05",X"2B",X"DD",X"75",X"04",X"DD",
		X"74",X"05",X"7D",X"B4",X"CC",X"CA",X"F4",X"DD",X"7E",X"01",X"6F",X"26",X"00",X"29",X"29",X"11",
		X"08",X"C1",X"19",X"23",X"23",X"DD",X"5E",X"06",X"DD",X"56",X"07",X"73",X"23",X"72",X"C9",X"CD",
		X"1A",X"F4",X"DD",X"23",X"CD",X"1A",X"F4",X"DD",X"2B",X"C9",X"DD",X"7E",X"0A",X"DD",X"86",X"08",
		X"4F",X"E6",X"0F",X"DD",X"77",X"0A",X"B9",X"C8",X"79",X"CB",X"2F",X"CB",X"2F",X"CB",X"2F",X"CB",
		X"2F",X"DD",X"86",X"06",X"DD",X"77",X"06",X"C9",X"DD",X"6E",X"0E",X"DD",X"66",X"0F",X"CB",X"46",
		X"28",X"2E",X"DD",X"6E",X"0C",X"DD",X"66",X"0D",X"CD",X"A5",X"F0",X"7D",X"B4",X"20",X"19",X"DD",
		X"CB",X"00",X"86",X"DD",X"36",X"06",X"00",X"DD",X"36",X"07",X"00",X"DD",X"36",X"08",X"00",X"DD",
		X"36",X"09",X"00",X"DD",X"36",X"02",X"00",X"C9",X"DD",X"73",X"0C",X"DD",X"72",X"0D",X"18",X"CE",
		X"4E",X"23",X"CD",X"A5",X"F0",X"DD",X"75",X"02",X"DD",X"74",X"03",X"CB",X"59",X"28",X"12",X"EB",
		X"CD",X"A5",X"F0",X"DD",X"75",X"08",X"DD",X"74",X"09",X"DD",X"36",X"0A",X"00",X"DD",X"36",X"0B",
		X"00",X"CB",X"51",X"28",X"18",X"EB",X"CD",X"A5",X"F0",X"DD",X"75",X"10",X"DD",X"74",X"11",X"DD",
		X"75",X"12",X"DD",X"74",X"13",X"DD",X"36",X"04",X"01",X"DD",X"36",X"05",X"00",X"CB",X"49",X"28",
		X"12",X"EB",X"CD",X"A5",X"F0",X"DD",X"75",X"06",X"DD",X"74",X"07",X"DD",X"36",X"0A",X"00",X"DD",
		X"36",X"0B",X"00",X"DD",X"73",X"0E",X"DD",X"72",X"0F",X"C9",X"DD",X"6E",X"10",X"DD",X"66",X"11",
		X"CD",X"A5",X"F0",X"7D",X"B4",X"20",X"08",X"DD",X"6E",X"12",X"DD",X"66",X"13",X"18",X"F1",X"DD",
		X"75",X"04",X"DD",X"74",X"05",X"DD",X"6E",X"01",X"26",X"00",X"29",X"29",X"01",X"08",X"C1",X"09",
		X"EB",X"7E",X"ED",X"A0",X"ED",X"A0",X"4F",X"DD",X"7E",X"01",X"FE",X"08",X"28",X"07",X"DD",X"75",
		X"10",X"DD",X"74",X"11",X"C9",X"13",X"13",X"CB",X"61",X"28",X"0C",X"3A",X"00",X"80",X"CB",X"7F",
		X"7E",X"23",X"28",X"03",X"32",X"00",X"A8",X"79",X"E6",X"0F",X"B7",X"28",X"0A",X"CB",X"3F",X"30",
		X"03",X"ED",X"A0",X"1B",X"13",X"18",X"F3",X"DD",X"75",X"10",X"DD",X"74",X"11",X"21",X"28",X"C1",
		X"CB",X"FE",X"C9",X"FD",X"36",X"07",X"08",X"FD",X"36",X"04",X"08",X"FD",X"36",X"05",X"03",X"FD",
		X"7E",X"00",X"3D",X"FE",X"12",X"38",X"04",X"D6",X"12",X"18",X"F8",X"87",X"5F",X"16",X"00",X"21",
		X"AB",X"F6",X"19",X"CD",X"A5",X"F0",X"7E",X"23",X"FE",X"FF",X"C8",X"CB",X"7F",X"28",X"07",X"E5",
		X"CD",X"9C",X"F5",X"E1",X"18",X"F0",X"CD",X"A5",X"F0",X"D5",X"E5",X"6F",X"26",X"00",X"29",X"29",
		X"E5",X"29",X"29",X"D1",X"19",X"11",X"30",X"C1",X"19",X"E5",X"DD",X"E1",X"E1",X"CD",X"A5",X"F0",
		X"DD",X"CB",X"00",X"C6",X"DD",X"77",X"01",X"DD",X"73",X"0C",X"DD",X"72",X"0D",X"DD",X"75",X"0E",
		X"DD",X"74",X"0F",X"CD",X"38",X"F4",X"CD",X"CA",X"F4",X"E1",X"18",X"BA",X"21",X"F3",X"F5",X"CB",
		X"47",X"28",X"1B",X"FD",X"CB",X"06",X"C6",X"FD",X"36",X"07",X"01",X"FD",X"36",X"04",X"01",X"21",
		X"27",X"F6",X"3A",X"00",X"80",X"CB",X"7F",X"28",X"05",X"3E",X"6D",X"32",X"00",X"A8",X"7E",X"23",
		X"B7",X"28",X"18",X"47",X"7E",X"23",X"4E",X"23",X"CD",X"A5",X"F0",X"D5",X"11",X"E0",X"FF",X"77",
		X"CB",X"DC",X"71",X"CB",X"9C",X"19",X"10",X"F7",X"E1",X"18",X"E3",X"7E",X"B7",X"C8",X"47",X"23",
		X"7E",X"23",X"4E",X"23",X"CD",X"A5",X"F0",X"77",X"CB",X"DC",X"71",X"CB",X"9C",X"23",X"10",X"F7",
		X"EB",X"18",X"E8",X"18",X"FD",X"1F",X"6D",X"97",X"18",X"FE",X"1F",X"6E",X"97",X"18",X"FE",X"1F",
		X"6F",X"97",X"18",X"FE",X"1F",X"70",X"97",X"18",X"0C",X"0B",X"72",X"97",X"04",X"00",X"1F",X"6D",
		X"95",X"04",X"00",X"1F",X"6E",X"95",X"04",X"00",X"1F",X"6F",X"95",X"04",X"00",X"1F",X"70",X"95",
		X"04",X"00",X"0B",X"92",X"95",X"00",X"00",X"16",X"FF",X"1D",X"4E",X"97",X"16",X"FF",X"1D",X"51",
		X"97",X"16",X"03",X"1D",X"45",X"97",X"16",X"03",X"1D",X"4D",X"97",X"16",X"03",X"1D",X"52",X"97",
		X"16",X"03",X"1D",X"5A",X"97",X"14",X"02",X"1D",X"26",X"97",X"14",X"02",X"1D",X"2C",X"97",X"14",
		X"02",X"1D",X"33",X"97",X"14",X"02",X"1D",X"39",X"97",X"12",X"01",X"1D",X"07",X"97",X"12",X"01",
		X"1D",X"0B",X"97",X"12",X"01",X"1D",X"14",X"97",X"12",X"01",X"1D",X"18",X"97",X"00",X"07",X"03",
		X"1D",X"46",X"97",X"07",X"03",X"1D",X"A6",X"94",X"07",X"03",X"1D",X"53",X"97",X"07",X"03",X"1D",
		X"B3",X"94",X"05",X"02",X"1D",X"27",X"97",X"05",X"02",X"1D",X"C7",X"94",X"05",X"02",X"1D",X"34",
		X"97",X"05",X"02",X"1D",X"D4",X"94",X"03",X"01",X"1D",X"08",X"97",X"03",X"01",X"1D",X"E8",X"94",
		X"03",X"01",X"1D",X"15",X"97",X"03",X"01",X"1D",X"F5",X"94",X"00",X"31",X"F7",X"31",X"F7",X"CF",
		X"F6",X"31",X"F7",X"31",X"F7",X"E9",X"F6",X"31",X"F7",X"31",X"F7",X"ED",X"F6",X"31",X"F7",X"31",
		X"F7",X"07",X"F7",X"31",X"F7",X"31",X"F7",X"17",X"F7",X"31",X"F7",X"31",X"F7",X"27",X"F7",X"06",
		X"47",X"F7",X"05",X"43",X"F7",X"04",X"3F",X"F7",X"03",X"3B",X"F7",X"02",X"37",X"F7",X"01",X"33",
		X"F7",X"00",X"4B",X"F7",X"08",X"4F",X"F7",X"80",X"FF",X"08",X"65",X"F7",X"FF",X"06",X"8D",X"F7",
		X"05",X"89",X"F7",X"04",X"85",X"F7",X"03",X"81",X"F7",X"02",X"7D",X"F7",X"01",X"69",X"F7",X"00",
		X"91",X"F7",X"08",X"95",X"F7",X"80",X"FF",X"00",X"99",X"F7",X"01",X"9D",X"F7",X"02",X"A1",X"F7",
		X"03",X"A5",X"F7",X"08",X"A9",X"F7",X"FF",X"00",X"AD",X"F7",X"01",X"B1",X"F7",X"02",X"B5",X"F7",
		X"03",X"B9",X"F7",X"08",X"BD",X"F7",X"FF",X"00",X"C1",X"F7",X"01",X"C5",X"F7",X"08",X"C9",X"F7",
		X"FF",X"81",X"FF",X"CD",X"F7",X"00",X"00",X"A3",X"F8",X"00",X"00",X"09",X"F9",X"00",X"00",X"6F",
		X"F9",X"00",X"00",X"D5",X"F9",X"00",X"00",X"3B",X"FA",X"00",X"00",X"A1",X"FA",X"00",X"00",X"BB",
		X"FA",X"FC",X"FA",X"FC",X"FA",X"FC",X"FA",X"FC",X"FA",X"FC",X"FA",X"FC",X"FA",X"FC",X"FA",X"FC",
		X"FA",X"09",X"FB",X"00",X"00",X"E9",X"FB",X"00",X"00",X"6D",X"FD",X"AC",X"FD",X"AC",X"FD",X"AC",
		X"FD",X"AC",X"FD",X"AC",X"FD",X"AC",X"FD",X"AC",X"FD",X"AC",X"FD",X"00",X"00",X"C9",X"FD",X"00",
		X"00",X"DF",X"FD",X"00",X"00",X"F5",X"FD",X"00",X"00",X"0B",X"FE",X"00",X"00",X"21",X"FE",X"00",
		X"00",X"37",X"FE",X"00",X"00",X"55",X"FE",X"00",X"00",X"6E",X"FC",X"00",X"00",X"78",X"FC",X"00",
		X"00",X"82",X"FC",X"00",X"00",X"8C",X"FC",X"00",X"00",X"BE",X"FC",X"00",X"00",X"0F",X"FD",X"00",
		X"00",X"19",X"FD",X"00",X"00",X"23",X"FD",X"00",X"00",X"2D",X"FD",X"00",X"00",X"4F",X"FD",X"00",
		X"00",X"57",X"FF",X"00",X"00",X"7D",X"FF",X"00",X"00",X"A8",X"FF",X"00",X"00",X"0E",X"66",X"00",
		X"18",X"00",X"51",X"F8",X"00",X"80",X"0C",X"20",X"00",X"00",X"00",X"1B",X"F8",X"0C",X"20",X"00",
		X"F0",X"00",X"43",X"F8",X"0C",X"18",X"00",X"00",X"00",X"1B",X"F8",X"0C",X"50",X"00",X"18",X"00",
		X"51",X"F8",X"08",X"A2",X"00",X"00",X"00",X"0E",X"14",X"00",X"10",X"00",X"43",X"F8",X"00",X"80",
		X"0C",X"14",X"00",X"F0",X"00",X"87",X"F8",X"08",X"10",X"00",X"00",X"00",X"0C",X"48",X"00",X"10",
		X"00",X"43",X"F8",X"0C",X"FF",X"FF",X"00",X"00",X"1B",X"F8",X"01",X"01",X"00",X"97",X"10",X"00",
		X"00",X"01",X"00",X"97",X"11",X"00",X"00",X"20",X"00",X"96",X"11",X"20",X"00",X"97",X"11",X"20",
		X"00",X"98",X"11",X"00",X"00",X"10",X"00",X"96",X"11",X"10",X"00",X"97",X"11",X"10",X"00",X"98",
		X"11",X"00",X"00",X"08",X"00",X"96",X"10",X"08",X"00",X"97",X"10",X"08",X"00",X"98",X"10",X"00",
		X"00",X"04",X"00",X"96",X"10",X"04",X"00",X"97",X"10",X"04",X"00",X"98",X"10",X"00",X"00",X"01",
		X"00",X"17",X"10",X"00",X"00",X"01",X"00",X"17",X"11",X"00",X"00",X"20",X"00",X"16",X"11",X"20",
		X"00",X"17",X"11",X"20",X"00",X"18",X"11",X"00",X"00",X"10",X"00",X"16",X"11",X"10",X"00",X"17",
		X"11",X"10",X"00",X"18",X"11",X"00",X"00",X"08",X"00",X"16",X"10",X"08",X"00",X"17",X"10",X"08",
		X"00",X"18",X"10",X"00",X"00",X"04",X"00",X"16",X"10",X"04",X"00",X"17",X"10",X"04",X"00",X"18",
		X"10",X"00",X"00",X"0E",X"0E",X"00",X"00",X"00",X"E7",X"F8",X"00",X"80",X"08",X"58",X"00",X"18",
		X"00",X"0C",X"20",X"00",X"00",X"00",X"D3",X"F8",X"0C",X"20",X"00",X"F0",X"00",X"D9",X"F8",X"0C",
		X"52",X"00",X"00",X"00",X"D3",X"F8",X"04",X"08",X"00",X"F5",X"F8",X"0C",X"64",X"00",X"F0",X"00",
		X"FB",X"F8",X"01",X"01",X"00",X"2F",X"12",X"00",X"00",X"08",X"00",X"2E",X"12",X"08",X"00",X"2F",
		X"12",X"08",X"00",X"30",X"12",X"00",X"00",X"04",X"00",X"2E",X"12",X"04",X"00",X"2F",X"12",X"04",
		X"00",X"30",X"12",X"00",X"00",X"01",X"00",X"AF",X"12",X"00",X"00",X"08",X"00",X"AE",X"12",X"08",
		X"00",X"AF",X"12",X"08",X"00",X"B0",X"12",X"00",X"00",X"0E",X"1C",X"00",X"00",X"00",X"4D",X"F9",
		X"00",X"80",X"08",X"4A",X"00",X"18",X"00",X"0C",X"20",X"00",X"00",X"00",X"39",X"F9",X"0C",X"20",
		X"00",X"F0",X"00",X"3F",X"F9",X"0C",X"52",X"00",X"00",X"00",X"39",X"F9",X"04",X"08",X"00",X"5B",
		X"F9",X"0C",X"4F",X"00",X"F0",X"00",X"61",X"F9",X"01",X"01",X"00",X"2F",X"13",X"00",X"00",X"08",
		X"00",X"2E",X"13",X"08",X"00",X"2F",X"13",X"08",X"00",X"30",X"13",X"00",X"00",X"04",X"00",X"2E",
		X"13",X"04",X"00",X"2F",X"13",X"04",X"00",X"30",X"13",X"00",X"00",X"01",X"00",X"AF",X"13",X"00",
		X"00",X"08",X"00",X"AE",X"13",X"08",X"00",X"AF",X"13",X"08",X"00",X"B0",X"13",X"00",X"00",X"0E",
		X"2A",X"00",X"00",X"00",X"B3",X"F9",X"00",X"80",X"08",X"3C",X"00",X"18",X"00",X"0C",X"20",X"00",
		X"00",X"00",X"9F",X"F9",X"0C",X"20",X"00",X"F0",X"00",X"A5",X"F9",X"0C",X"52",X"00",X"00",X"00",
		X"9F",X"F9",X"04",X"08",X"00",X"C1",X"F9",X"0C",X"3A",X"00",X"F0",X"00",X"C7",X"F9",X"01",X"01",
		X"00",X"2F",X"14",X"00",X"00",X"08",X"00",X"2E",X"14",X"08",X"00",X"2F",X"14",X"08",X"00",X"30",
		X"14",X"00",X"00",X"04",X"00",X"2E",X"14",X"04",X"00",X"2F",X"14",X"04",X"00",X"30",X"14",X"00",
		X"00",X"01",X"00",X"AF",X"14",X"00",X"00",X"08",X"00",X"AE",X"14",X"08",X"00",X"AF",X"14",X"08",
		X"00",X"B0",X"14",X"00",X"00",X"0E",X"38",X"00",X"00",X"00",X"19",X"FA",X"00",X"80",X"08",X"2E",
		X"00",X"18",X"00",X"0C",X"20",X"00",X"00",X"00",X"05",X"FA",X"0C",X"20",X"00",X"F0",X"00",X"0B",
		X"FA",X"0C",X"52",X"00",X"00",X"00",X"05",X"FA",X"04",X"08",X"00",X"27",X"FA",X"0C",X"25",X"00",
		X"F0",X"00",X"2D",X"FA",X"01",X"01",X"00",X"2F",X"15",X"00",X"00",X"08",X"00",X"2E",X"15",X"08",
		X"00",X"2F",X"15",X"08",X"00",X"30",X"15",X"00",X"00",X"04",X"00",X"2E",X"15",X"04",X"00",X"2F",
		X"15",X"04",X"00",X"30",X"15",X"00",X"00",X"01",X"00",X"AF",X"15",X"00",X"00",X"08",X"00",X"AE",
		X"15",X"08",X"00",X"AF",X"15",X"08",X"00",X"B0",X"15",X"00",X"00",X"0E",X"46",X"00",X"00",X"00",
		X"7F",X"FA",X"00",X"80",X"08",X"20",X"00",X"18",X"00",X"0C",X"20",X"00",X"00",X"00",X"6B",X"FA",
		X"0C",X"20",X"00",X"F0",X"00",X"71",X"FA",X"0C",X"52",X"00",X"00",X"00",X"6B",X"FA",X"04",X"08",
		X"00",X"8D",X"FA",X"0C",X"10",X"00",X"F0",X"00",X"93",X"FA",X"01",X"01",X"00",X"34",X"16",X"00",
		X"00",X"08",X"00",X"33",X"16",X"08",X"00",X"34",X"16",X"08",X"00",X"35",X"16",X"00",X"00",X"04",
		X"00",X"33",X"16",X"04",X"00",X"34",X"16",X"04",X"00",X"35",X"16",X"00",X"00",X"01",X"00",X"B4",
		X"16",X"00",X"00",X"08",X"00",X"B3",X"16",X"08",X"00",X"B4",X"16",X"08",X"00",X"B5",X"16",X"00",
		X"00",X"0E",X"05",X"00",X"00",X"00",X"B5",X"FA",X"10",X"80",X"08",X"30",X"00",X"18",X"00",X"08",
		X"FF",X"FF",X"00",X"00",X"01",X"01",X"00",X"2C",X"19",X"00",X"00",X"0E",X"F0",X"00",X"00",X"00",
		X"11",X"FB",X"90",X"60",X"02",X"40",X"00",X"90",X"70",X"02",X"10",X"00",X"8C",X"70",X"02",X"20",
		X"00",X"87",X"70",X"02",X"10",X"00",X"83",X"70",X"02",X"20",X"00",X"7E",X"70",X"02",X"40",X"00",
		X"7A",X"70",X"02",X"20",X"00",X"75",X"70",X"02",X"10",X"00",X"71",X"70",X"02",X"20",X"00",X"6C",
		X"70",X"02",X"10",X"00",X"68",X"70",X"02",X"20",X"00",X"63",X"70",X"01",X"06",X"20",X"00",X"CB",
		X"FB",X"63",X"68",X"02",X"20",X"00",X"63",X"70",X"01",X"06",X"FF",X"FF",X"DF",X"FB",X"63",X"68",
		X"01",X"70",X"00",X"1F",X"0B",X"60",X"04",X"14",X"24",X"34",X"10",X"00",X"1F",X"0B",X"63",X"C4",
		X"D4",X"E4",X"F4",X"48",X"00",X"1F",X"0B",X"63",X"04",X"14",X"24",X"34",X"28",X"00",X"1F",X"0B",
		X"63",X"C4",X"D4",X"E4",X"F4",X"10",X"00",X"1F",X"0A",X"64",X"CC",X"DC",X"EC",X"FC",X"30",X"00",
		X"1F",X"0A",X"63",X"08",X"18",X"28",X"38",X"10",X"00",X"1F",X"0A",X"61",X"0C",X"1C",X"2C",X"3C",
		X"20",X"00",X"1F",X"0A",X"61",X"08",X"18",X"28",X"38",X"10",X"00",X"1F",X"0A",X"61",X"0C",X"1C",
		X"2C",X"3C",X"20",X"00",X"1F",X"0A",X"61",X"08",X"18",X"28",X"38",X"08",X"00",X"1F",X"0A",X"61",
		X"0C",X"1C",X"2C",X"3C",X"08",X"00",X"13",X"0A",X"63",X"C8",X"D8",X"10",X"00",X"13",X"0A",X"63",
		X"0C",X"1C",X"20",X"00",X"13",X"0A",X"63",X"C8",X"D8",X"20",X"00",X"1F",X"0A",X"61",X"CC",X"DC",
		X"EC",X"FC",X"01",X"00",X"1F",X"0A",X"61",X"0C",X"1C",X"2C",X"3C",X"0F",X"00",X"10",X"0A",X"63",
		X"01",X"00",X"1F",X"0A",X"61",X"CC",X"DC",X"EC",X"FC",X"1F",X"00",X"10",X"0A",X"63",X"10",X"00",
		X"1F",X"0A",X"61",X"C8",X"D8",X"2C",X"3C",X"10",X"00",X"1F",X"0A",X"61",X"CC",X"DC",X"EC",X"FC",
		X"10",X"00",X"1F",X"0A",X"63",X"08",X"18",X"28",X"38",X"00",X"00",X"20",X"00",X"1F",X"0A",X"62",
		X"40",X"50",X"60",X"70",X"20",X"00",X"1F",X"0A",X"64",X"C0",X"D0",X"E0",X"F0",X"00",X"00",X"FF",
		X"FF",X"0F",X"0A",X"40",X"50",X"60",X"70",X"00",X"00",X"0E",X"C0",X"02",X"00",X"00",X"F8",X"FB",
		X"70",X"70",X"04",X"FF",X"FF",X"5B",X"FC",X"01",X"40",X"00",X"1F",X"0A",X"65",X"44",X"54",X"64",
		X"74",X"40",X"00",X"1F",X"0A",X"66",X"4C",X"5C",X"6C",X"7C",X"40",X"00",X"08",X"0A",X"B0",X"40",
		X"00",X"0F",X"0A",X"44",X"54",X"64",X"78",X"40",X"00",X"1F",X"0A",X"66",X"4C",X"5C",X"6C",X"B0",
		X"40",X"00",X"04",X"0A",X"A0",X"40",X"00",X"0F",X"0A",X"44",X"54",X"68",X"78",X"40",X"00",X"1F",
		X"0A",X"66",X"4C",X"5C",X"A0",X"B0",X"40",X"00",X"02",X"0A",X"90",X"40",X"00",X"0F",X"0A",X"44",
		X"58",X"68",X"78",X"40",X"00",X"1F",X"0A",X"66",X"4C",X"90",X"A0",X"B0",X"40",X"00",X"01",X"0A",
		X"80",X"40",X"00",X"0F",X"0A",X"48",X"58",X"68",X"78",X"00",X"00",X"40",X"00",X"1F",X"0A",X"66",
		X"80",X"90",X"A0",X"B0",X"40",X"00",X"0F",X"0A",X"48",X"58",X"68",X"78",X"00",X"00",X"0E",X"FF",
		X"FF",X"00",X"00",X"96",X"FC",X"60",X"80",X"01",X"0E",X"FF",X"FF",X"00",X"00",X"A0",X"FC",X"88",
		X"94",X"01",X"0E",X"FF",X"FF",X"00",X"00",X"AA",X"FC",X"94",X"7C",X"01",X"0E",X"FF",X"FF",X"00",
		X"00",X"B4",X"FC",X"70",X"98",X"01",X"D0",X"00",X"00",X"00",X"FF",X"FF",X"2C",X"19",X"00",X"00",
		X"90",X"01",X"00",X"00",X"FF",X"FF",X"2C",X"19",X"00",X"00",X"50",X"02",X"00",X"00",X"FF",X"FF",
		X"2C",X"19",X"00",X"00",X"10",X"03",X"00",X"00",X"FF",X"FF",X"2C",X"19",X"00",X"00",X"0E",X"40",
		X"00",X"00",X"00",X"CD",X"FC",X"70",X"70",X"04",X"FF",X"FF",X"D8",X"FC",X"01",X"40",X"00",X"1F",
		X"0A",X"65",X"44",X"54",X"64",X"74",X"00",X"00",X"20",X"00",X"1F",X"0A",X"69",X"4C",X"5C",X"6C",
		X"7C",X"20",X"00",X"08",X"0A",X"B0",X"20",X"00",X"04",X"0A",X"A0",X"20",X"00",X"02",X"0A",X"90",
		X"20",X"00",X"1F",X"0A",X"6A",X"48",X"58",X"68",X"78",X"08",X"00",X"01",X"0A",X"44",X"08",X"00",
		X"02",X"0A",X"54",X"08",X"00",X"04",X"0A",X"64",X"08",X"00",X"08",X"0A",X"74",X"00",X"00",X"0E",
		X"FF",X"FF",X"00",X"00",X"37",X"FD",X"60",X"80",X"01",X"0E",X"FF",X"FF",X"00",X"00",X"3D",X"FD",
		X"88",X"94",X"01",X"0E",X"FF",X"FF",X"00",X"00",X"43",X"FD",X"94",X"7C",X"01",X"0E",X"FF",X"FF",
		X"00",X"00",X"49",X"FD",X"70",X"98",X"01",X"FF",X"FF",X"2C",X"19",X"00",X"00",X"FF",X"FF",X"2C",
		X"19",X"00",X"00",X"FF",X"FF",X"2C",X"19",X"00",X"00",X"FF",X"FF",X"2C",X"19",X"00",X"00",X"0E",
		X"FF",X"FF",X"00",X"00",X"59",X"FD",X"70",X"70",X"01",X"40",X"00",X"1F",X"0A",X"6E",X"88",X"98",
		X"A8",X"B8",X"40",X"00",X"1F",X"0A",X"6F",X"8C",X"9C",X"AC",X"BC",X"00",X"00",X"0E",X"80",X"00",
		X"F0",X"00",X"87",X"F8",X"F0",X"80",X"0C",X"38",X"00",X"00",X"00",X"5F",X"F8",X"04",X"18",X"00",
		X"1B",X"F8",X"04",X"10",X"00",X"5F",X"F8",X"0C",X"20",X"00",X"F0",X"00",X"87",X"F8",X"0C",X"18",
		X"00",X"00",X"00",X"5F",X"F8",X"04",X"18",X"00",X"1B",X"F8",X"04",X"10",X"00",X"5F",X"F8",X"0C",
		X"50",X"00",X"F0",X"00",X"87",X"F8",X"08",X"50",X"00",X"00",X"00",X"01",X"0E",X"30",X"00",X"18",
		X"00",X"51",X"F8",X"00",X"80",X"0C",X"08",X"00",X"00",X"00",X"1B",X"F8",X"0C",X"30",X"00",X"E8",
		X"00",X"95",X"F8",X"08",X"08",X"00",X"00",X"00",X"01",X"0E",X"0E",X"00",X"00",X"00",X"D9",X"F8",
		X"00",X"80",X"08",X"58",X"00",X"10",X"00",X"0C",X"58",X"00",X"F0",X"00",X"FB",X"F8",X"01",X"0E",
		X"22",X"00",X"00",X"00",X"3F",X"F9",X"00",X"80",X"08",X"58",X"00",X"10",X"00",X"0C",X"58",X"00",
		X"F0",X"00",X"61",X"F9",X"01",X"0E",X"36",X"00",X"00",X"00",X"A5",X"F9",X"00",X"80",X"08",X"58",
		X"00",X"10",X"00",X"0C",X"58",X"00",X"F0",X"00",X"C7",X"F9",X"01",X"0E",X"4A",X"00",X"00",X"00",
		X"0B",X"FA",X"00",X"80",X"08",X"58",X"00",X"10",X"00",X"0C",X"58",X"00",X"F0",X"00",X"2D",X"FA",
		X"01",X"0E",X"5E",X"00",X"00",X"00",X"71",X"FA",X"00",X"80",X"08",X"58",X"00",X"10",X"00",X"0C",
		X"58",X"00",X"F0",X"00",X"93",X"FA",X"01",X"0E",X"08",X"00",X"00",X"00",X"B5",X"FA",X"E0",X"80",
		X"08",X"78",X"00",X"F0",X"00",X"08",X"60",X"00",X"00",X"00",X"08",X"10",X"00",X"F0",X"00",X"08",
		X"FF",X"FF",X"00",X"00",X"01",X"0E",X"80",X"00",X"00",X"00",X"9B",X"FE",X"90",X"60",X"02",X"20",
		X"00",X"90",X"70",X"02",X"10",X"00",X"8C",X"70",X"02",X"50",X"00",X"87",X"70",X"02",X"10",X"00",
		X"83",X"70",X"02",X"50",X"00",X"7E",X"70",X"02",X"10",X"00",X"7A",X"70",X"02",X"20",X"00",X"75",
		X"70",X"02",X"10",X"00",X"71",X"70",X"02",X"20",X"00",X"6C",X"70",X"02",X"10",X"00",X"68",X"70",
		X"02",X"10",X"00",X"63",X"70",X"04",X"FF",X"FF",X"32",X"FF",X"01",X"40",X"00",X"1F",X"0B",X"67",
		X"C4",X"D4",X"24",X"34",X"40",X"00",X"13",X"0B",X"63",X"04",X"14",X"20",X"00",X"1F",X"0A",X"64",
		X"08",X"18",X"28",X"38",X"10",X"00",X"1F",X"0A",X"61",X"0C",X"1C",X"2C",X"3C",X"10",X"00",X"1F",
		X"0A",X"61",X"08",X"18",X"28",X"38",X"20",X"00",X"1F",X"0A",X"68",X"84",X"94",X"A4",X"B4",X"20",
		X"00",X"0F",X"0A",X"08",X"18",X"28",X"38",X"10",X"00",X"1F",X"0A",X"61",X"0C",X"1C",X"2C",X"3C",
		X"20",X"00",X"1F",X"0A",X"61",X"08",X"18",X"28",X"38",X"10",X"00",X"1F",X"0A",X"68",X"84",X"94",
		X"A4",X"B4",X"20",X"00",X"0F",X"0A",X"08",X"18",X"28",X"38",X"10",X"00",X"1F",X"0A",X"61",X"0C",
		X"1C",X"2C",X"3C",X"20",X"00",X"1F",X"0A",X"61",X"08",X"18",X"28",X"38",X"10",X"00",X"1F",X"0A",
		X"61",X"0C",X"1C",X"2C",X"3C",X"20",X"00",X"1F",X"0A",X"61",X"08",X"18",X"28",X"38",X"10",X"00",
		X"1F",X"0A",X"61",X"C8",X"D8",X"2C",X"3C",X"10",X"00",X"1F",X"0A",X"61",X"08",X"18",X"28",X"38",
		X"00",X"00",X"10",X"00",X"1F",X"0A",X"63",X"CC",X"DC",X"EC",X"FC",X"08",X"00",X"1F",X"0A",X"63",
		X"08",X"18",X"28",X"38",X"30",X"00",X"1F",X"0A",X"68",X"84",X"94",X"A4",X"B4",X"28",X"00",X"0F",
		X"0A",X"08",X"18",X"28",X"38",X"00",X"00",X"0E",X"64",X"00",X"10",X"00",X"43",X"F8",X"00",X"80",
		X"0C",X"20",X"00",X"00",X"00",X"21",X"F8",X"0C",X"30",X"00",X"04",X"00",X"27",X"F8",X"0C",X"20",
		X"00",X"00",X"00",X"21",X"F8",X"0C",X"00",X"01",X"08",X"00",X"35",X"F8",X"01",X"0E",X"64",X"00",
		X"F0",X"00",X"87",X"F8",X"F0",X"80",X"0C",X"20",X"00",X"00",X"00",X"65",X"F8",X"0C",X"30",X"00",
		X"FC",X"00",X"6B",X"F8",X"0C",X"1A",X"00",X"00",X"00",X"65",X"F8",X"04",X"06",X"00",X"21",X"F8",
		X"0C",X"00",X"01",X"08",X"00",X"35",X"F8",X"01",X"0E",X"64",X"00",X"00",X"00",X"59",X"FD",X"70",
		X"70",X"02",X"6A",X"00",X"70",X"62",X"02",X"06",X"00",X"70",X"66",X"08",X"00",X"01",X"08",X"00",
		X"04",X"01",X"00",X"C6",X"FF",X"01",X"01",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"20",X"20",X"20",X"20",X"47",X"55",X"5A",X"5A",X"4C",X"45",X"52",X"20",X"20",X"20",X"20",
		X"20",X"31",X"39",X"38",X"33",X"20",X"43",X"6F",X"70",X"79",X"72",X"69",X"67",X"68",X"74",X"20",
		X"20",X"20",X"20",X"54",X"45",X"48",X"4B",X"41",X"4E",X"20",X"4C",X"54",X"44",X"2E",X"20",X"20");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
