library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity kick_sp_bits is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of kick_sp_bits is
	type rom is array(0 to  32767) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"E0",X"00",X"EE",X"00",X"0E",X"00",X"EE",X"00",X"00",X"00",
		X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"0E",X"00",X"00",X"0E",X"E0",X"00",X"00",
		X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"E0",X"00",X"00",X"00",X"0E",X"10",X"00",X"00",X"00",
		X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"11",X"00",X"00",X"0E",X"11",X"00",X"00",X"EE",
		X"11",X"00",X"00",X"E0",X"11",X"E0",X"00",X"00",X"11",X"EE",X"00",X"00",X"11",X"0E",X"EE",X"00",
		X"10",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",
		X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",
		X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",
		X"70",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"70",X"00",X"EE",X"00",
		X"00",X"0E",X"EE",X"00",X"00",X"EE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"E0",
		X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"0E",X"00",X"00",X"E0",X"0E",X"00",X"00",X"00",
		X"0E",X"E0",X"00",X"00",X"EE",X"0E",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",
		X"EE",X"00",X"00",X"00",X"EE",X"00",X"0E",X"00",X"EE",X"EE",X"E0",X"00",X"EE",X"EE",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"0E",X"EE",X"00",X"00",X"EE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"E0",
		X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"7E",X"00",X"00",X"E0",X"77",X"D0",X"88",X"00",
		X"77",X"D0",X"88",X"00",X"77",X"DE",X"88",X"00",X"77",X"D0",X"88",X"00",X"77",X"00",X"88",X"00",
		X"77",X"00",X"88",X"00",X"75",X"00",X"8E",X"00",X"77",X"2E",X"E8",X"00",X"77",X"2E",X"EE",X"EE",
		X"FF",X"33",X"77",X"77",X"FF",X"43",X"77",X"77",X"55",X"44",X"77",X"77",X"55",X"44",X"77",X"77",
		X"05",X"44",X"77",X"77",X"00",X"44",X"77",X"77",X"00",X"44",X"77",X"77",X"00",X"44",X"07",X"77",
		X"00",X"04",X"00",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"33",X"77",X"77",X"55",X"33",X"77",X"77",X"55",X"33",X"77",X"72",X"FF",X"33",X"77",X"72",
		X"55",X"33",X"77",X"72",X"55",X"33",X"77",X"22",X"05",X"00",X"77",X"22",X"00",X"00",X"07",X"22",
		X"00",X"40",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"55",X"00",X"00",X"44",X"FF",X"00",
		X"00",X"44",X"55",X"00",X"00",X"44",X"55",X"B0",X"00",X"44",X"FF",X"00",X"00",X"44",X"55",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"33",X"77",X"77",X"55",X"33",X"77",X"77",X"FF",X"33",X"B7",X"77",X"55",X"33",X"BB",X"77",
		X"55",X"33",X"BB",X"77",X"05",X"43",X"BB",X"22",X"00",X"43",X"BB",X"22",X"00",X"44",X"07",X"22",
		X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"BB",
		X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"44",X"BB",X"00",X"00",X"44",X"BB",
		X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AB",X"00",X"00",X"00",X"AB",X"00",X"00",X"00",X"AA",
		X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"B7",X"00",X"00",X"00",X"BB",
		X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"B6",X"00",X"00",X"44",X"66",X"00",X"00",X"44",X"BB",
		X"00",X"00",X"00",X"BA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",
		X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",
		X"00",X"00",X"00",X"B6",X"00",X"00",X"00",X"B6",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",
		X"00",X"00",X"00",X"AA",X"00",X"00",X"44",X"AB",X"00",X"00",X"44",X"AB",X"00",X"00",X"00",X"AA",
		X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",
		X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"40",X"00",X"01",X"11",
		X"40",X"00",X"07",X"11",X"44",X"00",X"77",X"77",X"44",X"00",X"77",X"77",X"44",X"05",X"77",X"77",
		X"44",X"33",X"77",X"77",X"44",X"33",X"77",X"77",X"44",X"33",X"77",X"77",X"05",X"33",X"77",X"77",
		X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",
		X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"77",X"00",X"00",X"DD",X"77",X"00",X"00",X"DD",X"77",
		X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",
		X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",
		X"00",X"B0",X"00",X"77",X"00",X"B0",X"00",X"77",X"00",X"B0",X"00",X"77",X"00",X"B0",X"00",X"77",
		X"00",X"B0",X"00",X"77",X"00",X"BB",X"00",X"77",X"00",X"0B",X"00",X"77",X"00",X"0B",X"00",X"77",
		X"00",X"BB",X"00",X"77",X"00",X"BB",X"00",X"77",X"00",X"BB",X"00",X"77",X"00",X"BB",X"00",X"77",
		X"00",X"BB",X"00",X"77",X"00",X"FF",X"00",X"77",X"00",X"FF",X"00",X"77",X"00",X"FF",X"00",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"E0",X"00",X"EE",X"00",X"0E",X"00",X"EE",X"00",X"00",X"00",
		X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"0E",X"00",X"00",X"0E",X"E0",X"00",X"00",
		X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"E0",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"EE",
		X"00",X"00",X"00",X"E0",X"00",X"E0",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"0E",X"EE",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"5F",X"22",X"E0",X"00",X"5F",X"22",X"0E",X"00",X"05",X"77",X"00",X"00",X"EE",X"77",X"00",X"00",
		X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"0E",X"00",X"00",X"0E",X"E0",X"00",X"00",
		X"0E",X"00",X"00",X"E0",X"0E",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"EE",
		X"00",X"00",X"00",X"EE",X"00",X"E0",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"0E",X"EE",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"EE",X"EE",X"EE",X"77",X"EE",X"0E",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",
		X"77",X"0E",X"00",X"00",X"EE",X"E0",X"00",X"00",X"EE",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",
		X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",
		X"00",X"00",X"00",X"EE",X"00",X"E0",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"0E",X"EE",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",
		X"00",X"0B",X"00",X"77",X"00",X"BB",X"00",X"77",X"00",X"BB",X"00",X"77",X"00",X"BB",X"00",X"77",
		X"00",X"BB",X"00",X"77",X"00",X"05",X"00",X"77",X"00",X"0F",X"00",X"77",X"00",X"04",X"00",X"70",
		X"00",X"04",X"00",X"70",X"05",X"34",X"00",X"70",X"05",X"33",X"77",X"77",X"55",X"33",X"77",X"77",
		X"FF",X"33",X"77",X"77",X"55",X"33",X"77",X"77",X"55",X"34",X"77",X"77",X"FF",X"44",X"77",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"B5",X"00",X"00",X"00",X"5F",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"F5",X"00",
		X"00",X"00",X"45",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"40",X"01",X"00",X"00",X"07",X"71",
		X"00",X"00",X"77",X"71",X"05",X"00",X"77",X"71",X"05",X"33",X"77",X"77",X"55",X"33",X"77",X"77",
		X"FF",X"33",X"77",X"77",X"55",X"33",X"77",X"77",X"55",X"33",X"77",X"77",X"CF",X"33",X"77",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"11",
		X"00",X"0B",X"00",X"11",X"00",X"BB",X"00",X"11",X"00",X"BB",X"00",X"11",X"00",X"BB",X"00",X"11",
		X"00",X"BF",X"00",X"11",X"00",X"5F",X"00",X"11",X"00",X"F5",X"00",X"11",X"00",X"54",X"00",X"11",
		X"00",X"04",X"00",X"11",X"00",X"04",X"00",X"11",X"00",X"00",X"07",X"11",X"00",X"00",X"07",X"71",
		X"00",X"00",X"77",X"77",X"05",X"03",X"77",X"77",X"05",X"33",X"77",X"77",X"55",X"33",X"77",X"77",
		X"FF",X"33",X"77",X"77",X"55",X"33",X"77",X"77",X"55",X"33",X"77",X"77",X"CF",X"33",X"77",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"0B",X"00",X"00",
		X"00",X"05",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"07",X"00",X"04",X"00",X"07",X"00",X"04",X"00",X"77",X"00",X"44",X"07",X"77",
		X"00",X"33",X"77",X"77",X"05",X"33",X"77",X"77",X"05",X"33",X"77",X"77",X"55",X"33",X"77",X"77",
		X"FF",X"33",X"77",X"77",X"FF",X"33",X"77",X"77",X"55",X"33",X"77",X"77",X"55",X"33",X"77",X"77",
		X"00",X"00",X"00",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",
		X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"D0",
		X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"5B",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"F5",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"4F",X"00",X"00",X"00",X"4F",X"00",
		X"00",X"00",X"40",X"00",X"00",X"44",X"00",X"07",X"00",X"44",X"00",X"77",X"00",X"44",X"00",X"77",
		X"00",X"44",X"00",X"77",X"05",X"44",X"00",X"77",X"55",X"44",X"00",X"77",X"FF",X"44",X"00",X"77",
		X"55",X"40",X"07",X"77",X"55",X"33",X"F7",X"77",X"FF",X"33",X"F7",X"77",X"55",X"33",X"F7",X"77",
		X"55",X"33",X"F7",X"77",X"FF",X"33",X"F7",X"77",X"55",X"33",X"F7",X"77",X"55",X"40",X"07",X"77",
		X"FF",X"44",X"00",X"11",X"55",X"44",X"00",X"11",X"05",X"44",X"00",X"11",X"00",X"44",X"00",X"11",
		X"00",X"44",X"00",X"11",X"00",X"44",X"00",X"01",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"00",
		X"BB",X"FF",X"00",X"00",X"00",X"55",X"00",X"11",X"00",X"FF",X"00",X"11",X"00",X"55",X"00",X"11",
		X"00",X"55",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"05",X"00",X"00",X"00",X"55",X"DD",X"00",X"00",X"DB",X"DD",X"00",X"00",X"DB",X"DD",
		X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",
		X"77",X"77",X"5B",X"00",X"77",X"77",X"FB",X"00",X"77",X"77",X"50",X"00",X"77",X"EE",X"E0",X"EE",
		X"7E",X"E0",X"0E",X"00",X"EE",X"00",X"0E",X"00",X"EE",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",
		X"0E",X"0E",X"00",X"00",X"0E",X"0E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",
		X"00",X"00",X"00",X"EE",X"00",X"E0",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"0E",X"EE",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"FB",X"D0",X"00",X"EE",X"FB",X"E0",X"00",X"EE",X"00",X"0E",X"00",X"EE",X"0D",X"00",X"00",
		X"EE",X"0D",X"00",X"00",X"EE",X"0D",X"00",X"00",X"EE",X"0E",X"E0",X"E0",X"0E",X"E0",X"E0",X"0E",
		X"0E",X"00",X"E0",X"00",X"0E",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",
		X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",
		X"00",X"00",X"00",X"EE",X"00",X"E0",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"0E",X"EE",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"0E",X"EE",X"00",X"70",X"EE",X"00",X"00",X"70",X"E0",X"00",X"00",X"77",X"00",X"00",X"EE",
		X"77",X"00",X"00",X"EE",X"77",X"00",X"00",X"EE",X"77",X"00",X"00",X"00",X"77",X"00",X"8E",X"00",
		X"77",X"00",X"8E",X"00",X"77",X"00",X"8E",X"00",X"77",X"00",X"8E",X"00",X"77",X"00",X"E8",X"00",
		X"77",X"E0",X"E8",X"0E",X"77",X"7E",X"E8",X"E0",X"77",X"70",X"F5",X"00",X"EE",X"70",X"5F",X"00",
		X"EE",X"7F",X"DD",X"00",X"EE",X"5F",X"DD",X"00",X"EE",X"55",X"DD",X"00",X"EE",X"F5",X"DD",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"0E",X"EE",X"00",X"00",X"EE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"EE",
		X"00",X"00",X"00",X"EE",X"30",X"00",X"00",X"EE",X"33",X"00",X"00",X"E0",X"33",X"00",X"00",X"00",
		X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"3E",X"00",X"DD",X"00",X"3E",X"00",X"DD",X"00",
		X"3E",X"00",X"DD",X"00",X"EE",X"00",X"DD",X"00",X"7E",X"E0",X"DD",X"00",X"77",X"7E",X"BB",X"00",
		X"77",X"77",X"FB",X"00",X"77",X"77",X"5F",X"00",X"77",X"77",X"FE",X"00",X"77",X"77",X"E8",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"0E",X"EE",X"00",X"00",X"EE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"EE",
		X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"E0",X"00",X"00",X"30",X"EE",X"00",X"00",X"3E",X"8E",X"00",X"00",X"3E",X"8E",X"00",X"00",
		X"3E",X"88",X"00",X"00",X"EE",X"88",X"00",X"00",X"EE",X"88",X"0E",X"00",X"7E",X"E8",X"0E",X"00",
		X"77",X"EE",X"E0",X"EE",X"77",X"77",X"50",X"00",X"77",X"77",X"FB",X"00",X"77",X"77",X"5B",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"BB",X"04",X"00",X"00",X"BB",X"44",X"00",X"00",X"BB",X"44",X"00",X"00",X"00",X"44",
		X"00",X"00",X"0B",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"44",X"BB",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"BB",
		X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"A0",
		X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",
		X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",
		X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"44",X"BB",
		X"55",X"53",X"77",X"77",X"FF",X"33",X"77",X"77",X"55",X"33",X"77",X"77",X"55",X"33",X"77",X"77",
		X"FF",X"33",X"77",X"77",X"55",X"00",X"77",X"22",X"05",X"00",X"07",X"22",X"00",X"40",X"07",X"22",
		X"00",X"40",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"40",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",
		X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",
		X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"40",X"00",X"00",
		X"00",X"40",X"07",X"22",X"05",X"00",X"07",X"22",X"55",X"00",X"77",X"22",X"FF",X"33",X"77",X"77",
		X"55",X"33",X"77",X"77",X"55",X"33",X"77",X"77",X"FF",X"33",X"77",X"77",X"55",X"53",X"77",X"77",
		X"55",X"44",X"77",X"77",X"55",X"44",X"77",X"77",X"FF",X"44",X"77",X"72",X"55",X"44",X"77",X"72",
		X"55",X"44",X"77",X"72",X"05",X"44",X"77",X"22",X"05",X"43",X"77",X"22",X"00",X"33",X"07",X"22",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"40",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",
		X"00",X"04",X"44",X"44",X"00",X"04",X"44",X"44",X"00",X"04",X"44",X"44",X"00",X"04",X"44",X"44",
		X"00",X"04",X"44",X"44",X"00",X"04",X"44",X"44",X"00",X"04",X"44",X"44",X"00",X"00",X"44",X"44",
		X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"40",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"44",X"00",X"77",X"00",X"44",X"00",X"77",X"00",X"44",X"00",X"77",X"00",X"44",X"00",X"77",
		X"00",X"44",X"03",X"77",X"00",X"44",X"33",X"77",X"00",X"44",X"33",X"77",X"00",X"44",X"33",X"77",
		X"00",X"44",X"33",X"77",X"00",X"44",X"33",X"77",X"00",X"44",X"53",X"70",X"00",X"44",X"35",X"00",
		X"00",X"44",X"53",X"00",X"00",X"44",X"33",X"00",X"00",X"43",X"33",X"00",X"00",X"33",X"33",X"00",
		X"00",X"33",X"33",X"00",X"00",X"33",X"33",X"00",X"00",X"33",X"33",X"00",X"00",X"3B",X"33",X"00",
		X"00",X"3A",X"34",X"00",X"00",X"33",X"34",X"44",X"00",X"BB",X"44",X"44",X"00",X"BB",X"44",X"44",
		X"04",X"BB",X"44",X"44",X"04",X"BB",X"44",X"44",X"04",X"AB",X"44",X"00",X"04",X"BB",X"44",X"00",
		X"04",X"AA",X"40",X"00",X"04",X"AA",X"00",X"00",X"04",X"4A",X"00",X"00",X"44",X"00",X"00",X"00",
		X"77",X"77",X"DD",X"00",X"77",X"77",X"DD",X"00",X"77",X"70",X"DD",X"00",X"77",X"00",X"DD",X"00",
		X"77",X"00",X"0D",X"0E",X"77",X"00",X"E0",X"EE",X"77",X"00",X"00",X"EE",X"77",X"00",X"00",X"E0",
		X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",
		X"00",X"EE",X"EE",X"00",X"00",X"EE",X"E0",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",
		X"55",X"B0",X"00",X"00",X"FF",X"00",X"00",X"00",X"55",X"BB",X"00",X"00",X"55",X"00",X"00",X"00",
		X"FF",X"BB",X"00",X"00",X"55",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"E0",
		X"00",X"00",X"0E",X"EE",X"00",X"00",X"0E",X"EE",X"00",X"00",X"0E",X"EE",X"00",X"0E",X"0E",X"0E",
		X"00",X"EE",X"0E",X"0E",X"00",X"EE",X"0E",X"00",X"00",X"E0",X"0E",X"00",X"00",X"00",X"0E",X"00",
		X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"0E",X"00",X"00",X"0E",X"E0",
		X"00",X"00",X"0E",X"E0",X"00",X"00",X"0E",X"00",X"00",X"E0",X"0E",X"00",X"00",X"0E",X"0E",X"00",
		X"00",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"EE",X"00",X"0E",X"00",
		X"EE",X"00",X"DE",X"00",X"EE",X"05",X"DD",X"00",X"EE",X"55",X"DD",X"00",X"77",X"5F",X"DD",X"EE",
		X"33",X"33",X"00",X"05",X"33",X"44",X"40",X"55",X"03",X"44",X"44",X"5F",X"03",X"44",X"44",X"F5",
		X"00",X"44",X"44",X"55",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"00",X"00",
		X"00",X"45",X"00",X"00",X"00",X"5F",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"5F",X"00",X"00",
		X"AA",X"BB",X"00",X"00",X"AA",X"BB",X"00",X"E0",X"AA",X"BB",X"00",X"0E",X"00",X"BB",X"00",X"0E",
		X"00",X"BB",X"44",X"EE",X"00",X"BA",X"44",X"EE",X"00",X"BA",X"44",X"E0",X"00",X"B6",X"44",X"00",
		X"00",X"B6",X"44",X"50",X"00",X"BB",X"44",X"0B",X"00",X"B0",X"04",X"BB",X"00",X"00",X"00",X"BB",
		X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"D0",X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",
		X"00",X"B0",X"D0",X"00",X"00",X"55",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"F5",X"00",X"00",
		X"00",X"57",X"00",X"00",X"00",X"57",X"00",X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",
		X"00",X"0E",X"EE",X"00",X"00",X"EE",X"EE",X"70",X"00",X"EE",X"0E",X"77",X"00",X"E0",X"07",X"77",
		X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"07",X"77",X"77",X"00",X"77",X"7E",X"70",
		X"00",X"77",X"7E",X"00",X"00",X"77",X"E7",X"E0",X"00",X"77",X"E7",X"EE",X"07",X"77",X"77",X"EE",
		X"77",X"77",X"70",X"EE",X"77",X"77",X"00",X"0E",X"77",X"77",X"00",X"00",X"77",X"37",X"00",X"EE",
		X"77",X"33",X"00",X"00",X"73",X"33",X"00",X"00",X"73",X"33",X"0E",X"00",X"73",X"33",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"40",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",
		X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",
		X"00",X"00",X"00",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",
		X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"40",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",
		X"00",X"04",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"FF",X"00",
		X"00",X"44",X"44",X"00",X"00",X"FF",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"05",
		X"00",X"44",X"44",X"55",X"00",X"44",X"44",X"05",X"00",X"44",X"44",X"00",X"00",X"44",X"45",X"00",
		X"00",X"44",X"55",X"00",X"00",X"44",X"55",X"00",X"00",X"44",X"55",X"00",X"00",X"55",X"55",X"00",
		X"00",X"05",X"55",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",
		X"00",X"06",X"66",X"00",X"00",X"66",X"66",X"00",X"00",X"6F",X"66",X"00",X"00",X"6F",X"66",X"00",
		X"00",X"FF",X"66",X"00",X"00",X"FF",X"66",X"00",X"00",X"F6",X"66",X"00",X"00",X"F6",X"66",X"06",
		X"00",X"66",X"66",X"66",X"00",X"66",X"66",X"0D",X"00",X"66",X"66",X"00",X"00",X"66",X"66",X"00",
		X"00",X"66",X"66",X"00",X"00",X"66",X"DD",X"00",X"00",X"66",X"DD",X"00",X"00",X"86",X"DD",X"00",
		X"00",X"06",X"DD",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"C0",X"00",X"CC",X"AA",X"CC",X"00",X"CA",X"AA",X"AC",
		X"00",X"AA",X"CA",X"CC",X"00",X"AA",X"CC",X"C0",X"00",X"AA",X"FC",X"C0",X"00",X"AA",X"CC",X"CC",
		X"00",X"AA",X"CC",X"AC",X"00",X"AA",X"CC",X"AC",X"00",X"AA",X"CC",X"CC",X"00",X"AA",X"CA",X"C0",
		X"00",X"AA",X"CC",X"C0",X"00",X"AA",X"FC",X"CC",X"00",X"AA",X"CC",X"AC",X"00",X"AA",X"CC",X"AC",
		X"00",X"AA",X"CC",X"CC",X"00",X"AA",X"CC",X"C0",X"00",X"AA",X"CA",X"CC",X"00",X"AA",X"AA",X"AC",
		X"00",X"CA",X"AA",X"AC",X"00",X"CC",X"AA",X"CC",X"00",X"00",X"CC",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"C0",X"00",X"CC",X"66",X"CC",X"00",X"C6",X"66",X"6C",
		X"00",X"66",X"C6",X"CC",X"00",X"66",X"CC",X"C0",X"00",X"66",X"FC",X"C0",X"00",X"66",X"CC",X"CC",
		X"00",X"66",X"CC",X"6C",X"00",X"66",X"CC",X"6C",X"00",X"66",X"CC",X"CC",X"00",X"66",X"C6",X"C0",
		X"00",X"66",X"CC",X"C0",X"00",X"66",X"FC",X"CC",X"00",X"66",X"CC",X"6C",X"00",X"66",X"CC",X"6C",
		X"00",X"66",X"CC",X"CC",X"00",X"66",X"CC",X"C0",X"00",X"66",X"C6",X"CC",X"00",X"66",X"66",X"6C",
		X"00",X"C6",X"66",X"6C",X"00",X"CC",X"66",X"CC",X"00",X"00",X"CC",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"C0",X"00",X"CC",X"BB",X"CC",X"00",X"CB",X"BB",X"BC",
		X"00",X"BB",X"CB",X"CC",X"00",X"BB",X"CC",X"C0",X"00",X"BB",X"FC",X"C0",X"00",X"BB",X"CC",X"CC",
		X"00",X"BB",X"CC",X"BC",X"00",X"BB",X"CC",X"BC",X"00",X"BB",X"CC",X"CC",X"00",X"BB",X"CB",X"C0",
		X"00",X"BB",X"CC",X"C0",X"00",X"BB",X"FC",X"CC",X"00",X"BB",X"CC",X"BC",X"00",X"BB",X"CC",X"BC",
		X"00",X"BB",X"CC",X"CC",X"00",X"BB",X"CC",X"C0",X"00",X"BB",X"CB",X"CC",X"00",X"BB",X"BB",X"BC",
		X"00",X"CB",X"BB",X"BC",X"00",X"CC",X"BB",X"CC",X"00",X"00",X"CC",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",
		X"00",X"0A",X"AA",X"00",X"00",X"AA",X"AA",X"00",X"00",X"AA",X"AA",X"00",X"00",X"AA",X"FF",X"00",
		X"00",X"AA",X"AA",X"00",X"00",X"FF",X"AA",X"00",X"00",X"FF",X"AA",X"00",X"00",X"AA",X"AA",X"0A",
		X"00",X"AA",X"AA",X"AA",X"00",X"AA",X"AA",X"0A",X"00",X"AA",X"AA",X"00",X"00",X"AA",X"A9",X"00",
		X"00",X"AA",X"99",X"00",X"00",X"AA",X"99",X"00",X"00",X"9A",X"99",X"00",X"00",X"A9",X"99",X"00",
		X"00",X"0A",X"99",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"7F",X"00",
		X"00",X"00",X"66",X"00",X"00",X"FF",X"66",X"00",X"00",X"00",X"64",X"00",X"00",X"00",X"04",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"05",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"0A",X"00",X"00",X"00",X"A4",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"00",X"45",X"00",X"00",X"FF",X"40",X"00",X"00",X"00",X"04",X"00",
		X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"40",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"65",X"00",
		X"00",X"04",X"64",X"00",X"00",X"0A",X"54",X"00",X"00",X"0A",X"04",X"00",X"00",X"00",X"05",X"00",
		X"00",X"05",X"05",X"00",X"00",X"05",X"05",X"00",X"00",X"00",X"05",X"00",X"00",X"AA",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"40",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",
		X"00",X"00",X"44",X"44",X"00",X"00",X"04",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",
		X"00",X"00",X"00",X"44",X"00",X"00",X"04",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",
		X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"40",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"00",X"00",X"00",X"44",X"00",X"40",X"00",X"44",X"00",X"40",X"00",X"44",X"00",X"44",
		X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",
		X"00",X"44",X"04",X"44",X"00",X"44",X"04",X"44",X"00",X"44",X"04",X"40",X"00",X"04",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"04",X"00",X"99",X"90",X"00",X"00",X"A9",X"99",X"00",X"00",X"9A",X"99",
		X"0A",X"09",X"9A",X"99",X"00",X"09",X"A9",X"99",X"00",X"09",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"09",X"99",X"99",X"00",X"09",X"A9",X"99",X"00",X"09",X"9A",X"99",X"00",X"00",X"9A",X"99",
		X"00",X"00",X"A9",X"99",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",
		X"00",X"04",X"00",X"00",X"00",X"44",X"00",X"40",X"00",X"44",X"00",X"40",X"00",X"44",X"00",X"44",
		X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"04",X"44",X"00",X"44",X"04",X"44",
		X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"44",X"00",X"44",X"44",X"40",X"00",X"04",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"66",X"60",
		X"00",X"06",X"AA",X"66",X"00",X"06",X"AA",X"A6",X"00",X"06",X"A6",X"A6",X"00",X"06",X"A6",X"A6",
		X"00",X"06",X"A6",X"A6",X"00",X"06",X"A6",X"A6",X"00",X"06",X"A6",X"A6",X"00",X"06",X"A6",X"66",
		X"00",X"00",X"66",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"00",X"06",X"AA",X"A6",
		X"00",X"06",X"AA",X"A6",X"00",X"06",X"AA",X"A6",X"00",X"06",X"6A",X"A6",X"00",X"06",X"66",X"A6",
		X"00",X"06",X"06",X"A6",X"00",X"00",X"00",X"A6",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"66",X"60",
		X"00",X"06",X"AA",X"66",X"00",X"06",X"AA",X"A6",X"00",X"06",X"A6",X"A6",X"00",X"06",X"A6",X"A6",
		X"00",X"06",X"A6",X"A6",X"00",X"06",X"A6",X"A6",X"00",X"06",X"A6",X"A6",X"00",X"06",X"A6",X"66",
		X"00",X"00",X"66",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"60",X"00",X"06",X"AA",X"66",
		X"00",X"06",X"AA",X"A6",X"00",X"06",X"00",X"A6",X"00",X"06",X"00",X"A6",X"00",X"06",X"00",X"A6",
		X"00",X"06",X"00",X"A6",X"00",X"06",X"AA",X"A6",X"00",X"06",X"AA",X"66",X"00",X"00",X"66",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"A6",X"00",X"06",X"66",X"A6",X"00",X"06",X"AA",X"A6",
		X"00",X"06",X"AA",X"A6",X"00",X"06",X"66",X"A6",X"00",X"00",X"00",X"A6",X"00",X"00",X"00",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"66",X"60",X"00",X"06",X"AA",X"66",
		X"00",X"06",X"AA",X"A6",X"00",X"06",X"A6",X"A6",X"00",X"06",X"A6",X"A6",X"00",X"06",X"A6",X"A6",
		X"00",X"06",X"A6",X"A6",X"00",X"06",X"A6",X"A6",X"00",X"06",X"A6",X"66",X"00",X"06",X"66",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"A6",X"00",X"06",X"66",X"A6",X"00",X"06",X"AA",X"A6",
		X"00",X"06",X"AA",X"A6",X"00",X"06",X"66",X"A6",X"00",X"00",X"00",X"A6",X"00",X"00",X"00",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"66",
		X"00",X"06",X"A6",X"A6",X"00",X"06",X"AA",X"A6",X"00",X"06",X"AA",X"A6",X"00",X"06",X"6A",X"A6",
		X"00",X"06",X"66",X"A6",X"00",X"06",X"06",X"A6",X"00",X"06",X"00",X"A6",X"00",X"06",X"00",X"A6",
		X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"A6",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"6A",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"00",X"A6",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"60",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"60",
		X"00",X"06",X"AA",X"66",X"00",X"06",X"AA",X"A6",X"00",X"06",X"AA",X"A6",X"00",X"06",X"AA",X"A6",
		X"00",X"06",X"AA",X"A6",X"00",X"06",X"AA",X"A6",X"00",X"06",X"66",X"A6",X"00",X"06",X"00",X"66",
		X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"A6",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"6A",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"00",X"A6",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"60",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"6A",X"00",
		X"00",X"00",X"6A",X"00",X"00",X"66",X"6A",X"66",X"00",X"AA",X"AA",X"A6",X"00",X"6A",X"AA",X"A6",
		X"00",X"66",X"0A",X"66",X"00",X"06",X"0A",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"0A",X"00",
		X"00",X"00",X"0A",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"6A",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"A6",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"6A",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"00",X"A6",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"60",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"66",X"60",
		X"00",X"06",X"AA",X"66",X"00",X"06",X"AA",X"A6",X"00",X"06",X"A6",X"A6",X"00",X"06",X"A6",X"A6",
		X"00",X"06",X"A6",X"A6",X"00",X"06",X"A6",X"A6",X"00",X"06",X"A6",X"A6",X"00",X"06",X"A6",X"66",
		X"00",X"00",X"66",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"A6",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"6A",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"00",X"A6",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"60",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"C0",X"00",X"CC",X"55",X"CC",X"00",X"C5",X"55",X"5C",
		X"00",X"55",X"C5",X"CC",X"00",X"55",X"CC",X"C0",X"00",X"55",X"FC",X"C0",X"00",X"55",X"CC",X"CC",
		X"00",X"55",X"CC",X"5C",X"00",X"55",X"CC",X"5C",X"00",X"55",X"CC",X"CC",X"00",X"55",X"C5",X"C0",
		X"00",X"55",X"CC",X"C0",X"00",X"55",X"FC",X"CC",X"00",X"55",X"CC",X"5C",X"00",X"55",X"CC",X"5C",
		X"00",X"55",X"CC",X"CC",X"00",X"55",X"CC",X"C0",X"00",X"55",X"C5",X"CC",X"00",X"55",X"55",X"5C",
		X"00",X"C5",X"55",X"5C",X"00",X"CC",X"55",X"CC",X"00",X"00",X"CC",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"0E",X"0E",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"22",X"00",
		X"E0",X"00",X"22",X"00",X"E0",X"00",X"22",X"00",X"EE",X"00",X"22",X"0E",X"EE",X"00",X"00",X"EE",
		X"0E",X"00",X"00",X"EE",X"0E",X"00",X"00",X"EE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",
		X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"E0",X"0E",X"00",X"00",X"EE",X"EE",X"00",
		X"00",X"EE",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",
		X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"D0",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"E0",X"00",
		X"00",X"EE",X"EE",X"00",X"00",X"E0",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"0E",X"00",X"00",X"EE",X"0E",X"00",X"00",X"EE",
		X"EE",X"00",X"00",X"EE",X"EE",X"22",X"00",X"0E",X"E0",X"22",X"00",X"00",X"E0",X"22",X"00",X"00",
		X"E0",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"0E",X"0E",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"00",X"00",X"EE",X"EE",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"E0",X"00",
		X"00",X"EE",X"EE",X"00",X"00",X"E0",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"0E",X"00",X"00",X"EE",X"0E",X"00",X"00",X"EE",
		X"EE",X"00",X"00",X"EE",X"EE",X"00",X"00",X"0E",X"E0",X"00",X"00",X"00",X"E0",X"00",X"88",X"00",
		X"70",X"00",X"88",X"00",X"75",X"00",X"88",X"00",X"05",X"E0",X"88",X"00",X"00",X"0E",X"8E",X"00",
		X"50",X"00",X"E0",X"00",X"50",X"00",X"22",X"00",X"55",X"EE",X"22",X"00",X"E5",X"EE",X"EE",X"EE",
		X"FF",X"34",X"77",X"77",X"FF",X"34",X"77",X"77",X"55",X"34",X"77",X"77",X"55",X"44",X"77",X"77",
		X"55",X"44",X"77",X"77",X"04",X"44",X"77",X"77",X"04",X"44",X"77",X"77",X"04",X"44",X"77",X"77",
		X"00",X"44",X"77",X"77",X"00",X"44",X"07",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"33",X"77",X"22",X"55",X"33",X"77",X"22",X"55",X"33",X"77",X"23",X"FF",X"33",X"77",X"23",
		X"55",X"33",X"77",X"23",X"54",X"33",X"77",X"23",X"54",X"03",X"77",X"23",X"04",X"03",X"77",X"20",
		X"04",X"00",X"BB",X"00",X"04",X"00",X"B7",X"00",X"00",X"44",X"B0",X"00",X"00",X"44",X"BB",X"00",
		X"00",X"44",X"5B",X"00",X"00",X"44",X"5B",X"00",X"00",X"44",X"BB",X"00",X"00",X"00",X"B0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"33",X"77",X"77",X"55",X"33",X"77",X"77",X"FF",X"33",X"77",X"77",X"55",X"33",X"77",X"77",
		X"55",X"33",X"B7",X"77",X"54",X"33",X"B7",X"20",X"54",X"33",X"77",X"20",X"04",X"35",X"77",X"20",
		X"04",X"04",X"77",X"00",X"00",X"44",X"07",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"40",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",
		X"00",X"00",X"00",X"BB",X"00",X"00",X"44",X"BB",X"00",X"00",X"44",X"BB",X"00",X"00",X"44",X"BB",
		X"00",X"00",X"44",X"AB",X"00",X"00",X"04",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"AA",
		X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"BB",
		X"00",X"00",X"04",X"6B",X"00",X"00",X"44",X"BB",X"00",X"00",X"44",X"B7",X"00",X"00",X"44",X"7B",
		X"00",X"00",X"44",X"BB",X"00",X"00",X"04",X"BB",X"00",X"00",X"00",X"BA",X"00",X"00",X"00",X"AA",
		X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"A0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BA",
		X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"6B",X"00",X"00",X"00",X"BB",X"00",X"00",X"04",X"BB",
		X"00",X"00",X"44",X"BB",X"00",X"00",X"44",X"AB",X"00",X"00",X"44",X"BB",X"00",X"00",X"44",X"AB",
		X"00",X"00",X"04",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"01",X"11",
		X"00",X"00",X"01",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"01",X"00",X"00",X"77",X"00",
		X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"70",X"40",X"53",X"77",X"77",X"44",X"55",X"77",X"77",
		X"44",X"33",X"77",X"77",X"44",X"33",X"77",X"77",X"44",X"33",X"77",X"77",X"55",X"33",X"77",X"77",
		X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",
		X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"77",X"00",X"00",X"DD",X"77",X"00",X"00",X"D0",X"77",
		X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",
		X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",
		X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",
		X"00",X"0B",X"00",X"77",X"00",X"0B",X"00",X"77",X"00",X"0B",X"00",X"77",X"00",X"B0",X"00",X"77",
		X"00",X"B0",X"00",X"77",X"00",X"BB",X"00",X"77",X"00",X"BB",X"00",X"77",X"00",X"BB",X"00",X"77",
		X"0B",X"BB",X"00",X"77",X"0B",X"55",X"00",X"77",X"00",X"55",X"00",X"77",X"00",X"55",X"00",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"0E",X"0E",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",
		X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"EE",X"00",X"00",X"0E",X"EE",X"00",X"00",X"EE",
		X"0E",X"00",X"00",X"EE",X"0E",X"00",X"00",X"EE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"0E",X"00",X"00",X"EE",X"EE",X"00",
		X"00",X"EE",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F5",X"EE",X"0D",X"00",X"EE",X"EE",X"DD",X"00",X"77",X"77",X"DD",X"00",X"77",X"75",X"0E",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",
		X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"EE",X"00",X"00",X"EE",X"EE",X"00",X"00",X"0E",
		X"0E",X"00",X"00",X"EE",X"0E",X"00",X"00",X"EE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"0E",X"00",X"00",X"EE",X"EE",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"EE",X"EE",X"EE",X"77",X"EE",X"00",X"00",X"77",X"0E",X"E0",X"00",X"77",X"E0",X"E0",X"00",
		X"00",X"08",X"0E",X"00",X"00",X"08",X"0E",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",
		X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"EE",X"00",X"00",X"0E",X"EE",X"00",X"00",X"0E",
		X"0E",X"0E",X"00",X"EE",X"0E",X"0E",X"00",X"EE",X"00",X"0E",X"00",X"E0",X"00",X"0E",X"00",X"00",
		X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"0E",X"00",X"00",X"EE",X"EE",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",
		X"00",X"B0",X"00",X"77",X"00",X"BB",X"00",X"77",X"00",X"BB",X"00",X"77",X"00",X"BB",X"00",X"77",
		X"00",X"FF",X"07",X"77",X"00",X"5F",X"07",X"77",X"00",X"5F",X"07",X"07",X"00",X"F5",X"07",X"00",
		X"00",X"44",X"77",X"00",X"50",X"44",X"77",X"00",X"50",X"44",X"77",X"21",X"55",X"44",X"77",X"21",
		X"FF",X"34",X"77",X"71",X"55",X"34",X"77",X"71",X"55",X"44",X"77",X"72",X"FF",X"44",X"77",X"72",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"B0",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"5B",X"00",X"00",X"B0",X"5B",X"00",X"00",X"B0",X"F0",X"00",
		X"00",X"B0",X"F0",X"01",X"00",X"B0",X"00",X"01",X"00",X"BB",X"07",X"11",X"00",X"BB",X"77",X"11",
		X"00",X"BB",X"77",X"11",X"50",X"BB",X"77",X"11",X"50",X"BB",X"77",X"11",X"55",X"3B",X"77",X"11",
		X"FF",X"35",X"77",X"77",X"55",X"35",X"77",X"77",X"55",X"35",X"77",X"77",X"FF",X"33",X"77",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"B0",X"00",X"00",
		X"0B",X"B0",X"00",X"10",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",
		X"00",X"50",X"00",X"11",X"00",X"F5",X"00",X"11",X"00",X"44",X"01",X"11",X"00",X"44",X"01",X"11",
		X"00",X"44",X"11",X"11",X"00",X"44",X"11",X"11",X"00",X"44",X"77",X"10",X"00",X"45",X"77",X"10",
		X"00",X"55",X"77",X"70",X"50",X"33",X"77",X"77",X"50",X"33",X"77",X"77",X"55",X"33",X"77",X"77",
		X"FF",X"33",X"77",X"77",X"55",X"33",X"77",X"77",X"55",X"33",X"77",X"77",X"FF",X"33",X"77",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"B0",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"F5",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"07",X"00",X"44",X"00",X"77",X"00",X"44",X"00",X"77",
		X"00",X"44",X"00",X"77",X"00",X"45",X"00",X"77",X"00",X"55",X"77",X"77",X"00",X"33",X"77",X"77",
		X"00",X"33",X"77",X"77",X"50",X"33",X"77",X"77",X"50",X"33",X"77",X"77",X"55",X"33",X"77",X"77",
		X"FF",X"33",X"77",X"77",X"FF",X"33",X"77",X"77",X"55",X"33",X"77",X"77",X"55",X"33",X"77",X"77",
		X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",
		X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"D0",X"00",X"00",X"DD",X"00",
		X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0B",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"5B",X"00",
		X"00",X"00",X"5B",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"50",X"07",X"00",X"00",X"00",X"07",
		X"00",X"44",X"00",X"77",X"00",X"44",X"00",X"77",X"00",X"44",X"00",X"77",X"04",X"44",X"00",X"77",
		X"44",X"44",X"00",X"77",X"44",X"44",X"00",X"77",X"54",X"40",X"07",X"77",X"F4",X"00",X"77",X"77",
		X"54",X"00",X"77",X"77",X"55",X"33",X"77",X"77",X"F3",X"35",X"77",X"77",X"53",X"55",X"77",X"77",
		X"53",X"55",X"77",X"77",X"F3",X"35",X"77",X"72",X"55",X"33",X"77",X"22",X"54",X"00",X"77",X"22",
		X"F4",X"00",X"77",X"22",X"54",X"40",X"07",X"22",X"44",X"44",X"07",X"11",X"44",X"44",X"00",X"11",
		X"04",X"44",X"00",X"11",X"00",X"44",X"00",X"11",X"00",X"44",X"00",X"11",X"00",X"44",X"00",X"01",
		X"00",X"04",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"04",X"00",X"00",X"00",X"54",X"00",X"00",
		X"BB",X"FF",X"00",X"11",X"0B",X"55",X"00",X"11",X"0B",X"FF",X"00",X"11",X"00",X"54",X"00",X"11",
		X"00",X"50",X"00",X"11",X"00",X"00",X"00",X"10",X"00",X"00",X"F1",X"00",X"00",X"00",X"51",X"00",
		X"00",X"00",X"5F",X"0D",X"00",X"00",X"FF",X"DD",X"00",X"00",X"F5",X"DD",X"00",X"00",X"BD",X"DD",
		X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",
		X"77",X"77",X"BD",X"00",X"77",X"77",X"BD",X"00",X"77",X"EE",X"DD",X"00",X"77",X"00",X"DD",X"E0",
		X"00",X"00",X"0D",X"EE",X"00",X"0E",X"00",X"00",X"0E",X"0E",X"E0",X"00",X"E0",X"E0",X"E0",X"00",
		X"E0",X"E0",X"0E",X"00",X"E0",X"00",X"0E",X"00",X"EE",X"00",X"00",X"0E",X"EE",X"00",X"00",X"0E",
		X"0E",X"00",X"00",X"EE",X"0E",X"00",X"00",X"EE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"0E",X"00",X"00",X"EE",X"EE",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"BB",X"00",X"00",X"EE",X"BD",X"00",X"00",X"33",X"BD",X"E0",X"00",X"33",X"DD",X"0E",X"00",
		X"33",X"DD",X"00",X"00",X"30",X"DD",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",
		X"E0",X"00",X"00",X"E0",X"E0",X"00",X"00",X"0E",X"EE",X"00",X"00",X"0E",X"EE",X"00",X"00",X"0E",
		X"0E",X"00",X"00",X"EE",X"0E",X"00",X"E0",X"EE",X"00",X"00",X"E0",X"E0",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"E0",X"0E",X"00",X"00",X"EE",X"EE",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"EE",X"EE",X"00",X"00",X"E0",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",
		X"00",X"00",X"E0",X"00",X"70",X"00",X"E0",X"E0",X"7E",X"08",X"E0",X"EE",X"7E",X"08",X"00",X"EE",
		X"77",X"08",X"80",X"0E",X"77",X"00",X"82",X"0E",X"77",X"00",X"82",X"0E",X"77",X"00",X"82",X"E0",
		X"77",X"00",X"82",X"00",X"77",X"00",X"88",X"00",X"77",X"E0",X"88",X"00",X"77",X"5E",X"58",X"00",
		X"77",X"5E",X"3E",X"00",X"77",X"F5",X"D0",X"00",X"77",X"F5",X"D0",X"00",X"37",X"BB",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"EE",X"EE",X"00",X"00",X"E0",X"0E",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"E0",X"0E",X"0E",X"00",X"EE",X"3E",X"0D",X"00",X"EE",
		X"EE",X"0D",X"00",X"0E",X"EE",X"0D",X"00",X"0E",X"E7",X"0D",X"22",X"00",X"E7",X"0D",X"22",X"00",
		X"E7",X"00",X"22",X"00",X"77",X"00",X"22",X"00",X"77",X"00",X"DD",X"00",X"77",X"00",X"DD",X"00",
		X"77",X"E0",X"DD",X"00",X"77",X"77",X"E0",X"00",X"77",X"77",X"88",X"00",X"77",X"77",X"88",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"EE",X"EE",X"00",X"00",X"E0",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"0E",X"00",X"00",X"EE",X"0E",X"00",X"00",X"EE",
		X"EE",X"00",X"00",X"0E",X"EE",X"00",X"00",X"0E",X"E0",X"80",X"0D",X"00",X"E0",X"E8",X"DD",X"00",
		X"E0",X"E8",X"DD",X"00",X"7E",X"8E",X"DD",X"00",X"70",X"8E",X"DD",X"00",X"77",X"88",X"DD",X"EE",
		X"77",X"80",X"DD",X"E0",X"77",X"EE",X"DD",X"00",X"77",X"77",X"BD",X"00",X"77",X"77",X"BD",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",
		X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",
		X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",
		X"00",X"00",X"B0",X"44",X"00",X"00",X"BB",X"44",X"00",X"00",X"BB",X"44",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"44",X"AA",X"00",X"00",X"44",X"BB",X"00",X"00",X"04",X"BB",X"00",X"00",X"00",X"BB",
		X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"0B",X"B0",
		X"00",X"00",X"0B",X"B0",X"00",X"00",X"4B",X"B0",X"00",X"04",X"4B",X"B0",X"00",X"04",X"4A",X"A5",
		X"53",X"57",X"77",X"7F",X"F3",X"37",X"77",X"75",X"53",X"37",X"77",X"75",X"53",X"37",X"77",X"7F",
		X"F3",X"37",X"77",X"75",X"50",X"07",X"72",X"05",X"40",X"07",X"72",X"00",X"40",X"07",X"72",X"00",
		X"40",X"07",X"70",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"04",X"40",X"00",X"00",X"04",X"40",X"00",X"00",
		X"04",X"40",X"00",X"00",X"04",X"40",X"00",X"00",X"04",X"40",X"00",X"00",X"04",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"0B",X"B0",X"00",X"00",X"0B",
		X"B0",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"B0",X"00",X"00",X"0B",X"B0",X"00",X"00",X"0B",
		X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",
		X"BB",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",
		X"BB",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"40",X"00",X"00",
		X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"77",X"00",
		X"04",X"00",X"77",X"20",X"54",X"00",X"77",X"20",X"55",X"00",X"77",X"20",X"FF",X"33",X"77",X"77",
		X"55",X"33",X"77",X"77",X"55",X"33",X"77",X"77",X"FF",X"33",X"77",X"77",X"55",X"35",X"77",X"77",
		X"55",X"44",X"77",X"22",X"55",X"44",X"77",X"22",X"FF",X"44",X"77",X"21",X"55",X"44",X"77",X"21",
		X"55",X"43",X"77",X"21",X"54",X"33",X"77",X"21",X"54",X"33",X"77",X"20",X"04",X"33",X"77",X"20",
		X"00",X"04",X"77",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"04",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"40",X"00",X"44",X"44",X"40",X"00",X"44",X"44",X"40",X"00",X"44",X"44",X"40",
		X"00",X"44",X"44",X"40",X"00",X"44",X"44",X"40",X"00",X"44",X"44",X"40",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"04",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"44",X"00",X"77",X"00",X"44",X"00",X"77",X"00",X"44",X"03",X"77",X"00",X"44",X"33",X"77",
		X"00",X"44",X"33",X"77",X"00",X"44",X"33",X"77",X"00",X"44",X"33",X"77",X"00",X"44",X"33",X"77",
		X"00",X"44",X"33",X"70",X"00",X"44",X"33",X"00",X"00",X"44",X"53",X"00",X"00",X"44",X"33",X"00",
		X"00",X"43",X"53",X"00",X"00",X"33",X"33",X"00",X"00",X"33",X"33",X"00",X"00",X"33",X"33",X"00",
		X"00",X"33",X"33",X"00",X"00",X"33",X"33",X"00",X"00",X"33",X"30",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"AB",X"00",X"00",X"00",X"AB",X"44",X"44",X"BB",X"BB",X"44",X"44",X"BB",X"BB",X"44",X"44",
		X"BB",X"BB",X"44",X"44",X"4B",X"BB",X"44",X"40",X"44",X"BB",X"44",X"00",X"44",X"BB",X"44",X"00",
		X"44",X"AA",X"00",X"00",X"44",X"AA",X"00",X"00",X"44",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",
		X"77",X"70",X"DD",X"0E",X"77",X"00",X"DD",X"EE",X"77",X"00",X"DD",X"EE",X"77",X"00",X"DD",X"E0",
		X"77",X"00",X"DD",X"E0",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",
		X"77",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"0E",X"0E",X"EE",X"00",
		X"0E",X"E0",X"EE",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",
		X"55",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"55",X"BB",X"00",X"00",X"55",X"00",X"00",X"00",
		X"FF",X"BB",X"00",X"00",X"5B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"B0",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"E0",X"00",X"EE",X"00",X"EE",X"00",X"E0",X"00",X"EE",
		X"00",X"E0",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"0E",
		X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",
		X"E0",X"E0",X"00",X"00",X"E0",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"0E",X"00",
		X"00",X"DD",X"0E",X"00",X"00",X"FD",X"E0",X"00",X"77",X"FD",X"D0",X"00",X"77",X"F5",X"DD",X"EE",
		X"33",X"33",X"00",X"BB",X"33",X"44",X"00",X"BB",X"33",X"44",X"44",X"BB",X"33",X"44",X"44",X"BB",
		X"33",X"44",X"44",X"BB",X"33",X"44",X"44",X"5B",X"03",X"44",X"40",X"0B",X"03",X"54",X"E0",X"00",
		X"00",X"F5",X"0E",X"00",X"00",X"5F",X"00",X"00",X"00",X"F5",X"00",X"0E",X"AA",X"55",X"00",X"0E",
		X"AA",X"BB",X"00",X"EE",X"AA",X"AB",X"00",X"EE",X"AA",X"AA",X"00",X"E0",X"AA",X"BA",X"00",X"E0",
		X"0B",X"BB",X"00",X"00",X"0B",X"AB",X"4E",X"00",X"0B",X"AB",X"44",X"00",X"0B",X"6B",X"44",X"00",
		X"0B",X"60",X"44",X"BB",X"0B",X"BA",X"44",X"BB",X"0B",X"AA",X"44",X"B0",X"00",X"0A",X"44",X"BB",
		X"00",X"00",X"04",X"BB",X"00",X"04",X"00",X"B0",X"00",X"44",X"00",X"BB",X"00",X"44",X"00",X"0B",
		X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",
		X"00",X"0D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"50",X"00",X"00",
		X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"77",X"00",
		X"00",X"EE",X"77",X"00",X"00",X"EE",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"7E",X"70",
		X"00",X"00",X"7E",X"70",X"00",X"77",X"E7",X"70",X"00",X"77",X"E7",X"00",X"00",X"77",X"77",X"00",
		X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"77",X"77",X"77",X"00",X"77",X"77",X"00",X"00",
		X"77",X"77",X"00",X"E0",X"77",X"77",X"00",X"E0",X"77",X"77",X"00",X"E0",X"77",X"77",X"00",X"EE",
		X"33",X"77",X"00",X"EE",X"33",X"37",X"00",X"EE",X"33",X"33",X"EE",X"EB",X"33",X"33",X"00",X"BE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"04",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"04",X"44",X"40",X"00",X"00",X"44",X"40",X"00",X"00",X"04",X"40",X"00",X"00",X"00",X"40",
		X"00",X"00",X"04",X"40",X"00",X"00",X"44",X"40",X"00",X"04",X"44",X"40",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"04",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",
		X"00",X"44",X"40",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"4F",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"EE",X"00",X"44",X"44",X"0E",X"00",X"44",X"45",X"0E",X"00",X"44",X"55",X"00",
		X"00",X"44",X"55",X"00",X"00",X"44",X"55",X"00",X"00",X"44",X"55",X"00",X"00",X"45",X"54",X"00",
		X"00",X"55",X"40",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",
		X"00",X"66",X"60",X"00",X"00",X"66",X"66",X"00",X"00",X"F6",X"66",X"00",X"00",X"FF",X"66",X"00",
		X"00",X"FF",X"66",X"00",X"00",X"66",X"66",X"00",X"00",X"66",X"66",X"00",X"00",X"66",X"66",X"00",
		X"00",X"66",X"66",X"EE",X"00",X"66",X"66",X"0E",X"00",X"66",X"66",X"0E",X"00",X"66",X"6D",X"00",
		X"00",X"66",X"DD",X"00",X"00",X"66",X"DD",X"00",X"00",X"66",X"DD",X"00",X"00",X"6D",X"D6",X"00",
		X"00",X"DD",X"60",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CA",X"AA",X"00",X"00",X"AA",X"AA",X"00",
		X"00",X"AC",X"AA",X"00",X"00",X"CC",X"AA",X"00",X"00",X"CF",X"AA",X"00",X"00",X"CF",X"AA",X"00",
		X"00",X"CF",X"AA",X"00",X"00",X"CC",X"AA",X"00",X"00",X"AC",X"AA",X"00",X"00",X"AC",X"AA",X"00",
		X"00",X"CC",X"AA",X"00",X"00",X"CF",X"AA",X"00",X"00",X"CF",X"AA",X"00",X"00",X"CF",X"AA",X"00",
		X"00",X"CC",X"AA",X"00",X"00",X"AC",X"AA",X"00",X"00",X"AC",X"AA",X"00",X"00",X"AA",X"AA",X"00",
		X"00",X"AA",X"AA",X"00",X"00",X"CA",X"AA",X"00",X"00",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"CC",X"CC",X"00",X"00",X"C6",X"66",X"00",X"00",X"66",X"66",X"00",
		X"00",X"6C",X"66",X"00",X"00",X"CC",X"66",X"00",X"00",X"CF",X"66",X"00",X"00",X"CF",X"66",X"00",
		X"00",X"CF",X"66",X"00",X"00",X"CC",X"66",X"00",X"00",X"6C",X"66",X"00",X"00",X"6C",X"66",X"00",
		X"00",X"CC",X"66",X"00",X"00",X"CF",X"66",X"00",X"00",X"CF",X"66",X"00",X"00",X"CF",X"66",X"00",
		X"00",X"CC",X"66",X"00",X"00",X"6C",X"66",X"00",X"00",X"6C",X"66",X"00",X"00",X"66",X"66",X"00",
		X"00",X"66",X"66",X"00",X"00",X"C6",X"66",X"00",X"00",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CB",X"BB",X"00",X"00",X"BB",X"BB",X"00",
		X"00",X"BC",X"BB",X"00",X"00",X"CC",X"BB",X"00",X"00",X"CF",X"BB",X"00",X"00",X"CF",X"BB",X"00",
		X"00",X"CF",X"BB",X"00",X"00",X"CC",X"BB",X"00",X"00",X"BC",X"BB",X"00",X"00",X"BC",X"BB",X"00",
		X"00",X"CC",X"BB",X"00",X"00",X"CF",X"BB",X"00",X"00",X"CF",X"BB",X"00",X"00",X"CF",X"BB",X"00",
		X"00",X"CC",X"BB",X"00",X"00",X"BC",X"BB",X"00",X"00",X"BC",X"BB",X"00",X"00",X"BB",X"BB",X"00",
		X"00",X"BB",X"BB",X"00",X"00",X"CB",X"BB",X"00",X"00",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",
		X"00",X"AA",X"A0",X"00",X"00",X"AA",X"AA",X"00",X"00",X"AA",X"AA",X"00",X"00",X"AF",X"AA",X"00",
		X"00",X"AF",X"AA",X"00",X"00",X"AA",X"AA",X"00",X"00",X"FA",X"AA",X"00",X"00",X"AA",X"AA",X"00",
		X"00",X"AA",X"AA",X"EE",X"00",X"AA",X"AA",X"0E",X"00",X"AA",X"A9",X"0E",X"00",X"AA",X"99",X"00",
		X"00",X"AA",X"99",X"00",X"00",X"AA",X"99",X"00",X"00",X"9A",X"99",X"00",X"00",X"A9",X"9A",X"00",
		X"00",X"99",X"A0",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"04",X"00",X"00",
		X"00",X"00",X"05",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",
		X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"A4",X"00",X"00",X"AA",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"0A",X"00",X"00",X"00",X"F0",X"50",X"00",X"00",X"05",X"40",X"00",
		X"00",X"50",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"54",X"00",X"00",
		X"00",X"00",X"0A",X"00",X"00",X"00",X"5A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",
		X"04",X"00",X"50",X"00",X"00",X"00",X"05",X"00",X"00",X"A5",X"00",X"00",X"00",X"A5",X"00",X"00",
		X"00",X"0A",X"A0",X"40",X"00",X"0F",X"00",X"04",X"00",X"4A",X"00",X"00",X"00",X"00",X"00",X"00",
		X"05",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"44",X"40",X"00",X"00",X"44",X"40",X"00",X"00",X"44",X"40",X"00",X"00",X"04",X"40",
		X"00",X"00",X"44",X"40",X"00",X"00",X"44",X"40",X"00",X"00",X"44",X"40",X"00",X"00",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"44",X"04",X"00",X"00",X"44",X"04",X"00",X"00",X"44",X"04",X"00",X"00",X"44",X"04",X"00",
		X"00",X"44",X"04",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"04",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"99",X"9A",X"00",X"00",X"99",X"A9",X"00",
		X"A0",X"99",X"A9",X"90",X"AA",X"99",X"9A",X"90",X"AA",X"99",X"99",X"90",X"A6",X"99",X"99",X"90",
		X"00",X"99",X"99",X"90",X"00",X"99",X"9A",X"90",X"00",X"99",X"A9",X"90",X"00",X"99",X"A9",X"00",
		X"00",X"99",X"9A",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"44",X"04",X"00",X"00",X"44",X"04",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"04",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"00",
		X"00",X"A6",X"AA",X"00",X"00",X"AA",X"AA",X"00",X"00",X"AA",X"66",X"00",X"00",X"AA",X"00",X"00",
		X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"6A",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"6A",X"00",X"00",X"00",X"AA",X"60",X"00",
		X"00",X"A6",X"60",X"00",X"00",X"A6",X"A6",X"00",X"00",X"A6",X"AA",X"00",X"00",X"A6",X"AA",X"00",
		X"00",X"AA",X"6A",X"00",X"00",X"6A",X"66",X"00",X"00",X"06",X"06",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"00",
		X"00",X"A6",X"AA",X"00",X"00",X"AA",X"AA",X"00",X"00",X"AA",X"66",X"00",X"00",X"AA",X"00",X"00",
		X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"6A",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"00",X"00",X"6A",X"AA",X"00",
		X"00",X"AA",X"AA",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",
		X"00",X"AA",X"00",X"00",X"00",X"AA",X"AA",X"00",X"00",X"6A",X"AA",X"00",X"00",X"66",X"66",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"00",X"00",X"AA",X"AA",X"00",
		X"00",X"AA",X"AA",X"00",X"00",X"6A",X"66",X"00",X"00",X"66",X"00",X"00",X"00",X"06",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"00",X"00",X"A6",X"AA",X"00",
		X"00",X"AA",X"AA",X"00",X"00",X"AA",X"66",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",
		X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"66",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"00",X"00",X"AA",X"AA",X"00",
		X"00",X"AA",X"AA",X"00",X"00",X"6A",X"66",X"00",X"00",X"66",X"00",X"00",X"00",X"06",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",
		X"00",X"6A",X"60",X"00",X"00",X"AA",X"66",X"00",X"00",X"AA",X"A6",X"00",X"00",X"AA",X"AA",X"00",
		X"00",X"AA",X"AA",X"00",X"00",X"AA",X"6A",X"00",X"00",X"AA",X"66",X"00",X"00",X"6A",X"06",X"00",
		X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"6A",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"A6",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"00",X"6A",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"06",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"00",
		X"00",X"6A",X"AA",X"00",X"00",X"AA",X"AA",X"00",X"00",X"AA",X"66",X"00",X"00",X"AA",X"60",X"00",
		X"00",X"AA",X"60",X"00",X"00",X"AA",X"60",X"00",X"00",X"AA",X"60",X"00",X"00",X"6A",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"6A",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"A6",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"00",X"6A",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"06",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"A6",X"00",
		X"00",X"00",X"A6",X"00",X"00",X"66",X"A6",X"00",X"00",X"AA",X"AA",X"00",X"00",X"AA",X"AA",X"00",
		X"00",X"AA",X"A6",X"00",X"00",X"6A",X"A6",X"00",X"00",X"66",X"A6",X"00",X"00",X"06",X"A6",X"00",
		X"00",X"00",X"A6",X"00",X"00",X"00",X"A6",X"00",X"00",X"00",X"A6",X"00",X"00",X"00",X"A6",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"6A",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"A6",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"00",X"6A",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"06",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"00",
		X"00",X"A6",X"AA",X"00",X"00",X"AA",X"AA",X"00",X"00",X"AA",X"66",X"00",X"00",X"AA",X"00",X"00",
		X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"6A",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"6A",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"A6",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"00",X"6A",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"06",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"CC",X"CC",X"00",X"00",X"C5",X"55",X"00",X"00",X"55",X"55",X"00",
		X"00",X"5C",X"55",X"00",X"00",X"CC",X"55",X"00",X"00",X"CF",X"55",X"00",X"00",X"CF",X"55",X"00",
		X"00",X"CF",X"55",X"00",X"00",X"CC",X"55",X"00",X"00",X"5C",X"55",X"00",X"00",X"5C",X"55",X"00",
		X"00",X"CC",X"55",X"00",X"00",X"CF",X"55",X"00",X"00",X"CF",X"55",X"00",X"00",X"CF",X"55",X"00",
		X"00",X"CC",X"55",X"00",X"00",X"5C",X"55",X"00",X"00",X"5C",X"55",X"00",X"00",X"55",X"55",X"00",
		X"00",X"55",X"55",X"00",X"00",X"C5",X"55",X"00",X"00",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"00",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"E0",X"00",X"0E",
		X"00",X"00",X"00",X"0E",X"00",X"00",X"E0",X"0E",X"00",X"00",X"0E",X"0E",X"00",X"00",X"00",X"EE",
		X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"0E",X"00",X"00",X"E0",X"E0",X"00",X"00",X"E0",
		X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",
		X"0E",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"EE",X"00",X"00",X"EE",X"E0",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",
		X"D0",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"EE",X"E0",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"0E",X"00",X"0E",X"00",X"00",X"00",
		X"0E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",
		X"E0",X"00",X"00",X"E0",X"0E",X"00",X"00",X"E0",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",
		X"00",X"00",X"00",X"EE",X"00",X"00",X"0E",X"0E",X"00",X"00",X"E0",X"0E",X"00",X"00",X"00",X"0E",
		X"00",X"E0",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"EE",X"00",X"00",X"0E",X"EE",X"EE",X"00",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"EE",X"E0",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"0E",X"00",X"0E",X"00",X"00",X"00",
		X"0E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",
		X"E0",X"00",X"00",X"E0",X"0E",X"00",X"00",X"E0",X"00",X"00",X"00",X"EE",X"0D",X"00",X"00",X"EE",
		X"0D",X"00",X"00",X"EE",X"0D",X"00",X"0E",X"0E",X"5D",X"00",X"E0",X"0E",X"DD",X"00",X"00",X"0E",
		X"DD",X"E0",X"00",X"0E",X"DD",X"0E",X"00",X"0E",X"BD",X"11",X"00",X"0E",X"BD",X"EE",X"EE",X"EE",
		X"44",X"44",X"77",X"77",X"44",X"44",X"77",X"77",X"44",X"44",X"77",X"77",X"44",X"44",X"77",X"77",
		X"44",X"44",X"77",X"77",X"44",X"44",X"77",X"77",X"44",X"44",X"77",X"77",X"44",X"44",X"77",X"70",
		X"44",X"44",X"77",X"70",X"00",X"44",X"77",X"00",X"00",X"44",X"00",X"00",X"00",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"77",X"22",X"44",X"33",X"77",X"22",X"44",X"33",X"77",X"33",X"44",X"33",X"77",X"33",
		X"44",X"33",X"77",X"33",X"44",X"33",X"77",X"33",X"44",X"33",X"77",X"30",X"44",X"33",X"77",X"00",
		X"44",X"00",X"70",X"00",X"44",X"00",X"7B",X"00",X"44",X"44",X"BB",X"00",X"44",X"44",X"B0",X"00",
		X"44",X"44",X"BB",X"00",X"44",X"44",X"BB",X"00",X"04",X"44",X"B0",X"00",X"04",X"00",X"BB",X"00",
		X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"77",X"77",X"33",X"33",X"77",X"77",X"44",X"33",X"77",X"77",X"44",X"33",X"77",X"77",
		X"44",X"35",X"77",X"77",X"44",X"5F",X"77",X"00",X"44",X"55",X"77",X"00",X"44",X"55",X"77",X"00",
		X"44",X"5F",X"77",X"00",X"44",X"F5",X"77",X"00",X"44",X"40",X"00",X"00",X"04",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BA",X"00",X"00",X"04",X"BA",X"00",X"00",X"04",X"BA",
		X"00",X"00",X"44",X"BB",X"00",X"00",X"44",X"BB",X"00",X"00",X"44",X"BB",X"00",X"00",X"44",X"BB",
		X"00",X"00",X"44",X"BB",X"00",X"00",X"44",X"AB",X"00",X"00",X"44",X"AA",X"00",X"00",X"04",X"A0",
		X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0A",X"00",X"00",X"04",X"0A",X"00",X"00",X"44",X"00",
		X"00",X"00",X"44",X"BB",X"00",X"00",X"44",X"BB",X"00",X"00",X"44",X"BB",X"00",X"00",X"44",X"BA",
		X"00",X"00",X"44",X"AA",X"00",X"00",X"44",X"AA",X"00",X"00",X"44",X"AA",X"00",X"00",X"04",X"AA",
		X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",
		X"00",X"00",X"00",X"BB",X"00",X"00",X"04",X"BB",X"00",X"00",X"44",X"AA",X"00",X"00",X"44",X"BB",
		X"00",X"00",X"44",X"BB",X"00",X"00",X"44",X"BB",X"00",X"00",X"44",X"AB",X"00",X"00",X"44",X"AA",
		X"00",X"00",X"44",X"A0",X"00",X"00",X"44",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"01",X"11",
		X"00",X"00",X"01",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",
		X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"77",X"11",
		X"00",X"00",X"77",X"11",X"00",X"00",X"77",X"01",X"00",X"33",X"77",X"77",X"00",X"33",X"77",X"77",
		X"40",X"33",X"77",X"77",X"45",X"33",X"77",X"77",X"33",X"33",X"77",X"77",X"33",X"33",X"77",X"77",
		X"00",X"00",X"DD",X"D0",X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"D0",
		X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"B0",X"00",X"00",X"B0",X"B0",X"00",X"00",
		X"BB",X"00",X"00",X"70",X"0B",X"00",X"00",X"70",X"0B",X"00",X"00",X"77",X"00",X"0B",X"00",X"77",
		X"00",X"B0",X"00",X"77",X"00",X"B0",X"00",X"77",X"0B",X"00",X"00",X"77",X"BB",X"00",X"00",X"77",
		X"B0",X"00",X"00",X"77",X"00",X"F0",X"00",X"77",X"00",X"F0",X"07",X"77",X"00",X"F0",X"07",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"00",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"E0",X"00",X"0E",
		X"00",X"00",X"00",X"0E",X"00",X"00",X"E0",X"0E",X"00",X"00",X"0E",X"0E",X"00",X"00",X"00",X"EE",
		X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"0E",X"00",X"00",X"E0",X"E0",X"00",X"00",X"E0",
		X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",
		X"0E",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"EE",X"00",X"00",X"EE",X"E0",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"BD",X"EE",X"D0",X"0E",X"DD",X"55",X"DD",X"0E",X"DD",X"7E",X"DD",X"0E",X"77",X"E5",X"00",X"0E",
		X"00",X"00",X"E0",X"0E",X"00",X"00",X"0E",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"EE",
		X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"0E",X"00",X"00",X"E0",X"E0",X"00",X"00",X"E0",
		X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",
		X"0E",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"EE",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"EE",X"EE",X"EE",X"77",X"88",X"00",X"0E",X"77",X"88",X"00",X"0E",X"00",X"88",X"00",X"0E",
		X"00",X"88",X"00",X"0E",X"00",X"88",X"00",X"0E",X"00",X"0E",X"E0",X"0E",X"00",X"0E",X"E0",X"EE",
		X"0E",X"E0",X"0E",X"EE",X"E0",X"E0",X"0E",X"EE",X"00",X"E0",X"00",X"E0",X"00",X"E0",X"00",X"E0",
		X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",
		X"0E",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"EE",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",
		X"00",X"00",X"07",X"70",X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",
		X"00",X"50",X"77",X"77",X"00",X"55",X"77",X"77",X"00",X"F5",X"77",X"77",X"00",X"45",X"77",X"77",
		X"00",X"40",X"77",X"77",X"05",X"43",X"77",X"07",X"03",X"43",X"77",X"11",X"33",X"44",X"77",X"11",
		X"33",X"44",X"77",X"11",X"33",X"44",X"77",X"11",X"33",X"44",X"77",X"22",X"33",X"44",X"77",X"22",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"B0",X"00",
		X"00",X"00",X"B0",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"11",X"00",X"04",X"00",X"11",X"00",X"04",X"77",X"11",X"00",X"B4",X"77",X"11",
		X"00",X"BB",X"77",X"11",X"05",X"BB",X"77",X"11",X"03",X"BB",X"77",X"11",X"33",X"BB",X"77",X"11",
		X"33",X"F5",X"77",X"77",X"33",X"F5",X"77",X"77",X"33",X"F5",X"77",X"77",X"33",X"44",X"77",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"B0",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"0B",X"00",X"01",X"10",X"00",X"00",X"01",X"11",
		X"0B",X"00",X"11",X"11",X"BB",X"00",X"11",X"11",X"B0",X"00",X"11",X"11",X"00",X"00",X"11",X"11",
		X"00",X"40",X"11",X"11",X"00",X"44",X"11",X"11",X"00",X"44",X"77",X"11",X"00",X"44",X"77",X"11",
		X"00",X"54",X"77",X"01",X"05",X"33",X"77",X"77",X"03",X"33",X"77",X"77",X"33",X"33",X"77",X"77",
		X"33",X"33",X"77",X"77",X"33",X"33",X"77",X"77",X"33",X"33",X"77",X"77",X"33",X"33",X"77",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"5F",X"00",X"00",X"00",X"5F",X"00",X"00",X"00",X"5F",X"00",X"00",X"00",X"44",X"00",X"07",
		X"00",X"44",X"00",X"77",X"00",X"44",X"00",X"77",X"00",X"44",X"00",X"77",X"00",X"44",X"00",X"77",
		X"00",X"44",X"00",X"77",X"00",X"44",X"00",X"77",X"00",X"54",X"77",X"77",X"00",X"33",X"77",X"77",
		X"00",X"33",X"77",X"77",X"05",X"33",X"77",X"77",X"03",X"33",X"77",X"77",X"33",X"33",X"77",X"77",
		X"33",X"33",X"77",X"77",X"33",X"33",X"77",X"77",X"33",X"33",X"77",X"72",X"33",X"33",X"77",X"22",
		X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",
		X"00",X"00",X"DD",X"DD",X"00",X"0D",X"DD",X"D0",X"00",X"0D",X"DD",X"00",X"00",X"0D",X"DD",X"00",
		X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"07",X"00",X"00",X"BB",X"07",
		X"00",X"00",X"B0",X"77",X"00",X"00",X"00",X"77",X"00",X"04",X"00",X"77",X"00",X"44",X"00",X"77",
		X"00",X"44",X"00",X"77",X"00",X"44",X"00",X"77",X"44",X"44",X"00",X"77",X"44",X"44",X"00",X"77",
		X"44",X"40",X"00",X"77",X"44",X"00",X"07",X"77",X"44",X"00",X"77",X"77",X"44",X"00",X"77",X"77",
		X"44",X"00",X"77",X"70",X"33",X"33",X"77",X"70",X"33",X"33",X"77",X"20",X"35",X"53",X"77",X"2E",
		X"35",X"53",X"77",X"EE",X"33",X"33",X"77",X"11",X"33",X"33",X"77",X"11",X"44",X"03",X"77",X"11",
		X"44",X"00",X"77",X"11",X"44",X"00",X"77",X"11",X"44",X"00",X"77",X"11",X"44",X"40",X"00",X"11",
		X"44",X"44",X"00",X"11",X"44",X"44",X"00",X"11",X"00",X"44",X"00",X"11",X"00",X"44",X"00",X"11",
		X"00",X"44",X"00",X"01",X"00",X"44",X"00",X"00",X"B0",X"44",X"00",X"00",X"BB",X"44",X"00",X"11",
		X"BB",X"44",X"00",X"11",X"BB",X"44",X"00",X"11",X"BB",X"40",X"00",X"11",X"BB",X"00",X"00",X"11",
		X"0B",X"00",X"01",X"11",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"DD",
		X"00",X"00",X"F5",X"DD",X"00",X"00",X"5F",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",
		X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"0D",X"DD",X"00",X"00",X"00",X"DD",
		X"77",X"75",X"D2",X"0E",X"77",X"7F",X"D2",X"0E",X"77",X"05",X"DD",X"0E",X"77",X"0E",X"DD",X"0E",
		X"00",X"E0",X"DD",X"EE",X"EE",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"EE",
		X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"E0",X"E0",X"00",X"00",X"E0",X"E0",
		X"E0",X"00",X"0E",X"00",X"E0",X"00",X"0E",X"00",X"EE",X"00",X"0E",X"00",X"0E",X"00",X"00",X"00",
		X"0E",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"EE",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3E",X"DD",X"00",X"0E",X"E3",X"DD",X"00",X"0E",X"33",X"DD",X"00",X"0E",X"33",X"D2",X"00",X"0E",
		X"30",X"D2",X"EE",X"0E",X"00",X"D2",X"00",X"0E",X"00",X"02",X"00",X"0E",X"00",X"00",X"00",X"EE",
		X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"0E",X"00",X"00",X"E0",X"E0",X"00",X"00",X"E0",
		X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",
		X"0E",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"EE",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"0E",X"00",X"0E",X"00",X"00",X"00",
		X"0E",X"00",X"00",X"00",X"EE",X"88",X"00",X"00",X"E0",X"88",X"00",X"00",X"E0",X"88",X"00",X"00",
		X"E0",X"88",X"00",X"E0",X"7E",X"88",X"20",X"E0",X"77",X"00",X"20",X"EE",X"77",X"00",X"20",X"EE",
		X"77",X"00",X"20",X"EE",X"77",X"00",X"80",X"0E",X"77",X"00",X"80",X"0E",X"77",X"00",X"EE",X"0E",
		X"77",X"30",X"00",X"0E",X"77",X"33",X"00",X"0E",X"77",X"33",X"00",X"0E",X"77",X"5D",X"00",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"0E",X"00",X"0E",X"00",X"00",X"00",
		X"0E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"DD",X"00",X"00",
		X"00",X"DD",X"00",X"E0",X"00",X"DD",X"00",X"E0",X"E0",X"DD",X"0E",X"EE",X"7E",X"DD",X"0E",X"EE",
		X"77",X"0E",X"E0",X"EE",X"77",X"0E",X"E0",X"0E",X"77",X"0E",X"00",X"0E",X"77",X"0E",X"00",X"0E",
		X"77",X"0E",X"00",X"0E",X"77",X"75",X"00",X"0E",X"77",X"77",X"00",X"0E",X"77",X"77",X"00",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"0E",X"00",X"0E",X"00",X"00",X"00",
		X"0E",X"00",X"00",X"00",X"EE",X"00",X"0E",X"00",X"E0",X"00",X"0E",X"00",X"E0",X"00",X"0E",X"00",
		X"00",X"00",X"E0",X"E0",X"00",X"00",X"E0",X"E0",X"00",X"00",X"D0",X"EE",X"00",X"00",X"DD",X"EE",
		X"00",X"00",X"DD",X"EE",X"00",X"00",X"DD",X"0E",X"EE",X"00",X"DD",X"0E",X"00",X"E0",X"DD",X"EE",
		X"77",X"0E",X"DD",X"0E",X"77",X"05",X"DD",X"0E",X"77",X"7F",X"D2",X"0E",X"77",X"75",X"D2",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",
		X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",
		X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"55",
		X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",
		X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"04",
		X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",
		X"00",X"00",X"00",X"44",X"00",X"00",X"05",X"44",X"00",X"00",X"B5",X"44",X"00",X"00",X"BF",X"04",
		X"00",X"00",X"B5",X"04",X"00",X"0B",X"05",X"00",X"00",X"0B",X"00",X"00",X"00",X"B0",X"00",X"00",
		X"00",X"00",X"44",X"BB",X"00",X"00",X"44",X"BA",X"00",X"00",X"44",X"AB",X"00",X"00",X"44",X"BB",
		X"00",X"00",X"04",X"B0",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"04",X"B0",
		X"00",X"00",X"44",X"BB",X"00",X"00",X"44",X"AB",X"00",X"00",X"44",X"BA",X"00",X"00",X"44",X"BB",
		X"33",X"55",X"77",X"77",X"33",X"53",X"77",X"77",X"33",X"33",X"77",X"77",X"33",X"33",X"77",X"77",
		X"44",X"33",X"77",X"77",X"44",X"03",X"77",X"00",X"44",X"00",X"77",X"00",X"44",X"00",X"77",X"00",
		X"44",X"00",X"77",X"00",X"44",X"00",X"77",X"00",X"44",X"00",X"00",X"00",X"04",X"00",X"00",X"00",
		X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"5F",X"00",X"00",X"00",
		X"BF",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",
		X"B0",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",
		X"B0",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",
		X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BF",X"00",X"00",X"00",
		X"5F",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"02",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",
		X"04",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"70",X"00",
		X"44",X"00",X"77",X"00",X"44",X"00",X"77",X"00",X"44",X"03",X"77",X"00",X"44",X"33",X"77",X"77",
		X"33",X"33",X"77",X"77",X"33",X"33",X"77",X"77",X"33",X"53",X"77",X"77",X"33",X"55",X"77",X"77",
		X"33",X"44",X"77",X"22",X"44",X"44",X"77",X"22",X"44",X"43",X"77",X"11",X"44",X"33",X"77",X"11",
		X"44",X"33",X"77",X"11",X"44",X"33",X"77",X"10",X"44",X"33",X"77",X"00",X"44",X"33",X"77",X"00",
		X"44",X"44",X"77",X"00",X"00",X"44",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"04",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"04",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"77",X"00",X"00",X"3F",X"77",X"00",X"00",X"3F",X"77",X"00",X"00",X"3F",X"77",
		X"00",X"00",X"3F",X"77",X"00",X"00",X"33",X"77",X"00",X"00",X"33",X"77",X"00",X"00",X"33",X"77",
		X"00",X"00",X"33",X"00",X"00",X"03",X"33",X"00",X"00",X"33",X"33",X"00",X"00",X"33",X"33",X"00",
		X"00",X"33",X"33",X"00",X"00",X"33",X"33",X"00",X"00",X"33",X"33",X"00",X"00",X"33",X"33",X"00",
		X"00",X"35",X"30",X"00",X"00",X"33",X"00",X"00",X"04",X"33",X"00",X"00",X"04",X"B3",X"00",X"00",
		X"AA",X"B3",X"00",X"00",X"AA",X"B3",X"44",X"44",X"BB",X"B3",X"44",X"44",X"6B",X"B3",X"44",X"44",
		X"B6",X"B3",X"44",X"44",X"6B",X"B3",X"44",X"00",X"BB",X"A4",X"44",X"00",X"4A",X"A0",X"00",X"00",
		X"44",X"A0",X"00",X"00",X"44",X"A0",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"0D",X"D0",X"E0",X"77",X"00",X"D0",X"00",X"77",X"00",X"D0",X"00",X"77",X"00",X"D0",X"00",
		X"77",X"00",X"D0",X"00",X"77",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"70",X"00",X"00",X"00",
		X"00",X"0E",X"0E",X"00",X"00",X"E0",X"EE",X"00",X"00",X"E0",X"EE",X"00",X"EE",X"00",X"E0",X"00",
		X"EE",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0B",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"B0",X"00",X"00",X"BB",X"00",X"00",X"00",
		X"BB",X"BB",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",
		X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",
		X"0E",X"00",X"00",X"EE",X"0E",X"00",X"00",X"EE",X"EE",X"00",X"00",X"EE",X"EE",X"00",X"00",X"0E",
		X"E0",X"00",X"00",X"0E",X"E0",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",
		X"00",X"00",X"0E",X"0E",X"00",X"0D",X"E0",X"0E",X"00",X"DD",X"E0",X"0E",X"00",X"DD",X"00",X"0E",
		X"00",X"DD",X"00",X"0E",X"07",X"DD",X"00",X"EE",X"77",X"DD",X"00",X"EE",X"77",X"DD",X"DE",X"EE",
		X"33",X"34",X"00",X"BE",X"33",X"44",X"00",X"EE",X"33",X"44",X"44",X"BB",X"33",X"44",X"44",X"EE",
		X"33",X"44",X"44",X"BB",X"33",X"44",X"44",X"EB",X"33",X"44",X"00",X"EE",X"33",X"43",X"00",X"EE",
		X"33",X"33",X"00",X"EE",X"03",X"55",X"E0",X"EE",X"03",X"5F",X"0E",X"E0",X"AA",X"F5",X"00",X"E0",
		X"AA",X"B5",X"00",X"00",X"BB",X"B0",X"00",X"00",X"BA",X"B4",X"00",X"00",X"AB",X"A4",X"00",X"00",
		X"AB",X"B4",X"00",X"00",X"BB",X"44",X"EE",X"00",X"BB",X"44",X"44",X"00",X"BB",X"44",X"44",X"0B",
		X"BB",X"04",X"45",X"BB",X"BB",X"00",X"45",X"00",X"BB",X"00",X"45",X"00",X"00",X"00",X"45",X"00",
		X"00",X"40",X"05",X"BB",X"00",X"40",X"00",X"0B",X"00",X"40",X"00",X"00",X"00",X"40",X"00",X"B0",
		X"00",X"40",X"00",X"BB",X"00",X"40",X"00",X"0B",X"00",X"40",X"00",X"00",X"00",X"04",X"00",X"00",
		X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",
		X"DB",X"DD",X"00",X"00",X"DB",X"0D",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"70",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"70",X"00",
		X"00",X"EE",X"77",X"00",X"00",X"EE",X"77",X"00",X"00",X"00",X"E7",X"00",X"00",X"00",X"E7",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"77",X"EE",X"00",X"0E",X"77",X"7E",X"00",X"0E",X"77",X"7E",X"00",
		X"0E",X"77",X"77",X"00",X"77",X"77",X"77",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",
		X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"33",X"77",X"00",X"00",
		X"33",X"7E",X"00",X"00",X"33",X"70",X"EE",X"B0",X"33",X"30",X"00",X"00",X"33",X"3E",X"00",X"0B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"04",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"04",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"4F",X"40",X"00",X"00",X"FF",X"44",X"00",
		X"00",X"44",X"44",X"00",X"04",X"44",X"45",X"00",X"04",X"44",X"45",X"00",X"04",X"44",X"45",X"00",
		X"04",X"44",X"55",X"00",X"04",X"44",X"55",X"00",X"04",X"44",X"55",X"00",X"04",X"44",X"55",X"E0",
		X"00",X"44",X"55",X"E0",X"00",X"44",X"54",X"E0",X"00",X"45",X"50",X"0E",X"00",X"55",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"60",X"00",X"00",X"F6",X"66",X"00",
		X"00",X"FF",X"66",X"00",X"00",X"66",X"66",X"00",X"00",X"66",X"66",X"00",X"00",X"66",X"66",X"00",
		X"00",X"66",X"66",X"00",X"00",X"66",X"66",X"00",X"00",X"66",X"6D",X"00",X"00",X"66",X"DD",X"E0",
		X"00",X"66",X"DD",X"E0",X"00",X"66",X"D6",X"E0",X"00",X"DD",X"60",X"0E",X"00",X"DD",X"00",X"00",
		X"00",X"DD",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"CC",X"CC",X"00",X"00",X"AA",X"AA",X"00",X"00",X"AA",X"AA",X"00",
		X"00",X"CC",X"AA",X"00",X"0C",X"FF",X"AA",X"00",X"0C",X"FF",X"AA",X"00",X"CC",X"FF",X"AA",X"00",
		X"CA",X"CC",X"AA",X"00",X"CA",X"CC",X"AA",X"00",X"CA",X"CC",X"AA",X"00",X"CA",X"CC",X"AA",X"00",
		X"CA",X"FF",X"AA",X"00",X"CA",X"FF",X"AA",X"00",X"CA",X"FF",X"AA",X"00",X"CA",X"CC",X"AA",X"00",
		X"CC",X"CC",X"AA",X"00",X"0C",X"CC",X"AA",X"00",X"0C",X"CC",X"AA",X"00",X"00",X"AA",X"AA",X"00",
		X"00",X"AA",X"AA",X"00",X"00",X"AA",X"AA",X"00",X"00",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"CC",X"CC",X"00",X"00",X"66",X"66",X"00",X"00",X"66",X"66",X"00",
		X"00",X"CC",X"66",X"00",X"0C",X"FF",X"66",X"00",X"0C",X"FF",X"66",X"00",X"CC",X"FF",X"66",X"00",
		X"C6",X"CC",X"66",X"00",X"C6",X"CC",X"66",X"00",X"C6",X"CC",X"66",X"00",X"C6",X"CC",X"66",X"00",
		X"C6",X"FF",X"66",X"00",X"C6",X"FF",X"66",X"00",X"C6",X"FF",X"66",X"00",X"C6",X"CC",X"66",X"00",
		X"CC",X"CC",X"66",X"00",X"0C",X"CC",X"66",X"00",X"0C",X"CC",X"66",X"00",X"00",X"66",X"66",X"00",
		X"00",X"66",X"66",X"00",X"00",X"66",X"66",X"00",X"00",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"CC",X"CC",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",
		X"00",X"CC",X"BB",X"00",X"0C",X"FF",X"BB",X"00",X"0C",X"FF",X"BB",X"00",X"CC",X"FF",X"BB",X"00",
		X"CB",X"CC",X"BB",X"00",X"CB",X"CC",X"BB",X"00",X"CB",X"CC",X"BB",X"00",X"CB",X"CC",X"BB",X"00",
		X"CB",X"FF",X"BB",X"00",X"CB",X"FF",X"BB",X"00",X"CB",X"FF",X"BB",X"00",X"CB",X"CC",X"BB",X"00",
		X"CC",X"CC",X"BB",X"00",X"0C",X"CC",X"BB",X"00",X"0C",X"CC",X"BB",X"00",X"00",X"BB",X"BB",X"00",
		X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"00",X"00",
		X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AF",X"A0",X"00",X"00",X"FF",X"AA",X"00",
		X"00",X"FF",X"AA",X"00",X"0A",X"AA",X"AA",X"00",X"0A",X"AA",X"AA",X"00",X"0A",X"AA",X"AA",X"00",
		X"0A",X"AA",X"A9",X"00",X"0A",X"AA",X"99",X"00",X"0A",X"AA",X"99",X"00",X"0A",X"AA",X"99",X"E0",
		X"00",X"AA",X"99",X"E0",X"00",X"A9",X"9A",X"E0",X"00",X"99",X"A0",X"0E",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"A9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"70",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"50",X"00",
		X"00",X"40",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"0F",X"05",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",
		X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"04",X"00",
		X"00",X"00",X"40",X"00",X"00",X"0A",X"00",X"00",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0A",X"A0",X"00",X"00",X"AA",X"05",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",
		X"00",X"00",X"05",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",
		X"00",X"A0",X"00",X"00",X"00",X"0A",X"A0",X"00",X"00",X"0A",X"AA",X"00",X"00",X"50",X"A0",X"00",
		X"00",X"45",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",
		X"04",X"44",X"04",X"00",X"00",X"54",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"A0",X"40",X"05",X"00",X"0A",X"00",
		X"45",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"04",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"04",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"04",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"04",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"44",X"00",X"00",X"40",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"09",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"A9",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"A9",X"00",X"BB",X"99",X"99",X"00",
		X"00",X"99",X"A9",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"A9",X"00",X"00",X"99",X"99",X"00",X"00",X"09",X"99",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"40",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",
		X"00",X"60",X"AA",X"00",X"00",X"60",X"AA",X"00",X"00",X"60",X"66",X"00",X"00",X"60",X"00",X"00",
		X"00",X"60",X"00",X"00",X"00",X"66",X"06",X"00",X"00",X"AA",X"06",X"00",X"00",X"AA",X"06",X"00",
		X"00",X"66",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"60",X"A6",X"00",
		X"00",X"60",X"AA",X"00",X"00",X"60",X"AA",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",
		X"00",X"60",X"AA",X"00",X"00",X"60",X"AA",X"00",X"00",X"60",X"66",X"00",X"00",X"60",X"00",X"00",
		X"00",X"60",X"00",X"00",X"00",X"66",X"06",X"00",X"00",X"AA",X"06",X"00",X"00",X"AA",X"06",X"00",
		X"00",X"66",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"00",X"00",X"AA",X"AA",X"00",
		X"00",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"00",X"00",X"AA",X"AA",X"00",X"00",X"66",X"66",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"00",X"00",X"AA",X"AA",X"00",
		X"00",X"AA",X"AA",X"00",X"00",X"AA",X"66",X"00",X"00",X"AA",X"00",X"00",X"00",X"6A",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"60",X"AA",X"00",
		X"00",X"60",X"AA",X"00",X"00",X"60",X"66",X"00",X"00",X"60",X"00",X"00",X"00",X"60",X"00",X"00",
		X"00",X"66",X"06",X"00",X"00",X"AA",X"06",X"00",X"00",X"AA",X"06",X"00",X"00",X"66",X"06",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"00",X"00",X"AA",X"AA",X"00",
		X"00",X"AA",X"AA",X"00",X"00",X"AA",X"66",X"00",X"00",X"AA",X"00",X"00",X"00",X"6A",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",
		X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"66",X"60",X"00",X"00",X"60",X"66",X"00",
		X"00",X"60",X"A6",X"00",X"00",X"66",X"AA",X"00",X"00",X"A6",X"AA",X"00",X"00",X"A6",X"6A",X"00",
		X"00",X"66",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"66",X"00",X"00",X"06",X"6A",X"00",
		X"00",X"06",X"AA",X"00",X"00",X"06",X"A6",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"60",X"00",
		X"00",X"00",X"66",X"00",X"00",X"06",X"A6",X"00",X"00",X"06",X"AA",X"00",X"00",X"06",X"6A",X"00",
		X"00",X"06",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"00",
		X"00",X"AA",X"AA",X"00",X"00",X"AA",X"AA",X"00",X"00",X"66",X"66",X"00",X"00",X"60",X"00",X"00",
		X"00",X"60",X"00",X"00",X"00",X"66",X"06",X"00",X"00",X"A6",X"06",X"00",X"00",X"A6",X"06",X"00",
		X"00",X"66",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"66",X"00",X"00",X"06",X"6A",X"00",
		X"00",X"06",X"AA",X"00",X"00",X"06",X"A6",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"60",X"00",
		X"00",X"00",X"66",X"00",X"00",X"06",X"A6",X"00",X"00",X"06",X"AA",X"00",X"00",X"06",X"6A",X"00",
		X"00",X"06",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"00",X"00",X"AA",X"AA",X"00",X"00",X"AA",X"AA",X"00",
		X"00",X"00",X"66",X"00",X"00",X"A0",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"6A",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"66",X"00",X"00",X"06",X"6A",X"00",
		X"00",X"06",X"AA",X"00",X"00",X"06",X"A6",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"60",X"00",
		X"00",X"00",X"66",X"00",X"00",X"06",X"A6",X"00",X"00",X"06",X"AA",X"00",X"00",X"06",X"6A",X"00",
		X"00",X"06",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",
		X"00",X"60",X"AA",X"00",X"00",X"60",X"AA",X"00",X"00",X"60",X"66",X"00",X"00",X"60",X"00",X"00",
		X"00",X"60",X"00",X"00",X"00",X"66",X"06",X"00",X"00",X"AA",X"06",X"00",X"00",X"AA",X"06",X"00",
		X"00",X"66",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"66",X"00",X"00",X"06",X"6A",X"00",
		X"00",X"06",X"AA",X"00",X"00",X"06",X"A6",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"60",X"00",
		X"00",X"00",X"66",X"00",X"00",X"06",X"A6",X"00",X"00",X"06",X"AA",X"00",X"00",X"06",X"6A",X"00",
		X"00",X"06",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"CC",X"CC",X"00",X"00",X"55",X"55",X"00",X"00",X"55",X"55",X"00",
		X"00",X"CC",X"55",X"00",X"0C",X"FF",X"55",X"00",X"0C",X"FF",X"55",X"00",X"CC",X"FF",X"55",X"00",
		X"C5",X"CC",X"55",X"00",X"C5",X"CC",X"55",X"00",X"C5",X"CC",X"55",X"00",X"C5",X"CC",X"55",X"00",
		X"C5",X"FF",X"55",X"00",X"C5",X"FF",X"55",X"00",X"C5",X"FF",X"55",X"00",X"C5",X"CC",X"55",X"00",
		X"CC",X"CC",X"55",X"00",X"0C",X"CC",X"55",X"00",X"0C",X"CC",X"55",X"00",X"00",X"55",X"55",X"00",
		X"00",X"55",X"55",X"00",X"00",X"55",X"55",X"00",X"00",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"EE",X"EE",X"E0",X"EE",X"EE",X"00",X"E0",X"00",X"0E",X"00",X"E0",X"00",X"0E",X"00",X"E0",
		X"00",X"0E",X"00",X"E0",X"00",X"0E",X"00",X"E0",X"00",X"0E",X"00",X"E0",X"00",X"0E",X"E0",X"00",
		X"0E",X"0E",X"0E",X"00",X"E0",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"E0",X"0E",X"00",X"00",
		X"EE",X"0E",X"0E",X"00",X"EE",X"0E",X"EE",X"00",X"0E",X"0E",X"E0",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"0E",X"0E",X"E0",X"00",X"EE",X"0E",X"EE",X"00",X"EE",X"0E",X"0E",X"00",
		X"E0",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"E0",X"0E",X"00",X"00",X"0E",X"0E",X"0E",X"00",
		X"00",X"0E",X"E0",X"00",X"00",X"0E",X"00",X"E0",X"00",X"0E",X"00",X"E0",X"00",X"0E",X"00",X"E0",
		X"00",X"0E",X"00",X"E0",X"00",X"0E",X"00",X"E0",X"EE",X"EE",X"00",X"E0",X"EE",X"EE",X"00",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"0E",X"0E",X"E0",X"00",X"EE",X"0E",X"EE",X"00",X"EE",X"0E",X"0E",X"00",
		X"E0",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"E0",X"0E",X"00",X"00",X"DD",X"0E",X"0E",X"00",
		X"DD",X"0E",X"E0",X"00",X"DD",X"0E",X"00",X"E0",X"DD",X"0E",X"00",X"E0",X"DD",X"0E",X"00",X"E0",
		X"D0",X"0E",X"00",X"E0",X"D0",X"0E",X"00",X"E0",X"D2",X"EE",X"00",X"E0",X"D2",X"EE",X"EE",X"E0",
		X"44",X"4F",X"77",X"77",X"44",X"4F",X"77",X"77",X"44",X"4F",X"77",X"77",X"44",X"4F",X"77",X"77",
		X"44",X"4F",X"77",X"77",X"44",X"4F",X"77",X"77",X"44",X"4F",X"77",X"77",X"44",X"40",X"77",X"00",
		X"40",X"40",X"77",X"00",X"00",X"40",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"3F",X"77",X"22",X"43",X"3F",X"77",X"22",X"43",X"3F",X"77",X"22",X"44",X"3F",X"77",X"22",
		X"44",X"3F",X"77",X"22",X"44",X"3F",X"77",X"00",X"44",X"3F",X"77",X"00",X"44",X"00",X"70",X"00",
		X"44",X"00",X"BB",X"00",X"44",X"00",X"B0",X"00",X"44",X"45",X"00",X"00",X"44",X"4F",X"00",X"00",
		X"44",X"55",X"BB",X"00",X"44",X"55",X"BB",X"00",X"44",X"4F",X"00",X"00",X"44",X"05",X"00",X"00",
		X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"3B",X"77",X"77",X"33",X"3B",X"77",X"77",X"43",X"3B",X"77",X"77",X"43",X"BB",X"77",X"77",
		X"44",X"BB",X"77",X"22",X"44",X"FB",X"77",X"00",X"44",X"5B",X"77",X"00",X"44",X"F0",X"77",X"00",
		X"44",X"50",X"70",X"00",X"44",X"00",X"70",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",
		X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"B0",X"00",X"00",X"4B",X"B0",
		X"00",X"00",X"4B",X"BB",X"00",X"00",X"4B",X"BB",X"00",X"00",X"4B",X"BB",X"00",X"00",X"4B",X"BB",
		X"00",X"00",X"4B",X"BB",X"00",X"00",X"4B",X"00",X"00",X"00",X"4B",X"00",X"00",X"00",X"40",X"00",
		X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"BB",X"00",X"00",X"40",X"BB",X"00",X"00",X"40",X"7B",
		X"00",X"00",X"4B",X"BB",X"00",X"00",X"4B",X"BB",X"00",X"00",X"4B",X"BB",X"00",X"00",X"4B",X"AB",
		X"00",X"00",X"4B",X"A0",X"00",X"00",X"4B",X"A0",X"00",X"00",X"4B",X"A0",X"00",X"00",X"4B",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",
		X"00",X"00",X"4B",X"00",X"00",X"00",X"4B",X"A0",X"00",X"00",X"4B",X"AB",X"00",X"00",X"4B",X"BB",
		X"00",X"00",X"4A",X"BB",X"00",X"00",X"4A",X"BB",X"00",X"00",X"4A",X"00",X"00",X"00",X"4A",X"00",
		X"00",X"00",X"4A",X"00",X"00",X"00",X"4A",X"00",X"00",X"00",X"4A",X"00",X"00",X"00",X"AA",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",
		X"00",X"00",X"11",X"10",X"00",X"00",X"11",X"10",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",
		X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",
		X"00",X"00",X"77",X"11",X"00",X"3F",X"77",X"11",X"00",X"3F",X"77",X"77",X"00",X"3F",X"77",X"77",
		X"50",X"3F",X"77",X"77",X"55",X"3F",X"77",X"77",X"33",X"3F",X"77",X"77",X"33",X"3F",X"77",X"77",
		X"00",X"00",X"DD",X"00",X"00",X"0D",X"DD",X"00",X"00",X"DD",X"DD",X"07",X"00",X"DD",X"DD",X"00",
		X"00",X"DD",X"DD",X"00",X"00",X"DD",X"77",X"00",X"00",X"0D",X"77",X"00",X"00",X"00",X"77",X"00",
		X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",
		X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",
		X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",
		X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"B0",X"B0",X"77",X"00",X"BB",X"00",X"77",X"70",
		X"2B",X"00",X"77",X"77",X"0B",X"00",X"77",X"77",X"BB",X"00",X"77",X"77",X"BB",X"00",X"77",X"77",
		X"BB",X"00",X"77",X"77",X"25",X"00",X"77",X"77",X"25",X"00",X"77",X"77",X"25",X"00",X"77",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"EE",X"EE",X"E0",X"EE",X"EE",X"00",X"E0",X"00",X"0E",X"00",X"E0",X"00",X"0E",X"00",X"E0",
		X"00",X"0E",X"00",X"E0",X"00",X"0E",X"00",X"E0",X"00",X"0E",X"00",X"E0",X"00",X"0E",X"E0",X"00",
		X"0E",X"0E",X"0E",X"00",X"E0",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"E0",X"0E",X"00",X"00",
		X"EE",X"0E",X"0E",X"00",X"EE",X"0E",X"EE",X"00",X"0E",X"0E",X"E0",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DE",X"EE",X"22",X"E0",X"DD",X"EE",X"22",X"E0",X"DD",X"0E",X"00",X"E0",X"77",X"5E",X"00",X"E0",
		X"00",X"0E",X"00",X"E0",X"00",X"0E",X"00",X"E0",X"00",X"0E",X"E0",X"E0",X"00",X"0E",X"0E",X"00",
		X"0E",X"0E",X"00",X"00",X"E0",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"E0",X"0E",X"00",X"00",
		X"EE",X"0E",X"0E",X"00",X"EE",X"0E",X"EE",X"00",X"00",X"0E",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"EE",X"EE",X"E0",X"7E",X"88",X"00",X"E0",X"00",X"88",X"00",X"E0",X"00",X"80",X"00",X"E0",
		X"00",X"22",X"00",X"E0",X"00",X"22",X"00",X"E0",X"0E",X"22",X"00",X"E0",X"E0",X"22",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"0E",X"00",
		X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",
		X"EE",X"00",X"0E",X"00",X"EE",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",
		X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"70",X"BB",X"00",X"77",X"70",
		X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",
		X"50",X"00",X"77",X"77",X"55",X"3F",X"77",X"77",X"33",X"3F",X"77",X"77",X"33",X"3F",X"77",X"77",
		X"33",X"4F",X"77",X"77",X"33",X"4F",X"77",X"77",X"33",X"44",X"77",X"27",X"34",X"44",X"77",X"27",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"B0",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"05",X"00",X"11",X"00",X"04",X"00",X"11",
		X"00",X"44",X"00",X"11",X"00",X"44",X"00",X"11",X"00",X"44",X"77",X"11",X"00",X"44",X"77",X"11",
		X"50",X"44",X"77",X"11",X"55",X"B3",X"77",X"11",X"33",X"B3",X"77",X"00",X"33",X"B3",X"77",X"00",
		X"33",X"F5",X"77",X"77",X"33",X"F5",X"77",X"77",X"33",X"F5",X"77",X"77",X"33",X"44",X"77",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0B",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"01",X"00",
		X"BB",X"00",X"11",X"00",X"BB",X"00",X"11",X"00",X"BB",X"00",X"11",X"00",X"BB",X"00",X"11",X"00",
		X"BB",X"00",X"11",X"00",X"BB",X"00",X"11",X"10",X"05",X"00",X"11",X"11",X"00",X"00",X"11",X"11",
		X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"40",X"71",X"11",X"00",X"44",X"77",X"11",
		X"50",X"44",X"77",X"11",X"55",X"3F",X"77",X"77",X"33",X"3F",X"77",X"77",X"33",X"3F",X"77",X"77",
		X"33",X"3F",X"77",X"77",X"33",X"3F",X"77",X"77",X"33",X"3F",X"77",X"77",X"33",X"3F",X"77",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"B0",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"40",X"00",X"77",
		X"00",X"40",X"00",X"77",X"00",X"40",X"00",X"77",X"00",X"40",X"00",X"77",X"00",X"40",X"00",X"77",
		X"00",X"40",X"00",X"77",X"00",X"40",X"00",X"77",X"00",X"40",X"00",X"77",X"00",X"30",X"77",X"77",
		X"50",X"3F",X"77",X"77",X"55",X"3F",X"77",X"77",X"33",X"3F",X"77",X"77",X"33",X"3F",X"77",X"77",
		X"33",X"3F",X"77",X"77",X"33",X"3F",X"77",X"22",X"33",X"3F",X"77",X"22",X"33",X"3F",X"77",X"27",
		X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"0D",X"DD",X"DD",X"00",X"0D",X"DD",X"DD",
		X"00",X"DD",X"DD",X"D0",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",
		X"00",X"DD",X"D0",X"00",X"00",X"0D",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"07",
		X"00",X"00",X"BB",X"77",X"00",X"00",X"B0",X"77",X"00",X"00",X"B0",X"77",X"00",X"05",X"00",X"77",
		X"00",X"0F",X"00",X"77",X"00",X"44",X"00",X"77",X"00",X"44",X"00",X"77",X"00",X"44",X"00",X"77",
		X"00",X"44",X"00",X"77",X"04",X"44",X"00",X"77",X"44",X"40",X"00",X"70",X"44",X"00",X"07",X"70",
		X"44",X"00",X"77",X"70",X"44",X"00",X"77",X"00",X"44",X"00",X"77",X"00",X"44",X"00",X"77",X"00",
		X"44",X"33",X"77",X"00",X"33",X"33",X"77",X"00",X"53",X"33",X"77",X"0E",X"55",X"33",X"77",X"EE",
		X"55",X"33",X"77",X"EE",X"53",X"33",X"77",X"EE",X"33",X"33",X"77",X"00",X"44",X"33",X"77",X"10",
		X"44",X"33",X"77",X"10",X"44",X"00",X"71",X"11",X"44",X"00",X"11",X"11",X"44",X"00",X"11",X"11",
		X"44",X"00",X"01",X"11",X"44",X"40",X"00",X"11",X"04",X"44",X"00",X"11",X"00",X"44",X"00",X"11",
		X"00",X"44",X"00",X"11",X"00",X"44",X"00",X"11",X"00",X"44",X"00",X"11",X"05",X"40",X"00",X"11",
		X"BB",X"40",X"00",X"11",X"BB",X"00",X"00",X"11",X"BB",X"00",X"11",X"11",X"BB",X"00",X"11",X"10",
		X"B0",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"10",X"DD",
		X"00",X"00",X"00",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"0D",X"DD",X"DD",X"00",X"0D",X"DD",X"DD",
		X"00",X"0D",X"DD",X"DD",X"00",X"0D",X"DD",X"DD",X"00",X"0D",X"DD",X"DD",X"00",X"0D",X"00",X"DD",
		X"77",X"55",X"20",X"E0",X"77",X"FF",X"20",X"E0",X"77",X"55",X"E0",X"E0",X"77",X"00",X"0E",X"E0",
		X"EE",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",
		X"0E",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"E0",X"00",
		X"EE",X"00",X"EE",X"00",X"EE",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"5F",X"DD",X"00",X"E0",X"35",X"DD",X"00",X"E0",X"30",X"DE",X"00",X"E0",X"00",X"2E",X"00",X"E0",
		X"00",X"2E",X"00",X"E0",X"00",X"2E",X"EE",X"E0",X"00",X"20",X"00",X"E0",X"00",X"00",X"00",X"00",
		X"0E",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",
		X"EE",X"00",X"EE",X"00",X"EE",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"EE",X"00",X"EE",X"00",X"EE",X"00",
		X"E0",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"88",X"00",X"00",
		X"00",X"88",X"00",X"00",X"00",X"88",X"00",X"00",X"E0",X"88",X"00",X"00",X"7E",X"08",X"00",X"00",
		X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"E0",X"77",X"0E",X"EE",X"E0",X"77",X"0E",X"00",X"E0",
		X"75",X"0D",X"00",X"E0",X"75",X"DD",X"00",X"E0",X"7F",X"DD",X"00",X"E0",X"5F",X"DD",X"00",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"EE",X"00",X"EE",X"00",X"0E",X"00",
		X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"0E",X"00",
		X"00",X"DD",X"0E",X"00",X"00",X"DD",X"E0",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",
		X"E0",X"2D",X"00",X"00",X"7E",X"2D",X"00",X"E0",X"77",X"25",X"00",X"E0",X"77",X"55",X"00",X"E0",
		X"77",X"5F",X"00",X"E0",X"77",X"FF",X"00",X"E0",X"77",X"75",X"00",X"E0",X"77",X"77",X"00",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"EE",X"00",X"EE",X"00",X"EE",X"00",
		X"E0",X"00",X"E0",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",
		X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",
		X"08",X"00",X"00",X"00",X"08",X"00",X"D0",X"E0",X"08",X"00",X"D0",X"E0",X"EE",X"00",X"D0",X"E0",
		X"77",X"00",X"0E",X"E0",X"77",X"55",X"E0",X"E0",X"77",X"FF",X"20",X"E0",X"77",X"55",X"20",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"B0",
		X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"40",
		X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",
		X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",
		X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"44",
		X"00",X"00",X"00",X"44",X"00",X"00",X"55",X"44",X"00",X"0B",X"55",X"44",X"00",X"BB",X"FF",X"44",
		X"00",X"B0",X"55",X"44",X"00",X"00",X"55",X"44",X"00",X"00",X"50",X"44",X"00",X"00",X"00",X"44",
		X"00",X"00",X"4B",X"AB",X"00",X"00",X"4B",X"BB",X"00",X"00",X"4B",X"B0",X"00",X"00",X"4B",X"00",
		X"00",X"00",X"40",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"40",X"00",
		X"00",X"00",X"4B",X"00",X"00",X"00",X"4B",X"B0",X"00",X"00",X"4B",X"BB",X"00",X"00",X"4B",X"AB",
		X"55",X"3F",X"77",X"77",X"35",X"3F",X"77",X"77",X"33",X"3F",X"77",X"77",X"33",X"3F",X"77",X"77",
		X"43",X"3F",X"77",X"00",X"44",X"3F",X"77",X"00",X"44",X"00",X"77",X"00",X"44",X"00",X"77",X"00",
		X"44",X"00",X"70",X"00",X"44",X"00",X"70",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",
		X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"04",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"04",X"00",X"00",X"00",
		X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",
		X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",
		X"B0",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",
		X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",
		X"F5",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",
		X"04",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",
		X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",
		X"44",X"00",X"70",X"00",X"44",X"00",X"77",X"00",X"44",X"3F",X"77",X"00",X"43",X"3F",X"77",X"77",
		X"33",X"3F",X"77",X"77",X"33",X"3F",X"77",X"77",X"35",X"3F",X"77",X"77",X"55",X"3F",X"77",X"77",
		X"44",X"4F",X"77",X"22",X"44",X"3F",X"77",X"22",X"44",X"3F",X"77",X"22",X"44",X"3F",X"77",X"22",
		X"44",X"3F",X"77",X"22",X"44",X"3F",X"77",X"00",X"44",X"3F",X"77",X"00",X"44",X"40",X"77",X"00",
		X"40",X"40",X"70",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"44",X"40",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"40",X"00",
		X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"24",X"00",X"77",X"77",X"24",X"00",X"77",X"77",X"24",X"00",X"77",X"77",X"24",X"00",X"77",X"77",
		X"24",X"00",X"77",X"77",X"24",X"00",X"F7",X"77",X"24",X"03",X"F7",X"77",X"24",X"03",X"F7",X"77",
		X"24",X"33",X"F7",X"77",X"24",X"33",X"F7",X"07",X"24",X"33",X"F7",X"07",X"24",X"33",X"F7",X"00",
		X"04",X"33",X"F7",X"00",X"04",X"33",X"30",X"00",X"44",X"33",X"30",X"00",X"44",X"53",X"00",X"00",
		X"44",X"55",X"00",X"00",X"43",X"53",X"00",X"00",X"43",X"33",X"00",X"00",X"43",X"33",X"00",X"00",
		X"43",X"33",X"00",X"00",X"BB",X"33",X"44",X"44",X"BB",X"34",X"44",X"44",X"6B",X"34",X"44",X"44",
		X"BB",X"44",X"44",X"44",X"6A",X"44",X"44",X"00",X"AA",X"44",X"40",X"00",X"AA",X"44",X"00",X"00",
		X"AA",X"04",X"00",X"00",X"4A",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"DD",X"00",X"00",X"77",X"0D",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",
		X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"E0",X"EE",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"EE",X"00",X"00",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",
		X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"EE",X"00",X"00",X"EE",X"EE",X"00",
		X"00",X"E0",X"EE",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",
		X"EE",X"00",X"00",X"00",X"E0",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"EE",
		X"E0",X"00",X"00",X"EE",X"0E",X"00",X"0E",X"EE",X"00",X"00",X"0E",X"EE",X"00",X"00",X"E0",X"EE",
		X"00",X"00",X"00",X"E0",X"00",X"D0",X"00",X"E0",X"00",X"DD",X"00",X"E0",X"00",X"DD",X"00",X"00",
		X"00",X"DD",X"00",X"00",X"77",X"DD",X"00",X"00",X"77",X"DD",X"00",X"00",X"75",X"DD",X"EE",X"00",
		X"33",X"44",X"00",X"00",X"33",X"44",X"44",X"BB",X"34",X"44",X"44",X"00",X"34",X"44",X"44",X"00",
		X"44",X"44",X"44",X"00",X"44",X"44",X"00",X"B0",X"44",X"44",X"00",X"BB",X"44",X"00",X"00",X"00",
		X"34",X"00",X"00",X"00",X"33",X"50",X"00",X"00",X"33",X"50",X"00",X"00",X"A3",X"00",X"E0",X"00",
		X"AB",X"00",X"0E",X"00",X"BB",X"00",X"00",X"00",X"BB",X"40",X"00",X"00",X"BB",X"44",X"00",X"00",
		X"66",X"44",X"00",X"00",X"66",X"44",X"EE",X"00",X"BB",X"44",X"5E",X"00",X"BB",X"44",X"55",X"00",
		X"BB",X"44",X"FF",X"00",X"BB",X"44",X"55",X"00",X"BB",X"00",X"5F",X"00",X"00",X"00",X"F5",X"00",
		X"00",X"00",X"F5",X"00",X"00",X"00",X"55",X"B0",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",X"DD",X"DD",X"00",X"00",
		X"BB",X"DD",X"00",X"00",X"BB",X"DD",X"00",X"00",X"B5",X"00",X"00",X"00",X"55",X"00",X"00",X"00",
		X"55",X"00",X"00",X"00",X"0F",X"77",X"00",X"00",X"05",X"77",X"00",X"00",X"00",X"77",X"00",X"00",
		X"00",X"EE",X"77",X"00",X"00",X"EE",X"77",X"00",X"0E",X"00",X"77",X"00",X"0E",X"00",X"77",X"00",
		X"EE",X"77",X"77",X"00",X"E0",X"77",X"77",X"00",X"E0",X"77",X"E7",X"00",X"E0",X"77",X"EE",X"00",
		X"E7",X"77",X"EE",X"00",X"77",X"77",X"EE",X"00",X"77",X"77",X"0E",X"00",X"77",X"7E",X"00",X"00",
		X"77",X"7E",X"00",X"00",X"77",X"E0",X"00",X"00",X"77",X"E0",X"00",X"00",X"33",X"00",X"00",X"00",
		X"33",X"00",X"EE",X"00",X"33",X"00",X"00",X"0B",X"33",X"00",X"00",X"B0",X"33",X"EE",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"44",X"40",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"40",X"00",
		X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"04",X"FF",X"00",X"00",X"44",X"FF",X"00",X"00",
		X"44",X"44",X"00",X"00",X"FF",X"44",X"50",X"00",X"44",X"44",X"50",X"00",X"44",X"44",X"55",X"00",
		X"44",X"44",X"55",X"00",X"44",X"44",X"55",X"00",X"44",X"44",X"50",X"00",X"44",X"44",X"40",X"00",
		X"44",X"44",X"00",X"00",X"54",X"45",X"00",X"00",X"05",X"55",X"00",X"00",X"00",X"55",X"00",X"E0",
		X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"06",X"66",X"00",X"00",X"06",X"66",X"00",X"00",
		X"66",X"66",X"00",X"00",X"66",X"66",X"60",X"00",X"66",X"66",X"60",X"00",X"6F",X"66",X"66",X"00",
		X"66",X"66",X"66",X"00",X"66",X"66",X"DD",X"00",X"66",X"66",X"D0",X"00",X"66",X"66",X"60",X"00",
		X"86",X"66",X"00",X"00",X"06",X"6D",X"00",X"00",X"08",X"DD",X"00",X"00",X"00",X"DD",X"00",X"E0",
		X"00",X"DD",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"CC",X"CC",X"00",X"00",X"AA",X"AA",X"00",X"0C",X"AA",X"AA",X"00",
		X"CC",X"CC",X"AA",X"00",X"CA",X"FF",X"CC",X"00",X"AA",X"FF",X"CC",X"00",X"AA",X"CC",X"AA",X"00",
		X"AA",X"CC",X"AA",X"00",X"AA",X"CC",X"AA",X"00",X"AA",X"CC",X"AA",X"00",X"AA",X"CC",X"CC",X"00",
		X"AA",X"FF",X"CC",X"00",X"AA",X"FF",X"AA",X"00",X"AA",X"CC",X"AA",X"00",X"AA",X"CC",X"AA",X"00",
		X"AA",X"CC",X"AA",X"00",X"AA",X"CC",X"CC",X"00",X"CA",X"CC",X"CC",X"00",X"CC",X"AA",X"AA",X"00",
		X"0C",X"AA",X"AA",X"00",X"00",X"AA",X"AA",X"00",X"00",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"CC",X"CC",X"00",X"00",X"66",X"66",X"00",X"0C",X"66",X"66",X"00",
		X"CC",X"CC",X"66",X"00",X"C6",X"FF",X"CC",X"00",X"66",X"FF",X"CC",X"00",X"66",X"CC",X"66",X"00",
		X"66",X"CC",X"66",X"00",X"66",X"CC",X"66",X"00",X"66",X"CC",X"66",X"00",X"66",X"CC",X"CC",X"00",
		X"66",X"FF",X"CC",X"00",X"66",X"FF",X"66",X"00",X"66",X"CC",X"66",X"00",X"66",X"CC",X"66",X"00",
		X"66",X"CC",X"66",X"00",X"66",X"CC",X"CC",X"00",X"C6",X"CC",X"CC",X"00",X"CC",X"66",X"66",X"00",
		X"0C",X"66",X"66",X"00",X"00",X"66",X"66",X"00",X"00",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"CC",X"CC",X"00",X"00",X"BB",X"BB",X"00",X"0C",X"BB",X"BB",X"00",
		X"CC",X"CC",X"BB",X"00",X"CB",X"FF",X"CC",X"00",X"BB",X"FF",X"CC",X"00",X"BB",X"CC",X"BB",X"00",
		X"BB",X"CC",X"BB",X"00",X"BB",X"CC",X"BB",X"00",X"BB",X"CC",X"BB",X"00",X"BB",X"CC",X"CC",X"00",
		X"BB",X"FF",X"CC",X"00",X"BB",X"FF",X"BB",X"00",X"BB",X"CC",X"BB",X"00",X"BB",X"CC",X"BB",X"00",
		X"BB",X"CC",X"BB",X"00",X"BB",X"CC",X"CC",X"00",X"CB",X"CC",X"CC",X"00",X"CC",X"BB",X"BB",X"00",
		X"0C",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"00",X"00",
		X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"0A",X"FF",X"00",X"00",X"AA",X"FF",X"00",X"00",
		X"AA",X"FA",X"00",X"00",X"AF",X"AA",X"A0",X"00",X"FF",X"AA",X"A0",X"00",X"AA",X"AA",X"9A",X"00",
		X"AA",X"AA",X"AA",X"00",X"AA",X"AA",X"9A",X"00",X"AA",X"AA",X"90",X"00",X"AA",X"AA",X"A0",X"00",
		X"AA",X"A9",X"00",X"00",X"AA",X"99",X"00",X"00",X"0A",X"99",X"00",X"00",X"00",X"99",X"00",X"E0",
		X"00",X"99",X"00",X"00",X"00",X"A9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"0A",X"05",X"00",
		X"00",X"70",X"50",X"00",X"00",X"4A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"06",X"55",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"40",X"A0",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"04",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"66",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"A6",X"00",X"00",X"00",X"F6",X"00",X"00",X"0F",X"F6",X"00",X"00",
		X"00",X"FA",X"00",X"00",X"00",X"0A",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",
		X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"04",X"00",X"F5",X"04",X"40",X"00",X"00",X"04",X"00",X"00",X"00",X"A4",X"00",X"00",
		X"00",X"A4",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"6A",X"00",X"00",X"00",X"F6",X"00",X"00",
		X"04",X"46",X"00",X"00",X"00",X"66",X"44",X"00",X"00",X"04",X"00",X"00",X"00",X"05",X"00",X"00",
		X"00",X"05",X"00",X"00",X"05",X"00",X"00",X"00",X"55",X"50",X"00",X"00",X"0A",X"50",X"00",X"00",
		X"0A",X"50",X"A0",X"00",X"0A",X"40",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"44",X"40",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"04",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"04",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"40",X"00",
		X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"04",X"00",X"44",X"00",
		X"04",X"00",X"44",X"00",X"04",X"40",X"44",X"00",X"04",X"40",X"44",X"00",X"04",X"40",X"44",X"00",
		X"04",X"44",X"44",X"00",X"04",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"40",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"99",X"00",X"00",X"9A",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"09",X"9A",X"99",X"00",X"B9",X"99",X"99",X"00",
		X"09",X"9A",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"9A",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"90",X"00",
		X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"04",X"00",X"44",X"00",
		X"04",X"00",X"44",X"00",X"04",X"00",X"44",X"00",X"04",X"44",X"44",X"00",X"04",X"44",X"44",X"00",
		X"04",X"44",X"44",X"00",X"04",X"44",X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"00",
		X"00",X"44",X"40",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"66",X"00",
		X"00",X"66",X"AA",X"00",X"00",X"6A",X"AA",X"00",X"00",X"6A",X"6A",X"00",X"00",X"6A",X"6A",X"00",
		X"00",X"6A",X"6A",X"00",X"00",X"6A",X"6A",X"00",X"00",X"AA",X"AA",X"00",X"00",X"AA",X"AA",X"00",
		X"00",X"66",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"66",X"06",X"00",X"00",X"AA",X"6A",X"00",X"00",X"AA",X"6A",X"00",
		X"00",X"66",X"6A",X"00",X"00",X"06",X"6A",X"00",X"00",X"06",X"6A",X"00",X"00",X"00",X"6A",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"66",X"00",
		X"00",X"66",X"AA",X"00",X"00",X"6A",X"AA",X"00",X"00",X"6A",X"6A",X"00",X"00",X"6A",X"6A",X"00",
		X"00",X"6A",X"6A",X"00",X"00",X"6A",X"6A",X"00",X"00",X"AA",X"AA",X"00",X"00",X"AA",X"AA",X"00",
		X"00",X"66",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"00",X"00",X"AA",X"AA",X"00",
		X"00",X"AA",X"AA",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"0A",X"00",
		X"00",X"00",X"0A",X"00",X"00",X"AA",X"AA",X"00",X"00",X"AA",X"AA",X"00",X"00",X"66",X"66",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"6A",X"00",X"00",X"66",X"6A",X"00",X"00",X"AA",X"AA",X"00",
		X"00",X"AA",X"AA",X"00",X"00",X"66",X"6A",X"00",X"00",X"A6",X"6A",X"00",X"00",X"A6",X"66",X"00",
		X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"66",X"00",X"00",X"66",X"AA",X"00",
		X"00",X"6A",X"AA",X"00",X"00",X"6A",X"6A",X"00",X"00",X"6A",X"6A",X"00",X"00",X"6A",X"6A",X"00",
		X"00",X"6A",X"6A",X"00",X"00",X"AA",X"AA",X"00",X"00",X"AA",X"AA",X"00",X"00",X"66",X"66",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"6A",X"00",X"00",X"66",X"6A",X"00",X"00",X"AA",X"AA",X"00",
		X"00",X"AA",X"AA",X"00",X"00",X"66",X"6A",X"00",X"00",X"A6",X"6A",X"00",X"00",X"A6",X"66",X"00",
		X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"00",
		X"00",X"AA",X"6A",X"00",X"00",X"AA",X"6A",X"00",X"00",X"66",X"6A",X"00",X"00",X"06",X"6A",X"00",
		X"00",X"00",X"6A",X"00",X"00",X"00",X"6A",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"60",X"00",X"00",X"A6",X"60",X"00",
		X"00",X"AA",X"60",X"00",X"00",X"6A",X"60",X"00",X"00",X"66",X"00",X"00",X"00",X"06",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"6A",X"60",X"00",X"00",X"AA",X"60",X"00",X"00",X"A6",X"60",X"00",
		X"00",X"66",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"00",
		X"00",X"AA",X"AA",X"00",X"00",X"AA",X"AA",X"00",X"00",X"66",X"6A",X"00",X"00",X"06",X"6A",X"00",
		X"00",X"06",X"6A",X"00",X"00",X"06",X"6A",X"00",X"00",X"06",X"AA",X"00",X"00",X"00",X"AA",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"60",X"00",X"00",X"A6",X"60",X"00",
		X"00",X"AA",X"60",X"00",X"00",X"6A",X"60",X"00",X"00",X"66",X"00",X"00",X"00",X"06",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"6A",X"60",X"00",X"00",X"AA",X"60",X"00",X"00",X"A6",X"60",X"00",
		X"00",X"66",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"06",X"66",X"66",X"00",X"06",X"AA",X"AA",X"00",X"06",X"AA",X"AA",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",
		X"00",X"AA",X"00",X"00",X"00",X"6A",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"06",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"60",X"00",X"00",X"A6",X"60",X"00",
		X"00",X"AA",X"60",X"00",X"00",X"6A",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"06",X"00",X"00",
		X"00",X"06",X"00",X"00",X"00",X"6A",X"60",X"00",X"00",X"AA",X"60",X"00",X"00",X"A6",X"60",X"00",
		X"00",X"66",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"66",X"00",
		X"00",X"66",X"AA",X"00",X"00",X"6A",X"AA",X"00",X"00",X"6A",X"6A",X"00",X"00",X"6A",X"6A",X"00",
		X"00",X"6A",X"6A",X"00",X"00",X"6A",X"6A",X"00",X"00",X"AA",X"AA",X"00",X"00",X"AA",X"AA",X"00",
		X"00",X"66",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"60",X"00",X"00",X"A6",X"60",X"00",
		X"00",X"AA",X"60",X"00",X"00",X"6A",X"60",X"00",X"00",X"66",X"00",X"00",X"00",X"06",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"6A",X"60",X"00",X"00",X"AA",X"60",X"00",X"00",X"A6",X"60",X"00",
		X"00",X"66",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"CC",X"CC",X"00",X"00",X"55",X"55",X"00",X"0C",X"55",X"55",X"00",
		X"CC",X"CC",X"55",X"00",X"C5",X"FF",X"CC",X"00",X"55",X"FF",X"CC",X"00",X"55",X"CC",X"55",X"00",
		X"55",X"CC",X"55",X"00",X"55",X"CC",X"55",X"00",X"55",X"CC",X"55",X"00",X"55",X"CC",X"CC",X"00",
		X"55",X"FF",X"CC",X"00",X"55",X"FF",X"55",X"00",X"55",X"CC",X"55",X"00",X"55",X"CC",X"55",X"00",
		X"55",X"CC",X"55",X"00",X"55",X"CC",X"CC",X"00",X"C5",X"CC",X"CC",X"00",X"CC",X"55",X"55",X"00",
		X"0C",X"55",X"55",X"00",X"00",X"55",X"55",X"00",X"00",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
