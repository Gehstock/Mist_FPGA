library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity tropical_spr_bit3 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of tropical_spr_bit3 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"07",X"0F",X"0F",X"07",X"06",X"02",X"00",X"00",X"00",X"00",X"01",X"0F",X"3F",X"7F",X"7F",
		X"E0",X"E0",X"F0",X"F0",X"F0",X"70",X"70",X"30",X"00",X"00",X"40",X"C0",X"F0",X"FC",X"FE",X"FE",
		X"7F",X"3F",X"0F",X"07",X"0E",X"00",X"02",X"00",X"00",X"00",X"08",X"5E",X"4F",X"4F",X"67",X"30",
		X"7E",X"7F",X"7D",X"70",X"70",X"00",X"F0",X"30",X"38",X"18",X"18",X"38",X"38",X"38",X"30",X"40",
		X"0E",X"06",X"06",X"06",X"03",X"03",X"01",X"01",X"01",X"01",X"01",X"03",X"03",X"03",X"01",X"01",
		X"20",X"20",X"20",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"70",X"30",X"30",X"30",X"F0",X"F0",
		X"00",X"00",X"00",X"03",X"07",X"0F",X"0F",X"0C",X"08",X"00",X"00",X"00",X"00",X"00",X"01",X"07",
		X"00",X"00",X"00",X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"60",X"60",X"00",X"C0",X"FC",X"FE",
		X"FF",X"FF",X"FF",X"EF",X"EF",X"EF",X"67",X"76",X"7F",X"37",X"37",X"1B",X"0B",X"01",X"00",X"00",
		X"F0",X"F8",X"F8",X"DC",X"8C",X"8E",X"86",X"00",X"C0",X"C0",X"C0",X"C0",X"E0",X"E0",X"70",X"F0",
		X"F1",X"03",X"01",X"21",X"78",X"7C",X"7C",X"3C",X"0C",X"06",X"02",X"03",X"07",X"07",X"0B",X"0B",
		X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"40",X"40",X"C0",X"C0",
		X"0F",X"1F",X"3F",X"3F",X"2F",X"07",X"07",X"03",X"01",X"00",X"03",X"07",X"0F",X"1F",X"3F",X"3B",
		X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"00",X"00",X"E0",X"F8",X"FC",X"FE",X"FE",
		X"7F",X"7E",X"3D",X"BD",X"BF",X"80",X"3C",X"BF",X"BF",X"BF",X"5F",X"07",X"07",X"27",X"27",X"33",
		X"60",X"36",X"37",X"18",X"18",X"00",X"00",X"00",X"C0",X"E0",X"E0",X"E0",X"EC",X"CC",X"CE",X"8E",
		X"E0",X"F0",X"F8",X"FC",X"7C",X"3C",X"0E",X"0E",X"0E",X"CF",X"CF",X"E7",X"73",X"39",X"1B",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"C0",
		X"00",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"F8",X"FC",X"FC",X"FC",X"FC",X"7C",X"38",X"18",X"00",X"10",X"7F",X"7F",X"7F",X"FF",X"DF",
		X"80",X"C0",X"E0",X"F0",X"F0",X"B9",X"1F",X"4F",X"E6",X"00",X"FE",X"FF",X"FF",X"5F",X"06",X"1E",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"F8",X"40",X"00",X"00",X"00",X"00",X"00",X"70",X"78",X"7C",
		X"60",X"F8",X"FC",X"FC",X"FE",X"3E",X"3F",X"1F",X"0F",X"07",X"83",X"D0",X"EC",X"3F",X"3F",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"60",X"E0",X"F0",X"F0",
		X"00",X"00",X"00",X"07",X"07",X"0F",X"0F",X"0F",X"0E",X"0C",X"00",X"00",X"00",X"00",X"38",X"7F",
		X"00",X"00",X"00",X"C0",X"E0",X"F0",X"F0",X"30",X"10",X"10",X"00",X"00",X"00",X"40",X"C0",X"F0",
		X"0F",X"1F",X"1F",X"3F",X"31",X"01",X"01",X"00",X"01",X"01",X"09",X"0B",X"1F",X"1F",X"1F",X"1F",
		X"FF",X"FF",X"FF",X"F7",X"F6",X"F6",X"E6",X"6E",X"FC",X"EC",X"E8",X"D0",X"80",X"00",X"80",X"98",
		X"03",X"03",X"03",X"03",X"02",X"02",X"02",X"02",X"01",X"01",X"01",X"01",X"02",X"02",X"02",X"02",
		X"84",X"08",X"08",X"00",X"04",X"14",X"34",X"2C",X"28",X"28",X"38",X"38",X"30",X"30",X"70",X"70",
		X"01",X"01",X"03",X"03",X"03",X"03",X"03",X"00",X"00",X"00",X"00",X"06",X"1F",X"3F",X"7F",X"7F",
		X"F0",X"F8",X"FC",X"FC",X"F8",X"E0",X"E0",X"80",X"00",X"00",X"00",X"10",X"F8",X"FC",X"FC",X"FC",
		X"03",X"37",X"76",X"0C",X"0C",X"00",X"01",X"03",X"0F",X"1F",X"1F",X"1F",X"5F",X"CF",X"C7",X"C3",
		X"7E",X"3E",X"5E",X"DC",X"4D",X"71",X"FB",X"FA",X"36",X"02",X"00",X"00",X"80",X"80",X"8C",X"98",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"03",
		X"0E",X"1E",X"1E",X"3C",X"3C",X"38",X"78",X"70",X"72",X"E6",X"E4",X"C4",X"CC",X"C8",X"88",X"98",
		X"1F",X"1F",X"3F",X"3F",X"3F",X"3F",X"3E",X"1E",X"1C",X"00",X"C8",X"FE",X"FE",X"FE",X"FF",X"FB",
		X"00",X"80",X"C0",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"07",X"1F",X"02",X"00",X"00",X"00",X"00",X"00",X"06",X"0E",X"1E",
		X"01",X"03",X"07",X"0F",X"0F",X"9D",X"F8",X"F2",X"67",X"02",X"1F",X"FF",X"FB",X"F0",X"F0",X"70",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"03",X"07",X"07",X"0F",X"0F",
		X"06",X"1F",X"3F",X"3F",X"7F",X"7F",X"FB",X"F7",X"EE",X"CC",X"D0",X"B0",X"60",X"E0",X"C0",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"01",X"02",X"07",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"90",X"90",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"90",X"90",X"90",X"90",X"90",X"80",X"80",X"80",
		X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"20",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",
		X"98",X"98",X"98",X"98",X"90",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"40",X"40",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"03",X"03",X"06",X"06",
		X"98",X"90",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"40",X"40",X"40",X"20",X"20",X"30",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"03",X"07",X"07",X"0E",X"0E",X"1E",X"1E",X"1E",
		X"C0",X"C0",X"C0",X"C0",X"40",X"60",X"60",X"30",X"30",X"38",X"38",X"1C",X"1C",X"1E",X"1E",X"1E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"A0",X"60",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"20",X"00",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"3F",X"0F",X"07",X"0E",X"00",X"02",X"00",X"00",X"00",X"08",X"5E",X"4F",X"4F",X"67",X"30",
		X"7E",X"7F",X"7D",X"70",X"70",X"00",X"F0",X"30",X"38",X"18",X"18",X"38",X"38",X"38",X"30",X"40",
		X"3F",X"3F",X"1F",X"06",X"01",X"07",X"0F",X"0F",X"0E",X"06",X"06",X"06",X"03",X"03",X"01",X"01",
		X"C0",X"68",X"68",X"18",X"10",X"30",X"30",X"20",X"20",X"20",X"20",X"60",X"60",X"60",X"60",X"60",
		X"01",X"01",X"00",X"02",X"02",X"02",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"70",X"70",X"70",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"0F",X"0F",X"0F",X"0E",X"0E",X"0E",X"06",X"07",X"07",X"03",X"03",X"01",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FD",X"F8",X"F8",X"78",X"60",X"FC",X"7C",X"7C",X"BC",X"BE",X"1E",X"07",X"0F",
		X"31",X"39",X"19",X"19",X"00",X"7E",X"7F",X"7F",X"3B",X"00",X"00",X"00",X"01",X"01",X"01",X"00",
		X"F0",X"F0",X"F0",X"E4",X"C4",X"0C",X"0C",X"1C",X"C4",X"0C",X"06",X"86",X"E2",X"F2",X"F2",X"F2",
		X"01",X"05",X"05",X"06",X"02",X"03",X"03",X"03",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",
		X"E0",X"E0",X"E0",X"E0",X"70",X"70",X"70",X"70",X"F8",X"F8",X"F8",X"F8",X"FC",X"FC",X"FC",X"FC",
		X"3B",X"1B",X"19",X"1D",X"0D",X"0C",X"09",X"1D",X"05",X"05",X"02",X"00",X"00",X"01",X"01",X"01",
		X"FB",X"F1",X"E9",X"E8",X"F8",X"00",X"E0",X"F8",X"FE",X"FF",X"FF",X"3F",X"3F",X"3E",X"3E",X"9C",
		X"10",X"06",X"FF",X"FF",X"7F",X"3E",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"1F",X"2F",X"C7",X"01",X"00",X"40",X"F0",X"FC",X"FF",X"3F",X"0F",X"01",X"00",X"00",X"00",
		X"1F",X"0F",X"07",X"01",X"04",X"06",X"03",X"03",X"03",X"01",X"01",X"01",X"00",X"00",X"00",X"00",
		X"C0",X"C0",X"E0",X"E0",X"E0",X"F0",X"30",X"F0",X"F8",X"F8",X"F8",X"FC",X"FC",X"FC",X"FE",X"7E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DF",X"DF",X"5F",X"4E",X"69",X"3B",X"31",X"18",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1E",X"0C",X"04",X"20",X"2C",X"1F",X"3F",X"7E",X"7E",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7E",X"7F",X"7F",X"7F",X"DF",X"C3",X"C0",X"00",X"30",X"3E",X"7F",X"7F",X"1F",X"0F",X"00",X"00",
		X"0F",X"07",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"F8",X"FC",X"7C",X"96",X"E6",X"7F",X"7F",X"3F",X"3F",X"1F",X"1F",X"0F",X"0F",X"07",X"07",
		X"FF",X"FF",X"FF",X"FF",X"1F",X"1F",X"1E",X"06",X"1F",X"1E",X"9E",X"BD",X"F8",X"F0",X"F8",X"F9",
		X"F8",X"FC",X"FC",X"7E",X"66",X"66",X"66",X"E2",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"80",
		X"1F",X"0F",X"47",X"41",X"47",X"6F",X"4F",X"E0",X"E1",X"C2",X"C2",X"C0",X"81",X"85",X"8D",X"8B",
		X"98",X"38",X"30",X"80",X"FC",X"FC",X"F8",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"04",X"04",X"04",X"0C",X"0C",X"0C",X"0C",X"1F",X"1F",X"1F",X"1F",X"3F",X"3F",X"3F",X"3F",
		X"60",X"60",X"E0",X"E0",X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",
		X"DF",X"CF",X"97",X"37",X"13",X"1C",X"7E",X"FE",X"CD",X"C0",X"C0",X"C0",X"E0",X"E0",X"E3",X"E6",
		X"B8",X"B8",X"B0",X"30",X"60",X"60",X"E0",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"C3",X"DF",X"8F",X"87",X"0C",X"10",X"00",X"40",X"C0",X"80",X"80",X"80",X"00",X"00",X"00",
		X"18",X"C4",X"FC",X"F8",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"03",X"07",X"04",X"04",X"0C",X"0C",X"0F",X"1F",X"1F",X"1F",X"3F",X"3F",X"3F",X"7F",X"7E",
		X"30",X"30",X"70",X"60",X"E0",X"E0",X"C0",X"C0",X"C0",X"80",X"80",X"80",X"00",X"00",X"00",X"00",
		X"FB",X"FB",X"F2",X"66",X"8C",X"98",X"14",X"20",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3E",X"7E",X"78",X"F8",X"F3",X"F1",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"60",X"60",X"00",X"60",X"E0",X"F4",X"FC",X"3C",X"3E",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"1E",X"3C",X"39",X"63",X"67",X"FE",X"FE",X"FC",X"FC",X"F8",X"F8",X"F0",X"F0",X"E0",X"E0",
		X"00",X"40",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"C0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"05",X"0B",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"C0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"03",X"04",X"0E",X"0F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"30",X"70",X"F0",X"70",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"03",X"02",X"14",X"16",X"1C",X"07",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"30",X"B0",X"F0",X"70",X"F0",X"F0",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"03",X"02",X"14",X"1E",X"0C",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"10",X"58",X"78",X"F8",X"38",X"78",X"F8",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"03",X"02",X"24",X"2E",X"3E",X"0C",X"03",X"00",
		X"00",X"00",X"00",X"00",X"20",X"00",X"18",X"5C",X"7C",X"FC",X"1C",X"3C",X"7C",X"F8",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"02",X"02",X"03",X"03",X"02",X"0C",X"5C",X"7E",X"3C",X"00",X"07",X"00",
		X"00",X"20",X"10",X"10",X"08",X"2A",X"2E",X"7E",X"FE",X"1E",X"7E",X"FE",X"7C",X"F8",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"03",X"03",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"50",X"30",X"F0",X"70",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"03",X"01",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"58",X"B8",X"78",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"02",X"03",X"01",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"58",X"58",X"B4",X"7C",X"7C",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"0C",X"05",X"06",X"06",X"06",X"0C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"38",X"58",X"98",X"B4",X"7C",X"FC",X"FC",X"FC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"18",X"09",X"0D",X"0D",X"0D",X"0D",X"19",X"00",
		X"00",X"00",X"00",X"00",X"08",X"10",X"38",X"5C",X"DA",X"9E",X"3E",X"FE",X"FE",X"FE",X"FC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"30",X"11",X"1B",X"5D",X"1D",X"1D",X"3D",X"19",X"00",
		X"00",X"00",X"08",X"08",X"18",X"30",X"6C",X"DC",X"9A",X"1A",X"7E",X"FE",X"FE",X"FE",X"F8",X"00",
		X"00",X"00",X"04",X"02",X"00",X"60",X"30",X"3B",X"3B",X"BD",X"9D",X"1D",X"3D",X"79",X"0B",X"00",
		X"08",X"08",X"18",X"10",X"78",X"EC",X"CC",X"9A",X"9A",X"3E",X"FE",X"FE",X"FE",X"FC",X"F8",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"02",X"60",X"A1",X"33",X"7B",X"7B",X"7D",X"3D",X"3D",X"3D",X"79",X"F9",X"13",X"00",
		X"0E",X"1C",X"7E",X"77",X"E3",X"87",X"8F",X"8E",X"AC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"02",X"02",X"00",X"00",X"00",X"00",X"01",X"00",X"00",
		X"02",X"00",X"C0",X"60",X"71",X"73",X"FB",X"FD",X"7D",X"7D",X"7C",X"7C",X"F8",X"F9",X"13",X"00",
		X"1F",X"3B",X"33",X"F1",X"E3",X"C7",X"83",X"83",X"AF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"00",
		X"00",X"40",X"40",X"C0",X"C0",X"A0",X"20",X"A0",X"E0",X"E0",X"E0",X"E0",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"00",X"40",X"20",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"02",X"02",
		X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"40",X"40",X"00",X"20",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"06",X"06",X"02",X"00",
		X"00",X"80",X"A0",X"A0",X"A0",X"80",X"80",X"00",X"00",X"40",X"40",X"60",X"30",X"30",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"02",X"02",X"06",X"06",X"02",X"00",
		X"90",X"80",X"80",X"80",X"80",X"00",X"40",X"40",X"60",X"20",X"30",X"30",X"18",X"18",X"10",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"03",X"02",X"06",X"06",X"06",X"0E",X"0C",X"04",X"00",
		X"80",X"80",X"80",X"00",X"40",X"40",X"40",X"60",X"20",X"20",X"30",X"30",X"38",X"18",X"10",X"00",
		X"02",X"02",X"06",X"04",X"0C",X"0C",X"1C",X"1C",X"1C",X"38",X"38",X"18",X"00",X"00",X"00",X"00",
		X"80",X"80",X"C0",X"40",X"60",X"60",X"70",X"70",X"70",X"38",X"38",X"30",X"00",X"00",X"00",X"00",
		X"02",X"06",X"06",X"06",X"0E",X"0E",X"1C",X"1C",X"3C",X"38",X"18",X"00",X"00",X"00",X"00",X"00",
		X"20",X"30",X"30",X"30",X"38",X"38",X"1C",X"1C",X"1E",X"1E",X"1C",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"90",X"90",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"0E",X"0E",X"1E",X"1C",X"3C",X"3C",X"7C",X"78",X"38",X"00",X"00",X"00",X"00",X"00",X"00",
		X"18",X"18",X"18",X"1C",X"1C",X"1E",X"0E",X"0F",X"0F",X"0E",X"0C",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"90",X"98",X"98",X"98",X"98",X"98",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3E",X"3E",X"7C",X"7C",X"7C",X"FC",X"F8",X"F8",X"78",X"38",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"1F",X"0F",X"0F",X"0F",X"0F",X"07",X"07",X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"80",X"80",X"C0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"C0",X"C8",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"C0",X"C0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"40",X"F0",X"3A",X"3A",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"48",X"20",X"00",X"00",X"08",X"04",X"0E",X"36",X"5D",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"50",X"B8",X"08",X"50",X"08",X"00",X"00",X"10",X"08",X"04",X"0E",X"0A",X"04",X"2C",X"72",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"20",X"18",X"10",X"08",X"00",X"00",X"00",X"06",X"14",X"18",X"12",X"2C",X"4E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"10",X"00",X"18",X"08",X"00",X"28",X"1C",X"04",X"52",X"F6",X"5C",X"FA",X"B2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"20",X"02",X"28",X"00",X"14",X"28",X"38",X"AC",X"F6",X"D2",X"64",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"02",X"02",X"04",X"07",
		X"00",X"00",X"03",X"1F",X"3F",X"7F",X"FF",X"83",X"83",X"81",X"00",X"7F",X"FF",X"FF",X"FC",X"F8",
		X"00",X"00",X"C0",X"F8",X"FC",X"FE",X"FF",X"81",X"81",X"81",X"00",X"FC",X"FE",X"FE",X"3E",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"40",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",
		X"00",X"00",X"00",X"03",X"0F",X"1F",X"1F",X"31",X"21",X"41",X"40",X"9F",X"BF",X"3F",X"3C",X"FC",
		X"00",X"00",X"7C",X"FF",X"FF",X"FF",X"FF",X"C0",X"C0",X"C0",X"00",X"FE",X"FF",X"FF",X"3F",X"1F",
		X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"60",X"60",X"20",X"20",X"40",X"40",X"40",X"40",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",
		X"00",X"00",X"00",X"00",X"03",X"07",X"0F",X"19",X"11",X"21",X"40",X"5F",X"BF",X"3F",X"38",X"F8",
		X"00",X"00",X"1F",X"FF",X"FF",X"FF",X"FF",X"C0",X"C0",X"C0",X"00",X"FE",X"FF",X"FF",X"7F",X"3F",
		X"00",X"00",X"80",X"C0",X"C0",X"E0",X"E0",X"60",X"60",X"20",X"20",X"40",X"40",X"40",X"40",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"07",
		X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"0D",X"09",X"11",X"20",X"5F",X"BF",X"3F",X"30",X"E0",
		X"00",X"00",X"07",X"3F",X"FF",X"FF",X"FF",X"C0",X"C0",X"C0",X"00",X"FE",X"FF",X"FF",X"FF",X"7F",
		X"00",X"00",X"E0",X"F0",X"F8",X"F8",X"F8",X"38",X"30",X"10",X"30",X"30",X"60",X"60",X"C0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"0C",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"0F",X"0B",X"33",X"40",X"BF",X"7F",X"7F",X"61",X"81",
		X"00",X"00",X"03",X"1F",X"FF",X"FF",X"FF",X"80",X"80",X"80",X"00",X"FC",X"FE",X"FE",X"FF",X"FF",
		X"00",X"00",X"F0",X"F8",X"FC",X"FC",X"FC",X"38",X"38",X"38",X"70",X"60",X"60",X"C0",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"06",X"08",X"30",X"7F",
		X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"1F",X"17",X"27",X"C0",X"7F",X"FF",X"FF",X"87",X"07",
		X"00",X"00",X"00",X"0F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"F8",X"FC",X"FD",X"FF",X"FE",
		X"00",X"00",X"F8",X"FE",X"FE",X"FE",X"FC",X"3C",X"3C",X"38",X"30",X"60",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"0C",X"10",X"7E",
		X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"0F",X"0F",X"37",X"40",X"FF",X"FF",X"FF",X"0F",X"07",
		X"00",X"00",X"00",X"07",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"F8",X"FD",X"FF",X"FE",X"F8",
		X"00",X"00",X"3F",X"FF",X"FF",X"FF",X"FF",X"1E",X"1C",X"38",X"60",X"C0",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"0F",X"11",X"E0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"0E",X"0E",X"1E",X"E0",X"FF",X"FF",X"FF",X"0F",X"07",
		X"00",X"00",X"00",X"01",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"F0",X"F9",X"FF",X"FE",X"F8",
		X"00",X"00",X"1F",X"FF",X"FF",X"FF",X"FF",X"0F",X"0F",X"1E",X"38",X"E0",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"80",X"E0",X"E0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"3B",X"C0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"01",X"0F",X"1F",X"1C",X"1C",X"60",X"FF",X"FF",X"FF",X"7F",X"3F",
		X"00",X"00",X"00",X"00",X"7F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"E0",X"F1",X"F7",X"FE",X"F8",
		X"00",X"00",X"07",X"7F",X"FF",X"FF",X"FF",X"0F",X"0F",X"0E",X"3C",X"F0",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"F0",X"F8",X"F8",X"F8",X"F0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"06",X"0E",X"0E",X"1F",X"1F",X"3F",X"7F",X"35",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E3",X"FE",
		X"14",X"0C",X"2C",X"38",X"30",X"18",X"78",X"58",X"18",X"18",X"1C",X"1C",X"1C",X"0C",X"EE",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"03",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"C0",X"00",
		X"00",X"04",X"28",X"3C",X"38",X"30",X"30",X"20",X"60",X"60",X"60",X"60",X"E0",X"C0",X"C0",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"7F",X"7B",X"77",X"BF",X"DF",X"77",X"AF",X"0C",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"FE",X"FE",X"EE",X"F5",X"FB",X"FE",X"F4",X"60",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"7F",X"7B",X"77",X"2F",X"DF",X"B7",X"5F",X"0C",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"FE",X"FE",X"EE",X"F5",X"FA",X"FC",X"FA",X"60",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"1F",X"3F",X"3F",X"37",X"27",X"23",X"60",X"70",X"20",X"00",X"10",
		X"00",X"00",X"00",X"00",X"E0",X"F8",X"FC",X"FC",X"F6",X"F2",X"F2",X"62",X"0E",X"0C",X"1C",X"78",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"0F",X"0F",X"07",X"06",X"02",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"F0",X"F0",X"F0",X"70",X"70",X"70",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"40",X"60",X"30",X"1F",X"0F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"08",X"00",X"18",X"F8",X"F0",X"20",X"20",
		X"00",X"00",X"00",X"00",X"03",X"07",X"0F",X"0F",X"07",X"0E",X"0B",X"00",X"00",X"00",X"00",X"18",
		X"00",X"00",X"00",X"00",X"E0",X"E0",X"F0",X"F0",X"F0",X"70",X"70",X"60",X"00",X"00",X"40",X"F8",
		X"60",X"3F",X"3F",X"1F",X"0F",X"00",X"01",X"03",X"02",X"06",X"06",X"02",X"02",X"07",X"07",X"03",
		X"60",X"F4",X"F4",X"78",X"08",X"00",X"20",X"60",X"60",X"60",X"E0",X"E0",X"60",X"60",X"60",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"06",X"00",X"08",X"08",
		X"0F",X"07",X"07",X"03",X"00",X"00",X"00",X"38",X"FD",X"FF",X"FF",X"1E",X"1D",X"0D",X"0D",X"2B",
		X"F0",X"F0",X"F0",X"F0",X"B0",X"00",X"00",X"40",X"C0",X"F0",X"F8",X"F8",X"FC",X"FC",X"DC",X"9C",
		X"00",X"00",X"03",X"07",X"07",X"03",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"00",X"00",
		X"00",X"40",X"00",X"00",X"20",X"A0",X"A0",X"A0",X"E0",X"E0",X"E0",X"E0",X"E0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"03",X"07",X"06",X"04",X"00",X"00",X"00",X"80",X"C0",X"60",X"30",X"18",
		X"3C",X"7C",X"EF",X"DD",X"9D",X"1B",X"38",X"33",X"37",X"3F",X"2E",X"24",X"03",X"41",X"41",X"80",
		X"18",X"10",X"20",X"F0",X"F8",X"78",X"F0",X"E0",X"C0",X"80",X"00",X"C0",X"A0",X"80",X"C0",X"C0",
		X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"01",X"01",X"01",X"03",X"03",X"03",X"03",X"03",X"01",
		X"1C",X"8C",X"8C",X"8C",X"88",X"88",X"98",X"18",X"10",X"30",X"30",X"30",X"E0",X"E0",X"E0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"0F",X"3C",
		X"07",X"07",X"07",X"03",X"00",X"01",X"01",X"00",X"03",X"03",X"01",X"30",X"F8",X"FF",X"FB",X"C7",
		X"80",X"C0",X"80",X"80",X"00",X"20",X"60",X"40",X"20",X"60",X"D0",X"30",X"F0",X"E0",X"C0",X"C0",
		X"06",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"0F",X"1F",
		X"FC",X"FE",X"7E",X"06",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"1F",X"3F",X"1F",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"0F",X"7F",X"FF",X"FE",X"FE",X"FC",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"07",X"0D",X"01",X"03",X"26",X"7F",X"CF",X"9F",X"3D",X"2C",X"07",X"21",X"18",X"03",X"00",
		X"00",X"00",X"00",X"B0",X"78",X"FC",X"DC",X"CE",X"E6",X"A2",X"01",X"00",X"C0",X"60",X"E0",X"70",
		X"27",X"33",X"33",X"33",X"17",X"1F",X"19",X"1C",X"0C",X"0C",X"0C",X"0E",X"06",X"06",X"07",X"07",
		X"90",X"A0",X"80",X"00",X"80",X"80",X"80",X"80",X"C0",X"C0",X"C0",X"40",X"60",X"60",X"E0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"04",X"06",X"03",X"01",X"02",X"01",X"00",X"00",X"04",X"0F",X"1B",X"13",X"17",X"25",
		X"78",X"08",X"88",X"D0",X"E0",X"E0",X"E0",X"A0",X"2E",X"5F",X"B7",X"F3",X"F8",X"EC",X"84",X"A0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"70",X"18",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"03",X"03",X"07",X"07",X"07",X"07",X"03",X"01",X"01",X"01",X"01",X"01",X"02",X"02",X"02",
		X"C1",X"C3",X"82",X"82",X"84",X"84",X"00",X"80",X"80",X"80",X"E0",X"E0",X"E0",X"F0",X"F0",X"F0",
		X"00",X"00",X"07",X"FF",X"FF",X"FE",X"38",X"70",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"1D",X"1F",X"1F",X"00",X"07",X"3F",X"FF",X"FF",X"7F",
		X"00",X"00",X"00",X"00",X"03",X"1F",X"FF",X"FC",X"E0",X"00",X"E3",X"FF",X"FC",X"F0",X"C0",X"00",
		X"04",X"06",X"06",X"07",X"07",X"07",X"03",X"07",X"03",X"03",X"53",X"0F",X"1F",X"0F",X"07",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"A0",X"C0",X"C8",X"D2",X"F8",X"F0",X"E8",X"F0",X"D8",
		X"04",X"06",X"06",X"07",X"07",X"07",X"03",X"03",X"13",X"07",X"0F",X"07",X"0F",X"9F",X"0F",X"07",
		X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"C8",X"D0",X"F8",X"D0",X"F0",X"F9",X"EC",X"B0",
		X"0C",X"0E",X"07",X"07",X"07",X"03",X"03",X"03",X"03",X"03",X"03",X"07",X"07",X"07",X"07",X"0F",
		X"00",X"00",X"00",X"80",X"C0",X"C0",X"E0",X"E0",X"F8",X"F2",X"F4",X"FC",X"FE",X"FD",X"F8",X"FC",
		X"0C",X"0E",X"07",X"07",X"07",X"03",X"03",X"03",X"03",X"03",X"03",X"07",X"07",X"07",X"07",X"07",
		X"00",X"00",X"00",X"80",X"C0",X"C0",X"E0",X"E0",X"F4",X"F0",X"FA",X"FC",X"FE",X"FC",X"F8",X"F4",
		X"03",X"03",X"03",X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"F8",X"F8",X"F8",X"FC",X"FC",X"FE",X"1E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"1F",X"1F",X"1F",X"3F",X"3F",X"7F",X"78",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"03",X"03",X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"F8",X"F8",X"F8",X"F8",X"FC",X"FE",X"1E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"3F",X"1F",X"1F",X"3F",X"3F",X"7F",X"78",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"07",X"07",X"07",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F8",X"FC",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"7F",X"3F",X"3F",X"7F",X"7F",X"FE",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"07",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"C1",X"C0",X"C0",X"C0",X"F0",X"F9",X"79",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"7F",X"7F",X"7E",X"FE",X"FC",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"3F",X"3F",X"3F",X"1F",X"1F",X"0F",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"07",X"01",X"01",X"01",X"C3",X"E7",X"E7",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FE",X"FC",X"FC",X"F8",X"F8",X"F0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FC",X"FC",X"FC",X"7C",X"7F",X"3F",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"1F",X"07",X"07",X"07",X"0F",X"9F",X"9E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"F8",X"F0",X"F0",X"E0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"F8",X"F8",X"F8",X"F8",X"FE",X"7F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"1F",X"0F",X"0F",X"0F",X"1F",X"3F",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"E0",X"E0",X"E0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"07",X"07",X"07",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"C0",X"C0",X"C0",X"C0",X"F8",X"FC",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"7F",X"1F",X"1F",X"1F",X"3F",X"FE",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"0F",X"0F",X"0F",X"07",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"81",X"80",X"80",X"C0",X"F0",X"F9",X"79",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"7F",X"7F",X"7E",X"FE",X"FC",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"04",X"0A",X"06",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"3F",X"FF",X"1F",X"3F",X"7F",X"C1",X"6C",X"2C",X"7E",X"3F",X"1F",X"3F",X"1F",X"08",
		X"86",X"8C",X"CC",X"C4",X"CC",X"8C",X"9C",X"1E",X"3F",X"F6",X"F4",X"0E",X"FD",X"D0",X"00",X"80",
		X"07",X"07",X"1F",X"0F",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"C0",X"E0",X"F0",X"80",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7C",X"F8",X"73",X"97",X"6F",X"0F",X"07",X"1F",X"3B",X"10",X"0B",X"1F",X"0F",X"07",X"0F",X"06",
		X"00",X"00",X"E0",X"E0",X"F1",X"F1",X"F1",X"E1",X"EB",X"0B",X"1C",X"37",X"E3",X"F0",X"80",X"40",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"80",X"C0",X"60",X"C0",X"A0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"07",X"1F",X"0F",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"F0",X"E0",X"80",
		X"03",X"23",X"63",X"F7",X"F7",X"F7",X"57",X"63",X"B3",X"3F",X"17",X"03",X"04",X"00",X"00",X"00",
		X"80",X"9C",X"FE",X"FF",X"FF",X"FF",X"FA",X"B5",X"CE",X"F8",X"B0",X"C0",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"07",X"0F",X"07",X"09",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"E0",X"F0",X"60",
		X"03",X"23",X"63",X"73",X"F7",X"F7",X"D7",X"67",X"33",X"2F",X"1B",X"07",X"03",X"00",X"00",X"00",
		X"80",X"9C",X"FE",X"FE",X"FF",X"FF",X"B8",X"B6",X"CE",X"FC",X"E8",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"03",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"04",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"00",X"00",X"00",X"00",
		X"1F",X"1F",X"1F",X"0F",X"07",X"0E",X"00",X"00",X"40",X"40",X"40",X"40",X"40",X"40",X"20",X"1F",
		X"F8",X"F8",X"78",X"78",X"70",X"08",X"08",X"0C",X"0C",X"1C",X"0C",X"08",X"00",X"00",X"00",X"E0",
		X"0F",X"07",X"37",X"72",X"30",X"28",X"70",X"30",X"38",X"1F",X"1F",X"0F",X"07",X"03",X"0B",X"04",
		X"F0",X"F0",X"FC",X"7E",X"72",X"06",X"0E",X"5E",X"FE",X"FC",X"F8",X"78",X"70",X"60",X"08",X"08",
		X"00",X"40",X"40",X"40",X"40",X"60",X"20",X"20",X"13",X"0F",X"0C",X"0C",X"0C",X"0E",X"0E",X"0F",
		X"0C",X"0C",X"1C",X"0C",X"00",X"00",X"00",X"00",X"E0",X"60",X"60",X"60",X"60",X"60",X"60",X"E0",
		X"00",X"00",X"00",X"18",X"7F",X"FF",X"3F",X"0F",X"0F",X"0F",X"00",X"02",X"02",X"00",X"00",X"40",
		X"00",X"00",X"40",X"F8",X"FE",X"FF",X"7C",X"70",X"70",X"70",X"00",X"60",X"48",X"08",X"18",X"18",
		X"00",X"00",X"04",X"04",X"04",X"04",X"04",X"04",X"06",X"06",X"07",X"07",X"07",X"07",X"07",X"07",
		X"20",X"60",X"E0",X"C0",X"E0",X"E0",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"E0",X"E0",X"E0",
		X"3F",X"7F",X"7F",X"7F",X"3F",X"0F",X"0F",X"00",X"07",X"02",X"02",X"00",X"00",X"41",X"47",X"43",
		X"FC",X"FE",X"FE",X"7F",X"7B",X"71",X"70",X"00",X"30",X"38",X"08",X"18",X"78",X"78",X"30",X"00",
		X"01",X"01",X"01",X"01",X"01",X"05",X"04",X"06",X"06",X"06",X"06",X"07",X"07",X"07",X"07",X"07",
		X"60",X"60",X"60",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"60",X"38",X"0C",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"13",X"0F",X"03",X"00",X"00",X"00",X"10",X"30",X"38",X"B8",X"98",X"C0",X"FF",X"FF",X"7F",X"1D",
		X"98",X"18",X"D8",X"18",X"30",X"30",X"30",X"30",X"10",X"58",X"D8",X"C8",X"08",X"08",X"08",X"C8",
		X"00",X"02",X"02",X"02",X"02",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"70",X"70",X"70",X"70",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"F8",X"FC",X"FC",X"7C",X"7C",X"7C",X"3C",X"18",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"06",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"01",X"03",X"03",X"07",X"07",X"E6",X"F8",X"F8",X"7C",X"2F",X"06",X"00",X"00",X"00",X"00",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"80",X"10",X"30",X"78",X"78",X"F8",X"38",X"7C",X"3E",X"3E",X"1E",
		X"09",X"09",X"09",X"09",X"19",X"19",X"1F",X"1F",X"3F",X"3F",X"3E",X"3E",X"3C",X"18",X"00",X"00",
		X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"70",X"40",X"00",X"00",X"00",X"00",X"02",X"06",X"64",X"01",X"80",X"92",X"07",X"06",X"06",X"06",
		X"0E",X"18",X"58",X"38",X"0D",X"07",X"0F",X"3D",X"FE",X"82",X"20",X"7C",X"FF",X"FF",X"7F",X"7F",
		X"80",X"00",X"20",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"E0",X"F0",X"F8",
		X"00",X"07",X"3F",X"7F",X"FF",X"FF",X"7E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"1F",X"3F",X"FF",X"F8",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FC",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"1F",X"0F",X"03",X"00",X"24",X"36",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"40",X"40",X"80",X"00",
		X"01",X"01",X"03",X"13",X"13",X"51",X"78",X"70",X"43",X"07",X"0F",X"0F",X"07",X"07",X"07",X"07",
		X"E0",X"E8",X"B0",X"F0",X"F4",X"C4",X"00",X"04",X"0C",X"2C",X"CC",X"88",X"08",X"18",X"90",X"90",
		X"03",X"03",X"03",X"03",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",X"FC",X"FC",X"FC",X"7C",X"7C",X"38",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"F0",X"F8",
		X"04",X"04",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"03",X"00",X"01",X"01",X"03",X"03",
		X"7C",X"8E",X"3E",X"1E",X"23",X"7F",X"EF",X"FD",X"FD",X"3C",X"80",X"C0",X"C0",X"E0",X"F1",X"E1",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"00",X"80",X"80",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"70",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"07",X"07",X"07",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"80",X"80",X"C0",X"E0",X"FC",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"7E",X"7E",X"FC",X"F0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"07",X"07",X"0F",X"0F",X"1E",X"37",X"1E",X"68",X"40",X"08",X"40",X"00",X"00",X"20",X"00",
		X"C0",X"E2",X"B0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"0F",X"0F",X"07",X"0D",X"1F",X"0C",X"18",X"14",X"20",X"00",X"00",X"10",X"80",X"00",X"00",
		X"E8",X"80",X"E0",X"A0",X"D2",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"3F",X"1F",X"3E",X"1E",X"77",X"18",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FA",X"F0",X"C0",X"E4",X"40",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"1F",X"3F",X"1F",X"6C",X"D8",X"12",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"F0",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
