module SN74LS393(
	input			A2,			//01
	input			CLR2,			//02	
	output		Q2A,			//03
	output		Q2B,			//04
	output		Q2C,			//05
	output		Q2D,			//06
	
	output		Q1D,			//03
	output		Q1C,			//09
	output		Q1B,			//10
	output		Q1A,			//11
	input			CLR1,			//12
	input			A1				//01
);

wire	SYNTHESIZED_WIRE_28;
wire	SYNTHESIZED_WIRE_29;
wire	SYNTHESIZED_WIRE_2;
wire	SYNTHESIZED_WIRE_3;
reg	DFF_9;
reg	SYNTHESIZED_WIRE_30;
reg	SYNTHESIZED_WIRE_31;
reg	SYNTHESIZED_WIRE_32;
reg	SYNTHESIZED_WIRE_33;
reg	SYNTHESIZED_WIRE_34;
wire	SYNTHESIZED_WIRE_35;
wire	SYNTHESIZED_WIRE_36;
wire	SYNTHESIZED_WIRE_6;
wire	SYNTHESIZED_WIRE_9;
wire	SYNTHESIZED_WIRE_12;
wire	SYNTHESIZED_WIRE_15;
wire	SYNTHESIZED_WIRE_18;
wire	SYNTHESIZED_WIRE_19;
reg	SYNTHESIZED_WIRE_37;
wire	SYNTHESIZED_WIRE_20;
reg	DFF_31;
wire	SYNTHESIZED_WIRE_23;
wire	SYNTHESIZED_WIRE_24;
wire	SYNTHESIZED_WIRE_27;

assign	Q2A = SYNTHESIZED_WIRE_33;
assign	Q2B = SYNTHESIZED_WIRE_34;
assign	Q2C = SYNTHESIZED_WIRE_37;
assign	Q2D = DFF_31;
assign	Q1D = DFF_9;
assign	Q1C = SYNTHESIZED_WIRE_32;
assign	Q1B = SYNTHESIZED_WIRE_30;
assign	Q1A = SYNTHESIZED_WIRE_31;




always@(posedge SYNTHESIZED_WIRE_29 or negedge SYNTHESIZED_WIRE_28)
begin
if (!SYNTHESIZED_WIRE_28)
	begin
	SYNTHESIZED_WIRE_31 <= 0;
	end
else
	begin
	SYNTHESIZED_WIRE_31 <= SYNTHESIZED_WIRE_2;
	end
end

assign	SYNTHESIZED_WIRE_27 = SYNTHESIZED_WIRE_3 ^ DFF_9;

assign	SYNTHESIZED_WIRE_3 = SYNTHESIZED_WIRE_30 & SYNTHESIZED_WIRE_31 & SYNTHESIZED_WIRE_32;

assign	SYNTHESIZED_WIRE_29 =  ~A1;

assign	SYNTHESIZED_WIRE_28 =  ~CLR1;

assign	SYNTHESIZED_WIRE_2 =  ~SYNTHESIZED_WIRE_31;

assign	SYNTHESIZED_WIRE_35 =  ~CLR2;

assign	SYNTHESIZED_WIRE_36 =  ~A2;

assign	SYNTHESIZED_WIRE_6 =  ~SYNTHESIZED_WIRE_33;

assign	SYNTHESIZED_WIRE_19 = SYNTHESIZED_WIRE_34 & SYNTHESIZED_WIRE_33;


always@(posedge SYNTHESIZED_WIRE_36 or negedge SYNTHESIZED_WIRE_35)
begin
if (!SYNTHESIZED_WIRE_35)
	begin
	SYNTHESIZED_WIRE_33 <= 0;
	end
else
	begin
	SYNTHESIZED_WIRE_33 <= SYNTHESIZED_WIRE_6;
	end
end


always@(posedge SYNTHESIZED_WIRE_36 or negedge SYNTHESIZED_WIRE_35)
begin
if (!SYNTHESIZED_WIRE_35)
	begin
	SYNTHESIZED_WIRE_34 <= 0;
	end
else
	begin
	SYNTHESIZED_WIRE_34 <= SYNTHESIZED_WIRE_9;
	end
end


always@(posedge SYNTHESIZED_WIRE_29 or negedge SYNTHESIZED_WIRE_28)
begin
if (!SYNTHESIZED_WIRE_28)
	begin
	SYNTHESIZED_WIRE_30 <= 0;
	end
else
	begin
	SYNTHESIZED_WIRE_30 <= SYNTHESIZED_WIRE_12;
	end
end


always@(posedge SYNTHESIZED_WIRE_36 or negedge SYNTHESIZED_WIRE_35)
begin
if (!SYNTHESIZED_WIRE_35)
	begin
	SYNTHESIZED_WIRE_37 <= 0;
	end
else
	begin
	SYNTHESIZED_WIRE_37 <= SYNTHESIZED_WIRE_15;
	end
end


always@(posedge SYNTHESIZED_WIRE_36 or negedge SYNTHESIZED_WIRE_35)
begin
if (!SYNTHESIZED_WIRE_35)
	begin
	DFF_31 <= 0;
	end
else
	begin
	DFF_31 <= SYNTHESIZED_WIRE_18;
	end
end

assign	SYNTHESIZED_WIRE_9 = SYNTHESIZED_WIRE_33 ^ SYNTHESIZED_WIRE_34;

assign	SYNTHESIZED_WIRE_15 = SYNTHESIZED_WIRE_19 ^ SYNTHESIZED_WIRE_37;

assign	SYNTHESIZED_WIRE_18 = SYNTHESIZED_WIRE_20 ^ DFF_31;

assign	SYNTHESIZED_WIRE_20 = SYNTHESIZED_WIRE_34 & SYNTHESIZED_WIRE_33 & SYNTHESIZED_WIRE_37;

assign	SYNTHESIZED_WIRE_12 = SYNTHESIZED_WIRE_31 ^ SYNTHESIZED_WIRE_30;


always@(posedge SYNTHESIZED_WIRE_29 or negedge SYNTHESIZED_WIRE_28)
begin
if (!SYNTHESIZED_WIRE_28)
	begin
	SYNTHESIZED_WIRE_32 <= 0;
	end
else
	begin
	SYNTHESIZED_WIRE_32 <= SYNTHESIZED_WIRE_23;
	end
end

assign	SYNTHESIZED_WIRE_23 = SYNTHESIZED_WIRE_24 ^ SYNTHESIZED_WIRE_32;

assign	SYNTHESIZED_WIRE_24 = SYNTHESIZED_WIRE_30 & SYNTHESIZED_WIRE_31;


always@(posedge SYNTHESIZED_WIRE_29 or negedge SYNTHESIZED_WIRE_28)
begin
if (!SYNTHESIZED_WIRE_28)
	begin
	DFF_9 <= 0;
	end
else
	begin
	DFF_9 <= SYNTHESIZED_WIRE_27;
	end
end


endmodule
