`define BUILD_DATE "190322"
`define BUILD_TIME "101029"
