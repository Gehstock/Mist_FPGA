library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity rom1t36 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of rom1t36 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"C2",X"27",X"19",X"2A",X"A7",X"7D",X"2A",X"C2",X"41",X"CD",X"C3",X"40",X"01",X"81",X"FE",X"7C",
		X"13",X"20",X"44",X"23",X"E1",X"4D",X"00",X"C9",X"C3",X"19",X"1B",X"C6",X"01",X"3E",X"D6",X"32",
		X"23",X"13",X"C2",X"0D",X"02",X"22",X"F3",X"C9",X"00",X"00",X"47",X"7E",X"77",X"1A",X"12",X"78",
		X"20",X"F5",X"CA",X"A7",X"17",X"E4",X"A6",X"C3",X"CA",X"76",X"03",X"3D",X"93",X"C3",X"3A",X"02",
		X"ED",X"C2",X"CD",X"1E",X"1F",X"92",X"1E",X"C3",X"C2",X"40",X"1F",X"54",X"92",X"CD",X"C9",X"1F",
		X"20",X"E6",X"32",X"3C",X"20",X"E6",X"51",X"C3",X"CD",X"1F",X"15",X"D2",X"D2",X"C3",X"3A",X"1D",
		X"51",X"C3",X"3A",X"02",X"20",X"E4",X"32",X"3C",X"3A",X"02",X"20",X"E5",X"32",X"3C",X"20",X"E5",
		X"32",X"3C",X"20",X"E3",X"51",X"C3",X"21",X"02",X"20",X"E4",X"51",X"C3",X"3A",X"02",X"20",X"E3",
		X"E4",X"32",X"21",X"20",X"21",X"C0",X"00",X"C9",X"21",X"00",X"32",X"97",X"20",X"E3",X"97",X"C9",
		X"E5",X"20",X"CD",X"D5",X"15",X"B4",X"E1",X"D1",X"00",X"00",X"11",X"00",X"20",X"B0",X"D3",X"2A",
		X"15",X"96",X"DE",X"C3",X"3A",X"15",X"20",X"E1",X"D6",X"3A",X"A7",X"20",X"D9",X"C2",X"CD",X"03",
		X"20",X"E0",X"CA",X"A7",X"04",X"EE",X"CC",X"C3",X"CA",X"A7",X"04",X"EE",X"A1",X"C3",X"3A",X"01",
		X"11",X"06",X"14",X"00",X"06",X"CD",X"11",X"15",X"3A",X"01",X"20",X"F6",X"0A",X"FE",X"D6",X"DA",
		X"B4",X"CD",X"3A",X"15",X"20",X"D6",X"01",X"FE",X"20",X"B0",X"F0",X"21",X"22",X"32",X"20",X"D3",
		X"15",X"96",X"32",X"97",X"20",X"D1",X"DA",X"32",X"1C",X"CA",X"C3",X"03",X"03",X"78",X"CD",X"00",
		X"20",X"E8",X"02",X"3E",X"32",X"00",X"20",X"F5",X"32",X"20",X"20",X"D7",X"D9",X"32",X"32",X"20",
		X"20",X"D2",X"02",X"3E",X"DD",X"32",X"32",X"20",X"05",X"3E",X"00",X"32",X"3E",X"20",X"32",X"10",
		X"32",X"01",X"20",X"D8",X"32",X"97",X"20",X"D6",X"20",X"CF",X"10",X"3E",X"D5",X"32",X"3E",X"20",
		X"97",X"13",X"F6",X"32",X"C3",X"20",X"08",X"EE",X"D0",X"32",X"00",X"20",X"00",X"00",X"66",X"C3",
		X"03",X"1C",X"9E",X"C3",X"D5",X"03",X"C3",X"C5",X"12",X"FE",X"94",X"C2",X"78",X"03",X"C2",X"A7",
		X"4E",X"CA",X"3E",X"03",X"47",X"20",X"E8",X"3A",X"02",X"C1",X"00",X"06",X"03",X"DB",X"08",X"E6",
		X"3E",X"20",X"C3",X"22",X"03",X"60",X"20",X"3E",X"A7",X"20",X"5E",X"CA",X"3D",X"03",X"E8",X"32",
		X"00",X"20",X"02",X"3E",X"E8",X"32",X"21",X"20",X"D3",X"B0",X"C3",X"01",X"05",X"89",X"DA",X"32",
		X"60",X"01",X"C3",X"00",X"03",X"8E",X"48",X"CD",X"20",X"EA",X"C3",X"34",X"16",X"41",X"00",X"00",
		X"D3",X"20",X"C3",X"01",X"00",X"C3",X"8D",X"21",X"C3",X"0B",X"00",X"F7",X"33",X"CA",X"3E",X"13",
		X"E6",X"7D",X"C3",X"1F",X"03",X"30",X"09",X"EB",X"5D",X"31",X"46",X"54",X"7E",X"23",X"47",X"B0",
		X"11",X"32",X"20",X"B0",X"E7",X"C3",X"21",X"02",X"FE",X"7C",X"C2",X"34",X"03",X"91",X"F0",X"21",
		X"0C",X"11",X"21",X"01",X"22",X"C0",X"0C",X"06",X"00",X"00",X"EB",X"22",X"22",X"20",X"20",X"DB",
		X"00",X"21",X"36",X"24",X"23",X"00",X"FE",X"7C",X"97",X"EF",X"CE",X"32",X"C9",X"22",X"04",X"D3",
		X"3E",X"00",X"D3",X"24",X"3A",X"01",X"20",X"AF",X"C2",X"40",X"03",X"CB",X"00",X"C9",X"00",X"00",
		X"C3",X"20",X"13",X"AE",X"32",X"97",X"20",X"AF",X"FF",X"FE",X"96",X"CA",X"3C",X"13",X"AF",X"32",
		X"E6",X"7B",X"5F",X"E0",X"C3",X"19",X"17",X"B3",X"00",X"3E",X"01",X"D3",X"50",X"C3",X"57",X"4A",
		X"C5",X"F3",X"E5",X"D5",X"C3",X"F5",X"02",X"37",X"31",X"F3",X"20",X"A0",X"C3",X"97",X"48",X"00",
		X"06",X"C5",X"0E",X"A0",X"0D",X"A0",X"1D",X"C2",X"1F",X"C3",X"C2",X"40",X"00",X"28",X"00",X"C9",
		X"77",X"1A",X"23",X"13",X"C3",X"05",X"00",X"13",X"05",X"00",X"04",X"D3",X"C5",X"C3",X"00",X"47",
		X"06",X"20",X"21",X"0C",X"20",X"A4",X"00",X"11",X"A1",X"32",X"32",X"20",X"20",X"A2",X"A3",X"32",
		X"CD",X"FB",X"09",X"43",X"00",X"00",X"D0",X"C3",X"EF",X"01",X"50",X"C3",X"CD",X"01",X"09",X"CB",
		X"21",X"40",X"08",X"06",X"21",X"EF",X"21",X"80",X"11",X"06",X"01",X"18",X"08",X"06",X"21",X"EF",
		X"06",X"EF",X"21",X"05",X"20",X"F6",X"21",X"EF",X"08",X"06",X"21",X"EF",X"21",X"C0",X"08",X"06",
		X"22",X"00",X"01",X"21",X"36",X"20",X"23",X"00",X"00",X"00",X"ED",X"22",X"3E",X"20",X"32",X"05",
		X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"7D",X"DA",X"24",X"00",X"7D",X"C6",X"CD",
		X"04",X"D3",X"AE",X"CD",X"3A",X"1E",X"20",X"F5",X"00",X"00",X"27",X"21",X"22",X"00",X"20",X"03",
		X"C2",X"02",X"00",X"98",X"39",X"C3",X"32",X"00",X"C2",X"A7",X"03",X"42",X"EF",X"3A",X"FE",X"20",
		X"C3",X"20",X"00",X"30",X"F5",X"3A",X"A7",X"20",X"20",X"E8",X"B9",X"C3",X"00",X"06",X"F5",X"32",
		X"A7",X"20",X"D3",X"C2",X"2A",X"00",X"20",X"A5",X"84",X"C3",X"C5",X"03",X"E5",X"D5",X"E2",X"3A",
		X"00",X"20",X"11",X"FE",X"EA",X"D2",X"01",X"00",X"D6",X"C3",X"2A",X"00",X"20",X"A9",X"01",X"78",
		X"01",X"00",X"2A",X"CD",X"A7",X"13",X"4A",X"C2",X"00",X"50",X"0E",X"FE",X"EA",X"D2",X"01",X"00",
		X"C1",X"D1",X"28",X"3E",X"31",X"C3",X"00",X"13",X"22",X"01",X"20",X"A5",X"40",X"CD",X"E1",X"0B",
		X"00",X"38",X"00",X"00",X"30",X"5D",X"18",X"00",X"00",X"2F",X"00",X"00",X"00",X"25",X"00",X"00",
		X"3E",X"82",X"13",X"00",X"2F",X"87",X"13",X"00",X"27",X"41",X"1A",X"00",X"35",X"01",X"1A",X"00",
		X"3E",X"FC",X"12",X"00",X"2F",X"95",X"12",X"00",X"28",X"FC",X"12",X"00",X"36",X"92",X"12",X"00",
		X"08",X"00",X"88",X"48",X"00",X"C8",X"01",X"00",X"28",X"F9",X"11",X"00",X"2F",X"92",X"11",X"00",
		X"C9",X"C1",X"A9",X"22",X"C3",X"20",X"03",X"7E",X"00",X"FE",X"FF",X"00",X"C2",X"FF",X"00",X"1B",
		X"C3",X"EF",X"00",X"45",X"75",X"21",X"C3",X"00",X"ED",X"21",X"11",X"20",X"01",X"3D",X"08",X"06",
		X"FE",X"20",X"C2",X"01",X"01",X"FF",X"E0",X"3A",X"09",X"03",X"00",X"00",X"00",X"00",X"F1",X"3A",
		X"3E",X"20",X"32",X"01",X"20",X"F5",X"C9",X"E1",X"A7",X"20",X"0C",X"CA",X"3D",X"06",X"E0",X"32",
		X"E0",X"3A",X"A7",X"20",X"95",X"C2",X"CD",X"01",X"3A",X"00",X"20",X"E2",X"C2",X"A7",X"01",X"B2",
		X"C3",X"20",X"01",X"A1",X"03",X"3E",X"8F",X"C3",X"05",X"DE",X"A1",X"C3",X"3D",X"01",X"E0",X"32",
		X"11",X"40",X"0B",X"98",X"17",X"21",X"C3",X"2F",X"3E",X"04",X"32",X"01",X"20",X"E2",X"08",X"CD",
		X"A7",X"20",X"F8",X"C2",X"CD",X"01",X"05",X"EC",X"01",X"D5",X"32",X"97",X"20",X"E2",X"E1",X"3A",
		X"02",X"AD",X"00",X"00",X"0D",X"CD",X"11",X"40",X"E0",X"3A",X"A7",X"20",X"CC",X"C2",X"C3",X"01",
		X"09",X"F1",X"73",X"CD",X"11",X"04",X"22",X"ED",X"0B",X"90",X"17",X"21",X"0E",X"2F",X"CD",X"08",
		X"08",X"11",X"0E",X"23",X"CD",X"F7",X"05",X"CF",X"50",X"0E",X"22",X"CD",X"21",X"02",X"21",X"08",
		X"32",X"3D",X"20",X"E1",X"CC",X"C3",X"00",X"01",X"01",X"3E",X"F5",X"32",X"C3",X"20",X"03",X"29",
		X"15",X"0E",X"11",X"04",X"DE",X"CD",X"C3",X"05",X"06",X"18",X"06",X"C9",X"0C",X"00",X"26",X"04",
		X"F1",X"CD",X"06",X"09",X"DF",X"06",X"C2",X"05",X"04",X"EE",X"00",X"21",X"C3",X"21",X"00",X"51",
		X"15",X"21",X"0E",X"2A",X"C3",X"0F",X"05",X"44",X"06",X"1D",X"0E",X"C9",X"C3",X"15",X"05",X"44",
		X"32",X"97",X"20",X"F5",X"53",X"C3",X"C2",X"05",X"01",X"3E",X"F5",X"32",X"C3",X"20",X"08",X"3F",
		X"C3",X"06",X"05",X"27",X"41",X"CD",X"D3",X"40",X"05",X"1E",X"AD",X"3A",X"A7",X"20",X"38",X"CA",
		X"40",X"CD",X"CD",X"0B",X"0B",X"48",X"22",X"C9",X"00",X"01",X"00",X"00",X"CD",X"00",X"0B",X"20",
		X"3E",X"20",X"32",X"01",X"20",X"CD",X"C9",X"E1",X"20",X"D3",X"CE",X"3A",X"3C",X"20",X"CE",X"32",
		X"06",X"12",X"CD",X"3A",X"A7",X"20",X"87",X"C2",X"32",X"00",X"22",X"CE",X"CD",X"32",X"C3",X"20",
		X"E6",X"01",X"CA",X"80",X"06",X"6E",X"32",X"97",X"3A",X"06",X"20",X"CE",X"61",X"C3",X"DB",X"05",
		X"77",X"FC",X"A5",X"C3",X"BC",X"18",X"B1",X"D2",X"20",X"CD",X"6E",X"C3",X"EB",X"06",X"E6",X"7E",
		X"B5",X"D2",X"2F",X"06",X"85",X"3C",X"E0",X"FE",X"2F",X"06",X"84",X"3C",X"02",X"FE",X"BD",X"C9",
		X"11",X"06",X"01",X"0C",X"C0",X"21",X"06",X"20",X"94",X"C9",X"A4",X"C3",X"95",X"06",X"AE",X"C3",
		X"E6",X"20",X"A7",X"01",X"C3",X"C0",X"19",X"5C",X"EF",X"0C",X"C8",X"C3",X"3D",X"05",X"EE",X"32",
		X"8F",X"CD",X"67",X"04",X"8D",X"CD",X"84",X"04",X"CB",X"CD",X"C3",X"09",X"04",X"BB",X"23",X"3E",
		X"3F",X"C3",X"00",X"08",X"1C",X"00",X"FF",X"38",X"C3",X"67",X"0C",X"AA",X"CD",X"0A",X"09",X"CB",
		X"FF",X"46",X"00",X"00",X"20",X"04",X"FF",X"FF",X"00",X"00",X"49",X"92",X"00",X"FF",X"62",X"00",
		X"07",X"A0",X"07",X"B0",X"07",X"C0",X"07",X"D0",X"07",X"60",X"07",X"76",X"07",X"80",X"07",X"90",
		X"40",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"40",X"01",X"00",X"40",X"FF",X"FF",X"40",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"20",X"50",X"88",X"FF",X"FF",X"50",X"88",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7C",X"10",X"10",X"FF",X"FF",X"10",X"10",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"08",X"14",X"22",X"FF",X"FF",X"14",X"22",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"04",X"04",X"FF",X"FF",X"04",X"04",X"00",
		X"04",X"FF",X"FF",X"04",X"04",X"04",X"04",X"FF",X"0E",X"1F",X"0E",X"FF",X"FF",X"0E",X"04",X"0E",
		X"1C",X"FF",X"FF",X"08",X"00",X"08",X"FF",X"FF",X"FF",X"04",X"00",X"04",X"FF",X"FF",X"1C",X"3E",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"38",X"7C",X"38",X"FF",X"FF",X"10",X"00",X"10",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"70",X"F8",X"70",X"FF",X"FF",X"20",X"00",X"20",
		X"00",X"40",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"E0",X"FC",X"00",X"07",X"E0",X"FF",X"FF",X"40",
		X"FF",X"00",X"00",X"80",X"FF",X"FF",X"FF",X"FF",X"E0",X"FE",X"03",X"3F",X"E0",X"FF",X"03",X"80",
		X"FF",X"01",X"00",X"00",X"00",X"01",X"FF",X"FF",X"80",X"F0",X"03",X"1F",X"80",X"FF",X"03",X"00",
		X"FF",X"02",X"00",X"00",X"00",X"02",X"FF",X"FF",X"00",X"80",X"07",X"0F",X"00",X"FF",X"07",X"00",
		X"FF",X"12",X"20",X"20",X"11",X"12",X"40",X"FF",X"80",X"40",X"0B",X"07",X"20",X"FF",X"01",X"00",
		X"86",X"CD",X"C3",X"0C",X"13",X"17",X"00",X"00",X"0C",X"C0",X"FF",X"08",X"11",X"FF",X"1C",X"B9",
		X"14",X"CD",X"3C",X"48",X"F6",X"32",X"C9",X"20",X"48",X"CD",X"C3",X"0B",X"00",X"F7",X"A0",X"FE",
		X"20",X"3E",X"EA",X"32",X"CD",X"20",X"40",X"3C",X"EA",X"3A",X"FE",X"20",X"DA",X"10",X"04",X"24",
		X"04",X"0B",X"45",X"CD",X"00",X"40",X"00",X"00",X"CD",X"00",X"48",X"14",X"F6",X"3A",X"C3",X"20",
		X"A7",X"20",X"40",X"CA",X"2A",X"04",X"20",X"A9",X"C8",X"C3",X"3A",X"18",X"20",X"E2",X"A5",X"2A",
		X"4E",X"D2",X"01",X"04",X"03",X"00",X"EB",X"CD",X"EF",X"3A",X"01",X"20",X"02",X"00",X"01",X"FE",
		X"A5",X"22",X"CD",X"20",X"0B",X"40",X"67",X"C3",X"3A",X"0B",X"20",X"E2",X"C2",X"A7",X"04",X"61",
		X"01",X"0C",X"0C",X"06",X"C0",X"21",X"EF",X"20",X"22",X"04",X"20",X"A9",X"48",X"CD",X"11",X"0B",
		X"04",X"75",X"C0",X"21",X"11",X"20",X"22",X"C0",X"C8",X"C3",X"06",X"18",X"DF",X"06",X"C2",X"05",
		X"D3",X"C9",X"DB",X"00",X"3E",X"01",X"6F",X"12",X"10",X"0E",X"22",X"CD",X"21",X"02",X"20",X"ED",
		X"D5",X"E5",X"80",X"11",X"19",X"00",X"D1",X"7E",X"30",X"E6",X"0F",X"0F",X"E6",X"B5",X"C9",X"0F",
		X"20",X"3E",X"01",X"D3",X"41",X"CD",X"C3",X"40",X"A7",X"E1",X"2A",X"C2",X"C3",X"19",X"1B",X"C6",
		X"38",X"C3",X"97",X"0B",X"EA",X"32",X"C3",X"20",X"00",X"4E",X"7E",X"23",X"00",X"BA",X"00",X"00",
		X"46",X"CD",X"00",X"40",X"3E",X"00",X"32",X"05",X"00",X"AF",X"ED",X"32",X"32",X"20",X"20",X"EE",
		X"88",X"CD",X"26",X"17",X"3A",X"20",X"22",X"00",X"22",X"00",X"3E",X"C9",X"32",X"01",X"20",X"DF",
		X"88",X"CD",X"C3",X"17",X"01",X"62",X"40",X"C3",X"CD",X"6F",X"18",X"8D",X"32",X"97",X"20",X"DF",
		X"46",X"41",X"CD",X"1A",X"41",X"3A",X"1A",X"46",X"11",X"48",X"20",X"A3",X"1A",X"46",X"3A",X"CD",
		X"46",X"20",X"CD",X"1A",X"41",X"4A",X"1A",X"46",X"3A",X"CD",X"21",X"41",X"20",X"AB",X"A3",X"11",
		X"4C",X"CD",X"CD",X"06",X"03",X"C6",X"06",X"3F",X"4A",X"CD",X"46",X"41",X"CD",X"1A",X"41",X"4A",
		X"21",X"04",X"30",X"17",X"70",X"11",X"CD",X"0B",X"00",X"00",X"00",X"00",X"3F",X"C3",X"0E",X"06",
		X"05",X"4A",X"CA",X"A7",X"06",X"38",X"2D",X"11",X"09",X"F1",X"AD",X"3A",X"FE",X"20",X"D2",X"02",
		X"06",X"30",X"74",X"11",X"21",X"0B",X"28",X"13",X"C3",X"09",X"06",X"28",X"F1",X"CD",X"C3",X"09",
		X"22",X"00",X"20",X"9F",X"C9",X"00",X"7A",X"C3",X"23",X"C3",X"31",X"06",X"20",X"9F",X"42",X"21",
		X"80",X"E6",X"6E",X"C2",X"11",X"06",X"20",X"B0",X"FE",X"06",X"D2",X"04",X"06",X"6E",X"FF",X"3E",
		X"FE",X"20",X"CA",X"01",X"05",X"BC",X"02",X"FE",X"D3",X"2A",X"CD",X"20",X"15",X"B4",X"CE",X"3A",
		X"3A",X"06",X"20",X"E3",X"3A",X"47",X"20",X"E4",X"C2",X"CA",X"21",X"05",X"29",X"9A",X"5F",X"C3",
		X"20",X"E6",X"A7",X"B0",X"A8",X"CA",X"C3",X"04",X"47",X"B0",X"E5",X"3A",X"B0",X"20",X"3A",X"47",
		X"C9",X"21",X"32",X"97",X"20",X"E6",X"80",X"21",X"00",X"98",X"32",X"97",X"20",X"E5",X"40",X"21",
		X"08",X"06",X"C9",X"EF",X"42",X"21",X"C3",X"3A",X"C9",X"21",X"A5",X"21",X"11",X"20",X"01",X"01",
		X"32",X"97",X"20",X"CE",X"71",X"C3",X"CD",X"06",X"05",X"86",X"83",X"21",X"C3",X"2B",X"05",X"86",
		X"01",X"0E",X"22",X"CD",X"C9",X"02",X"17",X"21",X"02",X"22",X"CE",X"21",X"11",X"20",X"22",X"CE",
		X"C3",X"09",X"05",X"F7",X"17",X"21",X"11",X"2F",X"11",X"2F",X"0B",X"90",X"08",X"0E",X"F1",X"CD",
		X"2E",X"15",X"03",X"11",X"0E",X"06",X"C3",X"09",X"0B",X"98",X"08",X"0E",X"F1",X"CD",X"21",X"09");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
