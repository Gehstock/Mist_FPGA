library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ps05 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ps05 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"7B",X"78",X"84",X"42",X"02",X"18",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"00",X"8B",X"78",X"00",X"FF",X"FE",X"00",X"00",X"00",X"01",X"02",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7B",X"28",
		X"28",X"E0",X"00",X"00",X"FD",X"00",X"80",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"00",X"00",X"00",X"00",X"03",X"80",X"28",X"00",X"02",X"00",X"00",X"CF",X"42",X"01",X"18",
		X"00",X"FE",X"00",X"00",X"E7",X"42",X"01",X"18",X"00",X"01",X"00",X"00",X"FE",X"42",X"01",X"12",
		X"13",X"43",X"00",X"01",X"00",X"FE",X"00",X"A0",X"32",X"19",X"43",X"00",X"03",X"00",X"FE",X"00",
		X"B0",X"78",X"23",X"43",X"00",X"03",X"00",X"FE",X"00",X"98",X"80",X"25",X"43",X"00",X"01",X"00",
		X"FE",X"00",X"A8",X"98",X"00",X"0A",X"00",X"FC",X"00",X"00",X"00",X"E4",X"48",X"01",X"08",X"00",
		X"00",X"FC",X"00",X"00",X"00",X"E4",X"48",X"01",X"08",X"00",X"00",X"00",X"FE",X"00",X"80",X"90",
		X"00",X"01",X"00",X"FE",X"00",X"80",X"90",X"00",X"03",X"00",X"FE",X"00",X"80",X"90",X"00",X"00",
		X"00",X"01",X"00",X"30",X"40",X"00",X"04",X"00",X"01",X"00",X"30",X"50",X"00",X"08",X"00",X"01",
		X"00",X"30",X"60",X"50",X"00",X"15",X"00",X"FC",X"00",X"00",X"00",X"E4",X"48",X"01",X"08",X"00",
		X"B2",X"47",X"01",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"E0",X"88",X"1A",X"46",X"02",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"30",X"E0",X"00",
		X"00",X"00",X"98",X"80",X"00",X"A8",X"98",X"00",X"B8",X"B0",X"00",X"C8",X"C8",X"00",X"D8",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"A0",X"90",X"00",X"B0",X"78",X"00",X"C0",X"60",X"00",X"D0",X"48",
		X"00",X"E0",X"30",X"00",X"00",X"00",X"00",X"01",X"68",X"F0",X"00",X"58",X"F0",X"00",X"40",X"F0",
		X"00",X"00",X"00",X"01",X"70",X"28",X"00",X"58",X"28",X"00",X"00",X"30",X"30",X"00",X"40",X"78",
		X"00",X"50",X"A8",X"00",X"58",X"58",X"00",X"48",X"38",X"00",X"00",X"00",X"00",X"00",X"01",X"03",
		X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"2E",X"00",X"00",X"02",X"2E",X"00",X"00",X"01",X"2E",
		X"00",X"91",X"44",X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"13",X"08",X"0B",X"13",X"1F",X"24",X"44",X"24",X"1F",X"7F",X"49",X"49",X"49",X"36",X"3E",X"41",
		X"41",X"41",X"22",X"7F",X"41",X"41",X"41",X"3E",X"7F",X"49",X"49",X"49",X"41",X"7F",X"48",X"48",
		X"48",X"40",X"3E",X"41",X"41",X"45",X"47",X"7F",X"08",X"08",X"08",X"7F",X"00",X"41",X"7F",X"41",
		X"00",X"02",X"01",X"01",X"01",X"7E",X"7F",X"08",X"14",X"22",X"41",X"7F",X"01",X"01",X"01",X"01",
		X"7F",X"20",X"18",X"20",X"7F",X"7F",X"10",X"08",X"04",X"7F",X"3E",X"41",X"41",X"41",X"3E",X"7F",
		X"48",X"48",X"48",X"30",X"3E",X"41",X"45",X"42",X"3D",X"7F",X"48",X"4C",X"4A",X"31",X"32",X"49",
		X"49",X"49",X"26",X"40",X"40",X"7F",X"40",X"40",X"7E",X"01",X"01",X"01",X"7E",X"7C",X"02",X"01",
		X"02",X"7C",X"7F",X"02",X"0C",X"02",X"7F",X"63",X"14",X"08",X"14",X"63",X"60",X"10",X"0F",X"10",
		X"60",X"43",X"45",X"49",X"51",X"61",X"00",X"00",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3E",X"45",X"49",X"51",X"3E",X"00",X"21",X"7F",X"01",X"00",X"23",X"45",X"49",X"49",X"31",X"42",
		X"41",X"49",X"59",X"66",X"0C",X"14",X"24",X"7F",X"04",X"72",X"51",X"51",X"51",X"4E",X"1E",X"29",
		X"49",X"49",X"46",X"40",X"47",X"48",X"50",X"60",X"36",X"49",X"49",X"49",X"36",X"31",X"49",X"49",
		X"4A",X"3C",X"08",X"14",X"22",X"41",X"00",X"00",X"41",X"22",X"14",X"08",X"14",X"14",X"14",X"14",
		X"14",X"22",X"14",X"7F",X"14",X"22",X"18",X"18",X"18",X"18",X"18",X"08",X"08",X"08",X"08",X"08",
		X"20",X"40",X"4D",X"50",X"20",X"00",X"00",X"79",X"00",X"79",X"00",X"00",X"00",X"00",X"0C",X"40",
		X"40",X"40",X"40",X"40",X"01",X"1C",X"3C",X"78",X"60",X"0F",X"14",X"12",X"07",X"02",X"11",X"04",
		X"03",X"08",X"13",X"1B",X"00",X"00",X"70",X"00",X"E8",X"00",X"E8",X"0B",X"F8",X"1B",X"F8",X"0B",
		X"F8",X"3F",X"F8",X"0F",X"F8",X"03",X"F8",X"00",X"F8",X"00",X"F8",X"00",X"F8",X"00",X"F8",X"00",
		X"F8",X"00",X"F0",X"00",X"70",X"00",X"70",X"00",X"70",X"00",X"60",X"00",X"60",X"00",X"F0",X"00",
		X"F8",X"01",X"60",X"00",X"03",X"3C",X"03",X"06",X"1F",X"1F",X"2F",X"6F",X"3F",X"1F",X"0F",X"0F",
		X"0F",X"0F",X"0E",X"04",X"0E",X"00",X"00",X"92",X"54",X"38",X"FE",X"38",X"54",X"92",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"34",X"1C",X"48",X"69",
		X"3B",X"3F",X"1E",X"0C",X"08",X"08",X"08",X"08",X"08",X"0C",X"1C",X"1E",X"3F",X"6B",X"49",X"08",
		X"18",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"0F",X"0F",X"0F",X"0F",X"0F",X"3F",X"3F",X"7F",X"FF",X"3F",X"3F",X"0F",X"0F",X"0F",X"06",
		X"36",X"0F",X"36",X"00",X"00",X"02",X"03",X"01",X"02",X"04",X"04",X"03",X"02",X"01",X"00",X"00",
		X"01",X"02",X"03",X"04",X"03",X"03",X"02",X"01",X"01",X"02",X"00",X"00",X"01",X"04",X"02",X"00",
		X"01",X"02",X"03",X"FF",X"FF",X"FF",X"D3",X"3C",X"7D",X"97",X"FF",X"7F",X"BB",X"FE",X"3B",X"E7",
		X"FC",X"1F",X"EF",X"F3",X"0D",X"E7",X"F9",X"04",X"FF",X"DF",X"02",X"EF",X"EC",X"03",X"6F",X"E6",
		X"60",X"F7",X"FF",X"10",X"F7",X"DF",X"09",X"DF",X"1F",X"3F",X"1F",X"0F",X"E4",X"BF",X"03",X"08",
		X"FF",X"01",X"10",X"FF",X"77",X"67",X"33",X"3F",X"77",X"7F",X"3F",X"9F",X"5B",X"FB",X"4F",X"9B",
		X"37",X"2F",X"6F",X"77",X"67",X"EF",X"FF",X"9F",X"DF",X"F7",X"F7",X"FF",X"01",X"FF",X"01",X"BF",
		X"01",X"7F",X"03",X"BF",X"03",X"FF",X"07",X"FB",X"0F",X"E7",X"0E",X"DF",X"1C",X"FB",X"37",X"73",
		X"7D",X"9F",X"7C",X"BB",X"7F",X"FF",X"77",X"FF",X"36",X"DF",X"3C",X"E7",X"1D",X"EF",X"0B",X"DF",
		X"0F",X"DB",X"07",X"E7",X"07",X"F5",X"03",X"F5",X"01",X"FF",X"01",X"FF",X"00",X"40",X"00",X"EF",
		X"01",X"20",X"00",X"DF",X"07",X"10",X"03",X"EF",X"07",X"90",X"04",X"F7",X"0F",X"7E",X"00",X"7F",
		X"9B",X"C7",X"00",X"4F",X"F2",X"81",X"19",X"9F",X"FD",X"03",X"07",X"BF",X"5F",X"0F",X"08",X"BF",
		X"FD",X"3C",X"00",X"5F",X"FF",X"7F",X"00",X"2F",X"F3",X"EF",X"01",X"DF",X"1F",X"DB",X"0F",X"FF",
		X"B7",X"7B",X"3C",X"FF",X"F9",X"71",X"FB",X"FF",X"FF",X"FF",X"FF",X"00",X"C4",X"20",X"38",X"00",
		X"01",X"C4",X"01",X"12",X"02",X"02",X"D5",X"01",X"0A",X"02",X"10",X"C4",X"01",X"38",X"02",X"02",
		X"C4",X"01",X"12",X"01",X"01",X"D5",X"01",X"0C",X"04",X"03",X"D8",X"01",X"10",X"04",X"06",X"C4",
		X"0A",X"38",X"07",X"06",X"C4",X"01",X"04",X"07",X"06",X"DE",X"02",X"04",X"07",X"04",X"C4",X"02",
		X"38",X"07",X"03",X"C4",X"01",X"12",X"06",X"03",X"D4",X"01",X"08",X"01",X"11",X"C4",X"0F",X"38",
		X"06",X"FF",X"0B",X"04",X"15",X"04",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"06",
		X"07",X"1F",X"37",X"3F",X"37",X"1F",X"1F",X"2F",X"27",X"0F",X"07",X"07",X"0E",X"06",X"04",X"04",
		X"06",X"0E",X"07",X"07",X"0F",X"27",X"2F",X"1F",X"1F",X"37",X"3F",X"37",X"1F",X"07",X"06",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"0D",X"12",X"04",X"11",X"13",X"1B",X"1B",X"02",
		X"0E",X"08",X"0D",X"3C",X"42",X"99",X"A5",X"A5",X"81",X"42",X"3C",X"13",X"00",X"08",X"13",X"0E",
		X"1B",X"02",X"0E",X"11",X"0F",X"0E",X"11",X"00",X"13",X"08",X"0E",X"0D",X"1B",X"1D",X"25",X"24",
		X"1C",X"20",X"20",X"20",X"10",X"10",X"40",X"40",X"40",X"80",X"00",X"00",X"20",X"20",X"10",X"20",
		X"40",X"80",X"00",X"20",X"10",X"40",X"80",X"40",X"20",X"10",X"00",X"40",X"20",X"80",X"20",X"40",
		X"10",X"81",X"80",X"82",X"44",X"08",X"08",X"18",X"1C",X"04",X"01",X"B0",X"83",X"19",X"15",X"6A",
		X"4C",X"D0",X"AA",X"C0",X"1F",X"68",X"3D",X"CC",X"1D",X"58",X"42",X"BC",X"8F",X"20",X"1B",X"D3",
		X"06",X"99",X"3A",X"20",X"08",X"B4",X"12",X"A1",X"22",X"10",X"00",X"10",X"01",X"C2",X"04",X"01",
		X"C4",X"03",X"03",X"03",X"28",X"10",X"38",X"10",X"28",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"00",X"24",X"10",X"2A",X"1C",X"10",X"0A",X"24",X"00",X"08",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"20",X"08",X"24",X"21",X"08",X"3A",X"A8",X"2C",X"64",X"54",X"6C",X"28",X"A9",X"38",
		X"20",X"22",X"48",X"51",X"12",X"08",X"44",X"00",X"00",X"06",X"0F",X"0F",X"1E",X"12",X"00",X"01",
		X"03",X"26",X"62",X"70",X"3C",X"38",X"91",X"01",X"0F",X"0F",X"0F",X"06",X"00",X"00",X"00",X"00",
		X"00",X"81",X"52",X"08",X"60",X"D1",X"82",X"28",X"42",X"10",X"18",X"5A",X"10",X"04",X"30",X"42",
		X"83",X"10",X"08",X"0A",X"20",X"44",X"C2",X"93",X"01",X"81",X"54",X"5C",X"3E",X"7C",X"1A",X"80",
		X"11",X"1A",X"C7",X"01",X"2A",X"04",X"18",X"C9",X"01",X"22",X"06",X"13",X"C9",X"01",X"1A",X"03",
		X"11",X"C9",X"01",X"1A",X"02",X"0E",X"C9",X"01",X"1A",X"04",X"0C",X"C9",X"01",X"1A",X"03",X"0A",
		X"C9",X"01",X"1A",X"01",X"08",X"C9",X"01",X"1A",X"02",X"15",X"C9",X"02",X"1A",X"05",X"FF",X"29",
		X"12",X"02",X"0E",X"11",X"04",X"1B",X"00",X"03",X"15",X"00",X"0D",X"02",X"04",X"1B",X"13",X"00",
		X"01",X"0B",X"04",X"29",X"29",X"04",X"17",X"13",X"11",X"00",X"28",X"21",X"1C",X"1C",X"1C",X"0F",
		X"0E",X"08",X"0D",X"13",X"29",X"15",X"2C",X"28",X"2C",X"2C",X"2C",X"1B",X"0F",X"0E",X"08",X"0D",
		X"13",X"13",X"2C",X"28",X"2C",X"2C",X"2C",X"1B",X"0F",X"0E",X"08",X"0D",X"13",X"11",X"2C",X"28",
		X"1D",X"1C",X"1C",X"1B",X"0F",X"0E",X"08",X"0D",X"13",X"0E",X"2C",X"28",X"1B",X"21",X"1C",X"1B",
		X"0F",X"0E",X"08",X"0D",X"13",X"0C",X"2C",X"28",X"1B",X"21",X"1C",X"1B",X"0F",X"0E",X"08",X"0D",
		X"13",X"0A",X"2C",X"28",X"1B",X"1F",X"1C",X"1B",X"0F",X"0E",X"08",X"0D",X"13",X"08",X"2C",X"28",
		X"1B",X"1D",X"1C",X"1B",X"0F",X"0E",X"08",X"0D",X"13",X"FF",X"91",X"24",X"12",X"5C",X"98",X"22",
		X"74",X"81",X"08",X"00",X"22",X"3B",X"12",X"00",X"01",X"03",X"13",X"39",X"29",X"19",X"88",X"80",
		X"46",X"8E",X"0C",X"18",X"00",X"00",X"65",X"30",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"00",X"08",X"00",X"74",X"0C",X"F0",X"0E",X"E0",X"05",X"E0",X"03",X"C0",X"03",X"E0",X"17",
		X"70",X"0E",X"38",X"7C",X"18",X"1C",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"0C",X"04",X"0E",X"3A",X"07",X"F8",X"02",X"F0",X"01",X"E0",X"03",X"E0",X"27",X"70",X"0E",
		X"70",X"78",X"30",X"18",X"38",X"08",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",
		X"30",X"00",X"00",X"00",X"39",X"08",X"FE",X"0C",X"FF",X"0F",X"0E",X"0B",X"71",X"04",X"70",X"04",
		X"30",X"00",X"30",X"00",X"30",X"00",X"30",X"00",X"00",X"00",X"30",X"00",X"30",X"00",X"30",X"00",
		X"30",X"00",X"70",X"04",X"71",X"04",X"0E",X"0B",X"FF",X"0F",X"FE",X"0C",X"39",X"08",X"00",X"00",
		X"30",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C4",X"21",X"F8",X"33",X"FC",X"3F",X"F8",X"1F",X"24",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",
		X"08",X"00",X"34",X"00",X"70",X"00",X"F0",X"01",X"E0",X"03",X"D0",X"03",X"80",X"03",X"00",X"27",
		X"00",X"3E",X"00",X"1C",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"15",X"00",X"0E",
		X"00",X"0E",X"00",X"0F",X"00",X"0E",X"00",X"1E",X"00",X"1E",X"00",X"1E",X"00",X"1E",X"00",X"06",
		X"00",X"06",X"00",X"06",X"00",X"0E",X"00",X"1C",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"10",
		X"80",X"2E",X"00",X"0F",X"80",X"07",X"C0",X"03",X"E0",X"03",X"F0",X"01",X"38",X"00",X"1C",X"00",
		X"18",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"12",X"FC",X"0F",X"FE",X"1F",X"E6",X"0F",X"C2",X"11",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",
		X"38",X"00",X"7C",X"00",X"E4",X"00",X"C0",X"01",X"C0",X"0B",X"C0",X"07",X"80",X"0F",X"00",X"0E",
		X"00",X"1C",X"00",X"10",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"0E",
		X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0E",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0E",
		X"00",X"1E",X"00",X"0E",X"00",X"0E",X"00",X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0C",X"00",X"18",X"00",X"38",X"00",X"1C",X"80",X"0F",X"C0",X"07",X"C0",X"03",X"E0",X"01",
		X"F0",X"00",X"74",X"01",X"08",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FB",X"00",
		X"FB",X"00",X"FB",X"00",X"FB",X"FB",X"00",X"FB",X"05",X"FB",X"05",X"00",X"05",X"05",X"00",X"05",
		X"FB",X"05",X"02",X"00",X"02",X"01",X"02",X"02",X"02",X"03",X"02",X"02",X"02",X"03",X"01",X"04",
		X"01",X"05",X"03",X"06",X"03",X"07",X"03",X"08",X"03",X"09",X"03",X"0A",X"03",X"0B",X"03",X"04",
		X"03",X"05",X"09",X"06",X"03",X"07",X"03",X"08",X"03",X"09",X"10",X"0A",X"03",X"0B",X"03",X"04",
		X"03",X"05",X"07",X"06",X"FF",X"04",X"05",X"15",X"06",X"03",X"07",X"06",X"08",X"03",X"09",X"10",
		X"0A",X"03",X"0B",X"03",X"04",X"03",X"05",X"03",X"06",X"03",X"07",X"03",X"08",X"03",X"09",X"08");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
