library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity bg_graphx_2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of bg_graphx_2 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"3F",X"CF",X"FF",X"EF",X"FF",X"AF",X"AF",X"AF",X"AF",
		X"6F",X"DF",X"6F",X"DF",X"EF",X"FF",X"CF",X"FF",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"FF",X"7F",X"0F",X"6F",X"FF",X"6F",X"CF",X"7F",
		X"CF",X"7F",X"CF",X"6F",X"FF",X"6F",X"FF",X"7F",X"8F",X"1F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"02",X"02",X"06",X"06",X"0E",X"0E",X"06",X"06",X"06",
		X"00",X"00",X"00",X"00",X"00",X"86",X"0E",X"CF",X"04",X"C8",X"00",X"4F",X"0F",X"C0",X"00",X"C0",
		X"00",X"00",X"00",X"00",X"01",X"09",X"0A",X"02",X"06",X"00",X"00",X"0F",X"0F",X"00",X"03",X"00",
		X"00",X"08",X"E0",X"02",X"F0",X"30",X"F4",X"74",X"04",X"C6",X"A6",X"87",X"A7",X"A6",X"A6",X"A6",
		X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"C2",X"00",X"C0",X"02",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"50",X"D0",X"50",X"D0",X"40",X"90",X"01",X"C0",X"F0",X"70",X"F0",X"30",X"E0",X"08",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"30",X"F0",X"FA",X"D0",X"B0",X"10",X"D0",
		X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"20",X"00",
		X"18",X"D0",X"D0",X"B0",X"F8",X"F0",X"F0",X"32",X"04",X"04",X"02",X"02",X"00",X"00",X"00",X"08",
		X"00",X"01",X"00",X"01",X"00",X"00",X"04",X"02",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"08",
		X"21",X"20",X"80",X"30",X"00",X"10",X"00",X"40",X"00",X"00",X"0C",X"1E",X"0E",X"0F",X"0F",X"0F",
		X"50",X"00",X"00",X"08",X"00",X"08",X"08",X"0C",X"0E",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0E",X"0B",X"0A",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"CF",
		X"C7",X"F5",X"E5",X"FF",X"6F",X"0F",X"EF",X"7F",X"6F",X"FF",X"6F",X"CF",X"6F",X"CF",X"6F",X"1F",
		X"0F",X"0A",X"0A",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"1F",X"0F",
		X"FF",X"35",X"F5",X"FF",X"FF",X"FF",X"0F",X"FF",X"AF",X"8F",X"AF",X"AF",X"FF",X"BF",X"6F",X"8F",
		X"60",X"10",X"62",X"C2",X"68",X"C1",X"6A",X"F0",X"E8",X"71",X"61",X"04",X"E0",X"F1",X"C0",X"F4",
		X"0C",X"C9",X"0A",X"0D",X"04",X"0D",X"04",X"0E",X"0D",X"0A",X"05",X"09",X"04",X"0A",X"05",X"0E",
		X"6F",X"8D",X"FD",X"BF",X"AF",X"A7",X"AF",X"8F",X"0F",X"FF",X"FF",X"FE",X"FF",X"FB",X"FF",X"3F",
		X"1F",X"0E",X"0D",X"0E",X"0F",X"0F",X"0F",X"0E",X"0E",X"0B",X"0F",X"0F",X"0D",X"0F",X"0F",X"0D",
		X"08",X"02",X"08",X"04",X"02",X"00",X"00",X"00",X"00",X"00",X"01",X"08",X"00",X"00",X"00",X"00",
		X"02",X"05",X"0B",X"02",X"F4",X"30",X"F9",X"F0",X"90",X"10",X"10",X"12",X"51",X"3E",X"70",X"B0",
		X"07",X"0E",X"0D",X"0D",X"0F",X"0B",X"0F",X"05",X"04",X"00",X"09",X"00",X"0D",X"42",X"08",X"00",
		X"0F",X"0B",X"87",X"06",X"0B",X"03",X"1D",X"03",X"11",X"0C",X"1B",X"82",X"9A",X"10",X"15",X"68",
		X"70",X"B0",X"50",X"31",X"13",X"13",X"93",X"17",X"FF",X"FF",X"FF",X"3F",X"0F",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"06",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"10",X"60",X"90",X"10",X"10",X"80",X"10",X"00",X"10",X"01",X"03",X"03",X"87",X"0F",X"0F",X"0F",
		X"00",X"01",X"02",X"41",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",
		X"0F",X"EF",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"EA",X"CB",X"FE",
		X"EF",X"FF",X"7F",X"8F",X"7F",X"FF",X"FF",X"FF",X"7F",X"FF",X"6F",X"CF",X"4F",X"C5",X"05",X"07",
		X"3F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"3F",X"0A",X"FA",X"0F",
		X"FF",X"FF",X"1F",X"EF",X"4F",X"8F",X"2F",X"9F",X"AF",X"8F",X"AF",X"AF",X"FF",X"B5",X"05",X"9F",
		X"0B",X"0D",X"4F",X"CF",X"6D",X"CD",X"76",X"FE",X"FD",X"FF",X"7F",X"FF",X"7B",X"8D",X"EF",X"F7",
		X"CF",X"FE",X"07",X"EF",X"06",X"0F",X"0F",X"07",X"0F",X"05",X"0F",X"0E",X"07",X"0B",X"0F",X"EE",
		X"0F",X"96",X"FB",X"B7",X"AD",X"AF",X"A5",X"8F",X"2B",X"9B",X"47",X"8D",X"1B",X"EB",X"F7",X"FF",
		X"F7",X"03",X"31",X"00",X"00",X"00",X"0B",X"08",X"00",X"05",X"09",X"09",X"00",X"02",X"38",X"03",
		X"0B",X"87",X"0F",X"CD",X"07",X"0A",X"0E",X"07",X"0B",X"05",X"0A",X"07",X"03",X"00",X"70",X"00",
		X"FF",X"83",X"FE",X"FD",X"03",X"0F",X"00",X"02",X"0E",X"80",X"22",X"C1",X"F0",X"F0",X"B0",X"F0",
		X"3F",X"0F",X"76",X"07",X"0B",X"04",X"0D",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"30",
		X"B1",X"30",X"F2",X"10",X"E1",X"10",X"F0",X"10",X"B0",X"10",X"B0",X"10",X"D0",X"10",X"D0",X"10",
		X"BF",X"FF",X"FE",X"F7",X"2F",X"CF",X"0F",X"8B",X"0B",X"0E",X"05",X"09",X"F0",X"F0",X"F0",X"80",
		X"73",X"0F",X"07",X"0F",X"0F",X"0F",X"07",X"07",X"0D",X"0B",X"00",X"08",X"00",X"C0",X"00",X"80",
		X"DF",X"1F",X"DB",X"17",X"BF",X"1B",X"BF",X"1B",X"F7",X"1C",X"EA",X"14",X"F0",X"10",X"B0",X"30",
		X"0F",X"3F",X"0B",X"0F",X"0F",X"0D",X"0E",X"07",X"0F",X"0D",X"0E",X"09",X"74",X"08",X"30",X"00",
		X"0F",X"0F",X"0F",X"0D",X"0F",X"07",X"0F",X"0F",X"0E",X"0F",X"0B",X"07",X"0E",X"0B",X"0B",X"0F",
		X"0D",X"07",X"0E",X"0D",X"0F",X"FF",X"0F",X"1E",X"0B",X"D5",X"0D",X"F7",X"0B",X"DD",X"0B",X"1E",
		X"0F",X"0B",X"0B",X"0F",X"0E",X"0F",X"0E",X"0F",X"0F",X"0F",X"0F",X"0B",X"0F",X"07",X"0E",X"0F",
		X"0F",X"0D",X"EB",X"0D",X"FF",X"1E",X"8F",X"FD",X"5D",X"C7",X"5F",X"1F",X"FB",X"5F",X"0F",X"7B",
		X"0F",X"1F",X"07",X"D3",X"01",X"F0",X"00",X"D0",X"01",X"13",X"01",X"F1",X"00",X"05",X"0F",X"0F",
		X"0B",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"0F",
		X"0F",X"7F",X"F6",X"50",X"50",X"10",X"50",X"C0",X"80",X"F0",X"F0",X"10",X"E0",X"00",X"05",X"0F",
		X"0F",X"0E",X"0C",X"08",X"0C",X"08",X"00",X"00",X"08",X"08",X"00",X"00",X"08",X"08",X"0C",X"0E",
		X"00",X"00",X"01",X"0B",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"C0",X"90",X"C0",X"F3",X"7F",X"7F",X"1F",X"EF",X"1F",X"CF",X"5F",X"8F",X"FF",X"FF",X"7F",X"FF",
		X"00",X"00",X"00",X"0C",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"F0",X"06",X"FF",X"0F",X"EF",X"1F",X"CF",X"1F",X"9F",X"1F",X"9F",X"1F",X"BF",X"1F",X"AF",X"1F",
		X"AF",X"AF",X"AF",X"AF",X"FF",X"EF",X"FF",X"CF",X"3F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"FF",X"CF",X"FF",X"EF",X"DF",X"6F",X"DF",X"6F",
		X"7F",X"CF",X"6F",X"FF",X"6F",X"0F",X"7F",X"FF",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"1F",X"8F",X"7F",X"FF",X"6F",X"FF",X"6F",X"CF",X"7F",X"CF",
		X"06",X"06",X"06",X"0E",X"0E",X"06",X"06",X"02",X"02",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"00",X"C0",X"0F",X"4F",X"00",X"C8",X"04",X"CF",X"0E",X"86",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"00",X"0F",X"0F",X"00",X"00",X"06",X"02",X"0A",X"09",X"01",X"00",X"00",X"00",X"00",
		X"A6",X"A6",X"A6",X"A7",X"87",X"A6",X"C6",X"04",X"74",X"F4",X"30",X"F0",X"02",X"E0",X"08",X"00",
		X"00",X"00",X"00",X"00",X"80",X"02",X"C0",X"00",X"C2",X"00",X"40",X"00",X"40",X"00",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"08",X"E0",X"30",X"F0",X"70",X"F0",X"C0",X"01",X"90",X"40",X"D0",X"50",X"D0",X"50",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",
		X"D0",X"10",X"B0",X"D0",X"FA",X"F0",X"30",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",
		X"00",X"20",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"01",X"00",X"00",X"00",
		X"08",X"00",X"00",X"00",X"02",X"02",X"04",X"04",X"32",X"F0",X"F0",X"F8",X"B0",X"D0",X"D0",X"18",
		X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"02",X"04",X"00",X"00",X"01",X"00",X"01",X"00",
		X"0F",X"0F",X"0F",X"0E",X"1E",X"0C",X"00",X"00",X"40",X"00",X"10",X"00",X"30",X"80",X"20",X"21",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0E",X"0C",X"08",X"08",X"00",X"08",X"00",X"00",X"50",
		X"CF",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0A",X"0B",X"0E",
		X"1F",X"6F",X"CF",X"6F",X"CF",X"6F",X"FF",X"6F",X"7F",X"EF",X"0F",X"6F",X"FF",X"E5",X"F5",X"C7",
		X"0F",X"1F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0A",X"0A",X"0F",
		X"8F",X"6F",X"BF",X"FF",X"AF",X"AF",X"8F",X"AF",X"FF",X"0F",X"FF",X"FF",X"FF",X"F5",X"35",X"FF",
		X"F4",X"C0",X"F1",X"E0",X"04",X"61",X"71",X"E8",X"F0",X"6A",X"C1",X"68",X"C2",X"62",X"10",X"60",
		X"0E",X"05",X"0A",X"04",X"09",X"05",X"0A",X"0D",X"0E",X"04",X"0D",X"04",X"0D",X"0A",X"C9",X"0C",
		X"3F",X"FF",X"FB",X"FF",X"FE",X"FF",X"FF",X"0F",X"8F",X"AF",X"A7",X"AF",X"BF",X"FD",X"8D",X"6F",
		X"0D",X"0F",X"0F",X"0D",X"0F",X"0F",X"0B",X"0E",X"0E",X"0F",X"0F",X"0F",X"0E",X"0D",X"0E",X"1F",
		X"00",X"00",X"00",X"00",X"08",X"01",X"00",X"00",X"00",X"00",X"00",X"02",X"04",X"08",X"02",X"08",
		X"B0",X"70",X"3E",X"51",X"12",X"10",X"10",X"90",X"F0",X"F9",X"30",X"F4",X"02",X"0B",X"05",X"02",
		X"00",X"08",X"42",X"0D",X"00",X"09",X"00",X"04",X"05",X"0F",X"0B",X"0F",X"0D",X"0D",X"0E",X"07",
		X"68",X"15",X"10",X"9A",X"82",X"1B",X"0C",X"11",X"03",X"1D",X"03",X"0B",X"06",X"87",X"0B",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"3F",X"FF",X"FF",X"FF",X"17",X"93",X"13",X"13",X"31",X"50",X"B0",X"70",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"06",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"87",X"03",X"03",X"01",X"10",X"00",X"10",X"80",X"10",X"10",X"90",X"60",X"10",
		X"07",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"41",X"02",X"01",X"00",
		X"FE",X"CB",X"EA",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"EF",X"0F",
		X"07",X"05",X"C5",X"4F",X"CF",X"6F",X"FF",X"7F",X"FF",X"FF",X"FF",X"7F",X"8F",X"7F",X"FF",X"EF",
		X"0F",X"FA",X"0A",X"3F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"3F",
		X"9F",X"05",X"B5",X"FF",X"AF",X"AF",X"8F",X"AF",X"9F",X"2F",X"8F",X"4F",X"EF",X"1F",X"FF",X"FF",
		X"F7",X"EF",X"8D",X"7B",X"FF",X"7F",X"FF",X"FD",X"FE",X"76",X"CD",X"6D",X"CF",X"4F",X"0D",X"0B",
		X"EE",X"0F",X"0B",X"07",X"0E",X"0F",X"05",X"0F",X"07",X"0F",X"0F",X"06",X"EF",X"07",X"FE",X"CF",
		X"FF",X"F7",X"EB",X"1B",X"8D",X"47",X"9B",X"2B",X"8F",X"A5",X"AF",X"AD",X"B7",X"FB",X"96",X"0F",
		X"03",X"38",X"02",X"00",X"09",X"09",X"05",X"00",X"08",X"0B",X"00",X"00",X"00",X"31",X"03",X"F7",
		X"00",X"70",X"00",X"03",X"07",X"0A",X"05",X"0B",X"07",X"0E",X"0A",X"07",X"CD",X"0F",X"87",X"0B",
		X"F0",X"B0",X"F0",X"F0",X"C1",X"22",X"80",X"0E",X"02",X"00",X"0F",X"03",X"FD",X"FE",X"83",X"FF",
		X"30",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"0D",X"04",X"0B",X"07",X"76",X"0F",X"3F",
		X"10",X"D0",X"10",X"D0",X"10",X"B0",X"10",X"B0",X"10",X"F0",X"10",X"E1",X"10",X"F2",X"30",X"B1",
		X"80",X"F0",X"F0",X"F0",X"09",X"05",X"0E",X"0B",X"8B",X"0F",X"CF",X"2F",X"F7",X"FE",X"FF",X"BF",
		X"80",X"00",X"C0",X"00",X"08",X"00",X"0B",X"0D",X"07",X"07",X"0F",X"0F",X"0F",X"07",X"0F",X"73",
		X"30",X"B0",X"10",X"F0",X"14",X"EA",X"1C",X"F7",X"1B",X"BF",X"1B",X"BF",X"17",X"DB",X"1F",X"DF",
		X"00",X"30",X"08",X"74",X"09",X"0E",X"0D",X"0F",X"07",X"0E",X"0D",X"0F",X"0F",X"0B",X"3F",X"0F",
		X"0F",X"0B",X"0B",X"0E",X"07",X"0B",X"0F",X"0E",X"0F",X"0F",X"07",X"0F",X"0D",X"0F",X"0F",X"0F",
		X"1E",X"0B",X"DD",X"0B",X"F7",X"0D",X"D5",X"0B",X"1E",X"0F",X"FF",X"0F",X"0D",X"0E",X"07",X"0D",
		X"0F",X"0E",X"07",X"0F",X"0B",X"0F",X"0F",X"0F",X"0F",X"0E",X"0F",X"0E",X"0F",X"0B",X"0B",X"0F",
		X"7B",X"0F",X"5F",X"FB",X"1F",X"5F",X"C7",X"5D",X"FD",X"8F",X"1E",X"FF",X"0D",X"EB",X"0D",X"0F",
		X"0F",X"0F",X"05",X"00",X"F1",X"01",X"13",X"01",X"D0",X"00",X"F0",X"01",X"D3",X"07",X"1F",X"0F",
		X"0F",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"0B",
		X"0F",X"05",X"00",X"E0",X"10",X"F0",X"F0",X"80",X"C0",X"50",X"10",X"50",X"50",X"F6",X"7F",X"0F",
		X"0E",X"0C",X"08",X"08",X"00",X"00",X"08",X"08",X"00",X"00",X"08",X"0C",X"08",X"0C",X"0E",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0B",X"01",X"00",X"00",
		X"FF",X"7F",X"FF",X"FF",X"8F",X"5F",X"CF",X"1F",X"EF",X"1F",X"7F",X"7F",X"F3",X"C0",X"90",X"C0",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0C",X"00",X"00",X"00",
		X"1F",X"AF",X"1F",X"BF",X"1F",X"9F",X"1F",X"9F",X"1F",X"CF",X"1F",X"EF",X"0F",X"FF",X"06",X"F0");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
