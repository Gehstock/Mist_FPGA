library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity fg_sp_graphx_3 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of fg_sp_graphx_3 is
	type rom is array(0 to  7167) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"3E",X"61",X"41",X"43",X"3E",X"1C",
		X"00",X"00",X"40",X"42",X"7F",X"7F",X"40",X"40",X"00",X"62",X"73",X"79",X"59",X"5D",X"4F",X"46",
		X"00",X"20",X"61",X"49",X"4D",X"4F",X"7B",X"31",X"00",X"18",X"1C",X"16",X"13",X"7F",X"7F",X"10",
		X"00",X"27",X"67",X"45",X"45",X"45",X"7D",X"38",X"00",X"3C",X"7E",X"4B",X"49",X"49",X"79",X"30",
		X"00",X"03",X"03",X"71",X"79",X"0D",X"07",X"03",X"00",X"36",X"4F",X"4D",X"59",X"59",X"76",X"30",
		X"00",X"06",X"4F",X"49",X"49",X"69",X"3F",X"1E",X"00",X"7C",X"7E",X"13",X"11",X"13",X"7E",X"7C",
		X"00",X"7F",X"7F",X"49",X"49",X"49",X"7F",X"36",X"00",X"1C",X"3E",X"63",X"41",X"41",X"63",X"22",
		X"00",X"7F",X"7F",X"41",X"41",X"63",X"3E",X"1C",X"00",X"00",X"7F",X"7F",X"49",X"49",X"49",X"41",
		X"00",X"7F",X"7F",X"09",X"09",X"09",X"09",X"01",X"00",X"1C",X"3E",X"63",X"41",X"49",X"79",X"79",
		X"00",X"7F",X"7F",X"08",X"08",X"08",X"7F",X"7F",X"00",X"00",X"41",X"41",X"7F",X"7F",X"41",X"41",
		X"00",X"20",X"60",X"40",X"40",X"40",X"7F",X"3F",X"00",X"7F",X"7F",X"18",X"3C",X"76",X"63",X"41",
		X"00",X"00",X"7F",X"7F",X"40",X"40",X"40",X"40",X"00",X"7F",X"7F",X"0E",X"1C",X"0E",X"7F",X"7F",
		X"00",X"7F",X"7F",X"0E",X"1C",X"38",X"7F",X"7F",X"00",X"3E",X"7F",X"41",X"41",X"41",X"7F",X"3E",
		X"00",X"7F",X"7F",X"11",X"11",X"11",X"1F",X"0E",X"00",X"3E",X"7F",X"41",X"51",X"71",X"3F",X"5E",
		X"00",X"7F",X"7F",X"11",X"31",X"79",X"6F",X"4E",X"00",X"26",X"6F",X"49",X"49",X"4B",X"7A",X"30",
		X"00",X"00",X"01",X"01",X"7F",X"7F",X"01",X"01",X"00",X"3F",X"7F",X"40",X"40",X"40",X"7F",X"3F",
		X"00",X"0F",X"1F",X"38",X"70",X"38",X"1F",X"0F",X"00",X"1F",X"7F",X"38",X"1C",X"38",X"7F",X"1F",
		X"00",X"63",X"77",X"3E",X"1C",X"3E",X"77",X"63",X"00",X"00",X"03",X"0F",X"78",X"78",X"0F",X"03",
		X"00",X"61",X"71",X"79",X"5D",X"4F",X"47",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"00",
		X"00",X"00",X"80",X"60",X"60",X"00",X"00",X"00",X"00",X"0C",X"02",X"A2",X"12",X"12",X"0C",X"00",
		X"00",X"00",X"BE",X"00",X"00",X"BE",X"00",X"00",X"7E",X"C3",X"99",X"A5",X"A5",X"81",X"C3",X"7E",
		X"00",X"FF",X"FF",X"C3",X"E7",X"7E",X"7E",X"FF",X"FF",X"DB",X"DB",X"DB",X"7E",X"FF",X"C3",X"C3",
		X"F7",X"76",X"7E",X"FF",X"C3",X"C3",X"FF",X"7E",X"7E",X"12",X"1E",X"00",X"7E",X"5A",X"5A",X"00",
		X"7E",X"12",X"1E",X"00",X"7E",X"12",X"1E",X"00",X"7E",X"5A",X"5A",X"00",X"7E",X"12",X"2E",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"C0",X"00",X"00",X"00",X"00",X"01",X"01",X"0F",X"01",X"01",X"00",X"0F",X"02",
		X"04",X"02",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"68",X"94",X"A8",X"40",X"00",
		X"00",X"00",X"10",X"0E",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"80",X"A0",X"80",X"00",X"00",X"20",X"00",X"50",X"00",X"00",X"20",X"80",X"80",X"80",X"00",
		X"00",X"03",X"1F",X"FF",X"FE",X"FC",X"F8",X"F9",X"F8",X"F9",X"FC",X"FE",X"FF",X"1F",X"03",X"00",
		X"00",X"00",X"00",X"10",X"08",X"00",X"22",X"00",X"08",X"00",X"20",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"02",X"15",X"2A",X"15",X"02",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"20",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"08",X"10",X"10",X"20",X"20",X"20",X"10",X"10",X"08",X"00",X"00",X"00",X"00",X"00",
		X"00",X"44",X"92",X"D6",X"92",X"D6",X"92",X"44",X"00",X"40",X"9A",X"82",X"8A",X"8A",X"9A",X"40",
		X"00",X"10",X"82",X"BA",X"82",X"BA",X"82",X"10",X"00",X"00",X"08",X"08",X"0A",X"08",X"08",X"00",
		X"00",X"00",X"00",X"2E",X"04",X"2E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"24",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"CC",X"E2",X"E0",X"20",X"20",X"20",X"60",X"64",X"E8",X"C0",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"24",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"08",X"00",X"02",X"80",X"E0",X"E0",X"E6",X"E0",X"00",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"24",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"40",X"68",X"68",X"28",X"24",X"20",X"20",X"60",X"E0",X"E0",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"4E",X"04",X"04",X"4E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"E0",X"EA",X"00",X"00",X"3A",X"30",X"20",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"4E",X"04",X"04",X"4E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"20",X"30",X"3A",X"00",X"00",X"EA",X"E0",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"20",X"30",X"30",X"00",X"00",X"00",X"E0",X"E0",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"E0",X"E0",X"00",X"00",X"00",X"30",X"30",X"20",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"4E",X"04",X"04",X"4E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"E0",X"EA",X"00",X"00",X"EA",X"E0",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"E0",X"E0",X"00",X"00",X"E0",X"E0",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"24",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"08",X"00",X"02",X"80",X"E0",X"E0",X"E6",X"E0",X"60",X"68",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"4E",X"04",X"04",X"4E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"E0",X"EA",X"00",X"00",X"2A",X"60",X"60",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"E0",X"E0",X"00",X"00",X"60",X"E0",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"4E",X"04",X"04",X"4E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"90",X"F0",X"F5",X"10",X"10",X"F5",X"F0",X"90",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"4E",X"04",X"04",X"4E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"90",X"F0",X"F5",X"10",X"10",X"F5",X"F0",X"90",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"40",X"20",X"00",X"00",X"20",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"90",X"F0",X"F5",X"10",X"10",X"F5",X"F0",X"90",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"06",X"0F",X"0F",X"0F",X"07",X"07",X"0F",X"0F",X"0F",X"06",X"00",X"00",X"00",
		X"00",X"00",X"FC",X"FE",X"C0",X"C0",X"80",X"80",X"80",X"C0",X"C0",X"FE",X"FC",X"00",X"00",X"00",
		X"00",X"00",X"00",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"00",X"00",X"00",
		X"00",X"00",X"30",X"60",X"C0",X"80",X"00",X"00",X"00",X"00",X"C0",X"E0",X"30",X"00",X"00",X"00",
		X"00",X"00",X"00",X"7F",X"FF",X"FD",X"FC",X"F8",X"F8",X"FC",X"FD",X"FF",X"7F",X"00",X"00",X"00",
		X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"00",
		X"00",X"00",X"0F",X"7F",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FF",X"7F",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0E",X"13",X"3F",X"FF",X"FF",X"FF",X"FE",X"FC",X"38",X"E0",X"00",X"00",X"00",
		X"80",X"80",X"80",X"9C",X"3E",X"2F",X"2F",X"2F",X"37",X"1B",X"0F",X"07",X"41",X"20",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"F8",X"FC",X"F2",X"FF",X"FF",X"FF",X"3F",X"1F",X"0E",
		X"00",X"08",X"10",X"10",X"20",X"00",X"03",X"0F",X"1F",X"1F",X"3F",X"3E",X"BF",X"BB",X"96",X"9C",
		X"00",X"00",X"00",X"00",X"F0",X"FC",X"FE",X"F3",X"FF",X"FF",X"F2",X"1C",X"00",X"00",X"00",X"00",
		X"00",X"10",X"20",X"40",X"03",X"0E",X"1B",X"37",X"3F",X"3F",X"1F",X"0E",X"80",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"1C",X"F2",X"FF",X"FF",X"F3",X"FE",X"FC",X"F0",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"80",X"0E",X"1B",X"2F",X"2F",X"3F",X"1F",X"0F",X"03",X"40",X"20",X"10",X"00",
		X"00",X"00",X"00",X"00",X"1C",X"FE",X"FF",X"FF",X"FF",X"FE",X"FC",X"F0",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"80",X"0E",X"1F",X"3F",X"3F",X"37",X"1B",X"0E",X"03",X"40",X"20",X"10",X"00",
		X"00",X"00",X"00",X"00",X"F0",X"DC",X"F6",X"FF",X"FF",X"FF",X"FE",X"1C",X"00",X"00",X"00",X"00",
		X"00",X"10",X"20",X"40",X"03",X"0F",X"1F",X"3F",X"3F",X"37",X"19",X"0E",X"80",X"80",X"80",X"80",
		X"00",X"E0",X"F0",X"F8",X"B8",X"A8",X"E8",X"F8",X"F0",X"F0",X"E0",X"E0",X"C0",X"80",X"60",X"80",
		X"00",X"00",X"01",X"83",X"83",X"87",X"47",X"1F",X"3F",X"7F",X"7F",X"7F",X"7D",X"33",X"1E",X"00",
		X"00",X"80",X"C0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",
		X"07",X"1F",X"3E",X"3D",X"7E",X"7D",X"FE",X"FC",X"FC",X"FC",X"FC",X"FE",X"FF",X"7E",X"7C",X"38",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"70",X"70",X"30",X"60",X"C0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"60",X"70",X"70",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"80",X"90",X"A4",X"00",X"80",X"90",X"A0",X"80",X"90",X"00",X"80",X"88",X"20",X"90",X"40",
		X"00",X"00",X"00",X"00",X"C0",X"E0",X"F8",X"D4",X"FC",X"E8",X"B8",X"70",X"00",X"00",X"00",X"00",
		X"40",X"40",X"80",X"80",X"0F",X"3D",X"7F",X"FE",X"FF",X"FF",X"7F",X"38",X"80",X"80",X"40",X"40",
		X"00",X"00",X"00",X"00",X"14",X"DE",X"F4",X"EF",X"B6",X"FC",X"E8",X"70",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"80",X"0C",X"1F",X"3C",X"3F",X"3F",X"1E",X"0F",X"03",X"80",X"80",X"80",X"80",
		X"E0",X"FC",X"7C",X"FE",X"BE",X"EF",X"FF",X"FF",X"B7",X"FF",X"FF",X"5E",X"FE",X"FC",X"F8",X"E0",
		X"21",X"47",X"4F",X"9F",X"9B",X"3E",X"37",X"3F",X"3D",X"BF",X"BB",X"9F",X"9F",X"8F",X"07",X"01",
		X"C0",X"E0",X"C0",X"C0",X"E0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"01",X"01",X"81",X"81",X"81",X"81",X"81",X"01",X"01",X"01",X"01",X"81",X"81",X"41",X"41",X"21",
		X"E0",X"F8",X"7C",X"FE",X"BE",X"EF",X"FF",X"FF",X"B7",X"FF",X"FF",X"5E",X"FE",X"FC",X"F8",X"E0",
		X"21",X"47",X"4F",X"9F",X"9B",X"3E",X"37",X"3F",X"3D",X"BF",X"BB",X"9F",X"9F",X"8F",X"07",X"01",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"E0",X"C0",X"C0",X"C0",X"C0",X"E0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"01",X"01",X"81",X"81",X"81",X"81",X"81",X"01",X"01",X"01",X"01",X"81",X"81",X"41",X"41",X"21",
		X"E0",X"F8",X"7C",X"FE",X"BE",X"EF",X"FF",X"FF",X"B7",X"FF",X"FF",X"5E",X"FE",X"FC",X"F8",X"E0",
		X"21",X"47",X"4F",X"9F",X"9B",X"3E",X"37",X"3F",X"3D",X"BF",X"BB",X"9F",X"9F",X"8F",X"07",X"01",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"01",X"01",X"81",X"81",X"81",X"81",X"81",X"01",X"01",X"01",X"01",X"81",X"81",X"41",X"41",X"21",
		X"00",X"C0",X"E0",X"F0",X"F0",X"F8",X"D8",X"F8",X"B8",X"F8",X"F8",X"F0",X"F0",X"E0",X"C0",X"00",
		X"87",X"9F",X"BB",X"7F",X"5F",X"FF",X"BF",X"FF",X"EF",X"FF",X"DF",X"7F",X"7F",X"BF",X"9F",X"87",
		X"00",X"00",X"00",X"80",X"80",X"C0",X"40",X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"00",X"00",X"00",
		X"58",X"BE",X"EF",X"7F",X"FF",X"FF",X"FF",X"FF",X"BE",X"FF",X"FF",X"FF",X"7F",X"FF",X"BE",X"58",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"60",X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F0",X"F0",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"80",X"88",X"00",X"A0",X"80",X"A0",X"00",X"88",X"80",X"A0",X"A0",X"88",X"00",X"A0",X"48",
		X"00",X"80",X"C0",X"F0",X"F0",X"E8",X"F8",X"78",X"F8",X"D8",X"F8",X"E0",X"F0",X"E0",X"80",X"00",
		X"20",X"47",X"9F",X"BF",X"3B",X"7F",X"7F",X"7F",X"7F",X"7B",X"7F",X"3F",X"BF",X"9E",X"47",X"20",
		X"00",X"E0",X"B8",X"F4",X"F8",X"FE",X"F4",X"FE",X"DA",X"FC",X"FE",X"FC",X"DC",X"F0",X"A0",X"00",
		X"80",X"80",X"87",X"8F",X"0F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"0F",X"8E",X"87",X"81",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"50",X"00",X"10",X"80",X"04",X"00",X"10",X"00",X"00",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"1C",X"3E",X"6E",X"6F",X"43",X"6F",X"3E",X"1C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"20",X"80",X"C0",X"68",X"E0",X"60",X"E4",X"C0",X"84",X"20",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"03",X"07",X"0D",X"0E",X"0D",X"0F",X"07",X"03",X"04",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"10",X"08",X"00",X"0C",X"08",X"06",X"06",X"0C",X"06",X"06",X"0C",X"0E",X"06",X"04",X"0E",
		X"0E",X"04",X"06",X"0E",X"0C",X"06",X"06",X"0C",X"06",X"06",X"08",X"0C",X"00",X"08",X"10",X"00",
		X"00",X"20",X"10",X"00",X"18",X"10",X"0C",X"0C",X"18",X"0C",X"0C",X"18",X"1C",X"0C",X"08",X"1C",
		X"1C",X"08",X"0C",X"1C",X"18",X"0C",X"0C",X"18",X"0C",X"0C",X"10",X"18",X"00",X"10",X"20",X"00",
		X"00",X"40",X"20",X"00",X"30",X"20",X"18",X"18",X"30",X"18",X"18",X"30",X"38",X"18",X"10",X"38",
		X"38",X"10",X"18",X"38",X"30",X"18",X"18",X"30",X"18",X"18",X"20",X"30",X"00",X"20",X"40",X"00",
		X"00",X"80",X"40",X"00",X"60",X"40",X"30",X"30",X"60",X"30",X"30",X"60",X"70",X"30",X"20",X"70",
		X"70",X"20",X"30",X"70",X"60",X"30",X"30",X"60",X"30",X"30",X"40",X"60",X"00",X"40",X"80",X"00",
		X"00",X"00",X"80",X"00",X"C0",X"80",X"60",X"60",X"C0",X"60",X"60",X"C0",X"E0",X"60",X"40",X"E0",
		X"E0",X"40",X"60",X"E0",X"C0",X"60",X"60",X"C0",X"60",X"60",X"80",X"C0",X"00",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"00",X"C0",X"C0",X"80",X"C0",X"C0",X"80",X"C0",X"C0",X"80",X"C0",
		X"C0",X"80",X"C0",X"C0",X"80",X"C0",X"C0",X"80",X"C0",X"C0",X"00",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"80",X"80",X"00",X"80",X"80",X"00",X"80",
		X"80",X"00",X"80",X"80",X"00",X"80",X"80",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"02",X"01",X"00",X"01",X"01",X"00",X"00",X"01",X"00",X"00",X"01",X"01",X"00",X"00",X"01",
		X"01",X"00",X"00",X"01",X"01",X"00",X"00",X"01",X"00",X"00",X"01",X"01",X"00",X"01",X"02",X"00",
		X"00",X"04",X"02",X"00",X"03",X"02",X"01",X"01",X"03",X"01",X"01",X"03",X"03",X"01",X"01",X"03",
		X"03",X"01",X"01",X"03",X"03",X"01",X"01",X"03",X"01",X"01",X"02",X"03",X"00",X"02",X"04",X"00",
		X"00",X"08",X"04",X"00",X"06",X"04",X"03",X"03",X"06",X"03",X"03",X"06",X"07",X"03",X"02",X"07",
		X"07",X"02",X"03",X"07",X"06",X"03",X"03",X"06",X"03",X"03",X"04",X"06",X"00",X"04",X"08",X"00",
		X"00",X"40",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"40",X"00",
		X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",
		X"00",X"01",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"01",X"00",
		X"00",X"02",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",
		X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"02",X"00",
		X"00",X"04",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",
		X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"04",X"00",
		X"00",X"08",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",
		X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"08",X"00",
		X"00",X"10",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",
		X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"10",X"00",
		X"00",X"20",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",
		X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"20",X"14",X"38",X"BA",X"7C",X"7E",X"FC",X"7C",X"7E",X"7C",X"FC",X"7C",X"FC",X"7E",
		X"7E",X"FC",X"7C",X"FC",X"7C",X"7E",X"7C",X"FC",X"7E",X"7C",X"BA",X"38",X"14",X"20",X"00",X"00",
		X"00",X"00",X"40",X"28",X"70",X"74",X"F8",X"FC",X"F8",X"F8",X"FC",X"F8",X"F8",X"F8",X"F8",X"FC",
		X"FC",X"F8",X"F8",X"F8",X"F8",X"FC",X"F8",X"F8",X"FC",X"F8",X"74",X"70",X"28",X"40",X"00",X"00",
		X"00",X"00",X"80",X"50",X"E0",X"E8",X"F0",X"F8",X"F0",X"F0",X"F8",X"F0",X"F0",X"F0",X"F0",X"F8",
		X"F8",X"F0",X"F0",X"F0",X"F0",X"F8",X"F0",X"F0",X"F8",X"F0",X"E8",X"E0",X"50",X"80",X"00",X"00",
		X"00",X"00",X"00",X"A0",X"C0",X"D0",X"E0",X"F0",X"E0",X"E0",X"F0",X"E0",X"E0",X"E0",X"E0",X"F0",
		X"F0",X"E0",X"E0",X"E0",X"E0",X"F0",X"E0",X"E0",X"F0",X"E0",X"D0",X"C0",X"A0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"40",X"80",X"A0",X"C0",X"E0",X"C0",X"C0",X"E0",X"C0",X"C0",X"C0",X"C0",X"E0",
		X"E0",X"C0",X"C0",X"C0",X"C0",X"E0",X"C0",X"C0",X"E0",X"C0",X"A0",X"80",X"40",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"00",X"40",X"80",X"C0",X"80",X"80",X"C0",X"80",X"80",X"80",X"80",X"C0",
		X"C0",X"80",X"80",X"80",X"80",X"C0",X"80",X"80",X"C0",X"80",X"40",X"00",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"80",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"80",
		X"80",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"80",X"00",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"01",X"01",X"03",X"01",X"01",X"01",X"03",X"01",X"03",X"01",
		X"01",X"03",X"01",X"03",X"01",X"01",X"01",X"03",X"01",X"01",X"02",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"01",X"05",X"03",X"03",X"07",X"03",X"03",X"03",X"07",X"03",X"07",X"03",
		X"03",X"07",X"03",X"07",X"03",X"03",X"03",X"07",X"03",X"03",X"05",X"01",X"00",X"01",X"00",X"00",
		X"00",X"00",X"02",X"01",X"03",X"0B",X"07",X"07",X"0F",X"07",X"07",X"07",X"0F",X"07",X"0F",X"07",
		X"07",X"0F",X"07",X"0F",X"07",X"07",X"07",X"0F",X"07",X"07",X"0B",X"03",X"01",X"02",X"00",X"00",
		X"00",X"00",X"04",X"02",X"07",X"17",X"0F",X"0F",X"1F",X"0F",X"0F",X"0F",X"1F",X"0F",X"1F",X"0F",
		X"0F",X"1F",X"0F",X"1F",X"0F",X"0F",X"0F",X"1F",X"0F",X"0F",X"17",X"07",X"02",X"04",X"00",X"00",
		X"00",X"00",X"08",X"05",X"0E",X"2E",X"1F",X"1F",X"3F",X"1F",X"1F",X"1F",X"3F",X"1F",X"3F",X"1F",
		X"1F",X"3F",X"1F",X"3F",X"1F",X"1F",X"1F",X"3F",X"1F",X"1F",X"2E",X"0E",X"05",X"08",X"00",X"00",
		X"00",X"00",X"10",X"0A",X"1C",X"5D",X"3E",X"3F",X"7E",X"3E",X"3F",X"3E",X"7E",X"3E",X"7E",X"3F",
		X"3F",X"7E",X"3E",X"7E",X"3E",X"3F",X"3E",X"7E",X"3F",X"3E",X"5D",X"1C",X"0A",X"10",X"00",X"00",
		X"00",X"00",X"FA",X"8A",X"90",X"B6",X"B6",X"F6",X"B6",X"F2",X"F6",X"F4",X"F6",X"F2",X"F4",X"F6",
		X"F2",X"F6",X"F6",X"F6",X"F2",X"F6",X"F4",X"F6",X"F2",X"F6",X"F4",X"B2",X"F8",X"C2",X"00",X"00",
		X"00",X"00",X"F4",X"14",X"20",X"6C",X"6C",X"EC",X"6C",X"E4",X"EC",X"E8",X"EC",X"E4",X"E8",X"EC",
		X"E4",X"EC",X"EC",X"EC",X"E4",X"EC",X"E8",X"EC",X"E4",X"EC",X"E8",X"64",X"F0",X"84",X"00",X"00",
		X"00",X"00",X"E8",X"28",X"40",X"D8",X"D8",X"D8",X"D8",X"C8",X"D8",X"D0",X"D8",X"C8",X"D0",X"D8",
		X"C8",X"D8",X"D8",X"D8",X"C8",X"D8",X"D0",X"D8",X"C8",X"D8",X"D0",X"C8",X"E0",X"08",X"00",X"00",
		X"00",X"00",X"D0",X"50",X"80",X"B0",X"B0",X"B0",X"B0",X"90",X"B0",X"A0",X"B0",X"90",X"A0",X"B0",
		X"90",X"B0",X"B0",X"B0",X"90",X"B0",X"A0",X"B0",X"90",X"B0",X"A0",X"90",X"C0",X"10",X"00",X"00",
		X"00",X"00",X"A0",X"A0",X"00",X"60",X"60",X"60",X"60",X"20",X"60",X"40",X"60",X"20",X"40",X"60",
		X"20",X"60",X"60",X"60",X"20",X"60",X"40",X"60",X"20",X"60",X"40",X"20",X"80",X"20",X"00",X"00",
		X"00",X"00",X"40",X"40",X"00",X"C0",X"C0",X"C0",X"C0",X"40",X"C0",X"80",X"C0",X"40",X"80",X"C0",
		X"40",X"C0",X"C0",X"C0",X"40",X"C0",X"80",X"C0",X"40",X"C0",X"80",X"40",X"00",X"40",X"00",X"00",
		X"00",X"00",X"80",X"80",X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"80",X"80",X"00",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"80",X"80",X"80",X"00",X"80",X"00",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",
		X"00",X"00",X"03",X"02",X"02",X"02",X"02",X"03",X"02",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"02",X"03",X"03",X"00",X"00",
		X"00",X"00",X"07",X"04",X"04",X"05",X"05",X"07",X"05",X"07",X"07",X"07",X"07",X"07",X"07",X"07",
		X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"05",X"07",X"06",X"00",X"00",
		X"00",X"00",X"0F",X"08",X"09",X"0B",X"0B",X"0F",X"0B",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0B",X"0F",X"0C",X"00",X"00",
		X"00",X"00",X"1F",X"11",X"12",X"16",X"16",X"1E",X"16",X"1E",X"1E",X"1E",X"1E",X"1E",X"1E",X"1E",
		X"1E",X"1E",X"1E",X"1E",X"1E",X"1E",X"1E",X"1E",X"1E",X"1E",X"1E",X"16",X"1F",X"18",X"00",X"00",
		X"00",X"00",X"3E",X"22",X"24",X"2D",X"2D",X"3D",X"2D",X"3C",X"3D",X"3D",X"3D",X"3C",X"3D",X"3D",
		X"3C",X"3D",X"3D",X"3D",X"3C",X"3D",X"3D",X"3D",X"3C",X"3D",X"3D",X"2C",X"3E",X"30",X"00",X"00",
		X"00",X"00",X"7D",X"45",X"48",X"5B",X"5B",X"7B",X"5B",X"79",X"7B",X"7A",X"7B",X"79",X"7A",X"7B",
		X"79",X"7B",X"7B",X"7B",X"79",X"7B",X"7A",X"7B",X"79",X"7B",X"7A",X"59",X"7C",X"61",X"00",X"00",
		X"D0",X"78",X"BC",X"FE",X"74",X"7A",X"FC",X"F8",X"7C",X"FA",X"FE",X"7C",X"3A",X"7C",X"F4",X"FE",
		X"FE",X"F4",X"7C",X"3A",X"7C",X"FE",X"FA",X"7C",X"F8",X"FC",X"7A",X"74",X"FE",X"BC",X"78",X"00",
		X"A0",X"F0",X"78",X"FC",X"E8",X"F4",X"F8",X"F0",X"F8",X"F4",X"FC",X"F8",X"74",X"F8",X"E8",X"FC",
		X"FC",X"E8",X"F8",X"74",X"F8",X"FC",X"F4",X"F8",X"F0",X"F8",X"F4",X"E8",X"FC",X"78",X"F0",X"00",
		X"40",X"E0",X"F0",X"F8",X"D0",X"E8",X"F0",X"E0",X"F0",X"E8",X"F8",X"F0",X"E8",X"F0",X"D0",X"F8",
		X"F8",X"D0",X"F0",X"E8",X"F0",X"F8",X"E8",X"F0",X"E0",X"F0",X"E8",X"D0",X"F8",X"F0",X"E0",X"00",
		X"80",X"C0",X"E0",X"F0",X"A0",X"D0",X"E0",X"C0",X"E0",X"D0",X"F0",X"E0",X"D0",X"E0",X"A0",X"F0",
		X"F0",X"A0",X"E0",X"D0",X"E0",X"F0",X"D0",X"E0",X"C0",X"E0",X"D0",X"A0",X"F0",X"E0",X"C0",X"00",
		X"00",X"80",X"C0",X"E0",X"40",X"A0",X"C0",X"80",X"C0",X"A0",X"E0",X"C0",X"A0",X"C0",X"40",X"E0",
		X"E0",X"40",X"C0",X"A0",X"C0",X"E0",X"A0",X"C0",X"80",X"C0",X"A0",X"40",X"E0",X"C0",X"80",X"00",
		X"00",X"00",X"80",X"C0",X"80",X"40",X"80",X"00",X"80",X"40",X"C0",X"80",X"40",X"80",X"80",X"C0",
		X"C0",X"80",X"80",X"40",X"80",X"C0",X"40",X"80",X"00",X"80",X"40",X"80",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"80",X"00",X"80",X"00",X"00",X"00",X"80",X"80",X"00",X"80",X"00",X"00",X"80",
		X"80",X"00",X"00",X"80",X"00",X"80",X"80",X"00",X"00",X"00",X"80",X"00",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"01",X"01",X"00",X"00",X"01",X"01",X"00",X"01",X"01",X"00",X"00",X"00",X"01",X"01",
		X"01",X"01",X"00",X"00",X"00",X"01",X"01",X"00",X"01",X"01",X"00",X"00",X"01",X"01",X"00",X"00",
		X"03",X"01",X"02",X"03",X"01",X"01",X"03",X"03",X"01",X"03",X"03",X"01",X"00",X"01",X"03",X"03",
		X"03",X"03",X"01",X"00",X"01",X"03",X"03",X"01",X"03",X"03",X"01",X"01",X"03",X"02",X"01",X"00",
		X"06",X"03",X"05",X"07",X"03",X"03",X"07",X"07",X"03",X"07",X"07",X"03",X"01",X"03",X"07",X"07",
		X"07",X"07",X"03",X"01",X"03",X"07",X"07",X"03",X"07",X"07",X"03",X"03",X"07",X"05",X"03",X"00",
		X"0D",X"07",X"0B",X"0F",X"07",X"07",X"0F",X"0F",X"07",X"0F",X"0F",X"07",X"03",X"07",X"0F",X"0F",
		X"0F",X"0F",X"07",X"03",X"07",X"0F",X"0F",X"07",X"0F",X"0F",X"07",X"07",X"0F",X"0B",X"07",X"00",
		X"1A",X"0F",X"17",X"1F",X"0E",X"0F",X"1F",X"1F",X"0F",X"1F",X"1F",X"0F",X"07",X"0F",X"1E",X"1F",
		X"1F",X"1E",X"0F",X"07",X"0F",X"1F",X"1F",X"0F",X"1F",X"1F",X"0F",X"0E",X"1F",X"17",X"0F",X"00",
		X"34",X"1E",X"2F",X"3F",X"1D",X"1E",X"3F",X"3E",X"1F",X"3E",X"3F",X"1F",X"0E",X"1F",X"3D",X"3F",
		X"3F",X"3D",X"1F",X"0E",X"1F",X"3F",X"3E",X"1F",X"3E",X"3F",X"1E",X"1D",X"3F",X"2F",X"1E",X"00",
		X"68",X"3C",X"5E",X"7F",X"3A",X"3D",X"7E",X"7C",X"3E",X"7D",X"7F",X"3E",X"1D",X"3E",X"7A",X"7F",
		X"7F",X"7A",X"3E",X"1D",X"3E",X"7F",X"7D",X"3E",X"7C",X"7E",X"3D",X"3A",X"7F",X"5E",X"3C",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
