library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ttag_bg_bits_2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ttag_bg_bits_2 is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"50",X"15",X"01",X"50",X"15",X"01",X"50",X"15",X"50",X"54",X"05",X"40",X"54",X"05",X"40",X"54",
		X"51",X"50",X"15",X"01",X"50",X"15",X"01",X"50",X"55",X"40",X"54",X"05",X"40",X"54",X"05",X"40",
		X"55",X"01",X"50",X"15",X"01",X"50",X"15",X"00",X"54",X"05",X"40",X"54",X"05",X"40",X"54",X"00",
		X"50",X"15",X"01",X"50",X"15",X"01",X"50",X"00",X"50",X"54",X"05",X"40",X"54",X"05",X"40",X"00",
		X"51",X"50",X"15",X"01",X"50",X"15",X"00",X"00",X"55",X"40",X"54",X"05",X"40",X"54",X"00",X"00",
		X"55",X"01",X"50",X"15",X"01",X"50",X"00",X"00",X"54",X"05",X"40",X"54",X"05",X"40",X"00",X"00",
		X"50",X"15",X"01",X"50",X"15",X"00",X"00",X"00",X"50",X"54",X"05",X"40",X"54",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"01",X"55",X"01",X"50",X"15",X"01",X"50",X"15",X"01",X"54",X"05",X"40",X"54",X"05",X"40",X"54",
		X"00",X"54",X"15",X"01",X"50",X"15",X"01",X"50",X"00",X"14",X"54",X"05",X"40",X"54",X"05",X"40",
		X"00",X"15",X"50",X"15",X"01",X"50",X"15",X"00",X"00",X"05",X"40",X"54",X"05",X"40",X"54",X"00",
		X"00",X"01",X"41",X"50",X"15",X"01",X"50",X"00",X"00",X"01",X"55",X"40",X"54",X"05",X"40",X"00",
		X"00",X"00",X"55",X"01",X"50",X"15",X"00",X"00",X"00",X"00",X"14",X"05",X"40",X"54",X"00",X"00",
		X"00",X"00",X"15",X"15",X"01",X"50",X"00",X"00",X"00",X"00",X"05",X"54",X"05",X"40",X"00",X"00",
		X"00",X"00",X"01",X"50",X"15",X"00",X"00",X"00",X"00",X"00",X"01",X"50",X"54",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"55",X"40",X"54",X"05",X"40",X"54",X"05",X"00",X"55",X"01",X"50",X"15",X"01",X"50",X"15",
		X"00",X"15",X"05",X"40",X"54",X"05",X"40",X"55",X"00",X"05",X"15",X"01",X"50",X"15",X"01",X"55",
		X"00",X"05",X"54",X"05",X"40",X"54",X"05",X"45",X"00",X"01",X"50",X"15",X"01",X"50",X"15",X"05",
		X"00",X"00",X"50",X"54",X"05",X"40",X"54",X"05",X"00",X"00",X"55",X"50",X"15",X"01",X"50",X"15",
		X"00",X"00",X"15",X"40",X"54",X"05",X"40",X"55",X"00",X"00",X"05",X"01",X"50",X"15",X"01",X"55",
		X"00",X"00",X"05",X"45",X"40",X"54",X"05",X"45",X"00",X"00",X"01",X"55",X"01",X"50",X"15",X"05",
		X"00",X"00",X"00",X"54",X"05",X"40",X"54",X"05",X"00",X"00",X"00",X"54",X"15",X"01",X"50",X"15",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"28",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"A0",X"20",X"00",X"00",X"00",
		X"00",X"00",X"00",X"20",X"28",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"2A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"54",X"05",X"40",X"54",X"05",X"40",X"55",X"00",X"55",X"01",X"50",X"15",X"01",X"50",X"15",X"00",
		X"55",X"40",X"54",X"05",X"40",X"54",X"54",X"00",X"51",X"50",X"15",X"01",X"50",X"15",X"50",X"00",
		X"50",X"54",X"05",X"40",X"54",X"05",X"50",X"00",X"50",X"15",X"01",X"50",X"15",X"05",X"40",X"00",
		X"54",X"05",X"40",X"54",X"05",X"45",X"00",X"00",X"55",X"01",X"50",X"15",X"01",X"55",X"00",X"00",
		X"55",X"40",X"54",X"05",X"40",X"54",X"00",X"00",X"51",X"50",X"15",X"01",X"50",X"50",X"00",X"00",
		X"50",X"54",X"05",X"40",X"54",X"50",X"00",X"00",X"50",X"15",X"01",X"50",X"15",X"40",X"00",X"00",
		X"54",X"05",X"40",X"54",X"05",X"00",X"00",X"00",X"55",X"01",X"50",X"15",X"15",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"54",X"05",X"40",X"54",X"05",X"40",X"55",X"00",X"15",X"01",X"50",X"15",X"01",X"50",X"15",X"00",
		X"05",X"40",X"54",X"05",X"40",X"54",X"54",X"00",X"01",X"50",X"15",X"01",X"50",X"15",X"50",X"00",
		X"00",X"54",X"05",X"40",X"54",X"05",X"50",X"00",X"00",X"15",X"01",X"50",X"15",X"05",X"40",X"00",
		X"00",X"05",X"40",X"54",X"05",X"45",X"00",X"00",X"00",X"01",X"50",X"15",X"01",X"55",X"00",X"00",
		X"00",X"00",X"54",X"05",X"40",X"54",X"00",X"00",X"00",X"00",X"15",X"01",X"50",X"50",X"00",X"00",
		X"00",X"00",X"05",X"40",X"55",X"50",X"00",X"00",X"00",X"00",X"01",X"50",X"15",X"40",X"00",X"00",
		X"00",X"00",X"00",X"54",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"15",X"15",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"54",X"05",X"40",X"54",X"05",X"40",X"54",X"05",X"15",X"01",X"50",X"15",X"01",X"50",X"15",X"05",
		X"05",X"40",X"54",X"05",X"40",X"54",X"05",X"45",X"01",X"50",X"15",X"01",X"50",X"15",X"01",X"55",
		X"00",X"54",X"05",X"40",X"54",X"05",X"40",X"55",X"00",X"15",X"01",X"50",X"15",X"01",X"50",X"15",
		X"00",X"05",X"40",X"54",X"05",X"40",X"54",X"05",X"00",X"01",X"50",X"15",X"01",X"50",X"15",X"05",
		X"00",X"00",X"54",X"05",X"40",X"54",X"05",X"45",X"00",X"00",X"15",X"01",X"50",X"15",X"01",X"55",
		X"00",X"00",X"05",X"40",X"54",X"05",X"40",X"55",X"00",X"00",X"01",X"50",X"15",X"01",X"50",X"15",
		X"00",X"00",X"00",X"54",X"05",X"40",X"54",X"05",X"00",X"00",X"00",X"15",X"01",X"50",X"15",X"05",
		X"2A",X"AA",X"CF",X"3C",X"F3",X"CF",X"AA",X"A8",X"20",X"96",X"F3",X"CF",X"3C",X"F3",X"82",X"58",
		X"20",X"AA",X"FC",X"F3",X"CF",X"3F",X"AA",X"58",X"20",X"96",X"CF",X"3C",X"F3",X"CF",X"82",X"58",
		X"2A",X"96",X"F3",X"CF",X"3C",X"F3",X"82",X"A8",X"20",X"96",X"33",X"33",X"33",X"33",X"82",X"08",
		X"A0",X"AA",X"CC",X"CC",X"CC",X"CC",X"AA",X"0A",X"08",X"82",X"33",X"33",X"33",X"33",X"82",X"08",
		X"02",X"82",X"CC",X"CC",X"CC",X"CC",X"82",X"20",X"AA",X"82",X"33",X"33",X"33",X"33",X"82",X"AA",
		X"25",X"62",X"CC",X"CC",X"CC",X"CC",X"82",X"58",X"25",X"5A",X"33",X"33",X"33",X"33",X"89",X"58",
		X"AA",X"AA",X"CC",X"0C",X"CC",X"00",X"AA",X"AA",X"02",X"56",X"33",X"03",X"03",X"33",X"80",X"95",
		X"02",X"56",X"C0",X"C0",X"0C",X"0C",X"80",X"95",X"AA",X"AA",X"00",X"00",X"00",X"00",X"AA",X"AA",
		X"51",X"50",X"15",X"01",X"50",X"00",X"00",X"00",X"55",X"40",X"54",X"05",X"40",X"00",X"00",X"00",
		X"55",X"01",X"50",X"15",X"00",X"00",X"00",X"00",X"54",X"05",X"40",X"54",X"00",X"00",X"00",X"00",
		X"50",X"15",X"01",X"50",X"00",X"00",X"00",X"00",X"50",X"54",X"05",X"40",X"00",X"00",X"00",X"00",
		X"51",X"50",X"15",X"00",X"00",X"00",X"00",X"00",X"55",X"40",X"54",X"00",X"00",X"00",X"00",X"00",
		X"55",X"01",X"50",X"00",X"00",X"00",X"00",X"00",X"54",X"05",X"40",X"00",X"00",X"00",X"00",X"00",
		X"50",X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"54",X"00",X"00",X"00",X"00",X"00",X"00",
		X"51",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"55",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"15",X"40",X"00",X"00",X"00",
		X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"40",X"00",X"00",X"00",X"00",
		X"00",X"00",X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"14",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"15",X"54",X"05",X"40",X"55",X"00",X"00",X"00",X"05",X"50",X"15",X"01",X"55",
		X"00",X"00",X"00",X"05",X"40",X"54",X"05",X"45",X"00",X"00",X"00",X"15",X"01",X"50",X"15",X"05",
		X"00",X"00",X"00",X"54",X"05",X"40",X"54",X"05",X"00",X"00",X"01",X"50",X"15",X"01",X"50",X"15",
		X"00",X"00",X"05",X"40",X"54",X"05",X"40",X"55",X"00",X"00",X"15",X"01",X"50",X"15",X"01",X"55",
		X"00",X"00",X"54",X"05",X"40",X"54",X"05",X"45",X"00",X"01",X"50",X"15",X"01",X"50",X"15",X"05",
		X"00",X"05",X"40",X"54",X"05",X"40",X"54",X"05",X"00",X"15",X"01",X"50",X"15",X"01",X"50",X"15",
		X"00",X"54",X"05",X"40",X"54",X"05",X"40",X"55",X"01",X"50",X"15",X"01",X"50",X"15",X"01",X"55",
		X"05",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"15",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"A8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"A8",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"A8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"A8",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"A8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"A8",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"A8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"A8",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"A8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"A8",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"A8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"A8",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"A8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"40",X"54",X"05",X"54",X"00",X"00",X"00",X"51",X"50",X"15",X"01",X"50",X"00",X"00",X"00",
		X"50",X"54",X"05",X"40",X"54",X"00",X"00",X"00",X"50",X"15",X"01",X"50",X"15",X"00",X"00",X"00",
		X"54",X"05",X"40",X"54",X"05",X"40",X"00",X"00",X"55",X"01",X"50",X"15",X"01",X"50",X"00",X"00",
		X"55",X"40",X"54",X"05",X"40",X"54",X"00",X"00",X"51",X"50",X"15",X"01",X"50",X"15",X"00",X"00",
		X"50",X"54",X"05",X"40",X"54",X"05",X"40",X"00",X"50",X"15",X"01",X"50",X"15",X"01",X"50",X"00",
		X"54",X"05",X"40",X"54",X"05",X"40",X"54",X"00",X"55",X"01",X"50",X"15",X"01",X"50",X"15",X"00",
		X"55",X"40",X"54",X"05",X"40",X"54",X"05",X"40",X"51",X"50",X"15",X"01",X"50",X"15",X"01",X"50",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"54",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"05",X"54",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"50",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"15",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"05",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"50",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"15",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"05",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"50",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"15",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"50",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"15",
		X"00",X"00",X"00",X"05",X"40",X"54",X"05",X"45",X"00",X"00",X"00",X"01",X"50",X"15",X"01",X"55",
		X"00",X"00",X"00",X"00",X"54",X"05",X"40",X"55",X"00",X"00",X"00",X"00",X"15",X"01",X"50",X"15",
		X"00",X"00",X"00",X"00",X"05",X"40",X"54",X"05",X"00",X"00",X"00",X"00",X"01",X"50",X"15",X"05",
		X"00",X"00",X"00",X"00",X"00",X"54",X"05",X"45",X"00",X"00",X"00",X"00",X"00",X"15",X"01",X"55",
		X"00",X"00",X"00",X"00",X"00",X"05",X"40",X"55",X"00",X"00",X"00",X"00",X"00",X"01",X"50",X"15",
		X"00",X"00",X"00",X"00",X"00",X"00",X"54",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"15",X"05",
		X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"45",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"15",
		X"0C",X"CC",X"CF",X"FC",X"FF",X"FF",X"FF",X"FF",X"00",X"33",X"33",X"CF",X"FF",X"FF",X"FF",X"FF",
		X"0C",X"CC",X"CC",X"F3",X"FF",X"FF",X"FF",X"FF",X"33",X"33",X"33",X"3C",X"FF",X"FF",X"FF",X"FF",
		X"0C",X"CC",X"CF",X"CF",X"FF",X"FF",X"FF",X"FF",X"00",X"33",X"30",X"F3",X"FF",X"FF",X"FF",X"FF",
		X"00",X"CC",X"CF",X"3C",X"FF",X"FF",X"FF",X"FF",X"33",X"30",X"33",X"CF",X"FF",X"FF",X"FF",X"FF",
		X"0C",X"CC",X"CC",X"F3",X"FF",X"FF",X"FF",X"FF",X"30",X"33",X"33",X"3C",X"FF",X"FF",X"FF",X"FF",
		X"0C",X"CC",X"0F",X"CF",X"FF",X"FF",X"FF",X"FF",X"30",X"33",X"30",X"F3",X"FF",X"FF",X"FF",X"FF",
		X"00",X"0C",X"CC",X"3C",X"FF",X"FF",X"FF",X"FF",X"03",X"33",X"33",X"CF",X"FF",X"FF",X"FF",X"FF",
		X"0C",X"CC",X"CC",X"F3",X"FF",X"FF",X"FF",X"FF",X"33",X"33",X"33",X"3C",X"FF",X"FF",X"FF",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"50",X"15",X"01",X"50",X"15",X"01",X"50",X"15",X"50",X"54",X"05",X"40",X"54",X"05",X"40",X"54",
		X"51",X"50",X"15",X"01",X"50",X"15",X"01",X"50",X"55",X"40",X"54",X"05",X"40",X"54",X"05",X"40",
		X"55",X"01",X"50",X"15",X"01",X"50",X"15",X"00",X"54",X"05",X"40",X"54",X"05",X"40",X"54",X"00",
		X"50",X"15",X"01",X"50",X"15",X"01",X"50",X"00",X"50",X"54",X"05",X"40",X"54",X"05",X"40",X"00",
		X"51",X"50",X"15",X"01",X"50",X"15",X"00",X"00",X"55",X"40",X"54",X"05",X"40",X"54",X"00",X"00",
		X"55",X"01",X"50",X"15",X"01",X"50",X"00",X"00",X"54",X"05",X"40",X"54",X"05",X"40",X"00",X"00",
		X"50",X"15",X"01",X"50",X"15",X"00",X"00",X"00",X"50",X"54",X"05",X"40",X"54",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"55",X"01",X"50",X"15",X"01",X"50",X"15",X"00",X"54",X"05",X"40",X"54",X"05",X"40",X"54",
		X"00",X"15",X"15",X"01",X"50",X"15",X"01",X"50",X"00",X"05",X"54",X"05",X"40",X"54",X"05",X"40",
		X"00",X"05",X"50",X"15",X"01",X"50",X"15",X"00",X"00",X"01",X"50",X"54",X"05",X"40",X"54",X"00",
		X"00",X"00",X"51",X"50",X"15",X"01",X"50",X"00",X"00",X"00",X"55",X"40",X"54",X"05",X"40",X"00",
		X"00",X"00",X"15",X"01",X"50",X"15",X"00",X"00",X"00",X"00",X"05",X"05",X"40",X"54",X"00",X"00",
		X"00",X"00",X"05",X"55",X"01",X"50",X"00",X"00",X"00",X"00",X"01",X"54",X"05",X"40",X"00",X"00",
		X"00",X"00",X"00",X"50",X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"54",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"55",X"01",X"50",X"15",X"01",X"50",X"15",X"00",X"54",X"05",X"40",X"54",X"05",X"40",X"55",
		X"00",X"15",X"15",X"01",X"50",X"15",X"01",X"55",X"00",X"05",X"54",X"05",X"40",X"54",X"05",X"45",
		X"00",X"05",X"50",X"15",X"01",X"50",X"15",X"05",X"00",X"01",X"50",X"54",X"05",X"40",X"54",X"05",
		X"00",X"00",X"51",X"50",X"15",X"01",X"50",X"15",X"00",X"00",X"55",X"40",X"54",X"05",X"40",X"55",
		X"00",X"00",X"15",X"01",X"50",X"15",X"01",X"55",X"00",X"00",X"05",X"05",X"40",X"54",X"05",X"45",
		X"00",X"00",X"05",X"55",X"01",X"50",X"15",X"05",X"00",X"00",X"01",X"54",X"05",X"40",X"54",X"05",
		X"00",X"00",X"00",X"50",X"15",X"01",X"50",X"15",X"00",X"00",X"00",X"54",X"54",X"05",X"40",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"A8",X"A0",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A8",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"80",X"00",X"00",X"00",X"00",X"00",
		X"02",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",
		X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"01",X"50",X"15",X"01",X"50",X"15",X"00",X"55",X"40",X"54",X"05",X"40",X"54",X"14",X"00",
		X"51",X"50",X"15",X"01",X"50",X"15",X"54",X"00",X"50",X"54",X"05",X"40",X"54",X"05",X"50",X"00",
		X"50",X"15",X"01",X"50",X"15",X"01",X"40",X"00",X"54",X"05",X"40",X"54",X"05",X"45",X"40",X"00",
		X"55",X"01",X"50",X"15",X"01",X"55",X"00",X"00",X"55",X"40",X"54",X"05",X"40",X"54",X"00",X"00",
		X"51",X"50",X"15",X"01",X"50",X"54",X"00",X"00",X"50",X"54",X"05",X"40",X"55",X"50",X"00",X"00",
		X"50",X"15",X"01",X"50",X"15",X"40",X"00",X"00",X"54",X"05",X"40",X"54",X"05",X"40",X"00",X"00",
		X"55",X"01",X"50",X"15",X"15",X"00",X"00",X"00",X"55",X"40",X"54",X"05",X"54",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"54",X"05",X"40",X"54",X"05",X"40",X"15",X"00",X"15",X"01",X"50",X"15",X"01",X"50",X"14",X"00",
		X"05",X"40",X"54",X"05",X"40",X"54",X"54",X"00",X"01",X"50",X"15",X"01",X"50",X"15",X"50",X"00",
		X"00",X"54",X"05",X"40",X"54",X"05",X"40",X"00",X"00",X"15",X"01",X"50",X"15",X"15",X"40",X"00",
		X"00",X"05",X"40",X"54",X"05",X"55",X"00",X"00",X"00",X"01",X"50",X"15",X"01",X"54",X"00",X"00",
		X"00",X"00",X"54",X"05",X"40",X"54",X"00",X"00",X"00",X"00",X"15",X"01",X"51",X"50",X"00",X"00",
		X"00",X"00",X"05",X"40",X"55",X"40",X"00",X"00",X"00",X"00",X"01",X"50",X"15",X"40",X"00",X"00",
		X"00",X"00",X"00",X"54",X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"15",X"14",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"54",X"05",X"40",X"54",X"05",X"40",X"54",X"05",X"15",X"01",X"50",X"15",X"01",X"50",X"15",X"05",
		X"05",X"40",X"54",X"05",X"40",X"54",X"05",X"45",X"01",X"50",X"15",X"01",X"50",X"15",X"01",X"55",
		X"00",X"54",X"05",X"40",X"54",X"05",X"40",X"55",X"00",X"15",X"01",X"50",X"15",X"01",X"50",X"15",
		X"00",X"05",X"40",X"54",X"05",X"40",X"54",X"05",X"00",X"01",X"50",X"15",X"01",X"50",X"15",X"05",
		X"00",X"00",X"54",X"05",X"40",X"54",X"05",X"45",X"00",X"00",X"15",X"01",X"50",X"15",X"01",X"55",
		X"00",X"00",X"05",X"40",X"54",X"05",X"40",X"55",X"00",X"00",X"01",X"50",X"15",X"01",X"50",X"15",
		X"00",X"00",X"00",X"54",X"05",X"40",X"54",X"05",X"00",X"00",X"00",X"15",X"01",X"50",X"15",X"05",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"30",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"CC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"30",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"CC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"CC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"30",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"CC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"0C",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"30",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"C0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"30",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"CC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"CC",
		X"51",X"50",X"15",X"01",X"50",X"00",X"00",X"00",X"55",X"40",X"54",X"05",X"40",X"00",X"00",X"00",
		X"55",X"01",X"50",X"15",X"00",X"00",X"00",X"00",X"54",X"05",X"40",X"54",X"00",X"00",X"00",X"00",
		X"50",X"15",X"01",X"50",X"00",X"00",X"00",X"00",X"50",X"54",X"05",X"40",X"00",X"00",X"00",X"00",
		X"51",X"50",X"15",X"00",X"00",X"00",X"00",X"00",X"55",X"40",X"54",X"00",X"00",X"00",X"00",X"00",
		X"55",X"01",X"50",X"00",X"00",X"00",X"00",X"00",X"54",X"05",X"40",X"00",X"00",X"00",X"00",X"00",
		X"50",X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"54",X"00",X"00",X"00",X"00",X"00",X"00",
		X"51",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"15",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"40",X"00",X"00",X"00",
		X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"40",X"00",X"00",X"00",X"00",
		X"00",X"00",X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"15",X"50",X"15",X"01",X"55",X"00",X"00",X"00",X"05",X"40",X"54",X"05",X"45",
		X"00",X"00",X"00",X"15",X"01",X"50",X"15",X"05",X"00",X"00",X"00",X"54",X"05",X"40",X"54",X"05",
		X"00",X"00",X"01",X"50",X"15",X"01",X"50",X"15",X"00",X"00",X"05",X"40",X"54",X"05",X"40",X"55",
		X"00",X"00",X"15",X"01",X"50",X"15",X"01",X"55",X"00",X"00",X"54",X"05",X"40",X"54",X"05",X"45",
		X"00",X"01",X"50",X"15",X"01",X"50",X"15",X"05",X"00",X"05",X"40",X"54",X"05",X"40",X"54",X"05",
		X"00",X"15",X"01",X"50",X"15",X"01",X"50",X"15",X"00",X"54",X"05",X"40",X"54",X"05",X"40",X"55",
		X"01",X"50",X"15",X"01",X"50",X"15",X"01",X"55",X"05",X"40",X"54",X"05",X"40",X"54",X"05",X"45",
		X"15",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"AA",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0A",X"AA",X"80",X"00",X"00",X"00",X"00",X"00",X"2A",X"AA",X"A0",X"00",X"00",
		X"00",X"00",X"00",X"2A",X"AA",X"A0",X"00",X"00",X"00",X"00",X"00",X"2A",X"AA",X"A0",X"00",X"00",
		X"00",X"00",X"00",X"2A",X"AA",X"A0",X"00",X"00",X"00",X"00",X"00",X"2A",X"AA",X"A0",X"00",X"00",
		X"00",X"00",X"00",X"2A",X"AA",X"A0",X"00",X"00",X"00",X"00",X"00",X"2A",X"AA",X"A0",X"00",X"00",
		X"00",X"00",X"00",X"0A",X"AA",X"80",X"00",X"00",X"00",X"00",X"00",X"02",X"AA",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"51",X"50",X"15",X"01",X"54",X"00",X"00",X"00",X"50",X"54",X"05",X"40",X"54",X"00",X"00",X"00",
		X"50",X"15",X"01",X"50",X"15",X"00",X"00",X"00",X"54",X"05",X"40",X"54",X"05",X"40",X"00",X"00",
		X"55",X"01",X"50",X"15",X"01",X"50",X"00",X"00",X"55",X"40",X"54",X"05",X"40",X"54",X"00",X"00",
		X"51",X"50",X"15",X"01",X"50",X"15",X"00",X"00",X"50",X"54",X"05",X"40",X"54",X"05",X"40",X"00",
		X"50",X"15",X"01",X"50",X"15",X"01",X"50",X"00",X"54",X"05",X"40",X"54",X"05",X"40",X"54",X"00",
		X"55",X"01",X"50",X"15",X"01",X"50",X"15",X"00",X"55",X"40",X"54",X"05",X"40",X"54",X"05",X"40",
		X"51",X"50",X"15",X"01",X"50",X"15",X"01",X"50",X"50",X"54",X"05",X"40",X"54",X"05",X"40",X"54",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"05",X"54",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"50",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"15",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"05",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"50",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"15",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"05",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"50",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"15",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"50",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"15",
		X"00",X"00",X"00",X"05",X"40",X"54",X"05",X"45",X"00",X"00",X"00",X"01",X"50",X"15",X"01",X"55",
		X"00",X"00",X"00",X"00",X"54",X"05",X"40",X"55",X"00",X"00",X"00",X"00",X"15",X"01",X"50",X"15",
		X"00",X"00",X"00",X"00",X"05",X"40",X"54",X"05",X"00",X"00",X"00",X"00",X"01",X"50",X"15",X"05",
		X"00",X"00",X"00",X"00",X"00",X"54",X"05",X"45",X"00",X"00",X"00",X"00",X"00",X"15",X"01",X"55",
		X"00",X"00",X"00",X"00",X"00",X"05",X"40",X"55",X"00",X"00",X"00",X"00",X"00",X"01",X"50",X"15",
		X"00",X"00",X"00",X"00",X"00",X"00",X"54",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"15",X"05",
		X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"45",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"15",
		X"82",X"08",X"20",X"00",X"00",X"00",X"00",X"00",X"AA",X"0A",X"A0",X"00",X"00",X"00",X"00",X"00",
		X"96",X"08",X"20",X"00",X"00",X"00",X"00",X"00",X"96",X"A8",X"20",X"00",X"00",X"00",X"00",X"00",
		X"96",X"08",X"20",X"00",X"00",X"00",X"00",X"00",X"96",X"08",X"20",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"95",X"60",X"25",X"60",X"20",X"25",X"60",X"20",
		X"95",X"60",X"25",X"60",X"20",X"25",X"60",X"20",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"82",X"02",X"02",X"02",X"56",X"02",X"02",X"02",X"82",X"02",X"02",X"02",X"56",X"02",X"02",X"02",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"80",X"25",X"60",X"20",X"20",X"20",X"25",X"60",
		X"80",X"25",X"60",X"20",X"20",X"20",X"25",X"60",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"20",X"00",X"00",X"00",X"0F",
		X"00",X"08",X"00",X"20",X"00",X"00",X"03",X"FF",X"00",X"08",X"00",X"20",X"00",X"00",X"FF",X"FF",
		X"00",X"02",X"00",X"80",X"00",X"3F",X"FF",X"FF",X"00",X"00",X"AA",X"00",X"0F",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"03",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"D5",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"FD",X"00",X"00",X"00",
		X"00",X"00",X"01",X"03",X"FD",X"00",X"00",X"00",X"00",X"00",X"0D",X"03",X"FD",X"03",X"C1",X"00",
		X"00",X"03",X"FD",X"03",X"FD",X"03",X"FD",X"00",X"00",X"FF",X"FD",X"03",X"FD",X"03",X"FD",X"00",
		X"3F",X"FF",X"FD",X"03",X"FD",X"03",X"FD",X"00",X"FF",X"FF",X"FD",X"03",X"FD",X"03",X"FD",X"00",
		X"FF",X"FF",X"FD",X"03",X"FD",X"03",X"FD",X"00",X"FF",X"FF",X"FD",X"03",X"FD",X"03",X"FD",X"00",
		X"FF",X"FF",X"FD",X"03",X"FD",X"03",X"FD",X"00",X"FD",X"5F",X"FD",X"03",X"FD",X"03",X"FD",X"00",
		X"54",X"03",X"FD",X"03",X"FD",X"03",X"FD",X"00",X"00",X"03",X"FD",X"03",X"FD",X"03",X"FD",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"3F",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"FF",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"2A",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"2A",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",
		X"2A",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"2A",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",
		X"2A",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"2A",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",
		X"2A",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"2A",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",
		X"2A",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"2A",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",
		X"2A",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"2A",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",
		X"2A",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"54",X"05",X"40",X"54",X"05",X"40",X"54",X"05",X"15",X"01",X"50",X"15",X"01",X"50",X"15",X"05",
		X"05",X"40",X"54",X"05",X"40",X"54",X"05",X"45",X"01",X"50",X"15",X"01",X"50",X"15",X"01",X"55",
		X"00",X"54",X"05",X"40",X"54",X"05",X"40",X"55",X"00",X"15",X"01",X"50",X"15",X"01",X"50",X"15",
		X"00",X"05",X"40",X"54",X"05",X"40",X"54",X"05",X"00",X"01",X"50",X"15",X"01",X"50",X"15",X"05",
		X"00",X"00",X"54",X"05",X"40",X"54",X"05",X"45",X"00",X"00",X"15",X"01",X"50",X"15",X"01",X"55",
		X"00",X"00",X"05",X"40",X"54",X"05",X"40",X"55",X"00",X"00",X"01",X"50",X"15",X"01",X"50",X"15",
		X"00",X"00",X"00",X"54",X"05",X"40",X"54",X"05",X"00",X"00",X"00",X"15",X"01",X"50",X"15",X"05",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"50",X"15",X"01",X"50",X"15",X"01",X"50",X"15",X"50",X"54",X"05",X"40",X"54",X"05",X"40",X"54",
		X"51",X"50",X"15",X"01",X"50",X"15",X"01",X"50",X"55",X"40",X"54",X"05",X"40",X"54",X"05",X"40",
		X"55",X"01",X"50",X"15",X"01",X"50",X"15",X"00",X"54",X"05",X"40",X"54",X"05",X"40",X"54",X"00",
		X"50",X"15",X"01",X"50",X"15",X"01",X"50",X"00",X"50",X"54",X"05",X"40",X"54",X"05",X"40",X"00",
		X"51",X"50",X"15",X"01",X"50",X"15",X"00",X"00",X"55",X"40",X"54",X"05",X"40",X"54",X"00",X"00",
		X"55",X"01",X"50",X"15",X"01",X"50",X"00",X"00",X"54",X"05",X"40",X"54",X"05",X"40",X"00",X"00",
		X"50",X"15",X"01",X"50",X"15",X"00",X"00",X"00",X"50",X"54",X"05",X"40",X"54",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"54",X"05",X"40",X"54",X"05",X"40",X"54",X"05",X"15",X"01",X"50",X"15",X"01",X"50",X"15",X"05",
		X"05",X"40",X"54",X"05",X"40",X"54",X"05",X"45",X"01",X"50",X"15",X"01",X"50",X"15",X"01",X"55",
		X"00",X"54",X"05",X"40",X"54",X"05",X"40",X"55",X"00",X"15",X"01",X"50",X"15",X"01",X"50",X"15",
		X"00",X"05",X"40",X"54",X"05",X"40",X"54",X"05",X"00",X"01",X"50",X"15",X"01",X"50",X"15",X"05",
		X"00",X"00",X"54",X"05",X"40",X"54",X"05",X"45",X"00",X"00",X"15",X"01",X"50",X"15",X"01",X"55",
		X"00",X"00",X"05",X"40",X"54",X"05",X"40",X"55",X"00",X"00",X"01",X"50",X"15",X"01",X"50",X"15",
		X"00",X"00",X"00",X"54",X"05",X"40",X"54",X"05",X"00",X"00",X"00",X"15",X"01",X"50",X"15",X"05",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"50",X"15",X"01",X"50",X"15",X"01",X"50",X"15",X"50",X"54",X"05",X"40",X"54",X"05",X"40",X"54",
		X"51",X"50",X"15",X"01",X"50",X"15",X"01",X"50",X"55",X"40",X"54",X"05",X"40",X"54",X"05",X"40",
		X"55",X"01",X"50",X"15",X"01",X"50",X"15",X"00",X"54",X"05",X"40",X"54",X"05",X"40",X"54",X"00",
		X"50",X"15",X"01",X"50",X"15",X"01",X"50",X"00",X"50",X"54",X"05",X"40",X"54",X"05",X"40",X"00",
		X"51",X"50",X"15",X"01",X"50",X"15",X"00",X"00",X"55",X"40",X"54",X"05",X"40",X"54",X"00",X"00",
		X"55",X"01",X"50",X"15",X"01",X"50",X"00",X"00",X"54",X"05",X"40",X"54",X"05",X"40",X"00",X"00",
		X"50",X"15",X"01",X"50",X"15",X"00",X"00",X"00",X"50",X"54",X"05",X"40",X"54",X"00",X"00",X"00",
		X"00",X"00",X"3F",X"FF",X"FF",X"FF",X"F5",X"40",X"03",X"D0",X"3F",X"FF",X"FF",X"FD",X"50",X"00",
		X"3F",X"D0",X"3F",X"FF",X"FF",X"54",X"00",X"00",X"3F",X"D0",X"3F",X"FF",X"D5",X"00",X"00",X"00",
		X"3F",X"D0",X"3F",X"F5",X"40",X"00",X"00",X"00",X"3F",X"D0",X"3F",X"D0",X"00",X"00",X"00",X"00",
		X"3F",X"D0",X"3F",X"D0",X"00",X"00",X"00",X"00",X"3F",X"D0",X"3F",X"D0",X"00",X"00",X"00",X"00",
		X"3F",X"D0",X"3F",X"D0",X"00",X"00",X"00",X"00",X"3F",X"D0",X"3F",X"D0",X"00",X"00",X"00",X"00",
		X"3F",X"D0",X"3F",X"D0",X"00",X"00",X"00",X"0F",X"3F",X"D0",X"3F",X"D0",X"00",X"00",X"0F",X"FF",
		X"3F",X"D0",X"3F",X"D0",X"00",X"0F",X"FF",X"FF",X"3F",X"D0",X"3F",X"F0",X"0F",X"FF",X"FF",X"FF",
		X"3F",X"D0",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"D0",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"03",X"FD",X"03",X"FD",X"03",X"FD",X"00",X"00",X"03",X"FD",X"03",X"FD",X"03",X"FD",X"00",
		X"00",X"03",X"FD",X"03",X"FD",X"03",X"FD",X"00",X"00",X"03",X"FD",X"03",X"FD",X"03",X"FD",X"00",
		X"00",X"03",X"FD",X"03",X"FD",X"03",X"FD",X"00",X"00",X"03",X"FD",X"03",X"FD",X"03",X"FD",X"00",
		X"00",X"03",X"FD",X"03",X"FD",X"03",X"FD",X"00",X"00",X"03",X"FD",X"03",X"FD",X"03",X"FD",X"00",
		X"00",X"0F",X"FD",X"03",X"FD",X"03",X"FD",X"00",X"0F",X"FF",X"FD",X"03",X"FD",X"03",X"FD",X"00",
		X"FF",X"FF",X"FD",X"03",X"FD",X"03",X"FD",X"00",X"FF",X"FF",X"FD",X"03",X"FD",X"03",X"FD",X"00",
		X"FF",X"FF",X"FD",X"03",X"FD",X"03",X"FD",X"00",X"FF",X"FF",X"F5",X"03",X"FD",X"03",X"FD",X"00",
		X"FF",X"F5",X"50",X"03",X"FD",X"03",X"FD",X"00",X"F5",X"50",X"00",X"03",X"FD",X"03",X"FD",X"00",
		X"00",X"00",X"3F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"3F",X"FF",X"FF",X"FC",X"00",X"00",
		X"00",X"00",X"3F",X"FF",X"FF",X"FF",X"D0",X"00",X"00",X"00",X"3F",X"FF",X"FF",X"FF",X"D0",X"00",
		X"00",X"00",X"3F",X"F5",X"7F",X"FF",X"D0",X"00",X"00",X"00",X"3F",X"D0",X"17",X"FF",X"D0",X"00",
		X"00",X"00",X"3F",X"D0",X"00",X"FF",X"D0",X"00",X"00",X"00",X"3F",X"D0",X"00",X"FF",X"D0",X"00",
		X"00",X"00",X"3F",X"D0",X"00",X"FF",X"D0",X"00",X"00",X"00",X"3F",X"D0",X"00",X"FF",X"D0",X"00",
		X"00",X"00",X"3F",X"D0",X"00",X"FF",X"D0",X"00",X"00",X"00",X"3D",X"50",X"00",X"FF",X"D0",X"00",
		X"00",X"00",X"54",X"00",X"00",X"FF",X"D0",X"00",X"00",X"00",X"00",X"00",X"03",X"FF",X"D0",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"D0",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"D0",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"05",X"40",X"54",X"05",X"45",X"00",X"00",X"00",X"01",X"50",X"15",X"01",X"55",
		X"00",X"00",X"00",X"00",X"54",X"05",X"40",X"55",X"00",X"00",X"00",X"00",X"15",X"01",X"50",X"15",
		X"00",X"00",X"00",X"00",X"05",X"40",X"54",X"05",X"00",X"00",X"00",X"00",X"01",X"50",X"15",X"05",
		X"00",X"00",X"00",X"00",X"00",X"54",X"05",X"45",X"00",X"00",X"00",X"00",X"00",X"15",X"01",X"55",
		X"00",X"00",X"00",X"00",X"00",X"05",X"40",X"55",X"00",X"00",X"00",X"00",X"00",X"01",X"50",X"15",
		X"00",X"00",X"00",X"00",X"00",X"00",X"54",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"15",X"05",
		X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"45",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"15",
		X"51",X"50",X"15",X"01",X"50",X"00",X"00",X"00",X"55",X"40",X"54",X"05",X"40",X"00",X"00",X"00",
		X"55",X"01",X"50",X"15",X"00",X"00",X"00",X"00",X"54",X"05",X"40",X"54",X"00",X"00",X"00",X"00",
		X"50",X"15",X"01",X"50",X"00",X"00",X"00",X"00",X"50",X"54",X"05",X"40",X"00",X"00",X"00",X"00",
		X"51",X"50",X"15",X"00",X"00",X"00",X"00",X"00",X"55",X"40",X"54",X"00",X"00",X"00",X"00",X"00",
		X"55",X"01",X"50",X"00",X"00",X"00",X"00",X"00",X"54",X"05",X"40",X"00",X"00",X"00",X"00",X"00",
		X"50",X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"54",X"00",X"00",X"00",X"00",X"00",X"00",
		X"51",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"05",X"40",X"54",X"05",X"45",X"00",X"00",X"00",X"01",X"50",X"15",X"01",X"55",
		X"00",X"00",X"00",X"00",X"54",X"05",X"40",X"55",X"00",X"00",X"00",X"00",X"15",X"01",X"50",X"15",
		X"00",X"00",X"00",X"00",X"05",X"40",X"54",X"05",X"00",X"00",X"00",X"00",X"01",X"50",X"15",X"05",
		X"00",X"00",X"00",X"00",X"00",X"54",X"05",X"45",X"00",X"00",X"00",X"00",X"00",X"15",X"01",X"55",
		X"00",X"00",X"00",X"00",X"00",X"05",X"40",X"55",X"00",X"00",X"00",X"00",X"00",X"01",X"50",X"15",
		X"00",X"00",X"00",X"00",X"00",X"00",X"54",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"15",X"05",
		X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"45",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",
		X"51",X"50",X"15",X"01",X"50",X"00",X"00",X"00",X"55",X"40",X"54",X"05",X"40",X"00",X"00",X"00",
		X"55",X"01",X"50",X"15",X"00",X"00",X"00",X"00",X"54",X"05",X"40",X"54",X"00",X"00",X"00",X"00",
		X"50",X"15",X"01",X"50",X"00",X"00",X"00",X"00",X"50",X"54",X"05",X"40",X"00",X"00",X"00",X"00",
		X"51",X"50",X"15",X"00",X"00",X"00",X"00",X"00",X"55",X"40",X"54",X"00",X"00",X"00",X"00",X"00",
		X"55",X"01",X"50",X"00",X"00",X"00",X"00",X"00",X"54",X"05",X"40",X"00",X"00",X"00",X"00",X"00",
		X"50",X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"54",X"00",X"00",X"00",X"00",X"00",X"00",
		X"51",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"D0",X"3F",X"FF",X"FF",X"FF",X"FF",X"F5",X"3F",X"D0",X"3F",X"FF",X"FF",X"FF",X"F5",X"50",
		X"3F",X"D0",X"3F",X"FF",X"FF",X"F5",X"50",X"00",X"3F",X"D0",X"3F",X"FF",X"F5",X"50",X"00",X"00",
		X"3F",X"D0",X"3F",X"F5",X"50",X"00",X"00",X"03",X"3F",X"D0",X"35",X"50",X"00",X"00",X"00",X"0F",
		X"3F",X"D0",X"10",X"00",X"00",X"0F",X"C0",X"3F",X"3F",X"D0",X"00",X"00",X"0F",X"FF",X"F0",X"3F",
		X"3F",X"D0",X"00",X"0F",X"FF",X"FF",X"FC",X"FF",X"3F",X"D0",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3F",X"D0",X"3F",X"FF",X"FF",X"FF",X"FF",X"FD",X"3F",X"D0",X"3F",X"FF",X"FF",X"FF",X"FF",X"F4",
		X"3F",X"D0",X"3F",X"FF",X"FF",X"F5",X"FF",X"D0",X"3F",X"D0",X"3F",X"FF",X"F5",X"50",X"3F",X"D0",
		X"3F",X"D0",X"3F",X"F5",X"50",X"00",X"3F",X"D0",X"3F",X"D0",X"3F",X"D0",X"00",X"00",X"3F",X"D0",
		X"50",X"00",X"01",X"03",X"FD",X"03",X"FD",X"00",X"00",X"00",X"0D",X"03",X"FD",X"03",X"FD",X"00",
		X"00",X"0F",X"FD",X"03",X"FD",X"03",X"FF",X"00",X"0F",X"FF",X"FD",X"03",X"FD",X"03",X"FF",X"FF",
		X"FF",X"FF",X"FD",X"03",X"FD",X"03",X"FF",X"FF",X"FF",X"FF",X"FD",X"03",X"FD",X"03",X"FF",X"FF",
		X"FF",X"FF",X"FD",X"03",X"FD",X"03",X"FF",X"FF",X"FF",X"FF",X"FD",X"03",X"FD",X"03",X"FF",X"FF",
		X"FF",X"FF",X"FD",X"03",X"FD",X"03",X"FF",X"FF",X"FD",X"5F",X"FD",X"03",X"FD",X"03",X"FF",X"55",
		X"54",X"03",X"FD",X"03",X"FD",X"03",X"55",X"00",X"00",X"03",X"FD",X"03",X"FD",X"05",X"00",X"00",
		X"00",X"03",X"FD",X"03",X"FD",X"00",X"00",X"00",X"00",X"03",X"FD",X"03",X"FD",X"00",X"00",X"FF",
		X"00",X"03",X"FD",X"03",X"FD",X"00",X"FF",X"FF",X"00",X"03",X"FD",X"03",X"FD",X"03",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"D0",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"D0",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"50",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"55",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"55",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"55",X"00",X"00",X"10",X"00",
		X"FF",X"FF",X"55",X"00",X"00",X"00",X"D0",X"00",X"FF",X"55",X"00",X"00",X"00",X"FF",X"D0",X"00",
		X"55",X"00",X"00",X"00",X"FF",X"FF",X"D0",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"D0",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"D0",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"D0",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"50",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"55",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"55",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"F5",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"15",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"55",
		X"54",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"15",X"00",X"00",X"00",X"00",X"00",X"01",X"55",
		X"05",X"40",X"00",X"00",X"00",X"00",X"05",X"45",X"01",X"50",X"00",X"00",X"00",X"00",X"05",X"55",
		X"00",X"54",X"00",X"00",X"00",X"00",X"15",X"55",X"00",X"15",X"00",X"00",X"00",X"00",X"54",X"15",
		X"00",X"05",X"40",X"00",X"00",X"00",X"54",X"05",X"00",X"01",X"50",X"00",X"00",X"01",X"55",X"05",
		X"00",X"00",X"54",X"00",X"00",X"05",X"45",X"45",X"00",X"00",X"15",X"00",X"00",X"05",X"01",X"55",
		X"00",X"00",X"05",X"40",X"00",X"15",X"40",X"55",X"00",X"00",X"01",X"50",X"00",X"55",X"50",X"15",
		X"00",X"00",X"00",X"54",X"00",X"50",X"54",X"05",X"00",X"00",X"00",X"15",X"01",X"50",X"15",X"05",
		X"54",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"05",
		X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"15",X"55",X"40",X"00",X"00",X"00",X"00",X"00",X"54",
		X"51",X"50",X"00",X"00",X"00",X"00",X"01",X"50",X"55",X"50",X"00",X"00",X"00",X"00",X"05",X"40",
		X"55",X"54",X"00",X"00",X"00",X"00",X"15",X"00",X"54",X"15",X"00",X"00",X"00",X"00",X"54",X"00",
		X"50",X"15",X"00",X"00",X"00",X"01",X"50",X"00",X"50",X"55",X"40",X"00",X"00",X"05",X"40",X"00",
		X"51",X"51",X"50",X"00",X"00",X"15",X"00",X"00",X"55",X"40",X"50",X"00",X"00",X"54",X"00",X"00",
		X"55",X"01",X"54",X"00",X"01",X"50",X"00",X"00",X"54",X"05",X"55",X"00",X"05",X"40",X"00",X"00",
		X"50",X"15",X"05",X"00",X"15",X"00",X"00",X"00",X"50",X"54",X"05",X"40",X"54",X"00",X"00",X"00",
		X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"15",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"55",
		X"54",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"15",X"00",X"00",X"00",X"00",X"00",X"01",X"55",
		X"05",X"40",X"00",X"00",X"00",X"00",X"05",X"45",X"01",X"50",X"00",X"00",X"00",X"00",X"05",X"55",
		X"00",X"54",X"00",X"00",X"00",X"00",X"15",X"55",X"00",X"15",X"00",X"00",X"00",X"00",X"54",X"15",
		X"00",X"05",X"40",X"00",X"00",X"00",X"54",X"05",X"00",X"01",X"50",X"00",X"00",X"01",X"55",X"05",
		X"00",X"00",X"54",X"00",X"00",X"05",X"45",X"45",X"00",X"00",X"15",X"00",X"00",X"05",X"01",X"55",
		X"00",X"00",X"05",X"40",X"00",X"15",X"40",X"55",X"00",X"00",X"01",X"50",X"00",X"55",X"50",X"15",
		X"00",X"00",X"00",X"54",X"00",X"50",X"54",X"05",X"00",X"00",X"00",X"15",X"01",X"50",X"15",X"05",
		X"54",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"05",
		X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"15",X"55",X"40",X"00",X"00",X"00",X"00",X"00",X"54",
		X"51",X"50",X"00",X"00",X"00",X"00",X"01",X"50",X"55",X"50",X"00",X"00",X"00",X"00",X"05",X"40",
		X"55",X"54",X"00",X"00",X"00",X"00",X"15",X"00",X"54",X"15",X"00",X"00",X"00",X"00",X"54",X"00",
		X"50",X"15",X"00",X"00",X"00",X"01",X"50",X"00",X"50",X"55",X"40",X"00",X"00",X"05",X"40",X"00",
		X"51",X"51",X"50",X"00",X"00",X"15",X"00",X"00",X"55",X"40",X"50",X"00",X"00",X"54",X"00",X"00",
		X"55",X"01",X"54",X"00",X"01",X"50",X"00",X"00",X"54",X"05",X"55",X"00",X"05",X"40",X"00",X"00",
		X"50",X"15",X"05",X"00",X"15",X"00",X"00",X"00",X"50",X"54",X"05",X"40",X"54",X"00",X"00",X"00",
		X"3F",X"D0",X"3F",X"D0",X"00",X"00",X"3F",X"D0",X"3F",X"D0",X"3F",X"D0",X"00",X"00",X"3F",X"D0",
		X"3F",X"D0",X"3F",X"D0",X"00",X"00",X"3F",X"D0",X"3F",X"D0",X"3F",X"D0",X"00",X"00",X"3F",X"D0",
		X"3F",X"D0",X"3F",X"F0",X"00",X"00",X"FF",X"F0",X"3F",X"D0",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3F",X"D0",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"D0",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3F",X"D0",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"D0",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3F",X"D0",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"D0",X"15",X"55",X"55",X"55",X"55",X"55",
		X"3F",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"D0",X"3F",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"03",X"FD",X"03",X"FD",X"03",X"FF",X"FF",X"00",X"03",X"FD",X"03",X"FD",X"03",X"FF",X"FF",
		X"00",X"03",X"FD",X"03",X"FD",X"03",X"FF",X"FF",X"00",X"03",X"FD",X"03",X"FD",X"03",X"FF",X"D5",
		X"00",X"03",X"FD",X"03",X"FD",X"03",X"FF",X"40",X"FF",X"FF",X"FD",X"03",X"FD",X"03",X"FF",X"40",
		X"FF",X"FF",X"FD",X"03",X"FD",X"03",X"FF",X"40",X"FF",X"FF",X"FD",X"03",X"FD",X"03",X"FF",X"40",
		X"FF",X"FF",X"FD",X"03",X"FD",X"03",X"FF",X"40",X"FF",X"FF",X"FD",X"03",X"FD",X"03",X"FF",X"40",
		X"FF",X"FF",X"FD",X"03",X"FD",X"03",X"FF",X"C0",X"55",X"55",X"55",X"03",X"FD",X"03",X"FF",X"FF",
		X"00",X"00",X"00",X"03",X"FD",X"03",X"FF",X"FF",X"00",X"00",X"00",X"03",X"FD",X"03",X"FF",X"FF",
		X"00",X"00",X"01",X"03",X"FD",X"03",X"FF",X"FF",X"00",X"00",X"0D",X"03",X"FD",X"05",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"D0",X"00",X"00",X"00",X"00",X"FF",X"55",X"3F",X"D0",X"00",X"00",X"00",X"00",
		X"55",X"00",X"3F",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"D0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"3F",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"D0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"3F",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"D0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"3F",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"D0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"3F",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"D0",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"3F",X"D0",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"D0",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"F0",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"05",X"45",X"54",X"05",X"45",X"00",X"00",X"00",X"01",X"55",X"15",X"01",X"55",
		X"00",X"00",X"00",X"00",X"55",X"05",X"40",X"55",X"00",X"00",X"00",X"00",X"15",X"01",X"50",X"15",
		X"00",X"00",X"00",X"00",X"05",X"40",X"54",X"05",X"00",X"00",X"00",X"00",X"01",X"50",X"15",X"05",
		X"00",X"00",X"00",X"00",X"00",X"54",X"05",X"45",X"00",X"00",X"00",X"00",X"00",X"15",X"01",X"55",
		X"00",X"00",X"00",X"00",X"00",X"05",X"40",X"55",X"00",X"00",X"00",X"00",X"00",X"01",X"50",X"15",
		X"00",X"00",X"00",X"00",X"00",X"00",X"54",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"15",X"05",
		X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"45",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"15",
		X"51",X"50",X"15",X"51",X"50",X"00",X"00",X"00",X"55",X"40",X"54",X"55",X"40",X"00",X"00",X"00",
		X"55",X"01",X"50",X"55",X"00",X"00",X"00",X"00",X"54",X"05",X"40",X"54",X"00",X"00",X"00",X"00",
		X"50",X"15",X"01",X"50",X"00",X"00",X"00",X"00",X"50",X"54",X"05",X"40",X"00",X"00",X"00",X"00",
		X"51",X"50",X"15",X"00",X"00",X"00",X"00",X"00",X"55",X"40",X"54",X"00",X"00",X"00",X"00",X"00",
		X"55",X"01",X"50",X"00",X"00",X"00",X"00",X"00",X"54",X"05",X"40",X"00",X"00",X"00",X"00",X"00",
		X"50",X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"54",X"00",X"00",X"00",X"00",X"00",X"00",
		X"51",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"05",X"45",X"54",X"05",X"45",X"00",X"00",X"00",X"01",X"55",X"15",X"01",X"55",
		X"00",X"00",X"00",X"00",X"55",X"05",X"40",X"55",X"00",X"00",X"00",X"00",X"15",X"01",X"50",X"15",
		X"00",X"00",X"00",X"00",X"05",X"40",X"54",X"05",X"00",X"00",X"00",X"00",X"01",X"50",X"15",X"05",
		X"00",X"00",X"00",X"00",X"00",X"54",X"05",X"45",X"00",X"00",X"00",X"00",X"00",X"15",X"01",X"55",
		X"00",X"00",X"00",X"00",X"00",X"05",X"40",X"55",X"00",X"00",X"00",X"00",X"00",X"01",X"50",X"15",
		X"00",X"00",X"00",X"00",X"00",X"00",X"54",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"15",X"05",
		X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"45",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"15",
		X"51",X"50",X"15",X"51",X"50",X"00",X"00",X"00",X"55",X"40",X"54",X"55",X"40",X"00",X"00",X"00",
		X"55",X"01",X"50",X"55",X"00",X"00",X"00",X"00",X"54",X"05",X"40",X"54",X"00",X"00",X"00",X"00",
		X"50",X"15",X"01",X"50",X"00",X"00",X"00",X"00",X"50",X"54",X"05",X"40",X"00",X"00",X"00",X"00",
		X"51",X"50",X"15",X"00",X"00",X"00",X"00",X"00",X"55",X"40",X"54",X"00",X"00",X"00",X"00",X"00",
		X"55",X"01",X"50",X"00",X"00",X"00",X"00",X"00",X"54",X"05",X"40",X"00",X"00",X"00",X"00",X"00",
		X"50",X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"54",X"00",X"00",X"00",X"00",X"00",X"00",
		X"51",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"D0",X"3F",X"FF",X"FF",X"FF",X"C0",X"00",X"3F",X"D0",X"3F",X"FF",X"FF",X"FF",X"F0",X"00",
		X"3F",X"D0",X"3F",X"FF",X"FF",X"FF",X"FC",X"0F",X"3F",X"D0",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3F",X"D0",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"D0",X"3F",X"F5",X"55",X"5F",X"FF",X"FF",
		X"3F",X"D0",X"3F",X"D0",X"00",X"07",X"FF",X"FF",X"3F",X"D0",X"3F",X"D0",X"00",X"01",X"FF",X"FF",
		X"3F",X"D0",X"3F",X"D0",X"00",X"00",X"3F",X"F5",X"3F",X"D0",X"3F",X"D0",X"00",X"00",X"3F",X"D0",
		X"3F",X"D0",X"3F",X"D0",X"00",X"00",X"3F",X"D0",X"3F",X"D0",X"3F",X"D0",X"00",X"00",X"3F",X"D0",
		X"3F",X"D0",X"3F",X"D0",X"00",X"00",X"3F",X"D0",X"3F",X"D0",X"3F",X"D0",X"00",X"00",X"3F",X"D0",
		X"3F",X"D0",X"3F",X"D0",X"00",X"00",X"3F",X"D0",X"3F",X"D0",X"3F",X"F0",X"00",X"00",X"FF",X"F0",
		X"00",X"0F",X"FD",X"03",X"FD",X"00",X"55",X"FF",X"0F",X"FF",X"FD",X"03",X"FD",X"00",X"00",X"55",
		X"FF",X"FF",X"FD",X"03",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FD",X"03",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"FD",X"03",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"F5",X"03",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"F5",X"50",X"03",X"FF",X"FF",X"FF",X"FF",X"F5",X"50",X"00",X"03",X"FF",X"FF",X"FF",X"FF",
		X"50",X"00",X"00",X"03",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"03",X"FF",X"55",X"FF",X"FF",
		X"00",X"00",X"00",X"03",X"FD",X"00",X"55",X"FF",X"00",X"00",X"00",X"03",X"FD",X"00",X"00",X"55",
		X"00",X"00",X"00",X"03",X"FD",X"0F",X"00",X"00",X"00",X"00",X"00",X"03",X"FD",X"0F",X"FF",X"00",
		X"00",X"00",X"00",X"03",X"FD",X"0F",X"FF",X"FF",X"00",X"00",X"01",X"03",X"FD",X"0F",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"10",X"00",
		X"55",X"FF",X"FF",X"FF",X"FF",X"FF",X"D0",X"00",X"00",X"55",X"FF",X"FF",X"FF",X"FF",X"D0",X"00",
		X"00",X"00",X"55",X"FF",X"FF",X"FF",X"D0",X"00",X"00",X"00",X"00",X"55",X"FF",X"FF",X"D0",X"00",
		X"FF",X"00",X"00",X"00",X"55",X"FF",X"D0",X"00",X"FF",X"FF",X"00",X"00",X"00",X"55",X"D0",X"00",
		X"FF",X"FF",X"FF",X"00",X"00",X"00",X"50",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"10",X"00",
		X"55",X"FF",X"FF",X"FF",X"FF",X"FF",X"D0",X"00",X"00",X"55",X"FF",X"FF",X"FF",X"FF",X"D0",X"00",
		X"00",X"00",X"55",X"FF",X"FF",X"FF",X"D0",X"00",X"FF",X"00",X"00",X"55",X"FF",X"FF",X"D0",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"15",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"15",
		X"54",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"01",X"55",
		X"55",X"40",X"00",X"00",X"00",X"00",X"01",X"45",X"51",X"50",X"00",X"00",X"00",X"00",X"05",X"55",
		X"50",X"54",X"00",X"00",X"00",X"00",X"15",X"55",X"50",X"15",X"00",X"00",X"00",X"00",X"14",X"15",
		X"54",X"05",X"40",X"00",X"00",X"00",X"54",X"05",X"55",X"01",X"50",X"00",X"00",X"01",X"55",X"05",
		X"55",X"40",X"54",X"00",X"00",X"01",X"45",X"45",X"51",X"50",X"15",X"00",X"00",X"05",X"41",X"55",
		X"50",X"54",X"05",X"40",X"00",X"15",X"40",X"55",X"50",X"15",X"01",X"50",X"00",X"15",X"50",X"15",
		X"54",X"05",X"40",X"54",X"00",X"54",X"54",X"05",X"55",X"01",X"50",X"15",X"01",X"50",X"15",X"05",
		X"54",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"54",X"00",X"00",X"00",X"00",X"00",X"00",X"05",
		X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"15",X"55",X"40",X"00",X"00",X"00",X"00",X"00",X"55",
		X"51",X"40",X"00",X"00",X"00",X"00",X"01",X"55",X"55",X"50",X"00",X"00",X"00",X"00",X"05",X"45",
		X"55",X"54",X"00",X"00",X"00",X"00",X"15",X"05",X"54",X"14",X"00",X"00",X"00",X"00",X"54",X"05",
		X"50",X"15",X"00",X"00",X"00",X"01",X"50",X"15",X"50",X"55",X"40",X"00",X"00",X"05",X"40",X"55",
		X"51",X"51",X"40",X"00",X"00",X"15",X"01",X"55",X"55",X"41",X"50",X"00",X"00",X"54",X"05",X"45",
		X"55",X"01",X"54",X"00",X"01",X"50",X"15",X"05",X"54",X"05",X"54",X"00",X"05",X"40",X"54",X"05",
		X"50",X"15",X"15",X"00",X"15",X"01",X"50",X"15",X"50",X"54",X"05",X"40",X"54",X"05",X"40",X"55",
		X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"15",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"15",
		X"54",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"01",X"55",
		X"55",X"40",X"00",X"00",X"00",X"00",X"01",X"45",X"51",X"50",X"00",X"00",X"00",X"00",X"05",X"55",
		X"50",X"54",X"00",X"00",X"00",X"00",X"15",X"55",X"50",X"15",X"00",X"00",X"00",X"00",X"14",X"15",
		X"54",X"05",X"40",X"00",X"00",X"00",X"54",X"05",X"55",X"01",X"50",X"00",X"00",X"01",X"55",X"05",
		X"55",X"40",X"54",X"00",X"00",X"01",X"45",X"45",X"51",X"50",X"15",X"00",X"00",X"05",X"41",X"55",
		X"50",X"54",X"05",X"40",X"00",X"15",X"40",X"55",X"50",X"15",X"01",X"50",X"00",X"15",X"50",X"15",
		X"54",X"05",X"40",X"54",X"00",X"54",X"54",X"05",X"55",X"01",X"50",X"15",X"01",X"50",X"15",X"05",
		X"54",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"54",X"00",X"00",X"00",X"00",X"00",X"00",X"05",
		X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"15",X"55",X"40",X"00",X"00",X"00",X"00",X"00",X"55",
		X"51",X"40",X"00",X"00",X"00",X"00",X"01",X"55",X"55",X"50",X"00",X"00",X"00",X"00",X"05",X"45",
		X"55",X"54",X"00",X"00",X"00",X"00",X"15",X"05",X"54",X"14",X"00",X"00",X"00",X"00",X"54",X"05",
		X"50",X"15",X"00",X"00",X"00",X"01",X"50",X"15",X"50",X"55",X"40",X"00",X"00",X"05",X"40",X"55",
		X"51",X"51",X"40",X"00",X"00",X"15",X"01",X"55",X"55",X"41",X"50",X"00",X"00",X"54",X"05",X"45",
		X"55",X"01",X"54",X"00",X"01",X"50",X"15",X"05",X"54",X"05",X"54",X"00",X"05",X"40",X"54",X"05",
		X"50",X"15",X"15",X"00",X"15",X"01",X"50",X"15",X"50",X"54",X"05",X"40",X"54",X"05",X"40",X"55",
		X"3F",X"D0",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"D0",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3F",X"D0",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"D0",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3F",X"D0",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"D0",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3F",X"D0",X"15",X"55",X"55",X"55",X"55",X"55",X"3F",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"D0",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"D0",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3F",X"D0",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"D0",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3F",X"D0",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"D0",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FD",X"03",X"FD",X"0F",X"FF",X"FF",X"FF",X"FF",X"FD",X"03",X"FD",X"0F",X"FF",X"FF",
		X"FF",X"FF",X"FD",X"03",X"FD",X"0F",X"FF",X"FF",X"FF",X"FF",X"FD",X"03",X"FD",X"0F",X"FF",X"FF",
		X"FF",X"FF",X"FD",X"03",X"FD",X"0F",X"FF",X"FF",X"FF",X"FF",X"FD",X"03",X"FD",X"0F",X"FF",X"FF",
		X"55",X"55",X"55",X"03",X"FD",X"0F",X"FF",X"FF",X"00",X"00",X"00",X"03",X"FD",X"0F",X"FF",X"FF",
		X"00",X"00",X"00",X"03",X"FD",X"0F",X"FF",X"FF",X"00",X"00",X"00",X"03",X"FD",X"0F",X"FF",X"FF",
		X"FF",X"FF",X"FD",X"03",X"FD",X"0F",X"FF",X"FF",X"FF",X"FF",X"FD",X"03",X"FD",X"0F",X"FF",X"FF",
		X"FF",X"FF",X"FD",X"03",X"FD",X"0F",X"FF",X"FF",X"FF",X"FF",X"FD",X"03",X"FD",X"0F",X"FF",X"FF",
		X"FF",X"FF",X"FD",X"05",X"7D",X"0F",X"FF",X"FF",X"FF",X"FF",X"FD",X"00",X"15",X"0F",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"55",X"FF",X"D0",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"55",X"D0",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"50",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"40",X"54",X"05",X"41",X"54",X"05",X"45",X"51",X"50",X"15",X"01",X"55",X"55",X"01",X"55",
		X"50",X"54",X"05",X"40",X"55",X"05",X"40",X"55",X"50",X"15",X"01",X"50",X"15",X"01",X"50",X"15",
		X"54",X"05",X"40",X"54",X"05",X"40",X"54",X"05",X"55",X"01",X"50",X"15",X"01",X"50",X"15",X"05",
		X"55",X"40",X"54",X"05",X"40",X"54",X"05",X"45",X"51",X"50",X"15",X"01",X"50",X"15",X"01",X"55",
		X"50",X"54",X"05",X"40",X"54",X"05",X"40",X"55",X"50",X"15",X"01",X"50",X"15",X"01",X"50",X"15",
		X"54",X"05",X"40",X"54",X"05",X"40",X"54",X"05",X"55",X"01",X"50",X"15",X"01",X"50",X"15",X"05",
		X"55",X"40",X"54",X"05",X"40",X"54",X"05",X"45",X"51",X"50",X"15",X"01",X"50",X"15",X"01",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"51",X"50",X"15",X"41",X"50",X"15",X"01",X"55",X"55",X"40",X"55",X"55",X"40",X"54",X"05",X"45",
		X"55",X"01",X"50",X"55",X"01",X"50",X"15",X"05",X"54",X"05",X"40",X"54",X"05",X"40",X"54",X"05",
		X"50",X"15",X"01",X"50",X"15",X"01",X"50",X"15",X"50",X"54",X"05",X"40",X"54",X"05",X"40",X"55",
		X"51",X"50",X"15",X"01",X"50",X"15",X"01",X"55",X"55",X"40",X"54",X"05",X"40",X"54",X"05",X"45",
		X"55",X"01",X"50",X"15",X"01",X"50",X"15",X"05",X"54",X"05",X"40",X"54",X"05",X"40",X"54",X"05",
		X"50",X"15",X"01",X"50",X"15",X"01",X"50",X"15",X"50",X"54",X"05",X"40",X"54",X"05",X"40",X"55",
		X"51",X"50",X"15",X"01",X"50",X"15",X"01",X"55",X"55",X"40",X"54",X"05",X"40",X"54",X"05",X"45",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"40",X"54",X"05",X"41",X"54",X"05",X"45",X"51",X"50",X"15",X"01",X"55",X"55",X"01",X"55",
		X"50",X"54",X"05",X"40",X"55",X"05",X"40",X"55",X"50",X"15",X"01",X"50",X"15",X"01",X"50",X"15",
		X"54",X"05",X"40",X"54",X"05",X"40",X"54",X"05",X"55",X"01",X"50",X"15",X"01",X"50",X"15",X"05",
		X"55",X"40",X"54",X"05",X"40",X"54",X"05",X"45",X"51",X"50",X"15",X"01",X"50",X"15",X"01",X"55",
		X"50",X"54",X"05",X"40",X"54",X"05",X"40",X"55",X"50",X"15",X"01",X"50",X"15",X"01",X"50",X"15",
		X"54",X"05",X"40",X"54",X"05",X"40",X"54",X"05",X"55",X"01",X"50",X"15",X"01",X"50",X"15",X"05",
		X"55",X"40",X"54",X"05",X"40",X"54",X"05",X"45",X"51",X"50",X"15",X"01",X"50",X"15",X"01",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"51",X"50",X"15",X"41",X"50",X"15",X"01",X"55",X"55",X"40",X"55",X"55",X"40",X"54",X"05",X"45",
		X"55",X"01",X"50",X"55",X"01",X"50",X"15",X"05",X"54",X"05",X"40",X"54",X"05",X"40",X"54",X"05",
		X"50",X"15",X"01",X"50",X"15",X"01",X"50",X"15",X"50",X"54",X"05",X"40",X"54",X"05",X"40",X"55",
		X"51",X"50",X"15",X"01",X"50",X"15",X"01",X"55",X"55",X"40",X"54",X"05",X"40",X"54",X"05",X"45",
		X"55",X"01",X"50",X"15",X"01",X"50",X"15",X"05",X"54",X"05",X"40",X"54",X"05",X"40",X"54",X"05",
		X"50",X"15",X"01",X"50",X"15",X"01",X"50",X"15",X"50",X"54",X"05",X"40",X"54",X"05",X"40",X"55",
		X"51",X"50",X"15",X"01",X"50",X"15",X"01",X"55",X"55",X"40",X"54",X"05",X"40",X"54",X"05",X"45",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"3F",X"D0",X"55",X"55",X"55",X"55",X"55",X"55",X"3F",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"D0",X"30",X"00",X"00",X"00",X"00",X"00",X"3F",X"D0",X"3F",X"F0",X"00",X"00",X"00",X"00",
		X"3F",X"D0",X"3F",X"FF",X"F0",X"00",X"00",X"00",X"3F",X"D0",X"3F",X"FF",X"FF",X"F0",X"00",X"00",
		X"3F",X"D0",X"3F",X"FF",X"FF",X"FF",X"F0",X"00",X"3F",X"D0",X"3F",X"FF",X"FF",X"FF",X"FF",X"F0",
		X"3F",X"D0",X"5F",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"D0",X"05",X"5F",X"FF",X"FF",X"FF",X"FF",
		X"3F",X"D0",X"00",X"05",X"5F",X"FF",X"FF",X"FF",X"3F",X"F0",X"00",X"00",X"05",X"5F",X"FF",X"FF",
		X"3F",X"FF",X"F0",X"00",X"00",X"05",X"5F",X"FF",X"3F",X"FF",X"FF",X"F0",X"00",X"00",X"05",X"5F",
		X"55",X"57",X"FD",X"00",X"00",X"0F",X"FF",X"FF",X"00",X"03",X"FD",X"0F",X"00",X"00",X"FF",X"FF",
		X"00",X"03",X"FD",X"0F",X"FF",X"00",X"00",X"FF",X"00",X"03",X"FD",X"0F",X"FF",X"FF",X"00",X"00",
		X"00",X"03",X"FD",X"0F",X"FF",X"FF",X"FF",X"00",X"00",X"03",X"FD",X"0F",X"FF",X"FF",X"FF",X"FF",
		X"00",X"03",X"FD",X"0F",X"FF",X"FF",X"FF",X"FF",X"00",X"03",X"FD",X"0F",X"FF",X"FF",X"FF",X"FF",
		X"00",X"03",X"FD",X"0F",X"FF",X"FF",X"FF",X"FF",X"00",X"03",X"FD",X"0F",X"FF",X"FF",X"FF",X"FF",
		X"F0",X"0F",X"FD",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"0F",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FD",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"0F",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FD",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"0F",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",
		X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"F0",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"F0",X"00",
		X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"F0",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"F0",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",
		X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"03",X"FF",
		X"FF",X"FF",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"FF",X"FF",X"FF",X"00",X"00",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"AA",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"2A",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"00",X"00",X"AA",X"A0",X"00",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"A0",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"00",
		X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"A0",X"00",X"FF",X"00",X"00",X"AA",X"AA",X"AA",X"A0",X"00",
		X"FF",X"FF",X"00",X"00",X"AA",X"AA",X"A0",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"AA",X"A0",X"00",
		X"FF",X"FF",X"FF",X"FC",X"00",X"00",X"A0",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",
		X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"F0",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"F0",X"00",
		X"FF",X"FF",X"FF",X"FF",X"CC",X"08",X"20",X"82",X"FF",X"FF",X"FF",X"FF",X"30",X"0A",X"A0",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"CC",X"C8",X"20",X"96",X"FF",X"FF",X"FF",X"FF",X"33",X"08",X"2A",X"96",
		X"FF",X"FF",X"FF",X"FF",X"C0",X"C8",X"25",X"96",X"FF",X"FF",X"FF",X"FF",X"00",X"0A",X"A5",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"AA",X"A8",X"25",X"82",X"FF",X"FF",X"FF",X"FF",X"98",X"0A",X"2A",X"82",
		X"FF",X"FF",X"FF",X"FF",X"98",X"09",X"A0",X"82",X"FF",X"FF",X"FF",X"FF",X"AA",X"AA",X"A0",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"80",X"80",X"88",X"96",X"FF",X"FF",X"FF",X"FF",X"80",X"80",X"82",X"96",
		X"FF",X"FF",X"FF",X"FF",X"AA",X"AA",X"AA",X"96",X"FF",X"FF",X"FF",X"FF",X"88",X"09",X"58",X"26",
		X"FF",X"FF",X"FF",X"FF",X"88",X"09",X"58",X"0A",X"FF",X"FF",X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"FF",X"FF",X"FF",X"F0",X"00",X"00",X"05",X"3F",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",X"00",
		X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",
		X"3F",X"F5",X"5F",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"D0",X"05",X"5F",X"FF",X"FF",X"FF",X"FF",
		X"3F",X"D0",X"00",X"05",X"5F",X"FF",X"FF",X"FF",X"3F",X"D0",X"00",X"00",X"05",X"5F",X"FF",X"FF",
		X"3F",X"D0",X"AA",X"00",X"00",X"05",X"5F",X"FF",X"3F",X"D0",X"AA",X"AA",X"00",X"00",X"05",X"5F",
		X"3F",X"D0",X"AA",X"AA",X"AA",X"00",X"00",X"05",X"3F",X"D0",X"AA",X"AA",X"AA",X"AA",X"00",X"00",
		X"3F",X"D0",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"3F",X"D0",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"3F",X"D0",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"3F",X"D0",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"5F",X"FF",X"FD",X"00",X"FF",X"FF",X"FF",X"FF",X"05",X"5F",X"FD",X"00",X"00",X"FF",X"FF",X"FF",
		X"00",X"05",X"5D",X"0F",X"00",X"00",X"FF",X"FF",X"00",X"00",X"05",X"0F",X"FF",X"00",X"00",X"FF",
		X"F0",X"00",X"00",X"0F",X"FF",X"FF",X"00",X"00",X"FF",X"F0",X"00",X"0F",X"FF",X"FF",X"FF",X"00",
		X"FF",X"FF",X"F1",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"0F",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FD",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"0F",X"FF",X"FF",X"FF",X"FF",
		X"5F",X"FF",X"FD",X"0F",X"FF",X"FF",X"FF",X"FF",X"05",X"5F",X"FD",X"0F",X"FF",X"FF",X"FF",X"FF",
		X"00",X"05",X"5D",X"0F",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"05",X"0F",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"00",X"00",X"0F",X"FF",X"FF",X"FF",X"FF",X"AA",X"AA",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"F0",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"F0",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"F0",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"F0",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",
		X"82",X"09",X"63",X"33",X"33",X"33",X"33",X"33",X"82",X"A9",X"60",X"CC",X"CC",X"CC",X"0C",X"CC",
		X"82",X"09",X"60",X"33",X"33",X"33",X"03",X"33",X"AA",X"0A",X"A0",X"CC",X"C0",X"CC",X"CC",X"CC",
		X"96",X"08",X"23",X"03",X"33",X"03",X"33",X"03",X"96",X"A8",X"20",X"00",X"00",X"00",X"00",X"00",
		X"96",X"08",X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"08",X"A0",X"25",X"60",X"20",X"20",X"20",
		X"82",X"0A",X"20",X"25",X"60",X"20",X"20",X"20",X"82",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"82",X"26",X"02",X"56",X"02",X"56",X"02",X"56",X"AA",X"96",X"02",X"56",X"02",X"56",X"02",X"56",
		X"96",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"98",X"25",X"60",X"20",X"20",X"25",X"60",X"20",
		X"A0",X"25",X"60",X"20",X"20",X"25",X"60",X"20",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"33",X"33",X"33",X"33",X"33",X"0A",X"A0",X"AA",X"CC",X"CC",X"CC",X"CC",X"CC",X"08",X"20",X"82",
		X"33",X"33",X"33",X"33",X"30",X"08",X"2A",X"82",X"C0",X"CC",X"CC",X"C0",X"CC",X"C8",X"25",X"82",
		X"33",X"30",X"30",X"33",X"03",X"0A",X"A5",X"AA",X"00",X"00",X"00",X"00",X"00",X"08",X"25",X"82",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"2A",X"82",X"20",X"25",X"60",X"25",X"60",X"26",X"20",X"82",
		X"20",X"25",X"60",X"25",X"60",X"25",X"A0",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"96",
		X"02",X"02",X"02",X"02",X"02",X"56",X"08",X"96",X"02",X"02",X"02",X"02",X"02",X"56",X"02",X"96",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"96",X"20",X"20",X"25",X"60",X"20",X"20",X"20",X"26",
		X"20",X"20",X"25",X"60",X"20",X"20",X"20",X"0A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FB",X"AA",X"FF",X"FF",X"EE",X"BF",X"FF",X"FF",X"FE",X"AA",X"FF",X"FF",X"FA",X"BF",X"FF",X"FF",
		X"FB",X"AA",X"FF",X"FF",X"EE",X"BF",X"FF",X"FF",X"FE",X"AA",X"FF",X"FF",X"FA",X"BF",X"FF",X"FF",
		X"FB",X"AA",X"FF",X"FF",X"EE",X"BF",X"FF",X"FF",X"FE",X"AA",X"FF",X"FF",X"FA",X"BF",X"FF",X"FF",
		X"FB",X"AA",X"FF",X"FF",X"EE",X"BF",X"FF",X"FF",X"FE",X"AA",X"FF",X"FF",X"FA",X"BF",X"FF",X"FF",
		X"FB",X"AA",X"FF",X"FF",X"EE",X"BF",X"FF",X"FF",X"FE",X"AA",X"FF",X"FF",X"FA",X"BF",X"FF",X"FF",
		X"FB",X"AA",X"FF",X"FF",X"EE",X"BF",X"FF",X"FF",X"FE",X"AA",X"FF",X"FF",X"FA",X"EA",X"AA",X"AA",
		X"FB",X"AA",X"FF",X"FF",X"EF",X"AA",X"AA",X"AA",X"FE",X"AA",X"FF",X"FF",X"FB",X"BB",X"BB",X"BB",
		X"FB",X"AA",X"FF",X"FF",X"EE",X"EE",X"EE",X"EE",X"FE",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FE",X"AF",X"FF",X"FF",X"AA",X"BF",X"FF",X"FF",X"FE",X"BB",X"FF",X"FF",X"AA",X"EF",
		X"FF",X"FF",X"FE",X"AF",X"FF",X"FF",X"AA",X"BF",X"FF",X"FF",X"FE",X"BB",X"FF",X"FF",X"AA",X"EF",
		X"FF",X"FF",X"FE",X"AF",X"FF",X"FF",X"AA",X"BF",X"FF",X"FF",X"FE",X"BB",X"FF",X"FF",X"AA",X"EF",
		X"FF",X"FF",X"FE",X"AF",X"FF",X"FF",X"AA",X"BF",X"FF",X"FF",X"FE",X"BB",X"FF",X"FF",X"AA",X"EF",
		X"FF",X"FF",X"FE",X"AF",X"FF",X"FF",X"AA",X"BF",X"FF",X"FF",X"FE",X"BB",X"FF",X"FF",X"AA",X"EF",
		X"FF",X"FF",X"FE",X"AF",X"FF",X"FF",X"AA",X"BF",X"AA",X"AA",X"AB",X"BB",X"FF",X"FF",X"AA",X"EF",
		X"AA",X"AA",X"AA",X"EF",X"FF",X"FF",X"AA",X"BF",X"BB",X"BB",X"BB",X"BB",X"FF",X"FF",X"AA",X"EF",
		X"EE",X"EE",X"EE",X"EF",X"FF",X"FF",X"AA",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"EF",
		X"82",X"08",X"20",X"C0",X"00",X"00",X"00",X"00",X"AA",X"0A",X"A3",X"00",X"00",X"00",X"00",X"00",
		X"82",X"A8",X"20",X"00",X"00",X"00",X"00",X"00",X"82",X"58",X"20",X"0C",X"00",X"00",X"00",X"00",
		X"82",X"58",X"20",X"00",X"00",X"00",X"00",X"00",X"AA",X"5A",X"A0",X"00",X"00",X"00",X"00",X"00",
		X"82",X"58",X"2A",X"AA",X"00",X"00",X"00",X"00",X"82",X"A8",X"A5",X"62",X"00",X"00",X"00",X"00",
		X"82",X"0A",X"25",X"62",X"00",X"00",X"00",X"00",X"AA",X"0A",X"AA",X"AA",X"00",X"00",X"00",X"00",
		X"96",X"22",X"02",X"56",X"00",X"00",X"00",X"00",X"96",X"82",X"02",X"56",X"00",X"00",X"00",X"00",
		X"96",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"00",X"98",X"25",X"60",X"22",X"00",X"00",X"00",X"00",
		X"A0",X"25",X"60",X"22",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"00",
		X"3F",X"D0",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"3F",X"D0",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"3F",X"D0",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"3F",X"D0",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"3F",X"D0",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"3F",X"D0",X"AA",X"00",X"00",X"AA",X"AA",X"AA",
		X"3F",X"D0",X"AA",X"AA",X"00",X"00",X"AA",X"AA",X"3F",X"D0",X"AA",X"AA",X"AA",X"00",X"00",X"AA",
		X"3F",X"D0",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"3F",X"D0",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",
		X"3F",X"D0",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"57",X"D0",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"01",X"50",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"00",X"02",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"02",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"00",X"00",X"FF",X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"FF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",
		X"AA",X"00",X"00",X"FF",X"FF",X"FF",X"F0",X"00",X"AA",X"AA",X"00",X"00",X"FF",X"FF",X"F0",X"00",
		X"AA",X"AA",X"AA",X"00",X"00",X"FF",X"F0",X"00",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"F0",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"00",
		X"AA",X"0A",X"A0",X"CC",X"FF",X"FF",X"FF",X"FF",X"82",X"09",X"63",X"F3",X"FF",X"FF",X"FF",X"FF",
		X"82",X"A9",X"60",X"CC",X"FF",X"FF",X"FF",X"FF",X"82",X"09",X"63",X"33",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"0A",X"A0",X"CF",X"FF",X"FF",X"FF",X"FF",X"82",X"08",X"23",X"33",X"FF",X"FF",X"FF",X"FF",
		X"82",X"A8",X"20",X"CC",X"FF",X"FF",X"FF",X"FF",X"82",X"08",X"23",X"33",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"0A",X"A0",X"CC",X"FF",X"FF",X"FF",X"FF",X"96",X"09",X"63",X"3F",X"FF",X"FF",X"FF",X"FF",
		X"96",X"A9",X"60",X"CF",X"FF",X"FF",X"FF",X"FF",X"96",X"09",X"63",X"33",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"0A",X"A0",X"CC",X"FF",X"FF",X"FF",X"FF",X"82",X"08",X"23",X"3F",X"FF",X"FF",X"FF",X"FF",
		X"82",X"A8",X"20",X"CC",X"FF",X"FF",X"FF",X"FF",X"82",X"08",X"23",X"33",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FB",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FB",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FB",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FB",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FB",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FB",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FB",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FB",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"EF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"EF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"EF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"EF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"EF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"EF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"EF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"EF",
		X"2A",X"AA",X"00",X"00",X"00",X"00",X"AA",X"A8",X"20",X"96",X"00",X"00",X"00",X"00",X"82",X"58",
		X"20",X"96",X"00",X"00",X"00",X"00",X"82",X"58",X"20",X"96",X"00",X"00",X"00",X"00",X"82",X"58",
		X"20",X"AA",X"00",X"00",X"00",X"00",X"82",X"A8",X"2A",X"82",X"00",X"00",X"00",X"00",X"82",X"08",
		X"A5",X"82",X"00",X"00",X"00",X"00",X"AA",X"0A",X"25",X"82",X"00",X"00",X"00",X"00",X"82",X"08",
		X"25",X"AA",X"00",X"00",X"00",X"00",X"82",X"08",X"AA",X"82",X"00",X"00",X"00",X"00",X"82",X"0A",
		X"08",X"82",X"00",X"00",X"00",X"00",X"AA",X"20",X"02",X"82",X"00",X"00",X"00",X"00",X"96",X"80",
		X"AA",X"82",X"00",X"00",X"00",X"00",X"96",X"AA",X"20",X"22",X"00",X"00",X"00",X"00",X"98",X"08",
		X"20",X"0A",X"00",X"00",X"00",X"00",X"A8",X"08",X"AA",X"AA",X"00",X"00",X"00",X"00",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"00",X"02",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"02",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"02",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"02",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FF",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"FF",X"FF",X"FF",X"00",X"00",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"AA",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"AA",
		X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"FF",X"00",X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"03",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"02",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"02",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"00",X"02",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"02",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"00",X"02",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"02",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"02",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"02",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FF",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"00",
		X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"A0",X"00",X"AA",X"00",X"00",X"AA",X"AA",X"AA",X"A0",X"00",
		X"AA",X"AA",X"00",X"00",X"AA",X"AA",X"A0",X"00",X"AA",X"AA",X"AA",X"00",X"00",X"AA",X"A0",X"00",
		X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"A0",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"00",
		X"02",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"00",X"00",X"02",X"AA",X"AA",X"AA",X"AA",X"A0",X"00",
		X"AA",X"00",X"02",X"AA",X"AA",X"AA",X"A0",X"00",X"AA",X"AA",X"00",X"02",X"AA",X"AA",X"A0",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FC",X"CA",X"A0",X"AA",X"FF",X"FF",X"FF",X"FF",X"33",X"09",X"60",X"82",
		X"FF",X"FF",X"FF",X"FF",X"CC",X"C9",X"6A",X"82",X"FF",X"FF",X"FF",X"FF",X"F3",X"09",X"60",X"82",
		X"FF",X"FF",X"FF",X"FF",X"CC",X"CA",X"A0",X"AA",X"FF",X"FF",X"FF",X"FF",X"33",X"08",X"20",X"96",
		X"FF",X"FF",X"FF",X"FF",X"CC",X"C8",X"2A",X"96",X"FF",X"FF",X"FF",X"FF",X"33",X"08",X"20",X"96",
		X"FF",X"FF",X"FF",X"FF",X"FC",X"CA",X"A0",X"AA",X"FF",X"FF",X"FF",X"FF",X"33",X"08",X"20",X"82",
		X"FF",X"FF",X"FF",X"FF",X"CC",X"C8",X"2A",X"82",X"FF",X"FF",X"FF",X"FF",X"33",X"08",X"25",X"82",
		X"FF",X"FF",X"FF",X"FF",X"CC",X"CA",X"A5",X"AA",X"FF",X"FF",X"FF",X"FF",X"33",X"08",X"25",X"82",
		X"FF",X"FF",X"FF",X"FF",X"FC",X"C8",X"2A",X"82",X"FF",X"FF",X"FF",X"FF",X"33",X"08",X"20",X"82",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"CC",X"C0",X"CC",X"C0",X"CC",X"CC",X"CC",X"CC",X"33",X"33",X"33",X"33",X"33",X"30",X"33",X"33",
		X"0C",X"CC",X"CC",X"CC",X"CC",X"CC",X"C0",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"25",X"60",X"20",X"08",X"08",X"09",X"58",X"08",
		X"25",X"60",X"20",X"08",X"08",X"09",X"58",X"08",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"02",X"02",X"00",X"95",X"80",X"95",X"80",X"80",X"02",X"02",X"00",X"95",X"80",X"95",X"80",X"80",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"20",X"25",X"60",X"08",X"08",X"08",X"09",X"58",
		X"20",X"25",X"60",X"08",X"08",X"08",X"09",X"58",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FB",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FB",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FB",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FB",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FB",X"AB",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FE",X"AE",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FB",X"BA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FE",X"EA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"FE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"EF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"EF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"EF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"EF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"EA",X"BF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"BA",X"EF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AE",X"BF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AB",X"EF",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BF",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"00",X"89",X"58",X"08",X"0A",
		X"00",X"00",X"00",X"00",X"89",X"58",X"08",X"26",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"96",
		X"00",X"00",X"00",X"00",X"95",X"80",X"96",X"96",X"00",X"00",X"00",X"00",X"95",X"80",X"98",X"96",
		X"00",X"00",X"00",X"00",X"AA",X"AA",X"A0",X"AA",X"00",X"00",X"00",X"00",X"88",X"08",X"A0",X"82",
		X"00",X"00",X"00",X"00",X"88",X"0A",X"20",X"82",X"00",X"00",X"00",X"00",X"AA",X"A8",X"2A",X"82",
		X"00",X"00",X"00",X"00",X"00",X"08",X"25",X"82",X"00",X"00",X"00",X"00",X"00",X"08",X"25",X"82",
		X"00",X"00",X"00",X"00",X"30",X"CA",X"A5",X"AA",X"00",X"00",X"00",X"00",X"00",X"08",X"25",X"82",
		X"00",X"00",X"00",X"00",X"30",X"08",X"2A",X"82",X"00",X"00",X"00",X"00",X"00",X"08",X"20",X"82",
		X"82",X"A8",X"20",X"00",X"00",X"00",X"00",X"00",X"82",X"08",X"2C",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"0A",X"A0",X"00",X"C0",X"00",X"00",X"0C",X"82",X"08",X"20",X"00",X"00",X"00",X"00",X"00",
		X"82",X"A8",X"20",X"00",X"00",X"0C",X"00",X"00",X"82",X"08",X"20",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"08",X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",X"96",X"08",X"88",X"08",X"09",X"56",X"02",X"02",
		X"96",X"AA",X"08",X"08",X"09",X"56",X"02",X"02",X"96",X"0A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"20",X"95",X"80",X"80",X"80",X"25",X"60",X"82",X"80",X"95",X"80",X"80",X"80",X"25",X"60",
		X"82",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"89",X"58",X"08",X"08",X"09",X"56",X"02",X"02",
		X"A5",X"58",X"08",X"08",X"09",X"56",X"02",X"02",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"08",X"2A",X"82",X"30",X"30",X"00",X"00",X"30",X"08",X"20",X"82",
		X"00",X"00",X"00",X"00",X"00",X"CA",X"A0",X"AA",X"00",X"03",X"00",X"30",X"00",X"08",X"20",X"96",
		X"00",X"C0",X"00",X"00",X"0C",X"08",X"2A",X"96",X"00",X"00",X"00",X"00",X"00",X"08",X"25",X"96",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"25",X"AA",X"02",X"02",X"56",X"02",X"56",X"02",X"25",X"82",
		X"02",X"02",X"56",X"02",X"56",X"00",X"A5",X"82",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A5",X"82",
		X"20",X"25",X"60",X"20",X"20",X"20",X"09",X"AA",X"20",X"25",X"60",X"20",X"20",X"20",X"02",X"82",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"82",X"02",X"02",X"02",X"02",X"02",X"56",X"00",X"22",
		X"02",X"02",X"02",X"02",X"02",X"56",X"00",X"0A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"0A",X"A3",X"00",X"00",X"00",X"00",X"00",X"82",X"09",X"60",X"00",X"00",X"00",X"00",X"00",
		X"82",X"A9",X"60",X"00",X"00",X"00",X"00",X"00",X"82",X"09",X"60",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"0A",X"A3",X"0F",X"00",X"00",X"00",X"00",X"96",X"08",X"20",X"00",X"00",X"00",X"00",X"00",
		X"96",X"A8",X"20",X"30",X"00",X"00",X"00",X"00",X"96",X"08",X"20",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"0A",X"A0",X"00",X"00",X"00",X"00",X"00",X"82",X"08",X"20",X"00",X"00",X"00",X"00",X"00",
		X"82",X"A8",X"20",X"C0",X"00",X"00",X"00",X"00",X"82",X"58",X"20",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"5A",X"A0",X"0C",X"00",X"00",X"00",X"00",X"82",X"58",X"20",X"00",X"00",X"00",X"00",X"00",
		X"82",X"A8",X"23",X"00",X"00",X"00",X"00",X"00",X"82",X"08",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"0A",X"A0",X"AA",X"00",X"00",X"00",X"00",X"00",X"09",X"60",X"82",
		X"00",X"00",X"00",X"00",X"30",X"09",X"6A",X"82",X"00",X"00",X"00",X"00",X"03",X"09",X"60",X"82",
		X"00",X"00",X"00",X"00",X"00",X"0A",X"A0",X"AA",X"00",X"00",X"00",X"00",X"00",X"08",X"20",X"96",
		X"00",X"00",X"00",X"00",X"00",X"C8",X"2A",X"96",X"00",X"00",X"00",X"00",X"00",X"C8",X"25",X"96",
		X"00",X"00",X"00",X"00",X"00",X"0A",X"A5",X"AA",X"00",X"00",X"00",X"00",X"00",X"08",X"25",X"82",
		X"00",X"00",X"00",X"00",X"03",X"08",X"2A",X"82",X"00",X"00",X"00",X"00",X"00",X"08",X"20",X"82",
		X"00",X"00",X"00",X"00",X"0C",X"0A",X"A0",X"AA",X"00",X"00",X"00",X"00",X"00",X"09",X"60",X"82",
		X"00",X"00",X"00",X"00",X"00",X"09",X"6A",X"82",X"00",X"00",X"00",X"00",X"00",X"09",X"60",X"82",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"00",X"30",X"00",X"00",X"C0",X"00",X"30",X"00",X"00",X"00",X"30",X"C0",X"00",
		X"30",X"00",X"F0",X"00",X"C0",X"30",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"20",X"20",X"20",X"09",X"58",X"09",X"58",X"08",
		X"20",X"20",X"20",X"09",X"58",X"09",X"58",X"08",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"02",X"56",X"00",X"80",X"80",X"80",X"80",X"80",X"02",X"56",X"00",X"80",X"80",X"80",X"80",X"80",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"20",X"20",X"25",X"58",X"09",X"58",X"09",X"58",
		X"20",X"20",X"25",X"58",X"09",X"58",X"09",X"58",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
