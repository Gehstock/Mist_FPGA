library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity cpu2_rom is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of cpu2_rom is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"31",X"80",X"8B",X"C3",X"85",X"00",X"FF",X"FF",X"87",X"30",X"05",X"24",X"18",X"02",X"FF",X"FF",
		X"85",X"6F",X"D0",X"24",X"C9",X"FF",X"FF",X"FF",X"77",X"23",X"10",X"FC",X"C9",X"FF",X"FF",X"FF",
		X"CF",X"7E",X"23",X"66",X"6F",X"E9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F5",X"E5",X"3A",X"3C",X"9B",X"A7",X"28",X"08",X"AF",X"32",
		X"3C",X"9B",X"E1",X"F1",X"ED",X"45",X"3E",X"01",X"32",X"3C",X"9B",X"32",X"22",X"68",X"AF",X"32",
		X"22",X"68",X"C3",X"B5",X"00",X"3E",X"01",X"32",X"22",X"68",X"CD",X"7F",X"06",X"21",X"40",X"8A",
		X"06",X"08",X"AF",X"DF",X"21",X"80",X"9A",X"36",X"00",X"11",X"81",X"9A",X"01",X"FF",X"00",X"ED",
		X"B0",X"21",X"E7",X"07",X"11",X"0A",X"9B",X"01",X"15",X"00",X"ED",X"B0",X"AF",X"32",X"22",X"68",
		X"31",X"80",X"8B",X"18",X"FB",X"21",X"20",X"9B",X"36",X"00",X"11",X"21",X"9B",X"01",X"0F",X"00",
		X"ED",X"B0",X"3A",X"57",X"86",X"CB",X"4F",X"28",X"3F",X"3A",X"CF",X"87",X"CB",X"67",X"28",X"10",
		X"21",X"80",X"9A",X"36",X"00",X"11",X"81",X"9A",X"01",X"27",X"00",X"ED",X"B0",X"C3",X"F5",X"02",
		X"AF",X"21",X"80",X"9A",X"06",X"0A",X"DF",X"21",X"96",X"9A",X"06",X"0A",X"DF",X"32",X"8E",X"9A",
		X"32",X"A4",X"9A",X"21",X"90",X"9A",X"06",X"03",X"DF",X"21",X"A6",X"9A",X"06",X"03",X"DF",X"32",
		X"94",X"9A",X"32",X"AA",X"9A",X"C3",X"D0",X"01",X"3A",X"33",X"9B",X"A7",X"28",X"09",X"21",X"80",
		X"9A",X"86",X"77",X"AF",X"32",X"33",X"9B",X"3A",X"81",X"9A",X"A7",X"28",X"0B",X"21",X"34",X"9B",
		X"36",X"01",X"CD",X"91",X"03",X"C3",X"E7",X"02",X"3A",X"88",X"9A",X"A7",X"28",X"0B",X"21",X"34",
		X"9B",X"36",X"08",X"CD",X"91",X"03",X"C3",X"E7",X"02",X"3A",X"82",X"9A",X"A7",X"28",X"0B",X"21",
		X"34",X"9B",X"36",X"02",X"CD",X"91",X"03",X"C3",X"E7",X"02",X"3A",X"83",X"9A",X"A7",X"28",X"0B",
		X"21",X"34",X"9B",X"36",X"03",X"CD",X"91",X"03",X"C3",X"E7",X"02",X"3A",X"94",X"9A",X"A7",X"28",
		X"0B",X"21",X"34",X"9B",X"36",X"14",X"CD",X"91",X"03",X"C3",X"E7",X"02",X"3A",X"87",X"9A",X"A7",
		X"28",X"0B",X"21",X"34",X"9B",X"36",X"07",X"CD",X"91",X"03",X"C3",X"E7",X"02",X"3A",X"84",X"9A",
		X"A7",X"28",X"0B",X"21",X"34",X"9B",X"36",X"04",X"CD",X"91",X"03",X"C3",X"E7",X"02",X"3A",X"85",
		X"9A",X"A7",X"28",X"0B",X"21",X"34",X"9B",X"36",X"05",X"CD",X"91",X"03",X"C3",X"E7",X"02",X"3A",
		X"91",X"9A",X"A7",X"28",X"10",X"21",X"34",X"9B",X"36",X"11",X"CD",X"91",X"03",X"3E",X"50",X"32",
		X"3B",X"9B",X"C3",X"D0",X"01",X"3A",X"3B",X"9B",X"3D",X"32",X"3B",X"9B",X"20",X"12",X"21",X"3B",
		X"9B",X"34",X"3A",X"92",X"9A",X"A7",X"28",X"08",X"21",X"34",X"9B",X"36",X"12",X"CD",X"91",X"03",
		X"21",X"34",X"9B",X"36",X"0F",X"3A",X"8F",X"9A",X"A7",X"28",X"0A",X"AF",X"32",X"8F",X"9A",X"CD",
		X"1A",X"03",X"C3",X"0F",X"02",X"3A",X"A5",X"9A",X"A7",X"28",X"06",X"CD",X"4E",X"03",X"C3",X"0F",
		X"02",X"21",X"34",X"9B",X"36",X"10",X"3A",X"90",X"9A",X"A7",X"28",X"0A",X"AF",X"32",X"90",X"9A",
		X"CD",X"1A",X"03",X"C3",X"0F",X"02",X"3A",X"A6",X"9A",X"A7",X"28",X"03",X"CD",X"4E",X"03",X"21",
		X"34",X"9B",X"36",X"0A",X"3A",X"8A",X"9A",X"A7",X"28",X"09",X"AF",X"32",X"8A",X"9A",X"CD",X"1A",
		X"03",X"18",X"3B",X"3A",X"A0",X"9A",X"A7",X"28",X"05",X"CD",X"4E",X"03",X"18",X"30",X"3A",X"8B",
		X"9A",X"A7",X"28",X"0B",X"21",X"34",X"9B",X"36",X"0B",X"CD",X"91",X"03",X"C3",X"5E",X"02",X"3A",
		X"8C",X"9A",X"A7",X"28",X"0B",X"21",X"34",X"9B",X"36",X"0C",X"CD",X"91",X"03",X"C3",X"5E",X"02",
		X"3A",X"8D",X"9A",X"A7",X"28",X"08",X"21",X"34",X"9B",X"36",X"0D",X"CD",X"91",X"03",X"21",X"34",
		X"9B",X"36",X"0E",X"3A",X"8E",X"9A",X"A7",X"28",X"09",X"AF",X"32",X"8E",X"9A",X"CD",X"1A",X"03",
		X"18",X"09",X"3A",X"A4",X"9A",X"A7",X"28",X"03",X"CD",X"4E",X"03",X"3A",X"89",X"9A",X"A7",X"28",
		X"1B",X"21",X"46",X"86",X"CB",X"46",X"28",X"09",X"AF",X"32",X"89",X"9A",X"32",X"9F",X"9A",X"18",
		X"0B",X"21",X"34",X"9B",X"36",X"09",X"CD",X"91",X"03",X"C3",X"C1",X"02",X"3A",X"86",X"9A",X"A7",
		X"28",X"1F",X"21",X"46",X"86",X"CB",X"46",X"20",X"07",X"21",X"01",X"84",X"CB",X"7E",X"28",X"09",
		X"AF",X"32",X"86",X"9A",X"32",X"9C",X"9A",X"18",X"08",X"21",X"34",X"9B",X"36",X"06",X"CD",X"91",
		X"03",X"3A",X"93",X"9A",X"A7",X"28",X"20",X"3A",X"57",X"86",X"CB",X"4F",X"C2",X"DF",X"02",X"21",
		X"01",X"84",X"CB",X"6E",X"20",X"09",X"AF",X"32",X"93",X"9A",X"32",X"A9",X"9A",X"18",X"08",X"21",
		X"34",X"9B",X"36",X"13",X"CD",X"91",X"03",X"3A",X"80",X"9A",X"A7",X"28",X"08",X"21",X"34",X"9B",
		X"36",X"00",X"CD",X"91",X"03",X"21",X"20",X"9B",X"11",X"10",X"68",X"01",X"10",X"00",X"ED",X"B0",
		X"3A",X"30",X"9B",X"32",X"05",X"68",X"3A",X"31",X"9B",X"32",X"0A",X"68",X"3A",X"32",X"9B",X"32",
		X"0F",X"68",X"AF",X"32",X"3C",X"9B",X"E1",X"F1",X"ED",X"45",X"21",X"96",X"9A",X"3A",X"34",X"9B",
		X"D7",X"34",X"21",X"34",X"9B",X"7E",X"87",X"86",X"21",X"54",X"07",X"D7",X"11",X"35",X"9B",X"01",
		X"03",X"00",X"ED",X"B0",X"21",X"36",X"9B",X"46",X"48",X"21",X"DB",X"9A",X"3A",X"35",X"9B",X"D7",
		X"AF",X"DF",X"41",X"21",X"AC",X"9A",X"3A",X"35",X"9B",X"D7",X"AF",X"DF",X"18",X"12",X"21",X"34",
		X"9B",X"7E",X"87",X"86",X"21",X"54",X"07",X"D7",X"11",X"35",X"9B",X"01",X"03",X"00",X"ED",X"B0",
		X"CD",X"D5",X"04",X"21",X"36",X"9B",X"35",X"28",X"0A",X"21",X"35",X"9B",X"34",X"21",X"37",X"9B",
		X"34",X"18",X"ED",X"3A",X"38",X"9B",X"A7",X"C8",X"AF",X"32",X"38",X"9B",X"21",X"96",X"9A",X"3A",
		X"34",X"9B",X"D7",X"36",X"00",X"21",X"0D",X"04",X"3A",X"34",X"9B",X"CF",X"5E",X"23",X"56",X"EB",
		X"E9",X"21",X"34",X"9B",X"7E",X"87",X"86",X"21",X"54",X"07",X"D7",X"11",X"35",X"9B",X"01",X"03",
		X"00",X"ED",X"B0",X"21",X"96",X"9A",X"3A",X"34",X"9B",X"D7",X"7E",X"A7",X"20",X"19",X"34",X"21",
		X"36",X"9B",X"46",X"48",X"21",X"DB",X"9A",X"3A",X"35",X"9B",X"D7",X"AF",X"DF",X"41",X"21",X"AC",
		X"9A",X"3A",X"35",X"9B",X"D7",X"AF",X"DF",X"CD",X"D5",X"04",X"21",X"36",X"9B",X"35",X"28",X"0A",
		X"21",X"35",X"9B",X"34",X"21",X"37",X"9B",X"34",X"18",X"ED",X"3A",X"38",X"9B",X"A7",X"C8",X"AF",
		X"32",X"38",X"9B",X"21",X"96",X"9A",X"3A",X"34",X"9B",X"D7",X"36",X"00",X"21",X"80",X"9A",X"3A",
		X"34",X"9B",X"D7",X"3A",X"34",X"9B",X"A7",X"28",X"12",X"FE",X"14",X"28",X"0E",X"36",X"00",X"21",
		X"0D",X"04",X"3A",X"34",X"9B",X"CF",X"5E",X"23",X"56",X"EB",X"E9",X"35",X"C9",X"37",X"04",X"38",
		X"04",X"37",X"04",X"37",X"04",X"C6",X"04",X"48",X"04",X"5F",X"04",X"6E",X"04",X"48",X"04",X"63",
		X"04",X"37",X"04",X"37",X"04",X"40",X"04",X"37",X"04",X"90",X"04",X"37",X"04",X"37",X"04",X"37",
		X"04",X"37",X"04",X"AB",X"04",X"37",X"04",X"C9",X"AF",X"32",X"94",X"9A",X"32",X"AA",X"9A",X"C9",
		X"AF",X"32",X"8D",X"9A",X"32",X"A3",X"9A",X"C9",X"AF",X"32",X"86",X"9A",X"32",X"89",X"9A",X"32",
		X"9C",X"9A",X"32",X"9F",X"9A",X"32",X"93",X"9A",X"32",X"A9",X"9A",X"3E",X"10",X"18",X"06",X"3E",
		X"0A",X"18",X"02",X"3E",X"0C",X"32",X"1B",X"9B",X"AF",X"32",X"A7",X"9A",X"18",X"07",X"AF",X"32",
		X"93",X"9A",X"32",X"A9",X"9A",X"21",X"8A",X"9A",X"11",X"8B",X"9A",X"01",X"08",X"00",X"36",X"00",
		X"ED",X"B0",X"21",X"A0",X"9A",X"11",X"A1",X"9A",X"01",X"08",X"00",X"36",X"00",X"ED",X"B0",X"C9",
		X"21",X"8A",X"9A",X"11",X"8B",X"9A",X"01",X"03",X"00",X"36",X"00",X"ED",X"B0",X"21",X"A0",X"9A",
		X"11",X"A1",X"9A",X"01",X"03",X"00",X"36",X"00",X"ED",X"B0",X"C9",X"21",X"8A",X"9A",X"11",X"8B",
		X"9A",X"01",X"06",X"00",X"36",X"00",X"ED",X"B0",X"21",X"A0",X"9A",X"11",X"A1",X"9A",X"01",X"06",
		X"00",X"36",X"00",X"ED",X"B0",X"C9",X"AF",X"32",X"86",X"9A",X"32",X"89",X"9A",X"32",X"9C",X"9A",
		X"32",X"9F",X"9A",X"18",X"99",X"21",X"AC",X"9A",X"3A",X"35",X"9B",X"D7",X"34",X"3A",X"35",X"9B",
		X"21",X"00",X"07",X"CF",X"5E",X"23",X"56",X"21",X"DB",X"9A",X"3A",X"35",X"9B",X"D7",X"7E",X"EB",
		X"D7",X"22",X"39",X"9B",X"7E",X"3C",X"CA",X"13",X"06",X"21",X"BD",X"07",X"3A",X"35",X"9B",X"D7",
		X"7E",X"A7",X"28",X"0D",X"3D",X"28",X"05",X"11",X"65",X"06",X"18",X"08",X"11",X"4B",X"06",X"18",
		X"03",X"11",X"31",X"06",X"2A",X"39",X"9B",X"7E",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"EB",X"CF",
		X"4E",X"23",X"46",X"EB",X"7E",X"E6",X"0F",X"28",X"07",X"CB",X"38",X"CB",X"19",X"3D",X"20",X"F9",
		X"3A",X"37",X"9B",X"A7",X"28",X"0D",X"3D",X"28",X"05",X"21",X"2B",X"9B",X"18",X"08",X"21",X"26",
		X"9B",X"18",X"03",X"21",X"21",X"9B",X"71",X"7E",X"0F",X"0F",X"0F",X"0F",X"23",X"77",X"23",X"70",
		X"7E",X"0F",X"0F",X"0F",X"0F",X"23",X"77",X"3A",X"37",X"9B",X"A7",X"28",X"0D",X"3D",X"28",X"05",
		X"11",X"2F",X"9B",X"18",X"08",X"11",X"2A",X"9B",X"18",X"03",X"11",X"25",X"9B",X"2A",X"39",X"9B",
		X"7E",X"D6",X"C0",X"28",X"4A",X"3A",X"35",X"9B",X"21",X"FC",X"07",X"D7",X"A7",X"28",X"21",X"3D",
		X"28",X"0F",X"21",X"AC",X"9A",X"3A",X"35",X"9B",X"D7",X"7E",X"FE",X"06",X"30",X"12",X"2F",X"18",
		X"33",X"21",X"AC",X"9A",X"3A",X"35",X"9B",X"D7",X"7E",X"FE",X"06",X"30",X"03",X"87",X"18",X"24",
		X"21",X"26",X"08",X"3A",X"35",X"9B",X"D7",X"7E",X"A7",X"28",X"17",X"47",X"21",X"AC",X"9A",X"3A",
		X"35",X"9B",X"D7",X"7E",X"90",X"38",X"0B",X"D6",X"0A",X"30",X"04",X"ED",X"44",X"18",X"05",X"AF",
		X"18",X"02",X"3E",X"0A",X"12",X"21",X"30",X"9B",X"3A",X"37",X"9B",X"D7",X"EB",X"21",X"93",X"07",
		X"3A",X"35",X"9B",X"D7",X"ED",X"A0",X"21",X"0A",X"9B",X"3A",X"34",X"9B",X"D7",X"7E",X"2A",X"39",
		X"9B",X"23",X"5E",X"16",X"00",X"21",X"00",X"00",X"06",X"08",X"CB",X"3F",X"30",X"01",X"19",X"CB",
		X"23",X"CB",X"12",X"10",X"F5",X"45",X"21",X"AC",X"9A",X"3A",X"35",X"9B",X"D7",X"78",X"BE",X"C0",
		X"21",X"DB",X"9A",X"3A",X"35",X"9B",X"D7",X"34",X"34",X"21",X"AC",X"9A",X"3A",X"35",X"9B",X"D7",
		X"36",X"00",X"C9",X"3A",X"37",X"9B",X"A7",X"28",X"0D",X"3D",X"28",X"05",X"21",X"2F",X"9B",X"18",
		X"08",X"21",X"2A",X"9B",X"18",X"03",X"21",X"25",X"9B",X"36",X"00",X"3E",X"01",X"32",X"38",X"9B",
		X"C9",X"50",X"81",X"00",X"89",X"26",X"91",X"C8",X"99",X"EC",X"A2",X"9D",X"AC",X"E0",X"B6",X"C0",
		X"C1",X"45",X"CD",X"7A",X"D9",X"69",X"E6",X"1C",X"F4",X"00",X"00",X"35",X"82",X"F2",X"89",X"27",
		X"92",X"D8",X"9A",X"0C",X"A4",X"CE",X"AD",X"23",X"B8",X"17",X"C3",X"B0",X"CE",X"FB",X"DA",X"01",
		X"E8",X"CC",X"F5",X"00",X"00",X"6E",X"80",X"11",X"88",X"29",X"90",X"BC",X"98",X"D0",X"A1",X"70",
		X"AB",X"A1",X"B5",X"6E",X"C0",X"DF",X"CB",X"FE",X"D7",X"D7",X"E4",X"72",X"F2",X"00",X"00",X"21",
		X"00",X"00",X"06",X"10",X"AF",X"86",X"2C",X"20",X"FC",X"24",X"10",X"F9",X"FE",X"AA",X"20",X"0C",
		X"3E",X"FF",X"32",X"01",X"8A",X"3A",X"01",X"8A",X"A7",X"20",X"FA",X"C9",X"3E",X"06",X"32",X"01",
		X"8A",X"18",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"50",X"08",X"9F",X"08",X"EE",X"08",X"31",X"09",X"31",X"09",X"4E",X"09",X"67",X"09",X"DC",X"09",
		X"51",X"0A",X"B2",X"0A",X"B2",X"0A",X"C9",X"0A",X"E2",X"0A",X"09",X"0B",X"36",X"0B",X"57",X"0B",
		X"62",X"0B",X"6D",X"0B",X"8E",X"0B",X"E5",X"0B",X"66",X"0C",X"77",X"0C",X"90",X"0C",X"90",X"0C",
		X"90",X"0C",X"A3",X"0C",X"BA",X"0C",X"E3",X"0C",X"0C",X"0D",X"35",X"0D",X"66",X"0D",X"73",X"0D",
		X"8C",X"0D",X"A5",X"0D",X"BE",X"0D",X"D7",X"0D",X"E2",X"0D",X"ED",X"0D",X"F8",X"0D",X"09",X"0E",
		X"62",X"0E",X"BB",X"0E",X"14",X"01",X"02",X"00",X"03",X"00",X"06",X"03",X"00",X"09",X"03",X"00",
		X"23",X"03",X"00",X"1A",X"03",X"00",X"21",X"02",X"00",X"16",X"03",X"00",X"03",X"03",X"00",X"1F",
		X"02",X"00",X"0D",X"01",X"02",X"19",X"01",X"02",X"11",X"01",X"02",X"0F",X"02",X"01",X"1D",X"02",
		X"01",X"15",X"01",X"00",X"0C",X"01",X"00",X"12",X"02",X"00",X"0E",X"01",X"01",X"26",X"01",X"00",
		X"27",X"03",X"00",X"02",X"00",X"05",X"03",X"00",X"04",X"02",X"00",X"05",X"05",X"02",X"04",X"05",
		X"04",X"06",X"02",X"01",X"02",X"03",X"04",X"03",X"03",X"00",X"01",X"05",X"02",X"02",X"02",X"02",
		X"00",X"01",X"05",X"05",X"02",X"04",X"02",X"02",X"02",X"02",X"02",X"00",X"05",X"00",X"01",X"00",
		X"00",X"01",X"00",X"00",X"01",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",
		X"01",X"00",X"00",X"00",X"01",X"02",X"00",X"00",X"01",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"02",X"00",X"00",X"00",X"00",X"08",X"10",X"0C",X"0C",X"08",X"06",X"10",X"0E",X"0C",
		X"10",X"02",X"04",X"02",X"04",X"02",X"04",X"02",X"10",X"04",X"08",X"0C",X"00",X"01",X"02",X"00",
		X"01",X"00",X"00",X"01",X"02",X"00",X"01",X"00",X"00",X"00",X"00",X"02",X"01",X"00",X"02",X"02",
		X"02",X"02",X"01",X"00",X"02",X"00",X"01",X"01",X"01",X"02",X"01",X"02",X"01",X"02",X"01",X"02",
		X"02",X"02",X"02",X"00",X"00",X"02",X"01",X"00",X"04",X"01",X"01",X"06",X"03",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"03",X"00",X"00",X"00",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"06",X"04",X"06",X"00",X"00",X"00",X"00",X"01",X"06",X"00",
		X"05",X"01",X"15",X"01",X"15",X"01",X"15",X"01",X"06",X"01",X"16",X"01",X"16",X"01",X"16",X"01",
		X"07",X"01",X"17",X"01",X"17",X"01",X"17",X"01",X"C0",X"01",X"15",X"01",X"15",X"01",X"15",X"01",
		X"15",X"01",X"C0",X"01",X"A6",X"01",X"C0",X"01",X"15",X"01",X"A6",X"02",X"15",X"01",X"35",X"01",
		X"A6",X"01",X"A6",X"01",X"A6",X"02",X"86",X"01",X"66",X"02",X"76",X"01",X"C0",X"01",X"16",X"01",
		X"C0",X"01",X"76",X"01",X"16",X"02",X"76",X"02",X"86",X"01",X"86",X"01",X"86",X"05",X"FF",X"06",
		X"01",X"16",X"01",X"16",X"01",X"16",X"01",X"07",X"01",X"17",X"01",X"17",X"01",X"17",X"01",X"08",
		X"01",X"18",X"01",X"18",X"01",X"18",X"01",X"C0",X"01",X"16",X"01",X"16",X"01",X"16",X"01",X"16",
		X"01",X"C0",X"01",X"A7",X"01",X"C0",X"01",X"16",X"01",X"A7",X"02",X"16",X"01",X"36",X"01",X"A7",
		X"01",X"A7",X"01",X"A7",X"02",X"87",X"01",X"67",X"02",X"77",X"01",X"C0",X"01",X"17",X"01",X"C0",
		X"01",X"77",X"01",X"17",X"02",X"77",X"02",X"87",X"01",X"87",X"01",X"87",X"05",X"FF",X"C0",X"0C",
		X"C0",X"01",X"18",X"01",X"38",X"01",X"58",X"01",X"68",X"01",X"18",X"01",X"68",X"01",X"18",X"01",
		X"68",X"01",X"18",X"01",X"68",X"01",X"18",X"01",X"68",X"01",X"18",X"01",X"68",X"01",X"18",X"01",
		X"68",X"01",X"18",X"01",X"68",X"01",X"18",X"01",X"48",X"01",X"18",X"01",X"48",X"01",X"18",X"01",
		X"48",X"01",X"18",X"01",X"48",X"01",X"18",X"01",X"58",X"01",X"18",X"01",X"58",X"01",X"18",X"05",
		X"FF",X"A6",X"01",X"B6",X"01",X"05",X"01",X"15",X"02",X"A6",X"01",X"B6",X"02",X"86",X"01",X"A6",
		X"02",X"66",X"01",X"86",X"02",X"56",X"01",X"66",X"03",X"65",X"02",X"66",X"04",X"FF",X"C0",X"03",
		X"18",X"02",X"C0",X"01",X"28",X"02",X"C0",X"01",X"38",X"02",X"C0",X"01",X"58",X"02",X"C0",X"01",
		X"68",X"04",X"C0",X"01",X"68",X"04",X"FF",X"A6",X"02",X"B6",X"01",X"15",X"02",X"A6",X"01",X"86",
		X"02",X"66",X"03",X"86",X"01",X"A6",X"02",X"36",X"01",X"16",X"02",X"C0",X"01",X"16",X"01",X"C0",
		X"01",X"16",X"04",X"A6",X"02",X"B6",X"01",X"15",X"02",X"A6",X"01",X"86",X"02",X"66",X"03",X"86",
		X"01",X"A6",X"02",X"16",X"01",X"36",X"02",X"C0",X"01",X"36",X"01",X"C0",X"01",X"36",X"04",X"B6",
		X"02",X"15",X"01",X"35",X"02",X"B6",X"01",X"A6",X"02",X"86",X"02",X"C0",X"01",X"86",X"01",X"A6",
		X"02",X"B6",X"01",X"15",X"02",X"A6",X"01",X"86",X"02",X"66",X"02",X"C0",X"01",X"66",X"01",X"86",
		X"02",X"A6",X"01",X"B6",X"02",X"86",X"01",X"66",X"02",X"56",X"03",X"36",X"01",X"56",X"02",X"16",
		X"01",X"66",X"02",X"C0",X"01",X"66",X"01",X"C0",X"01",X"66",X"04",X"FF",X"A7",X"02",X"B7",X"01",
		X"16",X"02",X"A7",X"01",X"87",X"02",X"67",X"03",X"87",X"01",X"A7",X"02",X"37",X"01",X"17",X"02",
		X"C0",X"01",X"17",X"01",X"C0",X"01",X"17",X"04",X"A7",X"02",X"B7",X"01",X"16",X"02",X"A7",X"01",
		X"87",X"02",X"67",X"03",X"87",X"01",X"A7",X"02",X"17",X"01",X"37",X"02",X"C0",X"01",X"37",X"01",
		X"C0",X"01",X"37",X"04",X"B7",X"02",X"16",X"01",X"36",X"02",X"B7",X"01",X"A7",X"02",X"87",X"02",
		X"C0",X"01",X"87",X"01",X"A7",X"02",X"B7",X"01",X"16",X"02",X"A7",X"01",X"87",X"02",X"67",X"02",
		X"C0",X"01",X"67",X"01",X"87",X"02",X"A7",X"01",X"B7",X"02",X"87",X"01",X"67",X"02",X"57",X"03",
		X"37",X"01",X"57",X"02",X"17",X"01",X"67",X"02",X"C0",X"01",X"67",X"01",X"C0",X"01",X"67",X"04",
		X"FF",X"C0",X"03",X"69",X"04",X"C0",X"01",X"69",X"03",X"C0",X"01",X"69",X"02",X"C0",X"01",X"69",
		X"04",X"C0",X"01",X"69",X"03",X"C0",X"01",X"69",X"02",X"C0",X"01",X"69",X"04",X"C0",X"01",X"89",
		X"03",X"C0",X"01",X"A9",X"02",X"C0",X"01",X"B9",X"04",X"C0",X"01",X"B9",X"03",X"C0",X"01",X"A9",
		X"02",X"C0",X"01",X"89",X"04",X"C0",X"01",X"A9",X"03",X"C0",X"01",X"B9",X"02",X"C0",X"01",X"A9",
		X"04",X"C0",X"01",X"89",X"03",X"C0",X"01",X"69",X"02",X"C0",X"01",X"89",X"04",X"C0",X"01",X"19",
		X"03",X"C0",X"01",X"B9",X"02",X"C0",X"01",X"A9",X"02",X"C0",X"01",X"89",X"01",X"C0",X"01",X"69",
		X"04",X"FF",X"B7",X"01",X"06",X"01",X"16",X"01",X"26",X"02",X"36",X"01",X"46",X"02",X"56",X"03",
		X"16",X"01",X"66",X"03",X"16",X"02",X"66",X"07",X"FF",X"67",X"02",X"C0",X"01",X"57",X"02",X"C0",
		X"01",X"47",X"02",X"C0",X"01",X"37",X"02",X"C0",X"01",X"27",X"02",X"C0",X"01",X"17",X"02",X"68",
		X"07",X"FF",X"05",X"01",X"55",X"01",X"15",X"01",X"65",X"01",X"25",X"01",X"75",X"01",X"35",X"01",
		X"85",X"01",X"45",X"01",X"95",X"01",X"55",X"01",X"A5",X"01",X"65",X"01",X"B5",X"01",X"B7",X"02",
		X"A7",X"02",X"97",X"02",X"87",X"02",X"C0",X"02",X"FF",X"08",X"01",X"38",X"01",X"28",X"01",X"58",
		X"01",X"48",X"01",X"78",X"01",X"68",X"01",X"96",X"01",X"88",X"01",X"B8",X"01",X"A8",X"01",X"17",
		X"01",X"07",X"01",X"37",X"01",X"27",X"01",X"57",X"01",X"47",X"01",X"77",X"01",X"67",X"01",X"97",
		X"01",X"87",X"01",X"B7",X"01",X"FF",X"05",X"01",X"15",X"01",X"05",X"01",X"B6",X"01",X"05",X"01",
		X"15",X"01",X"05",X"01",X"B6",X"01",X"06",X"01",X"16",X"01",X"06",X"01",X"B7",X"01",X"06",X"01",
		X"16",X"01",X"06",X"01",X"B7",X"01",X"FF",X"16",X"04",X"B5",X"01",X"55",X"01",X"A5",X"01",X"65",
		X"01",X"FF",X"09",X"01",X"18",X"01",X"27",X"01",X"36",X"01",X"45",X"04",X"FF",X"08",X"01",X"B9",
		X"01",X"08",X"01",X"18",X"01",X"08",X"01",X"B9",X"01",X"08",X"01",X"18",X"01",X"58",X"01",X"48",
		X"01",X"58",X"01",X"68",X"01",X"58",X"01",X"48",X"01",X"58",X"01",X"68",X"01",X"FF",X"06",X"01",
		X"16",X"01",X"16",X"01",X"16",X"02",X"16",X"01",X"16",X"01",X"16",X"01",X"16",X"01",X"16",X"01",
		X"16",X"01",X"16",X"02",X"16",X"01",X"16",X"01",X"16",X"01",X"A7",X"02",X"87",X"01",X"A7",X"02",
		X"87",X"01",X"A7",X"01",X"87",X"01",X"A7",X"04",X"87",X"04",X"97",X"01",X"A7",X"01",X"A7",X"01",
		X"A7",X"02",X"A7",X"01",X"A7",X"01",X"A7",X"01",X"A7",X"01",X"A7",X"01",X"A7",X"01",X"A7",X"02",
		X"A7",X"01",X"A7",X"01",X"A7",X"01",X"A7",X"02",X"87",X"01",X"A7",X"02",X"87",X"01",X"A7",X"01",
		X"87",X"01",X"16",X"08",X"FF",X"68",X"01",X"17",X"01",X"68",X"01",X"17",X"01",X"58",X"01",X"17",
		X"01",X"58",X"01",X"17",X"01",X"48",X"01",X"17",X"01",X"48",X"01",X"17",X"01",X"38",X"01",X"17",
		X"01",X"38",X"01",X"17",X"01",X"28",X"01",X"B8",X"01",X"28",X"01",X"B8",X"01",X"28",X"01",X"B8",
		X"01",X"28",X"01",X"B8",X"01",X"18",X"01",X"B8",X"01",X"18",X"01",X"B8",X"01",X"38",X"01",X"B8",
		X"01",X"58",X"01",X"B8",X"01",X"68",X"01",X"17",X"01",X"68",X"01",X"17",X"01",X"58",X"01",X"17",
		X"01",X"58",X"01",X"17",X"01",X"48",X"01",X"17",X"01",X"48",X"01",X"17",X"01",X"38",X"01",X"17",
		X"01",X"38",X"01",X"17",X"01",X"28",X"01",X"B8",X"01",X"28",X"01",X"B8",X"01",X"28",X"01",X"B8",
		X"01",X"28",X"01",X"B8",X"01",X"18",X"01",X"B8",X"01",X"18",X"01",X"B8",X"01",X"38",X"01",X"B8",
		X"01",X"58",X"01",X"B8",X"01",X"FF",X"26",X"01",X"36",X"01",X"66",X"01",X"A6",X"01",X"15",X"01",
		X"A6",X"01",X"66",X"01",X"36",X"01",X"FF",X"86",X"01",X"05",X"01",X"15",X"01",X"55",X"01",X"86",
		X"01",X"05",X"01",X"15",X"01",X"55",X"01",X"86",X"01",X"05",X"01",X"15",X"01",X"55",X"01",X"FF",
		X"66",X"01",X"86",X"01",X"A6",X"01",X"36",X"01",X"16",X"01",X"C0",X"01",X"35",X"01",X"C0",X"01",
		X"15",X"04",X"FF",X"0A",X"01",X"7A",X"01",X"29",X"01",X"99",X"01",X"48",X"01",X"B8",X"01",X"67",
		X"01",X"57",X"01",X"67",X"01",X"77",X"01",X"67",X"01",X"FF",X"16",X"01",X"06",X"01",X"B7",X"01",
		X"A7",X"01",X"B7",X"01",X"A7",X"01",X"97",X"01",X"87",X"01",X"97",X"01",X"87",X"01",X"77",X"01",
		X"67",X"01",X"77",X"01",X"67",X"01",X"57",X"01",X"47",X"01",X"37",X"01",X"B7",X"01",X"77",X"01",
		X"36",X"01",X"FF",X"77",X"01",X"67",X"01",X"57",X"01",X"47",X"01",X"57",X"01",X"47",X"01",X"37",
		X"01",X"27",X"01",X"37",X"01",X"27",X"01",X"17",X"01",X"07",X"01",X"17",X"01",X"07",X"01",X"B8",
		X"01",X"A8",X"01",X"98",X"01",X"57",X"01",X"17",X"01",X"97",X"01",X"FF",X"47",X"01",X"37",X"01",
		X"27",X"01",X"17",X"01",X"27",X"01",X"17",X"01",X"07",X"01",X"B8",X"01",X"07",X"01",X"B8",X"01",
		X"A8",X"01",X"98",X"01",X"A8",X"01",X"98",X"01",X"88",X"01",X"78",X"01",X"68",X"01",X"27",X"01",
		X"A8",X"01",X"67",X"01",X"FF",X"55",X"01",X"A5",X"01",X"55",X"01",X"A5",X"01",X"55",X"01",X"A5",
		X"01",X"55",X"01",X"A5",X"01",X"55",X"01",X"A5",X"01",X"55",X"01",X"A5",X"01",X"55",X"01",X"A5",
		X"01",X"55",X"01",X"A5",X"01",X"55",X"01",X"A5",X"01",X"55",X"01",X"A5",X"01",X"55",X"01",X"A5",
		X"01",X"55",X"01",X"A5",X"01",X"FF",X"09",X"04",X"19",X"04",X"29",X"04",X"39",X"04",X"49",X"04",
		X"39",X"04",X"FF",X"16",X"01",X"A7",X"01",X"A7",X"01",X"A7",X"01",X"26",X"01",X"A7",X"01",X"A7",
		X"01",X"A7",X"01",X"36",X"01",X"A7",X"01",X"A7",X"01",X"A7",X"05",X"FF",X"27",X"01",X"17",X"01",
		X"27",X"01",X"17",X"01",X"27",X"01",X"17",X"01",X"27",X"01",X"17",X"01",X"27",X"01",X"17",X"01",
		X"27",X"01",X"17",X"05",X"FF",X"16",X"01",X"16",X"01",X"A7",X"01",X"16",X"01",X"36",X"01",X"56",
		X"01",X"66",X"01",X"86",X"01",X"A6",X"01",X"A6",X"01",X"A6",X"01",X"A6",X"05",X"FF",X"68",X"01",
		X"18",X"02",X"18",X"01",X"68",X"01",X"18",X"02",X"18",X"01",X"68",X"01",X"18",X"02",X"18",X"02",
		X"18",X"01",X"18",X"01",X"18",X"01",X"FF",X"75",X"01",X"B5",X"01",X"34",X"01",X"64",X"01",X"75",
		X"02",X"FF",X"76",X"01",X"B6",X"01",X"35",X"01",X"65",X"01",X"76",X"02",X"FF",X"57",X"01",X"17",
		X"01",X"98",X"01",X"68",X"01",X"57",X"02",X"FF",X"55",X"01",X"65",X"01",X"95",X"01",X"A5",X"01",
		X"04",X"01",X"34",X"01",X"14",X"01",X"A5",X"01",X"FF",X"15",X"01",X"A6",X"01",X"15",X"01",X"25",
		X"01",X"A6",X"01",X"25",X"01",X"35",X"01",X"A6",X"01",X"35",X"01",X"25",X"01",X"A6",X"01",X"25",
		X"01",X"15",X"01",X"A6",X"01",X"15",X"01",X"05",X"01",X"A6",X"01",X"05",X"01",X"C0",X"02",X"26",
		X"01",X"C0",X"02",X"26",X"01",X"96",X"01",X"66",X"01",X"96",X"01",X"A6",X"01",X"66",X"01",X"A6",
		X"01",X"B6",X"01",X"66",X"01",X"B6",X"01",X"A6",X"01",X"66",X"01",X"A6",X"01",X"96",X"01",X"66",
		X"01",X"96",X"01",X"A6",X"01",X"66",X"01",X"A6",X"01",X"C0",X"02",X"26",X"01",X"C0",X"02",X"26",
		X"01",X"FF",X"A6",X"01",X"66",X"01",X"A6",X"01",X"A6",X"01",X"66",X"01",X"A6",X"01",X"A6",X"01",
		X"66",X"01",X"A6",X"01",X"A6",X"01",X"66",X"01",X"A6",X"01",X"A6",X"01",X"66",X"01",X"A6",X"01",
		X"A6",X"01",X"66",X"01",X"A6",X"01",X"C0",X"02",X"06",X"01",X"C0",X"02",X"06",X"01",X"66",X"01",
		X"06",X"01",X"66",X"01",X"66",X"01",X"16",X"01",X"66",X"01",X"66",X"01",X"26",X"01",X"66",X"01",
		X"66",X"01",X"16",X"01",X"66",X"01",X"66",X"01",X"06",X"01",X"66",X"01",X"66",X"01",X"16",X"01",
		X"66",X"01",X"C0",X"02",X"06",X"01",X"C0",X"02",X"06",X"01",X"FF",X"69",X"04",X"C0",X"01",X"69",
		X"03",X"C0",X"01",X"69",X"02",X"C0",X"01",X"69",X"04",X"C0",X"01",X"69",X"03",X"C0",X"01",X"69",
		X"02",X"C0",X"01",X"18",X"04",X"C0",X"01",X"18",X"03",X"C0",X"01",X"18",X"02",X"C0",X"01",X"18",
		X"04",X"C0",X"01",X"18",X"03",X"C0",X"01",X"18",X"02",X"C0",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C7");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
