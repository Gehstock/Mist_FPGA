library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_M4 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_M4 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"6C",X"C6",X"C6",X"FE",X"C6",X"C6",
		X"00",X"FC",X"C6",X"C6",X"FC",X"C6",X"C6",X"FC",X"00",X"3C",X"66",X"C0",X"C0",X"C0",X"66",X"3C",
		X"00",X"F8",X"CC",X"C6",X"C6",X"C6",X"CC",X"F8",X"00",X"FC",X"C0",X"C0",X"F8",X"C0",X"C0",X"FE",
		X"00",X"FE",X"C0",X"C0",X"FC",X"C0",X"C0",X"C0",X"00",X"3E",X"60",X"C0",X"CE",X"C6",X"66",X"3E",
		X"00",X"C6",X"C6",X"C6",X"FE",X"C6",X"C6",X"C6",X"00",X"FC",X"30",X"30",X"30",X"30",X"30",X"FC",
		X"00",X"06",X"06",X"06",X"06",X"06",X"C6",X"7C",X"00",X"C6",X"CC",X"D8",X"F0",X"F8",X"DC",X"CE",
		X"00",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"FE",X"00",X"C6",X"EE",X"FE",X"FE",X"D6",X"C6",X"C6",
		X"00",X"C6",X"E6",X"F6",X"FE",X"DE",X"CE",X"C6",X"00",X"7C",X"C6",X"C6",X"C6",X"C6",X"C6",X"7C",
		X"00",X"FC",X"C6",X"C6",X"C6",X"FC",X"C0",X"C0",X"00",X"FE",X"C0",X"C0",X"FE",X"C0",X"C3",X"C3",
		X"00",X"FC",X"C6",X"C6",X"CE",X"F8",X"DC",X"CE",X"00",X"78",X"CC",X"C0",X"7C",X"06",X"C6",X"7C",
		X"00",X"FC",X"30",X"30",X"30",X"30",X"30",X"30",X"00",X"C6",X"C6",X"C6",X"C6",X"C6",X"C6",X"7C",
		X"00",X"C6",X"C6",X"C6",X"EE",X"7C",X"38",X"10",X"00",X"C6",X"C6",X"D6",X"FE",X"FE",X"EE",X"C6",
		X"00",X"C4",X"C4",X"C0",X"C0",X"C0",X"C0",X"FE",X"00",X"CC",X"CC",X"CC",X"78",X"30",X"30",X"30",
		X"00",X"FE",X"0E",X"1C",X"38",X"70",X"E0",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"01",X"07",X"0E",X"0C",X"1F",X"7F",X"FF",X"C1",X"86",X"00",X"1E",X"FC",X"F8",X"F8",X"F0",
		X"01",X"03",X"07",X"0F",X"1F",X"1F",X"0F",X"07",X"E0",X"E0",X"C0",X"C0",X"80",X"80",X"00",X"00",
		X"03",X"03",X"07",X"07",X"0F",X"1F",X"7F",X"FF",X"FF",X"FE",X"FE",X"FC",X"FC",X"F8",X"F0",X"E0",
		X"F1",X"FB",X"FE",X"FC",X"F8",X"F0",X"C0",X"80",X"01",X"01",X"00",X"00",X"01",X"07",X"0F",X"01",
		X"01",X"07",X"1F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"F8",X"F8",X"F0",X"F0",X"E0",X"80",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"F0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"18",X"18",X"00",X"00",X"18",X"18",X"00",X"FC",X"FC",X"FC",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"0F",X"0F",X"07",X"03",X"03",X"01",X"00",X"00",X"FF",X"FF",X"FF",X"FC",X"F0",X"E0",X"C0",X"80",
		X"00",X"38",X"4C",X"C6",X"C6",X"C6",X"64",X"38",X"00",X"30",X"70",X"30",X"30",X"30",X"30",X"FC",
		X"00",X"7C",X"C6",X"0E",X"3C",X"78",X"E0",X"FE",X"00",X"7E",X"0C",X"18",X"3C",X"06",X"C6",X"7C",
		X"00",X"1C",X"3C",X"6C",X"CC",X"FE",X"0C",X"0C",X"00",X"FC",X"C0",X"FC",X"06",X"06",X"C6",X"7C",
		X"00",X"3C",X"60",X"C0",X"FC",X"C6",X"C6",X"7C",X"00",X"FE",X"C6",X"0C",X"18",X"30",X"30",X"30",
		X"00",X"78",X"C4",X"E4",X"78",X"9E",X"86",X"7C",X"00",X"7C",X"C6",X"C6",X"7E",X"06",X"0C",X"78",
		X"FE",X"FC",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"03",X"3F",X"7F",X"3F",
		X"80",X"00",X"00",X"00",X"80",X"C0",X"FC",X"FF",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",
		X"10",X"30",X"60",X"60",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"06",X"04",X"0C",X"08",
		X"F0",X"0E",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"20",X"10",X"08",X"04",
		X"04",X"02",X"02",X"02",X"01",X"01",X"01",X"01",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"F0",X"8E",X"81",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"F0",X"4E",X"41",X"40",X"40",X"40",X"80",X"80",X"40",X"40",X"40",X"80",X"80",X"80",X"80",X"80",
		X"F0",X"1E",X"21",X"20",X"20",X"20",X"40",X"40",X"20",X"20",X"40",X"40",X"40",X"80",X"80",X"80",
		X"F0",X"0E",X"09",X"08",X"10",X"10",X"10",X"20",X"10",X"10",X"20",X"20",X"40",X"40",X"80",X"80",
		X"F0",X"0E",X"03",X"04",X"04",X"08",X"08",X"10",X"08",X"10",X"10",X"20",X"20",X"40",X"80",X"80",
		X"F0",X"0E",X"01",X"01",X"02",X"02",X"04",X"08",X"04",X"08",X"10",X"10",X"20",X"40",X"40",X"80",
		X"F0",X"0E",X"01",X"00",X"00",X"01",X"02",X"04",X"00",X"00",X"80",X"40",X"A0",X"10",X"08",X"04",
		X"02",X"04",X"08",X"08",X"10",X"20",X"40",X"80",X"F0",X"0E",X"01",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"80",X"40",X"20",X"50",X"88",X"04",X"00",X"01",X"02",X"0C",X"10",X"20",X"40",X"80",
		X"84",X"02",X"02",X"02",X"01",X"01",X"01",X"01",X"00",X"00",X"80",X"40",X"20",X"10",X"28",X"44",
		X"00",X"00",X"01",X"02",X"0C",X"10",X"60",X"80",X"24",X"42",X"82",X"02",X"01",X"01",X"01",X"01",
		X"00",X"00",X"80",X"40",X"20",X"10",X"08",X"14",X"00",X"00",X"00",X"01",X"06",X"18",X"20",X"C0",
		X"0C",X"32",X"42",X"82",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"03",X"0C",X"30",X"C0",
		X"04",X"06",X"1A",X"62",X"81",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"03",X"1C",X"E0",
		X"04",X"02",X"02",X"0E",X"71",X"81",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"F8",
		X"04",X"02",X"02",X"02",X"03",X"3D",X"C1",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"04",X"02",X"02",X"02",X"01",X"01",X"3F",X"C1",X"01",X"01",X"01",X"01",X"02",X"02",X"02",X"04",
		X"04",X"08",X"10",X"20",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"0E",X"F0",
		X"FF",X"00",X"00",X"02",X"06",X"04",X"0C",X"08",X"FF",X"01",X"01",X"01",X"02",X"02",X"02",X"04",
		X"FF",X"00",X"00",X"02",X"06",X"04",X"0C",X"08",X"C1",X"3F",X"01",X"01",X"02",X"02",X"02",X"04",
		X"F8",X"07",X"00",X"02",X"06",X"04",X"0C",X"08",X"01",X"C1",X"3D",X"03",X"02",X"02",X"02",X"04",
		X"E0",X"1C",X"03",X"02",X"06",X"04",X"0C",X"08",X"01",X"01",X"81",X"71",X"0E",X"02",X"02",X"04",
		X"C0",X"30",X"0C",X"03",X"06",X"04",X"0C",X"08",X"01",X"01",X"01",X"81",X"62",X"1A",X"06",X"04",
		X"C0",X"20",X"18",X"06",X"07",X"04",X"0C",X"08",X"01",X"01",X"01",X"01",X"82",X"42",X"32",X"0C",
		X"80",X"60",X"10",X"0E",X"06",X"05",X"0C",X"08",X"01",X"01",X"01",X"01",X"02",X"82",X"42",X"24",
		X"14",X"08",X"10",X"20",X"40",X"80",X"00",X"00",X"80",X"40",X"20",X"12",X"0E",X"06",X"0D",X"08",
		X"01",X"01",X"01",X"01",X"02",X"02",X"02",X"84",X"44",X"28",X"10",X"20",X"40",X"80",X"00",X"00",
		X"80",X"40",X"20",X"12",X"0E",X"0C",X"0C",X"0A",X"01",X"00",X"00",X"00",X"00",X"01",X"0E",X"F0",
		X"04",X"88",X"50",X"20",X"40",X"80",X"00",X"00",X"80",X"40",X"40",X"22",X"16",X"14",X"0C",X"0C",
		X"04",X"02",X"01",X"00",X"00",X"01",X"0E",X"F0",X"04",X"08",X"10",X"A0",X"40",X"80",X"00",X"00",
		X"80",X"80",X"40",X"22",X"26",X"14",X"1C",X"08",X"08",X"04",X"02",X"02",X"01",X"01",X"0E",X"F0",
		X"80",X"80",X"40",X"42",X"26",X"24",X"1C",X"18",X"10",X"08",X"08",X"04",X"04",X"03",X"0E",X"F0",
		X"80",X"80",X"80",X"42",X"46",X"44",X"2C",X"28",X"20",X"10",X"10",X"10",X"08",X"09",X"0E",X"F0",
		X"80",X"80",X"80",X"82",X"86",X"44",X"4C",X"48",X"40",X"40",X"20",X"20",X"20",X"21",X"1E",X"F0",
		X"80",X"80",X"80",X"82",X"86",X"84",X"8C",X"88",X"80",X"80",X"40",X"40",X"40",X"41",X"4E",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"80",X"70",X"0F",X"20",X"10",X"08",X"04",X"02",X"01",X"00",X"00",
		X"80",X"80",X"80",X"80",X"40",X"40",X"40",X"20",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"81",X"71",X"0F",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"02",X"02",X"02",X"82",X"72",X"0F",X"01",X"01",X"01",X"01",X"01",X"02",X"02",X"02",
		X"02",X"02",X"04",X"04",X"04",X"84",X"78",X"0F",X"01",X"01",X"01",X"02",X"02",X"02",X"04",X"04",
		X"04",X"08",X"08",X"08",X"10",X"90",X"70",X"0F",X"01",X"01",X"02",X"02",X"04",X"04",X"08",X"08",
		X"08",X"10",X"10",X"20",X"20",X"C0",X"70",X"0F",X"01",X"01",X"02",X"04",X"04",X"08",X"08",X"10",
		X"10",X"20",X"40",X"40",X"80",X"80",X"70",X"0F",X"01",X"02",X"02",X"04",X"08",X"08",X"10",X"20",
		X"40",X"40",X"80",X"00",X"00",X"80",X"70",X"0F",X"20",X"10",X"08",X"05",X"02",X"01",X"00",X"00",
		X"01",X"02",X"04",X"08",X"10",X"10",X"20",X"40",X"80",X"00",X"00",X"00",X"00",X"80",X"70",X"0F",
		X"20",X"11",X"0A",X"04",X"02",X"01",X"00",X"00",X"01",X"02",X"04",X"08",X"30",X"40",X"80",X"00",
		X"80",X"80",X"80",X"80",X"40",X"40",X"40",X"21",X"22",X"14",X"08",X"04",X"02",X"01",X"00",X"00",
		X"01",X"06",X"08",X"30",X"40",X"80",X"00",X"00",X"80",X"80",X"80",X"80",X"40",X"41",X"42",X"24",
		X"28",X"10",X"08",X"04",X"02",X"01",X"00",X"00",X"03",X"04",X"18",X"60",X"80",X"00",X"00",X"00",
		X"80",X"80",X"80",X"80",X"41",X"42",X"4C",X"30",X"03",X"0C",X"30",X"C0",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"81",X"46",X"58",X"60",X"20",X"07",X"38",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"81",X"8E",X"70",X"40",X"40",X"20",X"1F",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"83",X"BC",X"C0",X"40",X"40",X"40",X"20",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"83",X"7C",X"80",X"80",X"40",X"40",X"40",X"20",X"20",X"40",X"40",X"40",X"80",X"80",X"80",X"80",
		X"00",X"00",X"01",X"02",X"04",X"08",X"10",X"20",X"0F",X"70",X"80",X"00",X"00",X"00",X"00",X"00",
		X"10",X"30",X"60",X"60",X"40",X"00",X"00",X"FF",X"20",X"40",X"40",X"40",X"80",X"80",X"80",X"FF",
		X"10",X"30",X"60",X"60",X"40",X"00",X"00",X"FF",X"20",X"40",X"40",X"40",X"80",X"80",X"FC",X"83",
		X"10",X"30",X"60",X"60",X"40",X"00",X"E0",X"1F",X"20",X"40",X"40",X"40",X"C0",X"BC",X"83",X"80",
		X"10",X"30",X"60",X"60",X"40",X"C0",X"38",X"07",X"20",X"40",X"40",X"70",X"8E",X"81",X"80",X"80",
		X"10",X"30",X"60",X"60",X"C0",X"30",X"0C",X"03",X"20",X"60",X"58",X"46",X"81",X"80",X"80",X"80",
		X"10",X"30",X"60",X"E0",X"60",X"18",X"04",X"03",X"30",X"4C",X"42",X"41",X"80",X"80",X"80",X"80",
		X"10",X"30",X"E0",X"60",X"70",X"08",X"06",X"01",X"24",X"42",X"41",X"40",X"80",X"80",X"80",X"80",
		X"00",X"00",X"01",X"02",X"04",X"08",X"10",X"28",X"10",X"B0",X"60",X"70",X"48",X"04",X"02",X"01",
		X"21",X"40",X"40",X"40",X"80",X"80",X"80",X"80",X"00",X"00",X"01",X"02",X"04",X"08",X"14",X"22",
		X"50",X"30",X"70",X"70",X"48",X"04",X"02",X"01",X"0F",X"70",X"80",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"01",X"02",X"04",X"0A",X"11",X"20",X"30",X"30",X"68",X"68",X"44",X"02",X"02",X"01",
		X"0F",X"70",X"80",X"00",X"00",X"80",X"40",X"20",X"00",X"00",X"01",X"02",X"05",X"08",X"10",X"20",
		X"10",X"38",X"68",X"64",X"44",X"02",X"01",X"01",X"0F",X"70",X"80",X"80",X"40",X"40",X"20",X"10",
		X"18",X"38",X"64",X"64",X"42",X"02",X"01",X"01",X"0F",X"70",X"C0",X"20",X"20",X"10",X"10",X"08",
		X"14",X"34",X"62",X"62",X"42",X"01",X"01",X"01",X"0F",X"70",X"90",X"10",X"08",X"08",X"08",X"04",
		X"12",X"32",X"62",X"61",X"41",X"01",X"01",X"01",X"0F",X"78",X"84",X"04",X"04",X"04",X"02",X"02",
		X"11",X"31",X"61",X"61",X"41",X"01",X"01",X"01",X"0F",X"72",X"82",X"02",X"02",X"02",X"01",X"01",
		X"F0",X"0E",X"61",X"60",X"00",X"00",X"00",X"00",X"F0",X"0E",X"01",X"00",X"00",X"60",X"60",X"00",
		X"F0",X"0E",X"01",X"00",X"06",X"06",X"00",X"00",X"00",X"00",X"80",X"40",X"20",X"10",X"C8",X"C4",
		X"04",X"62",X"62",X"02",X"01",X"01",X"01",X"01",X"04",X"02",X"02",X"02",X"01",X"61",X"61",X"01",
		X"04",X"02",X"02",X"02",X"01",X"0D",X"0D",X"01",X"01",X"61",X"61",X"01",X"02",X"02",X"02",X"04",
		X"01",X"0D",X"0D",X"01",X"02",X"02",X"02",X"04",X"01",X"01",X"01",X"01",X"02",X"62",X"62",X"04",
		X"C4",X"C8",X"10",X"20",X"40",X"80",X"00",X"00",X"00",X"06",X"06",X"00",X"00",X"01",X"0E",X"F0",
		X"00",X"60",X"60",X"00",X"00",X"01",X"0E",X"F0",X"00",X"00",X"00",X"00",X"60",X"61",X"0E",X"F0",
		X"00",X"06",X"06",X"00",X"00",X"80",X"70",X"0F",X"00",X"00",X"00",X"00",X"06",X"86",X"70",X"0F",
		X"00",X"60",X"60",X"00",X"00",X"80",X"70",X"0F",X"23",X"13",X"08",X"04",X"02",X"01",X"00",X"00",
		X"80",X"80",X"80",X"80",X"40",X"46",X"46",X"20",X"80",X"86",X"86",X"80",X"40",X"40",X"40",X"20",
		X"80",X"B0",X"B0",X"80",X"40",X"40",X"40",X"20",X"20",X"40",X"40",X"40",X"80",X"86",X"86",X"80",
		X"20",X"40",X"40",X"40",X"80",X"B0",X"B0",X"80",X"20",X"46",X"46",X"40",X"80",X"80",X"80",X"80",
		X"00",X"00",X"01",X"02",X"04",X"08",X"13",X"23",X"0F",X"70",X"80",X"00",X"00",X"60",X"60",X"00",
		X"0F",X"70",X"80",X"00",X"00",X"06",X"06",X"00",X"0F",X"70",X"86",X"06",X"00",X"00",X"00",X"00",
		X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",
		X"30",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"30",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"30",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"30",
		X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0C",
		X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
