-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

entity ROM_PGM_0 is
  port (
    CLK         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM_0 is


  type ROM_ARRAY is array(0 to 10087) of std_logic_vector(7 downto 0);
  constant ROM : ROM_ARRAY := (
    x"31",x"00",x"44",x"AF",x"C3",x"00",x"03",x"C3", -- 0x0000
    x"46",x"0B",x"55",x"50",x"4F",x"00",x"84",x"54", -- 0x0008
    x"77",x"23",x"10",x"FC",x"C9",x"06",x"C2",x"4C", -- 0x0010
    x"41",x"43",x"4B",x"4F",x"49",x"00",x"85",x"43", -- 0x0018
    x"C3",x"B4",x"04",x"45",x"00",x"10",x"00",x"05", -- 0x0020
    x"C3",x"0B",x"05",x"56",x"45",x"00",x"10",x"00", -- 0x0028
    x"85",x"42",x"49",x"4E",x"49",x"54",x"61",x"00", -- 0x0030
    x"C3",x"00",x"00",x"05",x"49",x"54",x"5E",x"00", -- 0x0038
    x"C3",x"00",x"10",x"41",x"4C",x"4F",x"C3",x"6A", -- 0x0040
    x"14",x"C3",x"7A",x"06",x"C3",x"EF",x"05",x"C3", -- 0x0048
    x"5C",x"03",x"C3",x"70",x"0C",x"C9",x"7B",x"15", -- 0x0050
    x"C3",x"BE",x"15",x"C3",x"46",x"0B",x"C3",x"F8", -- 0x0058
    x"0A",x"C3",x"6E",x"07",x"45",x"70",x"F5",x"AF", -- 0x0060
    x"32",x"01",x"70",x"08",x"3A",x"00",x"78",x"08", -- 0x0068
    x"C5",x"D5",x"E5",x"DD",x"E5",x"FD",x"E5",x"21", -- 0x0070
    x"00",x"43",x"11",x"00",x"58",x"01",x"80",x"00", -- 0x0078
    x"ED",x"B0",x"CD",x"FC",x"00",x"CD",x"CB",x"0C", -- 0x0080
    x"21",x"02",x"40",x"34",x"23",x"CD",x"77",x"05", -- 0x0088
    x"CD",x"D5",x"05",x"CD",x"46",x"00",x"CD",x"DD", -- 0x0090
    x"0A",x"CD",x"40",x"00",x"CD",x"85",x"06",x"3A", -- 0x0098
    x"10",x"40",x"F5",x"CB",x"47",x"28",x"05",x"CD", -- 0x00A0
    x"7D",x"05",x"18",x"0C",x"21",x"40",x"50",x"22", -- 0x00A8
    x"18",x"40",x"CD",x"92",x"07",x"CD",x"70",x"0B", -- 0x00B0
    x"F1",x"FD",x"E1",x"DD",x"E1",x"E1",x"D1",x"C1", -- 0x00B8
    x"3E",x"01",x"32",x"01",x"70",x"F1",x"C9",x"01", -- 0x00C0
    x"70",x"F1",x"C9",x"C1",x"3E",x"01",x"32",x"01", -- 0x00C8
    x"70",x"F1",x"C9",x"00",x"00",x"00",x"00",x"00", -- 0x00D0
    x"C3",x"3E",x"03",x"00",x"00",x"C3",x"FD",x"14", -- 0x00D8
    x"C3",x"C1",x"0B",x"C3",x"12",x"01",x"C3",x"53", -- 0x00E0
    x"01",x"C3",x"8E",x"01",x"C3",x"B1",x"01",x"00", -- 0x00E8
    x"C3",x"00",x"0D",x"C9",x"00",x"1A",x"C3",x"08", -- 0x00F0
    x"0A",x"C3",x"59",x"21",x"C3",x"E1",x"21",x"00", -- 0x00F8
    x"02",x"10",x"06",x"52",x"45",x"41",x"44",x"59", -- 0x0100
    x"40",x"50",x"4C",x"41",x"59",x"45",x"52",x"40", -- 0x0108
    x"31",x"FF",x"11",x"00",x"00",x"3A",x"14",x"40", -- 0x0110
    x"CB",x"5F",x"28",x"06",x"DD",x"21",x"00",x"41", -- 0x0118
    x"18",x"04",x"DD",x"21",x"00",x"42",x"DD",x"7E", -- 0x0120
    x"08",x"B7",x"28",x"18",x"21",x"4B",x"01",x"5F", -- 0x0128
    x"19",x"7E",x"07",x"07",x"07",x"4F",x"21",x"05", -- 0x0130
    x"43",x"71",x"23",x"23",x"7D",x"FE",x"3F",x"38", -- 0x0138
    x"F8",x"DD",x"7E",x"08",x"3C",x"E6",x"07",x"DD", -- 0x0140
    x"77",x"08",x"C9",x"00",x"20",x"40",x"60",x"80", -- 0x0148
    x"A0",x"C0",x"E0",x"3A",x"14",x"40",x"01",x"00", -- 0x0150
    x"00",x"11",x"40",x"50",x"CB",x"5F",x"28",x"05", -- 0x0158
    x"21",x"10",x"41",x"18",x"03",x"21",x"10",x"42", -- 0x0160
    x"7D",x"FE",x"FD",x"30",x"1E",x"7A",x"FE",x"54", -- 0x0168
    x"28",x"19",x"78",x"FE",x"FF",x"0E",x"10",x"28", -- 0x0170
    x"08",x"1A",x"4F",x"E6",x"FC",x"FE",x"30",x"20", -- 0x0178
    x"06",x"70",x"23",x"71",x"23",x"06",x"00",x"13", -- 0x0180
    x"04",x"18",x"DD",x"36",x"00",x"C9",x"3A",x"14", -- 0x0188
    x"40",x"11",x"40",x"50",x"CB",x"5F",x"28",x"05", -- 0x0190
    x"21",x"10",x"41",x"18",x"03",x"21",x"10",x"42", -- 0x0198
    x"7A",x"FE",x"54",x"C8",x"7E",x"47",x"B7",x"C8", -- 0x01A0
    x"13",x"10",x"FD",x"23",x"7E",x"12",x"23",x"18", -- 0x01A8
    x"EF",x"0E",x"00",x"21",x"01",x"43",x"CD",x"36", -- 0x01B0
    x"01",x"3A",x"01",x"40",x"E6",x"F0",x"32",x"01", -- 0x01B8
    x"40",x"AF",x"21",x"00",x"60",x"06",x"00",x"D7", -- 0x01C0
    x"21",x"00",x"68",x"D7",x"3E",x"FF",x"32",x"00", -- 0x01C8
    x"78",x"3A",x"14",x"40",x"CB",x"5F",x"28",x"0A", -- 0x01D0
    x"DD",x"21",x"00",x"41",x"FD",x"21",x"00",x"42", -- 0x01D8
    x"18",x"08",x"DD",x"21",x"00",x"42",x"FD",x"21", -- 0x01E0
    x"00",x"41",x"CB",x"7F",x"20",x"73",x"DD",x"7E", -- 0x01E8
    x"09",x"3D",x"B7",x"28",x"2E",x"DD",x"77",x"09", -- 0x01F0
    x"DD",x"7E",x"0A",x"FE",x"0F",x"28",x"01",x"3C", -- 0x01F8
    x"DD",x"77",x"0A",x"F5",x"DD",x"7E",x"05",x"FE", -- 0x0200
    x"1A",x"30",x"08",x"DD",x"34",x"05",x"21",x"00", -- 0x0208
    x"23",x"7E",x"47",x"F1",x"B8",x"DA",x"CC",x"02", -- 0x0210
    x"DD",x"7E",x"06",x"CB",x"A7",x"DD",x"77",x"06", -- 0x0218
    x"C3",x"CC",x"02",x"AF",x"32",x"10",x"40",x"CD", -- 0x0220
    x"49",x"00",x"3E",x"C0",x"CD",x"4C",x"00",x"11", -- 0x0228
    x"D0",x"02",x"E7",x"3E",x"80",x"CD",x"4C",x"00", -- 0x0230
    x"31",x"00",x"44",x"21",x"03",x"41",x"06",x"F8", -- 0x0238
    x"AF",x"D7",x"21",x"03",x"42",x"06",x"F8",x"D7", -- 0x0240
    x"21",x"00",x"43",x"06",x"80",x"D7",x"21",x"1C", -- 0x0248
    x"1F",x"22",x"05",x"41",x"22",x"05",x"42",x"CD", -- 0x0250
    x"49",x"00",x"AF",x"32",x"2F",x"40",x"C3",x"D8", -- 0x0258
    x"00",x"DD",x"7E",x"09",x"3D",x"B7",x"28",x"3B", -- 0x0260
    x"DD",x"77",x"09",x"DD",x"7E",x"0A",x"3C",x"DD", -- 0x0268
    x"77",x"0A",x"3A",x"14",x"40",x"EE",x"18",x"32", -- 0x0270
    x"14",x"40",x"CD",x"49",x"00",x"CD",x"00",x"25", -- 0x0278
    x"3E",x"E0",x"CD",x"4C",x"00",x"11",x"DD",x"02", -- 0x0280
    x"E7",x"3A",x"14",x"40",x"CB",x"5F",x"28",x"0E", -- 0x0288
    x"11",x"E6",x"02",x"E7",x"3E",x"C0",x"CD",x"4C", -- 0x0290
    x"00",x"CD",x"49",x"00",x"18",x"2E",x"11",x"F3", -- 0x0298
    x"02",x"18",x"F0",x"11",x"D0",x"02",x"E7",x"3E", -- 0x02A0
    x"C0",x"CD",x"4C",x"00",x"3A",x"14",x"40",x"CB", -- 0x02A8
    x"5F",x"28",x"06",x"11",x"E6",x"02",x"E7",x"18", -- 0x02B0
    x"03",x"11",x"F3",x"02",x"E7",x"3E",x"C0",x"CD", -- 0x02B8
    x"4C",x"00",x"CD",x"49",x"00",x"3A",x"14",x"40", -- 0x02C0
    x"CB",x"BF",x"18",x"A9",x"CD",x"12",x"01",x"C9", -- 0x02C8
    x"04",x"0C",x"08",x"47",x"41",x"4D",x"45",x"40", -- 0x02D0
    x"4F",x"56",x"45",x"52",x"FF",x"05",x"0C",x"0C", -- 0x02D8
    x"52",x"45",x"41",x"44",x"59",x"FF",x"05",x"0E", -- 0x02E0
    x"0A",x"50",x"4C",x"41",x"59",x"45",x"52",x"40", -- 0x02E8
    x"40",x"31",x"FF",x"05",x"0E",x"0A",x"50",x"4C", -- 0x02F0
    x"41",x"59",x"45",x"52",x"40",x"40",x"32",x"FF", -- 0x02F8
    x"08",x"3A",x"00",x"78",x"08",x"AF",x"32",x"01", -- 0x0300
    x"70",x"21",x"00",x"50",x"3E",x"10",x"06",x"00", -- 0x0308
    x"D7",x"D7",x"D7",x"D7",x"08",x"3A",x"00",x"78", -- 0x0310
    x"08",x"21",x"00",x"58",x"AF",x"D7",x"08",x"3A", -- 0x0318
    x"00",x"78",x"08",x"21",x"00",x"68",x"D7",x"21", -- 0x0320
    x"00",x"60",x"D7",x"08",x"3A",x"00",x"78",x"08", -- 0x0328
    x"21",x"00",x"70",x"D7",x"21",x"00",x"40",x"AF", -- 0x0330
    x"D7",x"D7",x"D7",x"06",x"F8",x"D7",x"3E",x"FF", -- 0x0338
    x"32",x"00",x"78",x"08",x"3A",x"00",x"78",x"08", -- 0x0340
    x"21",x"FF",x"FF",x"22",x"C0",x"40",x"3E",x"01", -- 0x0348
    x"32",x"01",x"70",x"11",x"00",x"04",x"E7",x"CD", -- 0x0350
    x"84",x"07",x"18",x"23",x"21",x"00",x"50",x"22", -- 0x0358
    x"18",x"40",x"21",x"50",x"40",x"06",x"30",x"D7", -- 0x0360
    x"3E",x"08",x"32",x"11",x"40",x"CD",x"6E",x"07", -- 0x0368
    x"3E",x"01",x"32",x"01",x"70",x"3E",x"E0",x"CD", -- 0x0370
    x"EF",x"05",x"C9",x"AF",x"32",x"0C",x"40",x"3A", -- 0x0378
    x"10",x"40",x"CB",x"D7",x"CB",x"C7",x"32",x"10", -- 0x0380
    x"40",x"CD",x"C1",x"0B",x"C3",x"00",x"1E",x"00", -- 0x0388
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0390
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0398
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03F8
    x"06",x"00",x"00",x"53",x"43",x"4F",x"52",x"45", -- 0x0400
    x"31",x"40",x"40",x"40",x"40",x"48",x"49",x"40", -- 0x0408
    x"53",x"43",x"4F",x"52",x"45",x"40",x"40",x"40", -- 0x0410
    x"40",x"53",x"43",x"4F",x"52",x"45",x"32",x"FF", -- 0x0418
    x"05",x"01",x"00",x"00",x"41",x"06",x"05",x"01", -- 0x0420
    x"0B",x"34",x"40",x"06",x"05",x"01",x"16",x"00", -- 0x0428
    x"42",x"06",x"03",x"14",x"0D",x"06",x"40",x"02", -- 0x0430
    x"06",x"10",x"0B",x"43",x"52",x"45",x"44",x"49", -- 0x0438
    x"54",x"FF",x"05",x"08",x"04",x"50",x"52",x"45", -- 0x0440
    x"53",x"53",x"40",x"31",x"40",x"50",x"4C",x"41", -- 0x0448
    x"59",x"45",x"52",x"40",x"42",x"55",x"54",x"54", -- 0x0450
    x"4F",x"4E",x"FF",x"05",x"08",x"02",x"50",x"55", -- 0x0458
    x"53",x"48",x"40",x"31",x"40",x"4F",x"52",x"40", -- 0x0460
    x"32",x"40",x"50",x"4C",x"41",x"59",x"45",x"52", -- 0x0468
    x"40",x"42",x"55",x"54",x"54",x"4F",x"4E",x"FF", -- 0x0470
    x"05",x"0C",x"04",x"49",x"4E",x"53",x"45",x"52", -- 0x0478
    x"54",x"40",x"41",x"4E",x"4F",x"54",x"48",x"45", -- 0x0480
    x"52",x"40",x"43",x"4F",x"49",x"4E",x"FF",x"03", -- 0x0488
    x"14",x"0A",x"46",x"52",x"45",x"45",x"40",x"50", -- 0x0490
    x"4C",x"41",x"59",x"FF",x"02",x"1E",x"04",x"40", -- 0x0498
    x"40",x"41",x"52",x"4D",x"40",x"40",x"40",x"40", -- 0x04A0
    x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"31", -- 0x04A8
    x"39",x"38",x"31",x"FF",x"F5",x"C5",x"D5",x"E5", -- 0x04B0
    x"D5",x"DD",x"E1",x"DD",x"7E",x"01",x"87",x"06", -- 0x04B8
    x"00",x"4F",x"FD",x"21",x"00",x"43",x"FD",x"09", -- 0x04C0
    x"FD",x"36",x"00",x"00",x"DD",x"7E",x"00",x"FD", -- 0x04C8
    x"77",x"01",x"DD",x"46",x"02",x"3E",x"1B",x"90", -- 0x04D0
    x"B7",x"CA",x"E7",x"04",x"21",x"40",x"50",x"01", -- 0x04D8
    x"20",x"00",x"09",x"3D",x"C2",x"E2",x"04",x"DD", -- 0x04E0
    x"4E",x"01",x"06",x"00",x"09",x"01",x"E0",x"FF", -- 0x04E8
    x"DD",x"23",x"DD",x"23",x"DD",x"23",x"DD",x"7E", -- 0x04F0
    x"00",x"FE",x"FF",x"28",x"09",x"D6",x"30",x"77", -- 0x04F8
    x"09",x"DD",x"23",x"C3",x"F6",x"04",x"E1",x"D1", -- 0x0500
    x"C1",x"F1",x"C9",x"F5",x"C5",x"D5",x"E5",x"D5", -- 0x0508
    x"DD",x"E1",x"DD",x"7E",x"01",x"87",x"06",x"00", -- 0x0510
    x"4F",x"FD",x"21",x"00",x"43",x"FD",x"09",x"FD", -- 0x0518
    x"36",x"00",x"00",x"DD",x"7E",x"00",x"FD",x"77", -- 0x0520
    x"01",x"DD",x"46",x"02",x"3E",x"1B",x"90",x"B7", -- 0x0528
    x"CA",x"40",x"05",x"FD",x"21",x"40",x"50",x"01", -- 0x0530
    x"20",x"00",x"FD",x"09",x"3D",x"C2",x"3A",x"05", -- 0x0538
    x"DD",x"4E",x"01",x"06",x"00",x"FD",x"09",x"01", -- 0x0540
    x"E0",x"FF",x"DD",x"56",x"05",x"DD",x"66",x"04", -- 0x0548
    x"DD",x"6E",x"03",x"CB",x"42",x"CA",x"62",x"05", -- 0x0550
    x"7E",x"E6",x"0F",x"FD",x"77",x"00",x"23",x"C3", -- 0x0558
    x"6C",x"05",x"7E",x"0F",x"0F",x"0F",x"0F",x"E6", -- 0x0560
    x"0F",x"FD",x"77",x"00",x"FD",x"09",x"15",x"C2", -- 0x0568
    x"53",x"05",x"E1",x"D1",x"C1",x"F1",x"C9",x"7E", -- 0x0570
    x"B7",x"C8",x"3C",x"77",x"C9",x"CD",x"70",x"0C", -- 0x0578
    x"3E",x"1C",x"32",x"0B",x"40",x"2A",x"18",x"40", -- 0x0580
    x"3A",x"05",x"40",x"47",x"CB",x"43",x"20",x"20", -- 0x0588
    x"E6",x"1F",x"11",x"00",x"00",x"5F",x"19",x"3A", -- 0x0590
    x"0B",x"40",x"47",x"7D",x"E6",x"1F",x"FE",x"03", -- 0x0598
    x"38",x"29",x"B8",x"30",x"26",x"7C",x"FE",x"53", -- 0x05A0
    x"30",x"13",x"36",x"32",x"22",x"18",x"40",x"C9", -- 0x05A8
    x"DD",x"A6",x"06",x"F5",x"DD",x"7E",x"05",x"32", -- 0x05B0
    x"0B",x"40",x"F1",x"18",x"D5",x"7D",x"FE",x"BF", -- 0x05B8
    x"38",x"E8",x"3A",x"10",x"40",x"CB",x"87",x"32", -- 0x05C0
    x"10",x"40",x"C9",x"11",x"16",x"00",x"7D",x"E6", -- 0x05C8
    x"F0",x"6F",x"19",x"18",x"D0",x"3A",x"00",x"40", -- 0x05D0
    x"5F",x"3A",x"01",x"40",x"57",x"0F",x"AB",x"5F", -- 0x05D8
    x"ED",x"57",x"83",x"AA",x"07",x"07",x"07",x"AA", -- 0x05E0
    x"83",x"32",x"05",x"40",x"C9",x"3E",x"80",x"32", -- 0x05E8
    x"03",x"40",x"3A",x"03",x"40",x"B7",x"C8",x"18", -- 0x05F0
    x"F9",x"21",x"02",x"50",x"3E",x"10",x"06",x"1E", -- 0x05F8
    x"D7",x"11",x"02",x"00",x"19",x"7C",x"FE",x"54", -- 0x0600
    x"20",x"F2",x"AF",x"21",x"02",x"43",x"06",x"7D", -- 0x0608
    x"D7",x"C9",x"AF",x"21",x"40",x"40",x"06",x"A0", -- 0x0610
    x"D7",x"21",x"02",x"43",x"06",x"7C",x"D7",x"08", -- 0x0618
    x"3A",x"00",x"78",x"08",x"21",x"02",x"58",x"06", -- 0x0620
    x"7C",x"D7",x"21",x"00",x"60",x"06",x"07",x"D7", -- 0x0628
    x"21",x"00",x"68",x"06",x"07",x"D7",x"3E",x"FF", -- 0x0630
    x"32",x"00",x"78",x"C9",x"3A",x"00",x"60",x"CB", -- 0x0638
    x"47",x"28",x"06",x"3E",x"01",x"32",x"08",x"40", -- 0x0640
    x"C9",x"3A",x"08",x"40",x"B7",x"C8",x"3A",x"07", -- 0x0648
    x"40",x"3C",x"32",x"07",x"40",x"AF",x"32",x"08", -- 0x0650
    x"40",x"3A",x"10",x"40",x"E6",x"18",x"B7",x"C0", -- 0x0658
    x"CD",x"7A",x"06",x"3A",x"10",x"40",x"CB",x"57", -- 0x0660
    x"C0",x"AF",x"32",x"0C",x"40",x"3E",x"04",x"32", -- 0x0668
    x"10",x"40",x"AF",x"32",x"03",x"40",x"CD",x"EC", -- 0x0670
    x"0B",x"C9",x"CD",x"F9",x"05",x"CD",x"12",x"06", -- 0x0678
    x"11",x"66",x"0C",x"E7",x"C9",x"CD",x"3C",x"06", -- 0x0680
    x"3A",x"10",x"40",x"47",x"E6",x"18",x"5F",x"3A", -- 0x0688
    x"06",x"40",x"4F",x"3A",x"07",x"40",x"81",x"B7", -- 0x0690
    x"C8",x"3A",x"0F",x"00",x"B7",x"20",x"08",x"3A", -- 0x0698
    x"06",x"40",x"B7",x"20",x"02",x"18",x"0C",x"3A", -- 0x06A0
    x"00",x"68",x"E6",x"C0",x"FE",x"C0",x"28",x"7C", -- 0x06A8
    x"B7",x"28",x"70",x"7B",x"B7",x"3A",x"07",x"40", -- 0x06B0
    x"20",x"05",x"FE",x"01",x"CC",x"33",x"07",x"FE", -- 0x06B8
    x"02",x"20",x"0A",x"79",x"3C",x"27",x"32",x"06", -- 0x06C0
    x"40",x"AF",x"32",x"07",x"40",x"3A",x"2F",x"40", -- 0x06C8
    x"B7",x"C0",x"3A",x"06",x"40",x"FE",x"01",x"28", -- 0x06D0
    x"68",x"FE",x"02",x"D4",x"59",x"07",x"21",x"40", -- 0x06D8
    x"40",x"AF",x"06",x"14",x"D7",x"11",x"38",x"04", -- 0x06E0
    x"E7",x"11",x"9C",x"04",x"E7",x"3E",x"2B",x"32", -- 0x06E8
    x"9E",x"53",x"11",x"32",x"04",x"EF",x"3A",x"00", -- 0x06F0
    x"40",x"CB",x"5F",x"28",x"18",x"21",x"0F",x"43", -- 0x06F8
    x"06",x"10",x"34",x"23",x"23",x"10",x"FB",x"CD", -- 0x0700
    x"EC",x"0B",x"CD",x"84",x"07",x"3A",x"00",x"60", -- 0x0708
    x"CB",x"67",x"C2",x"15",x"07",x"3E",x"01",x"31", -- 0x0710
    x"00",x"44",x"32",x"01",x"70",x"AF",x"32",x"04", -- 0x0718
    x"70",x"18",x"FE",x"3A",x"07",x"40",x"FE",x"01", -- 0x0720
    x"28",x"99",x"18",x"A1",x"3E",x"04",x"32",x"06", -- 0x0728
    x"40",x"18",x"9A",x"CB",x"48",x"C0",x"3A",x"2F", -- 0x0730
    x"40",x"B7",x"20",x"18",x"11",x"78",x"04",x"18", -- 0x0738
    x"12",x"11",x"42",x"04",x"3A",x"00",x"68",x"CB", -- 0x0740
    x"47",x"28",x"05",x"3E",x"40",x"32",x"13",x"40", -- 0x0748
    x"E7",x"18",x"8B",x"E7",x"AF",x"32",x"04",x"70", -- 0x0750
    x"C9",x"11",x"5B",x"04",x"3A",x"00",x"68",x"CB", -- 0x0758
    x"47",x"20",x"E8",x"CB",x"4F",x"28",x"EC",x"3E", -- 0x0760
    x"C0",x"32",x"13",x"40",x"18",x"E5",x"FD",x"21", -- 0x0768
    x"50",x"40",x"FD",x"36",x"00",x"10",x"FD",x"36", -- 0x0770
    x"01",x"E0",x"FD",x"36",x"05",x"0D",x"3E",x"26", -- 0x0778
    x"32",x"44",x"40",x"C9",x"3A",x"00",x"70",x"E6", -- 0x0780
    x"03",x"C6",x"01",x"32",x"09",x"41",x"32",x"09", -- 0x0788
    x"42",x"C9",x"CD",x"E2",x"07",x"3A",x"43",x"40", -- 0x0790
    x"32",x"7D",x"43",x"32",x"79",x"43",x"3A",x"44", -- 0x0798
    x"40",x"4F",x"3A",x"0F",x"40",x"B7",x"28",x"03", -- 0x07A0
    x"79",x"2F",x"4F",x"79",x"32",x"7F",x"43",x"D6", -- 0x07A8
    x"05",x"32",x"7B",x"43",x"CD",x"00",x"0D",x"C9", -- 0x07B0
    x"3A",x"10",x"40",x"E6",x"18",x"C8",x"CB",x"5F", -- 0x07B8
    x"28",x"05",x"21",x"09",x"41",x"18",x"03",x"21", -- 0x07C0
    x"09",x"42",x"7E",x"3D",x"B7",x"C8",x"47",x"21", -- 0x07C8
    x"DF",x"50",x"11",x"E0",x"FF",x"36",x"FC",x"19", -- 0x07D0
    x"10",x"FB",x"C9",x"21",x"00",x"00",x"22",x"43", -- 0x07D8
    x"40",x"C9",x"FD",x"21",x"43",x"40",x"CD",x"A6", -- 0x07E0
    x"08",x"3A",x"42",x"40",x"FE",x"FA",x"20",x"06", -- 0x07E8
    x"F5",x"AF",x"32",x"05",x"68",x"F1",x"B7",x"28", -- 0x07F0
    x"04",x"3C",x"32",x"42",x"40",x"3A",x"10",x"40", -- 0x07F8
    x"CB",x"4F",x"20",x"D7",x"CD",x"0D",x"09",x"3A", -- 0x0800
    x"50",x"40",x"B7",x"C8",x"3A",x"41",x"40",x"B7", -- 0x0808
    x"20",x"4E",x"3A",x"10",x"40",x"5F",x"3A",x"0F", -- 0x0810
    x"40",x"57",x"CB",x"53",x"C2",x"9F",x"08",x"3A", -- 0x0818
    x"42",x"40",x"B7",x"20",x"14",x"7A",x"B7",x"20", -- 0x0820
    x"05",x"3A",x"00",x"60",x"18",x"07",x"CB",x"63", -- 0x0828
    x"28",x"F7",x"3A",x"00",x"68",x"CB",x"67",x"20", -- 0x0830
    x"16",x"3A",x"50",x"40",x"C6",x"07",x"32",x"43", -- 0x0838
    x"40",x"3A",x"51",x"40",x"2F",x"D6",x"06",x"32", -- 0x0840
    x"44",x"40",x"AF",x"32",x"05",x"68",x"C9",x"3E", -- 0x0848
    x"01",x"32",x"41",x"40",x"32",x"05",x"68",x"CD", -- 0x0850
    x"75",x"08",x"3E",x"F8",x"32",x"42",x"40",x"C9", -- 0x0858
    x"3A",x"50",x"40",x"C6",x"07",x"32",x"43",x"40", -- 0x0860
    x"3A",x"44",x"40",x"FE",x"D8",x"30",x"2A",x"C6", -- 0x0868
    x"08",x"32",x"44",x"40",x"C9",x"3A",x"10",x"40", -- 0x0870
    x"CB",x"5F",x"28",x"06",x"FD",x"21",x"00",x"41", -- 0x0878
    x"18",x"04",x"FD",x"21",x"00",x"42",x"FD",x"34", -- 0x0880
    x"04",x"11",x"B7",x"0C",x"1A",x"FD",x"BE",x"04", -- 0x0888
    x"C0",x"FD",x"36",x"04",x"00",x"FD",x"34",x"0A", -- 0x0890
    x"C9",x"AF",x"32",x"41",x"40",x"18",x"9A",x"3E", -- 0x0898
    x"01",x"32",x"41",x"40",x"18",x"93",x"E5",x"D5", -- 0x08A0
    x"FD",x"7E",x"00",x"2F",x"CB",x"3F",x"CB",x"3F", -- 0x08A8
    x"CB",x"3F",x"FD",x"77",x"02",x"FD",x"7E",x"01", -- 0x08B0
    x"2F",x"CB",x"3F",x"CB",x"3F",x"CB",x"3F",x"FD", -- 0x08B8
    x"77",x"03",x"21",x"00",x"00",x"11",x"20",x"00", -- 0x08C0
    x"FD",x"7E",x"02",x"B7",x"28",x"04",x"19",x"3D", -- 0x08C8
    x"18",x"F9",x"11",x"00",x"50",x"FD",x"7E",x"03", -- 0x08D0
    x"5F",x"19",x"11",x"01",x"00",x"B7",x"ED",x"52", -- 0x08D8
    x"FD",x"75",x"04",x"FD",x"74",x"05",x"7E",x"FD", -- 0x08E0
    x"77",x"06",x"B7",x"D1",x"E1",x"C9",x"3A",x"00", -- 0x08E8
    x"40",x"4F",x"DD",x"7E",x"05",x"E6",x"3E",x"57", -- 0x08F0
    x"DD",x"36",x"05",x"0E",x"CD",x"11",x"0A",x"DD", -- 0x08F8
    x"36",x"04",x"00",x"C3",x"83",x"09",x"3E",x"01", -- 0x0900
    x"32",x"1D",x"40",x"18",x"35",x"CD",x"70",x"0B", -- 0x0908
    x"CD",x"91",x"0A",x"3A",x"41",x"40",x"B7",x"C8", -- 0x0910
    x"FD",x"21",x"43",x"40",x"CD",x"A6",x"08",x"DD", -- 0x0918
    x"21",x"56",x"40",x"06",x"07",x"C5",x"DD",x"66", -- 0x0920
    x"03",x"DD",x"6E",x"02",x"DD",x"7E",x"05",x"E6", -- 0x0928
    x"3E",x"FE",x"10",x"38",x"58",x"FE",x"16",x"38", -- 0x0930
    x"CD",x"DD",x"7E",x"04",x"E6",x"3F",x"FE",x"18", -- 0x0938
    x"38",x"4B",x"DD",x"7E",x"01",x"4F",x"3A",x"0F", -- 0x0940
    x"40",x"B7",x"FD",x"7E",x"01",x"20",x"01",x"2F", -- 0x0948
    x"C6",x"04",x"91",x"FE",x"18",x"30",x"36",x"DD", -- 0x0950
    x"4E",x"00",x"3A",x"50",x"40",x"D6",x"08",x"91", -- 0x0958
    x"C6",x"06",x"FE",x"0C",x"30",x"27",x"CD",x"99", -- 0x0960
    x"08",x"CD",x"A6",x"08",x"3A",x"1D",x"40",x"B7", -- 0x0968
    x"C2",x"EE",x"08",x"DD",x"7E",x"05",x"E6",x"80", -- 0x0970
    x"4F",x"CD",x"58",x"00",x"E5",x"16",x"50",x"CD", -- 0x0978
    x"11",x"0A",x"E1",x"3E",x"01",x"32",x"1C",x"40", -- 0x0980
    x"3E",x"F0",x"32",x"03",x"40",x"AF",x"32",x"1D", -- 0x0988
    x"40",x"C1",x"11",x"06",x"00",x"DD",x"19",x"10", -- 0x0990
    x"8C",x"2A",x"47",x"40",x"7E",x"FE",x"10",x"20", -- 0x0998
    x"05",x"2B",x"7E",x"FE",x"10",x"C8",x"57",x"D5", -- 0x09A0
    x"FE",x"30",x"28",x"3F",x"FE",x"2C",x"28",x"3B", -- 0x09A8
    x"FE",x"F8",x"28",x"37",x"3D",x"77",x"3E",x"01", -- 0x09B0
    x"32",x"1C",x"40",x"3E",x"FC",x"32",x"03",x"40", -- 0x09B8
    x"FD",x"7E",x"00",x"D6",x"08",x"67",x"3A",x"0F", -- 0x09C0
    x"40",x"B7",x"FD",x"7E",x"01",x"20",x"01",x"2F", -- 0x09C8
    x"D6",x"18",x"6F",x"0E",x"0E",x"CD",x"46",x"0B", -- 0x09D0
    x"CD",x"99",x"08",x"D1",x"7A",x"E6",x"FC",x"FE", -- 0x09D8
    x"F8",x"28",x"04",x"CD",x"15",x"0A",x"C9",x"CD", -- 0x09E0
    x"11",x"0A",x"C9",x"36",x"10",x"18",x"C7",x"DD", -- 0x09E8
    x"E5",x"DD",x"21",x"87",x"0C",x"DD",x"7E",x"00", -- 0x09F0
    x"BA",x"20",x"07",x"DD",x"7E",x"01",x"DD",x"E1", -- 0x09F8
    x"C9",x"C9",x"DD",x"23",x"DD",x"23",x"18",x"ED", -- 0x0A00
    x"3A",x"14",x"40",x"0E",x"00",x"FD",x"E5",x"18", -- 0x0A08
    x"0B",x"0E",x"01",x"18",x"02",x"0E",x"00",x"FD", -- 0x0A10
    x"E5",x"3A",x"10",x"40",x"E6",x"18",x"B7",x"28", -- 0x0A18
    x"4B",x"CB",x"5F",x"20",x"66",x"FD",x"21",x"00", -- 0x0A20
    x"42",x"CD",x"EF",x"09",x"CB",x"41",x"20",x"0D", -- 0x0A28
    x"32",x"A8",x"40",x"32",x"39",x"40",x"5F",x"AF", -- 0x0A30
    x"32",x"38",x"40",x"18",x"0D",x"32",x"38",x"40", -- 0x0A38
    x"32",x"A9",x"40",x"5F",x"AF",x"32",x"39",x"40", -- 0x0A40
    x"18",x"34",x"FD",x"7E",x"02",x"B7",x"83",x"27", -- 0x0A48
    x"FD",x"77",x"02",x"30",x"17",x"FD",x"7E",x"01", -- 0x0A50
    x"B7",x"3C",x"27",x"FD",x"77",x"01",x"30",x"0C", -- 0x0A58
    x"FD",x"7E",x"00",x"3C",x"B7",x"27",x"FD",x"77", -- 0x0A60
    x"00",x"FD",x"34",x"0A",x"FD",x"E1",x"3A",x"10", -- 0x0A68
    x"40",x"E6",x"18",x"B7",x"C8",x"11",x"BE",x"0C", -- 0x0A70
    x"E7",x"11",x"B8",x"0C",x"EF",x"C9",x"FD",x"7E", -- 0x0A78
    x"01",x"B7",x"83",x"27",x"FD",x"77",x"01",x"30", -- 0x0A80
    x"E3",x"18",x"D5",x"FD",x"21",x"00",x"41",x"18", -- 0x0A88
    x"98",x"E5",x"D5",x"C5",x"FD",x"7E",x"05",x"DD", -- 0x0A90
    x"77",x"01",x"FD",x"7E",x"00",x"DD",x"77",x"00", -- 0x0A98
    x"C6",x"10",x"2F",x"CB",x"3F",x"CB",x"3F",x"CB", -- 0x0AA0
    x"3F",x"4F",x"FD",x"7E",x"01",x"DD",x"77",x"03", -- 0x0AA8
    x"C6",x"08",x"CB",x"3F",x"CB",x"3F",x"CB",x"3F", -- 0x0AB0
    x"47",x"21",x"00",x"00",x"11",x"20",x"00",x"79", -- 0x0AB8
    x"B7",x"28",x"04",x"19",x"3D",x"18",x"F9",x"11", -- 0x0AC0
    x"00",x"50",x"78",x"5F",x"19",x"11",x"01",x"00", -- 0x0AC8
    x"B7",x"ED",x"52",x"FD",x"75",x"02",x"FD",x"74", -- 0x0AD0
    x"03",x"C1",x"D1",x"E1",x"C9",x"DD",x"21",x"40", -- 0x0AD8
    x"43",x"11",x"04",x"00",x"FD",x"21",x"50",x"40", -- 0x0AE0
    x"06",x"08",x"CD",x"91",x"0A",x"FD",x"19",x"DD", -- 0x0AE8
    x"19",x"FD",x"23",x"FD",x"23",x"10",x"F3",x"C9", -- 0x0AF0
    x"DD",x"E5",x"FD",x"E5",x"E5",x"C5",x"F5",x"21", -- 0x0AF8
    x"56",x"40",x"06",x"23",x"AF",x"D7",x"3A",x"05", -- 0x0B00
    x"40",x"FE",x"30",x"38",x"04",x"FE",x"D0",x"38", -- 0x0B08
    x"02",x"3E",x"80",x"67",x"2E",x"00",x"DD",x"21", -- 0x0B10
    x"40",x"0B",x"DD",x"4E",x"00",x"06",x"06",x"CD", -- 0x0B18
    x"46",x"0B",x"DD",x"7E",x"00",x"FD",x"77",x"04", -- 0x0B20
    x"FD",x"77",x"05",x"DD",x"23",x"7C",x"C6",x"10", -- 0x0B28
    x"67",x"10",x"EC",x"3A",x"10",x"40",x"CB",x"C7", -- 0x0B30
    x"F1",x"C1",x"E1",x"FD",x"E1",x"DD",x"E1",x"C9", -- 0x0B38
    x"18",x"1C",x"1C",x"1C",x"1C",x"20",x"C5",x"06", -- 0x0B40
    x"07",x"FD",x"21",x"56",x"40",x"11",x"06",x"00", -- 0x0B48
    x"FD",x"7E",x"00",x"B7",x"20",x"13",x"FD",x"7E", -- 0x0B50
    x"05",x"B7",x"20",x"0D",x"FD",x"74",x"00",x"FD", -- 0x0B58
    x"75",x"01",x"FD",x"71",x"05",x"C1",x"3E",x"01", -- 0x0B60
    x"C9",x"FD",x"19",x"10",x"E3",x"AF",x"C1",x"C9", -- 0x0B68
    x"FD",x"21",x"50",x"40",x"06",x"08",x"11",x"06", -- 0x0B70
    x"00",x"FD",x"7E",x"00",x"B7",x"28",x"30",x"FD", -- 0x0B78
    x"7E",x"05",x"E6",x"FE",x"FE",x"0E",x"20",x"27", -- 0x0B80
    x"FE",x"3C",x"28",x"28",x"3A",x"03",x"40",x"B7", -- 0x0B88
    x"20",x"0F",x"AF",x"FD",x"77",x"00",x"FD",x"77", -- 0x0B90
    x"01",x"FD",x"77",x"05",x"32",x"1C",x"40",x"18", -- 0x0B98
    x"0E",x"FE",x"FC",x"30",x"06",x"FD",x"36",x"05", -- 0x0BA0
    x"0E",x"18",x"04",x"FD",x"36",x"05",x"0F",x"FD", -- 0x0BA8
    x"19",x"10",x"C6",x"C9",x"3A",x"03",x"40",x"FE", -- 0x0BB0
    x"E8",x"20",x"F4",x"FD",x"36",x"05",x"3D",x"18", -- 0x0BB8
    x"EE",x"3A",x"00",x"40",x"4F",x"3A",x"14",x"40", -- 0x0BC0
    x"E6",x"1C",x"B7",x"C8",x"CB",x"57",x"20",x"1C", -- 0x0BC8
    x"CB",x"5F",x"20",x"25",x"21",x"02",x"42",x"79", -- 0x0BD0
    x"CB",x"61",x"20",x"10",x"11",x"5C",x"0C",x"E7", -- 0x0BD8
    x"11",x"66",x"0C",x"E7",x"CD",x"0F",x"0C",x"CD", -- 0x0BE0
    x"B8",x"07",x"C9",x"C9",x"11",x"20",x"04",x"EF", -- 0x0BE8
    x"11",x"26",x"04",x"EF",x"11",x"2C",x"04",x"EF", -- 0x0BF0
    x"C9",x"21",x"02",x"41",x"CB",x"61",x"20",x"EC", -- 0x0BF8
    x"11",x"52",x"0C",x"E7",x"11",x"66",x"0C",x"E7", -- 0x0C00
    x"CD",x"0F",x"0C",x"CD",x"B8",x"07",x"C9",x"3A", -- 0x0C08
    x"10",x"40",x"CB",x"5F",x"28",x"06",x"DD",x"21", -- 0x0C10
    x"00",x"41",x"18",x"04",x"DD",x"21",x"00",x"42", -- 0x0C18
    x"3A",x"34",x"40",x"06",x"03",x"DD",x"BE",x"00", -- 0x0C20
    x"38",x"16",x"05",x"3A",x"35",x"40",x"DD",x"BE", -- 0x0C28
    x"01",x"38",x"0D",x"05",x"3A",x"36",x"40",x"DD", -- 0x0C30
    x"BE",x"02",x"38",x"04",x"CD",x"F9",x"00",x"C9", -- 0x0C38
    x"DD",x"E5",x"E1",x"23",x"23",x"11",x"36",x"40", -- 0x0C40
    x"7E",x"12",x"2B",x"1B",x"10",x"FA",x"CD",x"F9", -- 0x0C48
    x"00",x"C9",x"05",x"01",x"00",x"40",x"40",x"40", -- 0x0C50
    x"40",x"40",x"40",x"FF",x"05",x"01",x"16",x"40", -- 0x0C58
    x"40",x"40",x"40",x"40",x"40",x"FF",x"07",x"1F", -- 0x0C60
    x"16",x"40",x"40",x"40",x"40",x"40",x"40",x"FF", -- 0x0C68
    x"AB",x"3A",x"14",x"40",x"E6",x"18",x"C8",x"1E", -- 0x0C70
    x"01",x"CB",x"5F",x"28",x"05",x"DD",x"21",x"00", -- 0x0C78
    x"41",x"C9",x"DD",x"21",x"00",x"42",x"C9",x"32", -- 0x0C80
    x"40",x"31",x"30",x"30",x"20",x"2F",x"40",x"2E", -- 0x0C88
    x"80",x"2D",x"60",x"2C",x"40",x"F8",x"09",x"F9", -- 0x0C90
    x"09",x"FA",x"09",x"FB",x"09",x"00",x"00",x"00", -- 0x0C98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0CA0
    x"00",x"50",x"01",x"10",x"02",x"11",x"04",x"12", -- 0x0CA8
    x"06",x"13",x"06",x"14",x"50",x"15",x"50",x"60", -- 0x0CB0
    x"07",x"1F",x"0C",x"38",x"40",x"04",x"07",x"1F", -- 0x0CB8
    x"02",x"48",x"49",x"54",x"40",x"56",x"41",x"4C", -- 0x0CC0
    x"55",x"45",x"FF",x"2A",x"00",x"40",x"23",x"22", -- 0x0CC8
    x"00",x"40",x"3A",x"10",x"40",x"B7",x"CC",x"EC", -- 0x0CD0
    x"0B",x"C9",x"04",x"32",x"01",x"40",x"C9",x"CB", -- 0x0CD8
    x"BF",x"18",x"F8",x"00",x"00",x"00",x"00",x"00", -- 0x0CE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0CE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0CF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0CF8
    x"FD",x"21",x"50",x"40",x"0E",x"FF",x"3A",x"10", -- 0x0D00
    x"40",x"47",x"E6",x"1C",x"B7",x"C8",x"CB",x"50", -- 0x0D08
    x"C2",x"CE",x"0D",x"0E",x"00",x"CB",x"58",x"28", -- 0x0D10
    x"05",x"CD",x"80",x"0D",x"18",x"0E",x"3A",x"0F", -- 0x0D18
    x"40",x"B7",x"20",x"05",x"CD",x"80",x"0D",x"18", -- 0x0D20
    x"03",x"CD",x"A6",x"0D",x"79",x"CD",x"43",x"0D", -- 0x0D28
    x"CD",x"46",x"0E",x"CD",x"62",x"0D",x"3A",x"32", -- 0x0D30
    x"40",x"B7",x"20",x"03",x"CD",x"62",x"0D",x"FD", -- 0x0D38
    x"71",x"04",x"C9",x"FD",x"7E",x"00",x"FE",x"14", -- 0x0D40
    x"30",x"02",x"CB",x"A1",x"FE",x"E2",x"38",x"02", -- 0x0D48
    x"CB",x"99",x"FD",x"7E",x"01",x"FE",x"A0",x"30", -- 0x0D50
    x"02",x"CB",x"B1",x"FE",x"E6",x"38",x"02",x"CB", -- 0x0D58
    x"A9",x"C9",x"CB",x"59",x"28",x"05",x"FD",x"34", -- 0x0D60
    x"00",x"18",x"07",x"CB",x"61",x"28",x"03",x"FD", -- 0x0D68
    x"35",x"00",x"CB",x"69",x"28",x"03",x"FD",x"34", -- 0x0D70
    x"01",x"CB",x"71",x"C8",x"FD",x"35",x"01",x"C9", -- 0x0D78
    x"3A",x"00",x"60",x"CB",x"57",x"28",x"02",x"CB", -- 0x0D80
    x"E1",x"CB",x"5F",x"28",x"02",x"CB",x"D9",x"CB", -- 0x0D88
    x"77",x"28",x"02",x"CB",x"E9",x"CB",x"7F",x"28", -- 0x0D90
    x"02",x"CB",x"F1",x"79",x"B7",x"28",x"04",x"06", -- 0x0D98
    x"01",x"79",x"C9",x"06",x"00",x"C9",x"3A",x"00", -- 0x0DA0
    x"68",x"CB",x"57",x"28",x"02",x"CB",x"E1",x"CB", -- 0x0DA8
    x"5F",x"28",x"02",x"CB",x"D9",x"CB",x"6F",x"28", -- 0x0DB0
    x"02",x"CB",x"E9",x"3A",x"00",x"60",x"CB",x"4F", -- 0x0DB8
    x"28",x"02",x"CB",x"F1",x"79",x"B7",x"28",x"03", -- 0x0DC0
    x"06",x"01",x"C9",x"06",x"00",x"C9",x"FD",x"4E", -- 0x0DC8
    x"04",x"FD",x"7E",x"00",x"FE",x"0C",x"30",x"02", -- 0x0DD0
    x"CB",x"F1",x"FE",x"E0",x"38",x"02",x"CB",x"B1", -- 0x0DD8
    x"FD",x"7E",x"01",x"FE",x"80",x"30",x"02",x"CB", -- 0x0DE0
    x"E9",x"FE",x"E0",x"38",x"02",x"CB",x"A9",x"3A", -- 0x0DE8
    x"00",x"40",x"CB",x"77",x"28",x"12",x"CB",x"71", -- 0x0DF0
    x"28",x"08",x"FD",x"34",x"00",x"FD",x"34",x"00", -- 0x0DF8
    x"18",x"06",x"FD",x"35",x"00",x"FD",x"35",x"00", -- 0x0E00
    x"CB",x"69",x"28",x"05",x"FD",x"34",x"01",x"18", -- 0x0E08
    x"03",x"FD",x"35",x"01",x"FD",x"71",x"04",x"C9", -- 0x0E10
    x"C5",x"7D",x"E6",x"1F",x"47",x"AF",x"C6",x"08", -- 0x0E18
    x"10",x"FC",x"57",x"7D",x"E6",x"E0",x"CB",x"3F", -- 0x0E20
    x"CB",x"3F",x"CB",x"3F",x"CB",x"3F",x"CB",x"3F", -- 0x0E28
    x"4F",x"7C",x"E6",x"03",x"CB",x"27",x"CB",x"27", -- 0x0E30
    x"CB",x"27",x"B1",x"47",x"AF",x"D6",x"08",x"10", -- 0x0E38
    x"FC",x"D6",x"1C",x"5F",x"C1",x"C9",x"FD",x"66", -- 0x0E40
    x"03",x"FD",x"6E",x"02",x"E5",x"23",x"11",x"20", -- 0x0E48
    x"00",x"7E",x"FE",x"10",x"28",x"09",x"CD",x"DA", -- 0x0E50
    x"0E",x"C6",x"10",x"FE",x"08",x"38",x"11",x"23", -- 0x0E58
    x"7E",x"2B",x"FE",x"10",x"28",x"0C",x"23",x"CD", -- 0x0E60
    x"DA",x"0E",x"C6",x"10",x"FE",x"08",x"30",x"02", -- 0x0E68
    x"CB",x"99",x"11",x"40",x"00",x"19",x"7E",x"FE", -- 0x0E70
    x"10",x"28",x"07",x"CD",x"DA",x"0E",x"FE",x"E8", -- 0x0E78
    x"30",x"0F",x"23",x"7E",x"2B",x"FE",x"10",x"28", -- 0x0E80
    x"0A",x"23",x"CD",x"DA",x"0E",x"FE",x"E8",x"38", -- 0x0E88
    x"02",x"CB",x"A1",x"2B",x"7E",x"FE",x"10",x"28", -- 0x0E90
    x"09",x"CD",x"E2",x"0E",x"FE",x"FE",x"38",x"02", -- 0x0E98
    x"CB",x"B1",x"11",x"E0",x"FF",x"19",x"7E",x"FE", -- 0x0EA0
    x"10",x"28",x"09",x"CD",x"E2",x"0E",x"FE",x"FE", -- 0x0EA8
    x"38",x"02",x"CB",x"B1",x"E1",x"11",x"20",x"00", -- 0x0EB0
    x"19",x"23",x"23",x"7E",x"FE",x"10",x"28",x"09", -- 0x0EB8
    x"CD",x"E2",x"0E",x"FE",x"0C",x"30",x"02",x"CB", -- 0x0EC0
    x"A9",x"11",x"20",x"00",x"19",x"7E",x"FE",x"10", -- 0x0EC8
    x"C8",x"CD",x"E2",x"0E",x"FE",x"0C",x"D0",x"CB", -- 0x0ED0
    x"A9",x"C9",x"CD",x"18",x"0E",x"7B",x"FD",x"96", -- 0x0ED8
    x"00",x"C9",x"CD",x"18",x"0E",x"7A",x"FD",x"96", -- 0x0EE0
    x"01",x"ED",x"53",x"90",x"40",x"32",x"92",x"40", -- 0x0EE8
    x"C9",x"B1",x"E1",x"11",x"20",x"00",x"19",x"23", -- 0x0EF0
    x"23",x"7E",x"FE",x"10",x"28",x"09",x"CD",x"20", -- 0x0EF8
    x"0F",x"FE",x"0C",x"30",x"02",x"CB",x"A9",x"11", -- 0x0F00
    x"20",x"00",x"19",x"7E",x"FE",x"10",x"C8",x"CD", -- 0x0F08
    x"20",x"0F",x"FE",x"0C",x"D0",x"CB",x"A9",x"C9", -- 0x0F10
    x"CD",x"56",x"0E",x"7B",x"FD",x"96",x"00",x"C9", -- 0x0F18
    x"CD",x"56",x"0E",x"7A",x"FD",x"96",x"01",x"ED", -- 0x0F20
    x"53",x"90",x"40",x"32",x"92",x"40",x"C9",x"00", -- 0x0F28
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F30
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F38
    x"0F",x"FE",x"0C",x"30",x"02",x"CB",x"A9",x"11", -- 0x0F40
    x"20",x"00",x"19",x"7E",x"FE",x"10",x"C8",x"CD", -- 0x0F48
    x"20",x"0F",x"FE",x"0C",x"D0",x"CB",x"A9",x"C9", -- 0x0F50
    x"CD",x"56",x"0E",x"7B",x"FD",x"96",x"00",x"C9", -- 0x0F58
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F60
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F68
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F78
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F80
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F88
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F90
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0FA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0FA8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0FB0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0FB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0FC0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0FC8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0FD0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0FD8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0FE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0FE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0FF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0FF8
    x"CD",x"45",x"15",x"CD",x"98",x"13",x"AF",x"21", -- 0x1000
    x"A0",x"40",x"06",x"04",x"D7",x"32",x"0C",x"40", -- 0x1008
    x"3A",x"10",x"40",x"E6",x"1C",x"C8",x"FD",x"21", -- 0x1010
    x"56",x"40",x"06",x"07",x"FD",x"7E",x"05",x"4F", -- 0x1018
    x"E6",x"3E",x"FE",x"10",x"CA",x"00",x"26",x"FE", -- 0x1020
    x"14",x"CA",x"8E",x"26",x"FE",x"12",x"CA",x"0C", -- 0x1028
    x"27",x"79",x"E6",x"3F",x"FE",x"18",x"38",x"09", -- 0x1030
    x"FE",x"30",x"38",x"10",x"FE",x"38",x"DA",x"BF", -- 0x1038
    x"11",x"11",x"06",x"00",x"FD",x"19",x"10",x"D4", -- 0x1040
    x"CD",x"7F",x"15",x"C9",x"3A",x"0C",x"40",x"3C", -- 0x1048
    x"32",x"0C",x"40",x"FD",x"7E",x"04",x"E6",x"3F", -- 0x1050
    x"FE",x"18",x"CA",x"19",x"14",x"FE",x"24",x"CA", -- 0x1058
    x"19",x"14",x"FE",x"28",x"CA",x"19",x"14",x"FD", -- 0x1060
    x"7E",x"FF",x"E6",x"3F",x"FE",x"18",x"38",x"1E", -- 0x1068
    x"FE",x"30",x"30",x"1A",x"FD",x"7E",x"05",x"E6", -- 0x1070
    x"80",x"B7",x"FD",x"7E",x"FB",x"FD",x"77",x"01", -- 0x1078
    x"FD",x"7E",x"FA",x"20",x"04",x"C6",x"10",x"18", -- 0x1080
    x"02",x"D6",x"10",x"FD",x"77",x"00",x"FD",x"7E", -- 0x1088
    x"01",x"FE",x"A0",x"30",x"08",x"FD",x"7E",x"04", -- 0x1090
    x"CB",x"BF",x"FD",x"77",x"04",x"FD",x"7E",x"01", -- 0x1098
    x"FE",x"E8",x"38",x"0D",x"FD",x"7E",x"04",x"CB", -- 0x10A0
    x"FF",x"FD",x"77",x"04",x"3E",x"01",x"32",x"13", -- 0x10A8
    x"40",x"79",x"E6",x"80",x"B7",x"FD",x"7E",x"00", -- 0x10B0
    x"C2",x"6F",x"11",x"5F",x"FD",x"7E",x"04",x"E6", -- 0x10B8
    x"3F",x"FE",x"18",x"28",x"1E",x"FE",x"24",x"28", -- 0x10C0
    x"1A",x"FE",x"28",x"28",x"16",x"3A",x"16",x"40", -- 0x10C8
    x"B7",x"20",x"49",x"FD",x"7E",x"FB",x"FD",x"77", -- 0x10D0
    x"01",x"FD",x"7E",x"FA",x"C6",x"10",x"FD",x"77", -- 0x10D8
    x"00",x"18",x"21",x"3A",x"12",x"40",x"B7",x"C4", -- 0x10E0
    x"31",x"11",x"FD",x"7E",x"00",x"FE",x"18",x"DC", -- 0x10E8
    x"31",x"11",x"FD",x"66",x"03",x"FD",x"6E",x"02", -- 0x10F0
    x"11",x"40",x"00",x"19",x"7E",x"FE",x"10",x"C4", -- 0x10F8
    x"31",x"11",x"18",x"18",x"FD",x"7E",x"05",x"E6", -- 0x1100
    x"FC",x"4F",x"3A",x"00",x"40",x"E6",x"18",x"CB", -- 0x1108
    x"3F",x"CB",x"3F",x"CB",x"3F",x"B1",x"FD",x"77", -- 0x1110
    x"05",x"C3",x"36",x"13",x"FD",x"35",x"00",x"FD", -- 0x1118
    x"35",x"00",x"18",x"E0",x"3E",x"01",x"32",x"16", -- 0x1120
    x"40",x"18",x"1C",x"AF",x"32",x"16",x"40",x"18", -- 0x1128
    x"16",x"FD",x"7E",x"04",x"5F",x"E6",x"3C",x"FE", -- 0x1130
    x"18",x"28",x"E9",x"FE",x"28",x"28",x"E5",x"FE", -- 0x1138
    x"20",x"28",x"E8",x"FE",x"2C",x"28",x"E4",x"7B", -- 0x1140
    x"E6",x"80",x"57",x"FD",x"7E",x"05",x"E6",x"80", -- 0x1148
    x"4F",x"7B",x"E6",x"7F",x"CB",x"7A",x"20",x"08", -- 0x1150
    x"CD",x"1C",x"12",x"B1",x"FD",x"77",x"05",x"C9", -- 0x1158
    x"CD",x"16",x"12",x"F5",x"FD",x"7E",x"01",x"D6", -- 0x1160
    x"08",x"FD",x"77",x"01",x"F1",x"18",x"EC",x"5F", -- 0x1168
    x"FD",x"7E",x"04",x"E6",x"3F",x"FE",x"18",x"28", -- 0x1170
    x"1F",x"FE",x"24",x"28",x"1B",x"FE",x"28",x"28", -- 0x1178
    x"17",x"3A",x"16",x"40",x"B7",x"20",x"2C",x"FD", -- 0x1180
    x"7E",x"FB",x"FD",x"77",x"01",x"FD",x"7E",x"FA", -- 0x1188
    x"D6",x"10",x"FD",x"77",x"00",x"C3",x"04",x"11", -- 0x1190
    x"3A",x"12",x"40",x"B7",x"C4",x"31",x"11",x"FD", -- 0x1198
    x"7E",x"00",x"FE",x"D8",x"D4",x"31",x"11",x"FD", -- 0x11A0
    x"66",x"03",x"FD",x"6E",x"02",x"7E",x"FE",x"10", -- 0x11A8
    x"C4",x"31",x"11",x"FD",x"34",x"00",x"FD",x"34", -- 0x11B0
    x"00",x"FD",x"7E",x"00",x"C3",x"04",x"11",x"3A", -- 0x11B8
    x"0C",x"40",x"3C",x"32",x"0C",x"40",x"3A",x"00", -- 0x11C0
    x"40",x"E6",x"02",x"6F",x"FD",x"7E",x"04",x"E6", -- 0x11C8
    x"80",x"B7",x"20",x"21",x"FD",x"7E",x"05",x"4F", -- 0x11D0
    x"E6",x"80",x"5F",x"79",x"E6",x"3F",x"FE",x"33", -- 0x11D8
    x"CA",x"64",x"12",x"FE",x"37",x"D2",x"64",x"12", -- 0x11E0
    x"CB",x"4D",x"CA",x"41",x"10",x"3C",x"B3",x"FD", -- 0x11E8
    x"77",x"05",x"C3",x"41",x"10",x"FD",x"7E",x"05", -- 0x11F0
    x"4F",x"E6",x"C0",x"5F",x"79",x"E6",x"3F",x"FE", -- 0x11F8
    x"30",x"CA",x"64",x"12",x"FE",x"34",x"CA",x"64", -- 0x1200
    x"12",x"CB",x"4D",x"CA",x"41",x"10",x"3D",x"B3", -- 0x1208
    x"FD",x"77",x"05",x"C3",x"41",x"10",x"DD",x"21", -- 0x1210
    x"44",x"12",x"18",x"04",x"DD",x"21",x"36",x"12", -- 0x1218
    x"C5",x"06",x"07",x"E6",x"FC",x"DD",x"BE",x"00", -- 0x1220
    x"28",x"07",x"DD",x"23",x"DD",x"23",x"10",x"F5", -- 0x1228
    x"C9",x"DD",x"7E",x"01",x"C1",x"C9",x"18",x"30", -- 0x1230
    x"1C",x"34",x"20",x"34",x"24",x"30",x"28",x"30", -- 0x1238
    x"2C",x"30",x"00",x"00",x"18",x"73",x"1C",x"77", -- 0x1240
    x"20",x"77",x"24",x"73",x"28",x"77",x"2C",x"77", -- 0x1248
    x"00",x"00",x"FD",x"7E",x"04",x"CB",x"FF",x"FD", -- 0x1250
    x"77",x"04",x"C9",x"FD",x"7E",x"04",x"CB",x"BF", -- 0x1258
    x"FD",x"77",x"04",x"C9",x"FD",x"7E",x"05",x"E6", -- 0x1260
    x"3F",x"FE",x"18",x"CC",x"52",x"12",x"FE",x"24", -- 0x1268
    x"CC",x"52",x"12",x"FE",x"28",x"CC",x"52",x"12", -- 0x1270
    x"FE",x"37",x"CC",x"5B",x"12",x"FE",x"33",x"CC", -- 0x1278
    x"5B",x"12",x"FD",x"7E",x"0A",x"E6",x"3F",x"FE", -- 0x1280
    x"19",x"38",x"18",x"FE",x"24",x"28",x"14",x"FE", -- 0x1288
    x"28",x"28",x"10",x"FE",x"38",x"30",x"0C",x"FD", -- 0x1290
    x"7E",x"00",x"FD",x"77",x"06",x"FD",x"7E",x"01", -- 0x1298
    x"FD",x"77",x"07",x"FD",x"7E",x"04",x"5F",x"E6", -- 0x12A0
    x"80",x"57",x"FD",x"7E",x"05",x"E6",x"80",x"4F", -- 0x12A8
    x"FD",x"7E",x"04",x"E6",x"3F",x"FE",x"18",x"28", -- 0x12B0
    x"0A",x"FE",x"24",x"28",x"06",x"FE",x"28",x"28", -- 0x12B8
    x"02",x"18",x"0C",x"FD",x"7E",x"00",x"32",x"1E", -- 0x12C0
    x"40",x"FD",x"7E",x"01",x"32",x"1F",x"40",x"FD", -- 0x12C8
    x"7E",x"0A",x"E6",x"3F",x"FE",x"19",x"38",x"2D", -- 0x12D0
    x"FE",x"24",x"28",x"29",x"FE",x"28",x"28",x"25", -- 0x12D8
    x"FE",x"38",x"30",x"21",x"3A",x"1E",x"40",x"FD", -- 0x12E0
    x"77",x"06",x"3A",x"1F",x"40",x"FD",x"77",x"07", -- 0x12E8
    x"FD",x"7E",x"0A",x"E6",x"3F",x"CB",x"7A",x"28", -- 0x12F0
    x"05",x"CD",x"16",x"12",x"18",x"03",x"CD",x"1C", -- 0x12F8
    x"12",x"B1",x"FD",x"77",x"0B",x"3A",x"12",x"40", -- 0x1300
    x"B7",x"20",x"1A",x"FD",x"7E",x"04",x"E6",x"3F", -- 0x1308
    x"B1",x"EE",x"80",x"FD",x"77",x"05",x"3A",x"1F", -- 0x1310
    x"40",x"CB",x"7A",x"20",x"02",x"C6",x"08",x"FD", -- 0x1318
    x"77",x"01",x"C3",x"41",x"10",x"FD",x"7E",x"05", -- 0x1320
    x"E6",x"3F",x"CB",x"7A",x"20",x"05",x"CD",x"1C", -- 0x1328
    x"12",x"18",x"DD",x"CD",x"16",x"12",x"FD",x"7E", -- 0x1330
    x"05",x"E6",x"3F",x"FE",x"18",x"CA",x"4B",x"13", -- 0x1338
    x"FE",x"24",x"28",x"07",x"FE",x"28",x"28",x"03", -- 0x1340
    x"C3",x"41",x"10",x"D9",x"DD",x"21",x"50",x"40", -- 0x1348
    x"06",x"08",x"DD",x"7E",x"05",x"E6",x"3C",x"FE", -- 0x1350
    x"18",x"28",x"0A",x"FE",x"24",x"28",x"06",x"FE", -- 0x1358
    x"28",x"28",x"02",x"18",x"28",x"DD",x"E5",x"E1", -- 0x1360
    x"FD",x"E5",x"D1",x"B7",x"ED",x"52",x"28",x"1D", -- 0x1368
    x"FD",x"66",x"01",x"FD",x"6E",x"00",x"DD",x"56", -- 0x1370
    x"01",x"DD",x"5E",x"00",x"B7",x"ED",x"52",x"20", -- 0x1378
    x"0C",x"FD",x"7E",x"05",x"E6",x"80",x"4F",x"3E", -- 0x1380
    x"30",x"A9",x"FD",x"77",x"05",x"11",x"08",x"00", -- 0x1388
    x"DD",x"19",x"10",x"BE",x"D9",x"C3",x"41",x"10", -- 0x1390
    x"3A",x"10",x"40",x"E6",x"1C",x"C8",x"CB",x"4F", -- 0x1398
    x"C0",x"FD",x"21",x"50",x"40",x"FD",x"7E",x"00", -- 0x13A0
    x"FE",x"10",x"D8",x"DD",x"21",x"56",x"40",x"11", -- 0x13A8
    x"06",x"00",x"06",x"07",x"DD",x"7E",x"05",x"E6", -- 0x13B0
    x"3F",x"FE",x"10",x"38",x"27",x"FE",x"16",x"38", -- 0x13B8
    x"0D",x"DD",x"7E",x"04",x"E6",x"3F",x"FE",x"18", -- 0x13C0
    x"38",x"1A",x"FE",x"3C",x"30",x"16",x"DD",x"7E", -- 0x13C8
    x"00",x"B7",x"28",x"10",x"FD",x"7E",x"00",x"D6", -- 0x13D0
    x"04",x"4F",x"DD",x"7E",x"00",x"91",x"C6",x"08", -- 0x13D8
    x"FE",x"10",x"38",x"08",x"11",x"06",x"00",x"DD", -- 0x13E0
    x"19",x"10",x"C9",x"C9",x"DD",x"7E",x"01",x"4F", -- 0x13E8
    x"FD",x"7E",x"01",x"C6",x"04",x"91",x"C6",x"08", -- 0x13F0
    x"FE",x"10",x"30",x"E8",x"3A",x"10",x"40",x"32", -- 0x13F8
    x"14",x"40",x"3E",x"01",x"32",x"1C",x"40",x"3E", -- 0x1400
    x"02",x"32",x"10",x"40",x"3E",x"E0",x"32",x"03", -- 0x1408
    x"40",x"3E",x"3D",x"FD",x"77",x"05",x"C3",x"B5", -- 0x1410
    x"17",x"FD",x"E5",x"DD",x"E5",x"D9",x"FD",x"E5", -- 0x1418
    x"DD",x"E1",x"3E",x"01",x"32",x"09",x"40",x"11", -- 0x1420
    x"06",x"00",x"DD",x"19",x"DD",x"7E",x"05",x"E6", -- 0x1428
    x"3F",x"FE",x"18",x"38",x"15",x"FE",x"30",x"30", -- 0x1430
    x"11",x"FD",x"6E",x"02",x"FD",x"66",x"03",x"DD", -- 0x1438
    x"5E",x"02",x"DD",x"56",x"03",x"B7",x"ED",x"52", -- 0x1440
    x"28",x"12",x"DD",x"E5",x"D1",x"21",x"7F",x"40", -- 0x1448
    x"ED",x"52",x"30",x"D3",x"D9",x"DD",x"E1",x"FD", -- 0x1450
    x"E1",x"C3",x"8E",x"10",x"FD",x"7E",x"05",x"E6", -- 0x1458
    x"80",x"EE",x"80",x"C6",x"30",x"FD",x"77",x"05", -- 0x1460
    x"18",x"E0",x"3A",x"13",x"40",x"CB",x"77",x"C8", -- 0x1468
    x"CB",x"B7",x"32",x"13",x"40",x"AF",x"32",x"10", -- 0x1470
    x"40",x"3E",x"01",x"32",x"2F",x"40",x"32",x"01", -- 0x1478
    x"70",x"31",x"00",x"44",x"AF",x"21",x"00",x"60", -- 0x1480
    x"06",x"00",x"D7",x"21",x"00",x"68",x"D7",x"21", -- 0x1488
    x"00",x"00",x"22",x"06",x"70",x"21",x"16",x"1F", -- 0x1490
    x"22",x"05",x"41",x"22",x"05",x"42",x"3E",x"01", -- 0x1498
    x"32",x"08",x"41",x"CD",x"49",x"00",x"3A",x"13", -- 0x14A0
    x"40",x"CB",x"7F",x"3A",x"06",x"40",x"20",x"0C", -- 0x14A8
    x"3D",x"27",x"32",x"06",x"40",x"3E",x"08",x"32", -- 0x14B0
    x"14",x"40",x"18",x"0B",x"3D",x"3D",x"27",x"32", -- 0x14B8
    x"06",x"40",x"3E",x"88",x"32",x"14",x"40",x"3A", -- 0x14C0
    x"13",x"40",x"3E",x"C0",x"CD",x"4C",x"00",x"11", -- 0x14C8
    x"00",x"01",x"E7",x"3E",x"80",x"CD",x"4C",x"00", -- 0x14D0
    x"CD",x"49",x"00",x"21",x"50",x"40",x"06",x"30", -- 0x14D8
    x"AF",x"D7",x"21",x"00",x"41",x"CD",x"61",x"27", -- 0x14E0
    x"21",x"00",x"42",x"CD",x"61",x"27",x"AF",x"32", -- 0x14E8
    x"0A",x"41",x"32",x"0A",x"42",x"3A",x"10",x"40", -- 0x14F0
    x"CB",x"C7",x"32",x"10",x"40",x"3E",x"80",x"CD", -- 0x14F8
    x"4C",x"00",x"CD",x"4F",x"00",x"3A",x"14",x"40", -- 0x1500
    x"32",x"10",x"40",x"3E",x"01",x"32",x"04",x"70", -- 0x1508
    x"3A",x"10",x"40",x"CB",x"47",x"20",x"23",x"21", -- 0x1510
    x"40",x"50",x"11",x"00",x"00",x"7E",x"E6",x"FC", -- 0x1518
    x"FE",x"30",x"20",x"01",x"1C",x"23",x"7C",x"FE", -- 0x1520
    x"54",x"20",x"F2",x"7B",x"32",x"0A",x"40",x"B7", -- 0x1528
    x"20",x"08",x"3A",x"10",x"40",x"CB",x"C7",x"32", -- 0x1530
    x"10",x"40",x"CD",x"F3",x"00",x"CD",x"98",x"13", -- 0x1538
    x"CD",x"E0",x"00",x"18",x"CB",x"3A",x"0C",x"40", -- 0x1540
    x"B7",x"C0",x"3A",x"10",x"40",x"E6",x"1C",x"B7", -- 0x1548
    x"C8",x"21",x"A0",x"40",x"7E",x"4F",x"23",x"7E", -- 0x1550
    x"81",x"4F",x"23",x"7E",x"81",x"B7",x"C0",x"3E", -- 0x1558
    x"FF",x"32",x"00",x"78",x"CD",x"5E",x"00",x"CD", -- 0x1560
    x"57",x"18",x"3E",x"06",x"32",x"0C",x"40",x"FD", -- 0x1568
    x"21",x"7A",x"40",x"FD",x"7E",x"04",x"FE",x"18", -- 0x1570
    x"D8",x"FE",x"2F",x"D0",x"C3",x"26",x"17",x"FD", -- 0x1578
    x"21",x"56",x"40",x"21",x"00",x"00",x"06",x"07", -- 0x1580
    x"FD",x"7E",x"04",x"E6",x"3F",x"FE",x"1C",x"28", -- 0x1588
    x"25",x"FE",x"20",x"28",x"21",x"FE",x"2C",x"28", -- 0x1590
    x"1D",x"FE",x"18",x"28",x"1D",x"FE",x"28",x"28", -- 0x1598
    x"19",x"11",x"06",x"00",x"FD",x"19",x"10",x"E0", -- 0x15A0
    x"7C",x"B7",x"C8",x"7D",x"B7",x"C0",x"21",x"56", -- 0x15A8
    x"40",x"06",x"2C",x"AF",x"D7",x"C9",x"26",x"01", -- 0x15B0
    x"18",x"E7",x"2E",x"01",x"18",x"E3",x"36",x"2E", -- 0x15B8
    x"D9",x"DD",x"66",x"00",x"DD",x"6E",x"01",x"0E", -- 0x15C0
    x"0E",x"CD",x"5B",x"00",x"DD",x"7E",x"04",x"E6", -- 0x15C8
    x"3F",x"32",x"24",x"40",x"DD",x"7E",x"FE",x"E6", -- 0x15D0
    x"3F",x"32",x"25",x"40",x"DD",x"7E",x"0A",x"E6", -- 0x15D8
    x"3F",x"32",x"26",x"40",x"21",x"24",x"40",x"7E", -- 0x15E0
    x"FE",x"20",x"28",x"1C",x"FE",x"2C",x"28",x"0E", -- 0x15E8
    x"FE",x"24",x"28",x"14",x"23",x"36",x"FF",x"23", -- 0x15F0
    x"CD",x"10",x"16",x"77",x"18",x"2A",x"23",x"CD", -- 0x15F8
    x"10",x"16",x"77",x"23",x"36",x"FF",x"18",x"20", -- 0x1600
    x"23",x"36",x"FF",x"23",x"36",x"FF",x"18",x"18", -- 0x1608
    x"7E",x"06",x"06",x"FD",x"21",x"22",x"16",x"FD", -- 0x1610
    x"BE",x"00",x"C8",x"FD",x"23",x"10",x"F8",x"3E", -- 0x1618
    x"FF",x"C9",x"18",x"1C",x"20",x"24",x"28",x"2C", -- 0x1620
    x"DD",x"E5",x"FD",x"E5",x"DD",x"21",x"61",x"17", -- 0x1628
    x"FD",x"21",x"8B",x"17",x"06",x"00",x"3A",x"24", -- 0x1630
    x"40",x"DD",x"BE",x"00",x"C2",x"3F",x"17",x"3A", -- 0x1638
    x"25",x"40",x"DD",x"BE",x"01",x"C2",x"3F",x"17", -- 0x1640
    x"3A",x"26",x"40",x"DD",x"BE",x"02",x"C2",x"3F", -- 0x1648
    x"17",x"FD",x"7E",x"00",x"32",x"21",x"40",x"FD", -- 0x1650
    x"7E",x"01",x"32",x"22",x"40",x"FD",x"7E",x"02", -- 0x1658
    x"32",x"23",x"40",x"FD",x"E1",x"DD",x"E1",x"DD", -- 0x1660
    x"7E",x"04",x"E6",x"80",x"5F",x"3A",x"21",x"40", -- 0x1668
    x"B7",x"CA",x"FE",x"16",x"FE",x"FF",x"28",x"34", -- 0x1670
    x"B3",x"DD",x"77",x"04",x"DD",x"7E",x"05",x"E6", -- 0x1678
    x"80",x"5F",x"3A",x"21",x"40",x"B3",x"DD",x"77", -- 0x1680
    x"05",x"CD",x"8E",x"16",x"18",x"1E",x"DD",x"7E", -- 0x1688
    x"04",x"E6",x"3F",x"FE",x"18",x"28",x"09",x"FE", -- 0x1690
    x"24",x"28",x"05",x"FE",x"28",x"28",x"01",x"C9", -- 0x1698
    x"DD",x"E5",x"DD",x"E5",x"FD",x"E1",x"CD",x"31", -- 0x16A0
    x"11",x"DD",x"E1",x"C9",x"3A",x"22",x"40",x"B7", -- 0x16A8
    x"28",x"55",x"57",x"FE",x"FF",x"28",x"16",x"DD", -- 0x16B0
    x"7E",x"FE",x"E6",x"80",x"5F",x"7A",x"B3",x"DD", -- 0x16B8
    x"77",x"FE",x"DD",x"7E",x"FF",x"E6",x"80",x"5F", -- 0x16C0
    x"7A",x"B3",x"DD",x"77",x"FF",x"3A",x"23",x"40", -- 0x16C8
    x"B7",x"28",x"42",x"FE",x"FF",x"28",x"25",x"57", -- 0x16D0
    x"DD",x"7E",x"0A",x"E6",x"80",x"5F",x"7A",x"B3", -- 0x16D8
    x"DD",x"77",x"0A",x"DD",x"7E",x"0B",x"E6",x"80", -- 0x16E0
    x"5F",x"7A",x"B3",x"DD",x"77",x"0B",x"DD",x"E5", -- 0x16E8
    x"D5",x"11",x"06",x"00",x"DD",x"19",x"CD",x"8E", -- 0x16F0
    x"16",x"D1",x"DD",x"E1",x"D9",x"C9",x"DD",x"E5", -- 0x16F8
    x"FD",x"E1",x"CD",x"26",x"17",x"18",x"A5",x"DD", -- 0x1700
    x"E5",x"FD",x"E1",x"11",x"FA",x"FF",x"FD",x"19", -- 0x1708
    x"CD",x"26",x"17",x"18",x"B8",x"DD",x"E5",x"FD", -- 0x1710
    x"E1",x"11",x"06",x"00",x"FD",x"19",x"CD",x"26", -- 0x1718
    x"17",x"C3",x"FC",x"16",x"FD",x"E1",x"FD",x"36", -- 0x1720
    x"00",x"00",x"FD",x"36",x"01",x"00",x"FD",x"36", -- 0x1728
    x"02",x"00",x"FD",x"36",x"03",x"00",x"FD",x"36", -- 0x1730
    x"04",x"00",x"FD",x"36",x"05",x"00",x"C9",x"04", -- 0x1738
    x"78",x"FE",x"10",x"20",x"0D",x"AF",x"21",x"56", -- 0x1740
    x"40",x"06",x"2C",x"D7",x"FD",x"E1",x"DD",x"E1", -- 0x1748
    x"D9",x"C9",x"DD",x"23",x"DD",x"23",x"DD",x"23", -- 0x1750
    x"FD",x"23",x"FD",x"23",x"FD",x"23",x"C3",x"36", -- 0x1758
    x"16",x"18",x"FF",x"1C",x"18",x"FF",x"20",x"18", -- 0x1760
    x"FF",x"2C",x"1C",x"FF",x"1C",x"1C",x"FF",x"20", -- 0x1768
    x"1C",x"FF",x"2C",x"20",x"FF",x"FF",x"24",x"FF", -- 0x1770
    x"FF",x"28",x"FF",x"1C",x"28",x"FF",x"20",x"28", -- 0x1778
    x"FF",x"2C",x"2C",x"18",x"FF",x"2C",x"1C",x"FF", -- 0x1780
    x"2C",x"28",x"FF",x"28",x"FF",x"FF",x"28",x"FF", -- 0x1788
    x"FF",x"24",x"FF",x"00",x"20",x"FF",x"18",x"20", -- 0x1790
    x"FF",x"24",x"20",x"FF",x"24",x"2C",x"FF",x"FF", -- 0x1798
    x"00",x"FF",x"FF",x"00",x"FF",x"18",x"00",x"FF", -- 0x17A0
    x"24",x"00",x"FF",x"00",x"00",x"24",x"FF",x"00", -- 0x17A8
    x"20",x"FF",x"00",x"00",x"FF",x"3A",x"10",x"40", -- 0x17B0
    x"E6",x"E3",x"32",x"10",x"40",x"31",x"00",x"44", -- 0x17B8
    x"3A",x"14",x"40",x"4F",x"3E",x"01",x"32",x"01", -- 0x17C0
    x"70",x"CB",x"51",x"20",x"03",x"32",x"03",x"68", -- 0x17C8
    x"3A",x"03",x"40",x"FE",x"E8",x"20",x"F9",x"3E", -- 0x17D0
    x"3D",x"32",x"55",x"40",x"3A",x"03",x"40",x"FE", -- 0x17D8
    x"F0",x"20",x"F9",x"3E",x"0E",x"32",x"55",x"40", -- 0x17E0
    x"AF",x"32",x"03",x"68",x"3A",x"0A",x"40",x"FE", -- 0x17E8
    x"28",x"30",x"08",x"3A",x"10",x"40",x"CB",x"CF", -- 0x17F0
    x"32",x"10",x"40",x"3E",x"80",x"32",x"02",x"40", -- 0x17F8
    x"3A",x"02",x"40",x"B7",x"20",x"FA",x"CD",x"82", -- 0x1800
    x"18",x"AF",x"32",x"04",x"70",x"3E",x"C0",x"CD", -- 0x1808
    x"4C",x"00",x"21",x"50",x"40",x"AF",x"06",x"2F", -- 0x1810
    x"D7",x"CD",x"E6",x"00",x"CD",x"49",x"00",x"CD", -- 0x1818
    x"EC",x"00",x"3E",x"C0",x"CD",x"4C",x"00",x"CD", -- 0x1820
    x"E9",x"00",x"3E",x"C0",x"CD",x"4C",x"00",x"3A", -- 0x1828
    x"0A",x"40",x"FE",x"28",x"30",x"08",x"3A",x"14", -- 0x1830
    x"40",x"CB",x"C7",x"32",x"14",x"40",x"CD",x"61", -- 0x1838
    x"00",x"CD",x"57",x"18",x"3E",x"C0",x"CD",x"4C", -- 0x1840
    x"00",x"3E",x"01",x"32",x"04",x"70",x"3A",x"14", -- 0x1848
    x"40",x"32",x"10",x"40",x"C3",x"10",x"15",x"3A", -- 0x1850
    x"14",x"40",x"CB",x"5F",x"28",x"06",x"DD",x"21", -- 0x1858
    x"00",x"41",x"18",x"04",x"DD",x"21",x"00",x"42", -- 0x1860
    x"21",x"46",x"43",x"DD",x"7E",x"0C",x"3C",x"E6", -- 0x1868
    x"07",x"DD",x"77",x"0C",x"7D",x"FE",x"60",x"D0", -- 0x1870
    x"DD",x"7E",x"0C",x"77",x"23",x"23",x"23",x"23", -- 0x1878
    x"18",x"F2",x"21",x"C0",x"53",x"7C",x"FE",x"4F", -- 0x1880
    x"C8",x"7E",x"E6",x"3C",x"FE",x"2C",x"E5",x"CC", -- 0x1888
    x"96",x"18",x"E1",x"2B",x"18",x"EF",x"56",x"E5", -- 0x1890
    x"DD",x"E5",x"CD",x"F6",x"00",x"CD",x"E0",x"00", -- 0x1898
    x"DD",x"E1",x"E1",x"36",x"FA",x"3A",x"14",x"40", -- 0x18A0
    x"CB",x"57",x"20",x"05",x"3E",x"01",x"32",x"03", -- 0x18A8
    x"68",x"3E",x"FC",x"CD",x"4C",x"00",x"36",x"FB", -- 0x18B0
    x"AF",x"32",x"03",x"68",x"3E",x"FC",x"CD",x"4C", -- 0x18B8
    x"00",x"36",x"10",x"C9",x"10",x"C9",x"FE",x"E8", -- 0x18C0
    x"38",x"13",x"3A",x"0C",x"40",x"B7",x"20",x"0B", -- 0x18C8
    x"CD",x"F6",x"16",x"3E",x"FF",x"32",x"00",x"78", -- 0x18D0
    x"C3",x"3E",x"10",x"CB",x"D1",x"3A",x"00",x"40", -- 0x18D8
    x"CB",x"77",x"20",x"0E",x"CB",x"61",x"FD",x"7E", -- 0x18E0
    x"00",x"20",x"03",x"93",x"18",x"01",x"83",x"FD", -- 0x18E8
    x"77",x"00",x"CB",x"51",x"FD",x"7E",x"01",x"28", -- 0x18F0
    x"03",x"93",x"18",x"01",x"83",x"FD",x"77",x"01", -- 0x18F8
    x"CB",x"51",x"FD",x"7E",x"05",x"28",x"0B",x"CB", -- 0x1900
    x"B7",x"FD",x"77",x"05",x"FD",x"71",x"04",x"C3", -- 0x1908
    x"3E",x"10",x"CB",x"F7",x"18",x"F3",x"3A",x"A2", -- 0x1910
    x"40",x"3C",x"32",x"A2",x"40",x"FD",x"7E",x"05", -- 0x1918
    x"E6",x"3F",x"FE",x"15",x"28",x"64",x"FD",x"7E", -- 0x1920
    x"04",x"E6",x"03",x"B7",x"20",x"02",x"3E",x"03", -- 0x1928
    x"4F",x"FD",x"7E",x"01",x"5F",x"FD",x"BE",x"0F", -- 0x1930
    x"38",x"38",x"3A",x"05",x"40",x"E6",x"0F",x"FE", -- 0x1938
    x"03",x"20",x"2F",x"FD",x"66",x"03",x"FD",x"6E", -- 0x1940
    x"02",x"11",x"20",x"00",x"19",x"7D",x"E6",x"1F", -- 0x1948
    x"FE",x"1C",x"30",x"0C",x"36",x"32",x"3E",x"FC", -- 0x1950
    x"32",x"00",x"40",x"3E",x"15",x"FD",x"77",x"05", -- 0x1958
    x"3A",x"10",x"40",x"CB",x"57",x"CA",x"3E",x"10", -- 0x1960
    x"FD",x"7E",x"01",x"2F",x"32",x"00",x"78",x"C3", -- 0x1968
    x"3E",x"10",x"F5",x"3A",x"10",x"40",x"CB",x"57", -- 0x1970
    x"F1",x"28",x"04",x"2F",x"32",x"00",x"78",x"7B", -- 0x1978
    x"81",x"FE",x"F0",x"30",x"12",x"FD",x"77",x"01", -- 0x1980
    x"18",x"E5",x"3A",x"00",x"40",x"B7",x"20",x"DF", -- 0x1988
    x"3E",x"14",x"FD",x"77",x"05",x"18",x"D8",x"CD", -- 0x1990
    x"F6",x"16",x"3E",x"FF",x"32",x"00",x"78",x"18", -- 0x1998
    x"CE",x"3A",x"A1",x"40",x"3C",x"32",x"A1",x"40", -- 0x19A0
    x"3A",x"00",x"40",x"5F",x"FD",x"7E",x"04",x"4F", -- 0x19A8
    x"E6",x"03",x"B7",x"20",x"02",x"3E",x"03",x"57", -- 0x19B0
    x"FD",x"7E",x"00",x"CB",x"61",x"20",x"03",x"82", -- 0x19B8
    x"18",x"01",x"92",x"FD",x"77",x"00",x"FE",x"08", -- 0x19C0
    x"38",x"CD",x"FE",x"F8",x"30",x"C9",x"CB",x"53", -- 0x19C8
    x"20",x"04",x"3E",x"12",x"18",x"02",x"3E",x"13", -- 0x19D0
    x"CB",x"61",x"28",x"02",x"CB",x"FF",x"FD",x"77", -- 0x19D8
    x"05",x"FD",x"66",x"03",x"FD",x"6E",x"02",x"23", -- 0x19E0
    x"11",x"20",x"00",x"19",x"7E",x"FE",x"10",x"28", -- 0x19E8
    x"02",x"36",x"FA",x"C3",x"3E",x"10",x"00",x"00", -- 0x19F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19F8
    x"FD",x"E5",x"DD",x"E5",x"CD",x"0C",x"1A",x"DD", -- 0x1A00
    x"E1",x"FD",x"E1",x"C9",x"FD",x"21",x"00",x"40", -- 0x1A08
    x"FD",x"7E",x"0C",x"B7",x"C8",x"FD",x"7E",x"00", -- 0x1A10
    x"4F",x"3A",x"10",x"40",x"FE",x"04",x"28",x"6C", -- 0x1A18
    x"FD",x"7E",x"10",x"CB",x"5F",x"28",x"06",x"DD", -- 0x1A20
    x"21",x"00",x"41",x"18",x"04",x"DD",x"21",x"00", -- 0x1A28
    x"42",x"DD",x"7E",x"04",x"FE",x"04",x"D8",x"DD", -- 0x1A30
    x"7E",x"0A",x"FE",x"10",x"38",x"05",x"3E",x"0E", -- 0x1A38
    x"DD",x"77",x"0A",x"47",x"DD",x"7E",x"01",x"5F", -- 0x1A40
    x"E6",x"0F",x"57",x"78",x"FE",x"0F",x"20",x"0C", -- 0x1A48
    x"CB",x"79",x"20",x"08",x"FD",x"34",x"01",x"CB", -- 0x1A50
    x"B9",x"FD",x"71",x"00",x"7A",x"B7",x"CA",x"52", -- 0x1A58
    x"1B",x"FE",x"02",x"28",x"17",x"FE",x"04",x"28", -- 0x1A60
    x"53",x"FE",x"08",x"28",x"0F",x"FE",x"A0",x"CA", -- 0x1A68
    x"7F",x"1B",x"FE",x"C0",x"CA",x"03",x"1B",x"FE", -- 0x1A70
    x"E0",x"28",x"41",x"C9",x"FD",x"34",x"01",x"CB", -- 0x1A78
    x"61",x"C8",x"3A",x"10",x"40",x"CB",x"57",x"20", -- 0x1A80
    x"0F",x"DD",x"7E",x"0A",x"21",x"00",x"21",x"CD", -- 0x1A88
    x"B6",x"1B",x"3A",x"A0",x"40",x"BA",x"C8",x"D0", -- 0x1A90
    x"3E",x"F0",x"C5",x"D5",x"67",x"2E",x"F0",x"0E", -- 0x1A98
    x"10",x"CD",x"5B",x"00",x"D1",x"C1",x"B7",x"C8", -- 0x1AA0
    x"7B",x"FE",x"01",x"28",x"05",x"CB",x"51",x"20", -- 0x1AA8
    x"01",x"1D",x"7B",x"C6",x"04",x"FD",x"77",x"04", -- 0x1AB0
    x"DD",x"34",x"04",x"C9",x"FD",x"34",x"01",x"CB", -- 0x1AB8
    x"41",x"C8",x"3A",x"05",x"40",x"FE",x"20",x"38", -- 0x1AC0
    x"04",x"FE",x"D0",x"38",x"02",x"C6",x"80",x"F5", -- 0x1AC8
    x"DD",x"7E",x"0A",x"21",x"1F",x"21",x"CD",x"B6", -- 0x1AD0
    x"1B",x"3A",x"A2",x"40",x"BA",x"28",x"22",x"30", -- 0x1AD8
    x"20",x"F1",x"C5",x"D5",x"67",x"2E",x"08",x"0E", -- 0x1AE0
    x"14",x"CD",x"5B",x"00",x"D1",x"E1",x"B7",x"C8", -- 0x1AE8
    x"7B",x"FE",x"01",x"28",x"05",x"CB",x"49",x"20", -- 0x1AF0
    x"01",x"1D",x"FD",x"73",x"04",x"DD",x"34",x"04", -- 0x1AF8
    x"C9",x"F1",x"C9",x"FD",x"34",x"01",x"CB",x"41", -- 0x1B00
    x"C8",x"FD",x"34",x"01",x"DD",x"7E",x"0A",x"21", -- 0x1B08
    x"3D",x"21",x"CD",x"B6",x"1B",x"3A",x"A1",x"40", -- 0x1B10
    x"BA",x"D0",x"3A",x"05",x"40",x"FE",x"20",x"38", -- 0x1B18
    x"04",x"FE",x"E0",x"38",x"02",x"C6",x"80",x"6F", -- 0x1B20
    x"C5",x"D5",x"CB",x"49",x"28",x"04",x"26",x"10", -- 0x1B28
    x"18",x"02",x"26",x"F0",x"0E",x"12",x"CD",x"5B", -- 0x1B30
    x"00",x"B7",x"D1",x"C1",x"C8",x"CB",x"49",x"20", -- 0x1B38
    x"07",x"FD",x"73",x"04",x"FD",x"34",x"04",x"C9", -- 0x1B40
    x"7B",x"C6",x"10",x"FD",x"73",x"04",x"FD",x"34", -- 0x1B48
    x"04",x"C9",x"FD",x"34",x"01",x"3A",x"A1",x"40", -- 0x1B50
    x"B7",x"C0",x"3A",x"51",x"40",x"FE",x"C0",x"D0", -- 0x1B58
    x"6F",x"3A",x"50",x"40",x"FE",x"80",x"30",x"06", -- 0x1B60
    x"26",x"10",x"0E",x"02",x"18",x"04",x"26",x"F0", -- 0x1B68
    x"0E",x"12",x"C5",x"0E",x"12",x"CD",x"5B",x"00", -- 0x1B70
    x"C1",x"B7",x"C8",x"FD",x"71",x"04",x"C9",x"FD", -- 0x1B78
    x"34",x"01",x"3A",x"0C",x"40",x"FE",x"02",x"D8", -- 0x1B80
    x"DD",x"7E",x"0A",x"FE",x"06",x"D8",x"3A",x"01", -- 0x1B88
    x"40",x"3C",x"32",x"01",x"40",x"3A",x"05",x"40", -- 0x1B90
    x"E6",x"7F",x"67",x"2E",x"08",x"0E",x"24",x"CD", -- 0x1B98
    x"5B",x"00",x"FD",x"36",x"04",x"24",x"DD",x"7E", -- 0x1BA0
    x"04",x"67",x"2E",x"08",x"0E",x"24",x"CD",x"5B", -- 0x1BA8
    x"00",x"FD",x"36",x"04",x"24",x"C9",x"47",x"7E", -- 0x1BB0
    x"B8",x"30",x"02",x"18",x"05",x"23",x"5E",x"23", -- 0x1BB8
    x"56",x"C9",x"23",x"23",x"23",x"18",x"F0",x"56", -- 0x1BC0
    x"C9",x"23",x"23",x"23",x"18",x"F0",x"C9",x"23", -- 0x1BC8
    x"23",x"23",x"18",x"F0",x"23",x"18",x"F0",x"18", -- 0x1BD0
    x"04",x"DD",x"21",x"00",x"41",x"DD",x"7E",x"0D", -- 0x1BD8
    x"B7",x"C0",x"3A",x"00",x"70",x"CB",x"5F",x"28", -- 0x1BE0
    x"05",x"3A",x"4E",x"1C",x"18",x"03",x"3A",x"4F", -- 0x1BE8
    x"1C",x"DD",x"BE",x"00",x"C0",x"DD",x"36",x"0D", -- 0x1BF0
    x"01",x"DD",x"36",x"0E",x"01",x"DD",x"34",x"09", -- 0x1BF8
    x"11",x"38",x"1C",x"E7",x"11",x"2A",x"1C",x"E7", -- 0x1C00
    x"3A",x"10",x"40",x"F5",x"AF",x"32",x"10",x"40", -- 0x1C08
    x"21",x"00",x"1D",x"22",x"C0",x"40",x"AF",x"32", -- 0x1C10
    x"00",x"40",x"3A",x"00",x"40",x"FE",x"80",x"20", -- 0x1C18
    x"F9",x"11",x"38",x"1C",x"E7",x"F1",x"32",x"10", -- 0x1C20
    x"40",x"C9",x"01",x"1F",x"04",x"42",x"4F",x"4E", -- 0x1C28
    x"55",x"53",x"40",x"42",x"41",x"53",x"45",x"FF", -- 0x1C30
    x"05",x"1F",x"00",x"40",x"40",x"40",x"40",x"40", -- 0x1C38
    x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40", -- 0x1C40
    x"40",x"40",x"40",x"40",x"40",x"FF",x"50",x"75", -- 0x1C48
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C50
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C58
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C60
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C68
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C78
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C80
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C88
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C90
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CA8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CB0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CC0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CC8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CD0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CD8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CF8
    x"00",x"20",x"20",x"30",x"30",x"40",x"40",x"50", -- 0x1D00
    x"50",x"80",x"80",x"70",x"70",x"50",x"50",x"FF", -- 0x1D08
    x"44",x"77",x"99",x"AA",x"D0",x"80",x"60",x"40", -- 0x1D10
    x"50",x"80",x"80",x"80",x"FF",x"00",x"00",x"00", -- 0x1D18
    x"AA",x"BB",x"CC",x"DD",x"AA",x"90",x"80",x"FF", -- 0x1D20
    x"40",x"FF",x"C0",x"B0",x"A0",x"90",x"80",x"FF", -- 0x1D28
    x"12",x"34",x"56",x"78",x"9A",x"BC",x"DE",x"F1", -- 0x1D30
    x"23",x"45",x"67",x"FF",x"AB",x"CD",x"FF",x"00", -- 0x1D38
    x"F0",x"DC",x"BA",x"98",x"76",x"54",x"32",x"12", -- 0x1D40
    x"34",x"FF",x"78",x"9A",x"FF",x"00",x"00",x"00", -- 0x1D48
    x"C3",x"10",x"43",x"3E",x"1A",x"01",x"22",x"45", -- 0x1D50
    x"C9",x"01",x"FF",x"10",x"22",x"83",x"FF",x"00", -- 0x1D58
    x"10",x"10",x"20",x"20",x"30",x"30",x"40",x"40", -- 0x1D60
    x"30",x"30",x"20",x"20",x"10",x"10",x"FF",x"00", -- 0x1D68
    x"50",x"60",x"70",x"80",x"90",x"A0",x"B0",x"A0", -- 0x1D70
    x"90",x"80",x"70",x"FF",x"50",x"FF",x"00",x"00", -- 0x1D78
    x"F0",x"E0",x"C0",x"D0",x"E0",x"F0",x"D0",x"C0", -- 0x1D80
    x"A0",x"D0",x"FF",x"E0",x"F0",x"FF",x"00",x"00", -- 0x1D88
    x"18",x"68",x"74",x"98",x"A0",x"98",x"74",x"68", -- 0x1D90
    x"36",x"38",x"FF",x"3C",x"3E",x"FF",x"00",x"00", -- 0x1D98
    x"10",x"80",x"20",x"A0",x"30",x"E0",x"40",x"80", -- 0x1DA0
    x"80",x"FF",x"70",x"68",x"60",x"20",x"20",x"FF", -- 0x1DA8
    x"22",x"33",x"45",x"67",x"65",x"55",x"F0",x"E0", -- 0x1DB0
    x"20",x"30",x"20",x"30",x"20",x"FF",x"00",x"00", -- 0x1DB8
    x"82",x"84",x"86",x"88",x"8A",x"8C",x"8E",x"90", -- 0x1DC0
    x"92",x"94",x"96",x"98",x"9A",x"9C",x"9E",x"FF", -- 0x1DC8
    x"F0",x"E8",x"E0",x"D8",x"D0",x"C8",x"C0",x"B8", -- 0x1DD0
    x"B0",x"A8",x"A0",x"E0",x"F0",x"F0",x"F0",x"FF", -- 0x1DD8
    x"30",x"50",x"70",x"80",x"70",x"60",x"50",x"40", -- 0x1DE0
    x"30",x"20",x"10",x"FF",x"00",x"00",x"00",x"00", -- 0x1DE8
    x"80",x"80",x"F0",x"D9",x"68",x"65",x"D6",x"D7", -- 0x1DF0
    x"D9",x"22",x"33",x"44",x"55",x"66",x"77",x"FF", -- 0x1DF8
    x"AF",x"32",x"10",x"40",x"3E",x"C0",x"CD",x"4C", -- 0x1E00
    x"00",x"21",x"00",x"70",x"AF",x"06",x"20",x"D7", -- 0x1E08
    x"3E",x"01",x"32",x"01",x"70",x"21",x"00",x"43", -- 0x1E10
    x"06",x"40",x"D7",x"3A",x"00",x"68",x"E6",x"C0", -- 0x1E18
    x"FE",x"C0",x"20",x"05",x"3E",x"02",x"32",x"06", -- 0x1E20
    x"40",x"11",x"7D",x"1F",x"E7",x"3E",x"C0",x"CD", -- 0x1E28
    x"4C",x"00",x"11",x"92",x"1F",x"E7",x"3E",x"C0", -- 0x1E30
    x"CD",x"4C",x"00",x"11",x"9E",x"1F",x"E7",x"3E", -- 0x1E38
    x"80",x"CD",x"4C",x"00",x"11",x"C2",x"1F",x"E7", -- 0x1E40
    x"3E",x"80",x"CD",x"4C",x"00",x"11",x"C8",x"1F", -- 0x1E48
    x"E7",x"11",x"B1",x"1F",x"E7",x"3E",x"80",x"CD", -- 0x1E50
    x"4C",x"00",x"11",x"E5",x"1F",x"E7",x"3E",x"2B", -- 0x1E58
    x"32",x"98",x"53",x"3E",x"80",x"CD",x"4C",x"00", -- 0x1E60
    x"11",x"F9",x"1F",x"E7",x"11",x"19",x"20",x"E7", -- 0x1E68
    x"11",x"35",x"20",x"E7",x"3E",x"C0",x"CD",x"4C", -- 0x1E70
    x"00",x"CD",x"49",x"00",x"3E",x"C0",x"CD",x"4C", -- 0x1E78
    x"00",x"11",x"43",x"20",x"E7",x"3E",x"C0",x"CD", -- 0x1E80
    x"4C",x"00",x"DD",x"21",x"5A",x"20",x"FD",x"21", -- 0x1E88
    x"50",x"40",x"06",x"04",x"DD",x"7E",x"00",x"FD", -- 0x1E90
    x"77",x"00",x"DD",x"7E",x"01",x"FD",x"77",x"01", -- 0x1E98
    x"DD",x"7E",x"02",x"FD",x"77",x"05",x"11",x"06", -- 0x1EA0
    x"00",x"FD",x"19",x"11",x"03",x"00",x"DD",x"19", -- 0x1EA8
    x"10",x"E2",x"FD",x"E5",x"11",x"66",x"20",x"E7", -- 0x1EB0
    x"FD",x"E1",x"FD",x"36",x"00",x"40",x"FD",x"36", -- 0x1EB8
    x"01",x"E0",x"FD",x"36",x"05",x"10",x"FD",x"E5", -- 0x1EC0
    x"11",x"72",x"20",x"E7",x"FD",x"E1",x"FD",x"36", -- 0x1EC8
    x"06",x"40",x"FD",x"36",x"07",x"C0",x"FD",x"36", -- 0x1ED0
    x"0B",x"12",x"FD",x"E5",x"11",x"79",x"20",x"E7", -- 0x1ED8
    x"FD",x"E1",x"FD",x"36",x"0C",x"40",x"FD",x"36", -- 0x1EE0
    x"0D",x"A0",x"FD",x"36",x"11",x"14",x"11",x"80", -- 0x1EE8
    x"20",x"E7",x"3E",x"32",x"32",x"E7",x"52",x"11", -- 0x1EF0
    x"87",x"20",x"E7",x"3E",x"F8",x"32",x"EB",x"52", -- 0x1EF8
    x"11",x"8F",x"20",x"E7",x"3E",x"10",x"CD",x"4C", -- 0x1F00
    x"00",x"CD",x"49",x"00",x"3E",x"C0",x"CD",x"4C", -- 0x1F08
    x"00",x"11",x"9A",x"20",x"E7",x"3E",x"C0",x"CD", -- 0x1F10
    x"4C",x"00",x"11",x"B0",x"20",x"E7",x"3E",x"C0", -- 0x1F18
    x"CD",x"4C",x"00",x"3A",x"0F",x"00",x"B7",x"CA", -- 0x1F20
    x"1C",x"25",x"3A",x"00",x"68",x"07",x"07",x"B7", -- 0x1F28
    x"28",x"06",x"11",x"D0",x"20",x"E7",x"18",x"04", -- 0x1F30
    x"11",x"C0",x"20",x"E7",x"3E",x"80",x"CD",x"4C", -- 0x1F38
    x"00",x"CD",x"49",x"00",x"3E",x"C0",x"CD",x"4C", -- 0x1F40
    x"00",x"CD",x"4F",x"00",x"3A",x"10",x"40",x"CB", -- 0x1F48
    x"C7",x"32",x"10",x"40",x"3A",x"10",x"40",x"CB", -- 0x1F50
    x"47",x"20",x"F9",x"3E",x"01",x"32",x"04",x"70", -- 0x1F58
    x"3E",x"04",x"32",x"10",x"40",x"32",x"14",x"40", -- 0x1F60
    x"3E",x"01",x"32",x"09",x"41",x"32",x"09",x"42", -- 0x1F68
    x"3E",x"08",x"32",x"0A",x"42",x"32",x"0A",x"41", -- 0x1F70
    x"CD",x"E0",x"00",x"18",x"FE",x"02",x"04",x"05", -- 0x1F78
    x"46",x"4F",x"4F",x"44",x"40",x"41",x"4E",x"44", -- 0x1F80
    x"40",x"46",x"55",x"4E",x"40",x"43",x"4F",x"52", -- 0x1F88
    x"50",x"FF",x"03",x"08",x"0A",x"50",x"52",x"45", -- 0x1F90
    x"53",x"45",x"4E",x"54",x"53",x"FF",x"04",x"0C", -- 0x1F98
    x"06",x"57",x"41",x"52",x"40",x"4F",x"46",x"40", -- 0x1FA0
    x"54",x"48",x"45",x"40",x"42",x"55",x"47",x"53", -- 0x1FA8
    x"FF",x"06",x"13",x"08",x"4D",x"55",x"53",x"48", -- 0x1FB0
    x"52",x"4F",x"4F",x"4D",x"40",x"4D",x"41",x"5A", -- 0x1FB8
    x"45",x"FF",x"05",x"0E",x"0C",x"4F",x"52",x"FF", -- 0x1FC0
    x"06",x"11",x"02",x"4D",x"4F",x"4E",x"53",x"54", -- 0x1FC8
    x"45",x"52",x"4F",x"55",x"53",x"40",x"4D",x"41", -- 0x1FD0
    x"4E",x"4F",x"55",x"56",x"45",x"52",x"53",x"40", -- 0x1FD8
    x"49",x"4E",x"40",x"41",x"FF",x"00",x"18",x"06", -- 0x1FE0
    x"41",x"52",x"4D",x"45",x"4E",x"49",x"41",x"40", -- 0x1FE8
    x"4C",x"54",x"44",x"40",x"31",x"39",x"38",x"31", -- 0x1FF0
    x"FF",x"07",x"1D",x"00",x"50",x"52",x"4F",x"47", -- 0x1FF8
    x"FF",x"41",x"4D",x"4D",x"49",x"4E",x"47",x"40", -- 0x2000
    x"54",x"4F",x"54",x"41",x"4C",x"4C",x"59",x"40", -- 0x2008
    x"4F",x"52",x"49",x"47",x"49",x"4E",x"41",x"4C", -- 0x2010
    x"FF",x"07",x"1E",x"02",x"55",x"4E",x"41",x"55", -- 0x2018
    x"54",x"48",x"4F",x"52",x"49",x"53",x"45",x"44", -- 0x2020
    x"40",x"44",x"55",x"50",x"4C",x"49",x"43",x"41", -- 0x2028
    x"54",x"49",x"4F",x"4E",x"FF",x"07",x"1F",x"09", -- 0x2030
    x"50",x"52",x"4F",x"48",x"49",x"42",x"49",x"54", -- 0x2038
    x"45",x"44",x"FF",x"07",x"03",x"04",x"53",x"43", -- 0x2040
    x"4F",x"52",x"45",x"40",x"41",x"44",x"56",x"41", -- 0x2048
    x"4E",x"43",x"45",x"40",x"54",x"41",x"42",x"4C", -- 0x2050
    x"45",x"FF",x"40",x"80",x"18",x"50",x"80",x"1C", -- 0x2058
    x"60",x"80",x"1C",x"70",x"80",x"20",x"00",x"07", -- 0x2060
    x"10",x"32",x"30",x"40",x"33",x"30",x"40",x"34", -- 0x2068
    x"30",x"FF",x"01",x"0B",x"15",x"39",x"30",x"30", -- 0x2070
    x"FF",x"00",x"10",x"15",x"31",x"30",x"30",x"FF", -- 0x2078
    x"00",x"14",x"15",x"36",x"30",x"30",x"FF",x"00", -- 0x2080
    x"19",x"15",x"35",x"30",x"30",x"30",x"FF",x"00", -- 0x2088
    x"1D",x"13",x"4D",x"59",x"53",x"54",x"45",x"52", -- 0x2090
    x"59",x"FF",x"03",x"06",x"04",x"4F",x"4E",x"45", -- 0x2098
    x"40",x"4F",x"52",x"40",x"54",x"57",x"4F",x"40", -- 0x20A0
    x"50",x"4C",x"41",x"59",x"45",x"52",x"53",x"FF", -- 0x20A8
    x"04",x"0A",x"07",x"49",x"4E",x"53",x"45",x"52", -- 0x20B0
    x"54",x"40",x"43",x"4F",x"49",x"4E",x"53",x"FF", -- 0x20B8
    x"05",x"18",x"07",x"4F",x"4E",x"45",x"40",x"50", -- 0x20C0
    x"4C",x"41",x"59",x"40",x"32",x"30",x"43",x"FF", -- 0x20C8
    x"05",x"18",x"07",x"4F",x"4E",x"45",x"40",x"50", -- 0x20D0
    x"4C",x"41",x"59",x"40",x"32",x"30",x"43",x"FF", -- 0x20D8
    x"3E",x"02",x"32",x"06",x"40",x"18",x"FE",x"00", -- 0x20E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x20E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x20F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x20F8
    x"00",x"01",x"01",x"01",x"01",x"01",x"03",x"02", -- 0x2100
    x"01",x"06",x"03",x"01",x"08",x"03",x"01",x"0C", -- 0x2108
    x"03",x"02",x"00",x"00",x"00",x"00",x"10",x"03", -- 0x2110
    x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2118
    x"02",x"01",x"02",x"03",x"01",x"04",x"02",x"02", -- 0x2120
    x"08",x"03",x"03",x"0A",x"03",x"03",x"00",x"00", -- 0x2128
    x"00",x"00",x"00",x"00",x"10",x"03",x"04",x"00", -- 0x2130
    x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"01", -- 0x2138
    x"04",x"00",x"02",x"01",x"0F",x"03",x"03",x"06", -- 0x2140
    x"01",x"03",x"10",x"01",x"03",x"00",x"00",x"00", -- 0x2148
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2150
    x"00",x"3A",x"10",x"40",x"E6",x"18",x"B7",x"C8", -- 0x2158
    x"CB",x"5F",x"20",x"06",x"DD",x"21",x"00",x"42", -- 0x2160
    x"18",x"04",x"DD",x"21",x"00",x"41",x"DD",x"7E", -- 0x2168
    x"0D",x"B7",x"C0",x"3A",x"00",x"70",x"CB",x"5F", -- 0x2170
    x"28",x"05",x"3A",x"DF",x"21",x"18",x"03",x"3A", -- 0x2178
    x"E0",x"21",x"DD",x"BE",x"00",x"C0",x"DD",x"36", -- 0x2180
    x"0D",x"01",x"DD",x"36",x"0E",x"01",x"DD",x"34", -- 0x2188
    x"09",x"11",x"C9",x"21",x"E7",x"11",x"BB",x"21", -- 0x2190
    x"E7",x"3A",x"10",x"40",x"F5",x"AF",x"32",x"10", -- 0x2198
    x"40",x"21",x"00",x"1D",x"22",x"C0",x"40",x"AF", -- 0x21A0
    x"32",x"00",x"40",x"3A",x"00",x"40",x"FE",x"80", -- 0x21A8
    x"20",x"F9",x"11",x"C9",x"21",x"E7",x"F1",x"32", -- 0x21B0
    x"10",x"40",x"C9",x"01",x"1F",x"04",x"42",x"4F", -- 0x21B8
    x"4E",x"55",x"53",x"40",x"42",x"41",x"53",x"45", -- 0x21C0
    x"FF",x"05",x"1F",x"00",x"40",x"40",x"40",x"40", -- 0x21C8
    x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40", -- 0x21D0
    x"40",x"40",x"40",x"40",x"40",x"40",x"FF",x"50", -- 0x21D8
    x"75",x"CD",x"00",x"1A",x"2A",x"C0",x"40",x"7C", -- 0x21E0
    x"FE",x"18",x"30",x"07",x"3E",x"FF",x"32",x"00", -- 0x21E8
    x"78",x"18",x"29",x"3A",x"C2",x"40",x"3C",x"32", -- 0x21F0
    x"C2",x"40",x"2A",x"C0",x"40",x"7E",x"FE",x"01", -- 0x21F8
    x"C8",x"32",x"00",x"78",x"FE",x"FF",x"28",x"14", -- 0x2200
    x"3A",x"C2",x"40",x"CB",x"57",x"C8",x"CB",x"97", -- 0x2208
    x"32",x"C2",x"40",x"7E",x"32",x"00",x"78",x"23", -- 0x2210
    x"22",x"C0",x"40",x"C9",x"2A",x"D0",x"22",x"22", -- 0x2218
    x"C0",x"40",x"3A",x"10",x"40",x"E6",x"18",x"20", -- 0x2220
    x"08",x"21",x"00",x"68",x"AF",x"06",x"00",x"D7", -- 0x2228
    x"C9",x"3A",x"A0",x"40",x"B7",x"20",x"3C",x"CD", -- 0x2230
    x"4C",x"22",x"3A",x"0C",x"40",x"DD",x"21",x"D1", -- 0x2238
    x"22",x"DD",x"BE",x"00",x"28",x"1B",x"DD",x"23", -- 0x2240
    x"DD",x"23",x"18",x"F5",x"3A",x"A2",x"40",x"B7", -- 0x2248
    x"C8",x"3A",x"C8",x"40",x"2F",x"FE",x"20",x"28", -- 0x2250
    x"04",x"32",x"00",x"78",x"C9",x"3E",x"FF",x"18", -- 0x2258
    x"F8",x"DD",x"7E",x"00",x"DD",x"21",x"00",x"68", -- 0x2260
    x"06",x"07",x"DD",x"77",x"00",x"CB",x"3F",x"DD", -- 0x2268
    x"23",x"10",x"F7",x"3A",x"A1",x"40",x"B7",x"28", -- 0x2270
    x"0C",x"3A",x"00",x"40",x"07",x"07",x"07",x"07", -- 0x2278
    x"32",x"00",x"78",x"18",x"16",x"3A",x"A0",x"40", -- 0x2280
    x"B7",x"28",x"10",x"3A",x"00",x"40",x"CB",x"5F", -- 0x2288
    x"28",x"04",x"3E",x"20",x"18",x"02",x"3E",x"40", -- 0x2290
    x"32",x"00",x"78",x"3A",x"A9",x"40",x"B7",x"28", -- 0x2298
    x"1E",x"DD",x"21",x"DF",x"22",x"DD",x"BE",x"00", -- 0x22A0
    x"28",x"08",x"DD",x"23",x"DD",x"23",x"DD",x"23", -- 0x22A8
    x"18",x"F3",x"DD",x"66",x"02",x"DD",x"6E",x"01", -- 0x22B0
    x"22",x"C0",x"40",x"AF",x"32",x"A9",x"40",x"3A", -- 0x22B8
    x"A8",x"40",x"FE",x"50",x"C0",x"AF",x"32",x"A8", -- 0x22C0
    x"40",x"21",x"A0",x"1D",x"22",x"C0",x"40",x"C9", -- 0x22C8
    x"01",x"01",x"01",x"02",x"02",x"03",x"03",x"04", -- 0x22D0
    x"13",x"05",x"33",x"06",x"FF",x"00",x"00",x"01", -- 0x22D8
    x"20",x"1D",x"02",x"40",x"1D",x"03",x"40",x"1D", -- 0x22E0
    x"04",x"50",x"1D",x"05",x"60",x"1D",x"06",x"70", -- 0x22E8
    x"1D",x"07",x"80",x"1D",x"08",x"90",x"1D",x"09", -- 0x22F0
    x"A0",x"1D",x"09",x"B0",x"1D",x"50",x"C0",x"1D", -- 0x22F8
    x"0F",x"A0",x"40",x"3C",x"32",x"A0",x"40",x"FD", -- 0x2300
    x"7E",x"04",x"4F",x"E6",x"03",x"B7",x"20",x"02", -- 0x2308
    x"3E",x"01",x"00",x"00",x"5F",x"FD",x"7E",x"05", -- 0x2310
    x"E6",x"3E",x"57",x"3A",x"00",x"40",x"CB",x"3F", -- 0x2318
    x"CB",x"3F",x"E6",x"01",x"B2",x"FD",x"77",x"05", -- 0x2320
    x"FD",x"7E",x"00",x"FE",x"20",x"30",x"04",x"CB", -- 0x2328
    x"E1",x"18",x"06",x"FE",x"E8",x"38",x"02",x"CB", -- 0x2330
    x"A1",x"FD",x"7E",x"01",x"FE",x"80",x"30",x"04", -- 0x2338
    x"CB",x"91",x"18",x"17",x"FE",x"E8",x"38",x"13", -- 0x2340
    x"3A",x"0C",x"40",x"B7",x"20",x"0B",x"CD",x"0A", -- 0x2348
    x"17",x"3E",x"FF",x"32",x"00",x"78",x"C3",x"3E", -- 0x2350
    x"10",x"CB",x"D1",x"3A",x"00",x"40",x"CB",x"77", -- 0x2358
    x"20",x"0E",x"CB",x"61",x"FD",x"7E",x"00",x"20", -- 0x2360
    x"03",x"93",x"18",x"01",x"83",x"FD",x"77",x"00", -- 0x2368
    x"CB",x"51",x"FD",x"7E",x"01",x"28",x"03",x"93", -- 0x2370
    x"18",x"01",x"83",x"FD",x"77",x"01",x"CB",x"51", -- 0x2378
    x"FD",x"7E",x"05",x"28",x"0B",x"CB",x"B7",x"FD", -- 0x2380
    x"77",x"05",x"FD",x"71",x"04",x"C3",x"3E",x"10", -- 0x2388
    x"CB",x"F7",x"18",x"F3",x"3A",x"A2",x"40",x"3C", -- 0x2390
    x"32",x"A2",x"40",x"FD",x"7E",x"01",x"32",x"00", -- 0x2398
    x"78",x"FD",x"7E",x"05",x"E6",x"3F",x"FE",x"15", -- 0x23A0
    x"28",x"50",x"FD",x"7E",x"04",x"E6",x"03",x"B7", -- 0x23A8
    x"20",x"02",x"3E",x"03",x"4F",x"FD",x"7E",x"01", -- 0x23B0
    x"5F",x"3A",x"05",x"40",x"E6",x"1F",x"FE",x"05", -- 0x23B8
    x"20",x"28",x"FD",x"7E",x"01",x"FE",x"30",x"38", -- 0x23C0
    x"21",x"FD",x"66",x"03",x"FD",x"6E",x"02",x"11", -- 0x23C8
    x"20",x"00",x"19",x"7D",x"E6",x"1F",x"FE",x"1D", -- 0x23D0
    x"D2",x"3E",x"10",x"36",x"32",x"3E",x"FC",x"32", -- 0x23D8
    x"00",x"40",x"3E",x"15",x"FD",x"77",x"05",x"C3", -- 0x23E0
    x"3E",x"10",x"7B",x"81",x"FE",x"80",x"38",x"01", -- 0x23E8
    x"3C",x"FE",x"F8",x"30",x"12",x"FD",x"77",x"01", -- 0x23F0
    x"18",x"ED",x"3A",x"00",x"40",x"B7",x"20",x"E7", -- 0x23F8
    x"3E",x"14",x"FD",x"77",x"05",x"18",x"E0",x"CD", -- 0x2400
    x"0A",x"17",x"3E",x"FF",x"32",x"00",x"78",x"18", -- 0x2408
    x"D6",x"3A",x"A1",x"40",x"3C",x"32",x"A1",x"40", -- 0x2410
    x"3A",x"00",x"40",x"5F",x"FD",x"7E",x"04",x"4F", -- 0x2418
    x"E6",x"03",x"B7",x"20",x"02",x"3E",x"03",x"57", -- 0x2420
    x"FD",x"7E",x"00",x"CB",x"61",x"20",x"03",x"82", -- 0x2428
    x"18",x"01",x"92",x"FD",x"77",x"00",x"FE",x"08", -- 0x2430
    x"38",x"CD",x"FE",x"F8",x"30",x"C9",x"CB",x"53", -- 0x2438
    x"20",x"04",x"3E",x"12",x"18",x"02",x"3E",x"13", -- 0x2440
    x"CB",x"61",x"28",x"02",x"CB",x"FF",x"FD",x"77", -- 0x2448
    x"05",x"FD",x"66",x"03",x"FD",x"6E",x"02",x"23", -- 0x2450
    x"11",x"20",x"00",x"19",x"7E",x"FE",x"10",x"28", -- 0x2458
    x"02",x"36",x"FA",x"C3",x"3E",x"10",x"03",x"03", -- 0x2460
    x"00",x"56",x"40",x"20",x"02",x"02",x"00",x"0C", -- 0x2468
    x"40",x"04",x"6F",x"3A",x"14",x"40",x"CB",x"67", -- 0x2470
    x"C8",x"3E",x"01",x"32",x"06",x"70",x"32",x"07", -- 0x2478
    x"70",x"C9",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2480
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2488
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2490
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2498
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x24A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x24A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x24B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x24B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x24C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x24C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x24D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x24D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x24E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x24E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x24F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x24F8
    x"3A",x"00",x"60",x"CB",x"6F",x"C8",x"3A",x"14", -- 0x2500
    x"40",x"CB",x"67",x"20",x"0B",x"AF",x"32",x"0F", -- 0x2508
    x"40",x"32",x"06",x"70",x"32",x"07",x"70",x"C9", -- 0x2510
    x"3E",x"01",x"18",x"F2",x"3E",x"C0",x"CD",x"4C", -- 0x2518
    x"00",x"11",x"36",x"25",x"E7",x"3E",x"C0",x"CD", -- 0x2520
    x"4C",x"00",x"11",x"4A",x"25",x"E7",x"3E",x"80", -- 0x2528
    x"CD",x"4C",x"00",x"C3",x"3C",x"1F",x"04",x"14", -- 0x2530
    x"04",x"46",x"49",x"52",x"53",x"54",x"40",x"43", -- 0x2538
    x"52",x"45",x"44",x"49",x"54",x"40",x"34",x"30", -- 0x2540
    x"43",x"FF",x"05",x"18",x"04",x"46",x"55",x"52", -- 0x2548
    x"54",x"48",x"45",x"52",x"40",x"43",x"52",x"45", -- 0x2550
    x"44",x"49",x"54",x"53",x"40",x"32",x"30",x"43", -- 0x2558
    x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2560
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2568
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2570
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2578
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2580
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2588
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2590
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2598
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x25A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x25A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x25B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x25B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x25C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x25C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x25D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x25D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x25E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x25E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x25F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x25F8
    x"3A",x"A0",x"40",x"3C",x"32",x"A0",x"40",x"FD", -- 0x2600
    x"7E",x"04",x"4F",x"E6",x"03",x"B7",x"20",x"02", -- 0x2608
    x"3E",x"02",x"5F",x"FD",x"7E",x"05",x"E6",x"FE", -- 0x2610
    x"57",x"3A",x"00",x"40",x"CB",x"3F",x"CB",x"3F", -- 0x2618
    x"E6",x"01",x"B2",x"FD",x"77",x"05",x"FD",x"7E", -- 0x2620
    x"00",x"FE",x"20",x"30",x"02",x"CB",x"E1",x"FE", -- 0x2628
    x"E8",x"38",x"02",x"CB",x"A1",x"FD",x"7E",x"01", -- 0x2630
    x"FE",x"80",x"30",x"02",x"CB",x"91",x"FE",x"E8", -- 0x2638
    x"38",x"13",x"3A",x"0C",x"40",x"B7",x"20",x"0B", -- 0x2640
    x"CD",x"26",x"17",x"3E",x"FF",x"32",x"00",x"78", -- 0x2648
    x"C3",x"41",x"10",x"CB",x"D1",x"3A",x"00",x"40", -- 0x2650
    x"CB",x"77",x"20",x"0E",x"CB",x"61",x"FD",x"7E", -- 0x2658
    x"00",x"20",x"03",x"93",x"18",x"01",x"83",x"FD", -- 0x2660
    x"77",x"00",x"CB",x"51",x"FD",x"7E",x"01",x"28", -- 0x2668
    x"03",x"93",x"18",x"01",x"83",x"FD",x"77",x"01", -- 0x2670
    x"CB",x"51",x"FD",x"7E",x"05",x"28",x"0B",x"CB", -- 0x2678
    x"B7",x"FD",x"77",x"05",x"FD",x"71",x"04",x"C3", -- 0x2680
    x"41",x"10",x"CB",x"F7",x"18",x"F3",x"3A",x"A2", -- 0x2688
    x"40",x"3C",x"32",x"A2",x"40",x"FD",x"7E",x"01", -- 0x2690
    x"2F",x"32",x"00",x"78",x"FD",x"7E",x"05",x"E6", -- 0x2698
    x"3F",x"FE",x"15",x"28",x"50",x"FD",x"7E",x"04", -- 0x26A0
    x"E6",x"03",x"B7",x"20",x"02",x"3E",x"02",x"4F", -- 0x26A8
    x"FD",x"7E",x"01",x"FE",x"80",x"38",x"01",x"3C", -- 0x26B0
    x"5F",x"3A",x"05",x"40",x"E6",x"1F",x"FE",x"04", -- 0x26B8
    x"20",x"27",x"FD",x"66",x"03",x"FD",x"6E",x"02", -- 0x26C0
    x"11",x"20",x"00",x"19",x"7D",x"E6",x"1F",x"FE", -- 0x26C8
    x"1B",x"30",x"10",x"FE",x"04",x"38",x"0C",x"36", -- 0x26D0
    x"32",x"3E",x"FC",x"32",x"00",x"40",x"3E",x"15", -- 0x26D8
    x"FD",x"77",x"05",x"FD",x"7E",x"01",x"C3",x"41", -- 0x26E0
    x"10",x"2F",x"7B",x"81",x"FE",x"F0",x"30",x"12", -- 0x26E8
    x"FD",x"77",x"01",x"18",x"F1",x"3A",x"00",x"40", -- 0x26F0
    x"B7",x"20",x"EB",x"3E",x"14",x"FD",x"77",x"05", -- 0x26F8
    x"18",x"E4",x"CD",x"26",x"17",x"3E",x"FF",x"32", -- 0x2700
    x"00",x"78",x"18",x"DA",x"3A",x"A1",x"40",x"3C", -- 0x2708
    x"32",x"A1",x"40",x"3A",x"00",x"40",x"5F",x"FD", -- 0x2710
    x"7E",x"04",x"4F",x"E6",x"03",x"B7",x"20",x"02", -- 0x2718
    x"3E",x"03",x"57",x"FD",x"7E",x"00",x"CB",x"61", -- 0x2720
    x"20",x"03",x"82",x"18",x"01",x"92",x"FD",x"77", -- 0x2728
    x"00",x"FE",x"08",x"38",x"CD",x"FE",x"F8",x"30", -- 0x2730
    x"C9",x"CB",x"53",x"20",x"04",x"3E",x"12",x"18", -- 0x2738
    x"02",x"3E",x"13",x"CB",x"61",x"28",x"02",x"CB", -- 0x2740
    x"FF",x"FD",x"77",x"05",x"FD",x"66",x"03",x"FD", -- 0x2748
    x"6E",x"02",x"23",x"11",x"20",x"00",x"19",x"7E", -- 0x2750
    x"FE",x"10",x"28",x"02",x"36",x"FA",x"C3",x"41", -- 0x2758
    x"10",x"AF",x"06",x"04",x"D7",x"C9",x"00",x"00"
  );

begin

  p_rom : process
  begin
    wait until rising_edge(CLK);
       DATA <= ROM(to_integer(unsigned(ADDR)));
  end process;
end RTL;
