library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity sound is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of sound is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"21",X"FF",X"FF",X"2D",X"20",X"FD",X"25",X"20",X"FA",X"DB",X"00",X"FE",X"F0",X"28",X"FA",X"3E",
		X"10",X"3D",X"20",X"FD",X"DB",X"00",X"FE",X"F0",X"28",X"EF",X"FE",X"F1",X"20",X"25",X"21",X"80",
		X"01",X"01",X"4F",X"06",X"DD",X"21",X"2A",X"00",X"18",X"4C",X"06",X"02",X"21",X"FF",X"FF",X"2D",
		X"20",X"FD",X"25",X"20",X"05",X"05",X"20",X"02",X"18",X"CF",X"DB",X"00",X"FE",X"F1",X"28",X"EF",
		X"C3",X"09",X"00",X"FE",X"F2",X"C2",X"5B",X"00",X"21",X"50",X"06",X"01",X"8F",X"10",X"DD",X"21",
		X"55",X"00",X"C3",X"76",X"00",X"DB",X"00",X"FE",X"F2",X"28",X"FA",X"FE",X"F3",X"C2",X"09",X"00",
		X"21",X"90",X"10",X"01",X"FF",X"17",X"DD",X"21",X"6D",X"00",X"C3",X"76",X"00",X"DB",X"00",X"FE",
		X"F3",X"28",X"FA",X"C3",X"09",X"00",X"50",X"59",X"7E",X"E6",X"F0",X"D3",X"00",X"3E",X"1B",X"3D",
		X"20",X"FD",X"7E",X"E6",X"0F",X"07",X"07",X"07",X"07",X"D3",X"00",X"3E",X"19",X"3D",X"20",X"FD",
		X"23",X"EB",X"ED",X"52",X"EB",X"20",X"DF",X"DD",X"E9",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",
		X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",
		X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",
		X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",
		X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",
		X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",
		X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",
		X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",
		X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",
		X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",
		X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",
		X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",
		X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",
		X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",
		X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",X"3A",X"00",
		X"88",X"89",X"88",X"88",X"88",X"88",X"88",X"98",X"99",X"99",X"88",X"98",X"88",X"88",X"88",X"88",
		X"89",X"99",X"98",X"98",X"88",X"88",X"87",X"88",X"87",X"78",X"9A",X"AA",X"89",X"88",X"98",X"87",
		X"78",X"78",X"77",X"8B",X"CB",X"87",X"88",X"A8",X"87",X"78",X"87",X"78",X"AC",X"C9",X"87",X"89",
		X"88",X"77",X"87",X"68",X"AD",X"C9",X"87",X"89",X"87",X"67",X"76",X"9C",X"CA",X"77",X"89",X"86",
		X"67",X"77",X"AD",X"C9",X"56",X"99",X"96",X"55",X"6E",X"EC",X"85",X"79",X"87",X"67",X"65",X"EE",
		X"C8",X"37",X"9A",X"75",X"76",X"8F",X"CB",X"53",X"88",X"95",X"56",X"4F",X"FA",X"A1",X"89",X"87",
		X"45",X"4D",X"F8",X"B2",X"5B",X"78",X"45",X"5E",X"F7",X"83",X"5C",X"76",X"65",X"5F",X"F8",X"70",
		X"8A",X"94",X"56",X"6F",X"C8",X"50",X"C7",X"83",X"37",X"DF",X"F8",X"05",X"E7",X"71",X"48",X"FF",
		X"63",X"0D",X"8A",X"51",X"3F",X"F6",X"A0",X"89",X"68",X"32",X"EF",X"4C",X"05",X"B5",X"73",X"3B",
		X"FA",X"D2",X"4D",X"4A",X"41",X"BF",X"FD",X"32",X"F4",X"98",X"0D",X"F0",X"F1",X"3D",X"3C",X"51",
		X"FF",X"3D",X"06",X"94",X"F6",X"0F",X"F9",X"A0",X"A5",X"7F",X"36",X"FF",X"F2",X"5B",X"29",X"F0",
		X"FC",X"0F",X"0E",X"24",X"FA",X"3F",X"FC",X"A0",X"D0",X"5F",X"0F",X"F0",X"F0",X"86",X"3A",X"F4",
		X"FF",X"8A",X"0D",X"26",X"D5",X"F8",X"4E",X"0A",X"46",X"A3",X"FA",X"2E",X"3A",X"83",X"E8",X"CF",
		X"0C",X"65",X"C3",X"BA",X"8F",X"07",X"61",X"B8",X"9D",X"6F",X"07",X"80",X"94",X"9E",X"8F",X"14",
		X"A0",X"C3",X"8B",X"5F",X"F6",X"80",X"F5",X"A8",X"0F",X"F6",X"E0",X"D7",X"6F",X"0F",X"F1",X"F0",
		X"A8",X"5C",X"2F",X"F1",X"E0",X"8C",X"6C",X"0F",X"F1",X"C0",X"AC",X"8B",X"0F",X"F4",X"A0",X"8B",
		X"CB",X"0F",X"F3",X"F0",X"98",X"9E",X"0F",X"F0",X"F0",X"BE",X"3D",X"0F",X"F0",X"F0",X"9F",X"27",
		X"2F",X"F0",X"E0",X"CF",X"A4",X"3F",X"F0",X"E0",X"AF",X"67",X"9F",X"F1",X"D0",X"6F",X"64",X"FF",
		X"F4",X"A0",X"BF",X"20",X"FF",X"07",X"42",X"CF",X"70",X"FF",X"0D",X"20",X"EE",X"70",X"FF",X"00",
		X"25",X"FB",X"43",X"FF",X"00",X"07",X"FD",X"31",X"FF",X"09",X"08",X"FB",X"45",X"FF",X"0F",X"00",
		X"F9",X"18",X"FF",X"0F",X"00",X"F2",X"37",X"FF",X"0F",X"06",X"F7",X"0C",X"FF",X"5F",X"0A",X"F4",
		X"0F",X"FF",X"0F",X"0F",X"F4",X"0F",X"FF",X"5D",X"0F",X"E7",X"0F",X"FF",X"2F",X"00",X"F3",X"0F",
		X"FF",X"7F",X"00",X"D0",X"0F",X"F0",X"0E",X"0D",X"F0",X"0F",X"F0",X"0C",X"0F",X"F0",X"0F",X"F0",
		X"0A",X"0F",X"C3",X"0F",X"F0",X"08",X"0F",X"F0",X"0F",X"F0",X"06",X"0F",X"F0",X"3F",X"F0",X"00",
		X"0F",X"A0",X"7F",X"F0",X"00",X"0F",X"F0",X"FF",X"F0",X"00",X"5F",X"60",X"FF",X"F0",X"40",X"0F",
		X"F0",X"FF",X"F0",X"F0",X"EF",X"00",X"FF",X"00",X"F0",X"0F",X"00",X"FF",X"00",X"F0",X"FF",X"05",
		X"FF",X"00",X"40",X"FF",X"07",X"FF",X"00",X"A0",X"FF",X"00",X"FF",X"00",X"01",X"F1",X"0F",X"FF",
		X"00",X"01",X"FF",X"00",X"FF",X"0F",X"06",X"F3",X"0F",X"FF",X"0F",X"00",X"F0",X"0F",X"FF",X"0F",
		X"FB",X"F0",X"0F",X"F0",X"0F",X"00",X"F0",X"0F",X"F0",X"0F",X"0F",X"F0",X"1F",X"F0",X"0D",X"0F",
		X"E0",X"5F",X"F0",X"0F",X"00",X"F0",X"0F",X"F0",X"0F",X"0F",X"F0",X"AF",X"F0",X"0F",X"0F",X"90",
		X"0F",X"F0",X"0E",X"0F",X"A0",X"0F",X"F0",X"0E",X"0F",X"E0",X"0F",X"F0",X"04",X"0F",X"E0",X"FF",
		X"F0",X"0D",X"0E",X"F0",X"BF",X"F0",X"0C",X"2F",X"F0",X"5F",X"F0",X"87",X"1C",X"F0",X"AF",X"F0",
		X"CD",X"2B",X"C0",X"3F",X"F0",X"08",X"AB",X"E2",X"1F",X"F6",X"61",X"1E",X"F2",X"6F",X"B0",X"5A",
		X"4A",X"F1",X"1F",X"F6",X"02",X"DE",X"B4",X"4F",X"FC",X"30",X"4D",X"E4",X"7F",X"F7",X"03",X"8A",
		X"B8",X"48",X"FF",X"00",X"5F",X"C7",X"76",X"FE",X"33",X"49",X"C8",X"74",X"FF",X"60",X"0D",X"DB",
		X"83",X"BF",X"96",X"27",X"7A",X"A6",X"FF",X"50",X"3C",X"BA",X"64",X"9F",X"FC",X"00",X"8F",X"D3",
		X"AE",X"88",X"57",X"68",X"96",X"8D",X"FD",X"10",X"6F",X"B5",X"93",X"9F",X"F0",X"0A",X"F8",X"88",
		X"CF",X"80",X"2B",X"C4",X"88",X"9F",X"F0",X"0C",X"E5",X"75",X"3F",X"F8",X"01",X"AA",X"B8",X"7F",
		X"F1",X"0A",X"C6",X"78",X"6F",X"F7",X"06",X"A8",X"77",X"6A",X"FF",X"30",X"16",X"B9",X"7D",X"FD",
		X"21",X"57",X"88",X"8C",X"FD",X"66",X"26",X"96",X"8A",X"BE",X"E8",X"03",X"88",X"77",X"DF",X"F9",
		X"02",X"55",X"6A",X"BF",X"FD",X"22",X"55",X"58",X"9C",X"FF",X"63",X"44",X"56",X"6C",X"FF",X"74",
		X"66",X"45",X"56",X"FF",X"BA",X"95",X"56",X"33",X"DD",X"9A",X"C9",X"69",X"42",X"BD",X"86",X"AC",
		X"9A",X"75",X"AA",X"64",X"8A",X"8B",X"A5",X"BB",X"85",X"77",X"59",X"A7",X"BD",X"A7",X"89",X"57",
		X"86",X"AA",X"87",X"B9",X"79",X"A7",X"79",X"75",X"98",X"7A",X"A9",X"9A",X"98",X"A7",X"67",X"79",
		X"9A",X"97",X"BA",X"89",X"89",X"88",X"66",X"A8",X"8A",X"AB",X"99",X"75",X"A8",X"68",X"9B",X"AA",
		X"87",X"B8",X"66",X"79",X"8A",X"87",X"BA",X"88",X"99",X"69",X"85",X"99",X"99",X"BC",X"79",X"85",
		X"88",X"86",X"8B",X"9C",X"95",X"88",X"87",X"99",X"6A",X"A8",X"77",X"87",X"AB",X"8A",X"97",X"77",
		X"76",X"8A",X"8C",X"BA",X"77",X"96",X"78",X"69",X"9A",X"A8",X"87",X"99",X"79",X"AA",X"78",X"86",
		X"79",X"88",X"AB",X"89",X"A9",X"97",X"77",X"88",X"78",X"97",X"AB",X"97",X"9B",X"88",X"86",X"67",
		X"88",X"9A",X"99",X"A8",X"89",X"98",X"99",X"79",X"A7",X"68",X"86",X"8A",X"9A",X"CA",X"98",X"86",
		X"78",X"78",X"A9",X"78",X"98",X"AA",X"77",X"A9",X"88",X"87",X"78",X"68",X"BA",X"99",X"87",X"89",
		X"67",X"AA",X"A9",X"87",X"79",X"88",X"A9",X"99",X"77",X"88",X"67",X"AA",X"AA",X"97",X"77",X"66",
		X"8A",X"BB",X"98",X"87",X"67",X"89",X"BB",X"98",X"87",X"67",X"78",X"AB",X"AA",X"A8",X"67",X"67",
		X"99",X"AA",X"A9",X"78",X"67",X"89",X"99",X"A9",X"89",X"77",X"88",X"88",X"A8",X"89",X"88",X"99",
		X"89",X"98",X"79",X"87",X"88",X"9A",X"A8",X"79",X"88",X"88",X"89",X"A8",X"78",X"88",X"99",X"89",
		X"A8",X"89",X"88",X"88",X"89",X"A9",X"89",X"98",X"77",X"78",X"A9",X"89",X"99",X"98",X"78",X"88",
		X"89",X"98",X"98",X"88",X"88",X"89",X"99",X"98",X"89",X"97",X"79",X"99",X"98",X"89",X"88",X"88",
		X"89",X"97",X"88",X"87",X"8A",X"98",X"99",X"88",X"87",X"89",X"98",X"98",X"99",X"87",X"89",X"98",
		X"88",X"88",X"87",X"89",X"A9",X"A9",X"88",X"66",X"69",X"99",X"9A",X"98",X"76",X"69",X"99",X"89",
		X"A8",X"97",X"7A",X"8A",X"78",X"77",X"98",X"89",X"A9",X"9A",X"88",X"98",X"79",X"87",X"88",X"88",
		X"A9",X"87",X"88",X"89",X"99",X"99",X"78",X"78",X"89",X"99",X"A9",X"88",X"87",X"89",X"98",X"99",
		X"88",X"88",X"8A",X"99",X"99",X"88",X"77",X"78",X"89",X"A9",X"89",X"88",X"88",X"88",X"99",X"89",
		X"88",X"88",X"88",X"99",X"88",X"88",X"88",X"88",X"98",X"89",X"98",X"89",X"89",X"99",X"89",X"97",
		X"88",X"89",X"AA",X"9A",X"98",X"88",X"88",X"98",X"89",X"98",X"89",X"88",X"98",X"89",X"98",X"89",
		X"88",X"88",X"89",X"98",X"88",X"77",X"88",X"88",X"98",X"78",X"87",X"88",X"78",X"99",X"89",X"98",
		X"89",X"88",X"99",X"88",X"99",X"99",X"99",X"99",X"88",X"87",X"88",X"88",X"88",X"88",X"88",X"88",
		X"98",X"89",X"88",X"98",X"78",X"88",X"88",X"88",X"77",X"77",X"88",X"79",X"98",X"99",X"99",X"AA",
		X"9A",X"AA",X"AA",X"AA",X"A9",X"99",X"98",X"98",X"88",X"88",X"78",X"87",X"78",X"78",X"88",X"78",
		X"98",X"89",X"99",X"AA",X"AB",X"BA",X"AA",X"AA",X"AA",X"AA",X"A9",X"99",X"88",X"87",X"66",X"54",
		X"45",X"34",X"43",X"34",X"44",X"56",X"67",X"89",X"9A",X"BB",X"BB",X"BB",X"AA",X"AB",X"A9",X"99",
		X"99",X"99",X"89",X"98",X"77",X"88",X"88",X"99",X"AA",X"AA",X"AA",X"AA",X"AA",X"BA",X"AA",X"AA",
		X"A9",X"AA",X"A9",X"99",X"99",X"87",X"78",X"87",X"66",X"66",X"66",X"66",X"66",X"66",X"67",X"78",
		X"88",X"88",X"88",X"99",X"99",X"99",X"99",X"88",X"89",X"88",X"88",X"89",X"88",X"88",X"88",X"99",
		X"9A",X"AA",X"AA",X"AA",X"AA",X"9A",X"A9",X"99",X"98",X"88",X"77",X"77",X"76",X"66",X"66",X"66",
		X"66",X"77",X"77",X"88",X"88",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"99",X"98",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"78",X"87",X"88",X"77",X"77",X"77",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"9A",X"AB",X"A9",X"88",X"78",X"89",X"99",X"98",X"87",X"77",
		X"78",X"88",X"87",X"77",X"77",X"76",X"8C",X"BD",X"C9",X"87",X"67",X"89",X"AA",X"99",X"77",X"77",
		X"89",X"99",X"98",X"88",X"88",X"88",X"88",X"87",X"77",X"77",X"79",X"DD",X"DC",X"87",X"66",X"8A",
		X"AA",X"98",X"87",X"78",X"89",X"99",X"98",X"88",X"88",X"88",X"87",X"77",X"77",X"66",X"9D",X"DC",
		X"C7",X"66",X"69",X"BB",X"A9",X"77",X"67",X"89",X"9A",X"98",X"87",X"77",X"78",X"87",X"66",X"66",
		X"7B",X"FB",X"E8",X"56",X"78",X"CB",X"B9",X"66",X"77",X"9A",X"9A",X"A9",X"87",X"67",X"78",X"87",
		X"55",X"58",X"EF",X"BD",X"66",X"78",X"AB",X"98",X"87",X"98",X"98",X"88",X"A8",X"98",X"77",X"66",
		X"55",X"56",X"8F",X"CB",X"A4",X"7A",X"8D",X"B8",X"86",X"6A",X"88",X"9A",X"89",X"76",X"65",X"66",
		X"65",X"8C",X"F7",X"E4",X"69",X"7C",X"C8",X"98",X"6C",X"7A",X"A6",X"97",X"77",X"55",X"45",X"7B",
		X"F8",X"D5",X"28",X"79",X"E8",X"BA",X"6A",X"87",X"86",X"88",X"66",X"44",X"49",X"FF",X"9D",X"06",
		X"67",X"DA",X"BB",X"8A",X"85",X"93",X"85",X"57",X"36",X"9F",X"FB",X"C1",X"66",X"6D",X"9C",X"A7",
		X"B7",X"78",X"56",X"44",X"46",X"CF",X"CD",X"71",X"85",X"9D",X"DE",X"97",X"63",X"84",X"75",X"35",
		X"5C",X"F8",X"F5",X"5A",X"3B",X"BB",X"E6",X"A4",X"57",X"43",X"12",X"7D",X"F9",X"F4",X"5A",X"4D",
		X"AA",X"C9",X"96",X"75",X"31",X"05",X"BF",X"D9",X"80",X"B5",X"DF",X"8D",X"89",X"45",X"43",X"21",
		X"7F",X"FF",X"F0",X"B5",X"7F",X"4E",X"79",X"93",X"70",X"00",X"4E",X"FF",X"F0",X"84",X"8F",X"4F",
		X"4B",X"64",X"60",X"30",X"9F",X"FF",X"90",X"C0",X"F6",X"BD",X"4C",X"09",X"02",X"46",X"FF",X"F9",
		X"0A",X"0F",X"7E",X"A6",X"70",X"80",X"33",X"CF",X"BF",X"09",X"1B",X"98",X"D6",X"A1",X"52",X"36",
		X"FE",X"FE",X"3A",X"49",X"99",X"D6",X"50",X"11",X"5F",X"FF",X"F9",X"C1",X"82",X"A8",X"79",X"18",
		X"0E",X"9E",X"CC",X"CA",X"86",X"A6",X"62",X"37",X"6E",X"F8",X"F4",X"B5",X"8B",X"6D",X"25",X"16",
		X"CE",X"DF",X"5C",X"2A",X"56",X"72",X"87",X"DF",X"8F",X"0D",X"0E",X"58",X"40",X"A6",X"F7",X"F1",
		X"B3",X"97",X"46",X"0D",X"7F",X"AF",X"17",X"29",X"56",X"53",X"DB",X"F9",X"F0",X"72",X"87",X"45",
		X"6A",X"FE",X"F3",X"80",X"93",X"63",X"AA",X"FF",X"F5",X"52",X"36",X"59",X"9E",X"FE",X"B7",X"61",
		X"31",X"5A",X"FF",X"FC",X"54",X"23",X"33",X"8C",X"FF",X"FA",X"63",X"22",X"25",X"AE",X"FE",X"D6",
		X"71",X"31",X"4A",X"CF",X"EF",X"59",X"04",X"02",X"AA",X"FD",X"F7",X"92",X"10",X"19",X"AF",X"CF",
		X"6B",X"03",X"12",X"A9",X"FC",X"F5",X"90",X"31",X"3A",X"BF",X"DF",X"69",X"12",X"02",X"9B",X"FD",
		X"F7",X"A1",X"30",X"57",X"DF",X"FF",X"8A",X"03",X"05",X"8E",X"FF",X"D9",X"60",X"10",X"78",X"FF",
		X"F9",X"A3",X"20",X"09",X"9F",X"DF",X"5B",X"03",X"02",X"7C",X"06",X"F8",X"90",X"20",X"06",X"EF",
		X"FF",X"97",X"01",X"05",X"8F",X"FF",X"DB",X"30",X"00",X"68",X"FF",X"FB",X"C2",X"30",X"36",X"AF",
		X"FE",X"C8",X"42",X"03",X"5D",X"DF",X"CF",X"55",X"02",X"37",X"ED",X"FC",X"E3",X"30",X"14",X"BF",
		X"FF",X"E8",X"50",X"00",X"5D",X"EF",X"CF",X"45",X"01",X"27",X"EE",X"FC",X"C4",X"40",X"14",X"AF",
		X"FF",X"F6",X"60",X"11",X"6C",X"EF",X"EC",X"63",X"11",X"39",X"DF",X"FF",X"67",X"02",X"07",X"CF",
		X"FF",X"C5",X"30",X"13",X"9C",X"FE",X"F5",X"60",X"11",X"7D",X"FF",X"FB",X"61",X"00",X"4A",X"EF",
		X"FF",X"44",X"01",X"38",X"DF",X"FF",X"85",X"00",X"06",X"CF",X"FF",X"E4",X"20",X"02",X"9F",X"FF",
		X"F7",X"60",X"00",X"6C",X"FF",X"FE",X"52",X"00",X"27",X"FF",X"FF",X"77",X"00",X"05",X"CF",X"FF",
		X"E6",X"10",X"03",X"8F",X"FF",X"F6",X"50",X"00",X"5C",X"FF",X"FB",X"60",X"00",X"5A",X"FF",X"FF",
		X"45",X"01",X"27",X"DF",X"FF",X"85",X"00",X"05",X"BF",X"FF",X"F5",X"20",X"02",X"8E",X"FF",X"F9",
		X"50",X"00",X"5B",X"FF",X"FF",X"62",X"00",X"37",X"EF",X"FF",X"85",X"00",X"05",X"BF",X"FF",X"E6",
		X"20",X"02",X"7D",X"FF",X"FA",X"50",X"00",X"5B",X"FF",X"FD",X"71",X"00",X"37",X"EF",X"FF",X"95",
		X"00",X"14",X"BE",X"FF",X"E7",X"10",X"03",X"7D",X"FF",X"FB",X"60",X"00",X"49",X"DF",X"FE",X"73",
		X"01",X"36",X"CF",X"FF",X"B6",X"10",X"14",X"9D",X"FF",X"F9",X"41",X"03",X"5B",X"EF",X"FD",X"72",
		X"00",X"48",X"CF",X"FF",X"A5",X"10",X"25",X"AD",X"FF",X"D8",X"31",X"24",X"8C",X"FF",X"EA",X"41",
		X"02",X"6B",X"FF",X"FB",X"62",X"01",X"59",X"EF",X"FD",X"73",X"01",X"38",X"DF",X"FF",X"93",X"00",
		X"26",X"CF",X"FF",X"A4",X"10",X"26",X"AF",X"FF",X"C6",X"10",X"15",X"9E",X"FF",X"D7",X"20",X"14",
		X"8D",X"FF",X"E9",X"30",X"13",X"7C",X"FF",X"FA",X"41",X"02",X"6B",X"FF",X"FB",X"51",X"02",X"5A",
		X"FF",X"FC",X"72",X"01",X"5A",X"EF",X"FC",X"73",X"12",X"59",X"DF",X"FC",X"83",X"11",X"48",X"DF",
		X"FD",X"84",X"11",X"38",X"CF",X"FD",X"94",X"21",X"37",X"BF",X"FE",X"95",X"21",X"37",X"BE",X"FE",
		X"A5",X"21",X"36",X"BE",X"FE",X"B6",X"31",X"36",X"AE",X"FF",X"B6",X"31",X"25",X"9D",X"FF",X"C8",
		X"42",X"25",X"9D",X"FF",X"C8",X"42",X"24",X"8C",X"FF",X"D9",X"52",X"24",X"7B",X"EF",X"DA",X"52",
		X"13",X"7B",X"EF",X"EA",X"62",X"13",X"6A",X"DF",X"EB",X"73",X"23",X"59",X"CF",X"FD",X"84",X"22",
		X"48",X"CF",X"FE",X"A5",X"21",X"36",X"AE",X"FE",X"B7",X"31",X"25",X"9D",X"FF",X"D9",X"42",X"24",
		X"7B",X"EF",X"EB",X"63",X"23",X"69",X"DF",X"FC",X"84",X"22",X"47",X"BE",X"FE",X"B7",X"32",X"35",
		X"9C",X"EE",X"D9",X"53",X"24",X"7A",X"CE",X"EB",X"85",X"33",X"57",X"AC",X"DD",X"A8",X"54",X"46",
		X"8A",X"CC",X"CA",X"75",X"55",X"78",X"AB",X"BB",X"A8",X"76",X"67",X"88",X"99",X"AA",X"98",X"87",
		X"77",X"78",X"8A",X"AB",X"A8",X"76",X"66",X"78",X"9B",X"CB",X"A8",X"76",X"55",X"78",X"AC",X"CB",
		X"97",X"65",X"56",X"7A",X"BC",X"CA",X"86",X"55",X"67",X"9A",X"BC",X"B9",X"75",X"56",X"78",X"AB",
		X"BA",X"98",X"76",X"78",X"99",X"99",X"88",X"88",X"89",X"99",X"98",X"77",X"78",X"9A",X"AA",X"A8",
		X"76",X"66",X"89",X"AB",X"BA",X"87",X"66",X"67",X"9A",X"BB",X"A9",X"87",X"66",X"78",X"9A",X"AA",
		X"98",X"77",X"78",X"89",X"99",X"98",X"88",X"88",X"98",X"88",X"88",X"88",X"89",X"99",X"98",X"77",
		X"77",X"89",X"9A",X"A9",X"87",X"77",X"88",X"9A",X"A9",X"98",X"77",X"78",X"9A",X"AA",X"98",X"77",
		X"77",X"89",X"AA",X"A9",X"87",X"77",X"88",X"9A",X"A9",X"88",X"77",X"88",X"99",X"99",X"98",X"88",
		X"88",X"89",X"99",X"98",X"88",X"88",X"89",X"99",X"98",X"88",X"88",X"89",X"99",X"98",X"88",X"88",
		X"89",X"99",X"98",X"88",X"88",X"89",X"99",X"99",X"88",X"88",X"88",X"99",X"99",X"88",X"88",X"88",
		X"99",X"99",X"98",X"88",X"88",X"88",X"88",X"88",X"88",X"99",X"99",X"88",X"87",X"88",X"89",X"99",
		X"99",X"88",X"77",X"88",X"99",X"99",X"98",X"77",X"78",X"89",X"99",X"98",X"87",X"77",X"88",X"99",
		X"99",X"88",X"88",X"88",X"99",X"99",X"98",X"88",X"88",X"89",X"99",X"98",X"88",X"88",X"89",X"99",
		X"98",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"99",X"88",X"88",
		X"88",X"88",X"99",X"99",X"98",X"88",X"88",X"88",X"99",X"98",X"88",X"88",X"88",X"88",X"99",X"99",
		X"88",X"88",X"88",X"88",X"99",X"98",X"88",X"88",X"88",X"89",X"99",X"98",X"88",X"88",X"88",X"89",
		X"98",X"88",X"88",X"88",X"88",X"89",X"98",X"88",X"88",X"88",X"88",X"88",X"89",X"99",X"98",X"88",
		X"88",X"88",X"99",X"99",X"88",X"88",X"88",X"89",X"99",X"99",X"88",X"88",X"88",X"99",X"99",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"89",X"88",X"88",X"88",
		X"88",X"99",X"98",X"88",X"88",X"88",X"88",X"99",X"88",X"88",X"88",X"88",X"99",X"98",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"89",X"99",X"88",X"88",X"88",X"88",X"98",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"99",X"99",X"88",X"88",X"88",X"88",X"99",X"99",X"88",
		X"88",X"88",X"89",X"99",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"89",X"88",X"88",X"88",X"88",X"88",X"98",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"89",X"89",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"98",X"88",X"89",X"98",X"89",X"88",
		X"88",X"89",X"89",X"89",X"99",X"87",X"88",X"89",X"88",X"88",X"89",X"89",X"88",X"88",X"89",X"99",
		X"88",X"88",X"88",X"88",X"98",X"88",X"98",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"89",X"99",
		X"98",X"88",X"88",X"89",X"89",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"99",X"99",X"98",X"88",X"98",X"98",X"88",X"88",X"88",X"99",X"99",X"99",X"99",X"98",
		X"88",X"77",X"77",X"78",X"89",X"9A",X"AA",X"AA",X"99",X"87",X"77",X"66",X"77",X"88",X"9A",X"AA",
		X"AA",X"A9",X"88",X"77",X"66",X"67",X"78",X"89",X"AA",X"BB",X"AA",X"99",X"87",X"66",X"66",X"67",
		X"78",X"9A",X"AB",X"BB",X"A9",X"87",X"76",X"66",X"66",X"78",X"89",X"AB",X"BB",X"BB",X"A9",X"87",
		X"66",X"66",X"67",X"78",X"9A",X"AB",X"BB",X"BA",X"98",X"77",X"66",X"66",X"67",X"77",X"99",X"AA",
		X"BB",X"BA",X"A9",X"87",X"76",X"66",X"67",X"78",X"89",X"AB",X"BB",X"BA",X"A8",X"97",X"87",X"87",
		X"88",X"88",X"77",X"77",X"78",X"89",X"AA",X"AA",X"A9",X"99",X"98",X"88",X"87",X"66",X"66",X"68",
		X"8A",X"BB",X"CB",X"B9",X"A8",X"97",X"87",X"87",X"77",X"66",X"67",X"79",X"9B",X"AC",X"BB",X"A9",
		X"88",X"87",X"87",X"87",X"76",X"76",X"77",X"99",X"BB",X"CB",X"BA",X"99",X"78",X"78",X"78",X"78",
		X"77",X"77",X"78",X"99",X"BA",X"CA",X"B9",X"98",X"87",X"88",X"78",X"78",X"77",X"67",X"78",X"9A",
		X"BB",X"CA",X"B9",X"A7",X"87",X"87",X"88",X"88",X"77",X"67",X"78",X"99",X"BA",X"CA",X"B8",X"97",
		X"87",X"87",X"88",X"78",X"77",X"66",X"77",X"99",X"CB",X"DA",X"C9",X"97",X"87",X"78",X"78",X"78",
		X"67",X"66",X"77",X"A8",X"CA",X"DA",X"B9",X"88",X"77",X"68",X"79",X"79",X"77",X"66",X"76",X"99",
		X"BC",X"CD",X"AB",X"79",X"68",X"68",X"88",X"88",X"87",X"75",X"57",X"6A",X"9D",X"BD",X"BB",X"97",
		X"86",X"86",X"87",X"98",X"88",X"66",X"56",X"77",X"B9",X"EA",X"E9",X"B8",X"77",X"68",X"69",X"79",
		X"89",X"86",X"65",X"67",X"7A",X"9D",X"AD",X"AA",X"97",X"86",X"86",X"87",X"98",X"88",X"66",X"56",
		X"77",X"9A",X"BD",X"BD",X"9B",X"69",X"67",X"77",X"88",X"98",X"97",X"76",X"56",X"87",X"BA",X"EB",
		X"DB",X"A9",X"68",X"57",X"68",X"88",X"A8",X"96",X"85",X"65",X"87",X"B9",X"EB",X"DB",X"A9",X"68",
		X"47",X"68",X"89",X"A9",X"A7",X"75",X"54",X"86",X"BA",X"EC",X"CD",X"8A",X"47",X"47",X"77",X"A8",
		X"B9",X"A7",X"75",X"44",X"57",X"8D",X"AF",X"AF",X"9A",X"65",X"65",X"77",X"8A",X"9C",X"9A",X"77",
		X"54",X"46",X"78",X"DA",X"FB",X"F9",X"A6",X"56",X"47",X"88",X"B9",X"C9",X"A7",X"65",X"33",X"37",
		X"6D",X"BF",X"ED",X"D7",X"A2",X"63",X"67",X"8B",X"BC",X"C9",X"95",X"63",X"33",X"48",X"8F",X"CF",
		X"DE",X"A7",X"72",X"43",X"68",X"AC",X"CC",X"C9",X"84",X"52",X"22",X"59",X"9F",X"DF",X"FD",X"C4",
		X"70",X"42",X"78",X"CB",X"FC",X"D8",X"85",X"33",X"12",X"47",X"AC",X"FD",X"FA",X"E5",X"52",X"14",
		X"59",X"BE",X"EF",X"BB",X"66",X"23",X"22",X"35",X"9B",X"EF",X"DF",X"8D",X"36",X"23",X"56",X"AC",
		X"DE",X"DB",X"96",X"53",X"34",X"34",X"58",X"BA",X"FB",X"FA",X"C8",X"55",X"24",X"68",X"CC",X"EE",
		X"CB",X"76",X"44",X"44",X"35",X"4B",X"8F",X"FD",X"F9",X"D5",X"54",X"24",X"68",X"DC",X"FD",X"BB",
		X"67",X"34",X"44",X"34",X"3A",X"7E",X"FD",X"F9",X"D7",X"44",X"24",X"67",X"CE",X"DF",X"BC",X"76",
		X"43",X"44",X"44",X"46",X"B9",X"FE",X"EF",X"9C",X"54",X"43",X"59",X"8E",X"DD",X"F8",X"B4",X"54",
		X"35",X"65",X"64",X"7A",X"8E",X"ED",X"F9",X"C6",X"55",X"45",X"88",X"CE",X"BE",X"8A",X"65",X"54",
		X"57",X"56",X"44",X"98",X"AF",X"BF",X"E9",X"C3",X"64",X"56",X"98",X"EB",X"CB",X"79",X"57",X"56",
		X"67",X"45",X"25",X"88",X"EF",X"FF",X"CB",X"85",X"44",X"37",X"7A",X"CB",X"DB",X"A8",X"76",X"66",
		X"55",X"33",X"25",X"99",X"FF",X"FF",X"DB",X"75",X"34",X"36",X"8A",X"DD",X"DC",X"A9",X"76",X"55",
		X"45",X"44",X"34",X"9A",X"EF",X"FF",X"DB",X"75",X"23",X"35",X"9A",X"DD",X"DD",X"A9",X"76",X"45",
		X"55",X"54",X"54",X"8B",X"CF",X"FF",X"FB",X"87",X"33",X"44",X"79",X"AE",X"CC",X"C8",X"86",X"54",
		X"55",X"65",X"55",X"59",X"AC",X"FF",X"EF",X"A9",X"64",X"34",X"47",X"AA",X"ED",X"DC",X"97",X"64",
		X"46",X"57",X"66",X"55",X"7A",X"AE",X"FE",X"FB",X"97",X"43",X"44",X"69",X"AD",X"ED",X"CA",X"76",
		X"54",X"56",X"67",X"66",X"55",X"8A",X"BF",X"FE",X"FA",X"85",X"32",X"44",X"8A",X"BE",X"EC",X"B8",
		X"65",X"55",X"68",X"78",X"75",X"44",X"8A",X"BF",X"FF",X"FB",X"85",X"31",X"43",X"8A",X"CE",X"FC",
		X"B9",X"56",X"45",X"68",X"79",X"76",X"54",X"5A",X"9D",X"FD",X"FC",X"A5",X"50",X"35",X"6B",X"CD",
		X"DE",X"9A",X"65",X"56",X"78",X"98",X"96",X"53",X"24",X"99",X"EF",X"EF",X"D9",X"56",X"13",X"56",
		X"AC",X"EC",X"EA",X"97",X"65",X"77",X"79",X"78",X"75",X"33",X"26",X"AB",X"FF",X"FF",X"D7",X"64",
		X"14",X"58",X"AD",X"CD",X"CA",X"88",X"66",X"77",X"88",X"77",X"64",X"32",X"26",X"BD",X"FF",X"FF",
		X"C7",X"32",X"01",X"57",X"BE",X"FE",X"EB",X"86",X"54",X"56",X"78",X"88",X"76",X"53",X"24",X"9D",
		X"FF",X"FF",X"E9",X"41",X"10",X"36",X"BD",X"FF",X"DB",X"85",X"34",X"46",X"8A",X"AA",X"96",X"54",
		X"22",X"49",X"EF",X"FF",X"FC",X"73",X"01",X"05",X"9E",X"FF",X"FB",X"95",X"52",X"56",X"8A",X"BA",
		X"88",X"55",X"44",X"35",X"7C",X"FF",X"FF",X"D8",X"62",X"13",X"48",X"AF",X"EF",X"C9",X"65",X"54",
		X"68",X"AA",X"BA",X"87",X"54",X"45",X"45",X"69",X"DE",X"FF",X"EC",X"87",X"43",X"56",X"8A",X"CB",
		X"B9",X"85",X"56",X"78",X"AB",X"AA",X"97",X"55",X"55",X"56",X"66",X"8B",X"EE",X"FF",X"DA",X"76",
		X"23",X"35",X"7A",X"CC",X"DB",X"A7",X"76",X"76",X"89",X"99",X"98",X"77",X"76",X"67",X"65",X"79",
		X"DE",X"FF",X"C9",X"65",X"23",X"47",X"AC",X"FE",X"C9",X"84",X"34",X"57",X"9C",X"CC",X"A9",X"76",
		X"65",X"55",X"66",X"56",X"8C",X"DE",X"FE",X"C9",X"74",X"33",X"67",X"9B",X"CC",X"BA",X"86",X"56",
		X"78",X"AA",X"BA",X"97",X"66",X"66",X"67",X"77",X"67",X"9E",X"EE",X"FD",X"95",X"53",X"34",X"8B",
		X"CE",X"EC",X"87",X"54",X"35",X"79",X"CC",X"CA",X"97",X"66",X"66",X"67",X"77",X"66",X"7A",X"DC",
		X"ED",X"D8",X"76",X"55",X"6A",X"AB",X"BC",X"97",X"65",X"54",X"79",X"BD",X"DD",X"A9",X"65",X"44",
		X"45",X"68",X"98",X"88",X"AD",X"CC",X"CD",X"97",X"66",X"55",X"89",X"AA",X"CB",X"98",X"77",X"67",
		X"89",X"AA",X"BA",X"98",X"87",X"77",X"76",X"66",X"66",X"66",X"AD",X"DD",X"DD",X"97",X"65",X"55",
		X"89",X"AA",X"BA",X"87",X"67",X"67",X"8A",X"BB",X"CB",X"96",X"65",X"55",X"67",X"78",X"88",X"76",
		X"9C",X"CD",X"DE",X"A7",X"55",X"44",X"79",X"BB",X"CB",X"97",X"55",X"56",X"69",X"BC",X"CC",X"B8",
		X"75",X"55",X"56",X"78",X"88",X"87",X"9C",X"DD",X"CD",X"B8",X"55",X"55",X"68",X"AB",X"BB",X"A8",
		X"66",X"67",X"78",X"AB",X"BA",X"A8",X"76",X"66",X"66",X"78",X"87",X"77",X"79",X"CD",X"DC",X"DA",
		X"85",X"56",X"67",X"8B",X"BB",X"A9",X"76",X"55",X"77",X"9B",X"DC",X"BA",X"87",X"55",X"56",X"67",
		X"89",X"98",X"87",X"8B",X"CC",X"BC",X"B8",X"65",X"66",X"78",X"BC",X"BA",X"98",X"66",X"57",X"89",
		X"9B",X"CB",X"A8",X"87",X"66",X"67",X"77",X"78",X"78",X"77",X"AC",X"DC",X"CC",X"A8",X"56",X"67",
		X"78",X"BB",X"A8",X"87",X"76",X"78",X"99",X"9B",X"BA",X"87",X"77",X"66",X"78",X"88",X"78",X"87",
		X"66",X"8C",X"DC",X"BC",X"B9",X"65",X"67",X"88",X"AB",X"A9",X"87",X"77",X"67",X"89",X"AA",X"AA",
		X"A8",X"88",X"87",X"67",X"77",X"66",X"78",X"88",X"79",X"CD",X"CA",X"BA",X"96",X"56",X"78",X"79",
		X"AA",X"98",X"88",X"87",X"77",X"88",X"89",X"9A",X"AA",X"99",X"87",X"66",X"66",X"66",X"78",X"99",
		X"89",X"AB",X"BB",X"AA",X"98",X"66",X"77",X"88",X"9A",X"A9",X"88",X"88",X"77",X"89",X"99",X"99",
		X"A9",X"99",X"98",X"87",X"76",X"66",X"66",X"78",X"9A",X"BC",X"CB",X"A9",X"87",X"66",X"68",X"99",
		X"AA",X"A9",X"87",X"77",X"77",X"89",X"AA",X"99",X"98",X"88",X"99",X"88",X"77",X"66",X"67",X"78",
		X"89",X"AB",X"CB",X"AA",X"98",X"77",X"78",X"89",X"9A",X"99",X"88",X"88",X"88",X"89",X"99",X"98",
		X"88",X"88",X"88",X"99",X"99",X"87",X"76",X"66",X"77",X"89",X"AA",X"BB",X"B9",X"98",X"77",X"77",
		X"89",X"9A",X"99",X"98",X"77",X"78",X"89",X"99",X"99",X"88",X"88",X"88",X"99",X"99",X"87",X"66",
		X"77",X"78",X"99",X"9A",X"AA",X"A9",X"98",X"88",X"78",X"88",X"99",X"99",X"98",X"88",X"88",X"89",
		X"99",X"99",X"88",X"88",X"88",X"99",X"99",X"88",X"87",X"77",X"78",X"88",X"88",X"99",X"9A",X"AA",
		X"99",X"88",X"77",X"78",X"99",X"99",X"99",X"88",X"88",X"88",X"99",X"99",X"98",X"88",X"88",X"88",
		X"89",X"99",X"99",X"98",X"87",X"77",X"77",X"78",X"89",X"99",X"AA",X"AA",X"98",X"87",X"77",X"78",
		X"88",X"88",X"88",X"98",X"88",X"88",X"99",X"98",X"88",X"87",X"89",X"AA",X"A9",X"76",X"66",X"8C",
		X"EC",X"96",X"44",X"68",X"DF",X"D8",X"63",X"46",X"8D",X"FC",X"76",X"43",X"7A",X"9D",X"D9",X"67",
		X"44",X"8A",X"8D",X"D9",X"66",X"35",X"A9",X"BE",X"B6",X"65",X"48",X"B8",X"DC",X"96",X"64",X"69",
		X"9A",X"EC",X"86",X"54",X"8B",X"8D",X"D8",X"56",X"46",X"A9",X"BE",X"A6",X"64",X"5A",X"A7",X"EB",
		X"77",X"64",X"7B",X"7D",X"E8",X"57",X"37",X"C8",X"AF",X"95",X"74",X"4A",X"A9",X"FA",X"46",X"64",
		X"BB",X"5F",X"D5",X"58",X"37",X"C6",X"EF",X"63",X"84",X"7D",X"6A",X"F9",X"37",X"56",X"B7",X"BF",
		X"83",X"66",X"8D",X"59",X"F9",X"45",X"78",X"C5",X"BF",X"75",X"65",X"9C",X"3A",X"F7",X"47",X"6A",
		X"C2",X"CF",X"63",X"84",X"AC",X"3D",X"F4",X"27",X"7B",X"A4",X"FE",X"42",X"68",X"BA",X"9F",X"93",
		X"26",X"BD",X"4B",X"F8",X"33",X"5B",X"C6",X"FC",X"44",X"56",X"E7",X"5F",X"C4",X"35",X"7C",X"5C",
		X"F7",X"46",X"4A",X"B2",X"FE",X"54",X"77",X"B5",X"7F",X"95",X"56",X"9B",X"2F",X"D5",X"47",X"9D",
		X"55",X"F8",X"25",X"8A",X"B5",X"FA",X"43",X"69",X"E6",X"9F",X"73",X"47",X"DA",X"4F",X"A5",X"52",
		X"5F",X"8E",X"E3",X"47",X"5B",X"78",X"F8",X"35",X"48",X"D5",X"FF",X"54",X"44",X"B9",X"CF",X"42",
		X"87",X"97",X"7F",X"B3",X"45",X"6D",X"7F",X"C5",X"75",X"4A",X"6F",X"F4",X"17",X"88",X"47",X"FA",
		X"35",X"48",X"B6",X"FC",X"55",X"78",X"93",X"FE",X"64",X"67",X"B5",X"CF",X"48",X"55",X"B9",X"6F",
		X"64",X"57",X"9A",X"5F",X"91",X"64",X"6D",X"3F",X"F0",X"34",X"7C",X"58",X"F6",X"53",X"2A",X"A4",
		X"F8",X"37",X"49",X"A1",X"FF",X"46",X"47",X"C5",X"AF",X"67",X"47",X"C6",X"5F",X"96",X"54",X"BB",
		X"0F",X"F2",X"81",X"3F",X"82",X"F9",X"64",X"1C",X"D1",X"AF",X"7E",X"00",X"FE",X"1F",X"A7",X"D0",
		X"4F",X"4A",X"F2",X"D0",X"0F",X"90",X"F8",X"CC",X"08",X"E3",X"FF",X"2F",X"00",X"F9",X"2F",X"8E",
		X"D0",X"8B",X"5B",X"F2",X"F0",X"2E",X"83",X"F8",X"F6",X"0A",X"A6",X"FF",X"3F",X"02",X"EB",X"4F",
		X"9E",X"A0",X"89",X"5F",X"F1",X"F0",X"0C",X"B5",X"FB",X"8E",X"08",X"95",X"BF",X"6E",X"60",X"9A",
		X"5F",X"F3",X"F0",X"28",X"4E",X"F6",X"9B",X"0A",X"87",X"8F",X"8F",X"10",X"95",X"BF",X"F2",X"F1",
		X"0B",X"8C",X"8D",X"AF",X"05",X"78",X"CF",X"99",X"60",X"DA",X"C5",X"C8",X"F0",X"08",X"4D",X"DF",
		X"8C",X"07",X"8F",X"48",X"DC",X"D0",X"90",X"D5",X"FE",X"64",X"0A",X"DA",X"2F",X"5F",X"40",X"83",
		X"6C",X"FF",X"C0",X"0F",X"79",X"DB",X"4F",X"07",X"60",X"BF",X"F3",X"F0",X"97",X"DA",X"D5",X"CB",
		X"0F",X"0D",X"6F",X"9E",X"40",X"77",X"F3",X"F7",X"F3",X"37",X"4B",X"5F",X"5F",X"00",X"9B",X"87",
		X"F3",X"F0",X"59",X"08",X"EF",X"7F",X"05",X"79",X"8C",X"F6",X"F0",X"84",X"28",X"EF",X"3F",X"03",
		X"77",X"BB",X"F5",X"F1",X"55",X"1B",X"CF",X"BF",X"03",X"6B",X"A8",X"F5",X"F3",X"46",X"36",X"EF",
		X"1F",X"02",X"3A",X"78",X"FB",X"E6",X"24",X"46",X"BF",X"7F",X"81",X"0D",X"09",X"FD",X"FA",X"03",
		X"60",X"BF",X"FB",X"F0",X"29",X"07",X"CF",X"AF",X"35",X"33",X"49",X"FB",X"F8",X"40",X"32",X"9F",
		X"FB",X"E4",X"16",X"06",X"CF",X"FF",X"61",X"30",X"99",X"ED",X"FA",X"64",X"26",X"3E",X"EE",X"B6",
		X"36",X"66",X"D7",X"F8",X"B5",X"47",X"5B",X"CB",X"6A",X"76",X"88",X"69",X"A9",X"C8",X"57",X"88",
		X"89",X"88",X"9B",X"79",X"A5",X"9A",X"88",X"A5",X"9A",X"87",X"87",X"9C",X"79",X"89",X"69",X"88",
		X"88",X"A8",X"C6",X"77",X"6B",X"98",X"9A",X"5A",X"65",X"A9",X"B8",X"A5",X"B6",X"68",X"9B",X"7C",
		X"89",X"77",X"49",X"E7",X"C7",X"88",X"95",X"7A",X"9D",X"99",X"76",X"55",X"BA",X"D9",X"B5",X"87",
		X"27",X"AE",X"EB",X"54",X"86",X"67",X"DD",X"C7",X"77",X"43",X"7C",X"FD",X"A5",X"67",X"55",X"7D",
		X"DC",X"D6",X"05",X"84",X"AE",X"DC",X"95",X"27",X"36",X"BF",X"FA",X"71",X"65",X"66",X"FD",X"FB",
		X"51",X"27",X"5B",X"FF",X"B8",X"32",X"44",X"7D",X"FF",X"B3",X"23",X"65",X"9F",X"FF",X"84",X"03",
		X"57",X"DF",X"F7",X"53",X"34",X"77",X"FF",X"D8",X"32",X"27",X"7B",X"FE",X"C7",X"30",X"69",X"5E",
		X"FE",X"75",X"03",X"77",X"9F",X"FD",X"61",X"15",X"78",X"CF",X"CB",X"70",X"09",X"94",X"FF",X"E6",
		X"20",X"38",X"B8",X"FF",X"D1",X"13",X"58",X"8D",X"FD",X"86",X"01",X"AA",X"6D",X"FC",X"83",X"03",
		X"AA",X"5F",X"FA",X"42",X"16",X"A7",X"AF",X"F9",X"51",X"19",X"A7",X"AF",X"E7",X"41",X"2A",X"A4",
		X"FF",X"B6",X"30",X"3D",X"A6",X"FF",X"85",X"30",X"5C",X"97",X"FF",X"62",X"02",X"9C",X"7B",X"FB",
		X"46",X"00",X"DD",X"6C",X"F8",X"44",X"03",X"CE",X"7E",X"F6",X"14",X"28",X"E9",X"4F",X"F2",X"64",
		X"0C",X"F6",X"5F",X"D1",X"94",X"0B",X"F7",X"5F",X"C0",X"64",X"6C",X"D3",X"6F",X"93",X"A1",X"3F",
		X"B1",X"BF",X"44",X"B0",X"5E",X"D0",X"BF",X"13",X"B3",X"7F",X"70",X"FF",X"07",X"80",X"BF",X"70",
		X"FF",X"2B",X"60",X"CD",X"52",X"FC",X"09",X"73",X"DB",X"32",X"F7",X"2B",X"37",X"F9",X"07",X"F7",
		X"4B",X"19",X"F7",X"18",X"F4",X"99",X"1B",X"A9",X"0A",X"F5",X"78",X"4B",X"C4",X"0F",X"F1",X"99",
		X"2D",X"B3",X"0F",X"F4",X"A5",X"6B",X"96",X"0F",X"E2",X"97",X"3D",X"C0",X"3F",X"82",X"F4",X"1F",
		X"90",X"AF",X"06",X"F0",X"3F",X"90",X"FF",X"0A",X"E0",X"AE",X"00",X"FF",X"0E",X"A0",X"DD",X"04",
		X"FF",X"2F",X"40",X"FA",X"0E",X"F1",X"6F",X"05",X"F1",X"0F",X"F0",X"CC",X"09",X"F0",X"3F",X"F4",
		X"C6",X"0D",X"F0",X"AF",X"45",X"E3",X"0F",X"40",X"FF",X"0C",X"C0",X"6F",X"00",X"FF",X"2C",X"70",
		X"9F",X"06",X"FF",X"3E",X"50",X"F9",X"0F",X"F0",X"8E",X"02",X"F4",X"0F",X"F0",X"B8",X"08",X"F0",
		X"1F",X"F2",X"B6",X"0E",X"C0",X"FF",X"F4",X"C1",X"1F",X"A0",X"FF",X"16",X"B0",X"4F",X"50",X"FF",
		X"09",X"B0",X"AF",X"08",X"FF",X"1B",X"50",X"CC",X"0F",X"F4",X"3B",X"30",X"FA",X"0F",X"F0",X"4E",
		X"06",X"F1",X"2F",X"F0",X"A9",X"0A",X"E0",X"9F",X"50",X"97",X"0C",X"E0",X"FF",X"20",X"D4",X"3E",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"97",X"01",X"05",X"8F",X"FF",X"DB",X"30",X"00",X"68",X"FF",X"FB",X"C2",X"30",X"36",X"AF",
		X"FE",X"C8",X"42",X"03",X"5D",X"DF",X"CF",X"55",X"02",X"37",X"ED",X"FC",X"E3",X"30",X"14",X"BF",
		X"FF",X"E8",X"50",X"00",X"5D",X"EF",X"CF",X"45",X"01",X"27",X"EE",X"FC",X"C4",X"40",X"14",X"AF",
		X"FF",X"F6",X"60",X"11",X"6C",X"EF",X"EC",X"63",X"11",X"39",X"DF",X"FF",X"67",X"02",X"07",X"CF",
		X"FF",X"C5",X"30",X"13",X"9C",X"FE",X"F5",X"60",X"11",X"7D",X"FF",X"FB",X"61",X"00",X"4A",X"EF",
		X"FF",X"44",X"01",X"38",X"DF",X"FF",X"85",X"00",X"06",X"CF",X"FF",X"E4",X"20",X"02",X"9F",X"FF",
		X"F7",X"60",X"00",X"6C",X"FF",X"FE",X"52",X"00",X"27",X"FF",X"FF",X"77",X"00",X"05",X"CF",X"FF",
		X"E6",X"10",X"03",X"8F",X"FF",X"F6",X"50",X"00",X"5C",X"FF",X"FB",X"60",X"00",X"5A",X"FF",X"FF",
		X"45",X"01",X"27",X"DF",X"FF",X"85",X"00",X"05",X"BF",X"FF",X"F5",X"20",X"02",X"8E",X"FF",X"F9",
		X"50",X"00",X"5B",X"FF",X"FF",X"62",X"00",X"37",X"EF",X"FF",X"85",X"00",X"05",X"BF",X"FF",X"E6",
		X"20",X"02",X"7D",X"FF",X"FA",X"50",X"00",X"5B",X"FF",X"FD",X"71",X"00",X"37",X"EF",X"FF",X"95",
		X"00",X"14",X"BE",X"FF",X"E7",X"10",X"03",X"7D",X"FF",X"FB",X"60",X"00",X"49",X"DF",X"FE",X"73",
		X"01",X"36",X"CF",X"FF",X"B6",X"10",X"14",X"9D",X"FF",X"F9",X"41",X"03",X"5B",X"EF",X"FD",X"72",
		X"00",X"48",X"CF",X"FF",X"A5",X"10",X"25",X"AD",X"FF",X"D8",X"31",X"24",X"8C",X"FF",X"EA",X"41",
		X"02",X"6B",X"FF",X"FB",X"62",X"01",X"59",X"EF",X"FD",X"73",X"01",X"38",X"DF",X"FF",X"93",X"00",
		X"26",X"CF",X"FF",X"A4",X"10",X"26",X"AF",X"FF",X"C6",X"10",X"15",X"9E",X"FF",X"D7",X"20",X"14",
		X"8D",X"FF",X"E9",X"30",X"13",X"7C",X"FF",X"FA",X"41",X"02",X"6B",X"FF",X"FB",X"51",X"02",X"5A",
		X"FF",X"FC",X"72",X"01",X"5A",X"EF",X"FC",X"73",X"12",X"59",X"DF",X"FC",X"83",X"11",X"48",X"DF",
		X"FD",X"84",X"11",X"38",X"CF",X"FD",X"94",X"21",X"37",X"BF",X"FE",X"95",X"21",X"37",X"BE",X"FE",
		X"A5",X"21",X"36",X"BE",X"FE",X"B6",X"31",X"36",X"AE",X"FF",X"B6",X"31",X"25",X"9D",X"FF",X"C8",
		X"42",X"25",X"9D",X"FF",X"C8",X"42",X"24",X"8C",X"FF",X"D9",X"52",X"24",X"7B",X"EF",X"DA",X"52",
		X"13",X"7B",X"EF",X"EA",X"62",X"13",X"6A",X"DF",X"EB",X"73",X"23",X"59",X"CF",X"FD",X"84",X"22",
		X"48",X"CF",X"FE",X"A5",X"21",X"36",X"AE",X"FE",X"B7",X"31",X"25",X"9D",X"FF",X"D9",X"42",X"24",
		X"7B",X"EF",X"EB",X"63",X"23",X"69",X"DF",X"FC",X"84",X"22",X"47",X"BE",X"FE",X"B7",X"32",X"35",
		X"9C",X"EE",X"D9",X"53",X"24",X"7A",X"CE",X"EB",X"85",X"33",X"57",X"AC",X"DD",X"A8",X"54",X"46",
		X"8A",X"CC",X"CA",X"75",X"55",X"78",X"AB",X"BB",X"A8",X"76",X"67",X"88",X"99",X"AA",X"98",X"87",
		X"77",X"78",X"8A",X"AB",X"A8",X"76",X"66",X"78",X"9B",X"CB",X"A8",X"76",X"55",X"78",X"AC",X"CB",
		X"97",X"65",X"56",X"7A",X"BC",X"CA",X"86",X"55",X"67",X"9A",X"BC",X"B9",X"75",X"56",X"78",X"AB",
		X"BA",X"98",X"76",X"78",X"99",X"99",X"88",X"88",X"89",X"99",X"98",X"77",X"78",X"9A",X"AA",X"A8",
		X"76",X"66",X"89",X"AB",X"BA",X"87",X"66",X"67",X"9A",X"BB",X"A9",X"87",X"66",X"78",X"9A",X"AA",
		X"98",X"77",X"78",X"89",X"99",X"98",X"88",X"88",X"98",X"88",X"88",X"88",X"89",X"99",X"98",X"77",
		X"77",X"89",X"9A",X"A9",X"87",X"77",X"88",X"9A",X"A9",X"98",X"77",X"78",X"9A",X"AA",X"98",X"77",
		X"77",X"89",X"AA",X"A9",X"87",X"77",X"88",X"9A",X"A9",X"88",X"77",X"88",X"99",X"99",X"98",X"88",
		X"88",X"89",X"99",X"98",X"88",X"88",X"89",X"99",X"98",X"88",X"88",X"89",X"99",X"98",X"88",X"88",
		X"89",X"99",X"98",X"88",X"88",X"89",X"99",X"99",X"88",X"88",X"88",X"99",X"99",X"88",X"88",X"88",
		X"99",X"99",X"98",X"88",X"88",X"88",X"88",X"88",X"88",X"99",X"99",X"88",X"87",X"88",X"89",X"99",
		X"99",X"88",X"77",X"88",X"99",X"99",X"98",X"77",X"78",X"89",X"99",X"98",X"87",X"77",X"88",X"99",
		X"99",X"88",X"88",X"88",X"99",X"99",X"98",X"88",X"88",X"89",X"99",X"98",X"88",X"88",X"89",X"99",
		X"98",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"99",X"88",X"88",
		X"88",X"88",X"99",X"99",X"98",X"88",X"88",X"88",X"99",X"98",X"88",X"88",X"88",X"88",X"99",X"99",
		X"88",X"88",X"88",X"88",X"99",X"98",X"88",X"88",X"88",X"89",X"99",X"98",X"88",X"88",X"88",X"89",
		X"98",X"88",X"88",X"88",X"88",X"89",X"98",X"88",X"88",X"88",X"88",X"88",X"89",X"99",X"98",X"88",
		X"88",X"88",X"99",X"99",X"88",X"88",X"88",X"89",X"99",X"99",X"88",X"88",X"88",X"99",X"99",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"89",X"88",X"88",X"88",
		X"88",X"99",X"98",X"88",X"88",X"88",X"88",X"99",X"88",X"88",X"88",X"88",X"99",X"98",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"89",X"99",X"88",X"88",X"88",X"88",X"98",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"99",X"99",X"88",X"88",X"88",X"88",X"99",X"99",X"88",
		X"88",X"88",X"89",X"99",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"89",X"88",X"88",X"88",X"88",X"88",X"98",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"89",X"89",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"98",X"88",X"89",X"98",X"89",X"88",
		X"88",X"89",X"89",X"89",X"99",X"87",X"88",X"89",X"88",X"88",X"89",X"89",X"88",X"88",X"89",X"99",
		X"88",X"88",X"88",X"88",X"98",X"88",X"98",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"89",X"99",
		X"98",X"88",X"88",X"89",X"89",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"99",X"99",X"98",X"88",X"98",X"98",X"88",X"88",X"88",X"99",X"99",X"99",X"99",X"98",
		X"88",X"77",X"77",X"78",X"89",X"9A",X"AA",X"AA",X"99",X"87",X"77",X"66",X"77",X"88",X"9A",X"AA",
		X"AA",X"A9",X"88",X"77",X"66",X"67",X"78",X"89",X"AA",X"BB",X"AA",X"99",X"87",X"66",X"66",X"67",
		X"78",X"9A",X"AB",X"BB",X"A9",X"87",X"76",X"66",X"66",X"78",X"89",X"AB",X"BB",X"BB",X"A9",X"87",
		X"66",X"66",X"67",X"78",X"9A",X"AB",X"BB",X"BA",X"98",X"77",X"66",X"66",X"67",X"77",X"99",X"AA",
		X"BB",X"BA",X"A9",X"87",X"76",X"66",X"67",X"78",X"89",X"AB",X"BB",X"BA",X"A8",X"97",X"87",X"87",
		X"88",X"88",X"77",X"77",X"78",X"89",X"AA",X"AA",X"A9",X"99",X"98",X"88",X"87",X"66",X"66",X"68",
		X"8A",X"BB",X"CB",X"B9",X"A8",X"97",X"87",X"87",X"77",X"66",X"67",X"79",X"9B",X"AC",X"BB",X"A9",
		X"88",X"87",X"87",X"87",X"76",X"76",X"77",X"99",X"BB",X"CB",X"BA",X"99",X"78",X"78",X"78",X"78",
		X"77",X"77",X"78",X"99",X"BA",X"CA",X"B9",X"98",X"87",X"88",X"78",X"78",X"77",X"67",X"78",X"9A",
		X"BB",X"CA",X"B9",X"A7",X"87",X"87",X"88",X"88",X"77",X"67",X"78",X"99",X"BA",X"CA",X"B8",X"97",
		X"87",X"87",X"88",X"78",X"77",X"66",X"77",X"99",X"CB",X"DA",X"C9",X"97",X"87",X"78",X"78",X"78",
		X"67",X"66",X"77",X"A8",X"CA",X"DA",X"B9",X"88",X"77",X"68",X"79",X"79",X"77",X"66",X"76",X"99",
		X"BC",X"CD",X"AB",X"79",X"68",X"68",X"88",X"88",X"87",X"75",X"57",X"6A",X"9D",X"BD",X"BB",X"97",
		X"86",X"86",X"87",X"98",X"88",X"66",X"56",X"77",X"B9",X"EA",X"E9",X"B8",X"77",X"68",X"69",X"79",
		X"89",X"86",X"65",X"67",X"7A",X"9D",X"AD",X"AA",X"97",X"86",X"86",X"87",X"98",X"88",X"66",X"56",
		X"77",X"9A",X"BD",X"BD",X"9B",X"69",X"67",X"77",X"88",X"98",X"97",X"76",X"56",X"87",X"BA",X"EB",
		X"DB",X"A9",X"68",X"57",X"68",X"88",X"A8",X"96",X"85",X"65",X"87",X"B9",X"EB",X"DB",X"A9",X"68",
		X"47",X"68",X"89",X"A9",X"A7",X"75",X"54",X"86",X"BA",X"EC",X"CD",X"8A",X"47",X"47",X"77",X"A8",
		X"B9",X"A7",X"75",X"44",X"57",X"8D",X"AF",X"AF",X"9A",X"65",X"65",X"77",X"8A",X"9C",X"9A",X"77",
		X"54",X"46",X"78",X"DA",X"FB",X"F9",X"A6",X"56",X"47",X"88",X"B9",X"C9",X"A7",X"65",X"33",X"37",
		X"6D",X"BF",X"ED",X"D7",X"A2",X"63",X"67",X"8B",X"BC",X"C9",X"95",X"63",X"33",X"48",X"8F",X"CF",
		X"DE",X"A7",X"72",X"43",X"68",X"AC",X"CC",X"C9",X"84",X"52",X"22",X"59",X"9F",X"DF",X"FD",X"C4",
		X"70",X"42",X"78",X"CB",X"FC",X"D8",X"85",X"33",X"12",X"47",X"AC",X"FD",X"FA",X"E5",X"52",X"14",
		X"59",X"BE",X"EF",X"BB",X"66",X"23",X"22",X"35",X"9B",X"EF",X"DF",X"8D",X"36",X"23",X"56",X"AC",
		X"DE",X"DB",X"96",X"53",X"34",X"34",X"58",X"BA",X"FB",X"FA",X"C8",X"55",X"24",X"68",X"CC",X"EE",
		X"CB",X"76",X"44",X"44",X"35",X"4B",X"8F",X"FD",X"F9",X"D5",X"54",X"24",X"68",X"DC",X"FD",X"BB",
		X"67",X"34",X"44",X"34",X"3A",X"7E",X"FD",X"F9",X"D7",X"44",X"24",X"67",X"CE",X"DF",X"BC",X"76",
		X"43",X"44",X"44",X"46",X"B9",X"FE",X"EF",X"9C",X"54",X"43",X"59",X"8E",X"DD",X"F8",X"B4",X"54",
		X"35",X"65",X"64",X"7A",X"8E",X"ED",X"F9",X"C6",X"55",X"45",X"88",X"CE",X"BE",X"8A",X"65",X"54",
		X"57",X"56",X"44",X"98",X"AF",X"BF",X"E9",X"C3",X"64",X"56",X"98",X"EB",X"CB",X"79",X"57",X"56",
		X"67",X"45",X"25",X"88",X"EF",X"FF",X"CB",X"85",X"44",X"37",X"7A",X"CB",X"DB",X"A8",X"76",X"66",
		X"55",X"33",X"25",X"99",X"FF",X"FF",X"DB",X"75",X"34",X"36",X"8A",X"DD",X"DC",X"A9",X"76",X"55",
		X"45",X"44",X"34",X"9A",X"EF",X"FF",X"DB",X"75",X"23",X"35",X"9A",X"DD",X"DD",X"A9",X"76",X"45",
		X"55",X"54",X"54",X"8B",X"CF",X"FF",X"FB",X"87",X"33",X"44",X"79",X"AE",X"CC",X"C8",X"86",X"54",
		X"55",X"65",X"55",X"59",X"AC",X"FF",X"EF",X"A9",X"64",X"34",X"47",X"AA",X"ED",X"DC",X"97",X"64",
		X"46",X"57",X"66",X"55",X"7A",X"AE",X"FE",X"FB",X"97",X"43",X"44",X"69",X"AD",X"ED",X"CA",X"76",
		X"54",X"56",X"67",X"66",X"55",X"8A",X"BF",X"FE",X"FA",X"85",X"32",X"44",X"8A",X"BE",X"EC",X"B8",
		X"65",X"55",X"68",X"78",X"75",X"44",X"8A",X"BF",X"FF",X"FB",X"85",X"31",X"43",X"8A",X"CE",X"FC",
		X"B9",X"56",X"45",X"68",X"79",X"76",X"54",X"5A",X"9D",X"FD",X"FC",X"A5",X"50",X"35",X"6B",X"CD",
		X"DE",X"9A",X"65",X"56",X"78",X"98",X"96",X"53",X"24",X"99",X"EF",X"EF",X"D9",X"56",X"13",X"56",
		X"AC",X"EC",X"EA",X"97",X"65",X"77",X"79",X"78",X"75",X"33",X"26",X"AB",X"FF",X"FF",X"D7",X"64",
		X"14",X"58",X"AD",X"CD",X"CA",X"88",X"66",X"77",X"88",X"77",X"64",X"32",X"26",X"BD",X"FF",X"FF",
		X"C7",X"32",X"01",X"57",X"BE",X"FE",X"EB",X"86",X"54",X"56",X"78",X"88",X"76",X"53",X"24",X"9D",
		X"FF",X"FF",X"E9",X"41",X"10",X"36",X"BD",X"FF",X"DB",X"85",X"34",X"46",X"8A",X"AA",X"96",X"54",
		X"22",X"49",X"EF",X"FF",X"FC",X"73",X"01",X"05",X"9E",X"FF",X"FB",X"95",X"52",X"56",X"8A",X"BA",
		X"88",X"55",X"44",X"35",X"7C",X"FF",X"FF",X"D8",X"62",X"13",X"48",X"AF",X"EF",X"C9",X"65",X"54",
		X"68",X"AA",X"BA",X"87",X"54",X"45",X"45",X"69",X"DE",X"FF",X"EC",X"87",X"43",X"56",X"8A",X"CB",
		X"B9",X"85",X"56",X"78",X"AB",X"AA",X"97",X"55",X"55",X"56",X"66",X"8B",X"EE",X"FF",X"DA",X"76",
		X"23",X"35",X"7A",X"CC",X"DB",X"A7",X"76",X"76",X"89",X"99",X"98",X"77",X"76",X"67",X"65",X"79",
		X"DE",X"FF",X"C9",X"65",X"23",X"47",X"AC",X"FE",X"C9",X"84",X"34",X"57",X"9C",X"CC",X"A9",X"76",
		X"65",X"55",X"66",X"56",X"8C",X"DE",X"FE",X"C9",X"74",X"33",X"67",X"9B",X"CC",X"BA",X"86",X"56",
		X"78",X"AA",X"BA",X"97",X"66",X"66",X"67",X"77",X"67",X"9E",X"EE",X"FD",X"95",X"53",X"34",X"8B",
		X"CE",X"EC",X"87",X"54",X"35",X"79",X"CC",X"CA",X"97",X"66",X"66",X"67",X"77",X"66",X"7A",X"DC",
		X"ED",X"D8",X"76",X"55",X"6A",X"AB",X"BC",X"97",X"65",X"54",X"79",X"BD",X"DD",X"A9",X"65",X"44",
		X"45",X"68",X"98",X"88",X"AD",X"CC",X"CD",X"97",X"66",X"55",X"89",X"AA",X"CB",X"98",X"77",X"67",
		X"89",X"AA",X"BA",X"98",X"87",X"77",X"76",X"66",X"66",X"66",X"AD",X"DD",X"DD",X"97",X"65",X"55",
		X"89",X"AA",X"BA",X"87",X"67",X"67",X"8A",X"BB",X"CB",X"96",X"65",X"55",X"67",X"78",X"88",X"76",
		X"9C",X"CD",X"DE",X"A7",X"55",X"44",X"79",X"BB",X"CB",X"97",X"55",X"56",X"69",X"BC",X"CC",X"B8",
		X"75",X"55",X"56",X"78",X"88",X"87",X"9C",X"DD",X"CD",X"B8",X"55",X"55",X"68",X"AB",X"BB",X"A8",
		X"66",X"67",X"78",X"AB",X"BA",X"A8",X"76",X"66",X"66",X"78",X"87",X"77",X"79",X"CD",X"DC",X"DA",
		X"85",X"56",X"67",X"8B",X"BB",X"A9",X"76",X"55",X"77",X"9B",X"DC",X"BA",X"87",X"55",X"56",X"67",
		X"89",X"98",X"87",X"8B",X"CC",X"BC",X"B8",X"65",X"66",X"78",X"BC",X"BA",X"98",X"66",X"57",X"89",
		X"9B",X"CB",X"A8",X"87",X"66",X"67",X"77",X"78",X"78",X"77",X"AC",X"DC",X"CC",X"A8",X"56",X"67",
		X"78",X"BB",X"A8",X"87",X"76",X"78",X"99",X"9B",X"BA",X"87",X"77",X"66",X"78",X"88",X"78",X"87",
		X"66",X"8C",X"DC",X"BC",X"B9",X"65",X"67",X"88",X"AB",X"A9",X"87",X"77",X"67",X"89",X"AA",X"AA",
		X"A8",X"88",X"87",X"67",X"77",X"66",X"78",X"88",X"79",X"CD",X"CA",X"BA",X"96",X"56",X"78",X"79",
		X"AA",X"98",X"88",X"87",X"77",X"88",X"89",X"9A",X"AA",X"99",X"87",X"66",X"66",X"66",X"78",X"99",
		X"89",X"AB",X"BB",X"AA",X"98",X"66",X"77",X"88",X"9A",X"A9",X"88",X"88",X"77",X"89",X"99",X"99");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
