library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity vid2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of vid2 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"38",X"7C",X"C2",X"82",X"86",X"7C",X"38",X"00",X"02",X"02",X"FE",X"FE",X"42",X"02",X"00",X"00",
		X"62",X"F2",X"BA",X"9A",X"9E",X"CE",X"46",X"00",X"8C",X"DE",X"F2",X"B2",X"92",X"86",X"04",X"00",
		X"08",X"FE",X"FE",X"C8",X"68",X"38",X"18",X"00",X"1C",X"BE",X"A2",X"A2",X"A2",X"E6",X"E4",X"00",
		X"0C",X"9E",X"92",X"92",X"D2",X"7E",X"3C",X"00",X"C0",X"E0",X"B0",X"9E",X"8E",X"C0",X"C0",X"00",
		X"0C",X"6E",X"9A",X"9A",X"B2",X"F2",X"6C",X"00",X"78",X"FC",X"96",X"92",X"92",X"F2",X"60",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"7E",X"C8",X"88",X"C8",X"7E",X"3E",X"00",
		X"6C",X"FE",X"92",X"92",X"92",X"FE",X"FE",X"00",X"44",X"C6",X"82",X"82",X"C6",X"7C",X"38",X"00",
		X"38",X"7C",X"C6",X"82",X"82",X"FE",X"FE",X"00",X"82",X"92",X"92",X"92",X"FE",X"FE",X"00",X"00",
		X"80",X"90",X"90",X"90",X"90",X"FE",X"FE",X"00",X"9E",X"9E",X"92",X"82",X"C6",X"7C",X"38",X"00",
		X"FE",X"FE",X"10",X"10",X"10",X"FE",X"FE",X"00",X"82",X"82",X"FE",X"FE",X"82",X"82",X"00",X"00",
		X"FC",X"FE",X"02",X"02",X"02",X"06",X"04",X"00",X"82",X"C6",X"6E",X"3C",X"18",X"FE",X"FE",X"00",
		X"02",X"02",X"02",X"02",X"FE",X"FE",X"00",X"00",X"FE",X"FE",X"70",X"38",X"70",X"FE",X"FE",X"00",
		X"FE",X"FE",X"1C",X"38",X"70",X"FE",X"FE",X"00",X"7C",X"FE",X"82",X"82",X"82",X"FE",X"7C",X"00",
		X"70",X"F8",X"88",X"88",X"88",X"FE",X"FE",X"00",X"7A",X"FC",X"8E",X"8A",X"82",X"FE",X"7C",X"00",
		X"72",X"F6",X"9E",X"8C",X"88",X"FE",X"FE",X"00",X"0C",X"5E",X"D2",X"92",X"92",X"F6",X"64",X"00",
		X"80",X"80",X"FE",X"FE",X"80",X"80",X"00",X"00",X"FC",X"FE",X"02",X"02",X"02",X"FE",X"FC",X"00",
		X"F0",X"F8",X"1C",X"0E",X"1C",X"F8",X"F0",X"00",X"F8",X"FE",X"1C",X"38",X"1C",X"FE",X"F8",X"00",
		X"C6",X"EE",X"7C",X"38",X"7C",X"EE",X"C6",X"00",X"C0",X"F0",X"1E",X"1E",X"F0",X"C0",X"00",X"00",
		X"C2",X"E2",X"F2",X"BA",X"9E",X"8E",X"86",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"00",X"00",
		X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"00",X"00",X"40",X"40",X"40",X"40",X"40",X"40",X"00",
		X"00",X"00",X"00",X"00",X"28",X"00",X"00",X"00",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",
		X"00",X"00",X"82",X"C6",X"6C",X"38",X"00",X"00",X"00",X"00",X"38",X"6C",X"C6",X"82",X"00",X"00",
		X"00",X"00",X"82",X"FE",X"FE",X"82",X"00",X"00",X"82",X"FE",X"FE",X"82",X"82",X"FE",X"FE",X"82",
		X"00",X"28",X"28",X"28",X"28",X"28",X"28",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"00",
		X"F6",X"F6",X"00",X"00",X"F6",X"F6",X"00",X"00",X"FA",X"FA",X"00",X"00",X"FA",X"FA",X"00",X"00",
		X"00",X"00",X"00",X"F6",X"F6",X"00",X"00",X"00",X"00",X"00",X"00",X"FA",X"FA",X"00",X"00",X"00",
		X"00",X"00",X"00",X"E0",X"C0",X"00",X"00",X"00",X"00",X"E0",X"C0",X"00",X"E0",X"C0",X"00",X"00",
		X"00",X"60",X"E0",X"00",X"60",X"E0",X"00",X"00",X"00",X"00",X"C0",X"00",X"C0",X"00",X"00",X"00",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"FF",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"FF",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"FF",
		X"00",X"00",X"00",X"00",X"06",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"06",X"00",X"00",
		X"38",X"28",X"3E",X"00",X"00",X"00",X"00",X"00",X"3E",X"00",X"3C",X"02",X"02",X"3C",X"00",X"0E",
		X"22",X"2A",X"3E",X"00",X"00",X"0E",X"3A",X"2A",X"22",X"3E",X"00",X"3E",X"08",X"10",X"3E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"22",X"A5",X"BD",X"81",X"42",X"3C",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"3C",X"42",X"81",X"A5",X"FE",X"C2",X"82",X"BA",X"44",X"44",X"28",X"10",
		X"10",X"28",X"44",X"44",X"AA",X"BA",X"82",X"C2",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"45",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A3",X"59",X"FD",X"FD",X"9D",X"8C",X"88",X"00",X"00",X"00",X"01",X"03",X"31",X"59",X"28",X"5C",
		X"00",X"00",X"00",X"00",X"80",X"78",X"FC",X"7F",X"00",X"00",X"07",X"0F",X"0E",X"09",X"07",X"00",
		X"40",X"A0",X"50",X"B0",X"D0",X"68",X"B8",X"50",X"3E",X"9E",X"AE",X"DA",X"CA",X"DE",X"CD",X"D1",
		X"3F",X"7B",X"F1",X"FB",X"7F",X"FF",X"FD",X"78",X"00",X"0C",X"1E",X"3F",X"3F",X"3E",X"3E",X"1C",
		X"B8",X"50",X"A8",X"50",X"B0",X"50",X"A0",X"40",X"D1",X"D1",X"CD",X"DE",X"DA",X"AA",X"BE",X"9E",
		X"7D",X"7F",X"FF",X"FE",X"7C",X"FE",X"7F",X"3F",X"1E",X"3C",X"3E",X"3E",X"3F",X"1E",X"0C",X"00",
		X"00",X"88",X"8C",X"9D",X"FD",X"FD",X"59",X"A3",X"AE",X"1C",X"6D",X"19",X"33",X"01",X"00",X"00",
		X"7F",X"FF",X"7E",X"BE",X"1C",X"00",X"00",X"00",X"00",X"07",X"09",X"0E",X"0F",X"07",X"00",X"00",
		X"45",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"3C",X"7E",X"52",X"4A",X"7E",X"3C",X"00",X"02",X"02",X"FE",X"FE",X"42",X"02",X"00",X"00",
		X"00",X"22",X"72",X"5A",X"4E",X"66",X"22",X"00",X"00",X"44",X"6E",X"7A",X"52",X"46",X"44",X"00",
		X"00",X"04",X"7E",X"7E",X"34",X"1C",X"0C",X"00",X"00",X"4C",X"5E",X"52",X"52",X"76",X"74",X"00",
		X"00",X"0C",X"5E",X"52",X"52",X"7E",X"3C",X"00",X"00",X"60",X"70",X"58",X"4E",X"46",X"40",X"00",
		X"00",X"2C",X"7E",X"52",X"52",X"7E",X"2C",X"00",X"00",X"38",X"7C",X"56",X"52",X"72",X"20",X"00",
		X"7E",X"7E",X"30",X"18",X"30",X"7E",X"7E",X"00",X"1E",X"20",X"20",X"1E",X"20",X"20",X"3E",X"00",
		X"01",X"01",X"01",X"FE",X"01",X"01",X"01",X"00",X"08",X"08",X"08",X"07",X"08",X"08",X"08",X"08",
		X"00",X"00",X"00",X"01",X"01",X"01",X"FE",X"00",X"08",X"08",X"08",X"08",X"08",X"08",X"07",X"00",
		X"00",X"00",X"00",X"07",X"08",X"08",X"08",X"08",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"3F",X"03",X"03",X"3F",X"FF",X"FF",X"A7",X"A7",X"1F",X"1F",X"FF",X"1F",X"A7",X"A7",
		X"00",X"00",X"00",X"00",X"1F",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"7F",X"3B",X"3B",X"3F",X"3D",X"7B",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"04",X"00",X"00",X"10",X"00",
		X"00",X"00",X"00",X"00",X"3F",X"60",X"40",X"40",X"40",X"40",X"40",X"60",X"3F",X"00",X"00",X"00",
		X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"28",X"38",X"FF",X"38",X"28",X"00",
		X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"C7",X"C7",X"C7",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"02",X"04",X"00",X"FF",X"06",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"03",X"02",X"FC",X"FC",X"02",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"24",X"00",X"00",X"24",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"3B",X"61",X"41",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"70",X"7C",X"7E",
		X"7E",X"7C",X"70",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"41",X"61",X"3B",X"03",
		X"FC",X"FC",X"F8",X"F8",X"F0",X"F0",X"60",X"60",X"50",X"88",X"50",X"20",X"50",X"88",X"50",X"20",
		X"50",X"88",X"50",X"20",X"50",X"88",X"50",X"20",X"60",X"60",X"F0",X"F0",X"F8",X"F8",X"FC",X"FC",
		X"00",X"3F",X"40",X"C0",X"C0",X"40",X"40",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"40",X"40",X"C0",X"C0",X"40",X"3F",X"00",X"00",X"FC",X"02",X"03",X"03",X"02",X"02",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"02",X"03",X"03",X"02",X"FC",X"00",
		X"00",X"08",X"0C",X"FC",X"FC",X"00",X"A4",X"A6",X"00",X"C0",X"E8",X"00",X"40",X"A0",X"F8",X"F8",
		X"A0",X"A0",X"B0",X"BF",X"BF",X"B0",X"A0",X"A0",X"1C",X"3E",X"7E",X"7C",X"F8",X"FC",X"FE",X"FE",
		X"FC",X"FE",X"FE",X"FC",X"F8",X"FC",X"FE",X"FE",X"FE",X"FC",X"FC",X"F8",X"7C",X"7E",X"3E",X"1C",
		X"00",X"1F",X"3F",X"70",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",
		X"60",X"60",X"60",X"60",X"70",X"3F",X"1F",X"00",X"06",X"06",X"0E",X"FE",X"FE",X"0E",X"06",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"F0",X"00",X"F0",X"40",X"40",X"E0",X"E0",
		X"00",X"04",X"04",X"FC",X"F8",X"00",X"A8",X"A8",X"E0",X"F8",X"7D",X"01",X"70",X"88",X"FE",X"FE",
		X"00",X"F0",X"F0",X"60",X"60",X"F0",X"F0",X"00",X"81",X"80",X"90",X"80",X"A0",X"A1",X"81",X"81",
		X"00",X"F8",X"FC",X"0E",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",
		X"06",X"06",X"06",X"06",X"0E",X"FC",X"F8",X"00",X"00",X"3C",X"42",X"42",X"42",X"42",X"42",X"42",
		X"42",X"42",X"42",X"42",X"42",X"42",X"3C",X"00",X"00",X"0F",X"0F",X"06",X"06",X"0F",X"0F",X"00",
		X"04",X"08",X"10",X"08",X"04",X"02",X"01",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"90",X"90",X"8A",X"80",X"40",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"81",X"00",X"00",X"18",X"18",X"00",X"00",X"81",X"00",X"00",X"04",X"0A",X"1F",X"17",X"0D",X"06",
		X"38",X"7C",X"C2",X"82",X"86",X"7C",X"38",X"00",X"02",X"02",X"FE",X"FE",X"42",X"02",X"00",X"00",
		X"62",X"F2",X"BA",X"9A",X"9E",X"CE",X"46",X"00",X"8C",X"DE",X"F2",X"B2",X"92",X"86",X"04",X"00",
		X"08",X"FE",X"FE",X"C8",X"68",X"38",X"18",X"00",X"1C",X"BE",X"A2",X"A2",X"A2",X"E6",X"E4",X"00",
		X"0C",X"9E",X"92",X"92",X"D2",X"7E",X"3C",X"00",X"C0",X"E0",X"B0",X"9E",X"8E",X"C0",X"C0",X"00",
		X"0C",X"6E",X"9A",X"9A",X"B2",X"F2",X"6C",X"00",X"78",X"FC",X"96",X"92",X"92",X"F2",X"60",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"7E",X"C8",X"88",X"C8",X"7E",X"3E",X"00",
		X"6C",X"FE",X"92",X"92",X"92",X"FE",X"FE",X"00",X"44",X"C6",X"82",X"82",X"C6",X"7C",X"38",X"00",
		X"38",X"7C",X"C6",X"82",X"82",X"FE",X"FE",X"00",X"82",X"92",X"92",X"92",X"FE",X"FE",X"00",X"00",
		X"80",X"90",X"90",X"90",X"90",X"FE",X"FE",X"00",X"9E",X"9E",X"92",X"82",X"C6",X"7C",X"38",X"00",
		X"FE",X"FE",X"10",X"10",X"10",X"FE",X"FE",X"00",X"82",X"82",X"FE",X"FE",X"82",X"82",X"00",X"00",
		X"FC",X"FE",X"02",X"02",X"02",X"06",X"04",X"00",X"82",X"C6",X"6E",X"3C",X"18",X"FE",X"FE",X"00",
		X"02",X"02",X"02",X"02",X"FE",X"FE",X"00",X"00",X"FE",X"FE",X"70",X"38",X"70",X"FE",X"FE",X"00",
		X"FE",X"FE",X"1C",X"38",X"70",X"FE",X"FE",X"00",X"7C",X"FE",X"82",X"82",X"82",X"FE",X"7C",X"00",
		X"70",X"F8",X"88",X"88",X"88",X"FE",X"FE",X"00",X"7A",X"FC",X"8E",X"8A",X"82",X"FE",X"7C",X"00",
		X"72",X"F6",X"9E",X"8C",X"88",X"FE",X"FE",X"00",X"0C",X"5E",X"D2",X"92",X"92",X"F6",X"64",X"00",
		X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"00",X"FC",X"FE",X"02",X"02",X"02",X"FE",X"FC",X"00",
		X"F0",X"F8",X"1C",X"0E",X"1C",X"F8",X"F0",X"00",X"F8",X"FE",X"1C",X"38",X"1C",X"FE",X"F8",X"00",
		X"C6",X"EE",X"7C",X"38",X"7C",X"EE",X"C6",X"00",X"C0",X"F0",X"1E",X"1E",X"F0",X"C0",X"00",X"00",
		X"C2",X"E2",X"F2",X"BA",X"9E",X"8E",X"86",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"00",X"00",
		X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"00",X"00",X"40",X"40",X"40",X"40",X"40",X"40",X"00",
		X"00",X"00",X"00",X"00",X"28",X"00",X"00",X"00",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",
		X"03",X"0F",X"1F",X"3F",X"3F",X"7F",X"7F",X"7F",X"C0",X"F0",X"F8",X"FC",X"FC",X"FE",X"FE",X"FE",
		X"00",X"03",X"0F",X"1F",X"3F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"F0",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"80",X"81",X"C7",
		X"7F",X"7F",X"3F",X"3F",X"1F",X"7F",X"FF",X"FF",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",X"E7",X"E3",X"E1",X"E0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C3",X"07",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FC",
		X"FF",X"FF",X"FF",X"FE",X"FC",X"FE",X"FF",X"FF",X"E0",X"C0",X"80",X"00",X"00",X"00",X"80",X"C0",
		X"07",X"0F",X"1F",X"1F",X"3F",X"1F",X"1F",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",
		X"FF",X"FF",X"FF",X"FC",X"F0",X"C0",X"00",X"00",X"F0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"E0",X"E1",X"E3",X"E7",X"EF",X"FF",X"FF",X"07",X"07",X"C3",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FC",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FC",X"00",X"00",X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"C0",X"E0",X"F0",X"F8",X"F8",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"F0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"FC",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"3F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FC",X"FC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"3F",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"00",
		X"F8",X"F8",X"F0",X"E0",X"C0",X"00",X"00",X"00",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"00",
		X"3F",X"3F",X"3E",X"7E",X"7C",X"7C",X"7C",X"7C",X"0F",X"06",X"00",X"03",X"07",X"0F",X"1F",X"1F",
		X"3E",X"3C",X"3E",X"3F",X"3F",X"1F",X"1F",X"0F",X"73",X"07",X"0F",X"0F",X"1F",X"1F",X"3F",X"3F",
		X"1F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7C",X"79",X"7F",X"7F",X"7F",X"00",X"00",X"00",X"01",X"07",
		X"3F",X"3F",X"3F",X"00",X"7F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"FF",X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"FF",X"01",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"01",X"00",X"00",X"80",X"8C",X"9F",X"BF",X"FF",X"FF",X"FF",X"BF",X"9F",X"8C",X"80",X"00",
		X"F8",X"F8",X"FF",X"FF",X"FF",X"00",X"7E",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"FE",X"F8",
		X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"00",
		X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",X"F8",X"F0",X"E0",X"40",X"00",X"80",X"C0",X"E0",X"E0",
		X"FC",X"FC",X"FC",X"7C",X"7C",X"78",X"F8",X"F0",X"C8",X"E0",X"F0",X"F0",X"F8",X"78",X"7C",X"7C",
		X"00",X"00",X"F8",X"F8",X"F8",X"F8",X"38",X"98",X"F8",X"F8",X"F8",X"F8",X"E0",X"80",X"00",X"00",
		X"FC",X"FC",X"FC",X"00",X"F8",X"F8",X"F8",X"F8",X"01",X"00",X"00",X"00",X"00",X"3F",X"3F",X"3F",
		X"3C",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"07",X"7C",X"7C",X"7C",X"7F",X"7F",X"7F",X"07",X"31",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"01",X"07",X"0F",X"3F",X"3F",X"3F",X"3F",X"02",
		X"3F",X"3F",X"0F",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"3C",X"3E",X"3F",X"3F",X"3F",
		X"FF",X"FF",X"3C",X"3C",X"3C",X"FF",X"FF",X"FF",X"7E",X"1C",X"C1",X"F3",X"FF",X"FF",X"FF",X"FF",
		X"78",X"78",X"78",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"78",X"78",X"78",X"78",X"78",X"78",
		X"FF",X"FF",X"F8",X"F0",X"E0",X"C0",X"80",X"00",X"E0",X"F0",X"F8",X"FF",X"FF",X"7F",X"7F",X"7F",
		X"00",X"3C",X"7E",X"52",X"4A",X"7E",X"3C",X"00",X"02",X"02",X"FE",X"FE",X"42",X"02",X"00",X"00",
		X"00",X"22",X"72",X"5A",X"4E",X"66",X"22",X"00",X"00",X"44",X"6E",X"7A",X"52",X"46",X"44",X"00",
		X"00",X"04",X"7E",X"7E",X"34",X"1C",X"0C",X"00",X"00",X"4C",X"5E",X"52",X"52",X"76",X"74",X"00",
		X"00",X"0C",X"5E",X"52",X"52",X"7E",X"3C",X"00",X"00",X"60",X"70",X"58",X"4E",X"46",X"40",X"00",
		X"00",X"2C",X"7E",X"52",X"52",X"7E",X"2C",X"00",X"00",X"38",X"7C",X"56",X"52",X"72",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"00",X"00",X"00",X"00",X"FC",X"FC",X"FC",
		X"7C",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"F0",X"F8",X"F8",X"F8",X"F8",X"F8",X"C0",X"9C",X"3C",
		X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"FC",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FC",X"FC",X"FC",X"FC",X"FC",X"7F",X"7F",X"1F",X"07",X"01",X"00",X"00",X"00",
		X"0F",X"0F",X"63",X"78",X"7E",X"7F",X"7F",X"7F",X"3F",X"3E",X"3C",X"3E",X"3F",X"3F",X"1F",X"1F",
		X"79",X"73",X"07",X"0F",X"0F",X"1F",X"1F",X"3F",X"07",X"1F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7C",
		X"7F",X"7F",X"7F",X"7F",X"00",X"00",X"00",X"01",X"1F",X"1F",X"0F",X"0F",X"00",X"7F",X"7F",X"7F",
		X"FF",X"FF",X"FF",X"FF",X"FE",X"78",X"78",X"78",X"BF",X"FF",X"FE",X"FC",X"39",X"83",X"E7",X"FF",
		X"00",X"00",X"01",X"00",X"00",X"80",X"8C",X"9F",X"FF",X"FF",X"FF",X"FF",X"BF",X"9F",X"8C",X"80",
		X"F8",X"F8",X"F8",X"FF",X"FF",X"FF",X"00",X"7E",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"FE",
		X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"F8",X"F8",X"E0",X"80",X"00",X"00",X"00",X"00",
		X"80",X"38",X"78",X"F8",X"F8",X"F8",X"F8",X"F8",X"7C",X"FC",X"FC",X"FC",X"7C",X"7C",X"78",X"F8",
		X"98",X"C8",X"E0",X"F0",X"F0",X"F8",X"78",X"7C",X"00",X"00",X"00",X"F8",X"F8",X"F8",X"F8",X"38",
		X"F8",X"F8",X"F8",X"F8",X"F8",X"E0",X"80",X"00",X"F8",X"F8",X"F0",X"F0",X"00",X"F8",X"F8",X"F8",
		X"3F",X"3F",X"3E",X"3E",X"3E",X"3E",X"3F",X"3F",X"00",X"00",X"03",X"07",X"0F",X"0F",X"1F",X"1F",
		X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"81",X"00",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"88",
		X"F8",X"7C",X"7C",X"7C",X"7C",X"7C",X"FC",X"FC",X"00",X"FC",X"FC",X"FC",X"FC",X"F0",X"F0",X"F0",
		X"C0",X"E0",X"F0",X"F0",X"F8",X"F8",X"FC",X"FC",X"F0",X"F0",X"F0",X"F0",X"60",X"00",X"00",X"80",
		X"00",X"00",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"80",
		X"F0",X"E0",X"00",X"00",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"E0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"E0",X"F8",X"F8",X"F8",X"F8",X"F8",X"F0",X"F0",X"E0",
		X"C0",X"C0",X"E0",X"E0",X"F0",X"F0",X"F8",X"F8",X"F0",X"F0",X"F0",X"F0",X"70",X"20",X"00",X"80",
		X"00",X"00",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"F0",X"60",X"00",X"00",X"80",X"C0",X"C0",X"E0",
		X"F0",X"F0",X"C0",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"60",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"28",X"38",X"FF",X"38",X"28",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"28",X"38",X"FF",X"38",X"28",X"00",
		X"A0",X"A0",X"B0",X"BF",X"BF",X"B0",X"A0",X"A0",X"1C",X"3E",X"7E",X"7C",X"F8",X"FC",X"FE",X"FE",
		X"FC",X"FE",X"FE",X"FC",X"F8",X"FC",X"FE",X"FE",X"FE",X"FC",X"FC",X"F8",X"7C",X"7E",X"3E",X"1C",
		X"00",X"1F",X"3F",X"70",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",
		X"60",X"60",X"60",X"60",X"70",X"3F",X"1F",X"00",X"06",X"06",X"0E",X"FE",X"FE",X"0E",X"06",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"F0",X"00",X"F0",X"40",X"40",X"E0",X"E0",
		X"00",X"04",X"04",X"FC",X"F8",X"00",X"A8",X"A8",X"E0",X"F8",X"7D",X"01",X"70",X"88",X"FE",X"FE",
		X"00",X"F0",X"F0",X"60",X"60",X"F0",X"F0",X"00",X"81",X"80",X"90",X"80",X"A0",X"A1",X"81",X"81",
		X"00",X"F8",X"FC",X"0E",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",
		X"06",X"06",X"06",X"06",X"0E",X"FC",X"F8",X"00",X"00",X"3C",X"42",X"42",X"42",X"42",X"42",X"42",
		X"42",X"42",X"42",X"42",X"42",X"42",X"3C",X"00",X"00",X"0F",X"0F",X"06",X"06",X"0F",X"0F",X"00",
		X"04",X"08",X"10",X"08",X"04",X"02",X"01",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"90",X"90",X"8A",X"80",X"40",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"81",X"00",X"00",X"18",X"18",X"00",X"00",X"81",X"00",X"00",X"04",X"0A",X"1F",X"17",X"0D",X"06");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
