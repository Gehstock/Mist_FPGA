/* Atari on an FPGA
Masters of Engineering Project
Cornell University, 2007
Daniel Beer
 TIA.h
Header file that contains useful definitions for the TIA module.
*/
`define CXM0P 7'h70
`define CXM1P 7'h71
`define CXP0FB 7'h72
`define CXP1FB 7'h73
`define CXM0FB 7'h74
`define CXM1FB 7'h75
`define CXBLPF 7'h76
`define CXPPMM 7'h77
`define INPT0 7'h78
`define INPT1 7'h79
`define INPT2 7'h7A
`define INPT3 7'h7B
`define INPT4 7'h7C
`define INPT5 7'h7D
`define VSYNC 7'h00
`define VBLANK 7'h01
`define WSYNC 7'h02
`define RSYNC 7'h03
`define NUSIZ0 7'h04
`define NUSIZ1 7'h05
`define COLUP0 7'h06
`define COLUP1 7'h07
`define COLUPF 7'h08
`define COLUBK 7'h09
`define CTRLPF 7'h0A
`define REFP0 7'h0B
`define REFP1 7'h0C
`define PF0 7'h0D
`define PF1 7'h0E
`define PF2 7'h0F
`define RESP0 7'h10
`define RESP1 7'h11
`define RESM0 7'h12
`define RESM1 7'h13
`define RESBL 7'h14
`define AUDC0 7'h15
`define AUDC1 7'h16
`define AUDF0 7'h17
`define AUDF1 7'h18
`define AUDV0 7'h19
`define AUDV1 7'h1A
`define GRP0 7'h1B
`define GRP1 7'h1C
`define ENAM0 7'h1D
`define ENAM1 7'h1E
`define ENABL 7'h1F
`define HMP0 7'h20
`define HMP1 7'h21
`define HMM0 7'h22
`define HMM1 7'h23
`define HMBL 7'h24
`define VDELP0 7'h25
`define VDELP1 7'h26
`define VDELBL 7'h27
`define RESMP0 7'h28
`define RESMP1 7'h29
`define HMOVE 7'h2A
`define HMCLR 7'h2B
`define CXCLR 7'h2C

`define CXM0P_7800 7'h40
`define CXM1P_7800 7'h41
`define CXP0FB_7800 7'h42
`define CXP1FB_7800 7'h43
`define CXM0FB_7800 7'h44
`define CXM1FB_7800 7'h45
`define CXBLPF_7800 7'h46
`define CXPPMM_7800 7'h47
`define INPT0_7800 7'h48
`define INPT1_7800 7'h49
`define INPT2_7800 7'h4A
`define INPT3_7800 7'h4B
`define INPT4_7800 7'h4C
`define INPT5_7800 7'h4D