library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity cclimber_tile_bit0 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of cclimber_tile_bit0 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"1F",X"3F",X"40",X"80",X"80",X"80",X"80",X"80",X"F8",X"FC",X"02",X"01",X"01",X"01",X"01",X"01",
		X"80",X"80",X"80",X"80",X"40",X"3F",X"1F",X"00",X"01",X"01",X"01",X"01",X"02",X"FC",X"F8",X"00",
		X"7D",X"65",X"65",X"7D",X"69",X"6D",X"6C",X"00",X"AC",X"AA",X"AA",X"AC",X"AA",X"AA",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FD",X"FB",X"F7",X"EE",X"FF",X"FF",X"FF",X"EF",X"DF",X"BF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FD",X"FB",X"F7",X"EF",X"FF",X"FF",X"FF",X"EF",X"DF",X"BF",X"7F",X"FF",X"FF",
		X"FF",X"FF",X"FE",X"FF",X"FB",X"FF",X"00",X"00",X"FF",X"FF",X"EF",X"DF",X"BF",X"FF",X"00",X"00",
		X"FF",X"FF",X"FE",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",
		X"FF",X"80",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"FF",X"F6",X"ED",X"DB",X"BF",X"EF",X"DF",X"BF",
		X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"80",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",
		X"FF",X"18",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"FF",X"01",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",
		X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",
		X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"18",X"FF",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"01",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"02",X"04",X"08",X"10",X"10",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"08",X"08",X"04",X"04",X"04",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"08",X"10",X"10",X"20",X"10",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"10",X"20",X"20",X"40",X"80",X"80",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"04",X"04",X"0B",X"10",X"20",X"20",X"20",X"C0",X"00",
		X"08",X"10",X"10",X"10",X"20",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"16",X"E0",X"00",X"02",X"04",X"08",X"08",X"10",X"E0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"21",X"16",X"08",X"00",X"00",X"00",X"00",X"1C",X"E2",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"02",X"01",X"20",X"10",X"08",X"00",X"00",X"00",X"00",X"08",X"90",X"A0",X"A0",X"40",X"16",
		X"00",X"0A",X"15",X"20",X"02",X"04",X"00",X"08",X"08",X"40",X"08",X"84",X"82",X"40",X"40",X"00",
		X"00",X"41",X"21",X"00",X"04",X"00",X"10",X"80",X"40",X"00",X"88",X"80",X"10",X"00",X"00",X"04",
		X"40",X"00",X"00",X"09",X"04",X"00",X"10",X"00",X"00",X"00",X"01",X"20",X"18",X"20",X"10",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C0",X"80",X"40",X"A0",X"C0",X"80",X"40",X"A0",
		X"1F",X"0F",X"17",X"0F",X"1F",X"0F",X"17",X"0F",X"FF",X"7D",X"7D",X"83",X"C7",X"D7",X"D7",X"FF",
		X"00",X"00",X"05",X"0E",X"1B",X"0C",X"00",X"00",X"00",X"E0",X"9A",X"6D",X"20",X"00",X"02",X"07",
		X"30",X"70",X"EC",X"30",X"0F",X"04",X"07",X"03",X"01",X"02",X"00",X"00",X"F5",X"2F",X"E6",X"C0",
		X"02",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"A0",X"E0",X"E0",X"C0",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"07",X"07",X"03",X"00",X"00",X"00",X"00",X"F0",X"E0",X"E0",X"C0",
		X"41",X"32",X"0D",X"30",X"50",X"00",X"A8",X"51",X"08",X"04",X"18",X"28",X"00",X"00",X"D2",X"25",
		X"22",X"45",X"00",X"00",X"0F",X"07",X"07",X"03",X"1A",X"05",X"00",X"00",X"F0",X"E0",X"E0",X"C0",
		X"00",X"00",X"05",X"05",X"07",X"0A",X"09",X"0D",X"80",X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"90",
		X"05",X"04",X"02",X"02",X"0F",X"07",X"07",X"03",X"90",X"90",X"A0",X"E0",X"F0",X"E0",X"E0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"0F",X"1D",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"70",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"0F",X"1F",X"3D",X"00",X"00",X"00",X"00",X"80",X"E0",X"F0",X"78",
		X"3F",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"0F",X"1F",X"3D",X"3E",X"1F",X"1F",X"00",X"80",X"E0",X"F0",X"78",X"F8",X"F0",X"F0",
		X"0F",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"1B",X"3F",X"3F",X"1F",X"1F",X"0F",X"03",X"E0",X"70",X"F8",X"F8",X"F0",X"F0",X"E0",X"80",
		X"1F",X"7F",X"FF",X"7F",X"3F",X"00",X"00",X"00",X"F0",X"FC",X"FE",X"FC",X"F8",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",
		X"00",X"08",X"08",X"04",X"02",X"00",X"00",X"00",X"00",X"10",X"10",X"20",X"60",X"C0",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"08",X"05",X"03",X"00",X"00",X"80",X"90",X"CC",X"82",X"BA",X"E9",
		X"09",X"0D",X"15",X"0A",X"02",X"01",X"00",X"00",X"F0",X"B5",X"65",X"E2",X"66",X"48",X"80",X"80",
		X"00",X"00",X"18",X"00",X"20",X"38",X"18",X"09",X"00",X"04",X"04",X"08",X"08",X"18",X"48",X"A0",
		X"12",X"24",X"02",X"03",X"33",X"04",X"00",X"00",X"22",X"E1",X"D1",X"61",X"02",X"1C",X"30",X"10",
		X"00",X"02",X"02",X"04",X"08",X"00",X"00",X"A0",X"00",X"08",X"80",X"10",X"40",X"10",X"0C",X"5C",
		X"09",X"46",X"00",X"34",X"0C",X"2C",X"04",X"00",X"80",X"31",X"08",X"12",X"0E",X"1C",X"11",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"80",X"80",X"80",X"80",X"00",X"C0",X"40",
		X"02",X"02",X"00",X"01",X"00",X"00",X"00",X"00",X"A0",X"40",X"80",X"40",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"02",X"05",X"18",X"1C",X"00",X"00",X"00",X"00",X"A0",X"40",X"30",X"08",X"10",X"00",X"00",X"00",
		X"00",X"00",X"00",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",
		X"00",X"00",X"00",X"08",X"10",X"00",X"00",X"00",X"00",X"20",X"00",X"12",X"00",X"00",X"00",X"00",
		X"00",X"80",X"C0",X"E0",X"E0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"FC",X"FF",X"FF",X"E1",X"E0",X"E0",X"E0",X"00",X"00",X"00",X"C0",X"F8",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"E0",X"C0",X"00",X"F0",X"FE",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"E0",X"C0",X"00",X"F0",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"38",X"F8",X"F0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"E0",X"C0",X"01",X"FF",X"FF",X"FF",X"E0",X"18",X"38",X"70",X"F0",X"E0",X"C0",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"81",X"C3",X"E7",X"00",X"00",X"00",X"60",X"F0",X"E0",X"C0",X"80",
		X"EF",X"FE",X"FC",X"F8",X"F0",X"E0",X"E0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"80",X"C0",X"E0",X"E0",X"E0",X"C0",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"FF",X"E7",X"EE",X"EC",X"E0",X"E0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"E0",X"C0",X"00",X"E0",X"F8",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"E0",X"C0",X"0E",X"E7",X"FB",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E7",X"E3",X"C7",X"1F",X"FE",X"FC",X"F0",X"E0",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0C",X"0E",X"8E",X"C6",X"E7",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EF",X"EE",X"DC",X"3C",X"F8",X"F0",X"E0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"E0",X"E0",X"F0",X"F0",X"78",X"3C",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"00",X"00",X"00",X"00",
		X"E0",X"E0",X"E0",X"F0",X"F0",X"70",X"78",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3C",X"1C",X"1C",X"0E",X"0E",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"E0",X"F8",X"FC",X"FE",X"3E",X"1F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"0E",X"1C",X"1C",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"E0",X"F8",X"FC",X"FE",X"3E",X"0F",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"1C",X"38",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"FF",X"FF",X"FF",X"FF",X"07",X"0E",X"1C",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",
		X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E3",X"FF",X"FF",X"FF",X"FB",X"E1",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"C0",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"FB",X"FD",X"FD",
		X"FF",X"FE",X"FC",X"FC",X"F8",X"F8",X"D8",X"8C",X"9F",X"07",X"03",X"79",X"84",X"82",X"81",X"81",
		X"8E",X"AF",X"AC",X"98",X"C8",X"FC",X"FC",X"FE",X"41",X"22",X"3C",X"7E",X"7F",X"3F",X"1E",X"20",
		X"FA",X"FD",X"FE",X"FF",X"FF",X"FF",X"FE",X"FC",X"40",X"78",X"8E",X"63",X"90",X"CC",X"03",X"00",
		X"F8",X"F8",X"F8",X"F8",X"FC",X"FC",X"FC",X"FE",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"01",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"83",X"E7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"1F",X"17",X"2B",X"55",X"2B",X"43",X"33",X"19",X"F0",X"F8",X"FC",X"FE",X"FE",X"FE",X"FF",X"FF",
		X"F8",X"7E",X"FF",X"7F",X"FF",X"7F",X"03",X"00",X"7F",X"3E",X"3E",X"FC",X"FC",X"F8",X"F0",X"E0",
		X"1F",X"17",X"2B",X"55",X"2B",X"55",X"07",X"00",X"F8",X"FE",X"FF",X"FF",X"FF",X"E7",X"03",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"0F",X"3F",X"7F",X"5F",X"15",X"15",X"04",
		X"1F",X"1F",X"37",X"5B",X"2D",X"57",X"07",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"E0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",
		X"0C",X"00",X"00",X"00",X"06",X"06",X"00",X"00",X"30",X"00",X"00",X"00",X"60",X"60",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",
		X"06",X"00",X"00",X"0C",X"0E",X"0E",X"00",X"00",X"0C",X"00",X"00",X"30",X"70",X"70",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"EF",X"DF",X"BF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F9",X"E0",X"C0",X"9E",X"21",X"41",X"81",X"81",X"FF",X"7F",X"3F",X"3F",X"1F",X"1F",X"1B",X"31",
		X"82",X"44",X"3C",X"7E",X"FE",X"FC",X"78",X"04",X"71",X"F5",X"35",X"19",X"13",X"3F",X"3F",X"7F",
		X"02",X"1E",X"71",X"C6",X"09",X"33",X"C0",X"00",X"5F",X"BF",X"7F",X"FF",X"FF",X"FF",X"7F",X"3F",
		X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"80",X"1F",X"1F",X"1F",X"1F",X"3F",X"3F",X"3F",X"7F",
		X"C1",X"E7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"C0",X"E0",X"E0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"FC",X"FF",X"FF",X"FF",X"0F",X"00",X"00",X"78",X"F8",X"FE",X"FF",X"FF",X"FE",X"7C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"00",X"00",X"00",X"00",X"06",X"06",X"00",X"00",
		X"00",X"00",X"00",X"00",X"06",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"60",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",
		X"06",X"00",X"00",X"00",X"06",X"06",X"00",X"00",X"60",X"00",X"00",X"00",X"60",X"60",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"AA",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"AA",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"18",X"18",X"18",X"18",X"3C",X"18",X"18",X"18",
		X"FF",X"80",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"80",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",
		X"FF",X"18",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"FF",X"01",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",
		X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",
		X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"18",X"FF",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"01",X"FF",
		X"81",X"81",X"81",X"81",X"81",X"81",X"E1",X"E1",X"81",X"81",X"81",X"81",X"81",X"81",X"B1",X"B1",
		X"81",X"81",X"81",X"81",X"E1",X"E1",X"81",X"81",X"81",X"81",X"81",X"81",X"B1",X"B1",X"81",X"81",
		X"81",X"81",X"E1",X"E1",X"81",X"81",X"81",X"81",X"81",X"81",X"B1",X"B1",X"81",X"81",X"81",X"81",
		X"E1",X"E1",X"81",X"81",X"81",X"81",X"81",X"81",X"B1",X"B1",X"81",X"81",X"81",X"81",X"81",X"81",
		X"42",X"42",X"42",X"42",X"42",X"42",X"72",X"72",X"42",X"42",X"42",X"42",X"42",X"42",X"5A",X"5A",
		X"42",X"42",X"42",X"42",X"72",X"72",X"42",X"42",X"42",X"42",X"42",X"42",X"5A",X"5A",X"42",X"42",
		X"42",X"42",X"72",X"72",X"42",X"42",X"42",X"42",X"42",X"42",X"5A",X"5A",X"42",X"42",X"42",X"42",
		X"72",X"72",X"42",X"42",X"42",X"42",X"42",X"42",X"5A",X"5A",X"42",X"42",X"42",X"42",X"42",X"42",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"24",X"24",X"24",X"24",X"24",X"24",X"3C",X"3C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"24",X"24",X"24",X"24",X"3C",X"3C",X"24",X"24",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"24",X"24",X"3C",X"3C",X"24",X"24",X"24",X"24",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"3C",X"24",X"24",X"24",X"24",X"24",X"24",
		X"99",X"99",X"99",X"99",X"99",X"99",X"F9",X"F9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"99",X"99",X"99",X"F9",X"F9",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"99",X"F9",X"F9",X"99",X"99",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F9",X"F9",X"99",X"99",X"99",X"99",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"02",X"03",X"02",X"03",X"03",X"03",X"00",X"C0",X"C0",X"40",X"C0",X"E0",X"E0",X"E0",X"00",
		X"01",X"06",X"08",X"10",X"20",X"00",X"01",X"00",X"80",X"60",X"10",X"08",X"04",X"00",X"B8",X"00",
		X"1F",X"1F",X"1F",X"0F",X"0F",X"0F",X"03",X"00",X"F8",X"F8",X"F8",X"F0",X"F0",X"F0",X"C0",X"00",
		X"02",X"03",X"03",X"01",X"00",X"00",X"00",X"06",X"40",X"C0",X"C0",X"80",X"00",X"00",X"00",X"60",
		X"0D",X"0D",X"0F",X"07",X"05",X"07",X"03",X"00",X"B0",X"B0",X"F0",X"E0",X"A0",X"E0",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"0F",X"0E",X"11",X"21",X"22",X"9C",X"E0",X"F0",X"F0",
		X"0B",X"0C",X"0D",X"0A",X"08",X"08",X"06",X"01",X"D0",X"10",X"50",X"90",X"10",X"10",X"60",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"0F",X"1D",X"00",X"00",X"AA",X"00",X"00",X"00",X"E0",X"70",X"00",X"00",X"AA",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"0F",X"1F",X"3D",X"00",X"00",X"00",X"00",X"80",X"E0",X"F0",X"78",
		X"3F",X"1F",X"00",X"00",X"AA",X"00",X"00",X"00",X"F8",X"F0",X"00",X"00",X"AA",X"00",X"00",X"00",
		X"00",X"03",X"0F",X"1F",X"3D",X"3E",X"1F",X"1F",X"00",X"80",X"E0",X"F0",X"78",X"F8",X"F0",X"F0",
		X"0F",X"03",X"00",X"00",X"AA",X"00",X"00",X"00",X"E0",X"80",X"00",X"00",X"AA",X"00",X"00",X"00",
		X"0F",X"1B",X"3F",X"3F",X"1F",X"1F",X"0F",X"03",X"E0",X"70",X"F8",X"F8",X"F0",X"F0",X"E0",X"80",
		X"1F",X"7F",X"FF",X"7F",X"BF",X"00",X"00",X"00",X"F0",X"FC",X"FE",X"FC",X"FA",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"0F",X"3C",X"F0",X"03",X"0F",X"3C",X"F0",X"C0",X"00",X"03",X"0F",
		X"C0",X"00",X"03",X"0F",X"3C",X"F0",X"C0",X"00",X"3C",X"F0",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"03",X"03",X"06",X"06",X"0C",X"0C",X"86",X"86",X"0C",X"0C",X"18",X"18",X"30",X"30",
		X"18",X"18",X"30",X"30",X"61",X"61",X"C3",X"C3",X"60",X"60",X"C0",X"C0",X"80",X"80",X"00",X"00",
		X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",
		X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"84",X"87",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"E0",
		X"C7",X"E4",X"78",X"30",X"00",X"00",X"00",X"00",X"F0",X"38",X"1E",X"0C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"20",X"E0",X"F0",
		X"07",X"84",X"84",X"C0",X"78",X"30",X"00",X"00",X"1E",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"80",X"C0",X"F0",X"F0",
		X"01",X"07",X"03",X"41",X"60",X"70",X"3E",X"1C",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"08",X"0C",X"07",X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"20",X"C0",X"80",X"80",
		X"01",X"01",X"00",X"00",X"08",X"0C",X"07",X"03",X"80",X"80",X"00",X"00",X"00",X"00",X"60",X"C0",
		X"F0",X"F8",X"FC",X"FE",X"FF",X"FF",X"FF",X"F7",X"0F",X"0F",X"0F",X"0F",X"0F",X"8F",X"CF",X"EF",
		X"F3",X"F1",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"FF",X"FF",X"FF",X"7F",X"3F",X"1F",X"0F",X"0F",
		X"39",X"39",X"39",X"01",X"01",X"39",X"39",X"39",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"CC",X"DE",
		X"39",X"39",X"39",X"39",X"39",X"39",X"39",X"39",X"FF",X"CF",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C7",
		X"1D",X"38",X"38",X"38",X"38",X"1D",X"1F",X"07",X"C7",X"E7",X"E7",X"E7",X"E7",X"C7",X"C7",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"78",X"FC",X"3C",X"1C",X"1C",X"1C",X"1C",X"1C",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"FE",X"FF",X"07",X"03",X"03",X"03",X"07",X"FF",X"00",X"00",X"80",X"C0",X"C0",X"C0",X"8E",X"0E",
		X"FF",X"07",X"03",X"03",X"03",X"07",X"FF",X"FE",X"0E",X"8E",X"CE",X"CE",X"CF",X"8F",X"07",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"39",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"FE",
		X"39",X"39",X"38",X"38",X"38",X"F9",X"B9",X"38",X"86",X"C0",X"F8",X"7C",X"0E",X"86",X"FE",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"8F",
		X"61",X"70",X"3E",X"1F",X"03",X"61",X"7F",X"3F",X"9D",X"18",X"00",X"0F",X"98",X"98",X"9F",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"87",X"C7",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"78",
		X"C7",X"E7",X"E7",X"E7",X"E7",X"E7",X"E7",X"E7",X"FC",X"3C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",
		X"07",X"1F",X"3F",X"7C",X"78",X"F0",X"F0",X"F0",X"C0",X"E0",X"F0",X"78",X"38",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"78",X"7C",X"3F",X"1F",X"07",X"00",X"01",X"01",X"39",X"79",X"F0",X"E0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"C7",X"C7",X"C7",X"C7",X"EE",X"FE",X"38",X"00",X"00",X"00",X"00",X"66",X"66",X"02",X"04",
		X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"00",X"38",X"38",X"38",X"38",X"FE",X"FE",X"38",
		X"70",X"70",X"70",X"70",X"70",X"7F",X"7F",X"7F",X"38",X"38",X"38",X"38",X"38",X"38",X"1E",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"3E",X"7F",X"F1",X"E0",X"F1",X"7F",X"3E",X"0C",X"E0",X"E0",X"E0",X"E0",X"E3",X"E3",X"E0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"42",X"42",X"42",X"42",X"42",X"42",X"42",X"42",X"42",X"42",X"42",X"42",X"42",X"42",X"42",X"42",
		X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"24",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
