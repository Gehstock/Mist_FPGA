library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity travusa_chr_bit1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of travusa_chr_bit1 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",
		X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"10",X"08",X"08",X"10",X"10",X"20",X"20",X"10",X"10",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"30",X"30",X"30",X"30",X"30",
		X"30",X"30",X"30",X"30",X"38",X"30",X"20",X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"00",
		X"00",X"00",X"00",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"48",X"FC",X"48",X"24",X"7E",X"24",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"44",X"82",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"82",X"44",X"38",X"00",X"80",X"40",X"20",X"10",X"08",X"04",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"16",X"0E",X"00",X"00",X"00",
		X"00",X"00",X"16",X"0E",X"00",X"00",X"16",X"0E",X"00",X"F8",X"FC",X"26",X"22",X"26",X"FC",X"F8",
		X"00",X"FE",X"FE",X"92",X"92",X"92",X"FE",X"6C",X"00",X"38",X"7C",X"C6",X"82",X"82",X"C6",X"44",
		X"00",X"FE",X"FE",X"82",X"82",X"C6",X"7C",X"38",X"00",X"FE",X"FE",X"92",X"92",X"92",X"82",X"80",
		X"00",X"FE",X"FE",X"12",X"12",X"12",X"12",X"02",X"00",X"38",X"7C",X"C6",X"82",X"92",X"F2",X"F2",
		X"00",X"FE",X"FE",X"10",X"10",X"10",X"FE",X"FE",X"00",X"82",X"82",X"FE",X"FE",X"82",X"82",X"00",
		X"00",X"40",X"C0",X"80",X"80",X"80",X"7E",X"7E",X"00",X"FE",X"FE",X"30",X"78",X"EC",X"C6",X"82",
		X"00",X"FE",X"FE",X"80",X"80",X"80",X"80",X"80",X"00",X"FE",X"FE",X"1C",X"38",X"1C",X"FE",X"FE",
		X"00",X"FE",X"FE",X"1C",X"38",X"70",X"FE",X"FE",X"00",X"7C",X"FE",X"82",X"82",X"82",X"FE",X"7C",
		X"00",X"FE",X"FE",X"22",X"22",X"22",X"3E",X"1C",X"00",X"7C",X"FE",X"82",X"A2",X"C2",X"7E",X"FC",
		X"00",X"FE",X"FE",X"22",X"62",X"F2",X"DE",X"9C",X"00",X"4C",X"DE",X"92",X"92",X"96",X"F4",X"60",
		X"00",X"02",X"02",X"FE",X"FE",X"02",X"02",X"00",X"00",X"7E",X"FE",X"80",X"80",X"80",X"FE",X"7E",
		X"00",X"1E",X"3E",X"70",X"E0",X"70",X"3E",X"1E",X"00",X"FE",X"FE",X"70",X"38",X"70",X"FE",X"FE",
		X"00",X"C6",X"EE",X"7C",X"38",X"7C",X"EE",X"C6",X"00",X"0E",X"1E",X"F0",X"F0",X"1E",X"0E",X"00",
		X"00",X"C6",X"E6",X"F6",X"DE",X"CE",X"C6",X"00",X"00",X"1E",X"04",X"1A",X"00",X"1C",X"04",X"18",
		X"84",X"58",X"20",X"10",X"08",X"F4",X"22",X"C0",X"3C",X"42",X"99",X"A5",X"A5",X"91",X"42",X"3C",
		X"00",X"1E",X"04",X"08",X"04",X"1E",X"00",X"90",X"40",X"20",X"10",X"08",X"04",X"F2",X"20",X"C0",
		X"F8",X"80",X"80",X"00",X"80",X"00",X"F0",X"48",X"48",X"F0",X"00",X"80",X"00",X"00",X"00",X"00",
		X"F8",X"80",X"80",X"00",X"80",X"00",X"38",X"40",X"80",X"40",X"38",X"80",X"00",X"00",X"00",X"00",
		X"F8",X"20",X"20",X"F8",X"00",X"70",X"88",X"88",X"70",X"00",X"78",X"80",X"80",X"78",X"00",X"80",
		X"90",X"A8",X"A8",X"40",X"00",X"08",X"F8",X"08",X"80",X"00",X"00",X"F8",X"80",X"80",X"00",X"80",
		X"70",X"88",X"88",X"00",X"F8",X"20",X"20",X"F8",X"00",X"F8",X"00",X"80",X"00",X"00",X"00",X"00",
		X"1F",X"02",X"04",X"1F",X"00",X"10",X"03",X"04",X"1C",X"04",X"13",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"C0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"EA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"38",X"7C",X"C2",X"82",X"86",X"7C",X"38",X"00",X"80",X"84",X"FE",X"FE",X"80",X"80",X"00",
		X"00",X"CC",X"E6",X"F2",X"B2",X"BA",X"9E",X"8C",X"00",X"40",X"C2",X"92",X"9A",X"9E",X"F6",X"62",
		X"00",X"30",X"38",X"2C",X"26",X"FE",X"FE",X"20",X"00",X"4E",X"CE",X"8A",X"8A",X"FA",X"70",X"00",
		X"00",X"78",X"FC",X"96",X"92",X"92",X"F2",X"60",X"00",X"06",X"06",X"E2",X"F2",X"1A",X"0E",X"06",
		X"00",X"6C",X"9E",X"9A",X"B2",X"B2",X"EC",X"60",X"00",X"0C",X"9E",X"92",X"92",X"D2",X"7E",X"3C",
		X"00",X"40",X"C0",X"80",X"80",X"80",X"FE",X"7E",X"00",X"7E",X"FE",X"80",X"80",X"80",X"FE",X"7E",
		X"00",X"FE",X"FE",X"1C",X"38",X"1C",X"FE",X"FE",X"00",X"FE",X"FE",X"22",X"22",X"22",X"3E",X"1C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"20",X"20",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"E3",X"C1",X"C1",X"C1",X"C3",X"E3",X"E7",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"3F",X"1F",X"0F",X"07",X"47",X"E3",X"73",X"E3",X"E3",X"B3",
		X"F7",X"E7",X"4F",X"1F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"F3",X"E0",X"E0",X"E2",X"C2",
		X"C7",X"C3",X"CB",X"CF",X"CF",X"E5",X"E5",X"E5",X"E1",X"E0",X"F0",X"F8",X"FC",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"73",X"34",X"37",X"43",X"81",X"80",X"00",X"00",X"FF",X"FE",X"FC",X"FC",X"FC",X"FC",X"FE",X"FE",
		X"FF",X"3F",X"3F",X"43",X"81",X"80",X"00",X"00",X"FF",X"FE",X"FC",X"FC",X"FC",X"FC",X"FE",X"FE",
		X"0F",X"03",X"01",X"00",X"00",X"80",X"A1",X"BF",X"FC",X"FC",X"FC",X"FC",X"FE",X"FF",X"FF",X"FF",
		X"0F",X"03",X"01",X"00",X"00",X"80",X"E1",X"FF",X"FC",X"FC",X"FC",X"FC",X"FE",X"FF",X"FF",X"FF",
		X"DC",X"DC",X"9C",X"DC",X"DE",X"DF",X"1F",X"BF",X"06",X"20",X"20",X"20",X"00",X"00",X"00",X"00",
		X"0E",X"17",X"1F",X"1E",X"1F",X"0F",X"0F",X"07",X"07",X"05",X"03",X"03",X"03",X"03",X"03",X"03",
		X"03",X"03",X"03",X"03",X"07",X"07",X"06",X"0E",X"0C",X"15",X"1D",X"19",X"1B",X"1B",X"1B",X"2B",
		X"3B",X"3B",X"3B",X"19",X"1D",X"1C",X"1E",X"0E",X"0C",X"0E",X"0E",X"06",X"0E",X"0E",X"0E",X"0E",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"7F",X"3F",X"BF",X"BF",X"BF",X"9F",X"DF",X"DF",X"9F",X"DF",X"DF",X"DF",X"DF",X"1F",X"BF",
		X"BF",X"BF",X"3F",X"7F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F3",X"F4",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",X"F2",X"F9",X"FC",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"FC",X"FD",X"FD",X"FD",X"F9",X"FA",X"FB",X"FB",X"73",X"F4",X"E7",X"EF",X"CF",X"DF",X"9B",X"8D",
		X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"BE",X"AF",X"9F",X"DF",X"DF",X"CB",X"ED",X"EF",X"EF",X"E7",
		X"F0",X"F0",X"F0",X"F0",X"C0",X"F0",X"F0",X"70",X"F0",X"F8",X"F8",X"E8",X"D8",X"FC",X"FC",X"7C",
		X"B4",X"F8",X"F8",X"F8",X"F8",X"F8",X"E8",X"F0",X"F0",X"F0",X"E0",X"E0",X"C0",X"C0",X"C0",X"80",
		X"80",X"80",X"80",X"80",X"80",X"40",X"C0",X"C0",X"C0",X"C0",X"C0",X"A0",X"E0",X"E0",X"E0",X"F0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F0",X"F0",X"F8",X"FC",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",X"FD",X"F9",X"79",X"1D",X"3D",X"2F",
		X"DF",X"9E",X"DC",X"DC",X"DC",X"DC",X"1E",X"BE",X"FF",X"3F",X"3F",X"43",X"80",X"80",X"00",X"00",
		X"FC",X"FC",X"FC",X"FC",X"FE",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3D",X"1C",X"0C",X"06",X"06",X"06",X"0E",X"1A",X"BF",X"BE",X"3C",X"7C",X"7C",X"7C",X"7E",X"FE",
		X"FF",X"3F",X"3F",X"43",X"81",X"80",X"00",X"00",X"FC",X"FC",X"FC",X"FC",X"FE",X"FF",X"FF",X"FF",
		X"F0",X"90",X"D0",X"F0",X"10",X"F0",X"F0",X"F0",X"07",X"03",X"01",X"00",X"00",X"40",X"C1",X"C5",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FE",X"70",X"38",X"70",X"FE",X"FE",
		X"00",X"FE",X"FE",X"10",X"10",X"10",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"F8",X"E0",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",
		X"F0",X"F0",X"60",X"60",X"C0",X"80",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"6F",X"3F",X"1F",X"17",X"1F",X"3F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"F0",X"C0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"1F",X"03",X"00",X"80",X"C0",X"E0",X"00",X"00",X"00",X"00",X"80",X"C0",X"60",X"F0",
		X"FE",X"FF",X"FF",X"FF",X"7D",X"3F",X"3F",X"FF",X"0F",X"00",X"00",X"01",X"E1",X"03",X"C6",X"EC",
		X"F0",X"F0",X"E0",X"E0",X"C0",X"80",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FE",X"E7",X"E7",X"E3",X"E0",X"F0",X"F8",X"FC",X"FE",X"FF",X"FF",X"87",X"0F",
		X"1F",X"3F",X"03",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"FF",X"FF",X"7F",X"3F",X"1F",
		X"1F",X"74",X"F0",X"C1",X"E1",X"C3",X"8F",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F3",X"F1",X"E1",X"DF",X"FF",X"FF",X"FF",X"7F",X"FF",X"BF",X"FF",X"FF",X"FF",X"CF",X"83",X"80",
		X"00",X"40",X"60",X"F0",X"FC",X"FE",X"FC",X"FE",X"3F",X"03",X"01",X"A0",X"F8",X"38",X"58",X"DC",
		X"DE",X"CF",X"87",X"07",X"1F",X"FF",X"FF",X"FF",X"0F",X"0F",X"0F",X"1F",X"1F",X"1F",X"3F",X"3F",
		X"7F",X"1F",X"0F",X"07",X"03",X"03",X"01",X"00",X"00",X"00",X"01",X"01",X"01",X"03",X"03",X"07",
		X"0C",X"08",X"08",X"1E",X"1F",X"1F",X"30",X"21",X"00",X"FE",X"FE",X"92",X"92",X"92",X"82",X"80",
		X"00",X"FE",X"FE",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"82",X"FE",X"FE",X"82",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"3F",X"FC",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"FF",X"FF",X"FF",X"FF",X"E7",X"42",X"00",
		X"FF",X"FF",X"F8",X"00",X"00",X"00",X"00",X"00",X"FE",X"E0",X"00",X"00",X"00",X"00",X"01",X"07",
		X"F3",X"38",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"7F",X"FF",X"FF",
		X"04",X"03",X"FB",X"FF",X"FF",X"FB",X"FC",X"E0",X"FF",X"FF",X"FF",X"FF",X"F8",X"E0",X"20",X"20",
		X"80",X"00",X"00",X"03",X"07",X"0F",X"1F",X"1F",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"FF",X"FE",X"FC",X"E0",X"80",X"01",X"03",X"0F",X"1F",X"FF",X"FF",X"FF",X"FE",X"F8",X"F8",
		X"FC",X"E0",X"E0",X"80",X"80",X"00",X"00",X"00",X"F8",X"C8",X"08",X"0B",X"37",X"F7",X"F7",X"F7",
		X"00",X"00",X"3F",X"FF",X"FF",X"F2",X"C0",X"00",X"3F",X"FE",X"FC",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"FF",
		X"E0",X"00",X"00",X"00",X"1F",X"FF",X"FF",X"FF",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"3F",X"FC",X"E0",X"00",X"00",X"01",X"0F",X"7F",
		X"FF",X"FF",X"F8",X"C0",X"00",X"00",X"00",X"00",X"00",X"01",X"0F",X"3F",X"F8",X"E0",X"80",X"00",
		X"03",X"0F",X"3F",X"FF",X"FE",X"F8",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",X"03",X"0F",X"3E",
		X"F8",X"E0",X"80",X"00",X"03",X"0F",X"3F",X"FF",X"FE",X"F8",X"E0",X"80",X"00",X"00",X"00",X"00",
		X"00",X"03",X"0F",X"3E",X"F8",X"E0",X"80",X"00",X"0E",X"1F",X"3F",X"1F",X"3F",X"7F",X"6F",X"1F",
		X"00",X"03",X"1F",X"FE",X"F0",X"80",X"00",X"00",X"07",X"3F",X"FF",X"FF",X"FC",X"E0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"7F",X"FC",X"C0",X"00",X"00",X"01",X"1F",X"FF",X"FF",X"FF",X"F0",
		X"00",X"03",X"0F",X"7E",X"F8",X"C0",X"00",X"00",X"07",X"7F",X"FF",X"FF",X"FC",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"1F",X"FE",X"F0",X"80",X"00",X"00",X"07",X"3F",X"FF",X"FF",X"FC",
		X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",
		X"C0",X"00",X"00",X"00",X"1F",X"FF",X"FF",X"FF",X"70",X"38",X"B8",X"DC",X"FC",X"F8",X"FC",X"FC",
		X"00",X"01",X"1F",X"FF",X"F0",X"00",X"00",X"00",X"07",X"7F",X"FF",X"FF",X"FC",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"01",X"7F",X"FF",X"C0",X"00",X"00",X"00",X"1F",X"FF",X"FF",X"FF",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"1F",X"FF",X"F0",X"00",X"00",X"00",X"07",X"FF",X"FF",X"FF",X"FC",
		X"FF",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"FC",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",X"3F",X"FF",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"0F",X"1E",X"38",X"70",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"0E",X"0C",X"1C",X"18",X"18",X"18",
		X"18",X"18",X"18",X"18",X"18",X"1C",X"1F",X"0F",X"00",X"00",X"00",X"00",X"03",X"0F",X"3F",X"FF",
		X"FE",X"78",X"60",X"00",X"00",X"00",X"00",X"00",X"80",X"E0",X"FC",X"3E",X"07",X"03",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"E0",X"60",X"70",X"70",X"30",X"38",X"18",X"18",
		X"1C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"FF",
		X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"3F",X"3D",X"18",X"01",X"0F",X"06",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FF",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"FF",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"80",X"F8",X"FF",X"0F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"F8",X"7F",X"0F",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"F8",X"3E",
		X"C0",X"E0",X"70",X"38",X"1C",X"0E",X"07",X"1E",X"C0",X"E0",X"70",X"38",X"1C",X"0E",X"FF",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"F0",X"7C",X"1F",X"07",X"00",X"00",X"00",X"00",
		X"00",X"80",X"FF",X"FF",X"00",X"00",X"00",X"00",X"07",X"00",X"03",X"0F",X"7E",X"F8",X"C0",X"00",
		X"0F",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"E0",X"F8",X"3E",X"0F",X"03",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"E0",X"F0",X"3C",X"1E",X"07",X"03",X"00",X"00",X"00",X"00",X"00",
		X"00",X"80",X"C0",X"F0",X"78",X"1E",X"0F",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",X"70",X"38",X"1C",X"0E",X"07",X"03",
		X"F4",X"70",X"40",X"E0",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",
		X"3E",X"FF",X"FF",X"FC",X"E0",X"00",X"00",X"00",X"00",X"01",X"0F",X"FF",X"FF",X"FF",X"F8",X"80",
		X"00",X"00",X"00",X"00",X"1F",X"FF",X"FF",X"FF",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"07",X"FF",X"FF",X"FF",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"1F",
		X"00",X"00",X"01",X"03",X"07",X"0F",X"1F",X"3E",X"7C",X"38",X"10",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"3F",X"FC",
		X"3F",X"1F",X"00",X"60",X"E0",X"C0",X"80",X"00",X"E0",X"F8",X"E0",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"3F",X"FE",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"3F",X"FE",X"E0",
		X"00",X"20",X"9C",X"83",X"A0",X"F8",X"FF",X"E1",X"80",X"FE",X"FF",X"FF",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"E0",X"E0",X"E0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"0F",X"3E",
		X"00",X"00",X"00",X"C1",X"33",X"03",X"01",X"20",X"0F",X"7F",X"F8",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"3F",X"FE",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"3F",X"FE",X"E0",X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"F0",X"F0",X"F8",X"F8",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"0F",X"7F",X"FF",X"FF",X"F8",X"C0",X"00",X"00",
		X"40",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"FE",X"E0",X"07",X"3F",X"FF",X"FF",X"FC",X"E0",
		X"03",X"3F",X"FE",X"E0",X"03",X"1F",X"FF",X"FF",X"FE",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"3F",X"FE",X"E0",X"01",X"0F",X"FF",X"FF",X"FF",X"F8",X"80",X"00",X"00",X"00",
		X"70",X"70",X"FC",X"FC",X"FF",X"7F",X"7F",X"07",X"00",X"07",X"7F",X"FF",X"FF",X"FC",X"C0",X"00",
		X"00",X"00",X"00",X"03",X"FF",X"FF",X"FF",X"FE",X"00",X"00",X"00",X"00",X"00",X"01",X"0F",X"7F",
		X"78",X"78",X"78",X"7B",X"33",X"A7",X"AF",X"FC",X"00",X"00",X"00",X"07",X"3F",X"FF",X"FF",X"FC",
		X"FF",X"FE",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"3F",X"FF",X"7F",X"7C",
		X"20",X"F0",X"F0",X"F8",X"F8",X"E0",X"80",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",
		X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7C",X"F8",X"F0",X"E0",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"01",X"E3",X"83",X"87",X"C7",X"5E",X"1E",X"7C",
		X"B0",X"D8",X"D8",X"5E",X"4E",X"6F",X"EF",X"E7",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"E0",
		X"CF",X"FF",X"F8",X"00",X"00",X"00",X"07",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FD",X"F9",X"7B",X"31",X"10",X"00",X"00",X"00",X"F7",X"F7",X"F7",X"F7",X"F0",X"60",X"20",X"00",
		X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"02",X"22",X"12",
		X"39",X"7F",X"7F",X"FF",X"FE",X"FE",X"FD",X"FF",X"C0",X"80",X"1E",X"7E",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"30",X"78",X"7C",X"FC",X"41",X"E9",X"27",X"33",X"FD",X"7B",X"3B",X"7B",
		X"FB",X"F1",X"FB",X"F3",X"FB",X"FF",X"FD",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"FC",X"FE",X"FF",X"FF",X"FF",X"FE",X"F4",X"F8",
		X"E9",X"1C",X"12",X"04",X"05",X"03",X"03",X"01",X"FE",X"7C",X"FF",X"79",X"33",X"C7",X"FF",X"FD",
		X"EF",X"5F",X"1F",X"BF",X"FF",X"ED",X"C0",X"F1",X"FE",X"EF",X"DF",X"3E",X"EC",X"B0",X"7C",X"E8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B8",X"04",X"71",X"39",X"10",X"00",X"00",X"00",
		X"E0",X"48",X"1C",X"F7",X"F8",X"6E",X"00",X"00",X"C0",X"00",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"07",X"3F",X"FF",X"FF",X"FC",X"E0",X"00",X"39",X"FF",X"FF",X"E0",X"00",X"00",X"00",
		X"FF",X"FF",X"FC",X"F0",X"80",X"00",X"00",X"00",X"01",X"01",X"03",X"1F",X"7F",X"FF",X"FF",X"FF",
		X"80",X"00",X"01",X"07",X"3F",X"FF",X"FF",X"FC",X"43",X"DF",X"BF",X"BF",X"BC",X"80",X"C0",X"41",
		X"00",X"00",X"00",X"00",X"11",X"1F",X"1F",X"7F",X"F8",X"E0",X"C0",X"00",X"01",X"0F",X"7F",X"FF",
		X"FF",X"F8",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"7F",X"FF",X"FF",X"C0",X"00",
		X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"FE",X"FE",X"22",X"62",X"F2",X"DE",X"9C",X"00",X"70",X"F8",X"A8",X"A8",X"B8",X"B0",X"00",
		X"08",X"7C",X"FC",X"88",X"C8",X"40",X"00",X"F6",X"F6",X"00",X"00",X"F8",X"F8",X"20",X"38",X"18",
		X"00",X"70",X"F8",X"A8",X"A8",X"B8",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"7F",X"FF",X"C0",
		X"00",X"00",X"01",X"1F",X"FF",X"F0",X"00",X"00",X"0F",X"3E",X"F8",X"E0",X"00",X"00",X"00",X"00",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"00",X"00",X"00",X"03",X"0F",X"3E",X"F8",X"E0",X"0F",X"3E",X"F8",X"E0",X"80",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"3F",X"07",X"3F",X"FC",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"3F",X"00",X"00",X"00",X"00",X"03",X"3F",X"FF",X"FF",
		X"0F",X"1F",X"3E",X"FC",X"F8",X"F0",X"E0",X"80",X"E0",X"C0",X"C0",X"40",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"0F",X"07",X"03",X"07",X"08",X"38",X"F8",X"F0",X"F0",X"F0",X"E0",X"E0",
		X"FE",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"1F",X"3E",X"FC",X"F8",X"F0",X"FF",X"FF",
		X"E0",X"C0",X"C0",X"42",X"03",X"03",X"FF",X"FF",X"00",X"00",X"00",X"00",X"80",X"E0",X"F8",X"FE",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"03",X"03",X"02",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"FF",X"FF",X"FF",X"F8",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",
		X"7F",X"7F",X"7F",X"3F",X"3F",X"3F",X"3F",X"1F",X"1F",X"1F",X"1F",X"0F",X"0F",X"0F",X"0F",X"07",
		X"F0",X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",X"FC",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"F9",X"F3",X"67",X"6F",X"7F",X"3F",X"3E",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"04",X"07",X"FC",X"FC",X"FC",X"FC",X"FE",X"FE",X"FE",X"FE",
		X"FF",X"FF",X"FC",X"80",X"00",X"00",X"00",X"00",X"3C",X"FC",X"FF",X"FF",X"FF",X"FF",X"07",X"03",
		X"00",X"C2",X"E7",X"FF",X"FF",X"FF",X"FF",X"FF",X"40",X"70",X"F9",X"FF",X"FF",X"FF",X"CF",X"03",
		X"40",X"70",X"F1",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"01",X"01",X"03",X"1F",X"3F",X"3F",X"3F",X"3F",
		X"03",X"9F",X"FF",X"FF",X"FC",X"C0",X"C0",X"C1",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"1F",
		X"CF",X"FF",X"FF",X"FF",X"F8",X"E0",X"E0",X"E0",X"1F",X"1F",X"1F",X"0F",X"0F",X"0F",X"0F",X"07",
		X"F0",X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",X"07",X"07",X"07",X"03",X"03",X"03",X"03",X"01",
		X"FC",X"FC",X"FC",X"FC",X"FE",X"FE",X"FE",X"FE",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",
		X"7F",X"7F",X"7F",X"3F",X"3F",X"3F",X"3F",X"1F",X"C0",X"C0",X"C0",X"C0",X"E0",X"E0",X"E0",X"E0",
		X"1F",X"1F",X"1F",X"0F",X"0F",X"0F",X"0F",X"07",X"F0",X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",
		X"07",X"07",X"07",X"03",X"03",X"03",X"03",X"01",X"80",X"00",X"00",X"00",X"00",X"3F",X"FF",X"FF",
		X"C1",X"E7",X"FF",X"FF",X"FF",X"FE",X"F0",X"00",X"00",X"00",X"01",X"7F",X"FF",X"FF",X"FF",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"3F",X"FF",X"FF",X"FF",X"FF",X"80",X"00",X"00",X"00",
		X"00",X"0F",X"FF",X"FF",X"FF",X"F8",X"00",X"00",X"00",X"00",X"01",X"0F",X"0F",X"7F",X"7F",X"FF",
		X"FE",X"FC",X"F8",X"00",X"00",X"00",X"03",X"1F",X"FF",X"FF",X"FE",X"F0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"0F",X"8F",X"FF",X"FF",X"FF",X"FE",X"F0",X"00",
		X"00",X"00",X"01",X"07",X"3F",X"FF",X"FF",X"FC",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"9F",X"FF",X"FF",X"FF",X"FF",X"80",X"00",X"00",X"01",
		X"0F",X"3F",X"FF",X"FF",X"F8",X"E0",X"00",X"00",X"00",X"01",X"01",X"03",X"0F",X"3F",X"FF",X"FF",
		X"FE",X"FC",X"F8",X"00",X"03",X"0F",X"7F",X"FF",X"FE",X"F8",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"03",X"0D",X"3F",X"FF",X"FF",X"FE",X"F0",X"80",X"00",X"03",X"1F",X"7F",X"FF",X"FE",X"F0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"13",X"3F",X"FF",X"FF",X"FE",X"F8",X"E0",X"80",X"00",X"07",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"55",X"FF",X"55",X"FF",X"55",X"FF",X"FF",
		X"FF",X"55",X"FF",X"55",X"FF",X"55",X"FF",X"FF",X"FC",X"4E",X"FF",X"4B",X"FF",X"4F",X"FF",X"FF",
		X"00",X"00",X"00",X"80",X"F8",X"80",X"80",X"00",X"FF",X"FD",X"FF",X"55",X"FF",X"55",X"FF",X"FF",
		X"FF",X"FD",X"FF",X"F5",X"FF",X"F5",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"E0",X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"B9",X"FF",X"B9",X"FF",X"B9",X"FF",X"B9",X"B9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"38",X"7C",X"FC",X"FC",X"7C",X"7C",X"38",X"FF",X"FF",X"FF",X"7F",X"7F",X"00",X"68",X"04",
		X"FE",X"FF",X"FE",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FE",X"FD",X"F8",X"F5",X"FF",X"55",
		X"78",X"DB",X"00",X"5B",X"00",X"5B",X"00",X"00",X"20",X"40",X"2E",X"40",X"2E",X"40",X"3E",X"9F",
		X"00",X"00",X"00",X"00",X"00",X"60",X"C0",X"80",X"6B",X"07",X"7F",X"7C",X"F8",X"80",X"80",X"00",
		X"E0",X"E0",X"E0",X"00",X"00",X"00",X"00",X"00",X"FF",X"4D",X"FC",X"4A",X"FE",X"4C",X"FC",X"4A",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"FE",X"4C",X"FC",X"4A",X"FE",X"4C",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"4D",X"FC",X"4A",X"FE",X"4C",X"FF",X"FF",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"00",X"FF",X"FF",X"55",X"FF",X"FF",X"55",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"24",X"FF",X"24",X"FF",X"24",X"FF",X"FF",
		X"FF",X"92",X"FF",X"92",X"FF",X"92",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"BE",X"BF",X"FB",X"FF",
		X"FE",X"FE",X"DE",X"F6",X"FE",X"DC",X"00",X"00",X"00",X"00",X"00",X"F6",X"BE",X"EA",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FA",X"BE",X"F6",X"00",X"00",X"00",X"00",X"00",X"00",X"78",X"00",
		X"F8",X"F8",X"E0",X"E0",X"E0",X"E0",X"E0",X"F8",X"00",X"FE",X"F6",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FE",X"FE",X"00",X"00",X"00",X"00",X"00",X"D6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"4F",X"FF",X"4B",X"FF",X"4F",X"FF",X"FF",
		X"FC",X"4C",X"FC",X"48",X"FE",X"4C",X"FF",X"FF",X"FE",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"FE",X"FC",X"F0",X"F0",X"E0",X"E0",X"C0",X"FF",X"FF",X"4D",X"FC",X"4A",X"FE",X"4C",X"FC",X"48",
		X"B8",X"78",X"37",X"F0",X"00",X"00",X"00",X"00",X"FE",X"4C",X"FC",X"4A",X"FE",X"4C",X"FF",X"FF",
		X"FF",X"FC",X"FF",X"24",X"FF",X"24",X"FF",X"FF",X"FE",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FC",X"FF",X"F4",X"FF",X"E4",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"60",X"C0",X"80",
		X"FF",X"FF",X"FF",X"55",X"FF",X"55",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"0F",X"F1",X"FF",X"82",X"7C",X"B9",X"D7",X"FF",X"FF",X"01",X"FF",X"FE",X"45",X"B9",X"D7",
		X"55",X"FF",X"FF",X"01",X"FE",X"45",X"B9",X"D7",X"00",X"00",X"F0",X"0F",X"F2",X"7D",X"2A",X"D7",
		X"00",X"00",X"00",X"F0",X"38",X"FF",X"B8",X"F8",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"FF",X"FF",X"03",X"05",X"0E",X"0F",X"00",X"00",X"2D",X"D5",X"BB",X"01",X"FF",X"F0",X"00",X"00",
		X"29",X"D5",X"BB",X"01",X"FF",X"00",X"00",X"00",X"29",X"D5",X"BB",X"01",X"FF",X"00",X"00",X"00",
		X"2A",X"D7",X"82",X"7F",X"F0",X"00",X"00",X"00",X"03",X"B7",X"03",X"B5",X"03",X"B7",X"03",X"FF",
		X"FE",X"FF",X"00",X"DB",X"00",X"DB",X"00",X"FF",X"00",X"B6",X"03",X"B5",X"03",X"B7",X"03",X"FF",
		X"FF",X"4F",X"FF",X"49",X"FF",X"4F",X"FF",X"49",X"FF",X"92",X"FF",X"92",X"FF",X"92",X"FF",X"FF",
		X"FC",X"4C",X"FC",X"4A",X"FC",X"4C",X"FF",X"FF",X"FF",X"4F",X"FF",X"4B",X"FF",X"4F",X"FF",X"FF",
		X"FE",X"FF",X"F0",X"FB",X"E0",X"EB",X"C0",X"FF",X"00",X"6D",X"00",X"6D",X"00",X"6D",X"00",X"FF",
		X"FF",X"FF",X"00",X"AA",X"00",X"AA",X"00",X"FF",X"FF",X"FC",X"FF",X"F4",X"FF",X"E4",X"FF",X"FF",
		X"FF",X"24",X"FF",X"24",X"FF",X"24",X"FF",X"FF",X"00",X"00",X"80",X"F0",X"FF",X"F0",X"80",X"00",
		X"00",X"00",X"00",X"10",X"1F",X"F0",X"80",X"00",X"FE",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"DB",X"00",X"DB",X"00",X"DB",X"00",X"FF",X"FF",X"FC",X"FF",X"24",X"FF",X"24",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"55",X"FF",X"FF",X"55",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"04",X"06",X"07",X"17",X"07",X"07",X"FE",X"FC",X"00",X"00",X"8F",X"FF",X"FF",X"FF",
		X"00",X"00",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"04",X"8F",X"FF",X"FF",X"FD",X"FD",X"FF",
		X"07",X"FF",X"FF",X"E1",X"80",X"20",X"48",X"F0",X"E0",X"F8",X"F0",X"B8",X"10",X"00",X"00",X"00",
		X"07",X"47",X"D7",X"DC",X"7C",X"78",X"60",X"40",X"FF",X"FF",X"FF",X"7F",X"0F",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FB",X"03",X"01",X"00",X"FF",X"FF",X"F9",X"F1",X"E1",X"E0",X"F0",X"58",
		X"E0",X"F0",X"C8",X"40",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"09",X"04",X"05",X"05",X"05",X"05",X"01",
		X"00",X"80",X"83",X"01",X"04",X"04",X"48",X"48",X"00",X"1C",X"62",X"81",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"20",X"C0",X"80",X"40",X"50",X"00",X"C0",X"C0",X"00",X"C0",X"C5",X"05",X"C5",
		X"48",X"44",X"44",X"44",X"08",X"18",X"40",X"40",X"00",X"00",X"E0",X"40",X"E0",X"00",X"C0",X"60",
		X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"E0",X"80",X"00",X"E0",X"80",X"00",
		X"00",X"00",X"00",X"00",X"81",X"62",X"1C",X"00",X"00",X"00",X"03",X"07",X"07",X"0E",X"0C",X"0C",
		X"00",X"E0",X"F8",X"FE",X"0F",X"07",X"03",X"03",X"0E",X"0E",X"0E",X"CE",X"C8",X"08",X"C8",X"CE",
		X"01",X"02",X"03",X"03",X"01",X"01",X"01",X"00",X"08",X"C8",X"C8",X"0C",X"CC",X"C4",X"08",X"0C",
		X"01",X"01",X"01",X"03",X"03",X"02",X"01",X"03",X"00",X"00",X"C0",X"20",X"00",X"C0",X"A0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0E",X"07",X"07",X"03",X"00",X"00",X"00",
		X"03",X"07",X"0F",X"FE",X"F9",X"E0",X"19",X"F8",X"00",X"40",X"A0",X"00",X"E0",X"00",X"E0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C1",X"01",X"C3",X"03",X"06",X"07",X"0C",X"0F",
		X"91",X"F0",X"20",X"E1",X"40",X"C0",X"80",X"80",X"E0",X"00",X"C0",X"20",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"B0",X"00",X"00",X"00",X"00",X"18",
		X"00",X"01",X"03",X"07",X"0C",X"1B",X"10",X"00",X"07",X"FB",X"FC",X"0F",X"FD",X"FD",X"78",X"00",
		X"00",X"00",X"D0",X"94",X"DC",X"EC",X"78",X"3C",X"01",X"18",X"1C",X"0C",X"0E",X"0E",X"0F",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"0C",X"0F",X"0F",X"6F",X"07",X"07",X"6F",
		X"18",X"00",X"9C",X"0E",X"6F",X"1F",X"0F",X"0F",X"0F",X"6F",X"6F",X"0F",X"6F",X"6F",X"0F",X"6F",
		X"1F",X"5F",X"0F",X"AF",X"0F",X"0F",X"0F",X"0F",X"00",X"60",X"90",X"10",X"90",X"60",X"00",X"00",
		X"0F",X"0F",X"9F",X"0E",X"0C",X"98",X"00",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"0F",X"0E",X"0E",X"0C",X"1C",X"19",X"01",X"30",X"F0",X"20",X"20",X"C0",X"C0",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"08",X"08",X"04",X"04",X"04",X"08",X"00",
		X"00",X"00",X"01",X"01",X"05",X"08",X"0D",X"4F",X"40",X"80",X"80",X"C0",X"00",X"00",X"00",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"0A",X"40",X"0E",X"00",X"0E",X"4C",
		X"FC",X"FF",X"FF",X"FF",X"FA",X"F7",X"F6",X"FB",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"10",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"0A",X"00",X"0E",X"0C",X"00",X"07",
		X"FF",X"FF",X"FE",X"FE",X"FC",X"F0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"CC",X"04",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"FE",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"0F",X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"C0",X"70",X"1C",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"C0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"1C",X"07",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"C0",X"F0",X"FC",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"7F",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"E0",X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"FF",X"FF",X"CF",X"83",X"83",X"83",X"83",X"83",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"0F",X"0F",
		X"EC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FE",X"FE",X"E3",X"E3",X"E3",X"E3",X"E3",X"E3",X"E3",X"E3",
		X"0F",X"0F",X"0F",X"0F",X"07",X"07",X"07",X"07",X"FE",X"FE",X"FE",X"FE",X"FF",X"FF",X"9F",X"07",
		X"FB",X"CF",X"83",X"83",X"83",X"83",X"83",X"E7",X"07",X"07",X"03",X"03",X"03",X"03",X"03",X"03",
		X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"07",X"07",X"07",X"07",X"C7",X"C7",X"C7",X"C7",
		X"01",X"01",X"01",X"FF",X"FF",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"E0",X"F0",X"F0",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"70",X"70",X"70",X"F0",X"F0",X"70",X"70",X"70",X"7E",X"1E",X"06",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"70",X"10",X"00",X"00",X"00",X"C0",X"C0",X"C0",X"FF",X"FF",X"C0",X"C0",X"C0",
		X"C7",X"C7",X"C7",X"C7",X"F7",X"9F",X"07",X"07",X"07",X"07",X"07",X"CF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"3F",X"0F",X"03",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"C0",X"C0",X"F0",X"FF",X"00",
		X"FF",X"30",X"FC",X"3F",X"00",X"3F",X"C0",X"00",X"FF",X"00",X"0F",X"F0",X"30",X"1C",X"07",X"00",
		X"FF",X"0C",X"07",X"01",X"00",X"00",X"00",X"00",X"FF",X"F0",X"FC",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"03",X"00",X"FF",X"00",X"00",X"00",X"00",X"FF",X"38",X"0E",X"03",X"00",X"00",X"00",X"00",
		X"FF",X"0C",X"07",X"01",X"00",X"C0",X"F0",X"FC",X"FF",X"C0",X"F0",X"FC",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F3",X"E0",X"E0",X"E0",X"E0",X"E0",X"F8",X"F8",
		X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"FE",X"F3",X"E0",X"E0",X"E0",X"E0",X"E0",X"F9",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"60",X"00",X"C1",X"FF",X"00",X"00",X"00",X"07",X"10",X"1C",X"1F",X"1F",
		X"00",X"40",X"40",X"40",X"60",X"60",X"60",X"70",X"70",X"70",X"78",X"78",X"78",X"7C",X"7C",X"7C",
		X"7E",X"7E",X"7E",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"C0",X"C0",X"C0",X"E0",X"E0",X"E0",X"F0",
		X"F0",X"F0",X"F8",X"F8",X"F8",X"FC",X"FC",X"FC",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"01",X"01",X"03",X"03",X"03",X"03",X"03",X"03",X"07",X"07",X"07",X"07",X"07",X"07",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"1F",X"1F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",
		X"07",X"07",X"07",X"07",X"07",X"07",X"03",X"01",X"FE",X"FE",X"7E",X"7C",X"3C",X"1C",X"1C",X"08",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"70",X"70",X"30",X"30",X"F0",X"F0",X"F0",
		X"7E",X"1E",X"06",X"00",X"00",X"FF",X"FF",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"10",X"40",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"03",X"0E",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"0E",X"1C",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"70",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"03",X"0F",X"1E",X"18",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"0E",X"1E",X"7C",
		X"F8",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"0F",X"1F",X"7E",X"F8",X"F0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"C0",X"C0",X"C0",X"C0",
		X"00",X"00",X"00",X"00",X"01",X"03",X"0F",X"1F",X"7F",X"FE",X"FC",X"F0",X"E0",X"80",X"00",X"00",
		X"00",X"01",X"03",X"0F",X"1F",X"7F",X"FF",X"FC",X"0F",X"1F",X"7F",X"FF",X"FE",X"F8",X"F0",X"C0",
		X"00",X"00",X"00",X"01",X"03",X"07",X"07",X"07",X"07",X"06",X"04",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"08",X"10",X"40",X"80",X"00",X"00",
		X"02",X"0E",X"1C",X"30",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"60",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"0F",X"1E",X"38",X"30",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"1C",X"7C",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",
		X"03",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"0E",X"1E",X"7E",X"FE",X"FC",X"F0",X"E0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"01",X"03",X"0F",X"1F",X"7F",X"7F",X"7E",X"7C",X"70",X"60",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"18",X"20",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"02",X"0E",X"18",X"10",X"00",X"02",X"0E",X"1C",X"70",X"60",X"00",X"00",X"00",
		X"40",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"0F",X"1E",X"78",X"F0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"70",X"F0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"1E",X"1C",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",
		X"F0",X"F0",X"F0",X"F0",X"E0",X"80",X"00",X"00",X"FF",X"FE",X"FC",X"F0",X"E0",X"80",X"00",X"00",
		X"01",X"03",X"07",X"07",X"07",X"07",X"07",X"04",X"00",X"02",X"08",X"10",X"00",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"08",X"00",X"0C",X"1C",X"70",X"E0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",
		X"C0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"1F",X"7E",X"7C",X"70",X"60",X"00",X"00",X"00",
		X"00",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"02",X"00",X"10",X"00",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"18",X"30",X"00",X"00",X"08",X"18",X"70",X"E0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"1C",X"7C",X"FC",X"00",X"00",X"00",X"08",X"18",X"78",X"F8",X"F8",
		X"0F",X"0F",X"0F",X"0F",X"0E",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",
		X"10",X"60",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"0E",X"1E",X"78",X"F0",X"C0",
		X"0F",X"0E",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"1C",X"7C",X"F8",X"F0",X"C0",
		X"00",X"00",X"01",X"03",X"0F",X"1F",X"1F",X"1C",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"02",X"00",X"10",X"20",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"18",X"70",X"40",X"00",X"00",X"10",X"70",X"E0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"00",X"00",X"00",X"00",X"08",X"18",X"78",X"F0",X"C0",
		X"0F",X"1E",X"1C",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"70",X"F0",X"F0",X"C0",
		X"08",X"18",X"78",X"F8",X"F8",X"F8",X"F0",X"C0",X"00",X"00",X"01",X"03",X"0F",X"1F",X"3F",X"3F",
		X"00",X"00",X"04",X"10",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"18",X"70",X"40",
		X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"04",X"00",X"00",X"00",X"00",X"10",X"70",X"F0",X"C0",
		X"0F",X"1E",X"7C",X"70",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"C0",X"C0",X"C0",
		X"03",X"07",X"07",X"07",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"80",
		X"FF",X"FF",X"10",X"08",X"08",X"04",X"04",X"04",X"04",X"04",X"04",X"08",X"08",X"10",X"20",X"C0",
		X"00",X"00",X"00",X"10",X"70",X"F0",X"F0",X"F0",X"1F",X"7F",X"FF",X"FF",X"FE",X"F8",X"F0",X"C0",
		X"10",X"70",X"F0",X"F0",X"F0",X"F0",X"F0",X"C0",X"00",X"00",X"01",X"03",X"0F",X"1F",X"7F",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"10",X"70",X"F0",X"03",X"FE",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0C",X"C0",X"F1",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"60",X"F8",X"FC",X"FC",X"FE",X"FF",X"FB",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",
		X"3F",X"3F",X"3F",X"3F",X"3E",X"38",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"03",X"07",X"07",X"07",X"07",X"07",X"07",X"06",X"04",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"D0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C5",X"F8",X"E0",X"C0",X"C0",X"DF",X"FF",X"FF",X"70",X"38",X"B8",X"DC",X"FC",X"F8",X"FC",X"FC",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"8F",X"FF",X"FF",X"FF",X"FD",X"FF",X"00",X"00",X"00",X"80",X"E0",X"F0",X"F8",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E7",X"F3",X"C9",X"40",X"20",X"00",X"00",X"00",
		X"80",X"E0",X"F8",X"70",X"38",X"10",X"00",X"00",X"00",X"1C",X"62",X"81",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"81",X"62",X"1C",X"00",X"00",X"E0",X"F8",X"FE",X"0F",X"07",X"03",X"03",
		X"01",X"02",X"03",X"03",X"01",X"01",X"01",X"00",X"01",X"01",X"01",X"03",X"03",X"02",X"01",X"03",
		X"03",X"07",X"0F",X"FE",X"F9",X"E0",X"19",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"80",X"80",X"C0",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"CC",X"04",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"3F",X"3F",X"7F",X"7F",X"7F",X"7F",
		X"00",X"F8",X"E4",X"F4",X"F2",X"FA",X"FA",X"FA",X"7F",X"7F",X"3F",X"0F",X"0D",X"00",X"00",X"00",
		X"FA",X"FA",X"BA",X"3A",X"10",X"10",X"00",X"00",X"00",X"00",X"04",X"7E",X"00",X"00",X"3C",X"42",
		X"00",X"64",X"42",X"52",X"4C",X"00",X"3C",X"42",X"00",X"2E",X"4A",X"4A",X"32",X"00",X"3C",X"42",
		X"00",X"02",X"62",X"1A",X"06",X"00",X"3C",X"42",X"7E",X"00",X"3C",X"42",X"42",X"3C",X"00",X"3C",
		X"42",X"3C",X"00",X"3C",X"42",X"42",X"3C",X"00",X"42",X"42",X"3C",X"00",X"3C",X"42",X"42",X"3C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"08",X"5B",X"7F",
		X"00",X"00",X"07",X"1F",X"38",X"00",X"58",X"FC",X"00",X"00",X"00",X"80",X"C0",X"40",X"00",X"30",
		X"18",X"18",X"30",X"B0",X"B0",X"30",X"70",X"70",X"7F",X"FF",X"FF",X"FD",X"7C",X"78",X"FA",X"F2",
		X"F8",X"D0",X"45",X"0F",X"1F",X"1E",X"3C",X"3C",X"18",X"0C",X"C4",X"E0",X"30",X"10",X"00",X"00",
		X"71",X"79",X"78",X"7A",X"3E",X"3E",X"2C",X"0C",X"F3",X"F3",X"E1",X"61",X"70",X"20",X"20",X"20",
		X"18",X"39",X"33",X"13",X"01",X"21",X"60",X"E0",X"F0",X"E0",X"F8",X"F0",X"FC",X"F0",X"A0",X"00",
		X"0C",X"0D",X"0F",X"0B",X"03",X"01",X"01",X"00",X"02",X"06",X"06",X"03",X"93",X"9B",X"9F",X"C9",
		X"A7",X"33",X"10",X"02",X"01",X"00",X"00",X"00",X"24",X"FE",X"CC",X"00",X"C0",X"E0",X"70",X"00",
		X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"07",X"07",X"1F",X"7F",X"F3",X"C0",X"C0",X"80",X"08",
		X"C0",X"F0",X"F8",X"3E",X"0F",X"07",X"03",X"21",X"00",X"00",X"00",X"00",X"80",X"E0",X"F0",X"B8",
		X"06",X"06",X"07",X"0F",X"0E",X"0E",X"0C",X"0C",X"00",X"01",X"00",X"00",X"08",X"00",X"40",X"01",
		X"00",X"08",X"00",X"00",X"20",X"02",X"00",X"00",X"1C",X"1C",X"0E",X"46",X"06",X"07",X"03",X"03",
		X"0E",X"0E",X"0E",X"0C",X"0C",X"0E",X"06",X"07",X"00",X"00",X"10",X"00",X"00",X"02",X"20",X"00",
		X"08",X"00",X"40",X"00",X"00",X"12",X"00",X"00",X"87",X"0F",X"0F",X"0F",X"47",X"07",X"07",X"0E",
		X"07",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"C7",X"EF",X"FF",X"78",X"00",X"00",
		X"40",X"00",X"90",X"F8",X"FC",X"7E",X"1F",X"03",X"0E",X"8E",X"0E",X"1C",X"3C",X"78",X"F0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"28",X"28",X"11",X"00",X"00",X"40",X"40",X"40",X"20",X"0F",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"10",X"80",X"E0",X"03",X"07",X"07",X"0F",X"0F",X"0F",X"19",X"0C",
		X"FF",X"FF",X"FF",X"EF",X"47",X"1F",X"BE",X"0C",X"F8",X"F8",X"FC",X"FC",X"FC",X"F4",X"29",X"78",
		X"04",X"36",X"E9",X"E3",X"F3",X"F1",X"F8",X"F8",X"04",X"61",X"F0",X"F2",X"FB",X"F9",X"7D",X"FF",
		X"F8",X"FC",X"9C",X"38",X"18",X"50",X"24",X"CC",X"78",X"11",X"0F",X"03",X"01",X"20",X"00",X"18",
		X"5F",X"17",X"87",X"1F",X"FF",X"0F",X"01",X"00",X"F8",X"FC",X"FE",X"FE",X"CE",X"84",X"C0",X"70",
		X"00",X"00",X"01",X"00",X"20",X"20",X"10",X"03",X"00",X"00",X"00",X"00",X"40",X"42",X"00",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"07",X"4F",X"1D",X"3F",X"7F",X"4F",X"6B",X"E6",
		X"FF",X"FF",X"FF",X"CF",X"C0",X"F1",X"07",X"3F",X"00",X"40",X"70",X"60",X"70",X"7E",X"77",X"7F",
		X"F0",X"7A",X"38",X"BC",X"BC",X"9D",X"DC",X"7E",X"83",X"C0",X"61",X"63",X"70",X"3F",X"3F",X"0F",
		X"3F",X"4E",X"FA",X"78",X"79",X"F2",X"FE",X"F8",X"7E",X"37",X"31",X"18",X"5C",X"07",X"11",X"00",
		X"03",X"82",X"FF",X"7D",X"30",X"18",X"C3",X"7E",X"FC",X"24",X"34",X"FC",X"1C",X"79",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"80",X"00",X"20",X"70",X"FE",X"7F",X"1F",X"0F",X"0B",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"C0",X"E0",X"80",X"80",X"9F",X"C7",X"21",X"18",X"00",X"00",
		X"41",X"E0",X"F8",X"FF",X"FF",X"7F",X"1F",X"07",X"D0",X"00",X"00",X"00",X"80",X"E0",X"F8",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"38",X"39",X"31",X"38",X"3E",X"3F",X"1F",
		X"FC",X"7E",X"1B",X"20",X"28",X"04",X"80",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"47",X"41",X"00",X"00",X"01",X"01",X"08",X"08",X"70",X"F0",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"00",X"01",X"03",X"03",X"07",X"3F",X"FF",X"FF",X"FF",X"C0",X"80",X"00",X"00",
		X"80",X"E0",X"F8",X"FC",X"7E",X"1F",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"06",X"0E",X"7C",X"7C",X"7C",X"FC",X"F8",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"07",X"03",X"03",X"03",X"03",X"01",X"01",X"80",X"C0",X"C0",X"C0",X"C0",X"E0",X"E0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"07",X"06",X"00",X"00",X"00",
		X"01",X"01",X"61",X"F1",X"61",X"01",X"01",X"01",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"FF",X"BF",X"9C",X"83",X"A0",X"F8",X"FF",X"E1",X"FE",X"FE",X"00",X"C1",X"33",X"03",X"01",X"20",
		X"0F",X"EF",X"E0",X"F0",X"F0",X"F8",X"F8",X"F8",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"20",
		X"FF",X"FF",X"00",X"00",X"01",X"00",X"20",X"10",X"FF",X"FF",X"7F",X"FF",X"FE",X"FE",X"FD",X"FF",
		X"E7",X"83",X"1E",X"7E",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"30",X"78",X"7C",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FD",X"F9",X"7B",X"31",X"10",X"00",X"FF",X"FF",
		X"F7",X"F7",X"F7",X"F7",X"F0",X"60",X"2F",X"8F",X"E0",X"C0",X"80",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"B8",X"04",X"71",X"39",X"10",X"00",X"C2",X"E7",
		X"E0",X"48",X"1C",X"F7",X"F8",X"6E",X"11",X"7F",X"C0",X"00",X"60",X"00",X"00",X"00",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
