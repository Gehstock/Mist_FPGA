library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_PGM_2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_PGM_2 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"3A",X"00",X"50",X"CB",X"77",X"20",X"04",X"21",X"2C",X"4C",X"C9",X"21",X"B0",X"42",X"11",X"20",
		X"81",X"CD",X"ED",X"01",X"C3",X"14",X"80",X"C0",X"50",X"28",X"F0",X"18",X"EA",X"05",X"71",X"00",
		X"0F",X"01",X"05",X"31",X"00",X"0F",X"01",X"05",X"11",X"00",X"0F",X"01",X"05",X"E0",X"00",X"0F",
		X"01",X"10",X"AF",X"CD",X"60",X"32",X"C3",X"DE",X"23",X"CD",X"3A",X"24",X"32",X"87",X"4C",X"11",
		X"87",X"4C",X"C9",X"7C",X"47",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"32",X"7F",X"4C",X"7D",X"0F",
		X"0F",X"0F",X"0F",X"E6",X"0F",X"4F",X"78",X"E6",X"0F",X"0F",X"0F",X"0F",X"0F",X"B1",X"32",X"7E",
		X"4C",X"C9",X"CD",X"0C",X"87",X"36",X"00",X"23",X"7D",X"A7",X"20",X"F9",X"C9",X"02",X"C3",X"00",
		X"08",X"0F",X"07",X"79",X"00",X"08",X"0F",X"07",X"4B",X"00",X"08",X"0F",X"02",X"93",X"00",X"08",
		X"0F",X"07",X"88",X"00",X"08",X"0F",X"07",X"4B",X"00",X"08",X"0F",X"02",X"33",X"00",X"08",X"0F",
		X"07",X"88",X"00",X"08",X"0F",X"07",X"4B",X"00",X"08",X"0F",X"02",X"D2",X"00",X"08",X"0F",X"07",
		X"00",X"00",X"08",X"02",X"07",X"D2",X"00",X"08",X"03",X"07",X"D2",X"00",X"08",X"03",X"07",X"D2",
		X"00",X"08",X"03",X"07",X"D2",X"00",X"08",X"03",X"07",X"D2",X"00",X"08",X"03",X"07",X"D2",X"00",
		X"08",X"03",X"10",X"21",X"00",X"00",X"22",X"03",X"4C",X"CD",X"9C",X"19",X"3E",X"10",X"CD",X"10",
		X"1D",X"21",X"E1",X"80",X"22",X"03",X"4C",X"21",X"16",X"87",X"CD",X"3F",X"87",X"3A",X"FD",X"4F",
		X"C9",X"07",X"A5",X"00",X"0A",X"0F",X"07",X"56",X"00",X"0A",X"0F",X"07",X"27",X"00",X"0A",X"0F",
		X"07",X"88",X"00",X"0A",X"0F",X"07",X"4B",X"00",X"0A",X"05",X"07",X"4B",X"00",X"0A",X"05",X"07",
		X"4B",X"00",X"0F",X"1F",X"10",X"FF",X"FF",X"F5",X"C5",X"47",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",
		X"FE",X"0A",X"30",X"10",X"77",X"78",X"E6",X"0F",X"FE",X"0A",X"30",X"0C",X"01",X"E0",X"FF",X"09",
		X"06",X"49",X"40",X"43",X"41",X"4E",X"40",X"4E",X"4F",X"54",X"40",X"52",X"55",X"4E",X"5B",X"5B",
		X"5B",X"FF",X"06",X"20",X"1A",X"E5",X"CD",X"07",X"81",X"E1",X"23",X"13",X"7B",X"32",X"C0",X"50",
		X"A7",X"C8",X"05",X"20",X"EF",X"C5",X"01",X"80",X"FF",X"09",X"C1",X"18",X"E5",X"02",X"D2",X"00",
		X"0D",X"0F",X"03",X"22",X"00",X"08",X"07",X"02",X"D2",X"00",X"0D",X"07",X"02",X"22",X"00",X"0D",
		X"07",X"03",X"93",X"00",X"08",X"07",X"03",X"22",X"00",X"08",X"07",X"03",X"D2",X"00",X"08",X"07",
		X"02",X"D2",X"00",X"0D",X"0F",X"03",X"22",X"00",X"08",X"07",X"02",X"D2",X"00",X"0D",X"07",X"02",
		X"22",X"00",X"0D",X"07",X"03",X"93",X"00",X"08",X"07",X"03",X"22",X"00",X"08",X"07",X"03",X"D2",
		X"00",X"08",X"07",X"02",X"62",X"00",X"0D",X"0F",X"03",X"62",X"00",X"08",X"07",X"02",X"62",X"00",
		X"0D",X"07",X"02",X"C1",X"00",X"0D",X"07",X"03",X"93",X"00",X"08",X"07",X"03",X"62",X"00",X"08",
		X"07",X"03",X"D2",X"00",X"08",X"07",X"02",X"62",X"00",X"0D",X"0F",X"03",X"62",X"00",X"08",X"07",
		X"02",X"62",X"00",X"0D",X"07",X"02",X"C1",X"00",X"0D",X"07",X"03",X"93",X"00",X"08",X"07",X"03",
		X"62",X"00",X"08",X"07",X"03",X"D2",X"00",X"08",X"07",X"02",X"E1",X"00",X"0D",X"0F",X"03",X"62",
		X"00",X"08",X"07",X"02",X"E1",X"00",X"0D",X"07",X"02",X"D2",X"00",X"0D",X"07",X"03",X"C3",X"00",
		X"08",X"07",X"03",X"62",X"00",X"08",X"07",X"03",X"D2",X"00",X"08",X"07",X"02",X"E1",X"00",X"0D",
		X"0F",X"03",X"62",X"00",X"08",X"07",X"02",X"E1",X"00",X"0D",X"07",X"02",X"D2",X"00",X"0D",X"07",
		X"03",X"C3",X"00",X"08",X"07",X"03",X"62",X"00",X"08",X"07",X"03",X"D2",X"00",X"08",X"07",X"02",
		X"22",X"00",X"0D",X"0F",X"03",X"B2",X"00",X"08",X"07",X"02",X"22",X"00",X"0D",X"07",X"02",X"B2",
		X"00",X"0D",X"07",X"03",X"44",X"00",X"08",X"07",X"03",X"B2",X"00",X"08",X"07",X"03",X"33",X"00",
		X"08",X"07",X"02",X"22",X"00",X"0D",X"0F",X"03",X"B2",X"00",X"08",X"07",X"02",X"22",X"00",X"0D",
		X"07",X"02",X"B2",X"00",X"0D",X"07",X"03",X"44",X"00",X"08",X"07",X"03",X"B2",X"00",X"08",X"07",
		X"03",X"33",X"00",X"08",X"07",X"02",X"D2",X"00",X"0D",X"0F",X"03",X"22",X"00",X"08",X"07",X"03",
		X"D2",X"00",X"08",X"07",X"02",X"22",X"00",X"0D",X"07",X"03",X"93",X"00",X"08",X"07",X"03",X"22",
		X"00",X"08",X"07",X"03",X"D2",X"00",X"08",X"07",X"02",X"D2",X"00",X"0D",X"0F",X"03",X"22",X"00",
		X"08",X"07",X"03",X"D2",X"00",X"08",X"07",X"02",X"22",X"00",X"0D",X"07",X"03",X"93",X"00",X"08",
		X"07",X"03",X"22",X"00",X"08",X"07",X"03",X"D2",X"00",X"08",X"07",X"02",X"62",X"00",X"0D",X"0F",
		X"03",X"62",X"00",X"08",X"07",X"03",X"D2",X"00",X"08",X"07",X"02",X"93",X"00",X"0D",X"07",X"03",
		X"93",X"00",X"08",X"07",X"03",X"62",X"00",X"08",X"07",X"03",X"D2",X"00",X"08",X"07",X"02",X"62",
		X"00",X"0D",X"0F",X"03",X"62",X"00",X"08",X"07",X"03",X"D2",X"00",X"08",X"07",X"02",X"93",X"00",
		X"0D",X"07",X"03",X"93",X"00",X"08",X"07",X"03",X"62",X"00",X"08",X"07",X"03",X"D2",X"00",X"08",
		X"07",X"02",X"E1",X"00",X"0D",X"0F",X"03",X"62",X"00",X"08",X"07",X"03",X"D2",X"00",X"08",X"07",
		X"02",X"62",X"00",X"0D",X"07",X"03",X"C3",X"00",X"08",X"07",X"03",X"62",X"00",X"08",X"07",X"03",
		X"D2",X"00",X"08",X"07",X"02",X"E1",X"00",X"0D",X"0F",X"03",X"62",X"00",X"08",X"07",X"03",X"D2",
		X"00",X"08",X"07",X"02",X"62",X"00",X"0D",X"07",X"03",X"C3",X"00",X"08",X"07",X"03",X"62",X"00",
		X"08",X"07",X"03",X"D2",X"00",X"08",X"07",X"02",X"22",X"00",X"0D",X"0F",X"03",X"B2",X"00",X"08",
		X"07",X"03",X"33",X"00",X"08",X"07",X"02",X"B2",X"00",X"0D",X"07",X"03",X"44",X"00",X"08",X"07",
		X"03",X"B2",X"00",X"08",X"07",X"03",X"33",X"00",X"08",X"07",X"02",X"22",X"00",X"0D",X"0F",X"03",
		X"B2",X"00",X"08",X"07",X"03",X"33",X"00",X"08",X"07",X"02",X"B2",X"00",X"0D",X"07",X"03",X"44",
		X"00",X"08",X"07",X"03",X"B2",X"00",X"08",X"07",X"03",X"33",X"00",X"08",X"07",X"10",X"D2",X"00",
		X"0F",X"0F",X"02",X"22",X"00",X"0F",X"0F",X"02",X"62",X"00",X"0F",X"0F",X"02",X"B2",X"00",X"0F",
		X"0F",X"10",X"03",X"44",X"00",X"08",X"0F",X"03",X"44",X"00",X"08",X"0F",X"03",X"C4",X"00",X"08",
		X"07",X"03",X"A5",X"00",X"08",X"0F",X"03",X"56",X"00",X"08",X"07",X"03",X"27",X"00",X"08",X"0F",
		X"03",X"27",X"00",X"08",X"07",X"03",X"56",X"00",X"08",X"07",X"03",X"27",X"00",X"08",X"07",X"03",
		X"56",X"00",X"08",X"07",X"03",X"A5",X"00",X"08",X"07",X"03",X"C4",X"00",X"08",X"07",X"03",X"44",
		X"00",X"08",X"0F",X"03",X"44",X"00",X"08",X"0F",X"03",X"C4",X"00",X"08",X"07",X"03",X"A5",X"00",
		X"08",X"0F",X"03",X"56",X"00",X"08",X"07",X"03",X"27",X"00",X"08",X"0F",X"03",X"27",X"00",X"08",
		X"07",X"03",X"56",X"00",X"08",X"07",X"03",X"27",X"00",X"08",X"07",X"03",X"88",X"00",X"08",X"07",
		X"03",X"79",X"00",X"08",X"07",X"03",X"88",X"00",X"08",X"07",X"03",X"79",X"00",X"08",X"0F",X"03",
		X"79",X"00",X"08",X"07",X"03",X"9A",X"00",X"08",X"07",X"03",X"6B",X"00",X"08",X"0F",X"03",X"6B",
		X"00",X"08",X"07",X"03",X"9A",X"00",X"08",X"07",X"03",X"6B",X"00",X"08",X"0F",X"03",X"6B",X"00",
		X"08",X"07",X"03",X"9A",X"00",X"08",X"07",X"03",X"6B",X"00",X"08",X"07",X"03",X"9A",X"00",X"08",
		X"07",X"03",X"79",X"00",X"08",X"07",X"03",X"88",X"00",X"08",X"07",X"03",X"27",X"00",X"08",X"0F",
		X"03",X"27",X"00",X"08",X"07",X"03",X"88",X"00",X"08",X"07",X"03",X"56",X"00",X"08",X"0F",X"03",
		X"56",X"00",X"08",X"07",X"03",X"27",X"00",X"08",X"07",X"03",X"56",X"00",X"08",X"07",X"03",X"A5",
		X"00",X"08",X"07",X"03",X"C4",X"00",X"08",X"07",X"03",X"55",X"00",X"08",X"07",X"03",X"A5",X"00",
		X"08",X"0F",X"03",X"A5",X"00",X"08",X"0F",X"03",X"44",X"00",X"08",X"0F",X"03",X"C4",X"00",X"0F",
		X"07",X"03",X"A5",X"00",X"08",X"0F",X"03",X"56",X"00",X"08",X"07",X"03",X"A5",X"00",X"08",X"07",
		X"03",X"C4",X"00",X"08",X"07",X"03",X"44",X"00",X"08",X"0F",X"03",X"C4",X"00",X"08",X"07",X"03",
		X"A5",X"00",X"08",X"0F",X"03",X"56",X"00",X"08",X"07",X"03",X"A5",X"00",X"08",X"07",X"03",X"56",
		X"00",X"08",X"07",X"03",X"27",X"00",X"08",X"0F",X"03",X"56",X"00",X"08",X"07",X"03",X"27",X"00",
		X"08",X"0F",X"03",X"56",X"00",X"08",X"07",X"03",X"A5",X"00",X"08",X"07",X"03",X"56",X"00",X"08",
		X"07",X"03",X"27",X"00",X"08",X"0F",X"03",X"88",X"00",X"08",X"07",X"03",X"79",X"00",X"08",X"0F",
		X"03",X"88",X"00",X"08",X"07",X"03",X"27",X"00",X"08",X"07",X"03",X"88",X"00",X"08",X"07",X"03",
		X"79",X"00",X"08",X"0F",X"03",X"6B",X"00",X"08",X"07",X"03",X"2E",X"00",X"08",X"0F",X"03",X"CC",
		X"00",X"08",X"07",X"03",X"6B",X"00",X"08",X"07",X"03",X"CC",X"00",X"08",X"07",X"03",X"2E",X"00",
		X"08",X"0F",X"03",X"2E",X"00",X"08",X"07",X"03",X"CC",X"00",X"08",X"0F",X"03",X"2E",X"00",X"08",
		X"07",X"03",X"CC",X"00",X"08",X"07",X"03",X"2E",X"00",X"08",X"07",X"03",X"6B",X"00",X"08",X"0F",
		X"03",X"88",X"00",X"08",X"0F",X"03",X"27",X"00",X"08",X"07",X"03",X"56",X"00",X"08",X"0F",X"03",
		X"27",X"00",X"08",X"07",X"03",X"A5",X"00",X"08",X"0F",X"03",X"44",X"00",X"08",X"0F",X"03",X"A5",
		X"00",X"08",X"0F",X"03",X"A5",X"00",X"08",X"0F",X"10",X"02",X"62",X"00",X"09",X"07",X"02",X"62",
		X"00",X"09",X"07",X"04",X"03",X"00",X"06",X"07",X"04",X"33",X"00",X"06",X"07",X"04",X"93",X"00",
		X"06",X"07",X"02",X"91",X"00",X"09",X"07",X"04",X"03",X"00",X"06",X"07",X"02",X"B2",X"00",X"09",
		X"07",X"02",X"62",X"00",X"09",X"07",X"02",X"62",X"00",X"09",X"07",X"04",X"03",X"00",X"06",X"07",
		X"04",X"33",X"00",X"06",X"07",X"04",X"93",X"00",X"06",X"07",X"02",X"91",X"00",X"09",X"07",X"04",
		X"03",X"00",X"06",X"07",X"02",X"B2",X"00",X"09",X"07",X"04",X"33",X"00",X"06",X"07",X"04",X"33",
		X"00",X"06",X"07",X"04",X"04",X"00",X"06",X"07",X"04",X"44",X"00",X"06",X"07",X"04",X"C4",X"00",
		X"06",X"07",X"04",X"44",X"00",X"06",X"07",X"04",X"04",X"00",X"06",X"07",X"04",X"93",X"00",X"06",
		X"07",X"04",X"33",X"00",X"06",X"07",X"04",X"33",X"00",X"06",X"07",X"04",X"04",X"00",X"06",X"07",
		X"04",X"44",X"00",X"06",X"07",X"04",X"C4",X"00",X"06",X"07",X"04",X"44",X"00",X"06",X"07",X"04",
		X"04",X"00",X"06",X"07",X"04",X"93",X"00",X"10",X"07",X"10",X"07",X"62",X"00",X"06",X"07",X"07",
		X"79",X"00",X"06",X"07",X"07",X"0C",X"00",X"06",X"07",X"07",X"79",X"00",X"06",X"07",X"07",X"2E",
		X"00",X"06",X"07",X"07",X"79",X"00",X"06",X"07",X"07",X"0C",X"00",X"06",X"07",X"07",X"79",X"00",
		X"06",X"07",X"07",X"62",X"00",X"06",X"07",X"07",X"79",X"00",X"06",X"07",X"07",X"0C",X"00",X"06",
		X"07",X"07",X"79",X"00",X"06",X"07",X"07",X"2E",X"00",X"06",X"07",X"07",X"79",X"00",X"06",X"07",
		X"07",X"0C",X"00",X"06",X"07",X"07",X"79",X"00",X"06",X"07",X"07",X"91",X"00",X"06",X"07",X"07",
		X"79",X"00",X"06",X"07",X"07",X"CC",X"00",X"06",X"07",X"07",X"79",X"00",X"06",X"07",X"07",X"FF",
		X"00",X"06",X"07",X"07",X"79",X"00",X"06",X"07",X"07",X"CC",X"00",X"06",X"07",X"07",X"79",X"00",
		X"06",X"07",X"07",X"91",X"00",X"06",X"07",X"07",X"79",X"00",X"06",X"07",X"07",X"CC",X"00",X"06",
		X"07",X"07",X"79",X"00",X"06",X"07",X"07",X"FF",X"00",X"06",X"07",X"07",X"79",X"00",X"06",X"07",
		X"07",X"CC",X"00",X"06",X"07",X"07",X"79",X"00",X"06",X"07",X"10",X"02",X"00",X"00",X"10",X"02",
		X"02",X"79",X"00",X"10",X"0F",X"02",X"A7",X"00",X"08",X"0F",X"07",X"4B",X"00",X"08",X"0F",X"07",
		X"88",X"00",X"08",X"0F",X"02",X"27",X"00",X"08",X"0F",X"07",X"4B",X"00",X"08",X"0F",X"07",X"CC",
		X"00",X"08",X"0F",X"02",X"9A",X"00",X"08",X"0F",X"07",X"88",X"00",X"08",X"0F",X"07",X"4B",X"00",
		X"08",X"0F",X"02",X"4B",X"00",X"08",X"03",X"07",X"4B",X"00",X"08",X"03",X"07",X"4B",X"00",X"08",
		X"03",X"02",X"4B",X"00",X"08",X"03",X"07",X"4B",X"00",X"08",X"03",X"07",X"4B",X"00",X"08",X"03",
		X"10",X"D2",X"00",X"08",X"03",X"10",X"CD",X"01",X"07",X"C3",X"C6",X"06",X"21",X"00",X"00",X"22",
		X"3A",X"4C",X"21",X"41",X"4C",X"C9",X"03",X"27",X"00",X"0A",X"0F",X"03",X"A7",X"00",X"0A",X"0F",
		X"03",X"88",X"00",X"0A",X"0F",X"03",X"79",X"00",X"0A",X"0F",X"03",X"4B",X"00",X"0A",X"05",X"03",
		X"4B",X"00",X"0A",X"05",X"03",X"4B",X"00",X"0A",X"0F",X"03",X"4B",X"00",X"0A",X"0F",X"10",X"CD",
		X"9C",X"19",X"3E",X"05",X"CD",X"10",X"1D",X"C3",X"DC",X"25",X"02",X"D2",X"00",X"0F",X"0F",X"03",
		X"88",X"00",X"0A",X"07",X"03",X"4B",X"00",X"0A",X"07",X"02",X"C1",X"00",X"0F",X"0F",X"03",X"88",
		X"00",X"0A",X"07",X"03",X"9A",X"00",X"0A",X"07",X"02",X"E1",X"00",X"0F",X"0F",X"03",X"79",X"00",
		X"0A",X"07",X"03",X"4B",X"00",X"0A",X"07",X"02",X"22",X"00",X"0F",X"0F",X"03",X"88",X"00",X"0A",
		X"07",X"03",X"9A",X"00",X"0A",X"07",X"02",X"D2",X"00",X"0F",X"0F",X"03",X"88",X"00",X"0A",X"07",
		X"03",X"4B",X"00",X"0A",X"07",X"02",X"C1",X"00",X"0F",X"0F",X"03",X"88",X"00",X"0A",X"07",X"03",
		X"9A",X"00",X"0A",X"07",X"02",X"E1",X"00",X"0F",X"0F",X"03",X"79",X"00",X"0A",X"07",X"03",X"4B",
		X"00",X"0A",X"07",X"02",X"22",X"00",X"0F",X"0F",X"03",X"88",X"00",X"0A",X"07",X"03",X"9A",X"00",
		X"0A",X"07",X"02",X"71",X"00",X"0F",X"05",X"02",X"D2",X"00",X"0F",X"05",X"02",X"71",X"00",X"0F",
		X"05",X"02",X"D2",X"00",X"0F",X"05",X"10",X"07",X"4B",X"00",X"1A",X"0F",X"07",X"4B",X"00",X"1A",
		X"07",X"07",X"CC",X"00",X"0A",X"07",X"07",X"2E",X"00",X"1A",X"0F",X"07",X"2E",X"00",X"1A",X"07",
		X"07",X"0F",X"00",X"0A",X"07",X"07",X"E0",X"10",X"1A",X"0F",X"07",X"E0",X"10",X"1A",X"07",X"07",
		X"0F",X"00",X"0A",X"07",X"07",X"E0",X"10",X"1A",X"07",X"07",X"0F",X"00",X"1A",X"07",X"07",X"2E",
		X"00",X"0A",X"07",X"07",X"CC",X"00",X"0A",X"07",X"07",X"4B",X"00",X"0A",X"0F",X"07",X"4B",X"00",
		X"0A",X"07",X"07",X"CC",X"00",X"0A",X"07",X"07",X"2E",X"00",X"0A",X"0F",X"07",X"2E",X"00",X"0A",
		X"07",X"07",X"0F",X"00",X"0A",X"07",X"07",X"E0",X"10",X"0A",X"0F",X"07",X"E0",X"10",X"0A",X"07",
		X"07",X"0F",X"00",X"0A",X"07",X"07",X"E0",X"10",X"0A",X"07",X"07",X"0F",X"00",X"0A",X"07",X"07",
		X"2E",X"00",X"0A",X"07",X"07",X"CC",X"00",X"0A",X"07",X"07",X"A5",X"00",X"1A",X"05",X"07",X"A5",
		X"00",X"1A",X"05",X"07",X"A5",X"00",X"1A",X"05",X"07",X"A5",X"00",X"1A",X"05",X"10",X"00",X"00",
		X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"0C",X"0E",X"6E",X"0E",X"0E",
		X"0E",X"0E",X"0E",X"0C",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0A",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"0A",X"00",X"70",X"00",X"00",
		X"B0",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"0F",X"8F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"08",X"00",X"00",X"00",X"00",
		X"D0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F9",X"F0",X"F0",X"F0",X"F0",X"BB",X"00",X"00",
		X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"8E",X"0E",X"0E",X"07",X"00",X"00",X"0F",X"0F",
		X"CF",X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",X"EB",X"E0",X"E0",X"E0",X"E0",X"BB",X"00",X"00",
		X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"0E",X"0E",
		X"BE",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0A",X"00",X"00",X"00",X"00",X"B8",X"00",X"00",
		X"0F",X"78",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"90",X"00",X"00",X"B6",X"00",X"00",
		X"0E",X"07",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A0",X"00",X"09",X"90",X"00",X"00",X"00",X"C0",X"E0",X"E0",X"B0",X"00",X"00",X"B6",X"00",X"00",
		X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"DD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"0F",X"0B",X"D0",X"F0",X"FF",X"FF",X"BF",X"0F",X"00",X"80",X"00",X"00",X"B6",X"00",X"00",
		X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"EE",X"0E",X"0B",X"C0",X"E0",X"EE",X"EE",X"BE",X"0E",X"00",X"60",X"00",X"00",X"B6",X"00",X"00",
		X"00",X"D0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"BA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0A",X"A0",X"00",X"08",X"00",X"A0",X"00",X"00",X"70",X"00",X"00",X"B6",X"00",X"00",
		X"00",X"C0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"B6",X"00",X"00",
		X"00",X"B8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"90",X"00",X"07",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"B6",X"00",X"00",
		X"00",X"A7",X"00",X"00",X"00",X"60",X"00",X"00",X"09",X"00",X"00",X"68",X"00",X"08",X"00",X"00",
		X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"F0",X"F0",X"B6",X"00",X"00",
		X"00",X"80",X"00",X"00",X"00",X"60",X"00",X"00",X"0B",X"00",X"00",X"D0",X"F0",X"F6",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"D0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"C0",X"E0",X"E0",X"B7",X"1E",X"22",
		X"42",X"09",X"89",X"43",X"09",X"C9",X"40",X"09",X"E2",X"42",X"08",X"E9",X"42",X"08",X"B4",X"41",
		X"08",X"F1",X"40",X"07",X"62",X"40",X"07",X"0C",X"42",X"07",X"49",X"41",X"06",X"A2",X"41",X"06",
		X"74",X"41",X"06",X"5B",X"41",X"05",X"29",X"43",X"05",X"62",X"43",X"05",X"00",X"00",X"04",X"C2",
		X"40",X"04",X"91",X"40",X"04",X"00",X"00",X"03",X"56",X"43",X"03",X"14",X"41",X"03",X"4E",X"40",
		X"02",X"42",X"41",X"02",X"00",X"00",X"02",X"AC",X"41",X"01",X"B1",X"40",X"01",X"00",X"00",X"01",
		X"BB",X"41",X"00",X"34",X"42",X"00",X"00",X"00",X"00",X"E5",X"21",X"00",X"20",X"22",X"85",X"4C",
		X"E1",X"C3",X"8B",X"20",X"06",X"7E",X"41",X"69",X"40",X"E6",X"41",X"E2",X"41",X"33",X"43",X"36",
		X"43",X"11",X"BF",X"8A",X"06",X"0E",X"21",X"CB",X"42",X"CD",X"B6",X"26",X"06",X"09",X"21",X"CD",
		X"42",X"CD",X"B6",X"26",X"3E",X"FF",X"CD",X"10",X"1D",X"CD",X"DC",X"25",X"C3",X"AF",X"01",X"53",
		X"45",X"45",X"40",X"59",X"4F",X"55",X"40",X"41",X"47",X"41",X"49",X"4E",X"3D",X"42",X"59",X"45",
		X"40",X"42",X"59",X"45",X"40",X"5B",X"CB",X"67",X"C0",X"3D",X"C9",X"02",X"D2",X"00",X"0D",X"0F",
		X"06",X"88",X"00",X"08",X"07",X"06",X"4B",X"00",X"08",X"07",X"02",X"22",X"00",X"0D",X"07",X"06",
		X"2E",X"00",X"08",X"07",X"06",X"88",X"00",X"08",X"07",X"06",X"A5",X"00",X"08",X"07",X"02",X"D2",
		X"00",X"0D",X"0F",X"06",X"88",X"00",X"08",X"07",X"06",X"4B",X"00",X"08",X"07",X"02",X"D2",X"00",
		X"0D",X"07",X"06",X"A5",X"00",X"08",X"07",X"02",X"B2",X"00",X"0D",X"07",X"06",X"A5",X"00",X"08",
		X"07",X"02",X"62",X"00",X"0D",X"0F",X"06",X"79",X"00",X"08",X"07",X"06",X"4B",X"00",X"08",X"07",
		X"02",X"C1",X"00",X"0D",X"07",X"06",X"2E",X"00",X"08",X"07",X"06",X"79",X"00",X"08",X"07",X"06",
		X"4B",X"00",X"08",X"07",X"02",X"62",X"00",X"0D",X"0F",X"06",X"79",X"00",X"08",X"07",X"06",X"4B",
		X"00",X"08",X"07",X"02",X"62",X"00",X"0D",X"07",X"06",X"A5",X"00",X"08",X"07",X"02",X"C1",X"00",
		X"0D",X"07",X"02",X"02",X"00",X"0D",X"07",X"02",X"22",X"00",X"0D",X"0F",X"06",X"88",X"00",X"08",
		X"07",X"06",X"9A",X"00",X"08",X"07",X"02",X"B2",X"00",X"0D",X"07",X"06",X"E0",X"10",X"08",X"07",
		X"06",X"88",X"00",X"08",X"07",X"06",X"9A",X"00",X"08",X"07",X"02",X"22",X"00",X"0D",X"0F",X"06",
		X"88",X"00",X"08",X"07",X"06",X"9A",X"00",X"08",X"07",X"02",X"B2",X"00",X"0D",X"07",X"06",X"E0",
		X"10",X"08",X"07",X"06",X"88",X"00",X"08",X"07",X"06",X"9A",X"00",X"08",X"07",X"02",X"D2",X"00",
		X"0D",X"0F",X"06",X"88",X"00",X"08",X"07",X"06",X"4B",X"00",X"08",X"07",X"02",X"22",X"00",X"0D",
		X"07",X"06",X"2E",X"00",X"08",X"07",X"06",X"88",X"00",X"08",X"07",X"06",X"A5",X"00",X"08",X"07",
		X"02",X"B2",X"00",X"0D",X"0F",X"06",X"88",X"00",X"08",X"07",X"06",X"9A",X"00",X"08",X"07",X"02",
		X"22",X"00",X"0D",X"07",X"06",X"E0",X"10",X"08",X"07",X"06",X"88",X"00",X"08",X"07",X"06",X"9A",
		X"00",X"08",X"07",X"02",X"D2",X"00",X"0D",X"0F",X"06",X"88",X"00",X"08",X"07",X"06",X"4B",X"00",
		X"08",X"07",X"02",X"22",X"00",X"0D",X"07",X"06",X"2E",X"00",X"08",X"07",X"06",X"88",X"00",X"08",
		X"07",X"06",X"A5",X"00",X"08",X"07",X"02",X"D2",X"00",X"0D",X"0F",X"06",X"88",X"00",X"08",X"07",
		X"06",X"4B",X"00",X"08",X"07",X"02",X"D2",X"00",X"0D",X"07",X"06",X"A5",X"00",X"08",X"07",X"02",
		X"B2",X"00",X"0D",X"07",X"06",X"A5",X"00",X"08",X"07",X"02",X"62",X"00",X"0D",X"0F",X"06",X"79",
		X"00",X"08",X"07",X"06",X"4B",X"00",X"08",X"07",X"02",X"C1",X"00",X"0D",X"07",X"06",X"2E",X"00",
		X"08",X"07",X"06",X"79",X"00",X"08",X"07",X"06",X"4B",X"00",X"08",X"07",X"02",X"62",X"00",X"0D",
		X"0F",X"06",X"79",X"00",X"08",X"07",X"06",X"4B",X"00",X"08",X"07",X"02",X"62",X"00",X"0D",X"07",
		X"06",X"A5",X"00",X"08",X"07",X"02",X"C1",X"00",X"0D",X"07",X"02",X"02",X"00",X"0D",X"07",X"02",
		X"22",X"00",X"0D",X"0F",X"06",X"88",X"00",X"08",X"07",X"06",X"9A",X"00",X"08",X"07",X"02",X"B2",
		X"00",X"0D",X"07",X"06",X"E0",X"10",X"08",X"07",X"06",X"88",X"00",X"08",X"07",X"06",X"9A",X"00",
		X"08",X"07",X"02",X"22",X"00",X"0D",X"0F",X"06",X"88",X"00",X"08",X"07",X"06",X"9A",X"00",X"08",
		X"07",X"02",X"B2",X"00",X"0D",X"07",X"06",X"E0",X"10",X"08",X"07",X"06",X"88",X"00",X"08",X"07",
		X"06",X"9A",X"00",X"08",X"07",X"02",X"D2",X"00",X"0D",X"0F",X"06",X"88",X"00",X"08",X"07",X"06",
		X"4B",X"00",X"08",X"07",X"02",X"22",X"00",X"0D",X"07",X"06",X"2E",X"00",X"08",X"07",X"06",X"88",
		X"00",X"08",X"07",X"06",X"A5",X"00",X"08",X"07",X"02",X"D2",X"00",X"0D",X"0F",X"06",X"0A",X"00",
		X"08",X"07",X"06",X"4B",X"00",X"08",X"07",X"02",X"D2",X"00",X"0D",X"07",X"06",X"2E",X"00",X"08",
		X"07",X"06",X"0A",X"00",X"08",X"07",X"06",X"4B",X"00",X"08",X"07",X"02",X"E1",X"00",X"0D",X"0F",
		X"06",X"79",X"00",X"08",X"07",X"06",X"4B",X"00",X"08",X"07",X"02",X"D2",X"00",X"0D",X"07",X"06",
		X"0F",X"00",X"08",X"07",X"06",X"79",X"00",X"08",X"07",X"06",X"4B",X"00",X"08",X"07",X"02",X"E1",
		X"00",X"0D",X"0F",X"06",X"79",X"00",X"08",X"07",X"06",X"4B",X"00",X"08",X"07",X"02",X"E1",X"00",
		X"0D",X"07",X"06",X"4B",X"00",X"08",X"07",X"02",X"02",X"00",X"0D",X"07",X"06",X"0C",X"00",X"08",
		X"07",X"02",X"22",X"00",X"0D",X"0F",X"06",X"88",X"00",X"08",X"07",X"06",X"9A",X"00",X"08",X"07",
		X"02",X"B2",X"00",X"0D",X"07",X"06",X"E0",X"10",X"08",X"07",X"06",X"88",X"00",X"08",X"07",X"06",
		X"9A",X"00",X"08",X"07",X"02",X"22",X"00",X"0D",X"0F",X"06",X"88",X"00",X"08",X"07",X"06",X"9A",
		X"00",X"08",X"07",X"02",X"22",X"00",X"0D",X"07",X"06",X"9A",X"00",X"08",X"07",X"02",X"02",X"00",
		X"0D",X"07",X"06",X"0A",X"00",X"08",X"07",X"02",X"E1",X"00",X"0D",X"0F",X"06",X"79",X"00",X"08",
		X"07",X"06",X"4B",X"00",X"08",X"07",X"02",X"D2",X"00",X"0D",X"07",X"06",X"0F",X"00",X"08",X"07",
		X"06",X"79",X"00",X"08",X"07",X"06",X"4B",X"00",X"08",X"07",X"02",X"E1",X"00",X"0D",X"0F",X"06",
		X"79",X"00",X"08",X"07",X"06",X"4B",X"00",X"08",X"07",X"02",X"E1",X"00",X"0D",X"07",X"06",X"4B",
		X"00",X"08",X"07",X"02",X"02",X"00",X"0D",X"07",X"06",X"0C",X"00",X"08",X"07",X"02",X"22",X"00",
		X"0D",X"0F",X"06",X"88",X"00",X"08",X"07",X"06",X"9A",X"00",X"08",X"07",X"02",X"B2",X"00",X"0D",
		X"07",X"06",X"E0",X"10",X"08",X"07",X"06",X"88",X"00",X"08",X"07",X"06",X"9A",X"00",X"08",X"07",
		X"02",X"22",X"00",X"0D",X"0F",X"06",X"88",X"00",X"08",X"07",X"06",X"9A",X"00",X"08",X"07",X"02",
		X"B2",X"00",X"0D",X"07",X"06",X"E0",X"10",X"08",X"07",X"06",X"88",X"00",X"08",X"07",X"06",X"9A",
		X"00",X"08",X"07",X"06",X"E0",X"10",X"08",X"1F",X"02",X"22",X"00",X"0D",X"0F",X"02",X"62",X"00",
		X"0D",X"0F",X"02",X"B2",X"00",X"0D",X"0F",X"10",X"07",X"88",X"00",X"08",X"0F",X"07",X"88",X"00",
		X"08",X"0F",X"07",X"79",X"00",X"08",X"0F",X"07",X"88",X"00",X"08",X"0F",X"07",X"27",X"00",X"08",
		X"0F",X"07",X"27",X"00",X"08",X"0F",X"07",X"56",X"00",X"08",X"0F",X"07",X"A5",X"00",X"08",X"0F",
		X"07",X"27",X"00",X"08",X"0F",X"07",X"27",X"00",X"08",X"0F",X"07",X"27",X"00",X"08",X"0F",X"07",
		X"A5",X"00",X"18",X"0F",X"07",X"C4",X"00",X"08",X"1F",X"07",X"00",X"00",X"08",X"1F",X"07",X"56",
		X"00",X"08",X"0F",X"07",X"56",X"00",X"08",X"0F",X"07",X"56",X"00",X"08",X"0F",X"07",X"27",X"00",
		X"08",X"0F",X"07",X"56",X"00",X"08",X"0F",X"07",X"A5",X"00",X"08",X"0F",X"07",X"C4",X"00",X"18",
		X"1F",X"07",X"88",X"00",X"08",X"0F",X"07",X"88",X"00",X"08",X"1F",X"07",X"79",X"00",X"08",X"0F",
		X"07",X"56",X"00",X"18",X"1F",X"07",X"00",X"00",X"08",X"1F",X"07",X"00",X"00",X"08",X"0F",X"07",
		X"88",X"00",X"18",X"0F",X"07",X"79",X"00",X"18",X"0F",X"07",X"88",X"00",X"18",X"0F",X"07",X"27",
		X"00",X"08",X"0F",X"07",X"27",X"00",X"08",X"0F",X"07",X"56",X"00",X"08",X"0F",X"07",X"A5",X"00",
		X"08",X"0F",X"07",X"27",X"00",X"08",X"0F",X"07",X"27",X"00",X"08",X"0F",X"07",X"27",X"00",X"08",
		X"0F",X"07",X"A5",X"00",X"08",X"0F",X"07",X"C4",X"00",X"18",X"1F",X"07",X"C4",X"00",X"08",X"1F",
		X"07",X"00",X"00",X"08",X"0F",X"07",X"56",X"00",X"18",X"0F",X"07",X"56",X"00",X"08",X"0F",X"07",
		X"27",X"00",X"08",X"0F",X"07",X"56",X"00",X"08",X"0F",X"07",X"A5",X"00",X"08",X"0F",X"07",X"C4",
		X"00",X"08",X"0F",X"07",X"C4",X"00",X"08",X"0F",X"07",X"A5",X"00",X"18",X"1F",X"07",X"A5",X"00",
		X"08",X"1F",X"07",X"00",X"00",X"08",X"1F",X"07",X"00",X"00",X"08",X"1F",X"07",X"79",X"00",X"08",
		X"0F",X"07",X"79",X"00",X"18",X"1F",X"07",X"79",X"00",X"08",X"0F",X"07",X"79",X"00",X"08",X"0F",
		X"07",X"9A",X"00",X"08",X"0F",X"07",X"4B",X"00",X"18",X"1F",X"07",X"9A",X"00",X"08",X"0F",X"07",
		X"9A",X"00",X"18",X"0F",X"07",X"9A",X"00",X"18",X"0F",X"07",X"79",X"00",X"08",X"0F",X"07",X"88",
		X"00",X"08",X"1F",X"07",X"88",X"00",X"08",X"1F",X"07",X"79",X"00",X"08",X"0F",X"07",X"79",X"00",
		X"18",X"0F",X"07",X"79",X"00",X"18",X"0F",X"07",X"79",X"00",X"08",X"0F",X"07",X"79",X"00",X"08",
		X"0F",X"07",X"9A",X"00",X"08",X"0F",X"07",X"4B",X"00",X"08",X"1F",X"07",X"9A",X"00",X"08",X"1F",
		X"07",X"79",X"00",X"08",X"1F",X"07",X"88",X"00",X"18",X"1F",X"07",X"88",X"00",X"08",X"1F",X"07",
		X"4B",X"00",X"08",X"1F",X"07",X"88",X"00",X"08",X"0F",X"07",X"79",X"00",X"08",X"0F",X"07",X"9A",
		X"00",X"08",X"0F",X"10",X"3A",X"40",X"4C",X"CB",X"47",X"21",X"4D",X"81",X"C0",X"C1",X"21",X"DB",
		X"8A",X"22",X"03",X"4C",X"21",X"38",X"8E",X"22",X"07",X"4C",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"CD",X"02",X"31",X"3E",X"F0",X"CD",X"C1",X"01",X"3E",X"FF",X"C3",X"C1",X"01",X"CD",X"16",X"90",
		X"C3",X"ED",X"03",X"C3",X"29",X"90",X"21",X"3F",X"4C",X"C3",X"65",X"80",X"3A",X"2D",X"4C",X"CB",
		X"47",X"21",X"00",X"00",X"C8",X"21",X"96",X"13",X"C9",X"CD",X"30",X"91",X"CD",X"16",X"90",X"21",
		X"46",X"43",X"11",X"56",X"90",X"06",X"18",X"CD",X"24",X"91",X"21",X"47",X"43",X"06",X"18",X"CD",
		X"24",X"91",X"3E",X"80",X"CD",X"66",X"91",X"01",X"0C",X"91",X"16",X"06",X"CD",X"D0",X"03",X"3E",
		X"50",X"C3",X"77",X"91",X"B8",X"7F",X"5C",X"5D",X"60",X"61",X"64",X"65",X"68",X"69",X"6C",X"6D",
		X"70",X"71",X"40",X"40",X"74",X"75",X"70",X"71",X"78",X"79",X"7C",X"7D",X"86",X"87",X"5E",X"5F",
		X"62",X"63",X"66",X"67",X"6A",X"6B",X"6E",X"6F",X"72",X"73",X"40",X"40",X"76",X"77",X"72",X"73",
		X"7A",X"7B",X"7E",X"7F",X"88",X"89",X"06",X"40",X"43",X"4F",X"49",X"4E",X"40",X"40",X"43",X"52",
		X"45",X"44",X"49",X"54",X"FF",X"FF",X"FF",X"FF",X"FF",X"06",X"4F",X"4E",X"4C",X"59",X"40",X"4F",
		X"4E",X"45",X"40",X"50",X"4C",X"41",X"59",X"45",X"52",X"FF",X"FF",X"FF",X"FF",X"FF",X"06",X"42",
		X"4F",X"4E",X"55",X"53",X"40",X"50",X"4C",X"41",X"59",X"45",X"52",X"40",X"40",X"30",X"30",X"30",
		X"30",X"FF",X"FF",X"FF",X"FF",X"13",X"4E",X"55",X"4D",X"42",X"45",X"52",X"40",X"43",X"52",X"41",
		X"53",X"48",X"40",X"56",X"84",X"85",X"40",X"31",X"3D",X"30",X"FF",X"FF",X"FF",X"13",X"43",X"4F",
		X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"40",X"31",X"39",X"38",X"33",X"3D",X"36",X"3D",X"FF",
		X"FF",X"FF",X"1C",X"42",X"59",X"40",X"48",X"41",X"4E",X"53",X"48",X"49",X"4E",X"40",X"47",X"4F",
		X"52",X"41",X"4B",X"55",X"40",X"26",X"50",X"45",X"4E",X"49",X"26",X"FF",X"86",X"90",X"ED",X"42",
		X"99",X"90",X"EF",X"42",X"AE",X"90",X"F2",X"42",X"C5",X"90",X"7C",X"43",X"DD",X"90",X"9D",X"43",
		X"F2",X"90",X"9E",X"43",X"1A",X"77",X"E7",X"13",X"3E",X"03",X"CD",X"C1",X"01",X"10",X"F5",X"C9",
		X"CD",X"6E",X"91",X"21",X"00",X"44",X"01",X"04",X"00",X"3E",X"0D",X"CF",X"C9",X"06",X"20",X"21",
		X"46",X"47",X"3E",X"09",X"CD",X"4F",X"91",X"3E",X"0D",X"CD",X"4F",X"91",X"10",X"F1",X"C9",X"E5",
		X"C5",X"0E",X"02",X"E5",X"06",X"18",X"77",X"E7",X"10",X"FC",X"E1",X"23",X"0D",X"20",X"F4",X"C1",
		X"E1",X"3E",X"05",X"C3",X"C1",X"01",X"CD",X"3D",X"91",X"3E",X"40",X"C3",X"C1",X"01",X"21",X"00",
		X"00",X"22",X"3A",X"4C",X"C3",X"00",X"01",X"21",X"06",X"E8",X"22",X"30",X"4C",X"22",X"32",X"4C",
		X"22",X"34",X"4C",X"22",X"36",X"4C",X"DD",X"21",X"C0",X"4C",X"DD",X"36",X"00",X"53",X"DD",X"36",
		X"02",X"A5",X"DD",X"36",X"04",X"FF",X"AF",X"00",X"00",X"00",X"3E",X"03",X"32",X"C8",X"4C",X"DD",
		X"21",X"C0",X"4C",X"06",X"03",X"C5",X"CD",X"B9",X"91",X"C1",X"DD",X"23",X"DD",X"23",X"10",X"F5",
		X"3A",X"C8",X"4C",X"A7",X"20",X"E9",X"C3",X"74",X"92",X"3E",X"01",X"CD",X"C1",X"01",X"DD",X"7E",
		X"01",X"A7",X"28",X"07",X"3D",X"DD",X"77",X"01",X"C3",X"23",X"92",X"DD",X"7E",X"00",X"A7",X"28",
		X"05",X"3D",X"DD",X"77",X"00",X"C9",X"CD",X"5F",X"92",X"3E",X"08",X"DD",X"77",X"01",X"DD",X"E5",
		X"E1",X"7D",X"D6",X"90",X"6F",X"00",X"7D",X"FE",X"30",X"28",X"20",X"FE",X"32",X"28",X"23",X"7E",
		X"FE",X"CE",X"20",X"07",X"CD",X"1D",X"92",X"23",X"C3",X"67",X"92",X"FE",X"FE",X"D8",X"DD",X"7E",
		X"09",X"CB",X"E7",X"DD",X"77",X"09",X"21",X"C8",X"4C",X"35",X"C9",X"7E",X"FE",X"BE",X"20",X"EB",
		X"18",X"E2",X"7E",X"FE",X"AE",X"20",X"E4",X"CD",X"1D",X"92",X"23",X"18",X"22",X"47",X"23",X"4E",
		X"C3",X"13",X"07",X"DD",X"E5",X"E1",X"7D",X"D6",X"90",X"6F",X"34",X"CD",X"42",X"92",X"FE",X"04",
		X"78",X"00",X"38",X"02",X"79",X"00",X"DD",X"E5",X"E1",X"11",X"32",X"03",X"19",X"77",X"C9",X"C3",
		X"70",X"92",X"7D",X"FE",X"30",X"28",X"0C",X"FE",X"32",X"28",X"0E",X"06",X"10",X"0E",X"14",X"DD",
		X"7E",X"01",X"C9",X"06",X"18",X"0E",X"1C",X"18",X"F6",X"06",X"70",X"0E",X"74",X"18",X"F0",X"DD",
		X"7E",X"09",X"CB",X"67",X"C8",X"E1",X"C9",X"36",X"01",X"11",X"00",X"04",X"19",X"36",X"06",X"C9",
		X"36",X"01",X"18",X"F5",X"3E",X"88",X"32",X"F6",X"4F",X"21",X"E6",X"00",X"22",X"34",X"4C",X"21",
		X"80",X"43",X"36",X"FE",X"E7",X"36",X"FF",X"0E",X"04",X"06",X"08",X"3A",X"35",X"4C",X"3D",X"32",
		X"35",X"4C",X"3E",X"05",X"CD",X"C1",X"01",X"10",X"F2",X"C5",X"2A",X"34",X"4C",X"CD",X"11",X"07",
		X"36",X"FE",X"E7",X"36",X"FF",X"C1",X"0D",X"20",X"E0",X"21",X"E6",X"00",X"22",X"34",X"4C",X"21",
		X"2C",X"0E",X"22",X"F6",X"4F",X"06",X"18",X"3A",X"35",X"4C",X"3D",X"32",X"35",X"4C",X"3E",X"01",
		X"CD",X"C1",X"01",X"78",X"E6",X"0F",X"FE",X"0B",X"0E",X"30",X"30",X"08",X"FE",X"06",X"0E",X"34",
		X"30",X"02",X"0E",X"2C",X"79",X"32",X"F6",X"4F",X"10",X"DD",X"3E",X"0F",X"CD",X"C1",X"01",X"18",
		X"21",X"3E",X"20",X"32",X"F6",X"4F",X"06",X"0A",X"3A",X"34",X"4C",X"3D",X"32",X"34",X"4C",X"3E",
		X"02",X"CD",X"C1",X"01",X"CB",X"50",X"3E",X"20",X"20",X"02",X"3E",X"24",X"32",X"F6",X"4F",X"10",
		X"E7",X"C9",X"CD",X"E1",X"92",X"3E",X"20",X"32",X"F6",X"4F",X"3E",X"20",X"CD",X"C1",X"01",X"3E",
		X"24",X"CD",X"9F",X"93",X"21",X"CE",X"E8",X"22",X"30",X"4C",X"21",X"3C",X"06",X"22",X"F2",X"4F",
		X"06",X"10",X"CD",X"7D",X"93",X"06",X"48",X"CD",X"8A",X"93",X"2A",X"30",X"4C",X"CD",X"11",X"07",
		X"23",X"36",X"01",X"3E",X"30",X"CD",X"C1",X"01",X"06",X"10",X"CD",X"A8",X"93",X"21",X"BE",X"E8",
		X"22",X"30",X"4C",X"06",X"30",X"CD",X"7D",X"93",X"06",X"48",X"CD",X"8A",X"93",X"2A",X"30",X"4C",
		X"CD",X"11",X"07",X"23",X"36",X"01",X"06",X"10",X"CD",X"B1",X"93",X"3E",X"20",X"32",X"F6",X"4F",
		X"21",X"AE",X"E8",X"22",X"30",X"4C",X"21",X"3C",X"06",X"22",X"F2",X"4F",X"06",X"58",X"CD",X"7D",
		X"93",X"06",X"70",X"CD",X"8A",X"93",X"3E",X"80",X"CD",X"C1",X"01",X"18",X"3D",X"3A",X"30",X"4C",
		X"3D",X"32",X"30",X"4C",X"CD",X"97",X"93",X"10",X"F4",X"C9",X"3A",X"31",X"4C",X"3D",X"32",X"31",
		X"4C",X"CD",X"97",X"93",X"10",X"F4",X"C9",X"C5",X"06",X"00",X"CD",X"45",X"35",X"C1",X"C9",X"32",
		X"F6",X"4F",X"3E",X"40",X"32",X"24",X"43",X"C9",X"CD",X"E8",X"92",X"3E",X"40",X"32",X"E4",X"42",
		X"C9",X"CD",X"E8",X"92",X"3E",X"40",X"32",X"A4",X"42",X"C9",X"2A",X"30",X"4C",X"CD",X"11",X"07",
		X"23",X"36",X"01",X"3E",X"80",X"CD",X"C1",X"01",X"3E",X"22",X"32",X"F6",X"4F",X"06",X"2F",X"18",
		X"1A",X"3A",X"34",X"4C",X"3C",X"32",X"34",X"4C",X"3E",X"02",X"CD",X"C1",X"01",X"CB",X"50",X"3E",
		X"26",X"20",X"02",X"3E",X"22",X"32",X"F6",X"4F",X"10",X"E7",X"C9",X"CD",X"D1",X"93",X"3E",X"20",
		X"32",X"F6",X"4F",X"06",X"10",X"3A",X"35",X"4C",X"3D",X"32",X"35",X"4C",X"3E",X"01",X"CD",X"C1",
		X"01",X"10",X"F2",X"3E",X"30",X"CD",X"C1",X"01",X"3E",X"24",X"32",X"F6",X"4F",X"21",X"D6",X"D0",
		X"22",X"30",X"4C",X"21",X"8C",X"0D",X"22",X"F2",X"4F",X"21",X"46",X"43",X"CD",X"4A",X"94",X"0E",
		X"0D",X"06",X"10",X"3A",X"30",X"4C",X"3D",X"32",X"30",X"4C",X"CD",X"97",X"93",X"10",X"F4",X"2A",
		X"30",X"4C",X"CD",X"56",X"94",X"CD",X"4A",X"94",X"0D",X"20",X"E6",X"3E",X"30",X"CD",X"C1",X"01",
		X"06",X"D8",X"CD",X"E8",X"92",X"3E",X"A0",X"C3",X"C1",X"01",X"36",X"40",X"E7",X"36",X"40",X"23",
		X"36",X"40",X"DF",X"36",X"40",X"C9",X"C5",X"CD",X"11",X"07",X"C1",X"C9",X"CD",X"ED",X"01",X"CD",
		X"FF",X"12",X"C9",X"3A",X"2D",X"4C",X"CB",X"47",X"C8",X"21",X"3C",X"4C",X"C3",X"EC",X"12",X"21",
		X"43",X"96",X"22",X"4C",X"4C",X"21",X"00",X"25",X"22",X"85",X"4C",X"21",X"83",X"94",X"3E",X"02",
		X"C3",X"85",X"20",X"00",X"00",X"0F",X"0C",X"0E",X"0E",X"0E",X"0C",X"0E",X"0E",X"6E",X"0E",X"0E",
		X"0E",X"0E",X"BE",X"0E",X"0E",X"0E",X"0C",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0C",X"0E",
		X"0E",X"0E",X"BB",X"00",X"00",X"0E",X"0A",X"00",X"00",X"00",X"0A",X"00",X"00",X"6F",X"0F",X"0F",
		X"0F",X"0F",X"AF",X"0F",X"0F",X"0F",X"0B",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"0B",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"7E",X"0E",X"0E",
		X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0B",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"0A",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"9A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0B",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"B8",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"D0",X"F0",X"F0",X"F9",X"F0",X"F0",
		X"F0",X"F0",X"FB",X"F0",X"F0",X"F0",X"B0",X"08",X"00",X"00",X"00",X"00",X"A8",X"00",X"00",X"00",
		X"00",X"00",X"B6",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"C9",X"E0",X"E0",X"EB",X"E0",X"E0",
		X"E0",X"E0",X"EB",X"E0",X"E0",X"E0",X"B0",X"07",X"00",X"00",X"00",X"00",X"A6",X"00",X"00",X"00",
		X"00",X"00",X"B6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BA",X"00",X"00",X"0B",X"00",X"00",
		X"00",X"00",X"0A",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"00",X"00",
		X"00",X"00",X"B6",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"A0",X"00",X"00",X"0A",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"B6",X"00",X"00",X"F0",X"F0",X"F0",X"FA",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"B0",X"06",X"00",X"00",X"09",X"90",X"00",X"00",X"B0",X"00",
		X"00",X"00",X"B6",X"00",X"00",X"E8",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"B0",X"07",X"00",X"00",X"0B",X"D0",X"F0",X"F0",X"B0",X"00",
		X"00",X"00",X"B6",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"0A",X"E0",X"E0",X"E0",X"B0",X"00",
		X"00",X"00",X"B6",X"00",X"00",X"07",X"90",X"00",X"00",X"00",X"B0",X"00",X"00",X"09",X"00",X"00",
		X"00",X"00",X"08",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",
		X"00",X"00",X"B6",X"00",X"00",X"00",X"D0",X"F0",X"F0",X"F0",X"D0",X"F0",X"F0",X"FB",X"F0",X"F0",
		X"F0",X"F0",X"F6",X"F0",X"F0",X"F0",X"D0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"D0",X"F0",
		X"F0",X"F0",X"B7",X"1E",X"81",X"43",X"09",X"C9",X"42",X"09",X"32",X"41",X"09",X"81",X"42",X"08",
		X"B3",X"42",X"08",X"6E",X"40",X"08",X"04",X"43",X"07",X"CE",X"42",X"07",X"86",X"40",X"07",X"A6",
		X"41",X"06",X"8E",X"43",X"06",X"56",X"43",X"06",X"41",X"43",X"05",X"C2",X"41",X"05",X"77",X"41",
		X"05",X"26",X"41",X"04",X"D2",X"41",X"04",X"5A",X"42",X"04",X"C6",X"42",X"03",X"D8",X"42",X"03",
		X"F8",X"40",X"03",X"C1",X"42",X"02",X"09",X"43",X"02",X"98",X"40",X"02",X"C6",X"40",X"01",X"26",
		X"42",X"01",X"8E",X"42",X"01",X"13",X"43",X"00",X"89",X"43",X"00",X"5A",X"41",X"00",X"09",X"09",
		X"08",X"08",X"07",X"07",X"06",X"06",X"05",X"05",X"21",X"BE",X"43",X"06",X"0A",X"11",X"9E",X"96",
		X"1A",X"77",X"E7",X"13",X"10",X"FA",X"C3",X"DE",X"1C",X"02",X"53",X"50",X"45",X"43",X"49",X"41",
		X"4C",X"40",X"40",X"40",X"40",X"40",X"40",X"FF",X"FF",X"FF",X"11",X"24",X"20",X"CD",X"17",X"20",
		X"11",X"B9",X"96",X"21",X"A4",X"41",X"C3",X"76",X"97",X"7E",X"FE",X"53",X"C2",X"30",X"25",X"E1",
		X"21",X"40",X"40",X"01",X"04",X"80",X"3E",X"40",X"CF",X"CD",X"51",X"97",X"21",X"89",X"42",X"11",
		X"BA",X"96",X"06",X"08",X"CD",X"B6",X"26",X"11",X"D5",X"23",X"06",X"05",X"CD",X"61",X"97",X"0E",
		X"33",X"CD",X"8E",X"97",X"06",X"0D",X"77",X"E7",X"3C",X"10",X"FB",X"0D",X"20",X"F3",X"3E",X"30",
		X"CD",X"10",X"1D",X"21",X"8C",X"42",X"11",X"6A",X"97",X"06",X"06",X"CD",X"B6",X"26",X"11",X"71",
		X"97",X"06",X"05",X"CD",X"B6",X"26",X"3E",X"55",X"CD",X"10",X"1D",X"21",X"7A",X"43",X"11",X"CF",
		X"23",X"CD",X"ED",X"01",X"11",X"69",X"97",X"21",X"BA",X"41",X"CD",X"ED",X"01",X"3E",X"99",X"32",
		X"7F",X"4C",X"3E",X"90",X"32",X"7E",X"4C",X"CD",X"D6",X"24",X"AF",X"32",X"FD",X"4C",X"C3",X"5B",
		X"24",X"21",X"06",X"9B",X"22",X"03",X"4C",X"21",X"00",X"9C",X"C3",X"9C",X"19",X"00",X"00",X"00",
		X"00",X"CD",X"B6",X"26",X"AF",X"3D",X"C9",X"10",X"1D",X"07",X"09",X"09",X"09",X"00",X"00",X"40",
		X"FF",X"50",X"4F",X"49",X"4E",X"54",X"CD",X"ED",X"01",X"21",X"44",X"43",X"11",X"82",X"97",X"C3",
		X"ED",X"01",X"06",X"09",X"09",X"08",X"08",X"07",X"07",X"06",X"06",X"05",X"05",X"FF",X"21",X"89",
		X"46",X"F5",X"3E",X"02",X"CD",X"10",X"1D",X"F1",X"C9",X"C2",X"24",X"27",X"E5",X"2B",X"56",X"C3",
		X"0F",X"27",X"00",X"00",X"00",X"00",X"CD",X"CB",X"9A",X"E5",X"21",X"B8",X"97",X"22",X"03",X"4C",
		X"21",X"F4",X"98",X"CD",X"9C",X"19",X"E1",X"C9",X"03",X"88",X"00",X"0C",X"0F",X"03",X"88",X"00",
		X"0C",X"0F",X"03",X"88",X"00",X"0C",X"0F",X"03",X"08",X"00",X"0C",X"0F",X"03",X"27",X"00",X"0C",
		X"0F",X"03",X"27",X"00",X"0C",X"0F",X"03",X"27",X"00",X"0C",X"0F",X"03",X"08",X"00",X"0C",X"0F",
		X"03",X"79",X"00",X"0C",X"0F",X"03",X"79",X"00",X"0C",X"0F",X"03",X"9A",X"00",X"0C",X"1F",X"03",
		X"79",X"00",X"0C",X"1F",X"03",X"56",X"00",X"0C",X"1F",X"03",X"88",X"00",X"0C",X"0F",X"03",X"88",
		X"00",X"0C",X"0F",X"03",X"88",X"00",X"0C",X"0F",X"03",X"08",X"00",X"0C",X"0F",X"03",X"27",X"00",
		X"0C",X"0F",X"03",X"27",X"00",X"0C",X"0F",X"03",X"27",X"00",X"0C",X"0F",X"03",X"08",X"00",X"0C",
		X"0F",X"03",X"79",X"00",X"0C",X"0F",X"03",X"79",X"00",X"0C",X"0F",X"03",X"79",X"00",X"0C",X"0F",
		X"03",X"9A",X"00",X"0C",X"0F",X"03",X"79",X"00",X"1C",X"1F",X"03",X"79",X"00",X"0C",X"0F",X"03",
		X"9A",X"00",X"0C",X"0F",X"03",X"4B",X"00",X"1C",X"1F",X"03",X"4B",X"00",X"0C",X"0F",X"03",X"4B",
		X"00",X"0C",X"07",X"03",X"4B",X"00",X"0C",X"07",X"03",X"CC",X"00",X"1C",X"1F",X"03",X"CC",X"00",
		X"0C",X"0F",X"03",X"9A",X"00",X"0C",X"07",X"03",X"4B",X"00",X"0C",X"07",X"03",X"CC",X"00",X"1C",
		X"1F",X"03",X"CC",X"00",X"0C",X"07",X"03",X"CC",X"00",X"0C",X"07",X"03",X"CC",X"00",X"0C",X"07",
		X"03",X"4B",X"00",X"0C",X"07",X"03",X"4B",X"00",X"0C",X"1F",X"03",X"27",X"00",X"0C",X"0F",X"03",
		X"88",X"00",X"0C",X"0F",X"03",X"79",X"00",X"0C",X"07",X"03",X"79",X"00",X"0C",X"0F",X"03",X"79",
		X"00",X"0C",X"07",X"03",X"79",X"00",X"0C",X"07",X"03",X"79",X"00",X"0C",X"0F",X"03",X"79",X"00",
		X"0C",X"07",X"03",X"9A",X"00",X"0C",X"07",X"03",X"79",X"00",X"0C",X"07",X"03",X"79",X"00",X"0C",
		X"07",X"03",X"9A",X"00",X"0C",X"07",X"03",X"79",X"00",X"1C",X"1F",X"03",X"88",X"00",X"0C",X"0F",
		X"03",X"88",X"00",X"0C",X"0F",X"03",X"79",X"00",X"0C",X"07",X"03",X"88",X"00",X"0C",X"07",X"03",
		X"08",X"00",X"0C",X"0F",X"03",X"88",X"00",X"1C",X"0F",X"03",X"88",X"00",X"0C",X"0F",X"03",X"00",
		X"00",X"0A",X"20",X"10",X"04",X"22",X"00",X"0C",X"0F",X"06",X"88",X"00",X"08",X"07",X"06",X"9A",
		X"00",X"08",X"07",X"04",X"22",X"00",X"0C",X"0F",X"04",X"02",X"00",X"0C",X"0F",X"04",X"C1",X"00",
		X"0C",X"0F",X"06",X"88",X"00",X"08",X"07",X"06",X"9A",X"00",X"08",X"07",X"04",X"C1",X"00",X"0C",
		X"0F",X"04",X"22",X"00",X"0C",X"0F",X"04",X"62",X"00",X"0C",X"0F",X"06",X"88",X"00",X"08",X"07",
		X"06",X"4B",X"00",X"08",X"07",X"04",X"62",X"00",X"0C",X"07",X"06",X"2E",X"00",X"08",X"07",X"06",
		X"88",X"00",X"08",X"07",X"06",X"4B",X"00",X"08",X"07",X"04",X"33",X"00",X"0C",X"0F",X"06",X"79",
		X"00",X"08",X"07",X"06",X"4B",X"00",X"08",X"07",X"04",X"33",X"00",X"0C",X"07",X"04",X"D2",X"00",
		X"0C",X"07",X"04",X"B2",X"00",X"0C",X"07",X"04",X"62",X"00",X"0C",X"07",X"04",X"22",X"00",X"0C",
		X"0F",X"06",X"88",X"00",X"08",X"07",X"06",X"9A",X"00",X"08",X"07",X"04",X"22",X"00",X"0C",X"0F",
		X"04",X"02",X"00",X"0C",X"0F",X"04",X"C1",X"00",X"0C",X"0F",X"06",X"88",X"00",X"08",X"07",X"06",
		X"9A",X"00",X"08",X"07",X"04",X"C1",X"00",X"0C",X"0F",X"04",X"22",X"00",X"0C",X"0F",X"04",X"62",
		X"00",X"0C",X"0F",X"06",X"88",X"00",X"08",X"07",X"06",X"4B",X"00",X"08",X"07",X"04",X"62",X"00",
		X"0C",X"07",X"06",X"2E",X"00",X"08",X"07",X"06",X"88",X"00",X"08",X"07",X"06",X"4B",X"00",X"08",
		X"07",X"04",X"33",X"00",X"0C",X"0F",X"06",X"79",X"00",X"08",X"07",X"06",X"4B",X"00",X"08",X"07",
		X"04",X"62",X"00",X"0C",X"0F",X"04",X"B2",X"00",X"0C",X"0F",X"04",X"D2",X"00",X"0C",X"0F",X"06",
		X"88",X"00",X"08",X"07",X"06",X"4B",X"00",X"08",X"07",X"04",X"D2",X"00",X"0C",X"07",X"06",X"2E",
		X"00",X"08",X"07",X"06",X"88",X"00",X"08",X"07",X"06",X"4B",X"00",X"08",X"07",X"04",X"33",X"00",
		X"0C",X"0F",X"06",X"79",X"00",X"08",X"07",X"06",X"4B",X"00",X"08",X"07",X"04",X"33",X"00",X"0C",
		X"07",X"06",X"FF",X"00",X"08",X"07",X"06",X"79",X"00",X"08",X"07",X"06",X"4B",X"00",X"08",X"07",
		X"04",X"22",X"00",X"0C",X"0F",X"06",X"88",X"00",X"08",X"07",X"06",X"9A",X"00",X"08",X"07",X"04",
		X"B2",X"00",X"0C",X"0F",X"04",X"22",X"00",X"0C",X"0F",X"04",X"C1",X"00",X"0C",X"0F",X"06",X"88",
		X"00",X"08",X"07",X"06",X"9A",X"00",X"08",X"07",X"04",X"C1",X"00",X"0C",X"0F",X"04",X"22",X"00",
		X"0C",X"0F",X"04",X"62",X"00",X"0C",X"0F",X"06",X"88",X"00",X"08",X"07",X"06",X"4B",X"00",X"08",
		X"07",X"04",X"62",X"00",X"0C",X"07",X"06",X"2E",X"00",X"08",X"07",X"06",X"88",X"00",X"08",X"07",
		X"06",X"4B",X"00",X"08",X"07",X"04",X"33",X"00",X"0C",X"0F",X"06",X"79",X"00",X"08",X"07",X"06",
		X"4B",X"00",X"08",X"07",X"04",X"33",X"00",X"0C",X"07",X"06",X"FF",X"00",X"08",X"07",X"06",X"79",
		X"00",X"08",X"07",X"06",X"4B",X"00",X"08",X"07",X"04",X"22",X"00",X"0C",X"0F",X"06",X"88",X"00",
		X"08",X"07",X"06",X"9A",X"00",X"08",X"07",X"04",X"33",X"00",X"0C",X"07",X"06",X"FF",X"00",X"08",
		X"07",X"06",X"79",X"00",X"08",X"07",X"06",X"4B",X"00",X"08",X"07",X"06",X"44",X"00",X"18",X"0F",
		X"06",X"44",X"00",X"08",X"0F",X"04",X"00",X"00",X"08",X"20",X"10",X"22",X"00",X"4D",X"3E",X"80",
		X"CD",X"10",X"1D",X"E5",X"CD",X"DC",X"25",X"E1",X"3E",X"80",X"C3",X"10",X"1D",X"3A",X"40",X"4C",
		X"3D",X"E6",X"07",X"C9",X"32",X"81",X"4C",X"AF",X"32",X"89",X"4C",X"C9",X"05",X"A0",X"00",X"0F",
		X"0F",X"10",X"21",X"00",X"9B",X"22",X"0B",X"4C",X"AF",X"32",X"02",X"4C",X"21",X"BE",X"4C",X"C9",
		X"05",X"27",X"00",X"1F",X"8F",X"10",X"07",X"C4",X"00",X"0F",X"07",X"07",X"0C",X"00",X"0F",X"07",
		X"07",X"9A",X"00",X"0F",X"07",X"07",X"0C",X"00",X"0F",X"07",X"07",X"2E",X"00",X"0F",X"07",X"07",
		X"0C",X"00",X"0F",X"07",X"07",X"9A",X"00",X"0F",X"07",X"07",X"0C",X"00",X"0F",X"07",X"07",X"84",
		X"00",X"0F",X"07",X"07",X"9A",X"00",X"0F",X"07",X"07",X"9A",X"00",X"0F",X"07",X"07",X"9A",X"00",
		X"0F",X"07",X"07",X"2E",X"00",X"0F",X"07",X"07",X"9A",X"00",X"0F",X"07",X"07",X"9A",X"00",X"0F",
		X"07",X"07",X"9A",X"00",X"0F",X"07",X"07",X"44",X"00",X"0F",X"07",X"07",X"9A",X"00",X"0F",X"07",
		X"07",X"9A",X"00",X"0F",X"07",X"07",X"9A",X"00",X"0F",X"07",X"07",X"2E",X"00",X"0F",X"07",X"07",
		X"9A",X"00",X"0F",X"07",X"07",X"9A",X"00",X"0F",X"07",X"07",X"9A",X"00",X"0F",X"07",X"07",X"04",
		X"00",X"0F",X"07",X"07",X"79",X"00",X"0F",X"07",X"07",X"9A",X"00",X"0F",X"07",X"07",X"79",X"00",
		X"0F",X"07",X"07",X"2E",X"00",X"0F",X"07",X"07",X"79",X"00",X"0F",X"07",X"07",X"9A",X"00",X"0F",
		X"07",X"07",X"79",X"00",X"0F",X"07",X"07",X"C1",X"00",X"0F",X"07",X"07",X"F8",X"00",X"0F",X"07",
		X"07",X"9A",X"00",X"0F",X"07",X"07",X"F8",X"00",X"0F",X"07",X"07",X"2E",X"00",X"0F",X"07",X"07",
		X"2E",X"00",X"0F",X"07",X"07",X"2E",X"00",X"0F",X"07",X"07",X"2E",X"00",X"0F",X"07",X"10",X"32",
		X"3F",X"4C",X"32",X"81",X"4C",X"C9",X"CD",X"99",X"36",X"C3",X"ED",X"13",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"07",X"62",X"00",X"1F",X"1F",X"07",X"62",X"00",X"0F",X"1F",X"07",X"42",X"00",X"1F",X"1F",X"07",
		X"42",X"00",X"0F",X"1F",X"07",X"22",X"00",X"1F",X"1F",X"07",X"22",X"00",X"0F",X"1F",X"07",X"02",
		X"00",X"1F",X"1F",X"07",X"02",X"00",X"0F",X"1F",X"07",X"C1",X"00",X"1F",X"1F",X"07",X"C1",X"00",
		X"0F",X"1F",X"10",X"02",X"00",X"0F",X"1F",X"10",X"02",X"00",X"0F",X"1F",X"07",X"C1",X"00",X"0F",
		X"1F",X"07",X"C1",X"00",X"0F",X"1F",X"07",X"C1",X"00",X"0F",X"1F",X"07",X"C1",X"00",X"0F",X"1F",
		X"10",X"FF",X"14",X"E1",X"41",X"09",X"A5",X"42",X"09",X"45",X"41",X"00",X"B6",X"42",X"06",X"00",
		X"00",X"04",X"00",X"00",X"02",X"89",X"41",X"07",X"BB",X"42",X"08",X"8C",X"42",X"02",X"0C",X"42",
		X"06",X"6C",X"41",X"04",X"0E",X"43",X"03",X"51",X"42",X"01",X"00",X"00",X"03",X"76",X"42",X"00",
		X"97",X"41",X"05",X"F7",X"40",X"07",X"5B",X"42",X"05",X"3B",X"42",X"01",X"3B",X"41",X"08",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
