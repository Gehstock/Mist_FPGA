library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_SND_1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_SND_1 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"DD",X"7E",X"01",X"FD",X"77",X"01",X"DD",X"7E",X"02",X"FD",X"77",X"02",X"FD",X"36",X"05",X"00",
		X"C3",X"62",X"0F",X"04",X"0F",X"0F",X"00",X"21",X"13",X"10",X"11",X"A8",X"80",X"01",X"04",X"00",
		X"ED",X"B0",X"CD",X"7F",X"03",X"3E",X"01",X"CD",X"92",X"04",X"0E",X"0C",X"CD",X"3C",X"04",X"21",
		X"50",X"00",X"CD",X"5C",X"04",X"AF",X"C9",X"DD",X"21",X"13",X"10",X"FD",X"21",X"A8",X"80",X"FD",
		X"7E",X"03",X"FE",X"00",X"28",X"02",X"18",X"1B",X"CD",X"76",X"04",X"11",X"09",X"00",X"19",X"CD",
		X"5C",X"04",X"FD",X"35",X"00",X"20",X"0A",X"DD",X"7E",X"00",X"FD",X"77",X"00",X"FD",X"36",X"03",
		X"01",X"AF",X"C9",X"FD",X"35",X"01",X"20",X"F9",X"DD",X"7E",X"01",X"FD",X"77",X"01",X"CD",X"76",
		X"04",X"23",X"CD",X"5C",X"04",X"FD",X"35",X"02",X"28",X"02",X"AF",X"C9",X"3E",X"FF",X"C9",X"03",
		X"0A",X"0A",X"00",X"21",X"7F",X"10",X"11",X"B0",X"80",X"01",X"04",X"00",X"ED",X"B0",X"CD",X"7F",
		X"03",X"3E",X"01",X"CD",X"92",X"04",X"0E",X"0C",X"CD",X"3C",X"04",X"21",X"50",X"00",X"CD",X"5C",
		X"04",X"AF",X"C9",X"DD",X"21",X"7F",X"10",X"FD",X"21",X"B0",X"80",X"FD",X"7E",X"03",X"FE",X"00",
		X"28",X"02",X"18",X"1B",X"CD",X"76",X"04",X"11",X"09",X"00",X"19",X"CD",X"5C",X"04",X"FD",X"35",
		X"00",X"20",X"0A",X"DD",X"7E",X"00",X"FD",X"77",X"00",X"FD",X"36",X"03",X"01",X"AF",X"C9",X"FD",
		X"35",X"01",X"20",X"F9",X"DD",X"7E",X"01",X"FD",X"77",X"01",X"CD",X"76",X"04",X"23",X"CD",X"5C",
		X"04",X"FD",X"35",X"02",X"28",X"02",X"AF",X"C9",X"3E",X"FF",X"C9",X"3A",X"B6",X"80",X"B7",X"20",
		X"20",X"AF",X"CD",X"92",X"04",X"CD",X"7F",X"03",X"3E",X"00",X"32",X"67",X"80",X"CD",X"43",X"09",
		X"3E",X"11",X"21",X"02",X"80",X"77",X"23",X"36",X"00",X"23",X"3C",X"77",X"23",X"36",X"00",X"AF",
		X"C9",X"3E",X"FF",X"C9",X"DD",X"21",X"44",X"80",X"C3",X"86",X"07",X"3A",X"B6",X"80",X"B7",X"20",
		X"F0",X"AF",X"CD",X"92",X"04",X"CD",X"7F",X"03",X"AF",X"C9",X"DD",X"21",X"4C",X"80",X"C3",X"86",
		X"07",X"DD",X"21",X"54",X"80",X"C3",X"86",X"07",X"3E",X"01",X"32",X"B6",X"80",X"3E",X"10",X"CD",
		X"6D",X"00",X"3E",X"11",X"CD",X"6D",X"00",X"3E",X"12",X"CD",X"6D",X"00",X"AF",X"CD",X"92",X"04",
		X"CD",X"7F",X"03",X"3E",X"01",X"32",X"43",X"80",X"CD",X"3B",X"07",X"AF",X"C9",X"DD",X"21",X"20",
		X"80",X"C3",X"7E",X"05",X"DD",X"21",X"20",X"80",X"CD",X"7E",X"05",X"FE",X"FF",X"C0",X"AF",X"32",
		X"B6",X"80",X"3E",X"FF",X"C9",X"3E",X"01",X"32",X"B6",X"80",X"3E",X"10",X"CD",X"6D",X"00",X"3E",
		X"11",X"CD",X"6D",X"00",X"3E",X"12",X"CD",X"6D",X"00",X"AF",X"CD",X"92",X"04",X"CD",X"7F",X"03",
		X"AF",X"C9",X"DD",X"21",X"28",X"80",X"C3",X"7E",X"05",X"DD",X"21",X"28",X"80",X"C3",X"68",X"11",
		X"DD",X"21",X"30",X"80",X"C3",X"7E",X"05",X"DD",X"21",X"30",X"80",X"C3",X"68",X"11",X"3E",X"01",
		X"32",X"B6",X"80",X"3E",X"10",X"CD",X"6D",X"00",X"3E",X"11",X"CD",X"6D",X"00",X"3E",X"12",X"CD",
		X"6D",X"00",X"AF",X"CD",X"92",X"04",X"CD",X"7F",X"03",X"3E",X"02",X"32",X"43",X"80",X"CD",X"3B",
		X"07",X"AF",X"C9",X"3E",X"01",X"32",X"B6",X"80",X"3E",X"10",X"CD",X"6D",X"00",X"3E",X"11",X"CD",
		X"6D",X"00",X"3E",X"12",X"CD",X"6D",X"00",X"AF",X"CD",X"92",X"04",X"CD",X"7F",X"03",X"3E",X"03",
		X"32",X"43",X"80",X"CD",X"3B",X"07",X"AF",X"C9",X"3E",X"01",X"32",X"B6",X"80",X"3E",X"10",X"CD",
		X"6D",X"00",X"3E",X"11",X"CD",X"6D",X"00",X"3E",X"12",X"CD",X"6D",X"00",X"AF",X"CD",X"92",X"04",
		X"CD",X"7F",X"03",X"3E",X"04",X"32",X"43",X"80",X"CD",X"3B",X"07",X"AF",X"C9",X"3E",X"01",X"32",
		X"B6",X"80",X"3E",X"10",X"CD",X"6D",X"00",X"3E",X"11",X"CD",X"6D",X"00",X"3E",X"12",X"CD",X"6D",
		X"00",X"AF",X"CD",X"92",X"04",X"CD",X"7F",X"03",X"3E",X"05",X"32",X"43",X"80",X"CD",X"3B",X"07",
		X"AF",X"C9",X"3E",X"01",X"32",X"B6",X"80",X"3E",X"10",X"CD",X"6D",X"00",X"3E",X"11",X"CD",X"6D",
		X"00",X"3E",X"12",X"CD",X"6D",X"00",X"AF",X"CD",X"92",X"04",X"CD",X"7F",X"03",X"3E",X"06",X"32",
		X"43",X"80",X"CD",X"3B",X"07",X"AF",X"C9",X"DD",X"21",X"20",X"80",X"CD",X"7E",X"05",X"B7",X"C8",
		X"3E",X"01",X"C9",X"3E",X"01",X"32",X"B6",X"80",X"3E",X"10",X"CD",X"6D",X"00",X"3E",X"11",X"CD",
		X"6D",X"00",X"3E",X"12",X"CD",X"6D",X"00",X"AF",X"CD",X"92",X"04",X"CD",X"7F",X"03",X"AF",X"C9",
		X"DD",X"21",X"28",X"80",X"C3",X"6B",X"12",X"DD",X"21",X"30",X"80",X"C3",X"6B",X"12",X"3E",X"01",
		X"32",X"B6",X"80",X"3E",X"10",X"CD",X"6D",X"00",X"3E",X"11",X"CD",X"6D",X"00",X"3E",X"12",X"CD",
		X"6D",X"00",X"AF",X"CD",X"92",X"04",X"CD",X"7F",X"03",X"3E",X"07",X"32",X"43",X"80",X"CD",X"3B",
		X"07",X"AF",X"C9",X"3E",X"01",X"32",X"B6",X"80",X"3E",X"10",X"CD",X"6D",X"00",X"3E",X"11",X"CD",
		X"6D",X"00",X"3E",X"12",X"CD",X"6D",X"00",X"AF",X"CD",X"92",X"04",X"CD",X"7F",X"03",X"3E",X"08",
		X"32",X"43",X"80",X"CD",X"3B",X"07",X"AF",X"C9",X"3E",X"01",X"32",X"B6",X"80",X"3E",X"10",X"CD",
		X"6D",X"00",X"3E",X"11",X"CD",X"6D",X"00",X"3E",X"12",X"CD",X"6D",X"00",X"AF",X"CD",X"92",X"04",
		X"CD",X"7F",X"03",X"3E",X"09",X"32",X"43",X"80",X"CD",X"3B",X"07",X"AF",X"C9",X"49",X"13",X"65",
		X"13",X"81",X"13",X"9D",X"13",X"B9",X"13",X"D2",X"13",X"EE",X"13",X"29",X"14",X"64",X"14",X"9F",
		X"14",X"B6",X"14",X"C7",X"14",X"D8",X"14",X"10",X"15",X"48",X"15",X"80",X"15",X"AB",X"15",X"D6",
		X"15",X"01",X"16",X"2C",X"16",X"57",X"16",X"82",X"16",X"DA",X"16",X"27",X"17",X"6F",X"17",X"B7",
		X"17",X"09",X"18",X"5B",X"18",X"88",X"18",X"B5",X"18",X"1F",X"0D",X"3F",X"06",X"5F",X"09",X"4D",
		X"2F",X"2F",X"5F",X"08",X"2F",X"5F",X"07",X"2F",X"5F",X"06",X"2F",X"5F",X"05",X"2F",X"5F",X"04",
		X"2F",X"5F",X"03",X"2F",X"FF",X"1F",X"0D",X"3F",X"06",X"5F",X"09",X"4A",X"2B",X"2B",X"5F",X"08",
		X"2B",X"5F",X"07",X"2B",X"5F",X"06",X"2B",X"5F",X"05",X"2B",X"5F",X"04",X"2B",X"5F",X"03",X"2B",
		X"FF",X"1F",X"0D",X"3F",X"06",X"5F",X"09",X"46",X"26",X"26",X"5F",X"08",X"26",X"5F",X"07",X"26",
		X"5F",X"06",X"26",X"5F",X"05",X"26",X"5F",X"04",X"26",X"5F",X"03",X"26",X"FF",X"1F",X"0C",X"3F",
		X"0B",X"5F",X"09",X"70",X"90",X"72",X"70",X"6E",X"6D",X"6E",X"70",X"90",X"72",X"70",X"6E",X"6D",
		X"6E",X"70",X"70",X"8E",X"8D",X"8E",X"B0",X"B0",X"FF",X"1F",X"06",X"3F",X"0B",X"5F",X"08",X"79",
		X"99",X"7A",X"79",X"77",X"75",X"77",X"79",X"99",X"7A",X"79",X"77",X"75",X"77",X"B0",X"A0",X"A0",
		X"A0",X"FF",X"1F",X"06",X"3F",X"0B",X"5F",X"08",X"70",X"90",X"72",X"70",X"6E",X"6D",X"6E",X"70",
		X"90",X"72",X"70",X"6E",X"6D",X"6E",X"70",X"70",X"8E",X"8D",X"8E",X"B0",X"B0",X"FF",X"1F",X"0E",
		X"3F",X"0C",X"5F",X"09",X"93",X"70",X"73",X"70",X"60",X"95",X"71",X"75",X"71",X"60",X"93",X"31",
		X"31",X"31",X"31",X"91",X"60",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"B0",X"93",X"70",
		X"73",X"70",X"60",X"95",X"71",X"75",X"71",X"60",X"93",X"31",X"31",X"31",X"31",X"91",X"60",X"30",
		X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"B0",X"FF",X"1F",X"0E",X"3F",X"0C",X"5F",X"08",X"90",
		X"6C",X"70",X"6C",X"60",X"91",X"6E",X"71",X"6E",X"60",X"91",X"2E",X"2E",X"2E",X"2E",X"8E",X"60",
		X"2C",X"2C",X"2C",X"2C",X"2C",X"2C",X"2C",X"2C",X"AC",X"90",X"6C",X"70",X"6C",X"60",X"91",X"6E",
		X"71",X"6E",X"60",X"91",X"2E",X"2E",X"2E",X"2E",X"8E",X"60",X"2C",X"2C",X"2C",X"2C",X"2C",X"2C",
		X"2C",X"2C",X"AC",X"FF",X"1F",X"08",X"3F",X"0C",X"5F",X"08",X"30",X"30",X"30",X"30",X"30",X"30",
		X"30",X"30",X"B0",X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"B1",X"90",X"AE",X"90",X"8C",
		X"8E",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"B0",X"31",X"31",X"31",X"31",X"31",X"31",
		X"31",X"31",X"B1",X"90",X"AE",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"B0",X"FF",X"1F",
		X"0E",X"3F",X"0F",X"5F",X"09",X"AE",X"92",X"80",X"92",X"80",X"93",X"92",X"90",X"8E",X"8D",X"8B",
		X"89",X"8B",X"AD",X"B0",X"AE",X"FF",X"1F",X"08",X"3F",X"0F",X"5F",X"09",X"A2",X"A9",X"A9",X"A4",
		X"AB",X"AB",X"A1",X"A9",X"A4",X"A2",X"FF",X"1F",X"08",X"3F",X"0F",X"5F",X"09",X"AE",X"AE",X"AE",
		X"A0",X"B0",X"B0",X"A0",X"AD",X"B3",X"B2",X"FF",X"1F",X"0E",X"3F",X"0C",X"5F",X"09",X"29",X"29",
		X"29",X"29",X"29",X"20",X"26",X"26",X"26",X"26",X"20",X"29",X"29",X"29",X"29",X"20",X"2E",X"2E",
		X"2E",X"2E",X"2E",X"20",X"29",X"29",X"29",X"29",X"20",X"2E",X"2E",X"2E",X"2E",X"20",X"32",X"32",
		X"32",X"32",X"32",X"20",X"2E",X"2E",X"2E",X"2E",X"20",X"32",X"32",X"32",X"32",X"20",X"B5",X"FF",
		X"1F",X"0E",X"3F",X"0C",X"5F",X"09",X"26",X"26",X"26",X"26",X"26",X"20",X"22",X"22",X"22",X"22",
		X"20",X"26",X"26",X"26",X"26",X"20",X"29",X"29",X"29",X"29",X"29",X"20",X"26",X"26",X"26",X"26",
		X"20",X"29",X"29",X"29",X"29",X"20",X"2E",X"2E",X"2E",X"2E",X"2E",X"20",X"29",X"29",X"29",X"29",
		X"20",X"2E",X"2E",X"2E",X"2E",X"20",X"B2",X"FF",X"1F",X"08",X"3F",X"0C",X"5F",X"07",X"29",X"29",
		X"29",X"29",X"29",X"20",X"26",X"26",X"26",X"26",X"20",X"29",X"29",X"29",X"29",X"20",X"2E",X"2E",
		X"2E",X"2E",X"2E",X"20",X"29",X"29",X"29",X"29",X"20",X"2E",X"2E",X"2E",X"2E",X"20",X"32",X"32",
		X"32",X"32",X"32",X"20",X"2E",X"2E",X"2E",X"2E",X"20",X"32",X"32",X"32",X"32",X"20",X"B5",X"FF",
		X"1F",X"0E",X"3F",X"0C",X"5F",X"09",X"95",X"97",X"3A",X"39",X"38",X"37",X"36",X"35",X"34",X"33",
		X"32",X"31",X"30",X"2F",X"2E",X"2D",X"2C",X"2B",X"2A",X"29",X"28",X"27",X"26",X"25",X"24",X"23",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"A2",X"A0",X"FF",X"1F",X"0B",X"3F",X"0C",X"5F",
		X"09",X"9B",X"9D",X"3D",X"3C",X"3B",X"3A",X"39",X"38",X"37",X"36",X"35",X"34",X"33",X"32",X"31",
		X"30",X"2F",X"2E",X"2D",X"2C",X"2B",X"2A",X"29",X"28",X"27",X"26",X"25",X"25",X"25",X"25",X"25",
		X"25",X"25",X"25",X"A5",X"A0",X"FF",X"1F",X"0B",X"3F",X"0C",X"5F",X"09",X"9B",X"9D",X"39",X"38",
		X"37",X"36",X"35",X"34",X"33",X"32",X"31",X"30",X"2F",X"2E",X"2D",X"2C",X"2B",X"2A",X"29",X"28",
		X"27",X"26",X"25",X"24",X"23",X"22",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"A1",X"A0",
		X"FF",X"1F",X"0E",X"3F",X"0B",X"5F",X"07",X"89",X"89",X"8D",X"8D",X"8E",X"8E",X"90",X"90",X"89",
		X"89",X"8D",X"8D",X"8B",X"8B",X"84",X"84",X"89",X"89",X"8D",X"8D",X"8E",X"8E",X"8F",X"8F",X"1F",
		X"0B",X"90",X"92",X"90",X"92",X"B0",X"90",X"92",X"90",X"92",X"B0",X"FF",X"1F",X"05",X"3F",X"0B",
		X"5F",X"07",X"83",X"8F",X"87",X"8F",X"88",X"8F",X"8A",X"8F",X"83",X"8F",X"87",X"8F",X"85",X"91",
		X"8A",X"91",X"83",X"8F",X"87",X"8F",X"88",X"8F",X"8A",X"8F",X"1F",X"08",X"90",X"92",X"90",X"92",
		X"B0",X"90",X"92",X"90",X"92",X"B0",X"FF",X"1F",X"05",X"3F",X"0B",X"5F",X"07",X"83",X"93",X"80",
		X"93",X"80",X"93",X"80",X"93",X"80",X"93",X"80",X"93",X"80",X"94",X"80",X"94",X"80",X"93",X"80",
		X"93",X"80",X"93",X"80",X"93",X"1F",X"02",X"90",X"92",X"90",X"92",X"B0",X"90",X"92",X"90",X"92",
		X"B0",X"FF",X"1F",X"0E",X"3F",X"0E",X"5F",X"07",X"A4",X"A8",X"AB",X"84",X"A8",X"AB",X"84",X"A8",
		X"AB",X"A9",X"AD",X"AD",X"84",X"A9",X"AD",X"84",X"A9",X"AD",X"A4",X"A8",X"AB",X"84",X"A8",X"AB",
		X"84",X"A8",X"AB",X"A9",X"A9",X"89",X"A9",X"29",X"29",X"29",X"29",X"29",X"29",X"29",X"29",X"A9",
		X"A0",X"C0",X"AD",X"AE",X"AD",X"AB",X"A9",X"AB",X"A9",X"A6",X"AB",X"8B",X"8D",X"8B",X"8B",X"A9",
		X"A8",X"A6",X"A4",X"A0",X"AD",X"AE",X"AD",X"AB",X"A9",X"AB",X"A9",X"A6",X"8B",X"8B",X"8B",X"8D",
		X"8B",X"8B",X"A9",X"88",X"88",X"86",X"86",X"A4",X"A0",X"FF",X"1F",X"05",X"3F",X"0E",X"5F",X"06",
		X"AA",X"B1",X"B1",X"8A",X"B1",X"B1",X"8A",X"B1",X"B1",X"A3",X"AF",X"AF",X"83",X"AF",X"AF",X"83",
		X"AF",X"AF",X"AA",X"B1",X"B1",X"8A",X"B1",X"B1",X"8A",X"B1",X"B1",X"A3",X"A3",X"88",X"A8",X"83",
		X"A3",X"83",X"83",X"85",X"85",X"A6",X"A7",X"B1",X"AB",X"B1",X"A7",X"AF",X"AC",X"AF",X"A5",X"AF",
		X"AC",X"AF",X"AA",X"B1",X"A5",X"B1",X"A7",X"B1",X"AB",X"B1",X"A7",X"AF",X"AC",X"AF",X"A5",X"AF",
		X"AC",X"AF",X"AA",X"B1",X"A5",X"B1",X"FF",X"1F",X"08",X"3F",X"0E",X"5F",X"06",X"A4",X"AE",X"AE",
		X"80",X"AE",X"AE",X"80",X"AE",X"AE",X"A0",X"AD",X"AD",X"80",X"AD",X"AD",X"80",X"AD",X"AD",X"A4",
		X"AE",X"AE",X"80",X"AE",X"AE",X"80",X"AE",X"AE",X"AD",X"AD",X"8E",X"AE",X"8D",X"E0",X"A0",X"AD",
		X"A0",X"AD",X"A0",X"AD",X"A0",X"AD",X"A0",X"AF",X"A0",X"AF",X"A0",X"AE",X"A0",X"AE",X"A0",X"AD",
		X"A0",X"AD",X"A0",X"AD",X"A0",X"AD",X"A0",X"AF",X"A0",X"AF",X"A0",X"AE",X"A0",X"AE",X"FF",X"1F",
		X"0E",X"3F",X"0B",X"5F",X"06",X"90",X"91",X"92",X"91",X"90",X"91",X"B2",X"8D",X"8B",X"8B",X"8D",
		X"AB",X"A0",X"8B",X"8D",X"90",X"8B",X"8D",X"90",X"8B",X"8B",X"8C",X"8C",X"8C",X"8D",X"A9",X"A0",
		X"90",X"91",X"92",X"91",X"90",X"91",X"B2",X"8D",X"8B",X"8B",X"8D",X"AD",X"A0",X"8B",X"8D",X"90",
		X"8B",X"8D",X"90",X"8B",X"8B",X"6C",X"60",X"6C",X"60",X"6B",X"6B",X"60",X"29",X"29",X"29",X"29",
		X"89",X"64",X"66",X"60",X"64",X"86",X"FF",X"1F",X"05",X"3F",X"0B",X"5F",X"05",X"83",X"8F",X"87",
		X"8F",X"83",X"8F",X"87",X"8F",X"85",X"8F",X"8C",X"8F",X"85",X"8F",X"8C",X"8F",X"8A",X"91",X"85",
		X"91",X"8A",X"91",X"85",X"87",X"88",X"92",X"8C",X"92",X"83",X"8F",X"87",X"8F",X"83",X"8F",X"87",
		X"8F",X"83",X"8F",X"87",X"8F",X"85",X"8F",X"8C",X"8F",X"85",X"8F",X"8C",X"8F",X"8A",X"91",X"85",
		X"91",X"8A",X"91",X"85",X"87",X"1F",X"08",X"6C",X"60",X"6C",X"60",X"6B",X"6B",X"60",X"29",X"29",
		X"29",X"29",X"89",X"64",X"66",X"60",X"64",X"86",X"FF",X"1F",X"08",X"3F",X"0B",X"5F",X"05",X"89",
		X"8D",X"80",X"8D",X"80",X"8D",X"80",X"8D",X"80",X"8F",X"80",X"8F",X"80",X"8F",X"80",X"8F",X"80",
		X"8E",X"80",X"8E",X"80",X"8E",X"A0",X"80",X"8E",X"80",X"8E",X"80",X"8D",X"80",X"8D",X"89",X"8D",
		X"80",X"8D",X"80",X"8D",X"80",X"8D",X"80",X"8F",X"80",X"8F",X"80",X"8F",X"80",X"8F",X"80",X"8E",
		X"80",X"8E",X"80",X"8E",X"A0",X"1F",X"02",X"5F",X"07",X"6C",X"60",X"6C",X"60",X"6B",X"6B",X"60",
		X"29",X"29",X"29",X"29",X"89",X"64",X"66",X"60",X"64",X"86",X"FF",X"1F",X"0B",X"3F",X"0E",X"5F",
		X"07",X"6B",X"69",X"86",X"8E",X"8E",X"6B",X"69",X"86",X"8E",X"8E",X"6B",X"69",X"86",X"8E",X"8B",
		X"8E",X"89",X"8D",X"8D",X"6B",X"69",X"89",X"8D",X"8D",X"6B",X"69",X"89",X"8D",X"8D",X"6B",X"69",
		X"89",X"8D",X"8B",X"8D",X"8E",X"8E",X"8E",X"FF",X"1F",X"0B",X"3F",X"0E",X"5F",X"06",X"6B",X"69",
		X"80",X"86",X"86",X"6B",X"69",X"80",X"86",X"86",X"6B",X"69",X"80",X"86",X"80",X"86",X"80",X"87",
		X"87",X"6B",X"69",X"80",X"87",X"87",X"6B",X"69",X"80",X"87",X"87",X"6B",X"69",X"80",X"87",X"80",
		X"87",X"80",X"86",X"86",X"FF",X"1F",X"05",X"3F",X"0E",X"5F",X"06",X"80",X"2E",X"2E",X"2E",X"2E",
		X"2E",X"2E",X"2E",X"2E",X"AE",X"80",X"2E",X"2E",X"2E",X"2E",X"2E",X"2E",X"2E",X"2E",X"AE",X"80",
		X"AE",X"AB",X"29",X"29",X"29",X"29",X"29",X"29",X"29",X"29",X"A9",X"80",X"29",X"29",X"29",X"29",
		X"29",X"29",X"29",X"29",X"A9",X"80",X"29",X"29",X"29",X"29",X"29",X"29",X"29",X"29",X"A9",X"80",
		X"A9",X"AB",X"2E",X"2E",X"2E",X"2E",X"2E",X"2E",X"2E",X"2E",X"AE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
