library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity wacko_bg_bits_2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of wacko_bg_bits_2 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"08",X"20",X"2A",X"A8",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"80",X"A8",X"00",
		X"A0",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"02",X"00",X"0A",X"00",X"2A",X"00",X"AA",X"02",X"AA",X"0A",X"AA",X"2A",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A5",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"80",X"00",X"A8",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"0A",X"00",X"0A",X"00",X"2A",X"00",X"AA",X"00",X"AA",
		X"02",X"AA",X"0A",X"AA",X"8A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FD",X"55",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",
		X"00",X"A8",X"02",X"AA",X"00",X"AA",X"00",X"0A",X"00",X"0A",X"00",X"2A",X"00",X"AA",X"00",X"AA",
		X"02",X"AA",X"0A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A5",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"02",X"00",X"0A",X"00",X"2A",X"00",X"AA",X"02",X"AA",
		X"0A",X"AA",X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A5",
		X"AA",X"95",X"A9",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"F5",X"55",X"55",X"57",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"2A",X"00",X"AA",X"80",X"AA",X"A0",X"AA",X"A8",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"A9",X"AA",X"A5",X"AA",X"95",X"AA",X"55",X"A9",X"55",X"A5",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"7F",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"05",X"50",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"05",X"50",
		X"00",X"00",X"05",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"05",X"50",
		X"00",X"00",X"15",X"50",X"10",X"50",X"00",X"50",X"15",X"50",X"14",X"00",X"14",X"10",X"15",X"50",
		X"00",X"00",X"15",X"50",X"10",X"50",X"00",X"50",X"05",X"40",X"00",X"50",X"10",X"50",X"15",X"50",
		X"00",X"00",X"00",X"50",X"14",X"50",X"14",X"50",X"15",X"54",X"00",X"50",X"00",X"50",X"00",X"50",
		X"00",X"00",X"15",X"50",X"14",X"10",X"14",X"00",X"15",X"50",X"00",X"50",X"10",X"50",X"15",X"50",
		X"00",X"00",X"15",X"54",X"14",X"14",X"14",X"00",X"15",X"54",X"14",X"14",X"14",X"14",X"15",X"54",
		X"00",X"00",X"15",X"50",X"14",X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"00",X"50",
		X"00",X"00",X"15",X"54",X"14",X"14",X"14",X"14",X"05",X"50",X"14",X"14",X"14",X"14",X"15",X"54",
		X"00",X"00",X"15",X"54",X"14",X"14",X"14",X"14",X"15",X"54",X"00",X"14",X"14",X"14",X"15",X"54",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"80",X"A0",X"A2",X"A8",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"AA",X"A0",X"AA",X"80",X"AA",X"80",X"AA",X"A0",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"95",X"A9",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"F5",X"5F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"05",X"50",X"14",X"14",X"14",X"14",X"14",X"14",X"15",X"54",X"14",X"14",X"14",X"14",
		X"00",X"00",X"15",X"54",X"14",X"14",X"14",X"14",X"15",X"50",X"14",X"14",X"14",X"14",X"15",X"54",
		X"00",X"00",X"15",X"54",X"14",X"14",X"14",X"00",X"14",X"00",X"14",X"14",X"14",X"14",X"15",X"54",
		X"00",X"00",X"15",X"50",X"14",X"54",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"54",X"15",X"50",
		X"00",X"00",X"15",X"54",X"14",X"14",X"14",X"00",X"15",X"40",X"14",X"00",X"14",X"14",X"15",X"54",
		X"00",X"00",X"15",X"54",X"14",X"14",X"14",X"00",X"15",X"40",X"14",X"00",X"14",X"00",X"14",X"00",
		X"00",X"00",X"15",X"54",X"14",X"14",X"14",X"00",X"14",X"54",X"14",X"14",X"14",X"14",X"15",X"54",
		X"00",X"00",X"14",X"14",X"14",X"14",X"14",X"14",X"15",X"54",X"14",X"14",X"14",X"14",X"14",X"14",
		X"00",X"00",X"05",X"50",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"05",X"50",
		X"00",X"00",X"01",X"54",X"00",X"50",X"00",X"50",X"00",X"50",X"14",X"50",X"14",X"50",X"15",X"50",
		X"00",X"00",X"14",X"10",X"14",X"50",X"15",X"50",X"15",X"00",X"15",X"50",X"14",X"50",X"14",X"50",
		X"00",X"00",X"14",X"00",X"14",X"00",X"14",X"00",X"14",X"00",X"14",X"14",X"14",X"14",X"15",X"54",
		X"00",X"00",X"54",X"54",X"55",X"54",X"51",X"14",X"51",X"14",X"50",X"14",X"50",X"14",X"50",X"14",
		X"00",X"00",X"50",X"14",X"54",X"14",X"55",X"14",X"55",X"54",X"51",X"54",X"50",X"54",X"50",X"14",
		X"00",X"00",X"15",X"54",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"15",X"54",
		X"00",X"00",X"15",X"54",X"14",X"14",X"14",X"14",X"15",X"54",X"14",X"00",X"14",X"00",X"14",X"00",
		X"00",X"00",X"55",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"51",X"50",X"51",X"54",X"55",X"54",
		X"00",X"00",X"15",X"54",X"14",X"14",X"14",X"14",X"15",X"50",X"14",X"14",X"14",X"14",X"14",X"14",
		X"00",X"00",X"15",X"54",X"14",X"14",X"14",X"00",X"15",X"54",X"00",X"14",X"14",X"14",X"15",X"54",
		X"00",X"00",X"15",X"54",X"15",X"54",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",
		X"00",X"00",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"15",X"54",
		X"00",X"00",X"14",X"04",X"14",X"04",X"14",X"04",X"14",X"14",X"14",X"50",X"15",X"40",X"15",X"00",
		X"00",X"00",X"50",X"14",X"50",X"14",X"50",X"14",X"51",X"14",X"51",X"14",X"55",X"54",X"54",X"54",
		X"00",X"00",X"50",X"14",X"54",X"54",X"15",X"50",X"05",X"40",X"15",X"50",X"54",X"54",X"50",X"14",
		X"00",X"00",X"14",X"14",X"14",X"14",X"15",X"54",X"05",X"50",X"01",X"40",X"01",X"40",X"01",X"40",
		X"00",X"00",X"15",X"54",X"14",X"14",X"00",X"50",X"01",X"40",X"05",X"00",X"14",X"14",X"15",X"54",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"01",X"AA",X"05",X"AA",X"15",
		X"AA",X"55",X"A9",X"55",X"A5",X"55",X"A5",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"F5",X"55",X"FD",X"55",X"FF",X"D5",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"05",X"50",X"05",X"54",X"15",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"F5",X"55",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"A9",
		X"0A",X"A9",X"0A",X"A5",X"02",X"A5",X"00",X"15",X"00",X"55",X"00",X"55",X"01",X"55",X"01",X"55",
		X"05",X"55",X"15",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"7F",X"55",X"5F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"54",X"01",X"54",X"05",X"54",X"05",
		X"55",X"05",X"55",X"15",X"55",X"15",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"57",X"FF",X"57",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"54",X"01",X"55",X"05",X"55",X"05",X"55",X"45",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"50",X"50",
		X"55",X"54",X"55",X"56",X"55",X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"FF",X"F5",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"0A",X"02",
		X"AA",X"8A",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"AA",X"A8",X"60",X"A0",X"50",X"20",X"50",X"00",
		X"54",X"00",X"55",X"00",X"55",X"40",X"55",X"50",X"55",X"54",X"55",X"54",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"40",X"00",X"40",X"00",X"50",X"00",X"55",X"00",X"55",X"40",X"55",X"54",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"7F",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"54",X"02",
		X"55",X"0A",X"55",X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"7F",X"57",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"02",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"0A",X"00",X"AA",
		X"02",X"AA",X"02",X"AA",X"0A",X"AA",X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"5A",X"AA",X"56",X"AA",X"55",X"AA",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"A0",X"0A",X"AA",X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"02",X"AA",
		X"0A",X"AA",X"0A",X"AA",X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A9",X"AA",X"A5",
		X"AA",X"95",X"AA",X"55",X"A9",X"55",X"A5",X"55",X"95",X"55",X"95",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"FD",X"55",X"F5",X"55",X"F5",X"55",X"FD",X"55",X"FF",X"FD",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"80",X"2A",X"A0",X"AA",X"A0",X"AA",X"A8",X"AA",X"A8",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"6A",X"A9",X"6A",X"A9",
		X"AA",X"A9",X"AA",X"A9",X"AA",X"AA",X"5A",X"AA",X"56",X"AA",X"56",X"AA",X"55",X"AA",X"55",X"AA",
		X"55",X"6A",X"55",X"56",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"2A",X"00",
		X"AA",X"80",X"AA",X"A8",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"A6",X"AA",X"A6",X"AA",X"96",X"AA",X"5A",X"AA",X"5A",X"A9",X"5A",X"65",X"5A",X"55",X"5A",
		X"55",X"56",X"55",X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"A5",X"56",X"AA",X"56",X"AA",X"AA",
		X"AA",X"AB",X"AA",X"BF",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"AA",X"A0",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A9",
		X"FF",X"D5",X"FF",X"55",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"D5",X"55",X"FD",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"5F",X"57",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"5F",X"55",X"FF",X"F5",X"FF",X"FD",X"FF",X"FF",X"FF",X"FF",
		X"F5",X"55",X"F5",X"55",X"FD",X"55",X"FF",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"D5",X"FD",X"55",X"FD",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"55",X"AA",X"55",X"AA",X"55",X"A9",X"55",X"A5",X"55",X"95",X"55",X"55",X"55",X"D5",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"0A",X"00",X"2A",
		X"A8",X"00",X"AA",X"A8",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A9",X"AA",X"A5",X"AA",X"95",
		X"00",X"15",X"00",X"55",X"00",X"55",X"01",X"55",X"05",X"55",X"15",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"A0",X"00",X"A8",X"00",
		X"00",X"00",X"00",X"00",X"A0",X"00",X"AA",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A9",X"6A",X"A9",X"55",X"A5",X"55",X"55",
		X"A0",X"00",X"A8",X"00",X"A8",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"80",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"6A",X"AA",X"56",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"6A",X"AA",X"5A",X"AA",
		X"56",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"6A",X"55",X"5A",X"55",X"56",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"28",X"00",X"AA",X"02",X"AA",X"0A",X"AA",X"8A",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"95",X"55",X"A5",X"55",X"A9",X"55",
		X"A9",X"55",X"A9",X"55",X"A9",X"55",X"A9",X"55",X"A5",X"55",X"A5",X"55",X"A5",X"55",X"A9",X"55",
		X"A6",X"AA",X"A9",X"AA",X"AA",X"6A",X"AA",X"9A",X"AA",X"96",X"AA",X"A5",X"AA",X"A5",X"AA",X"A5",
		X"AA",X"A9",X"AA",X"A9",X"AA",X"A9",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"A9",X"AA",X"A9",X"AA",X"A9",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"EA",X"AA",X"FA",X"AA",X"FA",X"AA",X"FA",X"AA",X"FE",X"BA",X"FF",X"FF",X"FF",X"FF",
		X"00",X"02",X"80",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"2A",X"80",X"AA",X"A0",X"AA",X"A8",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"FF",X"AA",X"BF",X"AA",X"AF",X"AA",X"AF",X"AA",X"AF",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",
		X"AA",X"AB",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"BF",X"AB",X"FF",X"BF",X"FF",X"AF",X"FF",X"AF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"AB",X"FF",X"AA",X"BF",X"AA",X"AF",X"AA",X"AF",X"AA",X"AB",X"AA",X"AB",X"AA",X"AB",
		X"AA",X"AB",X"AA",X"AB",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"AF",X"FF",X"AB",X"FE",X"AB",X"FA",X"AB",X"EA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"AA",X"BF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"FF",X"AF",X"FF",X"AF",X"FF",X"AB",X"FF",
		X"AA",X"FF",X"AA",X"FF",X"AA",X"FF",X"AA",X"FF",X"AA",X"FF",X"AB",X"FF",X"AB",X"FF",X"AB",X"FF",
		X"AA",X"BF",X"AA",X"AF",X"AA",X"AB",X"AA",X"AB",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"AA",X"FF",X"AA",X"FE",X"AA",X"FA",X"AA",X"FA",X"AA",X"FA",X"AA",X"FA",X"AA",
		X"EA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"EA",X"AA",X"AA",X"AA",
		X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FA",X"FF",X"FA",X"EA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"02",X"AA",X"0A",X"AA",X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FA",X"AA",X"EA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FE",X"FF",X"FA",X"FF",X"FA",X"FF",X"FA",X"FA",X"BA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"A0",X"CA",X"A0",X"CA",X"A0",X"2A",X"80",X"02",X"8E",X"02",X"A8",X"00",X"A0",X"C0",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FE",X"FF",X"FA",X"FF",X"FA",X"FF",X"FA",X"FF",X"EA",X"FF",X"EA",X"FF",X"AA",X"FF",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"05",X"50",X"14",X"14",X"11",X"44",X"11",X"04",X"11",X"04",X"11",X"44",X"14",X"14",X"05",X"50",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"00",X"FF",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"03",X"FF",X"03",X"FF",X"03",X"FF",X"03",X"FF",X"03",X"FF",X"03",X"FF",
		X"03",X"FF",X"03",X"FF",X"03",X"FF",X"03",X"FF",X"03",X"FF",X"03",X"FF",X"03",X"FF",X"03",X"FF",
		X"03",X"FF",X"03",X"FF",X"03",X"FF",X"03",X"FF",X"03",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"AA",X"56",X"AA",X"56",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"03",X"C0",X"03",X"C0",X"0F",X"C0",X"0F",
		X"C0",X"3F",X"C0",X"3F",X"C0",X"FF",X"C0",X"FF",X"C3",X"FF",X"C3",X"FF",X"CF",X"FF",X"CF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"56",X"AA",X"56",X"AA",X"56",X"AA",X"96",X"AA",X"96",X"AA",X"96",X"AA",X"56",X"AA",X"5A",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FC",X"FF",X"F0",X"FF",X"F0",X"FF",X"C0",X"FF",X"C0",X"FF",X"00",
		X"FF",X"00",X"FC",X"00",X"FC",X"00",X"F0",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"30",X"00",X"FC",X"00",X"FC",X"03",X"FC",X"03",X"FC",X"0F",X"FC",X"0F",X"FC",
		X"3F",X"FC",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"A6",X"AA",X"A6",X"AA",X"A5",X"AA",X"A5",X"AA",X"A5",X"6A",X"AF",X"6A",X"AF",X"FF",X"AB",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"FF",X"3F",X"FF",
		X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"0F",X"FF",X"0F",X"FF",X"00",X"00",X"00",X"00",
		X"A8",X"00",X"AA",X"00",X"AA",X"80",X"AA",X"A0",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"C0",X"03",X"C0",X"03",X"C0",X"0F",X"F0",X"0F",X"F0",X"3F",X"F0",X"3F",X"F0",X"FF",X"F0",X"FF",
		X"F3",X"FF",X"F3",X"FF",X"F3",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A5",X"AA",X"A9",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FF",X"FC",X"FF",X"F0",X"FF",X"F0",
		X"FF",X"C0",X"FF",X"C0",X"FF",X"00",X"FF",X"00",X"FC",X"00",X"F0",X"00",X"00",X"03",X"00",X"03",
		X"00",X"FF",X"03",X"FF",X"0F",X"FF",X"0F",X"FF",X"3F",X"FF",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"C0",X"FF",X"C0",X"FF",X"C0",X"FF",X"00",X"FC",X"00",X"FC",X"00",X"F0",X"03",X"F0",X"03",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"3F",X"FF",X"0F",X"FF",X"00",X"FF",X"00",X"3F",X"00",X"0F",X"00",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"2A",X"82",
		X"00",X"00",X"02",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"0F",X"FF",X"3F",X"FF",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FF",X"FC",X"FF",X"F0",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A9",X"AA",X"A5",X"AA",X"A5",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"F3",X"FF",X"C3",X"FF",X"03",X"FF",X"03",X"FF",X"03",X"FF",X"03",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"AA",X"55",X"AA",X"95",X"AA",X"96",X"AA",X"96",X"AA",X"96",X"AA",X"9A",X"AA",X"AA",X"AA",
		X"AA",X"A9",X"AA",X"A5",X"AA",X"95",X"AA",X"55",X"AA",X"56",X"A6",X"56",X"55",X"5A",X"5F",X"FA",
		X"00",X"00",X"00",X"02",X"00",X"0A",X"00",X"0A",X"00",X"2A",X"A0",X"AA",X"A2",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"FF",X"0F",X"FF",X"0F",X"FF",X"0F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",
		X"A0",X"0A",X"A0",X"3A",X"A0",X"0A",X"A8",X"2A",X"AB",X"0A",X"AC",X"0A",X"AC",X"0A",X"A0",X"0A",
		X"3F",X"FF",X"3F",X"FF",X"0F",X"FF",X"0F",X"FF",X"0F",X"FF",X"0F",X"FF",X"0F",X"FF",X"0F",X"FF",
		X"0F",X"FF",X"03",X"FF",X"03",X"FF",X"03",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"3F",X"00",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"F0",X"00",
		X"00",X"03",X"00",X"3F",X"03",X"FF",X"0F",X"FF",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"0A",X"00",X"2A",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"FF",X"0F",X"FF",X"03",X"FF",X"00",X"FF",
		X"00",X"2A",X"00",X"AA",X"02",X"AA",X"0A",X"AA",X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"6A",X"AA",X"56",X"AA",X"55",X"AA",X"55",X"6A",X"55",X"5A",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3F",X"FF",X"0F",X"FF",X"0F",X"FF",X"0F",X"FF",X"03",X"FF",X"00",X"FF",X"00",X"3F",X"00",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"0F",X"00",X"3F",
		X"00",X"02",X"00",X"0A",X"00",X"2A",X"00",X"AA",X"6A",X"AA",X"6A",X"AA",X"5A",X"AA",X"56",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"00",X"C0",X"00",X"F0",X"00",X"F0",X"00",X"FC",X"00",X"FC",X"00",X"FF",X"00",X"FF",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"00",X"FC",X"03",X"FF",
		X"54",X"00",X"55",X"00",X"55",X"40",X"55",X"50",X"55",X"54",X"55",X"54",X"55",X"55",X"55",X"55",
		X"C3",X"FF",X"F3",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"0F",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FC",X"3F",X"FC",X"0F",X"F0",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",
		X"03",X"F0",X"03",X"FC",X"0F",X"FF",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",
		X"FF",X"3F",X"FC",X"3F",X"FC",X"3F",X"F0",X"3F",X"F0",X"3F",X"C0",X"3F",X"00",X"3F",X"00",X"3F",
		X"FF",X"FF",X"FF",X"3F",X"FC",X"3F",X"FC",X"3F",X"30",X"3F",X"00",X"3F",X"00",X"3F",X"00",X"3F",
		X"FF",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FC",X"00",X"FC",X"00",X"FC",X"00",X"FC",X"00",X"FC",X"00",X"FC",X"00",X"FC",X"00",X"FC",X"00",
		X"FC",X"00",X"FC",X"00",X"FC",X"00",X"FC",X"00",X"FC",X"00",X"FC",X"03",X"FC",X"0F",X"FC",X"3F",
		X"FC",X"3F",X"FC",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"3F",X"FC",X"0F",X"FC",X"03",X"FC",X"00",X"FC",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"F0",X"00",X"FC",X"00",X"FF",X"00",X"FF",X"C0",X"FF",X"F0",X"FF",X"FC",X"FF",X"FC",X"FF",X"FF",
		X"D5",X"55",X"F5",X"55",X"FF",X"55",X"FF",X"55",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F0",X"00",X"C0",X"03",X"00",X"03",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"3F",X"00",X"3F",
		X"00",X"3F",X"00",X"3F",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"C0",X"FF",X"F0",X"FF",X"F0",X"FF",X"FC",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"3F",X"FF",X"0F",X"FC",X"03",X"F0",X"00",X"F0",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"56",X"AA",X"55",X"6A",X"55",X"5A",X"55",X"56",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"FF",
		X"C0",X"3F",X"C0",X"3F",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"FF",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FF",X"F0",X"FF",X"C0",
		X"FF",X"00",X"FF",X"00",X"FC",X"00",X"FC",X"00",X"FC",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"FF",X"00",X"C0",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FF",X"FC",X"FF",X"F0",X"FF",X"F0",X"FF",X"C0",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"03",X"FF",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"D5",X"55",X"F5",X"55",X"F5",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"5A",X"AA",X"56",X"AA",X"55",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"55",X"6A",X"55",X"6A",X"55",X"5A",X"55",X"5A",X"55",X"5A",X"55",X"5A",X"55",X"56",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"5D",X"55",X"5F",X"D7",X"57",X"FF",
		X"AA",X"AA",X"59",X"AA",X"55",X"6A",X"55",X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"5F",X"FD",X"7F",X"5F",X"FF",X"5F",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"6A",X"AA",X"5A",X"AA",X"56",X"AA",
		X"56",X"AA",X"56",X"AA",X"55",X"AA",X"55",X"6A",X"55",X"5A",X"55",X"56",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"55",X"6A",X"55",X"5A",X"55",X"5A",X"55",X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"57",X"55",X"5F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"A0",X"00",X"AA",X"00",X"AA",X"80",X"AA",X"A0",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"95",X"AA",X"A5",X"AA",X"A9",X"AA",X"A9",X"AA",X"A9",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"59",X"6A",X"55",X"5A",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"FD",X"55",X"FF",X"D5",
		X"00",X"0A",X"00",X"2A",X"00",X"AA",X"02",X"AA",X"0A",X"AA",X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"56",X"AA",X"5A",X"AA",X"5A",X"AA",X"6A",X"AA",X"6A",X"AA",X"6A",X"AA",X"5A",X"AA",X"5A",X"AA",
		X"5A",X"AA",X"5A",X"AA",X"56",X"AA",X"56",X"AA",X"96",X"AA",X"96",X"AA",X"96",X"AA",X"95",X"AA",
		X"A5",X"AA",X"A5",X"AA",X"A6",X"AA",X"96",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"6A",X"AA",X"6A",X"AA",X"5A",X"AA",X"5A",X"AA",X"55",X"5A",X"55",X"56",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"6A",X"A9",X"5A",X"AA",X"96",X"AA",X"A6",X"AA",X"A6",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"55",X"00",X"55",X"40",X"55",X"50",X"55",X"54",X"55",X"55",X"55",X"55",X"55",X"55",X"54",X"05",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"A5",X"AA",X"A9",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A9",X"AA",X"A9",X"AA",X"A5",
		X"AA",X"A5",X"AA",X"96",X"AA",X"5A",X"A9",X"6A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"6A",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",
		X"96",X"AA",X"96",X"AA",X"96",X"AA",X"56",X"AA",X"56",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"6A",
		X"55",X"AA",X"56",X"AA",X"56",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"6A",X"AA",
		X"AA",X"A5",X"AA",X"95",X"AA",X"95",X"AA",X"55",X"AA",X"55",X"A5",X"56",X"95",X"5A",X"55",X"AA",
		X"55",X"AA",X"5A",X"AA",X"6A",X"AA",X"AA",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"9A",X"AA",X"5A",X"A9",X"5A",X"A9",X"5A",X"AA",X"5A",X"AA",X"56",X"AA",X"96",
		X"AA",X"AA",X"AA",X"AB",X"AA",X"AF",X"AA",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"2A",X"A0",X"0A",X"A0",X"2A",X"A8",X"0A",
		X"95",X"AA",X"A5",X"AA",X"BF",X"AA",X"FF",X"AA",X"FE",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"A9",X"55",X"AA",X"55",X"AA",X"95",X"AA",X"A9",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"5A",X"AA",X"5A",X"AA",X"56",X"AA",X"56",X"AA",X"56",X"AA",X"56",X"AA",X"55",X"AA",X"95",X"AA",
		X"95",X"6A",X"A5",X"5A",X"AA",X"55",X"AA",X"95",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"6A",X"AA",X"6A",X"AA",X"6A",X"AA",X"56",X"AA",X"56",X"AA",X"5A",X"AA",X"6A",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"A9",X"AA",X"A5",X"EA",X"A7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",
		X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"A5",X"DA",X"A5",X"FF",X"F5",X"FF",X"FD",
		X"A9",X"55",X"A5",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"57",X"D5",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"AA",X"A0",X"AA",X"80",
		X"AA",X"00",X"AA",X"00",X"AA",X"02",X"AA",X"8A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AB",X"AA",X"AF",X"AA",X"BF",
		X"AB",X"FF",X"AA",X"FF",X"AA",X"BF",X"AA",X"BF",X"AA",X"AF",X"AA",X"AB",X"AA",X"AA",X"AA",X"AA",
		X"A8",X"0A",X"A0",X"02",X"80",X"02",X"80",X"00",X"00",X"00",X"00",X"08",X"00",X"08",X"00",X"28",
		X"08",X"28",X"08",X"28",X"0A",X"2A",X"2A",X"AA",X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AF",X"AA",X"FF",X"AF",X"FF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"2A",X"A0",X"0A",X"A0",X"0A",X"80",X"0A",X"00",X"02",X"00",
		X"00",X"00",X"0A",X"20",X"0A",X"A0",X"0A",X"A0",X"2A",X"A2",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AB",X"AB",X"FF",
		X"AA",X"AA",X"2A",X"A8",X"0A",X"A0",X"02",X"80",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"A0",X"02",X"A0",X"82",X"A0",X"A2",X"A8",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"82",X"82",
		X"85",X"56",X"A5",X"5A",X"AA",X"A8",X"8A",X"A0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"05",X"50",X"1A",X"68",X"6A",X"AA",X"5A",X"69",X"55",X"55",X"59",X"55",X"1A",X"94",X"05",X"50",
		X"01",X"40",X"06",X"A0",X"06",X"A0",X"05",X"50",X"29",X"68",X"C0",X"03",X"AA",X"AA",X"22",X"C8",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AF",X"AB",X"FF",X"AF",X"FF",X"BF",X"FF",
		X"A0",X"02",X"80",X"80",X"02",X"00",X"00",X"00",X"00",X"0B",X"C0",X"AA",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AB",X"AA",X"FF",X"AF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AF",X"AF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"AB",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AF",X"00",X"FF",X"F0",X"FF",X"01",X"FF",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"48",X"00",X"0F",X"08",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"42",X"80",X"00",X"0F",X"00",X"03",X"30",X"83",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"BF",X"3F",X"FF",X"00",X"03",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"00",X"A8",X"00",X"A0",X"00",X"A0",X"00",X"F0",X"00",X"FC",X"00",X"FF",X"FF",X"FF",X"FF",
		X"0A",X"AA",X"0A",X"AB",X"0F",X"FF",X"0F",X"FF",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"A0",X"AA",X"9F",X"AA",X"57",X"AA",X"55",X"A9",X"55",X"A9",X"55",X"A9",X"55",X"A5",X"55",
		X"AF",X"FF",X"AF",X"FF",X"AF",X"FF",X"BF",X"FF",X"BF",X"FF",X"BF",X"FF",X"BF",X"FF",X"BF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"2A",
		X"00",X"0A",X"3C",X"00",X"FF",X"00",X"FF",X"C0",X"FF",X"F5",X"5F",X"D5",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"A0",X"00",X"00",X"03",X"15",X"0F",X"55",X"7F",X"55",X"5D",X"5A",X"55",X"6A",X"55",X"6A",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"AB",X"FF",X"AF",X"FF",X"BF",X"BF",X"FF",X"AF",X"FF",X"AB",X"FF",X"AB",X"F7",X"FE",
		X"F5",X"FE",X"F5",X"FF",X"F5",X"EE",X"FD",X"EA",X"BF",X"EE",X"AA",X"FF",X"EA",X"BF",X"FA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"EA",X"AF",X"EA",X"AB",X"AA",X"AA",X"AA",X"AA",X"FA",X"AA",X"BA",X"AA",
		X"BA",X"AA",X"FE",X"AA",X"EE",X"AA",X"AE",X"AA",X"EE",X"A9",X"FE",X"A9",X"FA",X"AB",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"FA",X"AB",X"FE",X"FF",X"FE",X"FF",X"FA",X"FF",X"FA",X"FF",X"BA",X"FF",
		X"BF",X"FF",X"BA",X"FF",X"FA",X"FF",X"FF",X"BF",X"FA",X"BB",X"7A",X"FA",X"FB",X"EB",X"FF",X"AF",
		X"00",X"00",X"10",X"00",X"10",X"00",X"10",X"00",X"14",X"00",X"04",X"00",X"94",X"00",X"94",X"00",
		X"85",X"00",X"89",X"00",X"89",X"00",X"A9",X"00",X"A5",X"00",X"A4",X"00",X"A4",X"00",X"A4",X"02",
		X"A4",X"02",X"A4",X"02",X"94",X"02",X"90",X"02",X"90",X"02",X"94",X"0A",X"A4",X"0A",X"A4",X"0A",
		X"A4",X"0A",X"A4",X"0A",X"A5",X"0A",X"A9",X"2A",X"A9",X"2A",X"A9",X"2A",X"A8",X"AA",X"A8",X"AA",
		X"00",X"00",X"10",X"00",X"14",X"00",X"04",X"00",X"04",X"00",X"05",X"00",X"49",X"00",X"49",X"00",
		X"29",X"00",X"A9",X"00",X"A5",X"00",X"A4",X"00",X"A4",X"02",X"A4",X"02",X"A5",X"02",X"A9",X"02",
		X"A9",X"02",X"A9",X"0A",X"A9",X"0A",X"A5",X"0A",X"A4",X"0A",X"A4",X"0A",X"A4",X"0A",X"A4",X"0A",
		X"A9",X"0A",X"A9",X"0A",X"A9",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"50",X"00",X"14",X"00",X"04",X"00",X"04",X"02",
		X"05",X"02",X"61",X"02",X"61",X"02",X"A9",X"0A",X"A9",X"0A",X"A4",X"0A",X"A4",X"0A",X"A4",X"0A",
		X"A4",X"0A",X"A4",X"0A",X"A4",X"2A",X"A8",X"2A",X"A8",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"40",X"00",X"50",X"00",X"10",X"00",X"14",X"00",X"04",X"04",X"05",X"00",X"01",X"08",
		X"01",X"28",X"49",X"2A",X"48",X"2A",X"28",X"AA",X"A8",X"AA",X"A8",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"05",X"00",X"55",X"01",X"55",X"05",X"55",X"05",X"55",X"15",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
