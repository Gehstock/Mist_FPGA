library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity snd_prg is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of snd_prg is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"81",X"C7",X"0F",X"BC",X"77",X"F3",X"2F",X"23",X"E8",X"5D",X"85",X"A9",X"87",X"D8",X"40",X"D3",
		X"0B",X"49",X"8C",X"52",X"D1",X"88",X"1E",X"5A",X"A5",X"8D",X"5A",X"3E",X"05",X"8D",X"22",X"9C",
		X"43",X"D8",X"5D",X"14",X"D2",X"B6",X"D9",X"5B",X"22",X"D1",X"80",X"1E",X"5B",X"96",X"B8",X"6D",
		X"49",X"C4",X"8C",X"58",X"D4",X"3D",X"18",X"D5",X"C1",X"5D",X"31",X"E4",X"9D",X"48",X"81",X"8D",
		X"49",X"82",X"E5",X"B3",X"C2",X"1E",X"5A",X"82",X"D5",X"D8",X"5A",X"A6",X"C4",X"0D",X"23",X"E2",
		X"8A",X"7D",X"19",X"42",X"D9",X"5D",X"85",X"C9",X"58",X"C5",X"8D",X"59",X"A3",X"8E",X"59",X"81",
		X"98",X"10",X"93",X"F2",X"2E",X"3A",X"85",X"BB",X"69",X"B6",X"C2",X"2E",X"5B",X"01",X"89",X"C7",
		X"1D",X"13",X"E0",X"5C",X"10",X"1F",X"35",X"D0",X"3E",X"05",X"AC",X"49",X"94",X"A8",X"82",X"1C",
		X"97",X"D0",X"5C",X"20",X"B1",X"10",X"B9",X"61",X"F4",X"2D",X"21",X"D0",X"39",X"C5",X"0D",X"40",
		X"D2",X"3E",X"12",X"B3",X"C1",X"83",X"E3",X"0B",X"10",X"5D",X"95",X"C8",X"5C",X"95",X"2D",X"05",
		X"CA",X"35",X"DA",X"5B",X"A6",X"9B",X"6B",X"86",X"D2",X"3D",X"82",X"1E",X"13",X"1F",X"85",X"9B",
		X"5A",X"82",X"88",X"B7",X"BA",X"68",X"C3",X"1C",X"00",X"39",X"F5",X"8C",X"48",X"A0",X"28",X"B4",
		X"3F",X"85",X"C9",X"30",X"C5",X"BA",X"68",X"D4",X"2D",X"85",X"9D",X"15",X"D8",X"5A",X"09",X"4A",
		X"91",X"83",X"BA",X"7C",X"30",X"B2",X"A5",X"9A",X"87",X"AC",X"41",X"D0",X"5D",X"05",X"AC",X"25",
		X"BC",X"25",X"D9",X"5C",X"85",X"9C",X"34",X"D0",X"4B",X"A5",X"8D",X"50",X"D4",X"1D",X"14",X"D9",
		X"5A",X"94",X"A8",X"49",X"C3",X"1C",X"03",X"AB",X"42",X"BA",X"36",X"D8",X"31",X"CA",X"42",X"9C",
		X"38",X"C4",X"8A",X"29",X"08",X"97",X"9D",X"33",X"BC",X"34",X"CA",X"50",X"A0",X"92",X"0C",X"2A",
		X"23",X"D0",X"2A",X"B7",X"8B",X"14",X"AA",X"58",X"C1",X"4A",X"C3",X"3D",X"A5",X"8B",X"59",X"90",
		X"19",X"1C",X"23",X"D9",X"50",X"D1",X"5C",X"A5",X"9B",X"5A",X"01",X"90",X"89",X"38",X"A2",X"C2",
		X"4A",X"B9",X"71",X"F0",X"59",X"C2",X"2A",X"80",X"18",X"92",X"99",X"82",X"3C",X"B7",X"B5",X"A9",
		X"13",X"BB",X"51",X"C8",X"4A",X"80",X"81",X"00",X"C3",X"2D",X"82",X"2A",X"D2",X"5C",X"82",X"89",
		X"3B",X"B7",X"0C",X"28",X"92",X"08",X"A3",X"8F",X"32",X"CA",X"40",X"A8",X"4A",X"92",X"2E",X"05",
		X"CA",X"58",X"A0",X"29",X"B5",X"1D",X"95",X"1D",X"04",X"9D",X"25",X"C8",X"11",X"A1",X"89",X"3B",
		X"02",X"9A",X"20",X"05",X"F0",X"4B",X"92",X"1B",X"39",X"90",X"23",X"F9",X"69",X"B1",X"3A",X"95",
		X"A9",X"22",X"BD",X"50",X"B0",X"5C",X"95",X"A9",X"39",X"90",X"29",X"1B",X"97",X"1F",X"05",X"8C",
		X"01",X"1A",X"83",X"A8",X"18",X"95",X"C2",X"8A",X"4A",X"92",X"2B",X"93",X"3D",X"C4",X"2E",X"12",
		X"C0",X"28",X"A1",X"1B",X"69",X"B2",X"3B",X"A4",X"90",X"88",X"3B",X"C7",X"8B",X"16",X"BA",X"40",
		X"B0",X"39",X"B5",X"9A",X"30",X"D1",X"4B",X"93",X"0C",X"13",X"C8",X"48",X"C1",X"28",X"C1",X"4A",
		X"C4",X"2D",X"83",X"8A",X"84",X"8B",X"04",X"8C",X"12",X"98",X"A2",X"4C",X"95",X"9A",X"10",X"80",
		X"2B",X"02",X"98",X"08",X"99",X"58",X"E4",X"0B",X"06",X"BB",X"78",X"A9",X"50",X"C0",X"20",X"B1",
		X"00",X"99",X"79",X"C2",X"4C",X"83",X"9A",X"11",X"0C",X"12",X"9A",X"31",X"D1",X"2A",X"A2",X"1A",
		X"3B",X"96",X"8A",X"12",X"D8",X"24",X"D9",X"15",X"AB",X"48",X"92",X"9A",X"48",X"90",X"94",X"AA",
		X"59",X"90",X"10",X"A0",X"28",X"A8",X"68",X"F1",X"3B",X"A4",X"2B",X"93",X"98",X"8A",X"79",X"A2",
		X"00",X"AB",X"70",X"9A",X"32",X"F0",X"28",X"A2",X"0C",X"15",X"AB",X"40",X"A0",X"18",X"A1",X"3B",
		X"C3",X"5A",X"E3",X"19",X"B3",X"88",X"82",X"89",X"B3",X"7B",X"B4",X"18",X"D2",X"4C",X"94",X"0B",
		X"02",X"98",X"81",X"92",X"B8",X"7A",X"92",X"1E",X"23",X"E8",X"30",X"AA",X"33",X"CB",X"41",X"B0",
		X"18",X"2A",X"A2",X"18",X"B0",X"4A",X"85",X"AF",X"58",X"A1",X"2B",X"A4",X"2B",X"B4",X"19",X"A0",
		X"4A",X"A3",X"3F",X"03",X"AC",X"33",X"BC",X"32",X"BA",X"15",X"9B",X"28",X"21",X"F0",X"38",X"C1",
		X"28",X"B2",X"88",X"01",X"AB",X"72",X"E0",X"29",X"90",X"28",X"A8",X"20",X"9A",X"50",X"E2",X"1A",
		X"80",X"49",X"D1",X"49",X"D1",X"5A",X"B4",X"1B",X"83",X"8A",X"94",X"0A",X"92",X"19",X"B4",X"1C",
		X"82",X"3F",X"84",X"9A",X"12",X"8B",X"85",X"0C",X"03",X"9B",X"30",X"8B",X"03",X"08",X"C4",X"8B",
		X"15",X"BB",X"24",X"8C",X"20",X"01",X"C8",X"38",X"BB",X"72",X"F0",X"39",X"A0",X"20",X"99",X"28",
		X"92",X"9A",X"05",X"9A",X"28",X"09",X"C3",X"7D",X"03",X"A9",X"12",X"9C",X"20",X"09",X"18",X"D5",
		X"1A",X"C1",X"31",X"D8",X"10",X"39",X"F1",X"3A",X"A1",X"12",X"D8",X"48",X"C0",X"69",X"B1",X"39",
		X"B0",X"69",X"A1",X"08",X"08",X"19",X"A3",X"09",X"91",X"5D",X"95",X"0B",X"83",X"98",X"2B",X"83",
		X"A9",X"12",X"3D",X"C5",X"1B",X"A1",X"58",X"D1",X"20",X"A9",X"13",X"C9",X"6A",X"A3",X"1B",X"02",
		X"9B",X"52",X"F1",X"29",X"A0",X"29",X"80",X"A5",X"0D",X"11",X"0E",X"15",X"AB",X"40",X"A8",X"28",
		X"A4",X"8A",X"84",X"9C",X"24",X"AB",X"22",X"8E",X"13",X"AA",X"24",X"C9",X"59",X"B3",X"2B",X"94",
		X"8A",X"01",X"0A",X"94",X"8C",X"22",X"9B",X"22",X"8C",X"03",X"99",X"91",X"69",X"C1",X"3B",X"00",
		X"92",X"9B",X"27",X"8D",X"04",X"A9",X"39",X"99",X"26",X"BC",X"51",X"C8",X"30",X"D0",X"38",X"B0",
		X"31",X"AE",X"23",X"9D",X"13",X"9B",X"06",X"9A",X"12",X"B9",X"38",X"A2",X"5D",X"83",X"9B",X"23",
		X"AB",X"31",X"B1",X"19",X"4B",X"D3",X"4B",X"C3",X"29",X"B1",X"5A",X"A3",X"0A",X"10",X"B0",X"68",
		X"F0",X"49",X"A2",X"2C",X"08",X"11",X"9B",X"50",X"C1",X"10",X"C2",X"00",X"A0",X"12",X"E8",X"7B",
		X"00",X"00",X"A1",X"3E",X"03",X"8D",X"04",X"9A",X"12",X"98",X"09",X"03",X"C9",X"40",X"D2",X"3B",
		X"B5",X"8B",X"12",X"1D",X"02",X"89",X"89",X"58",X"A8",X"25",X"E8",X"38",X"A8",X"49",X"98",X"21",
		X"D0",X"39",X"98",X"12",X"AA",X"A7",X"99",X"38",X"B1",X"40",X"C9",X"22",X"9A",X"B3",X"7A",X"B3",
		X"39",X"D1",X"39",X"9D",X"41",X"B9",X"25",X"C0",X"01",X"98",X"08",X"29",X"B3",X"01",X"BE",X"42",
		X"D0",X"3A",X"B5",X"8A",X"13",X"BC",X"60",X"AA",X"40",X"C1",X"29",X"A3",X"0E",X"22",X"9B",X"84",
		X"2D",X"93",X"0A",X"02",X"8C",X"14",X"9D",X"13",X"0D",X"02",X"08",X"A9",X"48",X"8B",X"14",X"0C",
		X"84",X"99",X"00",X"0A",X"03",X"B3",X"A8",X"2F",X"06",X"8B",X"82",X"2B",X"A3",X"2A",X"C1",X"40",
		X"AE",X"34",X"BB",X"33",X"B9",X"82",X"8A",X"58",X"B8",X"41",X"C0",X"10",X"B2",X"4D",X"B7",X"0A",
		X"81",X"2C",X"00",X"18",X"92",X"B9",X"68",X"A8",X"22",X"E0",X"10",X"80",X"B1",X"69",X"C2",X"19",
		X"09",X"A5",X"0B",X"10",X"93",X"0B",X"E2",X"6A",X"A1",X"21",X"AD",X"33",X"CA",X"31",X"B8",X"28",
		X"2B",X"B6",X"18",X"D8",X"48",X"90",X"91",X"3D",X"01",X"0A",X"A2",X"59",X"F2",X"3A",X"C2",X"29",
		X"19",X"0B",X"47",X"F7",X"AF",X"7E",X"4B",X"28",X"80",X"80",X"0A",X"4C",X"3C",X"5C",X"5D",X"5D",
		X"5D",X"4A",X"A6",X"D5",X"C8",X"5D",X"40",X"D5",X"8D",X"58",X"D3",X"3E",X"85",X"AD",X"52",X"DA",
		X"51",X"CA",X"51",X"AD",X"42",X"9A",X"B6",X"09",X"8B",X"42",X"A0",X"AA",X"42",X"B1",X"0D",X"04",
		X"8A",X"21",X"D8",X"22",X"A9",X"22",X"E8",X"11",X"0A",X"81",X"29",X"E1",X"00",X"2A",X"80",X"04",
		X"E9",X"6A",X"00",X"08",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"88",X"08",X"08",
		X"00",X"88",X"08",X"81",X"92",X"A3",X"B3",X"C3",X"0C",X"5A",X"94",X"0B",X"B3",X"78",X"AB",X"81",
		X"24",X"20",X"10",X"9A",X"FA",X"D9",X"16",X"30",X"DB",X"16",X"0C",X"84",X"8C",X"22",X"E2",X"1D",
		X"39",X"95",X"D3",X"A1",X"8A",X"5C",X"5C",X"3B",X"4B",X"29",X"94",X"E5",X"D4",X"A8",X"4D",X"5A",
		X"A6",X"D0",X"5D",X"13",X"C8",X"4A",X"B5",X"0C",X"13",X"AC",X"32",X"AD",X"41",X"AB",X"24",X"9A",
		X"A5",X"09",X"99",X"40",X"90",X"B1",X"49",X"80",X"B8",X"41",X"B2",X"8C",X"03",X"1B",X"03",X"BD",
		X"13",X"2D",X"02",X"0D",X"81",X"02",X"99",X"01",X"2B",X"D1",X"00",X"20",X"A9",X"12",X"20",X"F9",
		X"1F",X"78",X"B2",X"80",X"80",X"08",X"80",X"08",X"08",X"08",X"80",X"08",X"80",X"08",X"80",X"08",
		X"08",X"09",X"29",X"1B",X"28",X"93",X"BB",X"60",X"C8",X"15",X"8B",X"B9",X"22",X"16",X"00",X"09",
		X"8D",X"AC",X"B2",X"73",X"2B",X"F9",X"42",X"BC",X"42",X"D0",X"3B",X"A7",X"A0",X"3F",X"3A",X"84",
		X"D4",X"C3",X"B3",X"B3",X"B4",X"D5",X"C4",X"C4",X"C3",X"99",X"4D",X"5B",X"84",X"C2",X"1D",X"48",
		X"C4",X"8B",X"31",X"D1",X"3B",X"B5",X"0B",X"85",X"8B",X"04",X"8B",X"95",X"89",X"91",X"3A",X"8B",
		X"24",X"98",X"B0",X"40",X"90",X"C0",X"22",X"A0",X"9B",X"14",X"1B",X"11",X"E8",X"13",X"8B",X"22",
		X"BC",X"10",X"30",X"B0",X"33",X"FA",X"10",X"83",X"8A",X"01",X"48",X"D9",X"10",X"A1",X"48",X"A8",
		X"11",X"6C",X"F7",X"98",X"80",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"09",
		X"19",X"09",X"28",X"92",X"B1",X"3A",X"B2",X"7A",X"C0",X"23",X"29",X"9A",X"A0",X"80",X"82",X"36",
		X"01",X"DE",X"A0",X"44",X"9C",X"95",X"1C",X"95",X"9B",X"58",X"B5",X"9A",X"5C",X"28",X"A6",X"C3",
		X"C4",X"B3",X"B3",X"C4",X"C4",X"C4",X"B3",X"B2",X"0C",X"5C",X"39",X"A5",X"B1",X"2D",X"21",X"C2",
		X"1C",X"12",X"AA",X"58",X"B1",X"3A",X"B4",X"1B",X"A5",X"1A",X"B3",X"3A",X"B9",X"60",X"9A",X"83",
		X"19",X"9B",X"24",X"88",X"9B",X"14",X"1B",X"2C",X"91",X"40",X"B2",X"8D",X"01",X"38",X"B2",X"2D",
		X"A2",X"83",X"0A",X"83",X"2F",X"91",X"88",X"30",X"A8",X"23",X"8E",X"91",X"0A",X"04",X"0A",X"80",
		X"21",X"20",X"FF",X"7A",X"08",X"18",X"80",X"88",X"00",X"80",X"80",X"80",X"80",X"80",X"89",X"18",
		X"09",X"19",X"01",X"A1",X"2C",X"13",X"9B",X"86",X"29",X"BB",X"A9",X"02",X"18",X"09",X"AA",X"B2",
		X"73",X"41",X"CE",X"83",X"3A",X"E2",X"3C",X"A4",X"1E",X"21",X"D3",X"8B",X"7B",X"29",X"95",X"D4",
		X"B4",X"C3",X"B4",X"C3",X"C4",X"B4",X"B2",X"99",X"5C",X"3A",X"83",X"D3",X"8B",X"49",X"93",X"AA",
		X"80",X"80",X"80",X"80",X"00",X"00",X"80",X"80",X"80",X"88",X"80",X"90",X"80",X"89",X"80",X"80",
		X"80",X"10",X"80",X"01",X"80",X"10",X"80",X"80",X"80",X"A0",X"90",X"90",X"A8",X"80",X"90",X"80",
		X"00",X"02",X"81",X"81",X"10",X"00",X"00",X"88",X"88",X"80",X"A9",X"89",X"89",X"80",X"80",X"80",
		X"80",X"01",X"11",X"02",X"01",X"00",X"80",X"80",X"98",X"99",X"A9",X"98",X"B8",X"80",X"80",X"80",
		X"03",X"03",X"03",X"01",X"12",X"10",X"00",X"98",X"8A",X"A9",X"A9",X"B8",X"C0",X"B8",X"80",X"81",
		X"20",X"31",X"21",X"22",X"21",X"11",X"80",X"88",X"A9",X"AA",X"BA",X"C8",X"B8",X"A9",X"00",X"20",
		X"13",X"24",X"14",X"23",X"12",X"11",X"88",X"9A",X"AA",X"CB",X"BA",X"D9",X"B8",X"A9",X"00",X"31",
		X"23",X"43",X"33",X"33",X"22",X"10",X"88",X"AA",X"BC",X"AE",X"8C",X"9A",X"A8",X"80",X"02",X"43",
		X"34",X"43",X"43",X"33",X"31",X"08",X"9B",X"BD",X"CB",X"CB",X"CB",X"AA",X"A8",X"03",X"24",X"36",
		X"33",X"52",X"33",X"42",X"21",X"89",X"BD",X"BD",X"BC",X"BC",X"BB",X"A9",X"90",X"22",X"53",X"36",
		X"23",X"34",X"33",X"41",X"10",X"9A",X"CD",X"BC",X"BC",X"BB",X"BB",X"98",X"02",X"43",X"44",X"34",
		X"24",X"34",X"32",X"21",X"8A",X"BE",X"BC",X"CB",X"BC",X"BA",X"A8",X"01",X"33",X"54",X"23",X"34",
		X"34",X"42",X"31",X"19",X"BC",X"CC",X"CA",X"BD",X"AB",X"99",X"81",X"23",X"34",X"42",X"33",X"44",
		X"34",X"32",X"18",X"9C",X"CC",X"BB",X"CC",X"BA",X"B9",X"81",X"23",X"35",X"32",X"43",X"34",X"43",
		X"43",X"00",X"AB",X"CD",X"BB",X"CB",X"CA",X"B9",X"81",X"22",X"42",X"42",X"33",X"43",X"44",X"33",
		X"11",X"AB",X"DC",X"BC",X"BC",X"BA",X"C9",X"80",X"12",X"33",X"42",X"34",X"33",X"54",X"23",X"20",
		X"8B",X"CC",X"BD",X"BB",X"CB",X"AA",X"90",X"12",X"24",X"35",X"13",X"33",X"43",X"43",X"42",X"19",
		X"AC",X"CC",X"BB",X"DA",X"BA",X"A9",X"00",X"23",X"43",X"34",X"33",X"44",X"34",X"32",X"20",X"9A",
		X"CD",X"BC",X"CA",X"BB",X"AA",X"A8",X"02",X"33",X"53",X"52",X"23",X"43",X"43",X"33",X"21",X"AD",
		X"CC",X"BC",X"BB",X"CA",X"A9",X"98",X"12",X"24",X"35",X"13",X"33",X"44",X"43",X"32",X"18",X"AD",
		X"CC",X"BB",X"CA",X"BB",X"A9",X"80",X"13",X"52",X"42",X"33",X"34",X"43",X"43",X"32",X"88",X"BE",
		X"BC",X"CB",X"BC",X"AB",X"98",X"00",X"13",X"34",X"34",X"34",X"24",X"33",X"33",X"21",X"09",X"AC",
		X"EB",X"CC",X"CB",X"BB",X"99",X"80",X"13",X"34",X"43",X"33",X"42",X"43",X"44",X"31",X"19",X"AB",
		X"FB",X"BB",X"CB",X"AA",X"AA",X"A9",X"11",X"44",X"34",X"34",X"32",X"44",X"34",X"21",X"09",X"AB",
		X"EB",X"CC",X"BA",X"AB",X"A8",X"00",X"13",X"43",X"34",X"34",X"33",X"44",X"33",X"32",X"08",X"AB",
		X"EC",X"CC",X"BB",X"C9",X"A8",X"80",X"01",X"23",X"34",X"43",X"32",X"43",X"43",X"43",X"21",X"8A",
		X"CC",X"CC",X"CB",X"CA",X"AA",X"88",X"11",X"23",X"34",X"33",X"52",X"43",X"33",X"33",X"41",X"8B",
		X"CD",X"CC",X"BB",X"BC",X"AB",X"98",X"12",X"42",X"33",X"43",X"43",X"53",X"33",X"23",X"20",X"BF",
		X"CB",X"CA",X"AB",X"CA",X"99",X"81",X"02",X"43",X"34",X"32",X"33",X"54",X"42",X"11",X"80",X"09",
		X"DD",X"CB",X"AB",X"BB",X"BA",X"91",X"33",X"43",X"43",X"52",X"33",X"33",X"33",X"74",X"29",X"CB",
		X"B9",X"8C",X"DC",X"AA",X"90",X"00",X"01",X"23",X"43",X"32",X"35",X"24",X"33",X"21",X"09",X"CC",
		X"BB",X"DD",X"CB",X"99",X"89",X"90",X"33",X"32",X"43",X"52",X"32",X"34",X"53",X"19",X"11",X"CC",
		X"CB",X"BD",X"BB",X"98",X"9A",X"02",X"22",X"43",X"52",X"23",X"35",X"32",X"53",X"20",X"0A",X"AB",
		X"FE",X"AA",X"AB",X"99",X"99",X"01",X"34",X"23",X"23",X"52",X"24",X"32",X"45",X"21",X"88",X"8A",
		X"FC",X"BA",X"AB",X"E9",X"00",X"80",X"22",X"22",X"32",X"33",X"32",X"64",X"30",X"16",X"0B",X"A0",
		X"AF",X"B9",X"AC",X"98",X"A9",X"02",X"21",X"23",X"33",X"52",X"23",X"52",X"15",X"30",X"10",X"8C",
		X"E9",X"9D",X"BA",X"A9",X"BA",X"81",X"22",X"33",X"52",X"33",X"34",X"35",X"34",X"31",X"85",X"2E",
		X"BA",X"AE",X"B9",X"0A",X"B0",X"10",X"22",X"23",X"24",X"22",X"42",X"13",X"37",X"30",X"31",X"F8",
		X"8C",X"A9",X"D9",X"AA",X"88",X"00",X"11",X"32",X"24",X"21",X"42",X"17",X"10",X"52",X"09",X"08",
		X"F9",X"BB",X"B9",X"B9",X"91",X"08",X"23",X"34",X"33",X"34",X"32",X"44",X"23",X"44",X"11",X"98",
		X"FD",X"0B",X"D9",X"99",X"89",X"81",X"12",X"13",X"23",X"22",X"42",X"35",X"22",X"41",X"15",X"C9",
		X"9D",X"AA",X"CA",X"AA",X"A9",X"00",X"22",X"34",X"33",X"34",X"23",X"78",X"51",X"06",X"91",X"C0",
		X"9B",X"99",X"EB",X"09",X"80",X"81",X"12",X"21",X"31",X"41",X"22",X"37",X"02",X"24",X"91",X"9F",
		X"8D",X"8A",X"B8",X"B0",X"91",X"01",X"12",X"23",X"34",X"22",X"52",X"32",X"70",X"49",X"8A",X"0D",
		X"9B",X"E8",X"AA",X"A1",X"A1",X"03",X"12",X"32",X"32",X"43",X"26",X"31",X"50",X"40",X"A3",X"CC",
		X"AB",X"AF",X"99",X"A9",X"88",X"11",X"12",X"33",X"23",X"42",X"25",X"16",X"12",X"31",X"3C",X"9F",
		X"0D",X"0D",X"89",X"98",X"88",X"01",X"11",X"21",X"21",X"32",X"23",X"32",X"57",X"10",X"38",X"C0",
		X"DA",X"C9",X"BB",X"0C",X"88",X"80",X"22",X"32",X"33",X"34",X"14",X"14",X"24",X"71",X"08",X"1D",
		X"99",X"BD",X"AA",X"B8",X"B9",X"20",X"23",X"34",X"23",X"23",X"24",X"25",X"25",X"50",X"29",X"AB",
		X"9D",X"AE",X"8C",X"99",X"88",X"01",X"11",X"22",X"22",X"22",X"32",X"34",X"70",X"42",X"59",X"8A",
		X"AC",X"AD",X"9C",X"A8",X"99",X"01",X"12",X"32",X"32",X"33",X"23",X"43",X"55",X"40",X"11",X"89",
		X"FA",X"9C",X"AB",X"C9",X"0A",X"00",X"22",X"32",X"33",X"23",X"42",X"33",X"56",X"11",X"41",X"A9",
		X"F8",X"C9",X"C8",X"9A",X"80",X"00",X"12",X"13",X"22",X"22",X"32",X"34",X"56",X"12",X"39",X"C8",
		X"AD",X"9C",X"CB",X"A9",X"A9",X"01",X"23",X"42",X"23",X"32",X"33",X"35",X"25",X"37",X"11",X"8A",
		X"D9",X"AD",X"AB",X"9C",X"88",X"81",X"21",X"23",X"13",X"33",X"22",X"52",X"35",X"40",X"78",X"09",
		X"AA",X"BC",X"BD",X"B9",X"99",X"80",X"22",X"23",X"34",X"22",X"32",X"43",X"16",X"13",X"45",X"98",
		X"99",X"DC",X"CA",X"AA",X"99",X"88",X"13",X"22",X"34",X"22",X"23",X"33",X"37",X"22",X"53",X"20",
		X"E9",X"9C",X"CB",X"AD",X"A8",X"80",X"11",X"12",X"22",X"32",X"23",X"33",X"54",X"16",X"32",X"0A",
		X"9B",X"EA",X"DC",X"A9",X"B8",X"80",X"11",X"23",X"23",X"33",X"33",X"34",X"42",X"72",X"22",X"48",
		X"AB",X"DA",X"DC",X"BB",X"9A",X"A1",X"11",X"33",X"33",X"42",X"33",X"34",X"25",X"41",X"44",X"99",
		X"3E",X"AA",X"CA",X"BA",X"AB",X"88",X"12",X"32",X"43",X"23",X"33",X"52",X"23",X"74",X"21",X"2A",
		X"9C",X"BE",X"BB",X"CA",X"BA",X"98",X"13",X"33",X"43",X"32",X"33",X"43",X"35",X"55",X"28",X"80",
		X"BB",X"F9",X"AD",X"9B",X"9A",X"10",X"11",X"23",X"32",X"33",X"33",X"35",X"34",X"72",X"13",X"AA",
		X"CB",X"BE",X"9D",X"A9",X"A8",X"00",X"21",X"23",X"22",X"33",X"23",X"34",X"53",X"72",X"11",X"0A",
		X"CA",X"DB",X"BD",X"B9",X"A9",X"91",X"32",X"33",X"33",X"42",X"23",X"33",X"44",X"73",X"11",X"1B",
		X"9B",X"FC",X"AC",X"AA",X"99",X"81",X"22",X"23",X"23",X"33",X"32",X"42",X"72",X"23",X"40",X"82",
		X"CB",X"FA",X"DA",X"AA",X"98",X"00",X"12",X"22",X"33",X"32",X"33",X"34",X"33",X"77",X"30",X"88",
		X"BA",X"BB",X"FB",X"BB",X"C9",X"80",X"12",X"23",X"33",X"33",X"24",X"23",X"26",X"35",X"42",X"3A",
		X"DA",X"BD",X"AC",X"BA",X"89",X"81",X"21",X"33",X"23",X"33",X"32",X"43",X"36",X"62",X"10",X"2A",
		X"8F",X"AC",X"AB",X"AC",X"89",X"81",X"21",X"31",X"32",X"23",X"23",X"35",X"25",X"27",X"10",X"82",
		X"C9",X"DB",X"BA",X"AE",X"90",X"80",X"11",X"12",X"22",X"22",X"22",X"24",X"54",X"85",X"11",X"89",
		X"AE",X"9B",X"BE",X"90",X"B9",X"00",X"12",X"13",X"22",X"32",X"33",X"26",X"32",X"37",X"14",X"89",
		X"8B",X"FA",X"AC",X"C9",X"80",X"80",X"02",X"12",X"22",X"22",X"23",X"31",X"55",X"42",X"33",X"99",
		X"CE",X"BB",X"CC",X"8B",X"A8",X"81",X"22",X"32",X"34",X"22",X"22",X"33",X"47",X"35",X"08",X"10",
		X"D9",X"CB",X"AB",X"E9",X"A0",X"81",X"02",X"13",X"22",X"22",X"32",X"34",X"34",X"70",X"07",X"91",
		X"9A",X"AA",X"EA",X"9A",X"98",X"98",X"12",X"22",X"32",X"32",X"33",X"34",X"34",X"74",X"00",X"01",
		X"D8",X"AD",X"9C",X"A9",X"B9",X"91",X"12",X"23",X"32",X"41",X"31",X"42",X"27",X"07",X"93",X"A0",
		X"A9",X"CA",X"BC",X"AA",X"99",X"00",X"22",X"24",X"22",X"32",X"23",X"36",X"26",X"84",X"05",X"B8",
		X"9B",X"9E",X"AA",X"B9",X"A0",X"81",X"21",X"33",X"33",X"33",X"43",X"42",X"53",X"44",X"31",X"9C",
		X"BB",X"FA",X"CA",X"AB",X"99",X"11",X"12",X"42",X"32",X"32",X"23",X"34",X"72",X"14",X"20",X"99",
		X"AF",X"BB",X"AB",X"F9",X"88",X"00",X"01",X"12",X"22",X"22",X"23",X"41",X"37",X"14",X"02",X"8B",
		X"8B",X"FA",X"BE",X"99",X"99",X"18",X"11",X"13",X"22",X"22",X"33",X"25",X"22",X"73",X"A6",X"0B",
		X"0A",X"CA",X"BD",X"8B",X"98",X"88",X"11",X"21",X"24",X"23",X"22",X"43",X"33",X"75",X"90",X"5A",
		X"99",X"AD",X"9B",X"C9",X"09",X"98",X"11",X"22",X"22",X"33",X"51",X"22",X"53",X"43",X"31",X"9D",
		X"9B",X"EC",X"BA",X"AA",X"A9",X"08",X"13",X"34",X"33",X"34",X"23",X"34",X"43",X"54",X"20",X"08",
		X"FB",X"A9",X"BC",X"BB",X"B9",X"90",X"13",X"43",X"24",X"23",X"23",X"53",X"13",X"74",X"80",X"09",
		X"AA",X"BF",X"BB",X"AB",X"B8",X"88",X"31",X"33",X"43",X"34",X"23",X"34",X"62",X"15",X"20",X"9B",
		X"CB",X"CA",X"BD",X"BB",X"91",X"18",X"02",X"33",X"33",X"53",X"23",X"33",X"46",X"42",X"80",X"8A",
		X"CB",X"CC",X"CB",X"A9",X"B9",X"80",X"03",X"33",X"44",X"33",X"32",X"55",X"41",X"81",X"21",X"8B",
		X"FB",X"9A",X"EB",X"A8",X"89",X"00",X"12",X"23",X"34",X"22",X"34",X"43",X"32",X"25",X"38",X"BD",
		X"BB",X"CD",X"CB",X"A0",X"98",X"88",X"23",X"33",X"42",X"33",X"63",X"42",X"01",X"34",X"0B",X"CC",
		X"BD",X"AA",X"BB",X"BB",X"A8",X"23",X"43",X"34",X"34",X"34",X"33",X"43",X"33",X"20",X"89",X"BF",
		X"FC",X"B9",X"A9",X"98",X"08",X"00",X"22",X"35",X"32",X"33",X"43",X"53",X"34",X"31",X"AC",X"CC",
		X"DA",X"9B",X"AB",X"B9",X"81",X"32",X"33",X"44",X"33",X"43",X"42",X"12",X"14",X"22",X"28",X"BF",
		X"EB",X"BB",X"BB",X"99",X"00",X"13",X"33",X"44",X"33",X"33",X"44",X"33",X"22",X"22",X"8B",X"FC",
		X"CC",X"BC",X"A9",X"98",X"00",X"02",X"13",X"34",X"43",X"33",X"43",X"43",X"31",X"18",X"BD",X"DD",
		X"BB",X"CB",X"A8",X"80",X"01",X"22",X"34",X"34",X"34",X"23",X"42",X"23",X"42",X"10",X"CD",X"DC",
		X"BB",X"BB",X"99",X"81",X"12",X"33",X"53",X"34",X"33",X"45",X"23",X"21",X"09",X"AD",X"CB",X"DA",
		X"CA",X"9A",X"A9",X"88",X"22",X"43",X"34",X"34",X"34",X"33",X"43",X"21",X"08",X"CD",X"CB",X"DA",
		X"BA",X"AA",X"A8",X"81",X"23",X"53",X"33",X"53",X"33",X"53",X"32",X"21",X"8B",X"CD",X"CB",X"CB",
		X"CB",X"AB",X"98",X"01",X"33",X"44",X"33",X"34",X"33",X"53",X"42",X"21",X"8A",X"BD",X"BD",X"CB",
		X"CB",X"AB",X"98",X"01",X"23",X"43",X"42",X"34",X"33",X"53",X"33",X"21",X"8A",X"DB",X"DC",X"BB",
		X"CB",X"BA",X"A9",X"82",X"33",X"53",X"34",X"34",X"23",X"52",X"33",X"21",X"8A",X"BE",X"BD",X"BC",
		X"BB",X"BB",X"A9",X"80",X"23",X"53",X"35",X"23",X"43",X"34",X"42",X"32",X"18",X"BD",X"CD",X"BB",
		X"CB",X"BB",X"90",X"02",X"24",X"33",X"43",X"33",X"43",X"42",X"33",X"32",X"09",X"CD",X"CB",X"DB",
		X"CB",X"B9",X"A9",X"01",X"14",X"23",X"42",X"33",X"43",X"35",X"33",X"43",X"20",X"9C",X"DB",X"DB",
		X"CB",X"BB",X"A9",X"80",X"22",X"35",X"33",X"33",X"44",X"24",X"33",X"52",X"10",X"9B",X"CD",X"BC",
		X"BC",X"BA",X"A9",X"80",X"12",X"34",X"43",X"23",X"34",X"35",X"33",X"33",X"19",X"AE",X"CB",X"CC",
		X"BA",X"BB",X"A9",X"01",X"14",X"24",X"33",X"33",X"43",X"44",X"34",X"32",X"08",X"BD",X"CB",X"DB",
		X"BC",X"AB",X"98",X"01",X"23",X"34",X"34",X"23",X"43",X"35",X"33",X"32",X"0A",X"CD",X"BD",X"BC",
		X"BB",X"AB",X"98",X"02",X"24",X"24",X"32",X"42",X"33",X"43",X"52",X"33",X"08",X"AD",X"CC",X"BC",
		X"CA",X"BA",X"A8",X"81",X"13",X"34",X"42",X"33",X"33",X"44",X"42",X"42",X"00",X"9C",X"BD",X"CA",
		X"CA",X"BA",X"A9",X"80",X"22",X"34",X"24",X"33",X"33",X"52",X"43",X"33",X"31",X"8C",X"CD",X"BC",
		X"BC",X"BB",X"AB",X"99",X"02",X"34",X"42",X"34",X"24",X"22",X"34",X"34",X"31",X"19",X"BD",X"CB",
		X"DB",X"CA",X"BA",X"A9",X"01",X"14",X"23",X"35",X"22",X"33",X"44",X"33",X"41",X"18",X"AD",X"BD",
		X"BB",X"CB",X"CA",X"A9",X"81",X"13",X"42",X"34",X"23",X"34",X"33",X"53",X"32",X"28",X"BC",X"CD",
		X"BC",X"BC",X"BB",X"AA",X"80",X"22",X"43",X"34",X"33",X"43",X"34",X"35",X"32",X"20",X"9C",X"CB",
		X"DB",X"CB",X"BB",X"BA",X"98",X"22",X"43",X"43",X"42",X"33",X"35",X"34",X"34",X"11",X"9A",X"BE",
		X"BC",X"BC",X"BB",X"AB",X"A8",X"02",X"35",X"24",X"32",X"24",X"23",X"43",X"43",X"31",X"0A",X"BE",
		X"CB",X"CB",X"BC",X"BB",X"A9",X"01",X"23",X"53",X"33",X"34",X"34",X"25",X"23",X"41",X"18",X"AC",
		X"CB",X"CB",X"CA",X"CB",X"A9",X"90",X"22",X"34",X"33",X"43",X"24",X"33",X"44",X"33",X"20",X"9B",
		X"DC",X"CB",X"CB",X"BC",X"BA",X"98",X"02",X"34",X"33",X"43",X"24",X"33",X"44",X"33",X"21",X"0A",
		X"CD",X"BC",X"BC",X"CA",X"BA",X"A9",X"81",X"23",X"43",X"34",X"34",X"23",X"43",X"43",X"32",X"19",
		X"AD",X"CC",X"BB",X"CC",X"BA",X"B9",X"90",X"22",X"35",X"32",X"42",X"33",X"52",X"42",X"31",X"10",
		X"AB",X"EB",X"CB",X"CC",X"AB",X"AA",X"88",X"21",X"34",X"34",X"24",X"23",X"34",X"34",X"32",X"18",
		X"8C",X"BD",X"CB",X"CB",X"BC",X"AA",X"98",X"11",X"23",X"61",X"33",X"33",X"44",X"24",X"22",X"10",
		X"8B",X"BE",X"BD",X"BB",X"BC",X"BA",X"98",X"82",X"32",X"62",X"24",X"22",X"34",X"33",X"33",X"31",
		X"9C",X"CC",X"BD",X"BC",X"BB",X"BB",X"99",X"01",X"24",X"42",X"34",X"34",X"33",X"43",X"33",X"12",
		X"99",X"DB",X"EB",X"BC",X"CA",X"BA",X"9A",X"00",X"13",X"43",X"43",X"35",X"23",X"43",X"32",X"20",
		X"0A",X"BD",X"DB",X"CB",X"CB",X"AB",X"AA",X"80",X"22",X"43",X"53",X"42",X"33",X"43",X"33",X"31",
		X"09",X"BC",X"EB",X"CC",X"BB",X"BB",X"CA",X"88",X"02",X"25",X"23",X"53",X"14",X"23",X"33",X"32",
		X"00",X"AB",X"EC",X"BD",X"BC",X"AA",X"BA",X"99",X"03",X"14",X"23",X"63",X"33",X"43",X"23",X"33",
		X"18",X"8C",X"CB",X"EB",X"BC",X"BC",X"A9",X"A9",X"01",X"23",X"35",X"42",X"42",X"33",X"33",X"33",
		X"18",X"9B",X"CD",X"BD",X"AC",X"BA",X"A9",X"8A",X"01",X"32",X"45",X"24",X"23",X"43",X"23",X"22",
		X"88",X"AB",X"DB",X"EA",X"BB",X"BD",X"98",X"A0",X"02",X"23",X"43",X"44",X"23",X"42",X"32",X"28",
		X"0A",X"9C",X"BE",X"BB",X"CA",X"AC",X"99",X"80",X"03",X"25",X"23",X"52",X"33",X"52",X"20",X"10",
		X"8A",X"AD",X"BC",X"CB",X"CA",X"AB",X"8A",X"88",X"40",X"34",X"51",X"33",X"42",X"42",X"22",X"10",
		X"09",X"BB",X"DC",X"BC",X"BB",X"BD",X"98",X"A8",X"02",X"13",X"35",X"34",X"23",X"52",X"22",X"11",
		X"19",X"8B",X"AC",X"CB",X"BD",X"AA",X"AA",X"A8",X"81",X"13",X"32",X"51",X"33",X"42",X"33",X"02",
		X"89",X"9A",X"CA",X"CB",X"CA",X"BB",X"CA",X"88",X"11",X"22",X"43",X"34",X"33",X"52",X"31",X"20",
		X"08",X"9B",X"BC",X"CB",X"BD",X"AA",X"9B",X"89",X"18",X"33",X"41",X"34",X"34",X"33",X"24",X"01",
		X"80",X"A9",X"CA",X"CA",X"BC",X"C9",X"A9",X"A0",X"81",X"21",X"24",X"33",X"23",X"32",X"31",X"21",
		X"89",X"8B",X"AB",X"BC",X"BB",X"C8",X"C9",X"89",X"12",X"03",X"12",X"43",X"33",X"32",X"32",X"10",
		X"80",X"9A",X"AB",X"CA",X"BC",X"BB",X"B9",X"99",X"00",X"20",X"32",X"23",X"33",X"32",X"31",X"11",
		X"09",X"89",X"AB",X"AC",X"9B",X"C9",X"A8",X"0B",X"38",X"12",X"12",X"40",X"32",X"21",X"21",X"08",
		X"0A",X"8A",X"AB",X"AB",X"9C",X"9A",X"08",X"A0",X"28",X"12",X"40",X"31",X"31",X"41",X"01",X"08",
		X"0A",X"99",X"BA",X"AB",X"9C",X"9A",X"08",X"08",X"00",X"30",X"33",X"12",X"21",X"30",X"10",X"19",
		X"89",X"9B",X"9A",X"AB",X"8C",X"9A",X"08",X"08",X"00",X"30",X"31",X"32",X"21",X"21",X"10",X"09",
		X"09",X"9A",X"9A",X"BA",X"9B",X"8A",X"98",X"08",X"10",X"23",X"03",X"12",X"20",X"30",X"28",X"08",
		X"09",X"9B",X"8A",X"BA",X"9B",X"8B",X"88",X"08",X"08",X"21",X"48",X"40",X"22",X"12",X"11",X"00",
		X"90",X"99",X"B8",X"BA",X"B8",X"B8",X"B8",X"80",X"81",X"20",X"31",X"21",X"22",X"13",X"01",X"80",
		X"80",X"A8",X"B9",X"B9",X"CA",X"88",X"08",X"00",X"02",X"08",X"00",X"00",X"28",X"08",X"00",X"08",
		X"18",X"08",X"00",X"88",X"18",X"88",X"08",X"08",X"08",X"08",X"08",X"09",X"19",X"08",X"08",X"08",
		X"80",X"90",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"88",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"81",X"91",X"90",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"A0",X"80",X"80",X"91",X"80",X"10",X"80",X"01",X"10",X"81",X"80",X"08",X"80",
		X"90",X"80",X"80",X"A0",X"10",X"81",X"80",X"08",X"80",X"9F",X"DA",X"98",X"02",X"54",X"54",X"53",
		X"32",X"1B",X"DB",X"CA",X"BB",X"FF",X"B8",X"11",X"37",X"38",X"88",X"AE",X"90",X"01",X"01",X"15",
		X"40",X"9B",X"E8",X"01",X"15",X"09",X"D8",X"00",X"32",X"BC",X"80",X"52",X"9E",X"80",X"13",X"9C",
		X"80",X"10",X"88",X"04",X"39",X"D9",X"80",X"07",X"8C",X"00",X"80",X"00",X"93",X"4E",X"83",X"0D",
		X"02",X"B4",X"A9",X"18",X"85",X"B8",X"00",X"19",X"03",X"C0",X"87",X"A1",X"90",X"98",X"4B",X"80",
		X"13",X"E8",X"5B",X"82",X"81",X"B2",X"B4",X"B2",X"1D",X"01",X"88",X"2A",X"7A",X"91",X"86",X"B8",
		X"84",X"9A",X"03",X"0D",X"08",X"07",X"9A",X"03",X"AA",X"08",X"04",X"A8",X"00",X"08",X"03",X"A9",
		X"81",X"19",X"83",X"19",X"A8",X"98",X"17",X"7C",X"C0",X"07",X"0A",X"C0",X"03",X"29",X"F8",X"00",
		X"04",X"0B",X"A0",X"00",X"14",X"8B",X"90",X"00",X"13",X"0A",X"98",X"10",X"11",X"77",X"9C",X"90",
		X"08",X"00",X"14",X"8B",X"A8",X"08",X"00",X"10",X"12",X"40",X"DB",X"98",X"00",X"00",X"01",X"23",
		X"38",X"AD",X"BB",X"A8",X"80",X"01",X"11",X"33",X"35",X"53",X"09",X"CF",X"AA",X"88",X"10",X"01",
		X"81",X"12",X"03",X"43",X"43",X"20",X"CD",X"CB",X"A8",X"88",X"08",X"08",X"12",X"23",X"13",X"32",
		X"14",X"23",X"33",X"32",X"18",X"08",X"89",X"9B",X"AB",X"CA",X"CA",X"B0",X"83",X"80",X"08",X"81",
		X"25",X"53",X"30",X"AD",X"DB",X"BA",X"02",X"61",X"08",X"89",X"AB",X"D9",X"01",X"61",X"8A",X"C8",
		X"90",X"12",X"53",X"54",X"42",X"1B",X"FC",X"A8",X"83",X"11",X"80",X"26",X"31",X"AF",X"C0",X"23",
		X"51",X"BF",X"A8",X"16",X"38",X"CC",X"81",X"42",X"9E",X"80",X"14",X"8C",X"91",X"22",X"BB",X"02",
		X"4A",X"B1",X"20",X"B0",X"25",X"BA",X"47",X"BA",X"11",X"B2",X"5C",X"83",X"AA",X"5B",X"10",X"A4",
		X"99",X"81",X"6C",X"80",X"39",X"A0",X"81",X"82",X"B0",X"49",X"80",X"A9",X"54",X"D9",X"31",X"D0",
		X"08",X"03",X"9C",X"02",X"1B",X"00",X"01",X"AB",X"17",X"3C",X"B8",X"03",X"69",X"D8",X"24",X"0E",
		X"80",X"20",X"A9",X"02",X"1A",X"A0",X"25",X"8C",X"90",X"34",X"8C",X"A0",X"02",X"32",X"8D",X"B9",
		X"02",X"45",X"0B",X"D8",X"81",X"02",X"20",X"99",X"BA",X"91",X"14",X"53",X"0B",X"DA",X"90",X"00",
		X"11",X"23",X"21",X"9B",X"DB",X"A8",X"00",X"11",X"22",X"32",X"21",X"8A",X"CB",X"AC",X"CC",X"A9",
		X"82",X"35",X"31",X"12",X"23",X"21",X"8C",X"FB",X"BC",X"A9",X"90",X"32",X"32",X"20",X"38",X"32",
		X"32",X"41",X"18",X"AC",X"A9",X"AB",X"9C",X"BB",X"C9",X"90",X"82",X"13",X"31",X"24",X"03",X"33",
		X"22",X"02",X"11",X"02",X"89",X"9A",X"AB",X"A9",X"99",X"98",X"A9",X"8B",X"89",X"91",X"80",X"10",
		X"03",X"84",X"03",X"11",X"81",X"12",X"12",X"09",X"CB",X"B9",X"98",X"A9",X"CB",X"0C",X"0B",X"09",
		X"AB",X"91",X"56",X"33",X"08",X"00",X"88",X"00",X"38",X"8C",X"BC",X"B0",X"35",X"34",X"30",X"9C",
		X"DA",X"15",X"40",X"AB",X"B9",X"01",X"11",X"13",X"2D",X"92",X"73",X"AF",X"D9",X"14",X"51",X"BC",
		X"B0",X"55",X"0D",X"A1",X"31",X"AC",X"84",X"2A",X"C0",X"41",X"C9",X"30",X"B0",X"39",X"88",X"A2",
		X"69",X"D0",X"49",X"92",X"A0",X"2C",X"87",X"A8",X"29",X"98",X"14",X"8E",X"03",X"9A",X"28",X"80",
		X"18",X"A8",X"03",X"09",X"C8",X"52",X"BD",X"13",X"1A",X"B9",X"35",X"8C",X"A3",X"68",X"C9",X"03",
		X"39",X"CA",X"03",X"58",X"BB",X"82",X"34",X"1C",X"CA",X"13",X"41",X"8D",X"A9",X"13",X"32",X"9C",
		X"AA",X"01",X"32",X"20",X"9B",X"C9",X"88",X"12",X"33",X"20",X"BC",X"CA",X"98",X"23",X"41",X"18",
		X"08",X"8A",X"BC",X"B8",X"13",X"42",X"38",X"09",X"08",X"09",X"BD",X"AA",X"01",X"43",X"21",X"08",
		X"00",X"08",X"09",X"0A",X"89",X"89",X"89",X"08",X"01",X"28",X"00",X"11",X"08",X"18",X"88",X"99",
		X"09",X"08",X"98",X"89",X"08",X"00",X"18",X"28",X"08",X"08",X"18",X"18",X"08",X"08",X"08",X"08",
		X"88",X"09",X"08",X"08",X"08",X"98",X"08",X"08",X"08",X"08",X"28",X"08",X"08",X"08",X"08",X"08",
		X"08",X"88",X"08",X"18",X"88",X"08",X"08",X"08",X"08",X"08",X"08",X"18",X"08",X"08",X"80",X"88",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"08",X"00",X"88",X"28",X"89",X"21",X"98",X"80",X"01",X"99",X"84",X"8A",X"D5",X"B6",X"0A",X"B8",
		X"34",X"29",X"AD",X"B9",X"02",X"35",X"31",X"10",X"99",X"AA",X"BC",X"AA",X"D9",X"AC",X"98",X"99",
		X"09",X"10",X"28",X"11",X"22",X"12",X"40",X"31",X"21",X"31",X"21",X"21",X"20",X"20",X"28",X"10",
		X"08",X"18",X"08",X"88",X"08",X"08",X"89",X"89",X"08",X"89",X"88",X"89",X"99",X"09",X"88",X"99",
		X"88",X"88",X"09",X"08",X"18",X"09",X"09",X"0A",X"89",X"A9",X"BC",X"BF",X"BB",X"BD",X"AC",X"AA",
		X"BB",X"BB",X"C9",X"88",X"11",X"44",X"35",X"43",X"34",X"43",X"33",X"43",X"33",X"33",X"43",X"33",
		X"43",X"34",X"13",X"31",X"40",X"11",X"08",X"90",X"A9",X"80",X"80",X"37",X"33",X"30",X"EF",X"CC",
		X"CB",X"BC",X"BA",X"BB",X"CB",X"AB",X"98",X"23",X"54",X"34",X"33",X"43",X"24",X"35",X"35",X"20",
		X"8B",X"BC",X"CB",X"CB",X"A9",X"88",X"12",X"34",X"36",X"43",X"20",X"9A",X"CD",X"BA",X"80",X"02",
		X"36",X"43",X"89",X"BC",X"AA",X"A9",X"81",X"37",X"52",X"8B",X"EA",X"01",X"04",X"30",X"AD",X"A0",
		X"03",X"40",X"AB",X"92",X"1D",X"A0",X"37",X"2B",X"D8",X"02",X"48",X"C9",X"03",X"3B",X"C8",X"33",
		X"CA",X"61",X"CA",X"12",X"3A",X"BA",X"03",X"3A",X"B7",X"9A",X"40",X"C3",X"8C",X"40",X"91",X"D8",
		X"18",X"5A",X"89",X"19",X"5B",X"3B",X"3B",X"4B",X"3C",X"3B",X"59",X"0D",X"18",X"38",X"9B",X"01",
		X"02",X"0B",X"14",X"8B",X"82",X"12",X"08",X"FD",X"06",X"88",X"A8",X"11",X"08",X"08",X"08",X"89",
		X"14",X"39",X"FB",X"87",X"0A",X"A0",X"21",X"88",X"82",X"88",X"89",X"35",X"0F",X"A0",X"50",X"C8",
		X"02",X"80",X"88",X"18",X"80",X"87",X"8E",X"81",X"38",X"D8",X"20",X"08",X"80",X"00",X"99",X"70",
		X"D8",X"12",X"8C",X"82",X"00",X"80",X"00",X"9A",X"62",X"CC",X"05",X"0A",X"A1",X"29",X"09",X"02",
		X"3F",X"4D",X"3B",X"15",X"9B",X"98",X"11",X"60",X"89",X"BB",X"80",X"10",X"11",X"11",X"23",X"53",
		X"18",X"AB",X"BB",X"AB",X"BE",X"BA",X"AA",X"98",X"00",X"13",X"24",X"23",X"43",X"33",X"33",X"33",
		X"42",X"23",X"22",X"21",X"20",X"11",X"89",X"99",X"AB",X"AB",X"BC",X"AD",X"AA",X"BB",X"CB",X"AC",
		X"AC",X"AA",X"BB",X"CB",X"BB",X"BB",X"B9",X"CB",X"A9",X"BB",X"8C",X"9A",X"9A",X"89",X"8A",X"08",
		X"88",X"08",X"00",X"08",X"11",X"18",X"11",X"28",X"21",X"48",X"31",X"30",X"33",X"12",X"12",X"48",
		X"21",X"30",X"21",X"21",X"11",X"10",X"20",X"18",X"10",X"18",X"18",X"08",X"08",X"08",X"08",X"08",
		X"08",X"89",X"08",X"98",X"09",X"88",X"0A",X"08",X"99",X"88",X"09",X"88",X"89",X"89",X"08",X"FF",
		X"08",X"88",X"08",X"08",X"19",X"19",X"08",X"08",X"08",X"80",X"09",X"08",X"88",X"08",X"08",X"08",
		X"00",X"08",X"18",X"00",X"08",X"09",X"08",X"00",X"00",X"18",X"08",X"88",X"18",X"10",X"08",X"10",
		X"12",X"0F",X"FF",X"A0",X"15",X"64",X"20",X"9E",X"DA",X"00",X"37",X"28",X"CC",X"80",X"35",X"8B",
		X"C0",X"25",X"8D",X"92",X"59",X"D0",X"50",X"D8",X"59",X"C4",X"1D",X"30",X"D5",X"A9",X"5D",X"4B",
		X"3B",X"2A",X"3C",X"5B",X"28",X"A3",X"9A",X"22",X"AA",X"01",X"20",X"08",X"08",X"8A",X"AB",X"17",
		X"8B",X"28",X"A4",X"B2",X"90",X"19",X"A0",X"28",X"08",X"A9",X"22",X"C1",X"0A",X"13",X"D8",X"10",
		X"09",X"8A",X"21",X"C2",X"A2",X"B8",X"21",X"84",X"9F",X"11",X"A2",X"B4",X"8A",X"31",X"B8",X"96",
		X"98",X"21",X"19",X"08",X"08",X"98",X"08",X"08",X"18",X"80",X"18",X"0A",X"0A",X"98",X"12",X"18",
		X"08",X"09",X"08",X"08",X"11",X"10",X"09",X"98",X"90",X"10",X"28",X"20",X"89",X"08",X"90",X"08",
		X"02",X"89",X"0A",X"89",X"18",X"10",X"08",X"20",X"08",X"08",X"88",X"00",X"11",X"29",X"18",X"08",
		X"89",X"38",X"08",X"08",X"08",X"01",X"A8",X"19",X"19",X"18",X"C3",X"8B",X"9A",X"A5",X"AA",X"18",
		X"D4",X"8B",X"A9",X"88",X"34",X"AF",X"48",X"A2",X"0C",X"5A",X"92",X"38",X"98",X"81",X"31",X"AF",
		X"C5",X"1E",X"38",X"A4",X"B4",X"B3",X"8C",X"59",X"A3",X"19",X"D1",X"31",X"99",X"80",X"B8",X"08",
		X"05",X"03",X"20",X"FF",X"01",X"30",X"E8",X"22",X"D0",X"28",X"B3",X"0D",X"4A",X"84",X"D2",X"90",
		X"2C",X"4B",X"3C",X"3B",X"3C",X"3B",X"5B",X"4B",X"2A",X"01",X"B6",X"B2",X"99",X"5B",X"10",X"A4",
		X"A9",X"6B",X"84",X"A8",X"3B",X"84",X"A9",X"21",X"D0",X"5B",X"81",X"2C",X"03",X"9B",X"07",X"A9",
		X"04",X"A9",X"03",X"8C",X"01",X"4C",X"88",X"31",X"D8",X"04",X"0C",X"80",X"31",X"D8",X"01",X"4B",
		X"A0",X"04",X"1D",X"90",X"13",X"1E",X"88",X"03",X"2C",X"A0",X"01",X"68",X"C8",X"80",X"24",X"8D",
		X"88",X"01",X"40",X"BB",X"00",X"04",X"38",X"EA",X"00",X"12",X"40",X"DA",X"80",X"02",X"42",X"AD",
		X"A0",X"00",X"25",X"19",X"CA",X"91",X"02",X"43",X"0B",X"F9",X"80",X"02",X"42",X"8A",X"CB",X"80",
		X"02",X"44",X"18",X"BD",X"B8",X"01",X"24",X"41",X"8A",X"CC",X"90",X"01",X"34",X"31",X"9A",X"EB",
		X"A0",X"02",X"34",X"41",X"89",X"CC",X"A9",X"01",X"23",X"43",X"18",X"AB",X"EB",X"A8",X"03",X"35",
		X"32",X"09",X"AC",X"CC",X"98",X"12",X"34",X"31",X"08",X"9B",X"DB",X"C9",X"01",X"34",X"33",X"10",
		X"99",X"BC",X"CC",X"A8",X"13",X"34",X"32",X"18",X"9A",X"BC",X"DB",X"A8",X"22",X"53",X"31",X"08",
		X"89",X"AB",X"DB",X"CA",X"02",X"43",X"33",X"10",X"98",X"AA",X"AD",X"CA",X"A8",X"33",X"52",X"30",
		X"08",X"09",X"99",X"9B",X"9D",X"90",X"23",X"22",X"10",X"08",X"09",X"09",X"89",X"99",X"0B",X"38",
		X"11",X"10",X"08",X"08",X"09",X"09",X"09",X"98",X"08",X"10",X"18",X"18",X"08",X"09",X"19",X"08",
		X"88",X"09",X"18",X"00",X"08",X"08",X"19",X"08",X"08",X"08",X"09",X"08",X"08",X"18",X"08",X"08",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"08",X"18",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"09",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C3",X"87",X"E0",X"02",X"00",X"00",X"20",X"00",X"00",X"00",X"30",X"00",X"30",X"00",X"20",X"00",
		X"20",X"00",X"30",X"00",X"30",X"00",X"20",X"00",X"40",X"00",X"30",X"00",X"30",X"00",X"20",X"00",
		X"60",X"00",X"30",X"00",X"30",X"00",X"20",X"00",X"80",X"00",X"30",X"00",X"30",X"00",X"20",X"00",
		X"A0",X"00",X"30",X"00",X"30",X"00",X"20",X"00",X"C0",X"00",X"30",X"00",X"30",X"00",X"00",X"00",
		X"1E",X"49",X"00",X"30",X"C0",X"00",X"20",X"00",X"20",X"00",X"30",X"3D",X"E0",X"00",X"E0",X"00",
		X"50",X"07",X"00",X"E0",X"00",X"00",X"D3",X"1F",X"94",X"03",X"05",X"00",X"01",X"09",X"E0",X"23",
		X"ED",X"00",X"7C",X"BA",X"C0",X"7D",X"BB",X"C9",X"A7",X"ED",X"52",X"23",X"C9",X"23",X"7C",X"B5",
		X"2B",X"C9",X"7D",X"02",X"03",X"7C",X"02",X"03",X"C9",X"1A",X"6F",X"13",X"1A",X"67",X"C9",X"DB",
		X"04",X"E6",X"80",X"32",X"FD",X"FE",X"C9",X"31",X"00",X"F6",X"CD",X"60",X"F0",X"CD",X"23",X"EB",
		X"31",X"00",X"F6",X"21",X"03",X"E0",X"06",X"5F",X"AF",X"77",X"23",X"10",X"FC",X"CD",X"CA",X"E0",
		X"AF",X"32",X"FD",X"FE",X"32",X"FE",X"FE",X"3A",X"04",X"E0",X"A7",X"CC",X"82",X"F2",X"06",X"01",
		X"CD",X"3D",X"F3",X"CD",X"B6",X"F2",X"06",X"01",X"CD",X"3D",X"F3",X"CD",X"B6",X"F2",X"0E",X"00",
		X"CD",X"80",X"F3",X"0E",X"00",X"CD",X"80",X"F3",X"18",X"C6",X"AF",X"32",X"03",X"E0",X"32",X"FD",
		X"FE",X"32",X"01",X"F6",X"21",X"05",X"E0",X"22",X"5D",X"E0",X"21",X"04",X"ED",X"22",X"5F",X"E0",
		X"06",X"4D",X"36",X"20",X"23",X"10",X"FB",X"21",X"3D",X"EB",X"CD",X"4E",X"F2",X"CD",X"1E",X"F1",
		X"FE",X"01",X"CA",X"36",X"E1",X"FE",X"02",X"CA",X"96",X"E1",X"FE",X"03",X"CA",X"36",X"E2",X"FE",
		X"04",X"CA",X"47",X"E2",X"FE",X"06",X"CA",X"D0",X"F0",X"FE",X"07",X"20",X"BD",X"21",X"85",X"EB",
		X"CD",X"4E",X"F2",X"CD",X"1E",X"F1",X"FE",X"01",X"CA",X"CE",X"EE",X"FE",X"02",X"CA",X"00",X"F7",
		X"FE",X"03",X"CA",X"00",X"F4",X"FE",X"04",X"CA",X"9F",X"ED",X"FE",X"05",X"CA",X"00",X"FB",X"FE",
		X"07",X"C2",X"0D",X"E1",X"18",X"94",X"21",X"3F",X"EB",X"0E",X"05",X"CD",X"FE",X"EA",X"CD",X"75",
		X"E2",X"CD",X"82",X"F2",X"21",X"20",X"EC",X"CD",X"4E",X"F2",X"CD",X"49",X"F1",X"CD",X"D3",X"EA",
		X"20",X"F8",X"21",X"22",X"EC",X"0E",X"04",X"CD",X"FE",X"EA",X"CD",X"12",X"EB",X"21",X"2D",X"EC",
		X"CD",X"4E",X"F2",X"CD",X"49",X"F1",X"CD",X"DD",X"EA",X"20",X"F8",X"38",X"26",X"21",X"2F",X"EC",
		X"0E",X"04",X"CD",X"FE",X"EA",X"CD",X"12",X"EB",X"21",X"47",X"EC",X"CD",X"4E",X"F2",X"CD",X"49",
		X"F1",X"CD",X"DD",X"EA",X"20",X"F8",X"38",X"0B",X"21",X"4F",X"EC",X"0E",X"02",X"CD",X"FE",X"EA",
		X"CD",X"12",X"EB",X"C3",X"19",X"E9",X"21",X"49",X"EB",X"0E",X"04",X"CD",X"FE",X"EA",X"CD",X"75",
		X"E2",X"CD",X"82",X"F2",X"21",X"5C",X"EC",X"CD",X"4E",X"F2",X"CD",X"49",X"F1",X"CD",X"D3",X"EA",
		X"20",X"EF",X"21",X"5E",X"EC",X"0E",X"04",X"CD",X"FE",X"EA",X"CD",X"12",X"EB",X"21",X"69",X"EC",
		X"CD",X"4E",X"F2",X"CD",X"1E",X"F1",X"FE",X"01",X"28",X"5F",X"FE",X"03",X"20",X"F5",X"21",X"7D",
		X"EC",X"0E",X"0C",X"CD",X"FE",X"EA",X"CD",X"82",X"F2",X"21",X"8A",X"EC",X"CD",X"4E",X"F2",X"CD",
		X"49",X"F1",X"CD",X"D3",X"EA",X"20",X"F8",X"CD",X"12",X"EB",X"CD",X"82",X"F2",X"21",X"93",X"EC",
		X"CD",X"4E",X"F2",X"CD",X"49",X"F1",X"3A",X"04",X"F8",X"CD",X"DD",X"EA",X"20",X"F5",X"38",X"26",
		X"21",X"22",X"EC",X"0E",X"04",X"CD",X"FE",X"EA",X"CD",X"12",X"EB",X"21",X"A9",X"EC",X"CD",X"4E",
		X"F2",X"CD",X"49",X"F1",X"CD",X"DD",X"EA",X"20",X"F8",X"38",X"0B",X"21",X"2F",X"EC",X"0E",X"04",
		X"CD",X"FE",X"EA",X"CD",X"12",X"EB",X"C3",X"99",X"E8",X"21",X"6B",X"EC",X"0E",X"0A",X"CD",X"FE",
		X"EA",X"CD",X"04",X"E3",X"18",X"B4",X"21",X"52",X"EB",X"0E",X"0A",X"CD",X"FE",X"EA",X"CD",X"75",
		X"E2",X"CD",X"04",X"E3",X"C3",X"19",X"E9",X"21",X"5D",X"EB",X"0E",X"07",X"CD",X"FE",X"EA",X"CD",
		X"75",X"E2",X"CD",X"04",X"E3",X"CD",X"82",X"F2",X"21",X"8A",X"EC",X"CD",X"4E",X"F2",X"CD",X"49",
		X"F1",X"CD",X"D3",X"EA",X"20",X"F8",X"21",X"7D",X"EC",X"01",X"0C",X"00",X"CD",X"FE",X"EA",X"CD",
		X"12",X"EB",X"C3",X"EA",X"E1",X"21",X"CD",X"EB",X"CD",X"4E",X"F2",X"CD",X"1E",X"F1",X"FE",X"07",
		X"28",X"1A",X"FE",X"06",X"28",X"23",X"FE",X"05",X"28",X"2C",X"FE",X"04",X"28",X"35",X"FE",X"03",
		X"28",X"3E",X"FE",X"02",X"28",X"47",X"FE",X"01",X"28",X"50",X"18",X"D9",X"3E",X"00",X"01",X"09",
		X"00",X"11",X"0B",X"EC",X"21",X"00",X"08",X"18",X"4C",X"3E",X"32",X"01",X"06",X"00",X"11",X"02",
		X"EC",X"21",X"20",X"00",X"18",X"3F",X"3E",X"34",X"01",X"06",X"00",X"11",X"F8",X"EB",X"21",X"00",
		X"02",X"18",X"32",X"3E",X"54",X"01",X"04",X"00",X"11",X"EE",X"EB",X"21",X"00",X"10",X"18",X"25",
		X"3E",X"54",X"01",X"04",X"10",X"11",X"E4",X"EB",X"21",X"00",X"20",X"18",X"18",X"3E",X"49",X"01",
		X"04",X"00",X"11",X"DA",X"EB",X"21",X"00",X"10",X"18",X"0B",X"3E",X"49",X"01",X"04",X"10",X"11",
		X"D0",X"EB",X"21",X"00",X"20",X"32",X"41",X"E0",X"22",X"45",X"E0",X"21",X"40",X"E0",X"70",X"EB",
		X"CD",X"FE",X"EA",X"C9",X"11",X"FF",X"FF",X"2A",X"5D",X"E0",X"73",X"23",X"72",X"23",X"22",X"5D",
		X"E0",X"21",X"03",X"E0",X"34",X"C9",X"21",X"00",X"00",X"22",X"4D",X"E0",X"7D",X"32",X"3F",X"E0",
		X"2A",X"05",X"E0",X"22",X"49",X"E0",X"22",X"4F",X"E0",X"3A",X"03",X"E0",X"C9",X"CD",X"33",X"E3",
		X"C3",X"B8",X"E3",X"CD",X"16",X"E3",X"FE",X"01",X"20",X"23",X"2A",X"49",X"E0",X"11",X"00",X"E0",
		X"CD",X"62",X"E0",X"38",X"07",X"21",X"FF",X"FF",X"22",X"49",X"E0",X"23",X"EB",X"2A",X"45",X"E0",
		X"22",X"47",X"E0",X"2B",X"19",X"22",X"4B",X"E0",X"3E",X"01",X"D8",X"AF",X"C9",X"FE",X"02",X"20",
		X"21",X"EB",X"2A",X"07",X"E0",X"22",X"4B",X"E0",X"CD",X"68",X"E0",X"38",X"EB",X"22",X"47",X"E0",
		X"EB",X"2A",X"45",X"E0",X"1B",X"CD",X"62",X"E0",X"3E",X"00",X"30",X"01",X"3C",X"32",X"3F",X"E0",
		X"AF",X"C9",X"EB",X"2A",X"07",X"E0",X"22",X"4B",X"E0",X"CD",X"68",X"E0",X"38",X"CA",X"22",X"47",
		X"E0",X"2A",X"09",X"E0",X"22",X"4D",X"E0",X"EB",X"2A",X"45",X"E0",X"2B",X"CD",X"62",X"E0",X"3E",
		X"01",X"38",X"DA",X"2A",X"47",X"E0",X"19",X"EB",X"2A",X"45",X"E0",X"CD",X"62",X"E0",X"3E",X"00",
		X"30",X"CB",X"3C",X"18",X"C8",X"CD",X"92",X"E4",X"A7",X"C0",X"21",X"05",X"E0",X"06",X"3A",X"36",
		X"00",X"23",X"10",X"FB",X"3A",X"3F",X"E0",X"A7",X"28",X"2E",X"2A",X"45",X"E0",X"11",X"00",X"10",
		X"CD",X"62",X"E0",X"3E",X"00",X"30",X"61",X"ED",X"5B",X"45",X"E0",X"2A",X"47",X"E0",X"2B",X"CD",
		X"62",X"E0",X"D2",X"F9",X"E4",X"44",X"4D",X"2A",X"4D",X"E0",X"09",X"DA",X"58",X"E3",X"CD",X"62",
		X"E0",X"3E",X"01",X"D0",X"AF",X"32",X"3F",X"E0",X"D5",X"2A",X"45",X"E0",X"11",X"00",X"10",X"CD",
		X"62",X"E0",X"D1",X"21",X"56",X"E0",X"3E",X"01",X"38",X"02",X"3E",X"07",X"77",X"01",X"05",X"E0",
		X"2A",X"47",X"E0",X"CD",X"72",X"E0",X"2A",X"4D",X"E0",X"CD",X"72",X"E0",X"EB",X"2A",X"45",X"E0",
		X"19",X"22",X"4D",X"E0",X"2A",X"49",X"E0",X"CD",X"72",X"E0",X"2A",X"4F",X"E0",X"CD",X"72",X"E0",
		X"21",X"56",X"E0",X"35",X"20",X"DA",X"AF",X"C9",X"01",X"05",X"E0",X"ED",X"5B",X"45",X"E0",X"2A",
		X"4D",X"E0",X"A7",X"ED",X"52",X"30",X"FC",X"7D",X"2F",X"5F",X"7C",X"2F",X"57",X"13",X"2A",X"47",
		X"E0",X"CD",X"62",X"E0",X"F5",X"28",X"08",X"38",X"06",X"ED",X"52",X"22",X"47",X"E0",X"EB",X"CD",
		X"72",X"E0",X"EB",X"2A",X"4D",X"E0",X"CD",X"72",X"E0",X"19",X"22",X"4D",X"E0",X"2A",X"49",X"E0",
		X"CD",X"72",X"E0",X"CD",X"6D",X"E0",X"28",X"01",X"19",X"22",X"49",X"E0",X"2A",X"4F",X"E0",X"CD",
		X"72",X"E0",X"CD",X"6D",X"E0",X"28",X"01",X"19",X"22",X"4F",X"E0",X"F1",X"3E",X"00",X"C8",X"30",
		X"AA",X"C9",X"CD",X"16",X"E3",X"11",X"FF",X"FF",X"ED",X"53",X"4F",X"E0",X"FE",X"01",X"20",X"0C",
		X"11",X"00",X"E0",X"CD",X"62",X"E0",X"DA",X"4C",X"E3",X"3E",X"01",X"C9",X"47",X"11",X"00",X"E0",
		X"CD",X"62",X"E0",X"38",X"07",X"21",X"FF",X"FF",X"22",X"49",X"E0",X"23",X"78",X"FE",X"02",X"EB",
		X"2A",X"07",X"E0",X"22",X"4F",X"E0",X"CA",X"4D",X"E3",X"2A",X"09",X"E0",X"22",X"4D",X"E0",X"3E",
		X"01",X"32",X"3F",X"E0",X"78",X"FE",X"03",X"CA",X"4D",X"E3",X"EB",X"2A",X"0B",X"E0",X"CD",X"68",
		X"E0",X"DA",X"58",X"E3",X"22",X"47",X"E0",X"EB",X"2A",X"49",X"E0",X"CD",X"6D",X"E0",X"C8",X"19",
		X"22",X"4B",X"E0",X"11",X"00",X"E0",X"CD",X"62",X"E0",X"3E",X"01",X"D0",X"AF",X"C9",X"3A",X"41",
		X"E0",X"FE",X"32",X"28",X"04",X"FE",X"34",X"20",X"03",X"AF",X"18",X"10",X"A7",X"20",X"04",X"3E",
		X"10",X"18",X"09",X"06",X"30",X"FE",X"49",X"28",X"02",X"06",X"20",X"78",X"32",X"43",X"E0",X"C9",
		X"3A",X"3F",X"E0",X"A7",X"28",X"14",X"21",X"07",X"E0",X"7E",X"23",X"66",X"6F",X"ED",X"5B",X"45",
		X"E0",X"06",X"FF",X"A7",X"ED",X"52",X"04",X"30",X"FA",X"78",X"32",X"51",X"E0",X"C9",X"CD",X"5E",
		X"E5",X"D5",X"11",X"10",X"27",X"1B",X"7A",X"B3",X"20",X"FB",X"D1",X"C9",X"11",X"C0",X"C0",X"3A",
		X"43",X"E0",X"E6",X"30",X"FE",X"20",X"30",X"03",X"50",X"18",X"01",X"58",X"B2",X"C9",X"F5",X"32",
		X"44",X"E0",X"06",X"82",X"FE",X"00",X"20",X"02",X"06",X"80",X"78",X"D3",X"03",X"F1",X"E6",X"C0",
		X"47",X"D5",X"CD",X"4C",X"E5",X"D3",X"02",X"3A",X"3F",X"E0",X"A7",X"3E",X"0E",X"28",X"01",X"AF",
		X"47",X"3A",X"40",X"E0",X"E6",X"10",X"B0",X"32",X"40",X"E0",X"B3",X"D3",X"05",X"D1",X"C9",X"3A",
		X"44",X"E0",X"E6",X"C0",X"47",X"D5",X"CD",X"4C",X"E5",X"47",X"7C",X"E6",X"0F",X"B0",X"D3",X"02",
		X"7D",X"D3",X"00",X"3A",X"40",X"E0",X"E6",X"0E",X"FE",X"0E",X"7C",X"28",X"17",X"E6",X"F0",X"47",
		X"3A",X"43",X"E0",X"E6",X"20",X"28",X"0A",X"3A",X"40",X"E0",X"E6",X"10",X"20",X"03",X"78",X"17",
		X"47",X"78",X"18",X"04",X"E6",X"10",X"F6",X"E0",X"0F",X"0F",X"0F",X"0F",X"47",X"3A",X"40",X"E0",
		X"E6",X"10",X"B0",X"E6",X"1F",X"32",X"40",X"E0",X"B3",X"D1",X"D3",X"05",X"C9",X"D5",X"C5",X"06",
		X"80",X"CD",X"4C",X"E5",X"47",X"7C",X"E6",X"0F",X"B0",X"D3",X"02",X"47",X"3A",X"40",X"E0",X"B3",
		X"D3",X"05",X"4F",X"ED",X"5B",X"58",X"E0",X"1B",X"7A",X"B3",X"20",X"FB",X"78",X"CD",X"0B",X"E6",
		X"D3",X"02",X"79",X"CD",X"0B",X"E6",X"D3",X"05",X"C1",X"D1",X"C9",X"CB",X"77",X"C0",X"E6",X"7F",
		X"C9",X"21",X"05",X"E0",X"4E",X"23",X"46",X"23",X"5E",X"23",X"56",X"23",X"7E",X"23",X"66",X"6F",
		X"EB",X"C9",X"3A",X"03",X"E0",X"FE",X"03",X"3E",X"00",X"C8",X"D5",X"E5",X"2A",X"45",X"E0",X"11",
		X"00",X"10",X"CD",X"62",X"E0",X"E1",X"D1",X"01",X"01",X"01",X"38",X"02",X"0E",X"07",X"C5",X"3E",
		X"40",X"CD",X"3E",X"E5",X"3A",X"40",X"E0",X"E6",X"10",X"32",X"40",X"E0",X"11",X"00",X"00",X"C1",
		X"3E",X"00",X"F5",X"C5",X"D5",X"CD",X"8B",X"E6",X"D1",X"C1",X"28",X"01",X"C5",X"04",X"0D",X"28",
		X"07",X"2A",X"45",X"E0",X"19",X"EB",X"18",X"EB",X"3E",X"C0",X"CD",X"3E",X"E5",X"F1",X"A7",X"C8",
		X"CD",X"DB",X"E7",X"21",X"C5",X"EC",X"CD",X"52",X"F2",X"F1",X"A7",X"28",X"0B",X"CD",X"DB",X"E7",
		X"21",X"C5",X"EC",X"CD",X"52",X"F2",X"18",X"F1",X"3E",X"80",X"C9",X"ED",X"4B",X"45",X"E0",X"EB",
		X"50",X"59",X"CD",X"8F",X"E5",X"23",X"3A",X"43",X"E0",X"E6",X"30",X"06",X"FF",X"20",X"01",X"04",
		X"DB",X"01",X"B8",X"C0",X"1B",X"7A",X"B3",X"20",X"E9",X"C9",X"3E",X"C0",X"CD",X"3E",X"E5",X"3E",
		X"40",X"CD",X"3E",X"E5",X"3A",X"40",X"E0",X"E6",X"10",X"32",X"40",X"E0",X"AF",X"32",X"5B",X"E0",
		X"21",X"00",X"00",X"22",X"56",X"E0",X"22",X"52",X"E0",X"21",X"51",X"E0",X"34",X"2A",X"4B",X"E0",
		X"7E",X"4F",X"23",X"B6",X"F5",X"3E",X"C0",X"CC",X"3E",X"E5",X"F1",X"C8",X"46",X"23",X"EB",X"CD",
		X"79",X"E0",X"22",X"4D",X"E0",X"13",X"CD",X"79",X"E0",X"22",X"49",X"E0",X"13",X"CD",X"79",X"E0",
		X"22",X"4F",X"E0",X"13",X"EB",X"22",X"4B",X"E0",X"C5",X"2A",X"4D",X"E0",X"CD",X"8F",X"E5",X"EB",
		X"2A",X"49",X"E0",X"CD",X"6D",X"E0",X"DB",X"01",X"28",X"0D",X"47",X"3A",X"54",X"E0",X"A7",X"78",
		X"28",X"05",X"77",X"23",X"22",X"49",X"E0",X"21",X"5B",X"E0",X"FE",X"FF",X"28",X"05",X"35",X"28",
		X"01",X"34",X"34",X"F5",X"2A",X"52",X"E0",X"85",X"6F",X"7C",X"CE",X"00",X"67",X"22",X"52",X"E0",
		X"F1",X"2A",X"4F",X"E0",X"BE",X"C4",X"19",X"E8",X"C1",X"28",X"04",X"AF",X"32",X"55",X"E0",X"2A",
		X"4D",X"E0",X"23",X"22",X"4D",X"E0",X"2A",X"4F",X"E0",X"CD",X"6D",X"E0",X"28",X"04",X"23",X"22",
		X"4F",X"E0",X"0B",X"78",X"B1",X"20",X"A1",X"3E",X"C0",X"CD",X"3E",X"E5",X"3A",X"5C",X"E0",X"A7",
		X"20",X"05",X"3A",X"5B",X"E0",X"A7",X"C0",X"F5",X"F5",X"CD",X"D8",X"E7",X"F1",X"21",X"BF",X"EC",
		X"CC",X"52",X"F2",X"F1",X"C8",X"3A",X"61",X"E0",X"A7",X"28",X"2B",X"06",X"02",X"CD",X"3D",X"F3",
		X"CD",X"B6",X"F2",X"06",X"02",X"CD",X"3D",X"F3",X"CD",X"B6",X"F2",X"06",X"02",X"CD",X"3D",X"F3",
		X"CD",X"B6",X"F2",X"AF",X"32",X"61",X"E0",X"0E",X"80",X"CD",X"80",X"F3",X"0E",X"80",X"CD",X"80",
		X"F3",X"0E",X"80",X"CD",X"80",X"F3",X"CD",X"D8",X"E7",X"CD",X"0C",X"F2",X"2A",X"4F",X"E0",X"CD",
		X"6D",X"E0",X"28",X"12",X"2A",X"56",X"E0",X"7C",X"B5",X"28",X"0B",X"21",X"CE",X"EC",X"CD",X"55",
		X"F2",X"2A",X"56",X"E0",X"18",X"09",X"21",X"D3",X"EC",X"CD",X"55",X"F2",X"2A",X"52",X"E0",X"CD",
		X"E6",X"E7",X"2A",X"56",X"E0",X"7C",X"B5",X"C9",X"3A",X"51",X"E0",X"47",X"3E",X"F8",X"C6",X"0A",
		X"10",X"FC",X"57",X"1E",X"11",X"C9",X"7C",X"F5",X"0F",X"0F",X"0F",X"0F",X"CD",X"0D",X"E8",X"CD",
		X"2A",X"F2",X"F1",X"CD",X"0D",X"E8",X"CD",X"2A",X"F2",X"7D",X"F5",X"0F",X"0F",X"0F",X"0F",X"CD",
		X"0D",X"E8",X"CD",X"2A",X"F2",X"F1",X"CD",X"0D",X"E8",X"CD",X"2A",X"F2",X"C9",X"E6",X"0F",X"FE",
		X"0A",X"30",X"03",X"F6",X"30",X"C9",X"C6",X"37",X"C9",X"4F",X"2A",X"4F",X"E0",X"CD",X"6D",X"E0",
		X"C8",X"2A",X"56",X"E0",X"23",X"22",X"56",X"E0",X"3A",X"55",X"E0",X"A7",X"C8",X"C5",X"3E",X"01",
		X"32",X"61",X"E0",X"3A",X"FE",X"FE",X"FE",X"12",X"38",X"23",X"CD",X"49",X"F1",X"C1",X"3A",X"04",
		X"F8",X"FE",X"0D",X"28",X"52",X"C5",X"AF",X"32",X"FE",X"FE",X"21",X"D8",X"EC",X"CD",X"72",X"F1",
		X"3A",X"51",X"E0",X"F6",X"30",X"CD",X"B8",X"F2",X"CD",X"B6",X"F2",X"18",X"0A",X"2B",X"7C",X"B5",
		X"20",X"05",X"CD",X"B6",X"F2",X"18",X"E3",X"06",X"02",X"CD",X"3D",X"F3",X"2A",X"4D",X"E0",X"CD",
		X"20",X"F3",X"06",X"02",X"CD",X"3D",X"F3",X"C1",X"79",X"CD",X"25",X"F3",X"06",X"03",X"CD",X"3D",
		X"F3",X"2A",X"4F",X"E0",X"7E",X"F5",X"CD",X"20",X"F3",X"06",X"02",X"CD",X"3D",X"F3",X"F1",X"CD",
		X"25",X"F3",X"CD",X"B6",X"F2",X"AF",X"C9",X"A7",X"C9",X"CD",X"B5",X"E3",X"A7",X"C0",X"CD",X"FE",
		X"E4",X"11",X"11",X"01",X"CD",X"85",X"F2",X"11",X"12",X"01",X"CD",X"85",X"F2",X"3E",X"01",X"32",
		X"5C",X"E0",X"32",X"54",X"E0",X"32",X"55",X"E0",X"21",X"05",X"E0",X"22",X"4B",X"E0",X"CD",X"20",
		X"E5",X"3A",X"3F",X"E0",X"A7",X"28",X"0C",X"2A",X"4B",X"E0",X"7E",X"23",X"B6",X"C8",X"CD",X"AA",
		X"E6",X"18",X"F4",X"06",X"07",X"D5",X"E5",X"2A",X"45",X"E0",X"11",X"00",X"10",X"CD",X"62",X"E0",
		X"E1",X"D1",X"30",X"02",X"06",X"01",X"C5",X"AF",X"32",X"5C",X"E0",X"32",X"54",X"E0",X"32",X"55",
		X"E0",X"CD",X"AA",X"E6",X"3A",X"5B",X"E0",X"A7",X"28",X"1A",X"32",X"5C",X"E0",X"32",X"54",X"E0",
		X"32",X"55",X"E0",X"2A",X"4B",X"E0",X"11",X"F8",X"FF",X"19",X"22",X"4B",X"E0",X"21",X"51",X"E0",
		X"35",X"CD",X"AA",X"E6",X"C1",X"10",X"CF",X"AF",X"C9",X"CD",X"2D",X"E3",X"A7",X"C0",X"CD",X"FE",
		X"E4",X"11",X"11",X"01",X"CD",X"85",X"F2",X"11",X"12",X"01",X"CD",X"85",X"F2",X"CD",X"22",X"E6",
		X"A7",X"C0",X"21",X"F9",X"EC",X"3A",X"03",X"E0",X"FE",X"03",X"C4",X"4E",X"F2",X"2A",X"49",X"E0",
		X"CD",X"6D",X"E0",X"3E",X"00",X"C8",X"2A",X"45",X"E0",X"11",X"00",X"08",X"CD",X"62",X"E0",X"D2",
		X"DA",X"E9",X"21",X"0E",X"00",X"22",X"58",X"E0",X"CD",X"11",X"E6",X"C5",X"3E",X"C0",X"CD",X"3E",
		X"E5",X"C1",X"CD",X"86",X"E9",X"23",X"13",X"0B",X"78",X"B1",X"20",X"F6",X"AF",X"32",X"54",X"E0",
		X"3C",X"32",X"55",X"E0",X"32",X"5C",X"E0",X"21",X"05",X"E0",X"22",X"4B",X"E0",X"AF",X"32",X"51",
		X"E0",X"CD",X"AA",X"E6",X"AF",X"C9",X"C5",X"1A",X"D5",X"5F",X"06",X"08",X"0E",X"01",X"7B",X"A1",
		X"57",X"28",X"2A",X"C5",X"D5",X"1E",X"05",X"3E",X"00",X"CD",X"5E",X"E5",X"CD",X"8F",X"E5",X"AF",
		X"D3",X"01",X"CD",X"C9",X"E9",X"7A",X"D3",X"01",X"CD",X"DD",X"E5",X"3E",X"40",X"CD",X"5E",X"E5",
		X"CD",X"8F",X"E5",X"DB",X"01",X"AA",X"28",X"03",X"1D",X"20",X"DC",X"D1",X"C1",X"79",X"07",X"4F",
		X"CD",X"CF",X"E9",X"05",X"20",X"C8",X"D1",X"C1",X"C9",X"D5",X"11",X"14",X"00",X"18",X"04",X"D5",
		X"11",X"1E",X"00",X"1B",X"7B",X"B2",X"20",X"FB",X"D1",X"C9",X"21",X"05",X"E0",X"22",X"4B",X"E0",
		X"CD",X"20",X"E5",X"3A",X"3F",X"E0",X"A7",X"CA",X"47",X"EA",X"3E",X"05",X"32",X"5A",X"E0",X"21",
		X"94",X"03",X"22",X"58",X"E0",X"2A",X"4B",X"E0",X"7E",X"4F",X"23",X"B6",X"C8",X"46",X"2B",X"E5",
		X"00",X"00",X"00",X"01",X"C0",X"00",X"04",X"00",X"C4",X"00",X"01",X"D0",X"C5",X"D0",X"09",X"90",
		X"CF",X"50",X"02",X"80",X"D1",X"D0",X"01",X"A0",X"D3",X"70",X"01",X"F0",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",
		X"F4",X"12",X"F4",X"3F",X"F4",X"59",X"F4",X"76",X"F5",X"33",X"F5",X"E1",X"F8",X"07",X"F8",X"18",
		X"F8",X"33",X"F8",X"48",X"F8",X"5D",X"F8",X"72",X"F8",X"87",X"F8",X"99",X"F8",X"AE",X"F8",X"D6",
		X"EA",X"80",X"EA",X"F5",X"EB",X"6A",X"EC",X"01",X"EC",X"7B",X"ED",X"75",X"EE",X"31",X"F2",X"15",
		X"66",X"B8",X"40",X"77",X"41",X"00",X"42",X"8E",X"43",X"00",X"45",X"00",X"6C",X"14",X"6D",X"14",
		X"6E",X"14",X"68",X"0A",X"69",X"0A",X"6A",X"0A",X"04",X"EE",X"20",X"40",X"6A",X"42",X"7E",X"68",
		X"0A",X"69",X"0A",X"6A",X"0A",X"04",X"D4",X"20",X"68",X"0A",X"69",X"0A",X"6A",X"0A",X"04",X"D4",
		X"20",X"40",X"4F",X"42",X"5E",X"68",X"0A",X"69",X"0A",X"6A",X"0A",X"04",X"9F",X"40",X"40",X"59",
		X"42",X"6A",X"68",X"0A",X"69",X"0A",X"6A",X"0A",X"04",X"B3",X"40",X"40",X"5E",X"42",X"77",X"68",
		X"0A",X"69",X"0A",X"6A",X"0A",X"04",X"BD",X"40",X"40",X"6A",X"42",X"7E",X"68",X"0A",X"69",X"0A",
		X"6A",X"0A",X"04",X"D4",X"20",X"40",X"5E",X"42",X"77",X"68",X"0A",X"69",X"0A",X"6A",X"0A",X"04",
		X"BD",X"60",X"67",X"07",X"FF",X"66",X"BC",X"40",X"7A",X"41",X"01",X"43",X"00",X"6C",X"14",X"6D",
		X"14",X"6E",X"14",X"68",X"0A",X"69",X"0A",X"02",X"BD",X"24",X"40",X"3E",X"68",X"0A",X"69",X"0A",
		X"02",X"9F",X"24",X"40",X"1C",X"68",X"0A",X"69",X"0A",X"02",X"6A",X"24",X"40",X"3E",X"68",X"0A",
		X"69",X"0A",X"02",X"77",X"24",X"42",X"7E",X"49",X"0A",X"68",X"0A",X"00",X"7E",X"24",X"68",X"0A",
		X"00",X"3E",X"24",X"42",X"77",X"49",X"0A",X"68",X"0A",X"00",X"1C",X"24",X"68",X"0A",X"00",X"3E",
		X"24",X"49",X"00",X"42",X"5E",X"68",X"0A",X"69",X"0A",X"00",X"7A",X"24",X"42",X"9F",X"68",X"0A",
		X"69",X"0A",X"00",X"DD",X"24",X"42",X"8E",X"68",X"0A",X"69",X"0A",X"00",X"A9",X"24",X"42",X"77",
		X"68",X"0A",X"69",X"0A",X"00",X"DD",X"64",X"67",X"03",X"FF",X"66",X"BC",X"6C",X"14",X"6D",X"14",
		X"6E",X"14",X"FE",X"EB",X"8D",X"FE",X"EB",X"8D",X"FE",X"EB",X"C6",X"FE",X"EB",X"C6",X"FE",X"EB",
		X"8D",X"FE",X"EB",X"8D",X"FE",X"EB",X"C6",X"FE",X"EB",X"C6",X"67",X"03",X"FF",X"41",X"00",X"43",
		X"00",X"42",X"EE",X"68",X"0A",X"69",X"0A",X"00",X"77",X"22",X"68",X"0A",X"69",X"0A",X"00",X"5E",
		X"22",X"68",X"0A",X"69",X"0A",X"00",X"59",X"22",X"42",X"3E",X"43",X"01",X"68",X"0A",X"69",X"0A",
		X"00",X"4F",X"22",X"42",X"1C",X"68",X"0A",X"69",X"0A",X"00",X"59",X"22",X"42",X"3E",X"68",X"0A",
		X"69",X"0A",X"00",X"4F",X"22",X"FD",X"43",X"00",X"42",X"D4",X"68",X"0A",X"69",X"0A",X"00",X"6A",
		X"22",X"68",X"0A",X"69",X"0A",X"00",X"59",X"22",X"68",X"0A",X"69",X"0A",X"00",X"4F",X"22",X"43",
		X"01",X"42",X"1C",X"68",X"0A",X"69",X"0A",X"00",X"47",X"22",X"43",X"00",X"42",X"FD",X"68",X"0A",
		X"69",X"0A",X"00",X"4F",X"22",X"43",X"01",X"42",X"1C",X"68",X"0A",X"69",X"0A",X"00",X"47",X"22",
		X"FD",X"67",X"BF",X"66",X"BC",X"41",X"00",X"40",X"1C",X"43",X"00",X"44",X"00",X"45",X"00",X"6C",
		X"14",X"6D",X"14",X"6E",X"14",X"68",X"0A",X"69",X"0A",X"02",X"8E",X"18",X"40",X"FD",X"41",X"00",
		X"68",X"0A",X"69",X"0A",X"02",X"7E",X"18",X"40",X"EE",X"68",X"0A",X"69",X"0A",X"02",X"77",X"18",
		X"40",X"D4",X"68",X"0A",X"69",X"0A",X"02",X"6A",X"18",X"40",X"BD",X"68",X"0A",X"69",X"0A",X"02",
		X"5E",X"18",X"40",X"FD",X"68",X"0A",X"69",X"0A",X"02",X"7E",X"18",X"40",X"EE",X"68",X"0A",X"69",
		X"0A",X"02",X"77",X"18",X"40",X"D4",X"68",X"0A",X"69",X"0A",X"02",X"6A",X"18",X"40",X"BD",X"68",
		X"0A",X"69",X"0A",X"02",X"5E",X"18",X"40",X"A8",X"68",X"0A",X"69",X"0A",X"02",X"54",X"18",X"40",
		X"9F",X"68",X"0A",X"69",X"0A",X"02",X"4F",X"18",X"67",X"03",X"FF",X"66",X"B8",X"40",X"47",X"41",
		X"00",X"42",X"B3",X"43",X"00",X"45",X"01",X"6C",X"14",X"6D",X"14",X"6E",X"14",X"68",X"0A",X"69",
		X"0A",X"6A",X"0A",X"04",X"65",X"20",X"40",X"59",X"42",X"8F",X"68",X"0A",X"69",X"0A",X"6A",X"0A",
		X"04",X"65",X"20",X"40",X"4F",X"42",X"77",X"68",X"0A",X"69",X"0A",X"6A",X"0A",X"04",X"65",X"20",
		X"40",X"59",X"42",X"6A",X"45",X"00",X"68",X"0A",X"69",X"0A",X"6A",X"0A",X"04",X"00",X"20",X"40",
		X"00",X"42",X"59",X"68",X"0A",X"69",X"0A",X"6A",X"0A",X"04",X"00",X"20",X"40",X"59",X"42",X"6A",
		X"45",X"01",X"68",X"0A",X"69",X"0A",X"6A",X"0A",X"04",X"1C",X"20",X"40",X"4F",X"42",X"77",X"45",
		X"00",X"68",X"0A",X"69",X"0A",X"6A",X"0A",X"04",X"00",X"20",X"40",X"59",X"42",X"6A",X"68",X"0A",
		X"69",X"0A",X"6A",X"0A",X"04",X"EE",X"20",X"40",X"47",X"42",X"B3",X"45",X"01",X"68",X"0A",X"69",
		X"0A",X"6A",X"0A",X"04",X"65",X"20",X"40",X"59",X"42",X"8E",X"68",X"0A",X"69",X"0A",X"6A",X"0A",
		X"04",X"65",X"20",X"40",X"4F",X"42",X"77",X"68",X"0A",X"69",X"0A",X"6A",X"0A",X"04",X"65",X"20",
		X"40",X"59",X"42",X"6A",X"45",X"00",X"68",X"0A",X"69",X"0A",X"04",X"00",X"20",X"40",X"00",X"42",
		X"59",X"68",X"0A",X"69",X"0A",X"04",X"00",X"20",X"40",X"59",X"42",X"6A",X"45",X"01",X"68",X"0A",
		X"69",X"0A",X"6A",X"0A",X"04",X"1C",X"20",X"40",X"4F",X"42",X"77",X"45",X"00",X"68",X"0A",X"69",
		X"0A",X"6A",X"0A",X"04",X"00",X"20",X"40",X"59",X"42",X"6A",X"68",X"0A",X"69",X"0A",X"6A",X"0A",
		X"04",X"EE",X"20",X"40",X"47",X"42",X"59",X"45",X"01",X"68",X"0A",X"69",X"0A",X"6A",X"0A",X"04",
		X"65",X"60",X"67",X"07",X"FF",X"66",X"BC",X"40",X"BD",X"41",X"00",X"43",X"00",X"48",X"0A",X"69",
		X"0A",X"02",X"77",X"16",X"02",X"00",X"16",X"40",X"B3",X"48",X"0A",X"69",X"0A",X"02",X"8E",X"16",
		X"02",X"00",X"16",X"48",X"00",X"49",X"0A",X"42",X"9F",X"68",X"0A",X"00",X"9F",X"2C",X"68",X"0A",
		X"00",X"8E",X"2C",X"49",X"00",X"40",X"BD",X"48",X"0A",X"69",X"0A",X"02",X"77",X"16",X"02",X"00",
		X"16",X"40",X"9F",X"48",X"0A",X"69",X"0A",X"02",X"8E",X"16",X"02",X"00",X"16",X"48",X"00",X"42",
		X"9F",X"49",X"0A",X"68",X"0A",X"00",X"9F",X"2C",X"68",X"0A",X"00",X"8E",X"2C",X"49",X"00",X"40",
		X"BD",X"68",X"0A",X"69",X"0A",X"02",X"8E",X"2C",X"40",X"9F",X"68",X"0A",X"69",X"0A",X"02",X"7E",
		X"2C",X"40",X"B3",X"68",X"0A",X"69",X"0A",X"02",X"77",X"2C",X"40",X"D4",X"68",X"0A",X"79",X"0D",
		X"02",X"6A",X"2C",X"40",X"EE",X"68",X"0A",X"69",X"0A",X"02",X"77",X"58",X"67",X"03",X"FF",X"66",
		X"B7",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"48",X"10",X"06",X"01",X"28",X"48",X"00",X"06",X"00",
		X"28",X"48",X"10",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"06",X"01",X"28",X"48",X"00",X"06",X"00",
		X"28",X"48",X"10",X"4B",X"03",X"4C",X"02",X"4D",X"09",X"06",X"01",X"28",X"48",X"00",X"06",X"01",
		X"28",X"4B",X"00",X"4C",X"00",X"4D",X"00",X"66",X"B7",X"67",X"08",X"66",X"B8",X"6C",X"28",X"6D",
		X"10",X"6E",X"14",X"FE",X"F0",X"19",X"FE",X"F1",X"B3",X"FE",X"F0",X"7D",X"FE",X"F0",X"E5",X"FE",
		X"F0",X"19",X"FE",X"F1",X"B3",X"FE",X"F0",X"7D",X"FE",X"F1",X"4C",X"FE",X"F0",X"19",X"FE",X"F1",
		X"B3",X"FE",X"F0",X"7D",X"FE",X"F0",X"E5",X"FE",X"F0",X"19",X"FE",X"F1",X"B3",X"FE",X"F0",X"7D",
		X"FE",X"F1",X"4C",X"40",X"96",X"48",X"0C",X"43",X"01",X"44",X"3C",X"45",X"00",X"6C",X"28",X"6D",
		X"10",X"6E",X"14",X"69",X"0B",X"6A",X"0A",X"02",X"2C",X"2D",X"44",X"43",X"69",X"0B",X"6A",X"0D",
		X"02",X"2C",X"2D",X"40",X"86",X"44",X"4B",X"48",X"0C",X"69",X"0B",X"6A",X"0A",X"02",X"2C",X"2D",
		X"44",X"43",X"69",X"0B",X"6A",X"0A",X"02",X"2C",X"2D",X"48",X"00",X"40",X"77",X"44",X"3C",X"68",
		X"0C",X"69",X"0B",X"6A",X"0A",X"02",X"0C",X"2D",X"40",X"86",X"44",X"43",X"68",X"0C",X"69",X"0B",
		X"6A",X"0A",X"02",X"2C",X"2D",X"40",X"96",X"44",X"4B",X"68",X"0C",X"69",X"0B",X"6A",X"0A",X"02",
		X"3E",X"2D",X"40",X"77",X"44",X"3C",X"68",X"0C",X"69",X"0B",X"6A",X"0A",X"02",X"2C",X"2D",X"40",
		X"86",X"44",X"43",X"48",X"0C",X"69",X"0B",X"6A",X"0A",X"02",X"0C",X"2D",X"44",X"4B",X"69",X"0B",
		X"6A",X"0A",X"02",X"0C",X"2D",X"48",X"00",X"40",X"B3",X"44",X"4F",X"6A",X"0A",X"68",X"0C",X"69",
		X"0B",X"02",X"65",X"2D",X"40",X"86",X"48",X"0C",X"44",X"4B",X"6A",X"0A",X"69",X"0B",X"02",X"0C",
		X"2D",X"44",X"43",X"69",X"0B",X"6A",X"0A",X"02",X"65",X"2D",X"44",X"4B",X"6A",X"0A",X"69",X"0B",
		X"02",X"3E",X"2D",X"44",X"4F",X"6A",X"0A",X"69",X"0B",X"02",X"2C",X"2D",X"48",X"00",X"43",X"00",
		X"44",X"43",X"6A",X"0A",X"69",X"0B",X"02",X"EE",X"2D",X"40",X"86",X"43",X"01",X"44",X"38",X"48",
		X"0C",X"69",X"0B",X"6A",X"0A",X"02",X"0C",X"2D",X"44",X"3C",X"6A",X"0A",X"69",X"0B",X"02",X"0C",
		X"2D",X"40",X"77",X"44",X"43",X"48",X"0C",X"69",X"0B",X"6A",X"0A",X"02",X"0C",X"2D",X"44",X"3C",
		X"6A",X"0A",X"69",X"0B",X"02",X"0C",X"2D",X"48",X"00",X"40",X"71",X"43",X"00",X"44",X"38",X"6A",
		X"0A",X"68",X"0C",X"69",X"0B",X"02",X"EE",X"2D",X"40",X"77",X"43",X"01",X"44",X"3C",X"6A",X"0A",
		X"68",X"0C",X"69",X"0B",X"02",X"0C",X"2D",X"40",X"86",X"44",X"43",X"6A",X"0A",X"68",X"0C",X"69",
		X"0B",X"02",X"2C",X"2D",X"40",X"96",X"44",X"4B",X"6A",X"0A",X"68",X"0C",X"69",X"0B",X"02",X"0C",
		X"2D",X"40",X"77",X"43",X"00",X"44",X"3C",X"6A",X"0A",X"68",X"0C",X"69",X"0B",X"02",X"EE",X"2D",
		X"40",X"71",X"44",X"38",X"6A",X"0A",X"68",X"0C",X"69",X"0B",X"02",X"EE",X"2D",X"40",X"77",X"44",
		X"3C",X"6A",X"0A",X"68",X"0C",X"69",X"0B",X"02",X"EE",X"2D",X"40",X"86",X"44",X"43",X"6A",X"0A",
		X"68",X"0C",X"69",X"0B",X"02",X"EE",X"2D",X"40",X"77",X"44",X"3C",X"48",X"0C",X"4A",X"0A",X"69",
		X"0B",X"02",X"EE",X"16",X"69",X"0B",X"02",X"E1",X"16",X"48",X"00",X"4A",X"00",X"40",X"86",X"44",
		X"38",X"6A",X"0A",X"68",X"0C",X"69",X"0B",X"02",X"EE",X"2D",X"40",X"96",X"43",X"01",X"44",X"3C",
		X"6A",X"0A",X"68",X"0C",X"69",X"0B",X"02",X"0C",X"2D",X"40",X"9F",X"44",X"43",X"6A",X"0A",X"68",
		X"0C",X"69",X"0B",X"02",X"2C",X"2D",X"FE",X"EE",X"3D",X"40",X"B3",X"48",X"0C",X"43",X"01",X"45",
		X"00",X"69",X"0B",X"02",X"65",X"16",X"43",X"00",X"02",X"00",X"16",X"43",X"01",X"44",X"59",X"6A",
		X"0A",X"69",X"0B",X"02",X"65",X"2D",X"40",X"9F",X"44",X"64",X"48",X"0C",X"69",X"0B",X"6A",X"0A",
		X"02",X"2C",X"2D",X"44",X"59",X"69",X"0B",X"6A",X"0A",X"02",X"65",X"2D",X"48",X"00",X"40",X"96",
		X"68",X"0C",X"69",X"0B",X"02",X"2C",X"2D",X"40",X"9F",X"44",X"4B",X"6A",X"0A",X"68",X"0C",X"69",
		X"0B",X"02",X"3E",X"2D",X"40",X"B3",X"44",X"4F",X"48",X"0C",X"69",X"0B",X"6A",X"0A",X"02",X"65",
		X"2D",X"44",X"4B",X"6A",X"0A",X"69",X"0B",X"02",X"3E",X"2D",X"48",X"00",X"FD",X"40",X"B3",X"48",
		X"0C",X"69",X"0B",X"02",X"65",X"16",X"43",X"00",X"02",X"00",X"16",X"43",X"01",X"44",X"59",X"6A",
		X"0A",X"69",X"0B",X"02",X"65",X"2D",X"40",X"9F",X"44",X"64",X"48",X"0C",X"69",X"0B",X"6A",X"0A",
		X"02",X"2C",X"2D",X"44",X"59",X"69",X"0B",X"6A",X"0A",X"02",X"65",X"2D",X"48",X"00",X"40",X"77",
		X"44",X"59",X"6A",X"0A",X"68",X"0C",X"69",X"0B",X"02",X"0C",X"2D",X"40",X"86",X"43",X"00",X"44",
		X"4F",X"6A",X"0A",X"68",X"0C",X"69",X"0B",X"02",X"EE",X"2D",X"40",X"96",X"43",X"01",X"44",X"4B",
		X"48",X"0C",X"69",X"0B",X"6A",X"0A",X"02",X"0C",X"2D",X"44",X"3C",X"6A",X"0A",X"69",X"0B",X"02",
		X"2C",X"2D",X"48",X"00",X"FD",X"40",X"9F",X"48",X"0C",X"43",X"01",X"44",X"43",X"4A",X"0A",X"69",
		X"0B",X"02",X"90",X"2D",X"69",X"0B",X"02",X"90",X"2D",X"48",X"00",X"4A",X"00",X"40",X"96",X"43",
		X"01",X"44",X"4B",X"6A",X"0A",X"68",X"0C",X"69",X"0B",X"02",X"DD",X"2D",X"40",X"C8",X"43",X"01",
		X"44",X"4F",X"48",X"0C",X"4A",X"0A",X"69",X"0B",X"02",X"90",X"2D",X"69",X"0B",X"02",X"90",X"2D",
		X"48",X"00",X"4A",X"00",X"40",X"B3",X"44",X"4B",X"68",X"0C",X"69",X"0B",X"6A",X"0A",X"02",X"90",
		X"2D",X"40",X"9F",X"43",X"01",X"44",X"43",X"48",X"0C",X"4A",X"0A",X"69",X"0B",X"02",X"DD",X"2D",
		X"43",X"01",X"69",X"0B",X"02",X"90",X"2D",X"48",X"00",X"4A",X"00",X"FD",X"40",X"9F",X"48",X"0C",
		X"43",X"01",X"44",X"43",X"4A",X"0A",X"69",X"0B",X"02",X"90",X"2D",X"69",X"0B",X"02",X"90",X"2D",
		X"48",X"00",X"4A",X"00",X"40",X"96",X"43",X"01",X"44",X"4B",X"68",X"0C",X"69",X"0B",X"6A",X"0A",
		X"02",X"DD",X"2D",X"40",X"86",X"43",X"01",X"44",X"4F",X"4A",X"0A",X"48",X"0C",X"69",X"0B",X"02",
		X"90",X"2D",X"69",X"0B",X"02",X"90",X"2D",X"48",X"00",X"4A",X"00",X"40",X"96",X"44",X"4B",X"6A",
		X"0A",X"68",X"0C",X"69",X"0B",X"02",X"90",X"2D",X"40",X"9F",X"44",X"43",X"48",X"0C",X"4A",X"0A",
		X"43",X"01",X"69",X"0B",X"02",X"DD",X"2D",X"43",X"01",X"69",X"0B",X"02",X"90",X"2D",X"48",X"00",
		X"4A",X"00",X"FD",X"40",X"B3",X"48",X"0C",X"43",X"01",X"69",X"0B",X"02",X"65",X"16",X"43",X"00",
		X"02",X"00",X"16",X"43",X"01",X"44",X"59",X"6A",X"0A",X"69",X"0B",X"02",X"65",X"2D",X"40",X"9F",
		X"44",X"64",X"48",X"0C",X"69",X"0B",X"6A",X"0A",X"02",X"2C",X"2D",X"44",X"59",X"6A",X"0A",X"69",
		X"0B",X"02",X"65",X"2D",X"48",X"00",X"40",X"86",X"68",X"0C",X"69",X"0B",X"02",X"0C",X"2D",X"40",
		X"96",X"44",X"4B",X"6A",X"0A",X"68",X"0C",X"69",X"0B",X"02",X"2C",X"2D",X"40",X"9F",X"44",X"4F",
		X"48",X"0C",X"69",X"0B",X"6A",X"0A",X"02",X"3E",X"2D",X"44",X"4B",X"69",X"0B",X"6A",X"0A",X"02",
		X"2C",X"2D",X"48",X"00",X"FD",X"67",X"BF",X"66",X"B8",X"40",X"77",X"41",X"00",X"42",X"00",X"43",
		X"00",X"45",X"01",X"6C",X"14",X"6D",X"14",X"6E",X"14",X"FE",X"F2",X"AB",X"FE",X"F3",X"C5",X"FE",
		X"F2",X"E8",X"FE",X"F3",X"2F",X"FE",X"F3",X"7E",X"FE",X"F3",X"C5",X"40",X"47",X"42",X"D4",X"68",
		X"0A",X"69",X"0A",X"6A",X"0A",X"04",X"65",X"30",X"40",X"4F",X"42",X"BD",X"68",X"0A",X"69",X"0A",
		X"6A",X"0A",X"04",X"65",X"30",X"40",X"47",X"48",X"0A",X"42",X"B3",X"49",X"0A",X"6A",X"0A",X"04",
		X"65",X"30",X"6A",X"0A",X"04",X"65",X"30",X"48",X"00",X"49",X"00",X"40",X"4F",X"42",X"BD",X"68",
		X"0A",X"69",X"0A",X"6A",X"0A",X"04",X"7A",X"30",X"40",X"59",X"42",X"B3",X"68",X"0A",X"69",X"0A",
		X"6A",X"0A",X"04",X"7A",X"30",X"40",X"6A",X"42",X"8E",X"49",X"0A",X"68",X"0A",X"6A",X"0A",X"04",
		X"A9",X"30",X"40",X"5E",X"68",X"0A",X"69",X"0A",X"04",X"A9",X"30",X"40",X"77",X"42",X"9F",X"68",
		X"0A",X"69",X"0A",X"6A",X"0A",X"04",X"DD",X"C0",X"67",X"07",X"FF",X"68",X"0A",X"69",X"0A",X"6A",
		X"0A",X"04",X"DD",X"30",X"6A",X"0A",X"04",X"DD",X"30",X"40",X"5E",X"68",X"0A",X"6A",X"0A",X"04",
		X"DD",X"30",X"6A",X"0A",X"04",X"DD",X"30",X"40",X"4F",X"68",X"0A",X"6A",X"0A",X"04",X"DD",X"30",
		X"6A",X"0A",X"04",X"DD",X"30",X"40",X"59",X"68",X"0A",X"6A",X"0A",X"04",X"DD",X"30",X"40",X"6A",
		X"68",X"0A",X"6A",X"0A",X"04",X"DD",X"30",X"FD",X"40",X"8E",X"42",X"9F",X"48",X"0A",X"45",X"02",
		X"49",X"0A",X"6A",X"0A",X"04",X"38",X"30",X"6A",X"0A",X"04",X"38",X"30",X"40",X"77",X"48",X"0A",
		X"6A",X"0A",X"04",X"38",X"30",X"6A",X"0A",X"04",X"38",X"30",X"49",X"00",X"40",X"5E",X"48",X"0A",
		X"6A",X"0A",X"04",X"38",X"30",X"6A",X"0A",X"04",X"38",X"30",X"48",X"00",X"40",X"6A",X"68",X"0A",
		X"6A",X"0A",X"04",X"38",X"30",X"40",X"77",X"68",X"0A",X"6A",X"0A",X"04",X"38",X"30",X"FD",X"40",
		X"6A",X"48",X"0A",X"6A",X"0A",X"04",X"38",X"30",X"42",X"9F",X"69",X"0A",X"6A",X"0A",X"04",X"38",
		X"30",X"42",X"B3",X"69",X"0A",X"6A",X"0A",X"04",X"38",X"30",X"48",X"00",X"40",X"8E",X"42",X"BD",
		X"48",X"0A",X"6A",X"0A",X"69",X"0A",X"04",X"38",X"30",X"42",X"B3",X"49",X"0A",X"6A",X"0A",X"04",
		X"38",X"30",X"6A",X"0A",X"04",X"38",X"30",X"49",X"00",X"42",X"BD",X"69",X"0A",X"6A",X"0A",X"04",
		X"38",X"30",X"48",X"00",X"42",X"D4",X"69",X"0A",X"6A",X"0A",X"04",X"38",X"30",X"FD",X"40",X"77",
		X"48",X"0A",X"42",X"BD",X"45",X"01",X"49",X"0A",X"6A",X"0A",X"04",X"DD",X"30",X"6A",X"0A",X"04",
		X"DD",X"30",X"40",X"5E",X"48",X"0A",X"6A",X"0A",X"04",X"DD",X"30",X"6A",X"0A",X"04",X"DD",X"30",
		X"49",X"00",X"40",X"4F",X"48",X"0A",X"6A",X"0A",X"04",X"DD",X"30",X"6A",X"0A",X"04",X"DD",X"30",
		X"48",X"00",X"40",X"59",X"68",X"0A",X"6A",X"0A",X"04",X"DD",X"30",X"40",X"6A",X"68",X"0A",X"6A",
		X"0A",X"04",X"DD",X"30",X"FD",X"48",X"0A",X"40",X"5E",X"6A",X"0A",X"04",X"DD",X"30",X"42",X"EE",
		X"69",X"0A",X"6A",X"0A",X"04",X"DD",X"30",X"42",X"BD",X"69",X"0A",X"6A",X"0A",X"04",X"DD",X"30",
		X"40",X"4F",X"48",X"0A",X"42",X"B3",X"69",X"0A",X"6A",X"0A",X"04",X"DD",X"30",X"42",X"9F",X"49",
		X"0A",X"6A",X"0A",X"04",X"DD",X"30",X"6A",X"0A",X"04",X"DD",X"30",X"49",X"00",X"42",X"B3",X"69",
		X"0A",X"6A",X"0A",X"04",X"DD",X"30",X"48",X"00",X"42",X"D4",X"69",X"0A",X"6A",X"0A",X"04",X"DD",
		X"30",X"FD",X"77",X"BF",X"76",X"BE",X"51",X"00",X"53",X"D4",X"58",X"0A",X"59",X"0A",X"10",X"B3",
		X"1A",X"52",X"B3",X"10",X"8E",X"1A",X"52",X"77",X"10",X"5E",X"40",X"52",X"D4",X"10",X"B3",X"1A",
		X"52",X"B3",X"10",X"8E",X"1A",X"52",X"77",X"10",X"5E",X"60",X"58",X"00",X"77",X"01",X"FF",X"77",
		X"BF",X"76",X"B8",X"50",X"70",X"52",X"6D",X"58",X"10",X"59",X"10",X"5A",X"10",X"5B",X"30",X"5C",
		X"04",X"5D",X"09",X"14",X"78",X"80",X"77",X"07",X"FF",X"76",X"BD",X"53",X"00",X"52",X"43",X"59",
		X"10",X"5B",X"04",X"5C",X"10",X"1D",X"09",X"20",X"52",X"53",X"59",X"10",X"1D",X"09",X"E0",X"52",
		X"00",X"59",X"00",X"77",X"02",X"FF",X"66",X"B8",X"4B",X"00",X"4C",X"00",X"4D",X"00",X"40",X"70",
		X"41",X"00",X"42",X"75",X"43",X"00",X"45",X"00",X"48",X"0A",X"49",X"0A",X"4A",X"0A",X"6C",X"00",
		X"6D",X"00",X"6E",X"00",X"04",X"77",X"10",X"40",X"74",X"42",X"78",X"04",X"7A",X"10",X"40",X"78",
		X"42",X"7C",X"04",X"79",X"10",X"40",X"7B",X"42",X"77",X"04",X"7F",X"10",X"40",X"80",X"42",X"86",
		X"04",X"87",X"10",X"40",X"84",X"42",X"88",X"04",X"8A",X"10",X"40",X"89",X"42",X"8E",X"04",X"8F",
		X"10",X"40",X"90",X"42",X"91",X"04",X"92",X"10",X"40",X"98",X"42",X"99",X"04",X"9A",X"10",X"40",
		X"A0",X"42",X"A1",X"04",X"A2",X"10",X"40",X"A8",X"42",X"A9",X"04",X"AA",X"10",X"40",X"B0",X"42",
		X"B1",X"04",X"B2",X"10",X"40",X"B8",X"42",X"B9",X"04",X"BA",X"10",X"40",X"C0",X"42",X"C1",X"04",
		X"C2",X"10",X"40",X"C8",X"42",X"C9",X"04",X"CA",X"10",X"40",X"D0",X"42",X"D1",X"04",X"D2",X"10",
		X"40",X"D8",X"42",X"D9",X"04",X"DA",X"10",X"40",X"E0",X"42",X"E1",X"04",X"E2",X"10",X"40",X"E8",
		X"42",X"E9",X"04",X"EA",X"10",X"40",X"F0",X"42",X"F1",X"04",X"F2",X"10",X"40",X"F8",X"42",X"F9",
		X"04",X"FA",X"10",X"40",X"FF",X"42",X"FF",X"04",X"FF",X"30",X"48",X"00",X"49",X"00",X"4A",X"00",
		X"67",X"07",X"FF",X"66",X"B8",X"4B",X"00",X"4C",X"00",X"4D",X"00",X"40",X"FF",X"41",X"00",X"42",
		X"FF",X"43",X"00",X"45",X"00",X"48",X"0A",X"49",X"0A",X"4A",X"0A",X"6C",X"00",X"6D",X"00",X"6E",
		X"00",X"04",X"FF",X"10",X"40",X"F8",X"42",X"F9",X"04",X"FA",X"10",X"40",X"F0",X"42",X"F1",X"04",
		X"F2",X"10",X"40",X"E8",X"42",X"E9",X"04",X"EA",X"10",X"40",X"E0",X"42",X"E1",X"04",X"E2",X"10",
		X"40",X"D8",X"42",X"D9",X"04",X"DA",X"10",X"40",X"D0",X"42",X"D1",X"04",X"D2",X"10",X"40",X"C8",
		X"42",X"C9",X"04",X"CA",X"10",X"40",X"C0",X"42",X"C1",X"04",X"C2",X"10",X"40",X"B8",X"42",X"B9",
		X"04",X"BA",X"10",X"40",X"B0",X"42",X"B1",X"04",X"B2",X"10",X"40",X"A8",X"42",X"A9",X"04",X"AA",
		X"10",X"40",X"A0",X"42",X"A1",X"04",X"A2",X"10",X"40",X"9E",X"42",X"9A",X"04",X"98",X"10",X"40",
		X"96",X"42",X"93",X"04",X"94",X"10",X"40",X"8E",X"42",X"8A",X"04",X"88",X"10",X"40",X"87",X"42",
		X"85",X"04",X"83",X"10",X"40",X"7E",X"42",X"77",X"04",X"75",X"10",X"40",X"75",X"42",X"7A",X"04",
		X"70",X"30",X"40",X"00",X"42",X"00",X"44",X"00",X"48",X"00",X"49",X"00",X"4A",X"00",X"67",X"07",
		X"FF",X"76",X"BD",X"50",X"00",X"51",X"00",X"53",X"00",X"59",X"0C",X"58",X"0C",X"12",X"11",X"05",
		X"12",X"12",X"05",X"12",X"13",X"05",X"12",X"14",X"05",X"12",X"15",X"05",X"12",X"16",X"05",X"12",
		X"17",X"05",X"12",X"18",X"05",X"12",X"19",X"05",X"12",X"1A",X"05",X"50",X"16",X"12",X"1B",X"05",
		X"50",X"17",X"12",X"1C",X"05",X"50",X"18",X"12",X"1D",X"05",X"50",X"19",X"12",X"1E",X"05",X"50",
		X"1A",X"12",X"1F",X"05",X"50",X"1B",X"12",X"20",X"05",X"50",X"1C",X"12",X"21",X"05",X"50",X"1D",
		X"12",X"22",X"05",X"50",X"1E",X"12",X"23",X"05",X"50",X"1F",X"12",X"24",X"05",X"12",X"25",X"05",
		X"12",X"26",X"05",X"12",X"27",X"05",X"12",X"28",X"05",X"12",X"29",X"05",X"12",X"2A",X"05",X"50",
		X"26",X"12",X"2B",X"05",X"50",X"27",X"12",X"2C",X"05",X"50",X"28",X"12",X"2D",X"05",X"50",X"29",
		X"12",X"2E",X"05",X"50",X"2A",X"12",X"2F",X"05",X"50",X"2B",X"12",X"30",X"05",X"50",X"2C",X"12",
		X"31",X"05",X"50",X"2D",X"12",X"32",X"05",X"50",X"2E",X"12",X"33",X"05",X"50",X"2F",X"12",X"34",
		X"05",X"12",X"35",X"05",X"12",X"36",X"05",X"12",X"37",X"05",X"12",X"38",X"05",X"12",X"39",X"05",
		X"12",X"3A",X"05",X"50",X"36",X"12",X"3B",X"05",X"50",X"37",X"12",X"3C",X"05",X"50",X"38",X"12",
		X"3D",X"05",X"50",X"39",X"12",X"3E",X"05",X"50",X"3A",X"12",X"3F",X"05",X"50",X"3B",X"12",X"40",
		X"05",X"50",X"3C",X"12",X"41",X"05",X"50",X"3D",X"12",X"42",X"05",X"50",X"3E",X"12",X"43",X"05",
		X"50",X"3F",X"12",X"44",X"05",X"12",X"45",X"05",X"12",X"46",X"05",X"12",X"47",X"05",X"12",X"48",
		X"05",X"12",X"49",X"05",X"12",X"4A",X"05",X"50",X"46",X"12",X"4B",X"05",X"50",X"47",X"12",X"4C",
		X"05",X"50",X"48",X"12",X"4D",X"05",X"50",X"49",X"12",X"4E",X"05",X"50",X"4A",X"12",X"4F",X"05",
		X"50",X"4B",X"12",X"50",X"05",X"50",X"04",X"12",X"51",X"05",X"50",X"4D",X"12",X"52",X"05",X"50",
		X"4E",X"12",X"53",X"05",X"50",X"4F",X"12",X"54",X"05",X"12",X"55",X"05",X"12",X"56",X"05",X"12",
		X"57",X"05",X"12",X"58",X"05",X"12",X"59",X"05",X"12",X"5A",X"05",X"50",X"56",X"12",X"5B",X"05",
		X"50",X"57",X"12",X"5C",X"05",X"50",X"58",X"12",X"5D",X"05",X"50",X"59",X"12",X"5E",X"05",X"50",
		X"5A",X"12",X"5F",X"05",X"50",X"5B",X"12",X"60",X"05",X"50",X"5C",X"12",X"61",X"05",X"50",X"5D",
		X"12",X"62",X"05",X"50",X"5E",X"12",X"63",X"05",X"50",X"5F",X"12",X"64",X"05",X"12",X"65",X"05",
		X"12",X"66",X"05",X"12",X"67",X"05",X"12",X"68",X"05",X"12",X"69",X"05",X"12",X"6A",X"05",X"50",
		X"66",X"12",X"6B",X"05",X"50",X"67",X"12",X"6C",X"05",X"50",X"68",X"12",X"6D",X"05",X"50",X"69",
		X"12",X"6E",X"05",X"50",X"6A",X"12",X"6F",X"05",X"50",X"6B",X"12",X"70",X"05",X"50",X"6C",X"12",
		X"71",X"05",X"50",X"6D",X"12",X"72",X"05",X"50",X"6E",X"12",X"73",X"05",X"50",X"6F",X"12",X"74",
		X"05",X"12",X"75",X"05",X"12",X"76",X"05",X"12",X"77",X"05",X"12",X"78",X"05",X"12",X"79",X"05",
		X"12",X"7A",X"05",X"50",X"76",X"12",X"7B",X"05",X"50",X"77",X"12",X"7C",X"05",X"50",X"78",X"12",
		X"7D",X"05",X"50",X"79",X"12",X"7E",X"05",X"50",X"7A",X"12",X"7F",X"05",X"50",X"7B",X"12",X"80",
		X"05",X"50",X"7C",X"12",X"81",X"05",X"50",X"7D",X"12",X"82",X"05",X"50",X"7E",X"12",X"83",X"05",
		X"50",X"7F",X"12",X"84",X"05",X"12",X"85",X"05",X"12",X"86",X"05",X"12",X"87",X"05",X"12",X"88",
		X"05",X"12",X"89",X"05",X"12",X"8A",X"05",X"50",X"86",X"12",X"8B",X"05",X"50",X"87",X"12",X"8C",
		X"05",X"50",X"88",X"12",X"8D",X"05",X"50",X"89",X"12",X"8E",X"05",X"50",X"8A",X"12",X"8F",X"80",
		X"59",X"00",X"58",X"00",X"77",X"03",X"FF",X"76",X"BF",X"50",X"00",X"51",X"00",X"52",X"00",X"53",
		X"00",X"58",X"00",X"59",X"00",X"77",X"BF",X"FF",X"76",X"B7",X"5B",X"03",X"5C",X"02",X"5D",X"09",
		X"58",X"10",X"16",X"01",X"28",X"58",X"00",X"16",X"00",X"28",X"77",X"08",X"5B",X"00",X"5C",X"00",
		X"5D",X"00",X"FF",X"76",X"7F",X"1E",X"01",X"04",X"1E",X"00",X"50",X"1E",X"01",X"04",X"1E",X"00",
		X"50",X"1E",X"01",X"04",X"1E",X"00",X"50",X"FF",X"76",X"7F",X"1E",X"02",X"04",X"1E",X"00",X"50",
		X"1E",X"02",X"04",X"1E",X"00",X"50",X"1E",X"02",X"04",X"1E",X"00",X"50",X"FF",X"76",X"7F",X"1E",
		X"04",X"04",X"1E",X"00",X"50",X"1E",X"04",X"04",X"1E",X"00",X"50",X"1E",X"04",X"04",X"1E",X"00",
		X"50",X"FF",X"76",X"7F",X"1E",X"08",X"04",X"1E",X"00",X"50",X"1E",X"08",X"04",X"1E",X"00",X"50",
		X"1E",X"08",X"04",X"1E",X"00",X"50",X"FF",X"76",X"BB",X"55",X"00",X"5A",X"0C",X"FE",X"F8",X"BD",
		X"14",X"00",X"E0",X"14",X"00",X"E0",X"FE",X"F8",X"87",X"76",X"BB",X"55",X"00",X"5A",X"0C",X"FE",
		X"F8",X"BD",X"FE",X"F8",X"BD",X"14",X"00",X"70",X"14",X"00",X"E0",X"FE",X"F8",X"99",X"76",X"BB",
		X"55",X"00",X"5A",X"0C",X"FE",X"F8",X"BD",X"14",X"00",X"A0",X"FE",X"F8",X"AE",X"14",X"4F",X"10",
		X"14",X"47",X"10",X"14",X"4F",X"10",X"14",X"47",X"10",X"14",X"4F",X"10",X"14",X"47",X"10",X"14",
		X"4F",X"10",X"14",X"00",X"10",X"FD",X"66",X"B8",X"41",X"00",X"43",X"00",X"45",X"00",X"40",X"6A",
		X"42",X"7E",X"6C",X"14",X"6D",X"14",X"6E",X"14",X"68",X"0C",X"69",X"0C",X"6A",X"0C",X"04",X"D4",
		X"1F",X"68",X"0C",X"69",X"0C",X"6A",X"0C",X"04",X"D4",X"1F",X"68",X"0C",X"69",X"0C",X"6A",X"0C",
		X"04",X"D4",X"1F",X"40",X"5E",X"42",X"77",X"68",X"0C",X"69",X"0C",X"6A",X"0C",X"04",X"BD",X"3E",
		X"68",X"0C",X"69",X"0C",X"6A",X"0C",X"04",X"BD",X"3E",X"68",X"0C",X"69",X"0C",X"6A",X"0C",X"04",
		X"BD",X"1F",X"40",X"6A",X"42",X"7E",X"68",X"0C",X"69",X"0C",X"6A",X"0C",X"04",X"D4",X"1F",X"68",
		X"0C",X"69",X"0C",X"6A",X"0C",X"04",X"D4",X"1F",X"68",X"0C",X"69",X"0C",X"6A",X"0C",X"04",X"D4",
		X"1F",X"40",X"5E",X"42",X"77",X"68",X"0C",X"69",X"0C",X"6A",X"0C",X"04",X"BD",X"63",X"67",X"07",
		X"FF",X"20",X"20",X"20",X"7C",X"20",X"4A",X"20",X"7C",X"20",X"20",X"20",X"7C",X"20",X"4C",X"20",
		X"7C",X"20",X"20",X"20",X"2B",X"2D",X"2D",X"2D",X"2B",X"2D",X"2D",X"2D",X"2B",X"2D",X"2D",X"2D",
		X"2B",X"20",X"20",X"20",X"7C",X"20",X"4D",X"20",X"7C",X"20",X"2C",X"20",X"7C",X"20",X"2E",X"20",
		X"7C",X"20",X"20",X"20",X"2B",X"2D",X"2D",X"2D",X"2B",X"2D",X"2D",X"2D",X"2B",X"2D",X"2D",X"2D",
		X"2B",X"20",X"20",X"20",X"50",X"3D",X"61",X"64",X"64",X"72",X"65",X"73",X"73",X"2B",X"31",X"30",
		X"30",X"30",X"48",X"20",X"3B",X"3D",X"61",X"64",X"64",X"72",X"65",X"73",X"73",X"2B",X"30",X"31",
		X"30",X"30",X"48",X"20",X"2F",X"3D",X"61",X"64",X"64",X"72",X"65",X"73",X"73",X"2D",X"30",X"31",
		X"30",X"30",X"48",X"20",X"73",X"70",X"61",X"63",X"65",X"3D",X"6E",X"65",X"78",X"74",X"20",X"62",
		X"79",X"74",X"65",X"20",X"52",X"20",X"3D",X"20",X"72",X"65",X"74",X"75",X"72",X"6E",X"20",X"20",
		X"20",X"20",X"20",X"20",X"4D",X"45",X"4D",X"4F",X"52",X"59",X"20",X"20",X"20",X"45",X"44",X"49",
		X"54",X"4F",X"52",X"20",X"00",X"06",X"00",X"10",X"FE",X"C9",X"CD",X"ED",X"F9",X"CD",X"FC",X"03",
		X"0F",X"8E",X"00",X"FF",X"BD",X"FB",X"93",X"86",X"BF",X"C6",X"07",X"BD",X"FB",X"D5",X"86",X"13",
		X"C6",X"0F",X"BD",X"FB",X"D5",X"86",X"3F",X"C6",X"17",X"BD",X"FB",X"D5",X"BD",X"FB",X"A8",X"7F",
		X"08",X"00",X"0F",X"BD",X"FB",X"43",X"96",X"BC",X"2B",X"07",X"BD",X"FD",X"DE",X"86",X"FF",X"97",
		X"BC",X"0E",X"CE",X"00",X"00",X"DF",X"D1",X"96",X"80",X"26",X"0B",X"DE",X"84",X"D6",X"8C",X"BD",
		X"FC",X"D9",X"DF",X"84",X"97",X"80",X"7C",X"00",X"D2",X"96",X"81",X"26",X"0B",X"DE",X"86",X"D6",
		X"8D",X"BD",X"FC",X"D9",X"DF",X"86",X"97",X"81",X"7C",X"00",X"D2",X"96",X"82",X"26",X"0B",X"DE",
		X"88",X"D6",X"8E",X"BD",X"FC",X"D9",X"DF",X"88",X"97",X"82",X"7C",X"00",X"D2",X"96",X"83",X"26",
		X"0B",X"DE",X"8A",X"D6",X"8F",X"BD",X"FC",X"D9",X"DF",X"8A",X"97",X"83",X"96",X"A8",X"27",X"08",
		X"7F",X"00",X"A8",X"C6",X"08",X"BD",X"FC",X"37",X"96",X"A9",X"27",X"08",X"7F",X"00",X"A9",X"C6",
		X"09",X"BD",X"FC",X"37",X"96",X"AA",X"27",X"08",X"7F",X"00",X"AA",X"C6",X"0A",X"BD",X"FC",X"37",
		X"96",X"AB",X"27",X"08",X"7F",X"00",X"AB",X"C6",X"18",X"BD",X"FC",X"50",X"96",X"AC",X"27",X"08",
		X"7F",X"00",X"AC",X"C6",X"19",X"BD",X"FC",X"50",X"96",X"AD",X"27",X"08",X"7F",X"00",X"AD",X"C6",
		X"1A",X"BD",X"FC",X"50",X"96",X"BE",X"16",X"9A",X"D8",X"0F",X"97",X"D8",X"C6",X"0F",X"BD",X"FB",
		X"DB",X"7E",X"FA",X"22",X"96",X"C1",X"B7",X"08",X"01",X"96",X"C2",X"B7",X"08",X"02",X"7C",X"00",
		X"BD",X"96",X"BF",X"4C",X"97",X"BF",X"44",X"24",X"32",X"DE",X"C3",X"09",X"27",X"1E",X"DF",X"C3",
		X"DE",X"C7",X"A6",X"00",X"44",X"44",X"44",X"44",X"97",X"C1",X"DE",X"C5",X"09",X"27",X"15",X"DF",
		X"C5",X"DE",X"C9",X"A6",X"00",X"44",X"44",X"44",X"44",X"97",X"C2",X"3B",X"86",X"01",X"9A",X"BE",
		X"97",X"BE",X"20",X"E6",X"86",X"02",X"9A",X"BE",X"97",X"BE",X"3B",X"96",X"C7",X"81",X"20",X"25",
		X"09",X"DE",X"C7",X"A6",X"00",X"97",X"C1",X"08",X"DF",X"C7",X"96",X"C9",X"81",X"20",X"25",X"09",
		X"DE",X"C9",X"A6",X"00",X"97",X"C2",X"08",X"DF",X"C9",X"96",X"BF",X"84",X"0E",X"26",X"CC",X"7C",
		X"00",X"C0",X"3B",X"96",X"C0",X"27",X"3E",X"7A",X"00",X"C0",X"96",X"80",X"27",X"06",X"4C",X"27",
		X"03",X"7A",X"00",X"80",X"96",X"81",X"27",X"06",X"4C",X"27",X"03",X"7A",X"00",X"81",X"96",X"82",
		X"27",X"06",X"4C",X"27",X"03",X"7A",X"00",X"82",X"96",X"83",X"27",X"06",X"4C",X"27",X"03",X"7A",
		X"00",X"83",X"CE",X"00",X"06",X"A6",X"AD",X"27",X"09",X"4A",X"26",X"04",X"6C",X"A7",X"A6",X"B3",
		X"A7",X"AD",X"09",X"26",X"F0",X"39",X"B7",X"08",X"00",X"C6",X"0E",X"BD",X"FC",X"1D",X"84",X"3F",
		X"97",X"BC",X"3B",X"CE",X"FF",X"FF",X"DF",X"00",X"C6",X"4F",X"08",X"86",X"00",X"A7",X"80",X"08",
		X"5A",X"26",X"FA",X"86",X"13",X"97",X"D8",X"39",X"BD",X"FB",X"C0",X"86",X"BF",X"97",X"BB",X"C6",
		X"FF",X"D7",X"82",X"D7",X"83",X"D7",X"B1",X"D7",X"B2",X"D7",X"B3",X"C6",X"17",X"7E",X"FB",X"DB",
		X"86",X"BF",X"97",X"BA",X"C6",X"FF",X"D7",X"80",X"D7",X"81",X"D7",X"AE",X"D7",X"AF",X"D7",X"B0",
		X"C6",X"07",X"7E",X"FB",X"DB",X"7C",X"00",X"BD",X"20",X"04",X"0F",X"7F",X"00",X"BD",X"37",X"36",
		X"C1",X"10",X"2A",X"19",X"86",X"0D",X"97",X"03",X"D7",X"02",X"C6",X"08",X"D7",X"03",X"5C",X"32",
		X"97",X"02",X"96",X"BD",X"27",X"FC",X"D7",X"03",X"5A",X"D7",X"03",X"33",X"39",X"86",X"15",X"97",
		X"03",X"C4",X"0F",X"D7",X"02",X"C6",X"10",X"20",X"E3",X"37",X"20",X"E4",X"37",X"86",X"15",X"97",
		X"03",X"C4",X"0F",X"D7",X"02",X"C6",X"14",X"20",X"0D",X"C1",X"10",X"2A",X"EF",X"37",X"86",X"0D",
		X"97",X"03",X"D7",X"02",X"C6",X"0C",X"4F",X"97",X"03",X"97",X"00",X"D7",X"03",X"96",X"02",X"5F",
		X"D7",X"03",X"5A",X"D7",X"00",X"33",X"39",X"0F",X"BD",X"FC",X"1D",X"C6",X"09",X"7F",X"00",X"BD",
		X"84",X"1F",X"81",X"10",X"2A",X"08",X"4A",X"81",X"07",X"2B",X"03",X"BD",X"FC",X"09",X"0E",X"39",
		X"0F",X"BD",X"FC",X"0C",X"C6",X"11",X"20",X"E5",X"17",X"84",X"0F",X"81",X"08",X"2A",X"08",X"A6",
		X"94",X"AB",X"98",X"A7",X"94",X"20",X"67",X"CB",X"38",X"DE",X"CD",X"A6",X"05",X"36",X"DE",X"D1",
		X"AB",X"94",X"A7",X"94",X"32",X"2B",X"0C",X"24",X"02",X"6C",X"98",X"BD",X"FB",X"DA",X"5C",X"A6",
		X"94",X"20",X"4B",X"25",X"F6",X"6A",X"98",X"20",X"F2",X"6F",X"8C",X"DE",X"CD",X"C1",X"A0",X"2B",
		X"02",X"08",X"08",X"08",X"08",X"08",X"C1",X"C0",X"2B",X"08",X"17",X"84",X"0F",X"81",X"08",X"2B",
		X"01",X"08",X"86",X"01",X"39",X"DF",X"CD",X"DE",X"D1",X"6A",X"90",X"27",X"DC",X"C1",X"A0",X"2A",
		X"10",X"C4",X"1F",X"A6",X"94",X"36",X"DE",X"CD",X"A6",X"03",X"BD",X"FB",X"DA",X"0E",X"32",X"08",
		X"39",X"C1",X"C0",X"2A",X"93",X"A6",X"90",X"44",X"A6",X"94",X"25",X"02",X"A6",X"98",X"C4",X"1F",
		X"BD",X"FB",X"DA",X"0E",X"DE",X"CD",X"A6",X"04",X"39",X"26",X"CA",X"DF",X"CD",X"E6",X"00",X"2A",
		X"03",X"7E",X"FD",X"90",X"C4",X"3F",X"C1",X"20",X"2A",X"11",X"A6",X"01",X"BD",X"FB",X"DA",X"0E",
		X"E6",X"00",X"08",X"08",X"58",X"2B",X"E4",X"A6",X"00",X"08",X"39",X"C4",X"1F",X"17",X"84",X"0F",
		X"26",X"31",X"A6",X"01",X"97",X"CE",X"A6",X"02",X"97",X"CD",X"BD",X"FD",X"D1",X"DC",X"CD",X"04",
		X"DD",X"CD",X"E6",X"00",X"C4",X"1F",X"5C",X"5C",X"BD",X"FD",X"D1",X"7C",X"00",X"CE",X"26",X"03",
		X"7C",X"00",X"CD",X"BD",X"FD",X"D1",X"CB",X"07",X"86",X"09",X"BD",X"FB",X"DB",X"0E",X"E6",X"00",
		X"08",X"20",X"BF",X"80",X"08",X"2B",X"29",X"DD",X"CF",X"84",X"03",X"C1",X"10",X"2B",X"02",X"8B",
		X"03",X"16",X"A6",X"01",X"CE",X"00",X"00",X"3A",X"D6",X"CF",X"C1",X"04",X"2A",X"0B",X"A6",X"B4",
		X"A7",X"AE",X"DE",X"CD",X"D6",X"D0",X"7E",X"FC",X"EA",X"A7",X"B4",X"DE",X"CD",X"7E",X"FC",X"F0",
		X"4C",X"27",X"17",X"5C",X"C1",X"10",X"2A",X"09",X"96",X"BA",X"A4",X"01",X"97",X"BA",X"7E",X"FC",
		X"EC",X"96",X"BB",X"A4",X"01",X"97",X"BB",X"7E",X"FC",X"EC",X"C1",X"10",X"2A",X"09",X"96",X"BA",
		X"AA",X"01",X"97",X"BA",X"7E",X"FC",X"EC",X"96",X"BB",X"AA",X"01",X"97",X"BB",X"7E",X"FC",X"EC",
		X"C1",X"F0",X"2A",X"17",X"A6",X"01",X"EE",X"02",X"3C",X"DE",X"D1",X"E7",X"8C",X"4C",X"A7",X"90",
		X"32",X"A7",X"94",X"32",X"A7",X"98",X"DE",X"CD",X"86",X"01",X"39",X"5C",X"27",X"12",X"DE",X"D1",
		X"5C",X"26",X"10",X"DC",X"CD",X"A7",X"9C",X"E7",X"A0",X"DE",X"CD",X"EE",X"01",X"86",X"01",X"39",
		X"86",X"FF",X"39",X"A6",X"9C",X"E6",X"A0",X"DD",X"CD",X"DE",X"CD",X"08",X"08",X"08",X"86",X"01",
		X"39",X"96",X"CE",X"BD",X"FB",X"DA",X"5C",X"96",X"CD",X"BD",X"FB",X"DB",X"5C",X"39",X"26",X"06",
		X"BD",X"FB",X"93",X"7E",X"FB",X"A8",X"81",X"10",X"2B",X"03",X"7E",X"FE",X"5B",X"81",X"07",X"2A",
		X"35",X"97",X"CB",X"96",X"D8",X"8A",X"01",X"16",X"C4",X"FE",X"D7",X"D8",X"C6",X"0F",X"BD",X"FB",
		X"DB",X"86",X"05",X"7F",X"00",X"BD",X"D6",X"BD",X"27",X"FC",X"4A",X"26",X"F6",X"D6",X"CB",X"58",
		X"58",X"CE",X"EA",X"00",X"3A",X"3C",X"EE",X"00",X"DF",X"C7",X"38",X"EE",X"02",X"DF",X"C3",X"96",
		X"BE",X"84",X"02",X"97",X"BE",X"39",X"97",X"CC",X"96",X"D8",X"8A",X"02",X"16",X"C4",X"FD",X"D7",
		X"D8",X"C6",X"0F",X"BD",X"FB",X"DB",X"86",X"05",X"7F",X"00",X"BD",X"D6",X"BD",X"27",X"FC",X"4A",
		X"26",X"F6",X"D6",X"CC",X"58",X"58",X"CE",X"EA",X"00",X"3A",X"3C",X"EE",X"00",X"DF",X"C9",X"38",
		X"EE",X"02",X"DF",X"C5",X"96",X"BE",X"84",X"01",X"97",X"BE",X"39",X"16",X"58",X"CE",X"EA",X"30",
		X"3A",X"EE",X"00",X"81",X"20",X"2B",X"22",X"7E",X"FE",X"6E",X"81",X"15",X"2A",X"34",X"3C",X"36",
		X"BD",X"FB",X"93",X"BD",X"FB",X"A8",X"32",X"38",X"97",X"A4",X"DF",X"84",X"7F",X"00",X"80",X"7F",
		X"00",X"8C",X"C6",X"B8",X"DA",X"BA",X"D7",X"BA",X"39",X"81",X"13",X"2A",X"DD",X"81",X"1F",X"27",
		X"DD",X"DF",X"88",X"97",X"A6",X"7F",X"00",X"82",X"7F",X"00",X"8E",X"86",X"78",X"9A",X"BB",X"97",
		X"BB",X"39",X"81",X"18",X"2A",X"E7",X"DF",X"8A",X"97",X"A7",X"7F",X"00",X"83",X"7F",X"00",X"8F",
		X"86",X"78",X"9A",X"BB",X"97",X"BB",X"39",X"81",X"15",X"2A",X"E7",X"DF",X"86",X"7F",X"00",X"8D",
		X"7F",X"00",X"81",X"86",X"B8",X"9A",X"BA",X"97",X"BA",X"39",X"06",X"91",X"68",X"F6",X"06",X"91",
		X"68",X"F6",X"06",X"91",X"68",X"F6",X"06",X"91",X"68",X"F6",X"06",X"91",X"68",X"F6",X"06",X"91",
		X"68",X"F6",X"06",X"91",X"68",X"F6",X"06",X"91",X"68",X"F6",X"06",X"91",X"68",X"F6",X"06",X"91",
		X"68",X"F6",X"06",X"91",X"68",X"F6",X"06",X"91",X"68",X"F6",X"06",X"91",X"68",X"00",X"00",X"00",
		X"09",X"0A",X"0C",X"0D",X"0F",X"10",X"12",X"13",X"15",X"16",X"18",X"19",X"1B",X"1C",X"1E",X"1F",
		X"23",X"24",X"26",X"27",X"29",X"2A",X"2C",X"2D",X"2F",X"30",X"32",X"33",X"35",X"36",X"38",X"39",
		X"22",X"5A",X"38",X"30",X"22",X"3B",X"3B",X"20",X"20",X"64",X"65",X"74",X"61",X"20",X"69",X"73",
		X"20",X"20",X"2D",X"2D",X"2D",X"2D",X"48",X"20",X"74",X"6F",X"20",X"2D",X"2D",X"2D",X"2D",X"48",
		X"45",X"4E",X"44",X"48",X"45",X"58",X"3E",X"3E",X"20",X"50",X"61",X"72",X"61",X"6D",X"74",X"65",
		X"72",X"20",X"65",X"72",X"72",X"6F",X"72",X"20",X"3C",X"3C",X"0D",X"00",X"44",X"55",X"4D",X"50",
		X"20",X"4C",X"49",X"53",X"54",X"20",X"50",X"41",X"47",X"45",X"20",X"3D",X"20",X"F6",X"06",X"0D",
		X"0D",X"00",X"06",X"91",X"68",X"F6",X"06",X"91",X"68",X"F6",X"06",X"91",X"68",X"F6",X"06",X"91",
		X"68",X"F6",X"06",X"91",X"68",X"F6",X"06",X"91",X"68",X"F6",X"06",X"91",X"68",X"F6",X"06",X"91",
		X"68",X"F6",X"06",X"91",X"68",X"F6",X"06",X"91",X"68",X"F6",X"06",X"91",X"68",X"F6",X"06",X"91",
		X"68",X"F6",X"06",X"91",X"68",X"F6",X"06",X"91",X"68",X"F6",X"06",X"91",X"68",X"F6",X"06",X"91",
		X"68",X"F6",X"06",X"91",X"68",X"F6",X"06",X"91",X"68",X"F6",X"06",X"91",X"68",X"F6",X"06",X"91",
		X"68",X"F6",X"06",X"91",X"68",X"F6",X"06",X"91",X"68",X"F6",X"06",X"91",X"68",X"F6",X"06",X"91",
		X"68",X"F6",X"06",X"91",X"68",X"F6",X"06",X"91",X"68",X"F6",X"06",X"91",X"68",X"F6",X"06",X"91",
		X"68",X"F6",X"00",X"00",X"00",X"00",X"06",X"91",X"68",X"F6",X"06",X"91",X"68",X"F6",X"06",X"91",
		X"FA",X"00",X"FA",X"00",X"FA",X"00",X"FA",X"00",X"FB",X"86",X"FA",X"00",X"FA",X"D4",X"FA",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
