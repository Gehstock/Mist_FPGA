library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_E1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_E1 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"C6",X"C6",X"20",X"53",X"3D",X"A5",X"C6",X"D0",X"03",X"4C",X"AE",X"3B",X"20",X"8C",X"3B",X"90",
		X"0A",X"20",X"38",X"3D",X"24",X"BB",X"10",X"03",X"20",X"53",X"3D",X"20",X"72",X"3D",X"4C",X"B7",
		X"37",X"20",X"D3",X"3A",X"A9",X"01",X"85",X"00",X"20",X"2E",X"3D",X"E6",X"B8",X"20",X"08",X"36",
		X"A2",X"06",X"20",X"C0",X"39",X"95",X"68",X"B5",X"41",X"30",X"1A",X"B5",X"A1",X"F0",X"05",X"D6",
		X"A1",X"4C",X"73",X"38",X"B5",X"41",X"30",X"0D",X"A9",X"00",X"95",X"A1",X"A9",X"F7",X"35",X"A0",
		X"95",X"A0",X"4C",X"73",X"38",X"95",X"20",X"A0",X"00",X"94",X"C7",X"B5",X"A0",X"29",X"08",X"D0",
		X"0E",X"A9",X"01",X"95",X"80",X"A9",X"08",X"15",X"A0",X"95",X"A0",X"A9",X"0F",X"85",X"CF",X"A9",
		X"10",X"95",X"A1",X"A4",X"CF",X"F0",X"0B",X"8A",X"D0",X"0A",X"A5",X"B8",X"29",X"03",X"D0",X"04",
		X"C6",X"CF",X"84",X"42",X"B5",X"C7",X"F0",X"1A",X"95",X"69",X"D6",X"C7",X"A0",X"02",X"B5",X"A0",
		X"30",X"04",X"A0",X"02",X"D0",X"06",X"29",X"10",X"D0",X"02",X"A0",X"FE",X"98",X"18",X"75",X"99",
		X"95",X"99",X"B5",X"A0",X"10",X"28",X"A5",X"B8",X"29",X"03",X"D0",X"22",X"20",X"03",X"3B",X"C9",
		X"F9",X"10",X"02",X"95",X"69",X"C9",X"00",X"18",X"30",X"0C",X"75",X"80",X"D0",X"0E",X"B5",X"80",
		X"F0",X"0A",X"A9",X"FF",X"D0",X"06",X"75",X"80",X"D0",X"02",X"A9",X"01",X"95",X"80",X"B5",X"80",
		X"4A",X"4A",X"4A",X"85",X"BC",X"B5",X"B1",X"B4",X"A0",X"30",X"0C",X"B5",X"99",X"4A",X"4A",X"4A",
		X"4A",X"4A",X"09",X"88",X"4C",X"07",X"39",X"A8",X"0A",X"85",X"BE",X"B9",X"C4",X"3D",X"A8",X"A9",
		X"00",X"18",X"65",X"BC",X"88",X"D0",X"FA",X"4A",X"4A",X"4A",X"38",X"E5",X"BE",X"10",X"02",X"A9",
		X"00",X"C9",X"10",X"30",X"02",X"A9",X"0F",X"95",X"91",X"A9",X"04",X"B4",X"80",X"10",X"02",X"A9",
		X"03",X"85",X"BC",X"B5",X"99",X"29",X"F8",X"85",X"BE",X"B5",X"81",X"29",X"F8",X"38",X"E5",X"BE",
		X"F0",X"1F",X"30",X"10",X"C9",X"10",X"30",X"02",X"95",X"69",X"A9",X"00",X"38",X"E5",X"BC",X"85",
		X"BC",X"4C",X"3A",X"39",X"C9",X"F8",X"10",X"02",X"95",X"69",X"A5",X"BC",X"18",X"75",X"81",X"95",
		X"81",X"20",X"42",X"3A",X"20",X"35",X"3C",X"E0",X"00",X"D0",X"0C",X"C6",X"D0",X"D0",X"08",X"C6",
		X"D3",X"F0",X"15",X"A5",X"D1",X"85",X"D0",X"CA",X"CA",X"30",X"03",X"4C",X"32",X"38",X"2C",X"00",
		X"10",X"30",X"FB",X"85",X"44",X"4C",X"28",X"38",X"A9",X"00",X"85",X"00",X"85",X"BB",X"85",X"BE",
		X"A5",X"DD",X"4A",X"F0",X"04",X"A9",X"40",X"85",X"BB",X"A9",X"02",X"85",X"BF",X"A2",X"06",X"B5",
		X"A0",X"29",X"03",X"95",X"A0",X"CA",X"CA",X"10",X"F6",X"A2",X"06",X"A9",X"F0",X"95",X"68",X"35",
		X"91",X"95",X"91",X"9D",X"60",X"00",X"20",X"1B",X"3D",X"20",X"9F",X"3C",X"CA",X"CA",X"10",X"EB",
		X"A9",X"00",X"85",X"42",X"85",X"44",X"2C",X"00",X"10",X"30",X"FB",X"2C",X"00",X"10",X"10",X"FB",
		X"E6",X"B8",X"A5",X"BB",X"10",X"01",X"60",X"C6",X"BE",X"D0",X"CE",X"C6",X"BF",X"D0",X"CA",X"60",
		X"B5",X"A0",X"30",X"7D",X"B5",X"C7",X"F0",X"04",X"29",X"03",X"D0",X"66",X"A9",X"00",X"85",X"BC",
		X"A9",X"08",X"85",X"BD",X"B5",X"A8",X"18",X"69",X"F8",X"4A",X"4A",X"4A",X"18",X"65",X"BC",X"85",
		X"BC",X"A9",X"00",X"85",X"BE",X"65",X"BD",X"85",X"BD",X"B5",X"A9",X"18",X"69",X"FB",X"29",X"F8",
		X"0A",X"26",X"BE",X"0A",X"26",X"BE",X"18",X"65",X"BC",X"85",X"BC",X"A5",X"BE",X"65",X"BD",X"85",
		X"BD",X"B5",X"99",X"29",X"F8",X"85",X"C0",X"A0",X"00",X"B1",X"BC",X"4A",X"B0",X"02",X"29",X"6F",
		X"0A",X"29",X"E0",X"38",X"E5",X"C0",X"29",X"F8",X"F0",X"18",X"4A",X"4A",X"4A",X"4A",X"18",X"2C",
		X"35",X"3B",X"F0",X"07",X"09",X"F0",X"69",X"FE",X"4C",X"2D",X"3A",X"69",X"02",X"18",X"75",X"99",
		X"95",X"99",X"B5",X"80",X"18",X"69",X"01",X"DD",X"CC",X"3D",X"90",X"03",X"BD",X"CC",X"3D",X"95",
		X"80",X"60",X"86",X"BC",X"B5",X"80",X"F0",X"59",X"4A",X"4A",X"4A",X"85",X"BE",X"B5",X"81",X"4A",
		X"4A",X"4A",X"AA",X"86",X"C0",X"BD",X"E0",X"3D",X"F0",X"20",X"AA",X"20",X"A4",X"3A",X"A6",X"BC",
		X"A5",X"C2",X"18",X"75",X"88",X"95",X"88",X"A5",X"C3",X"75",X"A8",X"A0",X"10",X"C9",X"10",X"90",
		X"06",X"C9",X"F8",X"90",X"03",X"A0",X"F8",X"98",X"95",X"A8",X"A6",X"C0",X"BD",X"D8",X"3D",X"F0",
		X"20",X"AA",X"20",X"A4",X"3A",X"A6",X"BC",X"A5",X"C2",X"18",X"75",X"89",X"95",X"89",X"A5",X"C3",
		X"75",X"A9",X"A0",X"12",X"C9",X"12",X"90",X"06",X"C9",X"DF",X"90",X"03",X"A0",X"DE",X"98",X"95",
		X"A9",X"A6",X"BC",X"60",X"86",X"BF",X"8A",X"10",X"04",X"49",X"FF",X"AA",X"E8",X"A9",X"00",X"85",
		X"C2",X"85",X"C3",X"A5",X"C2",X"18",X"65",X"BE",X"85",X"C2",X"90",X"02",X"E6",X"C3",X"CA",X"D0",
		X"F2",X"A5",X"BF",X"10",X"0D",X"A9",X"00",X"38",X"E5",X"C2",X"85",X"C2",X"A9",X"00",X"E5",X"C3",
		X"85",X"C3",X"60",X"A0",X"00",X"A5",X"63",X"4A",X"6A",X"90",X"0C",X"C8",X"2A",X"90",X"08",X"C8",
		X"A5",X"62",X"4A",X"4A",X"90",X"01",X"C8",X"B9",X"C8",X"3D",X"85",X"D0",X"85",X"D1",X"A9",X"00",
		X"85",X"D2",X"85",X"CF",X"85",X"42",X"A9",X"64",X"85",X"D3",X"85",X"20",X"85",X"22",X"85",X"24",
		X"85",X"26",X"60",X"B5",X"80",X"4A",X"4A",X"4A",X"4A",X"0A",X"A8",X"B5",X"B1",X"4A",X"4A",X"90",
		X"01",X"C8",X"B5",X"40",X"30",X"05",X"B9",X"00",X"3E",X"D0",X"03",X"B9",X"20",X"3E",X"18",X"B4",
		X"B1",X"84",X"BC",X"46",X"BC",X"B0",X"04",X"4A",X"4A",X"4A",X"4A",X"29",X"0F",X"2C",X"35",X"3B",
		X"F0",X"02",X"09",X"F0",X"60",X"08",X"84",X"C2",X"A8",X"B9",X"58",X"3E",X"85",X"BE",X"B9",X"59",
		X"3E",X"85",X"BF",X"A5",X"60",X"29",X"03",X"48",X"86",X"C0",X"0A",X"0A",X"0A",X"85",X"C4",X"68",
		X"0A",X"18",X"65",X"C4",X"18",X"65",X"C0",X"AA",X"BD",X"82",X"3E",X"85",X"C0",X"BD",X"83",X"3E",
		X"85",X"C1",X"A0",X"00",X"B1",X"C0",X"F0",X"23",X"A6",X"C2",X"10",X"02",X"09",X"80",X"29",X"BF",
		X"A2",X"00",X"81",X"BE",X"A5",X"C2",X"18",X"65",X"BE",X"85",X"BE",X"A9",X"00",X"24",X"C2",X"10",
		X"02",X"A9",X"FF",X"65",X"BF",X"85",X"BF",X"C8",X"4C",X"64",X"3B",X"60",X"18",X"2C",X"00",X"18",
		X"10",X"05",X"A5",X"D2",X"D0",X"0A",X"60",X"A9",X"04",X"A4",X"D2",X"85",X"D2",X"F0",X"04",X"60",
		X"C6",X"D2",X"60",X"A4",X"B9",X"C8",X"C0",X"0A",X"90",X"02",X"A0",X"00",X"84",X"B9",X"A0",X"21",
		X"A9",X"A0",X"99",X"00",X"08",X"A9",X"20",X"99",X"5E",X"0B",X"88",X"10",X"F3",X"A9",X"0A",X"20",
		X"C4",X"3B",X"A5",X"B9",X"0A",X"85",X"BE",X"0A",X"18",X"65",X"BE",X"A8",X"86",X"C4",X"A2",X"00",
		X"B9",X"01",X"28",X"95",X"BC",X"C8",X"E8",X"E0",X"06",X"D0",X"F5",X"A2",X"00",X"A0",X"00",X"C0",
		X"00",X"D0",X"0C",X"A9",X"06",X"20",X"19",X"3C",X"A9",X"02",X"20",X"19",X"3C",X"A0",X"0F",X"A1",
		X"BC",X"48",X"4A",X"4A",X"4A",X"4A",X"20",X"19",X"3C",X"68",X"20",X"19",X"3C",X"E6",X"BE",X"D0",
		X"04",X"E6",X"BF",X"F0",X"0C",X"88",X"85",X"44",X"E6",X"BC",X"D0",X"D3",X"E6",X"BD",X"4C",X"DF",
		X"3B",X"A6",X"C4",X"A9",X"00",X"85",X"DE",X"38",X"60",X"29",X"0F",X"4A",X"AA",X"BD",X"40",X"3E",
		X"2C",X"34",X"3C",X"D0",X"02",X"09",X"00",X"69",X"00",X"A2",X"00",X"81",X"C0",X"E6",X"C0",X"D0",
		X"02",X"E6",X"C1",X"60",X"02",X"B5",X"A0",X"10",X"66",X"A5",X"B9",X"0A",X"0A",X"0A",X"0A",X"85",
		X"BC",X"B5",X"D5",X"0A",X"29",X"1C",X"C9",X"10",X"D0",X"08",X"A0",X"A0",X"A9",X"05",X"85",X"BC",
		X"D0",X"08",X"18",X"65",X"BC",X"A8",X"A9",X"04",X"85",X"BC",X"B5",X"A9",X"29",X"F0",X"85",X"C4",
		X"B5",X"A8",X"4A",X"4A",X"4A",X"4A",X"29",X"0F",X"05",X"C4",X"85",X"C4",X"B9",X"43",X"28",X"C5",
		X"C4",X"F0",X"07",X"C8",X"C6",X"BC",X"D0",X"F4",X"F0",X"25",X"F8",X"18",X"A9",X"02",X"75",X"D5",
		X"95",X"D5",X"A9",X"00",X"75",X"D6",X"95",X"D6",X"D8",X"A4",X"D4",X"D9",X"D6",X"00",X"90",X"0F",
		X"F0",X"02",X"B0",X"09",X"B5",X"D5",X"D9",X"D5",X"00",X"90",X"04",X"F0",X"02",X"86",X"D4",X"BC",
		X"48",X"3E",X"84",X"BC",X"BC",X"49",X"3E",X"84",X"BD",X"A0",X"00",X"B5",X"91",X"10",X"22",X"E0",
		X"03",X"90",X"0F",X"A9",X"1C",X"20",X"01",X"3D",X"A9",X"1D",X"20",X"01",X"3D",X"A9",X"1E",X"4C",
		X"01",X"3D",X"A9",X"9C",X"20",X"01",X"3D",X"A9",X"9D",X"20",X"01",X"3D",X"A9",X"9E",X"4C",X"01",
		X"3D",X"E4",X"D4",X"D0",X"15",X"A9",X"18",X"24",X"B8",X"D0",X"0F",X"A9",X"20",X"20",X"01",X"3D",
		X"A9",X"20",X"20",X"01",X"3D",X"A9",X"20",X"4C",X"01",X"3D",X"B5",X"D6",X"20",X"FA",X"3C",X"B5",
		X"D5",X"4A",X"4A",X"4A",X"4A",X"20",X"FA",X"3C",X"B5",X"D5",X"29",X"0F",X"09",X"30",X"1D",X"50",
		X"3E",X"91",X"BC",X"A5",X"BC",X"18",X"7D",X"51",X"3E",X"85",X"BC",X"BD",X"51",X"3E",X"10",X"04",
		X"A9",X"FF",X"D0",X"02",X"A9",X"00",X"65",X"BD",X"85",X"BD",X"60",X"B5",X"A8",X"95",X"90",X"B5",
		X"A9",X"95",X"98",X"B5",X"A0",X"10",X"06",X"B5",X"91",X"29",X"0F",X"95",X"91",X"60",X"A2",X"06",
		X"20",X"1B",X"3D",X"CA",X"CA",X"10",X"F9",X"60",X"A2",X"02",X"A5",X"61",X"4A",X"B0",X"02",X"A2",
		X"04",X"86",X"C3",X"A0",X"01",X"A9",X"04",X"20",X"36",X"3B",X"A6",X"C3",X"A0",X"FF",X"A9",X"08",
		X"4C",X"36",X"3B",X"A0",X"01",X"A2",X"00",X"A9",X"02",X"20",X"36",X"3B",X"A0",X"FF",X"A2",X"00",
		X"A9",X"06",X"20",X"36",X"3B",X"A5",X"C6",X"09",X"30",X"8D",X"05",X"0A",X"09",X"80",X"8D",X"59",
		X"09",X"60",X"A5",X"DE",X"C5",X"DD",X"D0",X"01",X"60",X"A5",X"60",X"29",X"03",X"85",X"BC",X"A8",
		X"B9",X"6A",X"3E",X"A0",X"01",X"A2",X"08",X"20",X"36",X"3B",X"A4",X"BC",X"B9",X"6E",X"3E",X"A0",
		X"FF",X"A2",X"08",X"20",X"36",X"3B",X"06",X"BC",X"A4",X"BC",X"B9",X"72",X"3E",X"85",X"BC",X"B9",
		X"73",X"3E",X"85",X"BD",X"B9",X"7A",X"3E",X"85",X"BE",X"B9",X"7B",X"3E",X"85",X"BF",X"A5",X"DD",
		X"85",X"DE",X"4A",X"C9",X"04",X"90",X"02",X"A9",X"04",X"09",X"30",X"A0",X"00",X"91",X"BC",X"09",
		X"80",X"91",X"BE",X"60",X"0C",X"08",X"06",X"05",X"26",X"38",X"4B",X"5E",X"A0",X"D0",X"90",X"C0",
		X"80",X"B0",X"70",X"A0",X"00",X"00",X"00",X"00",X"EA",X"EA",X"EC",X"EE",X"F0",X"F4",X"F8",X"FC",
		X"00",X"04",X"08",X"0C",X"10",X"12",X"14",X"16",X"16",X"16",X"14",X"12",X"10",X"0C",X"08",X"04",
		X"00",X"FC",X"F8",X"F4",X"F0",X"EE",X"EC",X"EA",X"EA",X"EA",X"EC",X"EE",X"F0",X"F4",X"F8",X"FC",
		X"71",X"11",X"62",X"11",X"43",X"11",X"25",X"21",X"04",X"21",X"F3",X"21",X"E2",X"31",X"D1",X"41",
		X"D0",X"41",X"CF",X"32",X"BE",X"12",X"BE",X"13",X"AE",X"03",X"9D",X"F2",X"9D",X"E2",X"9C",X"D1",
		X"00",X"00",X"EF",X"FF",X"CF",X"FF",X"AE",X"FF",X"9E",X"FF",X"9D",X"EF",X"9D",X"EF",X"9C",X"EF",
		X"9C",X"EF",X"9B",X"DE",X"9B",X"DE",X"9A",X"CE",X"9A",X"BE",X"99",X"BD",X"99",X"AC",X"99",X"AB",
		X"20",X"60",X"A0",X"E0",X"22",X"62",X"A2",X"E2",X"08",X"08",X"19",X"08",X"77",X"0B",X"66",X"0B",
		X"C0",X"FF",X"80",X"FF",X"40",X"01",X"00",X"01",X"A9",X"09",X"06",X"0A",X"87",X"0A",X"58",X"09",
		X"D7",X"08",X"04",X"0B",X"06",X"0B",X"5B",X"08",X"59",X"08",X"0A",X"0C",X"0C",X"0C",X"0E",X"10",
		X"10",X"10",X"03",X"0B",X"12",X"0B",X"06",X"0B",X"11",X"0B",X"5C",X"08",X"4D",X"08",X"59",X"08",
		X"4E",X"08",X"7E",X"3F",X"88",X"3F",X"9D",X"3F",X"E4",X"3E",X"B2",X"3F",X"44",X"3F",X"1D",X"3F",
		X"30",X"3F",X"E4",X"3E",X"CC",X"3F",X"55",X"3F",X"F2",X"3E",X"07",X"3F",X"E4",X"3E",X"E2",X"3F",
		X"AA",X"3E",X"BF",X"3E",X"D1",X"3E",X"E4",X"3E",X"69",X"3F",X"20",X"53",X"45",X"43",X"4F",X"4E",
		X"44",X"53",X"20",X"55",X"4E",X"54",X"49",X"4C",X"20",X"53",X"54",X"41",X"52",X"54",X"00",X"31",
		X"20",X"43",X"4F",X"49",X"4E",X"20",X"50",X"45",X"52",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",
		X"00",X"32",X"20",X"43",X"4F",X"49",X"4E",X"53",X"20",X"50",X"45",X"52",X"20",X"50",X"4C",X"41",
		X"59",X"45",X"52",X"00",X"52",X"41",X"4D",X"20",X"4F",X"4B",X"20",X"52",X"4F",X"4D",X"20",X"4F",
		X"4B",X"00",X"31",X"20",X"4D",X"4F",X"4E",X"45",X"44",X"41",X"20",X"50",X"4F",X"52",X"20",X"4A",
		X"55",X"47",X"41",X"44",X"4F",X"52",X"00",X"32",X"20",X"4D",X"4F",X"4E",X"45",X"44",X"41",X"53",
		X"20",X"50",X"4F",X"52",X"20",X"4A",X"55",X"47",X"41",X"44",X"4F",X"52",X"00",X"31",X"20",X"50",
		X"49",X"45",X"43",X"45",X"20",X"50",X"41",X"52",X"20",X"4A",X"4F",X"55",X"45",X"55",X"52",X"00",
		X"32",X"20",X"50",X"49",X"45",X"43",X"45",X"53",X"20",X"50",X"41",X"52",X"20",X"4A",X"4F",X"55",
		X"45",X"55",X"52",X"00",X"20",X"53",X"45",X"43",X"4F",X"4E",X"44",X"45",X"53",X"20",X"44",X"45",
		X"50",X"41",X"52",X"54",X"00",X"20",X"53",X"45",X"47",X"55",X"4E",X"44",X"4F",X"53",X"20",X"44",
		X"45",X"20",X"45",X"53",X"50",X"45",X"52",X"41",X"00",X"43",X"52",X"45",X"44",X"49",X"54",X"20",
		X"46",X"4F",X"52",X"20",X"20",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"53",X"00",X"20",X"53",
		X"45",X"4B",X"55",X"4E",X"44",X"45",X"4E",X"00",X"31",X"20",X"4D",X"55",X"45",X"4E",X"5A",X"45",
		X"20",X"50",X"52",X"4F",X"20",X"53",X"50",X"49",X"45",X"4C",X"45",X"52",X"00",X"32",X"20",X"4D",
		X"55",X"45",X"4E",X"5A",X"45",X"20",X"50",X"52",X"4F",X"20",X"53",X"50",X"49",X"45",X"4C",X"45",
		X"52",X"00",X"20",X"53",X"50",X"49",X"45",X"4C",X"45",X"52",X"20",X"48",X"41",X"42",X"45",X"4E",
		X"20",X"47",X"55",X"54",X"53",X"43",X"48",X"52",X"49",X"46",X"54",X"00",X"43",X"52",X"45",X"44",
		X"49",X"54",X"20",X"50",X"4F",X"55",X"52",X"20",X"20",X"20",X"4A",X"4F",X"55",X"45",X"55",X"52",
		X"53",X"00",X"20",X"20",X"4A",X"55",X"47",X"41",X"44",X"4F",X"52",X"45",X"53",X"20",X"41",X"56",
		X"45",X"4E",X"54",X"41",X"4A",X"41",X"4E",X"00",X"82",X"00",X"0A",X"35",X"27",X"35",X"27",X"35");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
