library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity silverland_big_sprite_tile_bit0 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of silverland_big_sprite_tile_bit0 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"06",X"1A",X"60",X"80",
		X"00",X"00",X"00",X"00",X"7F",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"03",X"03",
		X"06",X"78",X"40",X"00",X"81",X"01",X"00",X"80",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"FF",X"7F",X"00",X"00",X"00",X"00",X"03",X"03",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"C0",X"00",X"01",X"81",X"00",X"40",X"7F",X"06",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"60",X"1A",X"06",X"02",X"00",X"00",X"00",
		X"00",X"00",X"00",X"40",X"60",X"58",X"06",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"60",X"1E",X"02",X"00",X"81",X"80",X"00",X"03",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"C0",X"C0",X"00",X"00",X"00",X"00",X"FE",X"FF",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"80",X"81",X"00",X"02",X"1E",X"60",
		X"C0",X"C0",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FE",X"00",X"00",X"00",X"00",
		X"01",X"06",X"58",X"60",X"40",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"20",X"30",X"18",X"00",X"00",X"00",X"00",X"C0",X"E0",X"70",X"38",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1C",X"0E",X"07",X"03",X"01",X"00",X"00",X"00",X"1C",X"0E",X"07",X"83",X"C1",X"E1",X"73",X"3F",
		X"00",X"00",X"1F",X"90",X"C0",X"80",X"00",X"00",X"00",X"01",X"FF",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1D",X"08",X"00",X"30",X"20",X"20",X"20",X"20",
		X"00",X"00",X"00",X"00",X"01",X"00",X"10",X"38",X"00",X"00",X"00",X"80",X"C0",X"E0",X"70",X"38",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"70",
		X"1C",X"0E",X"07",X"03",X"01",X"00",X"00",X"00",X"1C",X"0E",X"04",X"80",X"00",X"00",X"00",X"00",
		X"04",X"06",X"06",X"07",X"03",X"03",X"01",X"01",X"20",X"38",X"18",X"1C",X"0C",X"8E",X"86",X"C7",
		X"38",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C3",X"E3",X"63",X"7F",X"3F",X"38",X"00",X"C0",
		X"10",X"98",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"81",X"83",X"83",X"81",X"81",
		X"00",X"00",X"08",X"18",X"0C",X"8E",X"86",X"C7",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"C3",X"E3",X"61",X"71",X"21",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",
		X"20",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0F",X"0F",
		X"30",X"30",X"30",X"30",X"30",X"30",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"09",X"61",X"40",X"40",X"40",X"80",X"80",X"0C",
		X"90",X"06",X"02",X"02",X"02",X"01",X"01",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"01",X"02",X"02",X"04",X"04",X"08",X"1C",X"00",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",
		X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"80",X"40",X"40",X"20",X"20",X"10",X"38",X"00",
		X"80",X"C0",X"C0",X"E0",X"60",X"70",X"30",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"07",X"06",X"0E",X"0C",X"1C",
		X"18",X"1C",X"0C",X"0E",X"06",X"07",X"03",X"03",X"E0",X"40",X"80",X"80",X"80",X"00",X"01",X"81",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C1",X"18",X"38",X"30",X"70",X"60",X"E0",X"C0",X"C0",
		X"03",X"03",X"02",X"06",X"06",X"00",X"00",X"00",X"80",X"C0",X"C0",X"E0",X"00",X"00",X"30",X"38",
		X"81",X"03",X"03",X"03",X"00",X"00",X"0C",X"1C",X"80",X"80",X"00",X"60",X"60",X"20",X"20",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"1C",X"0C",X"0E",X"04",X"00",X"00",X"00",
		X"18",X"38",X"30",X"70",X"20",X"00",X"00",X"00",X"10",X"10",X"10",X"08",X"08",X"1C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0E",X"0C",X"1C",X"18",
		X"00",X"00",X"00",X"20",X"70",X"30",X"38",X"18",X"00",X"00",X"1C",X"08",X"08",X"10",X"10",X"10",
		X"00",X"00",X"00",X"06",X"06",X"02",X"03",X"03",X"38",X"30",X"00",X"00",X"E0",X"C0",X"C0",X"80",
		X"1C",X"0C",X"00",X"00",X"03",X"03",X"03",X"81",X"20",X"20",X"20",X"60",X"60",X"00",X"80",X"80",
		X"03",X"03",X"07",X"06",X"0E",X"0C",X"1C",X"18",X"81",X"01",X"00",X"80",X"80",X"80",X"40",X"E0",
		X"C1",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"E0",X"60",X"70",X"30",X"38",X"18",
		X"38",X"30",X"70",X"60",X"E0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"0C",X"0E",X"06",X"07",X"03",X"03",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"60",X"10",X"10",X"08",X"08",X"04",X"04",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"20",X"10",X"28",X"74",
		X"02",X"01",X"01",X"00",X"01",X"01",X"00",X"01",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"E0",
		X"00",X"00",X"00",X"01",X"01",X"02",X"02",X"06",X"72",X"A1",X"80",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"C0",X"C0",X"40",X"60",X"00",X"A0",X"10",X"10",X"08",X"08",X"04",X"04",X"02",
		X"06",X"00",X"00",X"00",X"00",X"01",X"03",X"00",X"00",X"00",X"40",X"70",X"F8",X"F8",X"7C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"01",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"08",X"04",X"04",X"02",X"02",X"02",X"02",X"20",X"10",X"08",X"08",X"04",X"04",X"04",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"02",X"02",X"00",X"02",X"02",X"00",X"02",X"04",X"04",X"04",X"00",X"04",X"04",X"00",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"04",X"02",X"02",X"02",
		X"00",X"00",X"00",X"10",X"08",X"04",X"04",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"01",X"01",X"01",X"00",X"01",X"01",X"00",
		X"04",X"02",X"02",X"02",X"00",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"00",X"08",X"08",X"00",X"08",X"00",X"00",X"10",X"00",X"10",X"10",X"00",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"04",X"02",X"02",X"02",
		X"00",X"00",X"00",X"10",X"08",X"04",X"04",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"01",X"01",X"01",X"00",X"01",X"01",X"00",
		X"04",X"02",X"02",X"02",X"00",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"08",X"04",X"04",X"02",X"02",X"02",X"02",X"20",X"10",X"08",X"08",X"04",X"04",X"04",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"02",X"02",X"00",X"02",X"02",X"00",X"02",X"04",X"04",X"04",X"00",X"04",X"04",X"00",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"08",X"04",X"04",X"02",X"01",X"01",X"00",X"00",X"10",X"08",X"08",X"04",X"02",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"00",X"01",X"01",X"00",X"01",X"00",X"02",X"02",X"00",X"02",X"02",X"00",X"02",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"84",X"82",X"81",X"80",X"40",X"40",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"20",X"10",X"08",X"04",X"02",X"02",X"00",X"20",X"10",X"08",X"08",X"08",X"08",X"04",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"08",X"08",X"00",X"08",X"08",X"08",X"00",X"10",X"10",X"10",X"00",X"10",X"10",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"08",X"00",X"08",X"00",X"08",X"00",X"00",X"10",X"10",X"00",X"10",X"00",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"84",X"82",X"81",X"80",X"40",X"40",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"20",X"10",X"08",X"04",X"02",X"02",X"00",X"20",X"10",X"08",X"08",X"08",X"08",X"04",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"08",X"04",X"04",X"02",X"01",X"01",X"00",X"00",X"10",X"08",X"08",X"04",X"02",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"00",X"01",X"01",X"00",X"01",X"00",X"02",X"02",X"00",X"02",X"02",X"00",X"02",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
