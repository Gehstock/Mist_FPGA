library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity prom_palette_ic40 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(6 downto 0);
	data : out std_logic_vector(2 downto 0)
);
end entity;

architecture prom of prom_palette_ic40 is
	type rom is array(0 to  127) of std_logic_vector(2 downto 0);
	signal rom_data: rom := (
		"000","000","000","000","000","000","000","000","010","010","100","010","101","010","010","010",
		"000","001","010","000","010","001","001","001","000","001","001","001","110","100","100","100",
		"000","000","000","000","000","000","000","000","100","001","001","011","011","011","001","000",
		"010","101","101","001","001","001","111","000","110","111","111","101","101","101","011","111",
		"000","000","000","000","000","000","000","000","010","010","100","010","001","001","001","001",
		"000","001","010","000","010","010","010","010","000","001","001","001","100","100","100","100",
		"000","000","000","000","000","000","000","000","100","001","001","100","100","100","011","100",
		"010","101","101","101","101","101","111","000","101","111","111","011","011","011","101","111");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
