library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity travusa_chr_bit2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of travusa_chr_bit2 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"B0",X"B8",X"A8",X"E8",X"68",X"00",X"00",X"08",X"7C",X"FC",X"88",X"C8",X"40",X"00",
		X"00",X"00",X"F8",X"F8",X"08",X"F8",X"F0",X"00",X"60",X"F0",X"90",X"F0",X"7C",X"FC",X"00",X"00",
		X"00",X"00",X"F8",X"F8",X"20",X"38",X"18",X"00",X"60",X"F0",X"90",X"F0",X"7C",X"FC",X"00",X"00",
		X"00",X"08",X"7C",X"FC",X"88",X"C8",X"40",X"00",X"00",X"FC",X"FC",X"10",X"F0",X"E0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"38",X"7C",X"C2",X"82",X"86",X"7C",X"38",X"00",X"80",X"84",X"FE",X"FE",X"80",X"80",X"00",
		X"00",X"CC",X"E6",X"F2",X"B2",X"BA",X"9E",X"8C",X"00",X"40",X"C2",X"92",X"9A",X"9E",X"F6",X"62",
		X"00",X"30",X"38",X"2C",X"26",X"FE",X"FE",X"20",X"00",X"4E",X"CE",X"8A",X"8A",X"FA",X"70",X"00",
		X"00",X"78",X"FC",X"96",X"92",X"92",X"F2",X"60",X"00",X"06",X"06",X"E2",X"F2",X"1A",X"0E",X"06",
		X"00",X"6C",X"9E",X"9A",X"B2",X"B2",X"EC",X"60",X"00",X"0C",X"9E",X"92",X"92",X"D2",X"7E",X"3C",
		X"00",X"00",X"00",X"44",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"C0",X"80",X"80",X"80",X"FE",X"7E",X"00",X"7E",X"FE",X"80",X"80",X"80",X"FE",X"7E",
		X"00",X"FE",X"FE",X"1C",X"38",X"1C",X"FE",X"FE",X"00",X"FE",X"FE",X"22",X"22",X"22",X"3E",X"1C",
		X"FF",X"FF",X"F3",X"3E",X"00",X"FF",X"FF",X"00",X"FF",X"FF",X"F9",X"67",X"00",X"9F",X"FF",X"00",
		X"3F",X"9F",X"9B",X"8E",X"00",X"DC",X"BF",X"00",X"FC",X"FE",X"CE",X"72",X"00",X"FE",X"F8",X"00",
		X"FF",X"FF",X"F3",X"C9",X"81",X"00",X"0C",X"5C",X"1C",X"0C",X"89",X"80",X"C4",X"E1",X"E9",X"FF",
		X"7F",X"3F",X"1F",X"57",X"23",X"03",X"81",X"85",X"A0",X"B0",X"F0",X"F8",X"78",X"EA",X"E8",X"B0",
		X"F0",X"E1",X"41",X"03",X"03",X"07",X"8F",X"3F",X"FC",X"E0",X"C0",X"80",X"84",X"4F",X"0F",X"0F",
		X"07",X"03",X"0B",X"8F",X"8F",X"45",X"05",X"05",X"81",X"A0",X"80",X"C0",X"E0",X"E4",X"F8",X"FE",
		X"E7",X"C3",X"81",X"29",X"39",X"7C",X"7C",X"5E",X"F6",X"F6",X"FE",X"FE",X"FE",X"FE",X"FA",X"FE",
		X"FF",X"FF",X"FF",X"FF",X"FD",X"FD",X"FF",X"FF",X"FF",X"FB",X"F9",X"FD",X"FF",X"FF",X"FF",X"FF",
		X"03",X"C4",X"C7",X"BF",X"19",X"30",X"00",X"00",X"FF",X"FF",X"FF",X"FC",X"FC",X"FC",X"FE",X"FE",
		X"FF",X"FF",X"CF",X"BF",X"19",X"30",X"00",X"00",X"3F",X"1F",X"1F",X"1C",X"3C",X"7C",X"FE",X"FE",
		X"3F",X"7F",X"19",X"30",X"00",X"00",X"21",X"3F",X"FC",X"FC",X"FC",X"FC",X"FC",X"FE",X"FE",X"FE",
		X"3F",X"7F",X"19",X"30",X"00",X"80",X"E1",X"FF",X"FC",X"FC",X"FC",X"FC",X"FE",X"FF",X"FF",X"FF",
		X"CC",X"C4",X"84",X"C4",X"C2",X"C3",X"03",X"87",X"21",X"1F",X"1B",X"0E",X"00",X"DC",X"BF",X"00",
		X"0E",X"17",X"1F",X"1E",X"1F",X"0F",X"0F",X"07",X"07",X"05",X"03",X"03",X"03",X"03",X"03",X"03",
		X"03",X"03",X"03",X"03",X"07",X"07",X"06",X"0E",X"0C",X"14",X"1C",X"18",X"18",X"18",X"18",X"28",
		X"38",X"38",X"38",X"18",X"1C",X"1C",X"1E",X"0E",X"0C",X"0E",X"0E",X"06",X"0E",X"0E",X"0E",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"1F",X"17",X"03",X"83",X"83",X"87",X"87",X"CF",X"CF",X"87",X"C7",X"C7",X"C3",X"C3",X"03",X"87",
		X"87",X"8F",X"0F",X"0F",X"1F",X"1F",X"0F",X"0F",X"3F",X"1F",X"1F",X"1F",X"3F",X"7F",X"FF",X"FF",
		X"FF",X"7F",X"3F",X"3F",X"3F",X"7F",X"7F",X"3F",X"3F",X"1F",X"1F",X"0F",X"0F",X"0F",X"2F",X"3F",
		X"83",X"C4",X"C7",X"E7",X"E7",X"A7",X"87",X"87",X"82",X"C1",X"C0",X"C0",X"E8",X"F8",X"F8",X"F8",
		X"F0",X"E1",X"E1",X"E1",X"E1",X"C2",X"C3",X"83",X"03",X"04",X"07",X"0F",X"0F",X"1F",X"1B",X"0D",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3E",X"2F",X"1F",X"1F",X"1F",X"0B",X"0D",X"0F",X"0F",X"07",
		X"F0",X"F0",X"F0",X"F0",X"C0",X"F0",X"F0",X"70",X"F0",X"F8",X"F8",X"E8",X"D8",X"FC",X"FC",X"7C",
		X"B4",X"F8",X"F8",X"F8",X"F8",X"F8",X"E8",X"F0",X"F0",X"F0",X"E0",X"E0",X"C0",X"C0",X"C0",X"80",
		X"80",X"80",X"80",X"80",X"80",X"40",X"C0",X"C0",X"C0",X"C0",X"C0",X"A0",X"E0",X"E0",X"E0",X"F0",
		X"FE",X"FE",X"FF",X"FF",X"FF",X"FE",X"FE",X"FF",X"FE",X"FE",X"FC",X"FC",X"FC",X"FE",X"FE",X"FE",
		X"FF",X"FF",X"FE",X"FE",X"FC",X"FC",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"BF",X"9F",X"DF",X"FF",
		X"80",X"20",X"E0",X"70",X"F8",X"F8",X"FC",X"FC",X"7E",X"7E",X"7C",X"F8",X"68",X"0C",X"0C",X"0E",
		X"CF",X"87",X"C7",X"C4",X"C0",X"C0",X"02",X"86",X"FC",X"E0",X"C2",X"BC",X"18",X"30",X"00",X"00",
		X"FC",X"7C",X"3C",X"3C",X"3E",X"7F",X"7F",X"3F",X"30",X"7C",X"18",X"30",X"00",X"00",X"00",X"00",
		X"3E",X"1E",X"0A",X"00",X"00",X"00",X"00",X"00",X"87",X"8F",X"0F",X"0C",X"1C",X"1C",X"0E",X"0E",
		X"FF",X"FF",X"C3",X"BD",X"19",X"30",X"00",X"00",X"FC",X"7C",X"3C",X"3C",X"3E",X"7F",X"7F",X"3F",
		X"00",X"80",X"C0",X"E0",X"00",X"E0",X"E0",X"E0",X"37",X"7F",X"19",X"30",X"00",X"00",X"01",X"05",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",
		X"F0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FE",X"F8",X"C0",X"00",X"00",X"00",
		X"E0",X"C0",X"40",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"E0",
		X"80",X"C7",X"EF",X"E7",X"EF",X"CF",X"9E",X"80",X"FF",X"FC",X"E0",X"80",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FC",X"F0",X"80",X"00",X"C0",X"1C",X"7E",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"FE",X"FF",X"1F",X"03",X"00",X"80",X"C0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E2",X"FF",X"FE",X"FE",X"7C",X"3C",X"39",X"FB",X"0F",X"00",X"00",X"00",X"60",X"00",X"00",X"90",
		X"E0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FE",X"FC",X"F1",X"F7",X"7F",X"3F",
		X"81",X"CF",X"E7",X"F2",X"E7",X"E7",X"E3",X"E0",X"F0",X"F8",X"F8",X"E0",X"FC",X"FF",X"87",X"00",
		X"1F",X"3F",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"03",X"FE",X"7E",X"3E",X"1C",
		X"19",X"10",X"30",X"C1",X"81",X"02",X"0C",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"37",X"E0",X"06",
		X"F3",X"F1",X"E1",X"DF",X"FF",X"FF",X"FF",X"7F",X"7F",X"1F",X"7F",X"7F",X"7F",X"4F",X"03",X"00",
		X"00",X"00",X"00",X"C0",X"E0",X"E8",X"FC",X"FE",X"3C",X"03",X"01",X"20",X"78",X"30",X"10",X"10",
		X"D8",X"CC",X"86",X"00",X"03",X"FF",X"3E",X"00",X"F7",X"F7",X"F7",X"E1",X"E8",X"EE",X"CF",X"DE",
		X"80",X"E7",X"F3",X"F9",X"FD",X"FC",X"FE",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"FC",X"FD",X"F9",
		X"F0",X"F0",X"F0",X"E0",X"E8",X"EE",X"C0",X"C0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"F8",X"FE",X"F7",X"FB",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F3",X"3B",X"FB",X"FB",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"03",X"37",X"F7",
		X"00",X"04",X"07",X"7F",X"FF",X"FD",X"7F",X"7F",X"0F",X"7F",X"7B",X"3B",X"BF",X"9F",X"DF",X"DF",
		X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"6E",X"EE",X"E7",X"F7",X"37",
		X"E7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"09",X"15",X"74",X"F6",
		X"00",X"00",X"00",X"1F",X"FB",X"DD",X"BF",X"FF",X"00",X"1F",X"53",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"07",X"3F",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"07",X"1F",X"7F",X"FF",
		X"00",X"00",X"00",X"00",X"01",X"07",X"1F",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"07",X"1F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"07",X"1F",X"7F",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"01",X"07",X"1F",X"7F",X"FF",X"0E",X"1B",X"39",X"10",X"09",X"01",X"04",X"00",
		X"00",X"00",X"00",X"01",X"0F",X"7F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"03",X"1F",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",
		X"00",X"00",X"00",X"01",X"07",X"3F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"03",X"3F",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"30",X"18",X"18",X"0C",X"54",X"80",X"AC",X"04",
		X"00",X"00",X"00",X"00",X"0F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"03",X"3F",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"07",X"1F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"01",X"07",X"0F",X"1F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"07",X"07",X"07",
		X"07",X"07",X"07",X"07",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"F8",X"FC",X"FE",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"C0",X"C0",X"E0",X"E0",
		X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"04",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"F0",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"80",X"F0",X"FE",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",
		X"00",X"00",X"80",X"C0",X"E0",X"F0",X"F8",X"E0",X"00",X"00",X"80",X"C0",X"E0",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"E0",X"F8",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"F8",X"FF",X"FC",X"F0",X"80",X"00",X"00",X"00",
		X"F0",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"C0",X"F0",X"FC",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",X"F8",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"80",X"E0",X"F0",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"F0",X"F8",X"FC",
		X"10",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"00",X"00",X"0F",X"1F",X"1F",X"3F",X"7F",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"1F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"1F",
		X"00",X"60",X"FC",X"FF",X"FF",X"FF",X"DF",X"A1",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"C0",X"F0",X"F0",X"88",X"04",X"00",X"00",X"07",X"7F",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"01",X"1F",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"C0",X"00",X"60",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"80",X"00",X"00",X"07",X"3F",X"FF",X"FF",
		X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"1F",X"F8",X"C0",X"00",X"00",X"03",X"1F",
		X"00",X"00",X"01",X"1F",X"FF",X"FF",X"FF",X"FF",X"01",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"01",X"1F",X"FF",X"FF",X"00",X"00",X"00",X"07",X"7F",X"FF",X"FF",X"FF",
		X"06",X"01",X"01",X"60",X"00",X"18",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"3F",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"00",X"00",X"00",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"00",X"01",X"CF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"83",
		X"00",X"00",X"20",X"A0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"70",X"F8",X"F0",X"F0",X"C0",X"40",X"18",X"00",
		X"00",X"00",X"00",X"00",X"04",X"08",X"01",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"21",X"80",X"40",X"00",X"00",X"00",X"00",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"12",X"7A",X"7C",
		X"38",X"6C",X"42",X"00",X"30",X"68",X"C1",X"C1",X"00",X"00",X"1E",X"72",X"F9",X"A8",X"00",X"06",
		X"00",X"00",X"00",X"00",X"30",X"78",X"2C",X"04",X"7D",X"FD",X"7F",X"FC",X"FC",X"78",X"78",X"F8",
		X"80",X"C0",X"80",X"80",X"40",X"00",X"00",X"00",X"03",X"07",X"0E",X"1A",X"08",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"04",X"84",X"C0",X"41",X"01",X"02",X"00",X"00",
		X"E8",X"1C",X"12",X"04",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"03",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"EF",X"FE",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FE",X"FF",X"FF",X"E7",X"FF",X"FE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BF",X"2F",X"6E",X"78",X"00",X"00",X"40",X"40",
		X"FF",X"FF",X"FF",X"FF",X"EF",X"E7",X"16",X"70",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FC",X"EE",X"FE",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"FF",X"FF",X"00",X"01",X"07",X"1F",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"1F",X"00",X"01",X"07",X"1F",X"7F",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"1F",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"C0",X"E0",X"E0",X"E0",
		X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",X"FC",X"FC",X"FE",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"E0",X"F0",X"FC",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",X"EF",X"EB",X"EF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",X"FB",X"FB",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FB",X"FB",X"B3",X"D7",X"F7",X"03",X"01",X"00",
		X"FF",X"FF",X"FF",X"BF",X"7D",X"FB",X"FE",X"00",X"BF",X"9F",X"DF",X"DF",X"DF",X"87",X"01",X"00",
		X"BF",X"BF",X"F6",X"FC",X"F9",X"83",X"3F",X"7F",X"7F",X"7F",X"7F",X"7F",X"3F",X"1F",X"0F",X"07",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"07",X"07",X"03",X"03",X"03",X"03",X"03",X"03",
		X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"FE",X"FE",X"FF",X"FF",X"C0",X"FF",X"FF",X"FF",
		X"FF",X"7F",X"7E",X"78",X"00",X"C0",X"C0",X"C0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"80",X"80",X"80",X"80",X"80",X"80",X"C0",X"C0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"C0",X"C0",X"C0",X"E0",X"E0",X"E0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F8",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"F8",X"FC",X"FC",X"FC",X"FC",X"FE",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"7F",X"77",X"6F",X"7C",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"F3",X"FB",X"9B",X"FA",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"F3",X"FE",X"7C",
		X"78",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"77",X"37",X"BC",X"A0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"F7",X"F3",X"3B",X"FB",X"FA",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FE",X"FE",X"FE",X"FF",X"F3",X"FF",X"7C",
		X"78",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FC",X"EF",X"6F",X"7C",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"ED",X"ED",X"E7",X"F4",X"70",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"55",X"FF",X"55",X"FF",X"55",X"FF",X"FF",
		X"FF",X"55",X"FF",X"55",X"FF",X"55",X"FF",X"00",X"FC",X"4A",X"FF",X"4B",X"FD",X"4B",X"FC",X"00",
		X"00",X"00",X"00",X"80",X"F8",X"80",X"00",X"00",X"01",X"01",X"FF",X"55",X"FF",X"55",X"FF",X"FF",
		X"01",X"01",X"0F",X"05",X"1F",X"15",X"3F",X"00",X"00",X"00",X"FF",X"55",X"FF",X"55",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"B8",X"EF",X"01",X"00",X"0F",X"04",X"1F",X"04",X"3F",X"00",
		X"B9",X"EF",X"B9",X"EF",X"B9",X"E7",X"00",X"00",X"FF",X"92",X"FF",X"92",X"FF",X"92",X"FF",X"00",
		X"00",X"10",X"38",X"38",X"38",X"38",X"10",X"00",X"00",X"00",X"00",X"80",X"80",X"F8",X"FC",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"01",X"03",X"07",X"0F",X"FF",X"55",
		X"87",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"C0",X"80",X"D1",X"BF",X"D1",X"BF",X"C1",X"60",
		X"00",X"00",X"80",X"C0",X"E0",X"80",X"00",X"00",X"FC",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"4A",X"FF",X"4B",X"FD",X"4B",X"FF",X"4B",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"00",X"FD",X"4B",X"FF",X"4B",X"FD",X"4B",X"FC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"4A",X"FF",X"4B",X"FD",X"4B",X"FC",X"00",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"00",X"00",X"55",X"FF",X"FF",X"55",X"FF",X"00",
		X"E0",X"E0",X"E0",X"00",X"00",X"00",X"00",X"00",X"FF",X"24",X"FF",X"24",X"FF",X"24",X"FF",X"00",
		X"FF",X"92",X"FF",X"92",X"FF",X"92",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"80",
		X"FF",X"07",X"07",X"07",X"07",X"07",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"A0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"4A",X"FF",X"4B",X"FD",X"4B",X"FC",X"00",
		X"FC",X"4A",X"FF",X"49",X"FD",X"4B",X"FC",X"00",X"01",X"01",X"FF",X"55",X"FF",X"55",X"FF",X"FF",
		X"FF",X"55",X"FF",X"55",X"FF",X"55",X"FF",X"FF",X"FF",X"55",X"FF",X"55",X"FF",X"55",X"FF",X"00",
		X"01",X"01",X"0F",X"05",X"1F",X"15",X"3F",X"00",X"FC",X"4A",X"FF",X"4B",X"FD",X"4B",X"FF",X"49",
		X"F8",X"F8",X"FF",X"F8",X"F0",X"00",X"00",X"00",X"FD",X"4B",X"FF",X"4B",X"FD",X"4B",X"FC",X"00",
		X"01",X"00",X"FF",X"24",X"FF",X"24",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"0F",X"04",X"1F",X"04",X"3F",X"00",X"00",X"00",X"80",X"C0",X"E0",X"80",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"55",X"FF",X"55",X"FF",X"55",X"FF",X"FF",X"00",X"55",X"FF",X"55",X"FF",X"55",X"FF",X"00",
		X"FF",X"55",X"FF",X"55",X"FF",X"55",X"FF",X"00",X"01",X"01",X"FF",X"55",X"FF",X"55",X"FF",X"FF",
		X"F5",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"55",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"F0",X"F8",X"FF",X"F8",X"F8",X"00",X"00",X"00",X"00",X"00",X"2A",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",X"00",X"FC",X"48",X"FC",X"4A",X"FC",X"48",X"FC",X"00",
		X"01",X"00",X"FF",X"24",X"FF",X"24",X"FF",X"00",X"FC",X"4A",X"FF",X"4B",X"FD",X"4B",X"FC",X"00",
		X"00",X"B2",X"03",X"B5",X"01",X"B3",X"03",X"B5",X"00",X"6D",X"00",X"6D",X"00",X"6D",X"00",X"00",
		X"00",X"B2",X"03",X"B5",X"01",X"B3",X"00",X"00",X"01",X"B3",X"03",X"B5",X"01",X"B3",X"00",X"00",
		X"01",X"00",X"0F",X"04",X"1F",X"04",X"3F",X"00",X"FF",X"92",X"FF",X"92",X"FF",X"92",X"FF",X"00",
		X"00",X"00",X"FF",X"55",X"FF",X"55",X"FF",X"00",X"00",X"03",X"00",X"0B",X"00",X"1B",X"00",X"00",
		X"00",X"DB",X"00",X"DB",X"00",X"DB",X"00",X"00",X"00",X"00",X"80",X"E0",X"E0",X"00",X"00",X"00",
		X"00",X"00",X"80",X"E0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"24",X"FF",X"24",X"FF",X"24",X"FF",X"00",X"00",X"03",X"00",X"DB",X"00",X"DB",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"AA",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"FF",X"ED",X"FC",X"FC",X"00",X"00",X"00",X"00",X"8F",X"E7",X"75",X"00",
		X"00",X"00",X"1F",X"E1",X"FC",X"CE",X"E3",X"F8",X"00",X"00",X"81",X"E0",X"70",X"30",X"30",X"11",
		X"03",X"FD",X"80",X"00",X"00",X"00",X"00",X"C0",X"20",X"B8",X"90",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"BC",X"28",X"23",X"83",X"87",X"9F",X"BF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"80",X"40",X"60",X"10",X"08",
		X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"12",X"0A",X"1A",X"1A",X"1A",X"18",
		X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"0C",X"12",X"1A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"12",X"1A",X"1A",
		X"80",X"A0",X"20",X"20",X"30",X"20",X"80",X"B0",X"00",X"06",X"E9",X"46",X"E0",X"0F",X"C8",X"60",
		X"00",X"00",X"00",X"28",X"00",X"10",X"54",X"10",X"CF",X"09",X"E6",X"80",X"0F",X"ED",X"88",X"00",
		X"1E",X"08",X"1E",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"04",X"08",X"08",X"01",X"12",X"12",
		X"E0",X"18",X"06",X"01",X"F0",X"08",X"04",X"04",X"10",X"10",X"10",X"10",X"14",X"14",X"14",X"10",
		X"06",X"05",X"04",X"04",X"02",X"02",X"02",X"03",X"14",X"14",X"14",X"12",X"12",X"1A",X"16",X"12",
		X"02",X"02",X"02",X"04",X"04",X"05",X"06",X"04",X"E0",X"F0",X"38",X"D8",X"F8",X"38",X"58",X"38",
		X"00",X"00",X"00",X"00",X"00",X"40",X"90",X"A8",X"12",X"11",X"18",X"18",X"1C",X"1F",X"0F",X"0F",
		X"04",X"08",X"F0",X"01",X"06",X"1F",X"E6",X"07",X"F8",X"B8",X"58",X"F8",X"18",X"F8",X"18",X"38",
		X"48",X"00",X"D0",X"00",X"F0",X"00",X"E0",X"40",X"1E",X"1E",X"1C",X"1C",X"19",X"18",X"03",X"00",
		X"46",X"07",X"C7",X"06",X"87",X"03",X"01",X"00",X"19",X"F8",X"38",X"D8",X"38",X"F0",X"E0",X"00",
		X"20",X"80",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",
		X"00",X"01",X"03",X"47",X"6C",X"3B",X"70",X"00",X"07",X"FB",X"FF",X"0D",X"FF",X"FF",X"79",X"00",
		X"00",X"C0",X"E0",X"E4",X"E4",X"F4",X"F8",X"70",X"07",X"06",X"07",X"03",X"03",X"03",X"03",X"01",
		X"00",X"00",X"3F",X"3F",X"DF",X"DF",X"0F",X"E0",X"30",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"00",X"00",X"08",X"38",X"1C",X"38",X"08",X"00",X"01",X"00",X"01",X"01",X"01",X"01",X"01",X"01",
		X"F8",X"00",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FE",X"FD",X"FB",X"02",X"FB",X"00",X"00",X"40",X"80",X"60",X"80",X"00",X"F0",
		X"01",X"03",X"03",X"03",X"03",X"07",X"07",X"07",X"D2",X"F5",X"E6",X"ED",X"CA",X"CA",X"89",X"89",
		X"00",X"80",X"60",X"00",X"80",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"07",X"0F",
		X"00",X"00",X"02",X"06",X"06",X"0F",X"0F",X"4F",X"A0",X"70",X"70",X"20",X"80",X"C0",X"80",X"F0",
		X"00",X"00",X"00",X"00",X"08",X"1C",X"1C",X"08",X"1F",X"11",X"15",X"5F",X"11",X"1F",X"11",X"53",
		X"F0",X"EC",X"D8",X"D8",X"B4",X"A8",X"A8",X"B4",X"00",X"00",X"00",X"C0",X"F0",X"F8",X"F8",X"C0",
		X"00",X"06",X"03",X"00",X"00",X"00",X"00",X"00",X"1F",X"11",X"35",X"3F",X"71",X"73",X"FF",X"07",
		X"B8",X"D8",X"DC",X"EC",X"F0",X"F0",X"F4",X"FC",X"00",X"00",X"00",X"08",X"1C",X"1C",X"08",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"18",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"E1",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"F0",X"FC",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"3F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"F0",X"FC",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"9F",X"9F",X"9F",X"8F",X"CF",X"CF",X"CF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CF",X"CF",X"C7",X"E7",X"E7",X"E7",X"E7",X"E7",
		X"FF",X"FF",X"CF",X"E3",X"FB",X"FB",X"FB",X"FB",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"F0",X"F0",
		X"E3",X"F3",X"F3",X"F3",X"F3",X"F3",X"F1",X"F9",X"DB",X"C3",X"C3",X"C3",X"C3",X"C3",X"C3",X"C3",
		X"F0",X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",X"F9",X"F9",X"F9",X"F9",X"F8",X"FC",X"9C",X"C4",
		X"C3",X"C3",X"E3",X"FB",X"FB",X"FB",X"FB",X"FF",X"F8",X"F8",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"FF",X"FF",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"F4",X"F4",X"F4",X"F6",X"B6",X"86",X"86",X"86",
		X"FE",X"FE",X"FE",X"FF",X"FF",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"0F",X"03",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"80",X"E0",X"FF",X"FF",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"7F",X"1F",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F8",X"F8",X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"3F",X"3F",X"1F",X"1F",X"3F",X"3F",X"3F",
		X"86",X"87",X"87",X"87",X"87",X"87",X"C7",X"F6",X"F6",X"F6",X"F6",X"FC",X"FC",X"FC",X"FC",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"C0",X"00",X"3C",X"8E",X"E0",X"00",
		X"FF",X"0F",X"E3",X"38",X"00",X"FF",X"00",X"00",X"FF",X"C0",X"FF",X"00",X"0F",X"03",X"00",X"00",
		X"FF",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"70",X"1C",X"FF",X"00",X"00",X"00",X"00",
		X"01",X"FC",X"FF",X"FF",X"00",X"00",X"00",X"00",X"E0",X"3F",X"0F",X"03",X"00",X"00",X"00",X"00",
		X"FF",X"03",X"00",X"00",X"00",X"C0",X"F0",X"FC",X"FF",X"C0",X"F0",X"FC",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F3",X"F8",X"FE",X"FE",X"FE",X"FE",X"F6",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F8",X"FE",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"8F",X"63",X"00",X"01",X"07",X"FF",X"FF",X"FF",X"C7",X"F0",X"FC",X"FC",X"FC",
		X"FF",X"BF",X"BF",X"BF",X"9F",X"9F",X"9F",X"8F",X"8F",X"8F",X"87",X"87",X"87",X"83",X"83",X"83",
		X"81",X"81",X"81",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"3F",X"3F",X"3F",X"1F",X"1F",X"1F",X"0F",
		X"0F",X"0F",X"07",X"07",X"07",X"03",X"03",X"03",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"3F",X"3F",X"3F",X"3F",X"1F",X"1F",X"1F",X"1F",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",
		X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",
		X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FE",X"07",X"07",X"87",X"87",X"C7",X"E7",X"E7",X"F7",
		X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"F8",X"F8",X"F8",X"F8",X"78",X"78",X"F8",
		X"7F",X"1F",X"07",X"FF",X"FF",X"00",X"00",X"00",X"F8",X"F8",X"F8",X"7F",X"1F",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"07",X"07",X"07",X"07",X"03",X"03",X"03",X"03",X"01",X"01",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"3F",X"0F",X"03",X"00",X"3F",X"0F",X"03",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"04",X"00",X"20",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"00",X"00",X"60",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"70",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"E0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"03",X"0F",X"0C",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"60",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",
		X"0F",X"1E",X"7C",X"F0",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"0F",X"1F",X"7E",X"FC",X"F0",X"E0",X"80",X"00",X"00",
		X"00",X"00",X"01",X"03",X"0F",X"1F",X"7F",X"FC",X"03",X"0F",X"1F",X"3F",X"3E",X"38",X"30",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"08",X"18",X"78",X"F8",X"F8",X"F8",X"F0",X"E0",X"80",X"00",X"00",
		X"01",X"03",X"0F",X"1F",X"7F",X"FF",X"FF",X"FC",X"1F",X"7F",X"FF",X"FF",X"FE",X"F8",X"F0",X"C0",
		X"00",X"00",X"01",X"03",X"0F",X"1F",X"7F",X"FF",X"00",X"00",X"04",X"00",X"20",X"00",X"00",X"00",
		X"01",X"00",X"00",X"40",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"0F",X"1C",
		X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"C0",X"C0",
		X"00",X"00",X"00",X"01",X"03",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",
		X"1C",X"7C",X"FC",X"F0",X"E0",X"80",X"00",X"00",X"03",X"0F",X"1F",X"7F",X"FE",X"F8",X"F0",X"C0",
		X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"04",X"00",X"40",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"01",X"00",X"00",X"60",X"C0",X"01",X"00",X"00",X"00",X"80",X"80",X"00",X"00",
		X"38",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"03",X"0F",X"0F",X"0C",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"60",X"E0",X"E0",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"0F",X"0F",
		X"0F",X"0E",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"08",X"18",X"78",X"F8",X"F8",X"F8",X"00",X"00",X"04",X"00",X"60",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"04",X"03",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"78",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",
		X"0E",X"1E",X"7C",X"F0",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"0F",X"1F",X"3C",
		X"38",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"00",X"00",
		X"7F",X"7E",X"7C",X"70",X"60",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"60",X"00",X"00",X"00",
		X"00",X"00",X"01",X"03",X"02",X"00",X"40",X"C0",X"03",X"06",X"04",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"0E",X"1C",X"78",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"1C",X"7C",X"F0",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"0F",X"1F",X"7C",
		X"00",X"00",X"01",X"03",X"03",X"03",X"03",X"00",X"00",X"01",X"03",X"07",X"07",X"07",X"07",X"04",
		X"10",X"70",X"F0",X"F0",X"F0",X"F0",X"F0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"0C",
		X"08",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"00",X"00",
		X"00",X"10",X"70",X"F0",X"E0",X"80",X"00",X"00",X"01",X"03",X"03",X"03",X"02",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"E0",X"E0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"03",X"0F",X"1F",X"7F",X"7F",X"7C",X"78",X"60",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"02",X"0E",X"1E",X"7E",X"FE",X"00",X"00",X"0C",X"00",X"40",X"00",X"00",X"00",
		X"00",X"00",X"01",X"03",X"06",X"00",X"00",X"80",X"03",X"0E",X"0C",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"1C",X"00",X"01",X"03",X"07",X"06",X"00",X"00",X"00",
		X"00",X"00",X"60",X"E0",X"E0",X"80",X"00",X"00",X"01",X"03",X"0F",X"0F",X"0E",X"08",X"00",X"00",
		X"07",X"07",X"07",X"07",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"C0",
		X"00",X"02",X"08",X"00",X"40",X"80",X"00",X"00",X"00",X"00",X"01",X"03",X"06",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"18",X"00",X"01",X"03",X"0F",X"0E",X"08",X"00",X"00",
		X"00",X"00",X"00",X"80",X"80",X"80",X"00",X"00",X"01",X"03",X"0F",X"1F",X"3E",X"38",X"30",X"00",
		X"00",X"08",X"18",X"78",X"F8",X"F8",X"F0",X"C0",X"0F",X"1F",X"7F",X"7F",X"7E",X"78",X"70",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"03",X"0F",X"0F",X"0F",X"0F",X"0F",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0E",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"03",X"0F",X"0F",X"0F",X"0F",X"02",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"0F",X"1F",X"7F",X"FF",X"FF",X"FF",X"FC",
		X"00",X"00",X"10",X"70",X"F0",X"F0",X"F0",X"F0",X"C0",X"F1",X"F3",X"FF",X"F3",X"FD",X"F1",X"FD",
		X"00",X"60",X"78",X"FC",X"7C",X"FE",X"7F",X"7F",X"00",X"00",X"00",X"00",X"00",X"02",X"0E",X"1E",
		X"7F",X"FF",X"FF",X"FF",X"FE",X"F8",X"F0",X"C0",X"7E",X"FE",X"FE",X"FE",X"FE",X"F8",X"F0",X"C0",
		X"40",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"00",X"01",X"03",X"0F",X"1F",X"7F",X"FF",X"FF",
		X"00",X"00",X"00",X"08",X"18",X"78",X"F8",X"F8",X"F8",X"F8",X"F8",X"F0",X"E0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"F0",X"B1",X"AD",X"A1",X"80",X"00",X"0E",X"3F",X"D5",
		X"FE",X"7E",X"7C",X"3C",X"38",X"BF",X"FF",X"55",X"30",X"18",X"18",X"0C",X"54",X"80",X"AC",X"04",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"8F",X"C4",X"60",X"30",X"30",X"11",X"00",X"00",X"00",X"00",X"E0",X"30",X"18",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"41",X"81",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"A0",X"B8",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"18",X"06",X"01",X"F0",X"08",X"64",X"94",
		X"06",X"E5",X"54",X"E4",X"02",X"A2",X"52",X"03",X"F2",X"02",X"F2",X"64",X"F4",X"05",X"66",X"94",
		X"64",X"08",X"F0",X"01",X"06",X"1F",X"E6",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"01",X"03",X"03",X"81",X"C0",X"80",X"F0",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"C2",X"F7",X"FF",X"FA",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F1",X"F3",X"1B",X"09",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"20",X"20",X"40",X"40",X"40",X"40",
		X"00",X"18",X"3C",X"3C",X"7E",X"7E",X"7E",X"7E",X"40",X"40",X"00",X"30",X"12",X"1F",X"07",X"00",
		X"7E",X"7E",X"3E",X"BE",X"D8",X"D8",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"5B",X"7F",
		X"00",X"00",X"07",X"1F",X"38",X"00",X"58",X"FC",X"00",X"00",X"00",X"80",X"C0",X"40",X"00",X"30",
		X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"7F",X"FF",X"FF",X"FD",X"7C",X"78",X"FA",X"F2",
		X"F8",X"D0",X"45",X"0F",X"1F",X"1E",X"3C",X"3C",X"18",X"0C",X"C4",X"E0",X"30",X"10",X"00",X"00",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"F3",X"F3",X"E1",X"61",X"70",X"20",X"20",X"20",
		X"18",X"39",X"33",X"13",X"01",X"21",X"60",X"E0",X"F0",X"E0",X"F8",X"F0",X"FC",X"F0",X"A0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"06",X"06",X"03",X"13",X"1B",X"0B",X"01",
		X"A7",X"33",X"10",X"02",X"01",X"00",X"00",X"00",X"24",X"FE",X"CC",X"00",X"C0",X"E0",X"70",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"3F",X"3F",X"7F",X"F7",
		X"00",X"00",X"00",X"C0",X"F0",X"F8",X"FC",X"DE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",
		X"01",X"01",X"00",X"00",X"01",X"01",X"03",X"03",X"FF",X"FE",X"FF",X"FF",X"F7",X"FF",X"BF",X"FE",
		X"FF",X"F7",X"FF",X"FF",X"DF",X"FD",X"FF",X"FF",X"E0",X"E0",X"F0",X"B8",X"F8",X"F8",X"FC",X"FC",
		X"01",X"01",X"01",X"03",X"03",X"01",X"01",X"00",X"FF",X"FF",X"EF",X"FF",X"FF",X"FD",X"DF",X"FF",
		X"F7",X"FF",X"BF",X"FF",X"FF",X"ED",X"FF",X"FF",X"78",X"F0",X"F0",X"F0",X"B8",X"F8",X"F8",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"38",X"10",X"00",X"00",X"00",X"00",
		X"BF",X"FF",X"6F",X"07",X"03",X"01",X"00",X"00",X"F0",X"70",X"F0",X"E0",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"18",X"18",X"00",X"00",X"00",X"00",X"20",X"20",X"00",X"0F",X"65",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"E0",X"00",X"01",X"03",X"03",X"01",X"00",X"06",X"33",
		X"FF",X"B8",X"FF",X"FF",X"FD",X"FF",X"7F",X"FF",X"38",X"F8",X"2C",X"8C",X"C4",X"E8",X"F0",X"F0",
		X"7A",X"78",X"77",X"5F",X"0E",X"6E",X"27",X"07",X"FF",X"FF",X"FF",X"FD",X"FC",X"5E",X"EE",X"FC",
		X"F8",X"FC",X"FC",X"FC",X"FC",X"BC",X"D8",X"30",X"07",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FF",X"7F",X"E2",X"00",X"00",X"00",X"00",X"00",X"04",X"0E",X"1A",X"36",X"7E",X"3C",X"00",
		X"00",X"00",X"00",X"00",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"60",X"20",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"0E",X"0F",X"1F",X"3B",X"17",X"1F",
		X"EF",X"F7",X"7F",X"3F",X"FF",X"FF",X"FF",X"FF",X"00",X"40",X"70",X"F8",X"7C",X"7E",X"7B",X"5F",
		X"0F",X"C5",X"F7",X"73",X"53",X"72",X"33",X"01",X"61",X"33",X"9E",X"9C",X"8F",X"C0",X"FF",X"FF",
		X"DF",X"BF",X"0F",X"8F",X"86",X"6C",X"E0",X"F0",X"01",X"08",X"0E",X"07",X"03",X"00",X"00",X"00",
		X"EF",X"7D",X"00",X"82",X"CF",X"E7",X"3C",X"00",X"B0",X"D8",X"C8",X"00",X"E1",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"03",X"3B",X"7F",X"00",X"00",X"50",X"F8",X"FF",X"FF",X"F7",X"F6",
		X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"7F",X"7F",X"7F",X"3F",X"1F",X"07",X"01",X"00",
		X"CE",X"E3",X"F8",X"FC",X"EF",X"FF",X"FD",X"FF",X"C0",X"E0",X"C0",X"00",X"80",X"80",X"F8",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DE",X"D7",X"F0",X"F0",X"F8",X"FE",X"73",X"7F",
		X"BC",X"FE",X"FC",X"5E",X"14",X"00",X"80",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3E",X"1F",X"07",X"01",X"00",X"00",X"00",X"00",X"70",X"F0",X"E0",X"F0",X"20",X"00",X"00",X"00",
		X"00",X"00",X"03",X"07",X"0F",X"1F",X"1F",X"3F",X"07",X"FF",X"FF",X"F0",X"C0",X"80",X"00",X"00",
		X"80",X"E0",X"F8",X"3C",X"7E",X"1F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"3E",X"7E",X"0C",X"0C",X"0C",X"1C",X"18",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"07",X"03",X"03",X"03",X"03",X"00",X"00",X"80",X"C0",X"C0",X"C0",X"C0",X"E0",X"60",X"60",
		X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",
		X"00",X"60",X"FC",X"FF",X"FF",X"FF",X"DF",X"A1",X"00",X"00",X"00",X"C0",X"F0",X"F0",X"88",X"04",
		X"00",X"00",X"00",X"00",X"C0",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"78",X"7E",X"38",X"6C",X"42",X"00",X"30",X"68",X"C1",X"C1",
		X"00",X"00",X"1E",X"72",X"F9",X"A8",X"00",X"06",X"00",X"00",X"00",X"00",X"30",X"78",X"2C",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"60",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"40",X"21",X"80",X"40",X"00",X"00",X"0F",X"8F",X"80",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"C2",X"E7",
		X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
