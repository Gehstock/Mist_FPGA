-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

entity ROM_PGM_1 is
  port (
    CLK         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM_1 is


  type ROM_ARRAY is array(0 to 16383) of std_logic_vector(7 downto 0);
  constant ROM : ROM_ARRAY := (
    x"C3",x"01",x"01",x"00",x"00",x"00",x"00",x"00", -- 0x0000
    x"77",x"23",x"10",x"FC",x"C9",x"00",x"00",x"00", -- 0x0008
    x"85",x"6F",x"8C",x"95",x"67",x"7E",x"C9",x"00", -- 0x0010
    x"78",x"87",x"D7",x"5F",x"23",x"56",x"EB",x"C9", -- 0x0018
    x"E1",x"87",x"D7",x"5F",x"23",x"56",x"EB",x"E9", -- 0x0020
    x"ED",x"B0",x"AF",x"32",x"C0",x"50",x"C9",x"00", -- 0x0028
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0030
    x"C3",x"68",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0038
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0040
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0048
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0050
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0058
    x"00",x"00",x"00",x"00",x"00",x"00",x"ED",x"45", -- 0x0060
    x"F3",x"F5",x"DD",x"E5",x"E5",x"D5",x"C5",x"AF", -- 0x0068
    x"32",x"00",x"50",x"32",x"C0",x"50",x"2A",x"00", -- 0x0070
    x"4C",x"23",x"22",x"00",x"4C",x"3E",x"00",x"B7", -- 0x0078
    x"C2",x"EE",x"00",x"21",x"53",x"4C",x"11",x"F2", -- 0x0080
    x"4F",x"01",x"0C",x"00",x"EF",x"11",x"04",x"00", -- 0x0088
    x"19",x"11",x"62",x"50",x"01",x"0C",x"00",x"EF", -- 0x0090
    x"3A",x"1B",x"4C",x"3C",x"32",x"1B",x"4C",x"E6", -- 0x0098
    x"01",x"28",x"1C",x"2A",x"51",x"4C",x"ED",x"5B", -- 0x00A0
    x"61",x"4C",x"22",x"FA",x"4F",x"ED",x"53",x"6A", -- 0x00A8
    x"50",x"2A",x"5F",x"4C",x"ED",x"5B",x"6F",x"4C", -- 0x00B0
    x"22",x"FC",x"4F",x"ED",x"53",x"6C",x"50",x"3A", -- 0x00B8
    x"50",x"4C",x"B7",x"28",x"14",x"AF",x"32",x"1C", -- 0x00C0
    x"4C",x"AF",x"32",x"50",x"4C",x"CD",x"DD",x"0C", -- 0x00C8
    x"CD",x"DC",x"0C",x"CD",x"B7",x"0C",x"CD",x"92", -- 0x00D0
    x"07",x"CD",x"AF",x"12",x"AF",x"32",x"C0",x"50", -- 0x00D8
    x"3E",x"01",x"32",x"00",x"50",x"C1",x"D1",x"E1", -- 0x00E0
    x"DD",x"E1",x"F1",x"FB",x"ED",x"4D",x"21",x"51", -- 0x00E8
    x"4C",x"11",x"F0",x"4F",x"01",x"10",x"00",x"EF", -- 0x00F0
    x"11",x"60",x"50",x"01",x"10",x"00",x"EF",x"18", -- 0x00F8
    x"BE",x"F3",x"31",x"F0",x"4F",x"ED",x"56",x"3E", -- 0x0100
    x"FF",x"D3",x"00",x"AF",x"21",x"00",x"50",x"01", -- 0x0108
    x"08",x"08",x"CF",x"AF",x"32",x"C0",x"50",x"21", -- 0x0110
    x"00",x"4C",x"06",x"BE",x"CF",x"CF",x"CF",x"CF", -- 0x0118
    x"3E",x"0F",x"32",x"4C",x"4C",x"32",x"4D",x"4C", -- 0x0120
    x"21",x"0D",x"4C",x"11",x"0E",x"4C",x"01",x"0C", -- 0x0128
    x"00",x"36",x"30",x"EF",x"AF",x"12",x"32",x"13", -- 0x0130
    x"4C",x"21",x"CE",x"FA",x"22",x"02",x"4C",x"21", -- 0x0138
    x"40",x"50",x"06",x"40",x"CF",x"3E",x"01",x"32", -- 0x0140
    x"00",x"50",x"FB",x"AF",x"32",x"C0",x"50",x"32", -- 0x0148
    x"48",x"4C",x"32",x"49",x"4C",x"32",x"4A",x"4C", -- 0x0150
    x"3E",x"01",x"32",x"1D",x"4C",x"3E",x"68",x"32", -- 0x0158
    x"1E",x"4C",x"3E",x"00",x"32",x"1F",x"4C",x"3E", -- 0x0160
    x"01",x"32",x"20",x"4C",x"AF",x"32",x"24",x"4C", -- 0x0168
    x"32",x"22",x"4C",x"3E",x"FF",x"32",x"25",x"4C", -- 0x0170
    x"AF",x"32",x"50",x"4C",x"32",x"48",x"4C",x"32", -- 0x0178
    x"49",x"4C",x"32",x"4A",x"4C",x"3E",x"01",x"CD", -- 0x0180
    x"A2",x"12",x"CD",x"24",x"0F",x"3A",x"0B",x"4C", -- 0x0188
    x"B7",x"20",x"14",x"21",x"D9",x"11",x"11",x"BC", -- 0x0190
    x"43",x"0E",x"01",x"CD",x"93",x"0B",x"CD",x"83", -- 0x0198
    x"0B",x"3A",x"0B",x"4C",x"B7",x"28",x"F7",x"21", -- 0x01A0
    x"BD",x"11",x"11",x"BC",x"43",x"0E",x"01",x"CD", -- 0x01A8
    x"93",x"0B",x"CD",x"83",x"0B",x"3A",x"09",x"4C", -- 0x01B0
    x"E6",x"20",x"28",x"F6",x"3A",x"0B",x"4C",x"3D", -- 0x01B8
    x"32",x"0B",x"4C",x"3E",x"02",x"CD",x"A2",x"12", -- 0x01C0
    x"3E",x"00",x"32",x"2F",x"4C",x"3E",x"05",x"32", -- 0x01C8
    x"27",x"4C",x"21",x"0D",x"4C",x"11",x"0E",x"4C", -- 0x01D0
    x"01",x"05",x"00",x"36",x"30",x"EF",x"AF",x"12", -- 0x01D8
    x"3A",x"2F",x"4C",x"CD",x"1B",x"0D",x"AF",x"32", -- 0x01E0
    x"24",x"4C",x"CD",x"E2",x"26",x"AF",x"32",x"2B", -- 0x01E8
    x"4C",x"3A",x"30",x"4C",x"3C",x"32",x"30",x"4C", -- 0x01F0
    x"3E",x"01",x"32",x"0A",x"4C",x"CD",x"83",x"0B", -- 0x01F8
    x"CD",x"83",x"0B",x"CD",x"83",x"0B",x"AF",x"32", -- 0x0200
    x"0A",x"4C",x"CD",x"83",x"0B",x"3A",x"2E",x"4C", -- 0x0208
    x"3C",x"FE",x"06",x"38",x"0F",x"CD",x"3C",x"0B", -- 0x0210
    x"3A",x"39",x"4C",x"B7",x"20",x"05",x"3E",x"02", -- 0x0218
    x"32",x"2B",x"4C",x"AF",x"32",x"2E",x"4C",x"3A", -- 0x0220
    x"31",x"4C",x"32",x"33",x"4C",x"3A",x"32",x"4C", -- 0x0228
    x"32",x"34",x"4C",x"3A",x"04",x"4C",x"32",x"31", -- 0x0230
    x"4C",x"3A",x"05",x"4C",x"32",x"32",x"4C",x"ED", -- 0x0238
    x"5B",x"1D",x"4C",x"7A",x"C6",x"10",x"57",x"CD", -- 0x0240
    x"4B",x"0C",x"20",x"0E",x"ED",x"5B",x"1D",x"4C", -- 0x0248
    x"1C",x"7A",x"C6",x"10",x"57",x"CD",x"4B",x"0C", -- 0x0250
    x"28",x"41",x"3A",x"2C",x"4C",x"FE",x"00",x"28", -- 0x0258
    x"1E",x"3A",x"1F",x"4C",x"E6",x"02",x"28",x"08", -- 0x0260
    x"3A",x"31",x"4C",x"2F",x"E6",x"02",x"20",x"0D", -- 0x0268
    x"3A",x"31",x"4C",x"E6",x"FB",x"F6",x"02",x"32", -- 0x0270
    x"31",x"4C",x"32",x"26",x"4C",x"18",x"1C",x"3A", -- 0x0278
    x"1F",x"4C",x"E6",x"02",x"20",x"08",x"3A",x"31", -- 0x0280
    x"4C",x"2F",x"E6",x"04",x"20",x"0D",x"3A",x"31", -- 0x0288
    x"4C",x"E6",x"FD",x"F6",x"04",x"32",x"31",x"4C", -- 0x0290
    x"32",x"26",x"4C",x"3A",x"24",x"4C",x"B7",x"28", -- 0x0298
    x"06",x"3A",x"25",x"4C",x"32",x"31",x"4C",x"3A", -- 0x02A0
    x"31",x"4C",x"CB",x"4F",x"20",x"6F",x"F6",x"04", -- 0x02A8
    x"32",x"31",x"4C",x"32",x"26",x"4C",x"32",x"25", -- 0x02B0
    x"4C",x"3A",x"1F",x"4C",x"CB",x"4F",x"20",x"10", -- 0x02B8
    x"3A",x"31",x"4C",x"F6",x"02",x"32",x"31",x"4C", -- 0x02C0
    x"32",x"26",x"4C",x"32",x"25",x"4C",x"18",x"45", -- 0x02C8
    x"D6",x"04",x"E6",x"0F",x"32",x"1F",x"4C",x"FE", -- 0x02D0
    x"0E",x"20",x"3A",x"ED",x"5B",x"1D",x"4C",x"1D", -- 0x02D8
    x"CD",x"3A",x"0C",x"20",x"2B",x"ED",x"5B",x"1D", -- 0x02E0
    x"4C",x"1D",x"7A",x"C6",x"08",x"57",x"CD",x"3A", -- 0x02E8
    x"0C",x"20",x"1D",x"ED",x"5B",x"1D",x"4C",x"1D", -- 0x02F0
    x"7A",x"C6",x"0F",x"57",x"CD",x"3A",x"0C",x"20", -- 0x02F8
    x"0F",x"3A",x"1D",x"4C",x"3D",x"32",x"1D",x"4C", -- 0x0300
    x"FE",x"FF",x"20",x"11",x"3C",x"32",x"1D",x"4C", -- 0x0308
    x"3E",x"02",x"32",x"1F",x"4C",x"3A",x"1F",x"4C", -- 0x0310
    x"F6",x"02",x"32",x"1F",x"4C",x"3A",x"31",x"4C", -- 0x0318
    x"CB",x"57",x"20",x"70",x"F6",x"02",x"32",x"31", -- 0x0320
    x"4C",x"32",x"26",x"4C",x"32",x"25",x"4C",x"3A", -- 0x0328
    x"1F",x"4C",x"CB",x"4F",x"28",x"10",x"3A",x"31", -- 0x0330
    x"4C",x"F6",x"04",x"32",x"31",x"4C",x"32",x"26", -- 0x0338
    x"4C",x"32",x"25",x"4C",x"18",x"46",x"C6",x"04", -- 0x0340
    x"E6",x"0F",x"32",x"1F",x"4C",x"20",x"3D",x"ED", -- 0x0348
    x"5B",x"1D",x"4C",x"1C",x"1C",x"CD",x"3A",x"0C", -- 0x0350
    x"20",x"2D",x"ED",x"5B",x"1D",x"4C",x"1C",x"1C", -- 0x0358
    x"7A",x"C6",x"08",x"57",x"CD",x"3A",x"0C",x"20", -- 0x0360
    x"1E",x"ED",x"5B",x"1D",x"4C",x"1C",x"1C",x"7A", -- 0x0368
    x"C6",x"0F",x"57",x"CD",x"3A",x"0C",x"20",x"0F", -- 0x0370
    x"3A",x"1D",x"4C",x"3C",x"FE",x"1B",x"32",x"1D", -- 0x0378
    x"4C",x"20",x"11",x"3D",x"32",x"1D",x"4C",x"3E", -- 0x0380
    x"0C",x"32",x"1F",x"4C",x"3A",x"1F",x"4C",x"E6", -- 0x0388
    x"FD",x"32",x"1F",x"4C",x"3A",x"32",x"4C",x"CB", -- 0x0390
    x"57",x"20",x"25",x"3A",x"24",x"4C",x"B7",x"20", -- 0x0398
    x"1F",x"AF",x"32",x"23",x"4C",x"3E",x"01",x"32", -- 0x03A0
    x"24",x"4C",x"3E",x"FC",x"32",x"22",x"4C",x"3A", -- 0x03A8
    x"1E",x"4C",x"32",x"28",x"4C",x"3A",x"31",x"4C", -- 0x03B0
    x"32",x"25",x"4C",x"3E",x"01",x"32",x"2A",x"4C", -- 0x03B8
    x"3A",x"24",x"4C",x"B7",x"CA",x"BB",x"04",x"3C", -- 0x03C0
    x"32",x"24",x"4C",x"ED",x"5B",x"22",x"4C",x"3A", -- 0x03C8
    x"1E",x"4C",x"83",x"32",x"1E",x"4C",x"3A",x"24", -- 0x03D0
    x"4C",x"E6",x"01",x"28",x"0D",x"7B",x"CB",x"7F", -- 0x03D8
    x"20",x"04",x"FE",x"04",x"30",x"04",x"3C",x"32", -- 0x03E0
    x"22",x"4C",x"3A",x"22",x"4C",x"CB",x"7F",x"C2", -- 0x03E8
    x"53",x"04",x"FE",x"03",x"38",x"5D",x"ED",x"5B", -- 0x03F0
    x"1D",x"4C",x"7A",x"C6",x"10",x"57",x"CD",x"1B", -- 0x03F8
    x"0C",x"28",x"20",x"AF",x"32",x"22",x"4C",x"32", -- 0x0400
    x"24",x"4C",x"3A",x"1E",x"4C",x"E6",x"F8",x"32", -- 0x0408
    x"1E",x"4C",x"3A",x"28",x"4C",x"C6",x"18",x"5F", -- 0x0410
    x"3A",x"1E",x"4C",x"BB",x"38",x"05",x"3E",x"02", -- 0x0418
    x"32",x"2B",x"4C",x"ED",x"5B",x"1D",x"4C",x"1C", -- 0x0420
    x"7A",x"C6",x"10",x"57",x"CD",x"1B",x"0C",x"28", -- 0x0428
    x"20",x"AF",x"32",x"22",x"4C",x"32",x"24",x"4C", -- 0x0430
    x"3A",x"1E",x"4C",x"E6",x"F8",x"32",x"1E",x"4C", -- 0x0438
    x"3A",x"28",x"4C",x"C6",x"18",x"5F",x"3A",x"1E", -- 0x0440
    x"4C",x"BB",x"38",x"05",x"3E",x"02",x"32",x"2B", -- 0x0448
    x"4C",x"18",x"56",x"ED",x"5B",x"1D",x"4C",x"15", -- 0x0450
    x"CD",x"3A",x"0C",x"20",x"0B",x"ED",x"5B",x"1D", -- 0x0458
    x"4C",x"1C",x"15",x"CD",x"3A",x"0C",x"28",x"41", -- 0x0460
    x"3A",x"22",x"4C",x"CB",x"7F",x"28",x"3A",x"AF", -- 0x0468
    x"32",x"22",x"4C",x"3E",x"FF",x"32",x"25",x"4C", -- 0x0470
    x"32",x"26",x"4C",x"3A",x"1E",x"4C",x"3D",x"E6", -- 0x0478
    x"78",x"C6",x"08",x"32",x"1E",x"4C",x"ED",x"5B", -- 0x0480
    x"1D",x"4C",x"7A",x"C6",x"10",x"57",x"D5",x"CD", -- 0x0488
    x"1B",x"0C",x"D1",x"20",x"06",x"1C",x"CD",x"1B", -- 0x0490
    x"0C",x"28",x"0E",x"AF",x"32",x"24",x"4C",x"32", -- 0x0498
    x"22",x"4C",x"3E",x"FF",x"32",x"25",x"4C",x"18", -- 0x04A0
    x"43",x"3A",x"23",x"4C",x"3C",x"32",x"23",x"4C", -- 0x04A8
    x"FE",x"11",x"38",x"38",x"3E",x"FF",x"32",x"25", -- 0x04B0
    x"4C",x"18",x"31",x"3A",x"24",x"4C",x"B7",x"20", -- 0x04B8
    x"2B",x"ED",x"5B",x"1D",x"4C",x"7A",x"C6",x"10", -- 0x04C0
    x"57",x"D5",x"CD",x"1B",x"0C",x"D1",x"20",x"1C", -- 0x04C8
    x"1C",x"CD",x"1B",x"0C",x"20",x"16",x"AF",x"32", -- 0x04D0
    x"22",x"4C",x"3E",x"FF",x"32",x"25",x"4C",x"3E", -- 0x04D8
    x"01",x"32",x"24",x"4C",x"3A",x"1E",x"4C",x"C6", -- 0x04E0
    x"10",x"32",x"28",x"4C",x"ED",x"5B",x"1D",x"4C", -- 0x04E8
    x"CB",x"23",x"CB",x"23",x"CB",x"23",x"ED",x"4B", -- 0x04F0
    x"1F",x"4C",x"D5",x"79",x"E6",x"0C",x"1F",x"D1", -- 0x04F8
    x"83",x"32",x"29",x"4C",x"ED",x"5B",x"1D",x"4C", -- 0x0500
    x"CB",x"23",x"CB",x"23",x"CB",x"23",x"ED",x"4B", -- 0x0508
    x"1F",x"4C",x"CB",x"49",x"28",x"04",x"79",x"EE", -- 0x0510
    x"0C",x"4F",x"3E",x"00",x"CD",x"D5",x"0B",x"DD", -- 0x0518
    x"21",x"71",x"4C",x"06",x"01",x"3A",x"41",x"4C", -- 0x0520
    x"B7",x"28",x"21",x"4F",x"C5",x"DD",x"5E",x"01", -- 0x0528
    x"CB",x"23",x"CB",x"23",x"CB",x"23",x"DD",x"56", -- 0x0530
    x"02",x"DD",x"4E",x"00",x"78",x"06",x"01",x"CD", -- 0x0538
    x"D5",x"0B",x"C1",x"11",x"07",x"00",x"DD",x"19", -- 0x0540
    x"04",x"0D",x"20",x"E0",x"DD",x"21",x"8D",x"4C", -- 0x0548
    x"3A",x"42",x"4C",x"B7",x"28",x"21",x"4F",x"C5", -- 0x0550
    x"DD",x"5E",x"01",x"CB",x"23",x"CB",x"23",x"CB", -- 0x0558
    x"23",x"DD",x"56",x"02",x"DD",x"4E",x"00",x"78", -- 0x0560
    x"06",x"01",x"CD",x"D5",x"0B",x"C1",x"11",x"07", -- 0x0568
    x"00",x"DD",x"19",x"04",x"0D",x"20",x"E0",x"78", -- 0x0570
    x"FE",x"08",x"28",x"0C",x"11",x"F0",x"F0",x"DD", -- 0x0578
    x"4E",x"00",x"CD",x"D5",x"0B",x"04",x"18",x"EF", -- 0x0580
    x"3E",x"01",x"32",x"50",x"4C",x"3A",x"24",x"4C", -- 0x0588
    x"B7",x"20",x"43",x"ED",x"5B",x"1D",x"4C",x"7A", -- 0x0590
    x"C6",x"10",x"57",x"CD",x"0F",x"0C",x"FE",x"68", -- 0x0598
    x"38",x"12",x"FE",x"A0",x"30",x"0E",x"3C",x"77", -- 0x05A0
    x"E6",x"07",x"20",x"08",x"36",x"03",x"CB",x"D4", -- 0x05A8
    x"3A",x"36",x"4C",x"77",x"ED",x"5B",x"1D",x"4C", -- 0x05B0
    x"1C",x"7A",x"C6",x"10",x"57",x"CD",x"0F",x"0C", -- 0x05B8
    x"FE",x"68",x"38",x"12",x"FE",x"A0",x"30",x"0E", -- 0x05C0
    x"3C",x"77",x"E6",x"07",x"20",x"08",x"36",x"03", -- 0x05C8
    x"CB",x"D4",x"3A",x"36",x"4C",x"77",x"ED",x"5B", -- 0x05D0
    x"1D",x"4C",x"CD",x"7A",x"0A",x"1C",x"CD",x"7A", -- 0x05D8
    x"0A",x"7A",x"C6",x"08",x"57",x"CD",x"7A",x"0A", -- 0x05E0
    x"1D",x"CD",x"7A",x"0A",x"7A",x"C6",x"07",x"57", -- 0x05E8
    x"CD",x"7A",x"0A",x"1C",x"CD",x"7A",x"0A",x"DD", -- 0x05F0
    x"21",x"71",x"4C",x"3A",x"41",x"4C",x"B7",x"28", -- 0x05F8
    x"61",x"47",x"DD",x"7E",x"03",x"DD",x"86",x"06", -- 0x0600
    x"DD",x"77",x"03",x"1F",x"1F",x"1F",x"DD",x"77", -- 0x0608
    x"01",x"DD",x"7E",x"03",x"DD",x"BE",x"04",x"38", -- 0x0610
    x"05",x"DD",x"BE",x"05",x"38",x"08",x"DD",x"7E", -- 0x0618
    x"06",x"2F",x"3C",x"DD",x"77",x"06",x"DD",x"7E", -- 0x0620
    x"03",x"E6",x"06",x"87",x"4F",x"DD",x"7E",x"00", -- 0x0628
    x"E6",x"F0",x"B1",x"DD",x"77",x"00",x"DD",x"CB", -- 0x0630
    x"06",x"7E",x"28",x"08",x"DD",x"7E",x"00",x"EE", -- 0x0638
    x"0E",x"DD",x"77",x"00",x"DD",x"5E",x"03",x"DD", -- 0x0640
    x"56",x"02",x"2A",x"1D",x"4C",x"3A",x"29",x"4C", -- 0x0648
    x"6F",x"CD",x"FA",x"09",x"38",x"05",x"3E",x"02", -- 0x0650
    x"32",x"2B",x"4C",x"11",x"07",x"00",x"DD",x"19", -- 0x0658
    x"10",x"A0",x"DD",x"21",x"8D",x"4C",x"3A",x"42", -- 0x0660
    x"4C",x"B7",x"CA",x"2C",x"07",x"47",x"DD",x"7E", -- 0x0668
    x"06",x"B7",x"28",x"11",x"3A",x"2F",x"4C",x"FE", -- 0x0670
    x"07",x"28",x"04",x"FE",x"0B",x"20",x"06",x"11", -- 0x0678
    x"0E",x"0A",x"CD",x"26",x"0A",x"DD",x"7E",x"02", -- 0x0680
    x"DD",x"86",x"06",x"DD",x"77",x"02",x"DD",x"BE", -- 0x0688
    x"04",x"38",x"05",x"DD",x"BE",x"05",x"38",x"4A", -- 0x0690
    x"DD",x"7E",x"06",x"2F",x"3C",x"DD",x"77",x"06", -- 0x0698
    x"3A",x"2F",x"4C",x"FE",x"07",x"28",x"37",x"FE", -- 0x06A0
    x"0B",x"28",x"33",x"FE",x"0D",x"28",x"13",x"FE", -- 0x06A8
    x"04",x"28",x"02",x"18",x"2D",x"3A",x"3C",x"4C", -- 0x06B0
    x"B7",x"20",x"27",x"3E",x"00",x"DD",x"77",x"06", -- 0x06B8
    x"18",x"20",x"DD",x"7E",x"03",x"C6",x"40",x"DD", -- 0x06C0
    x"77",x"03",x"1F",x"1F",x"1F",x"DD",x"77",x"01", -- 0x06C8
    x"AF",x"DD",x"77",x"02",x"DD",x"7E",x"06",x"2F", -- 0x06D0
    x"3C",x"DD",x"77",x"06",x"18",x"04",x"AF",x"32", -- 0x06D8
    x"42",x"4C",x"3A",x"30",x"4C",x"E6",x"03",x"20", -- 0x06E0
    x"23",x"DD",x"7E",x"00",x"FE",x"20",x"38",x"1C", -- 0x06E8
    x"FE",x"A0",x"38",x"13",x"C6",x"04",x"DD",x"77", -- 0x06F0
    x"00",x"E6",x"0C",x"FE",x"00",x"20",x"0D",x"DD", -- 0x06F8
    x"7E",x"00",x"D6",x"10",x"DD",x"77",x"00",x"EE", -- 0x0700
    x"04",x"DD",x"77",x"00",x"DD",x"5E",x"03",x"DD", -- 0x0708
    x"56",x"02",x"2A",x"1D",x"4C",x"3A",x"29",x"4C", -- 0x0710
    x"6F",x"CD",x"FA",x"09",x"38",x"05",x"3E",x"02", -- 0x0718
    x"32",x"2B",x"4C",x"11",x"07",x"00",x"DD",x"19", -- 0x0720
    x"05",x"C2",x"6E",x"06",x"3A",x"07",x"4C",x"E6", -- 0x0728
    x"20",x"28",x"0A",x"3A",x"05",x"4C",x"E6",x"60", -- 0x0730
    x"20",x"03",x"C3",x"58",x"01",x"3A",x"2B",x"4C", -- 0x0738
    x"B7",x"CA",x"ED",x"01",x"FE",x"01",x"28",x"1C", -- 0x0740
    x"3E",x"40",x"32",x"4E",x"4C",x"3A",x"27",x"4C", -- 0x0748
    x"3D",x"32",x"27",x"4C",x"C2",x"E0",x"01",x"AF", -- 0x0750
    x"32",x"47",x"4C",x"32",x"24",x"4C",x"CD",x"19", -- 0x0758
    x"09",x"C3",x"58",x"01",x"AF",x"32",x"24",x"4C", -- 0x0760
    x"3A",x"39",x"4C",x"B7",x"28",x"11",x"32",x"4A", -- 0x0768
    x"4C",x"CD",x"83",x"0B",x"CD",x"3C",x"0B",x"11", -- 0x0770
    x"14",x"0A",x"CD",x"26",x"0A",x"18",x"E5",x"3A", -- 0x0778
    x"2F",x"4C",x"3C",x"32",x"2F",x"4C",x"FE",x"14", -- 0x0780
    x"DA",x"E0",x"01",x"AF",x"32",x"2F",x"4C",x"C3", -- 0x0788
    x"E0",x"01",x"3A",x"2F",x"4C",x"FE",x"12",x"C0", -- 0x0790
    x"11",x"14",x"00",x"CD",x"6D",x"0B",x"CB",x"D4", -- 0x0798
    x"11",x"14",x"00",x"7E",x"FE",x"18",x"20",x"34", -- 0x07A0
    x"7E",x"FE",x"18",x"20",x"24",x"36",x"0F",x"2C", -- 0x07A8
    x"14",x"18",x"F5",x"01",x"E1",x"FF",x"09",x"15", -- 0x07B0
    x"1D",x"7E",x"FE",x"18",x"28",x"EA",x"18",x"1C", -- 0x07B8
    x"7E",x"FE",x"18",x"20",x"EE",x"36",x"0F",x"01", -- 0x07C0
    x"20",x"00",x"09",x"1D",x"FA",x"DC",x"07",x"18", -- 0x07C8
    x"EF",x"01",x"1F",x"00",x"09",x"15",x"1D",x"7E", -- 0x07D0
    x"FE",x"18",x"28",x"E9",x"21",x"A4",x"47",x"36", -- 0x07D8
    x"0F",x"2E",x"84",x"36",x"0F",x"DD",x"21",x"71", -- 0x07E0
    x"4C",x"3A",x"41",x"4C",x"B7",x"28",x"31",x"47", -- 0x07E8
    x"DD",x"5E",x"03",x"DD",x"56",x"02",x"CB",x"3B", -- 0x07F0
    x"CB",x"3B",x"CB",x"3B",x"CB",x"3A",x"CB",x"3A", -- 0x07F8
    x"CB",x"3A",x"CD",x"6D",x"0B",x"CB",x"D4",x"CD", -- 0x0800
    x"0B",x"09",x"2C",x"CD",x"0B",x"09",x"11",x"E0", -- 0x0808
    x"FF",x"19",x"CD",x"0B",x"09",x"2D",x"CD",x"0B", -- 0x0810
    x"09",x"11",x"07",x"00",x"DD",x"19",x"10",x"D0", -- 0x0818
    x"DD",x"21",x"8D",x"4C",x"3A",x"42",x"4C",x"B7", -- 0x0820
    x"CA",x"5E",x"08",x"47",x"DD",x"5E",x"03",x"DD", -- 0x0828
    x"56",x"02",x"CB",x"3B",x"CB",x"3B",x"CB",x"3B", -- 0x0830
    x"CB",x"3A",x"CB",x"3A",x"CB",x"3A",x"CD",x"6D", -- 0x0838
    x"0B",x"CB",x"D4",x"CD",x"0B",x"09",x"2C",x"CD", -- 0x0840
    x"0B",x"09",x"11",x"E0",x"FF",x"19",x"CD",x"0B", -- 0x0848
    x"09",x"2D",x"CD",x"0B",x"09",x"11",x"07",x"00", -- 0x0850
    x"DD",x"19",x"05",x"C2",x"2C",x"08",x"3A",x"2F", -- 0x0858
    x"4C",x"FE",x"12",x"C0",x"11",x"14",x"00",x"CD", -- 0x0860
    x"6D",x"0B",x"CB",x"D4",x"11",x"14",x"00",x"01", -- 0x0868
    x"20",x"00",x"7E",x"FE",x"16",x"28",x"13",x"FE", -- 0x0870
    x"0F",x"20",x"16",x"36",x"18",x"2C",x"14",x"18", -- 0x0878
    x"F1",x"7E",x"FE",x"16",x"28",x"F5",x"FE",x"0F", -- 0x0880
    x"20",x"07",x"36",x"18",x"09",x"1D",x"F2",x"81", -- 0x0888
    x"08",x"DD",x"21",x"71",x"4C",x"3A",x"41",x"4C", -- 0x0890
    x"B7",x"28",x"31",x"47",x"DD",x"5E",x"03",x"DD", -- 0x0898
    x"56",x"02",x"CB",x"3B",x"CB",x"3B",x"CB",x"3B", -- 0x08A0
    x"CB",x"3A",x"CB",x"3A",x"CB",x"3A",x"CD",x"6D", -- 0x08A8
    x"0B",x"CB",x"D4",x"CD",x"12",x"09",x"2C",x"CD", -- 0x08B0
    x"12",x"09",x"11",x"E0",x"FF",x"19",x"CD",x"12", -- 0x08B8
    x"09",x"2D",x"CD",x"12",x"09",x"11",x"07",x"00", -- 0x08C0
    x"DD",x"19",x"10",x"D0",x"DD",x"21",x"8D",x"4C", -- 0x08C8
    x"3A",x"42",x"4C",x"B7",x"CA",x"0A",x"09",x"47", -- 0x08D0
    x"DD",x"5E",x"03",x"DD",x"56",x"02",x"CB",x"3B", -- 0x08D8
    x"CB",x"3B",x"CB",x"3B",x"CB",x"3A",x"CB",x"3A", -- 0x08E0
    x"CB",x"3A",x"CD",x"6D",x"0B",x"CB",x"D4",x"CD", -- 0x08E8
    x"12",x"09",x"2C",x"CD",x"12",x"09",x"11",x"E0", -- 0x08F0
    x"FF",x"19",x"CD",x"12",x"09",x"2D",x"CD",x"12", -- 0x08F8
    x"09",x"11",x"07",x"00",x"DD",x"19",x"05",x"C2", -- 0x0900
    x"D8",x"08",x"C9",x"7E",x"FE",x"0F",x"C0",x"36", -- 0x0908
    x"16",x"C9",x"7E",x"FE",x"18",x"C8",x"36",x"0F", -- 0x0910
    x"C9",x"AF",x"32",x"50",x"4C",x"CD",x"83",x"0B", -- 0x0918
    x"11",x"00",x"00",x"06",x"1C",x"D5",x"C5",x"CD", -- 0x0920
    x"6D",x"0B",x"06",x"10",x"AF",x"36",x"03",x"CB", -- 0x0928
    x"D4",x"77",x"CB",x"94",x"2C",x"10",x"F6",x"C1", -- 0x0930
    x"D1",x"1C",x"10",x"E9",x"CD",x"CB",x"0E",x"3E", -- 0x0938
    x"60",x"32",x"1E",x"4C",x"CD",x"83",x"0B",x"ED", -- 0x0940
    x"5F",x"11",x"00",x"00",x"06",x"1C",x"D5",x"C5", -- 0x0948
    x"F5",x"CD",x"6D",x"0B",x"F1",x"06",x"10",x"CB", -- 0x0950
    x"D4",x"77",x"2C",x"10",x"FA",x"C1",x"D1",x"1C", -- 0x0958
    x"10",x"EC",x"21",x"20",x"46",x"3A",x"1E",x"4C", -- 0x0960
    x"47",x"3E",x"60",x"90",x"1F",x"1F",x"1F",x"E6", -- 0x0968
    x"1F",x"3C",x"47",x"3E",x"01",x"77",x"2C",x"10", -- 0x0970
    x"FC",x"ED",x"4B",x"1E",x"4C",x"3E",x"61",x"91", -- 0x0978
    x"1F",x"1F",x"1F",x"E6",x"1F",x"57",x"1E",x"0C", -- 0x0980
    x"CD",x"6D",x"0B",x"36",x"17",x"CB",x"D4",x"36", -- 0x0988
    x"01",x"11",x"5D",x"70",x"01",x"14",x"01",x"3E", -- 0x0990
    x"02",x"CD",x"D5",x"0B",x"11",x"60",x"60",x"01", -- 0x0998
    x"00",x"01",x"3E",x"01",x"CD",x"D5",x"0B",x"11", -- 0x09A0
    x"5E",x"00",x"ED",x"4B",x"1E",x"4C",x"3E",x"61", -- 0x09A8
    x"91",x"57",x"01",x"18",x"01",x"3E",x"00",x"CD", -- 0x09B0
    x"D5",x"0B",x"3A",x"1E",x"4C",x"3D",x"32",x"1E", -- 0x09B8
    x"4C",x"F5",x"CB",x"3F",x"CB",x"3F",x"32",x"4A", -- 0x09C0
    x"4C",x"F1",x"C2",x"44",x"09",x"11",x"00",x"00", -- 0x09C8
    x"06",x"1C",x"AF",x"D5",x"C5",x"F5",x"CD",x"6D", -- 0x09D0
    x"0B",x"F1",x"06",x"10",x"CB",x"D4",x"77",x"2C", -- 0x09D8
    x"10",x"FA",x"C1",x"D1",x"1C",x"10",x"EC",x"21", -- 0x09E0
    x"20",x"46",x"06",x"0C",x"3E",x"01",x"77",x"2C", -- 0x09E8
    x"10",x"FC",x"06",x"FA",x"CD",x"83",x"0B",x"10", -- 0x09F0
    x"FB",x"C9",x"7D",x"C6",x"06",x"BB",x"D8",x"7B", -- 0x09F8
    x"C6",x"06",x"BD",x"D8",x"7C",x"C6",x"0F",x"BA", -- 0x0A00
    x"D8",x"7A",x"C6",x"0F",x"BC",x"C9",x"00",x"00", -- 0x0A08
    x"01",x"00",x"00",x"00",x"08",x"00",x"00",x"00", -- 0x0A10
    x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00", -- 0x0A18
    x"00",x"05",x"02",x"00",x"00",x"00",x"E5",x"C5", -- 0x0A20
    x"21",x"12",x"4C",x"01",x"00",x"06",x"1A",x"86", -- 0x0A28
    x"81",x"77",x"0E",x"00",x"FE",x"3A",x"38",x"04", -- 0x0A30
    x"D6",x"0A",x"77",x"0C",x"2B",x"13",x"10",x"EE", -- 0x0A38
    x"21",x"0D",x"4C",x"11",x"14",x"4C",x"06",x"06", -- 0x0A40
    x"1A",x"BE",x"28",x"0E",x"30",x"10",x"21",x"0D", -- 0x0A48
    x"4C",x"11",x"14",x"4C",x"01",x"06",x"00",x"EF", -- 0x0A50
    x"18",x"04",x"23",x"13",x"10",x"EA",x"CD",x"AE", -- 0x0A58
    x"0E",x"C1",x"E1",x"C9",x"CD",x"83",x"0B",x"3A", -- 0x0A60
    x"40",x"50",x"E6",x"20",x"20",x"F6",x"C9",x"CD", -- 0x0A68
    x"83",x"0B",x"3A",x"40",x"50",x"E6",x"20",x"28", -- 0x0A70
    x"F6",x"C9",x"D5",x"CD",x"0F",x"0C",x"D1",x"FE", -- 0x0A78
    x"18",x"D8",x"FE",x"20",x"DA",x"10",x"0B",x"FE", -- 0x0A80
    x"30",x"D8",x"FE",x"40",x"DA",x"10",x"0B",x"FE", -- 0x0A88
    x"FE",x"D2",x"16",x"0B",x"FE",x"DE",x"38",x"05", -- 0x0A90
    x"FE",x"E0",x"DA",x"16",x"0B",x"FE",x"44",x"28", -- 0x0A98
    x"42",x"FE",x"45",x"28",x"3E",x"FE",x"46",x"C0", -- 0x0AA0
    x"36",x"47",x"7B",x"FE",x"11",x"38",x"23",x"3A", -- 0x0AA8
    x"8D",x"4C",x"C6",x"08",x"32",x"8D",x"4C",x"3E", -- 0x0AB0
    x"04",x"32",x"93",x"4C",x"E5",x"D5",x"21",x"E2", -- 0x0AB8
    x"41",x"AF",x"77",x"11",x"E0",x"FF",x"19",x"77", -- 0x0AC0
    x"CB",x"D4",x"77",x"AF",x"ED",x"52",x"77",x"D1", -- 0x0AC8
    x"E1",x"C9",x"E5",x"D5",x"21",x"AB",x"41",x"AF", -- 0x0AD0
    x"77",x"2C",x"77",x"CB",x"D4",x"77",x"2D",x"77", -- 0x0AD8
    x"D1",x"E1",x"C9",x"36",x"03",x"CB",x"D4",x"3A", -- 0x0AE0
    x"36",x"4C",x"77",x"3A",x"3C",x"4C",x"3D",x"32", -- 0x0AE8
    x"3C",x"4C",x"D5",x"11",x"1A",x"0A",x"CD",x"26", -- 0x0AF0
    x"0A",x"D1",x"3E",x"02",x"32",x"4F",x"4C",x"3A", -- 0x0AF8
    x"2F",x"4C",x"FE",x"04",x"C0",x"3A",x"3C",x"4C", -- 0x0B00
    x"B7",x"C0",x"3E",x"01",x"32",x"93",x"4C",x"C9", -- 0x0B08
    x"3E",x"02",x"32",x"2B",x"4C",x"C9",x"3A",x"3C", -- 0x0B10
    x"4C",x"B7",x"C0",x"D5",x"3A",x"29",x"4C",x"C6", -- 0x0B18
    x"05",x"1F",x"1F",x"1F",x"E6",x"1F",x"5F",x"3A", -- 0x0B20
    x"1E",x"4C",x"C6",x"08",x"57",x"CD",x"0F",x"0C", -- 0x0B28
    x"D1",x"E6",x"DE",x"FE",x"DE",x"C0",x"3E",x"01", -- 0x0B30
    x"32",x"2B",x"4C",x"C9",x"3A",x"39",x"4C",x"B7", -- 0x0B38
    x"28",x"25",x"3D",x"32",x"39",x"4C",x"1F",x"1F", -- 0x0B40
    x"1F",x"E6",x"1F",x"C6",x"04",x"5F",x"16",x"11", -- 0x0B48
    x"CD",x"6D",x"0B",x"3A",x"39",x"4C",x"E6",x"07", -- 0x0B50
    x"C6",x"60",x"77",x"E6",x"07",x"FE",x"07",x"C0", -- 0x0B58
    x"11",x"E0",x"FF",x"19",x"36",x"A0",x"C9",x"21", -- 0x0B60
    x"31",x"43",x"36",x"A0",x"C9",x"7A",x"C6",x"A0", -- 0x0B68
    x"6F",x"26",x"43",x"7B",x"11",x"E0",x"FF",x"B7", -- 0x0B70
    x"C8",x"1F",x"30",x"01",x"19",x"EB",x"29",x"EB", -- 0x0B78
    x"C3",x"77",x"0B",x"E5",x"2A",x"00",x"4C",x"AF", -- 0x0B80
    x"32",x"C0",x"50",x"3A",x"00",x"4C",x"BD",x"28", -- 0x0B88
    x"F6",x"E1",x"C9",x"7E",x"23",x"B7",x"C8",x"C6", -- 0x0B90
    x"80",x"12",x"CB",x"D2",x"79",x"12",x"7B",x"D6", -- 0x0B98
    x"20",x"5F",x"CB",x"92",x"7A",x"DE",x"00",x"57", -- 0x0BA0
    x"C3",x"93",x"0B",x"7C",x"CD",x"B0",x"0B",x"7D", -- 0x0BA8
    x"F5",x"1F",x"1F",x"1F",x"1F",x"CD",x"B9",x"0B", -- 0x0BB0
    x"F1",x"E6",x"0F",x"FE",x"0A",x"38",x"02",x"C6", -- 0x0BB8
    x"07",x"C6",x"B0",x"E5",x"D5",x"F5",x"CD",x"6D", -- 0x0BC0
    x"0B",x"F1",x"77",x"CB",x"D4",x"36",x"12",x"CB", -- 0x0BC8
    x"94",x"D1",x"1C",x"E1",x"C9",x"F5",x"3E",x"F0", -- 0x0BD0
    x"BA",x"20",x"03",x"BB",x"28",x"2C",x"F1",x"3C", -- 0x0BD8
    x"D5",x"ED",x"5B",x"1C",x"4C",x"BB",x"38",x"03", -- 0x0BE0
    x"32",x"1C",x"4C",x"E6",x"07",x"87",x"5F",x"16", -- 0x0BE8
    x"00",x"21",x"51",x"4C",x"19",x"D1",x"71",x"23", -- 0x0BF0
    x"70",x"23",x"D5",x"11",x"0E",x"00",x"19",x"D1", -- 0x0BF8
    x"3E",x"EE",x"93",x"77",x"23",x"3E",x"00",x"92", -- 0x0C00
    x"77",x"C9",x"F1",x"3C",x"D5",x"18",x"DC",x"7A", -- 0x0C08
    x"1F",x"1F",x"1F",x"E6",x"1F",x"57",x"CD",x"6D", -- 0x0C10
    x"0B",x"7E",x"C9",x"CD",x"0F",x"0C",x"FE",x"05", -- 0x0C18
    x"38",x"14",x"FE",x"18",x"38",x"12",x"FE",x"20", -- 0x0C20
    x"38",x"0C",x"FE",x"30",x"38",x"0A",x"FE",x"48", -- 0x0C28
    x"38",x"04",x"FE",x"A0",x"38",x"02",x"AF",x"C9", -- 0x0C30
    x"B7",x"C9",x"CD",x"0F",x"0C",x"FE",x"20",x"38", -- 0x0C38
    x"04",x"FE",x"30",x"38",x"02",x"AF",x"C9",x"3E", -- 0x0C40
    x"01",x"B7",x"C9",x"CD",x"0F",x"0C",x"FE",x"48", -- 0x0C48
    x"38",x"04",x"FE",x"60",x"38",x"02",x"AF",x"C9", -- 0x0C50
    x"3E",x"01",x"B7",x"C9",x"32",x"36",x"4C",x"F5", -- 0x0C58
    x"AF",x"32",x"50",x"4C",x"CD",x"83",x"0B",x"F1", -- 0x0C60
    x"F3",x"E5",x"D5",x"C5",x"F5",x"21",x"00",x"40", -- 0x0C68
    x"11",x"01",x"40",x"01",x"00",x"04",x"36",x"03", -- 0x0C70
    x"ED",x"B0",x"01",x"40",x"00",x"36",x"00",x"ED", -- 0x0C78
    x"B0",x"01",x"80",x"03",x"77",x"ED",x"B0",x"36", -- 0x0C80
    x"00",x"01",x"3F",x"00",x"ED",x"B0",x"FB",x"CD", -- 0x0C88
    x"83",x"0B",x"F3",x"11",x"00",x"10",x"06",x"10", -- 0x0C90
    x"D5",x"C5",x"CD",x"6D",x"0B",x"11",x"E0",x"FF", -- 0x0C98
    x"CB",x"D4",x"06",x"20",x"36",x"00",x"19",x"10", -- 0x0CA0
    x"FB",x"C1",x"D1",x"14",x"10",x"EA",x"CD",x"69", -- 0x0CA8
    x"12",x"F1",x"C1",x"D1",x"E1",x"FB",x"C9",x"3A", -- 0x0CB0
    x"3C",x"4C",x"B7",x"C0",x"ED",x"5F",x"21",x"D8", -- 0x0CB8
    x"0C",x"E6",x"03",x"5F",x"16",x"00",x"19",x"7E", -- 0x0CC0
    x"2A",x"3F",x"4C",x"CB",x"D4",x"77",x"2C",x"77", -- 0x0CC8
    x"11",x"E0",x"FF",x"19",x"77",x"2D",x"77",x"C9", -- 0x0CD0
    x"09",x"11",x"14",x"17",x"C9",x"DD",x"2A",x"37", -- 0x0CD8
    x"4C",x"DD",x"7E",x"02",x"B7",x"C8",x"47",x"DD", -- 0x0CE0
    x"5E",x"00",x"DD",x"56",x"01",x"CD",x"6D",x"0B", -- 0x0CE8
    x"DD",x"7E",x"05",x"32",x"2C",x"4C",x"FE",x"00", -- 0x0CF0
    x"3A",x"30",x"4C",x"28",x"01",x"2F",x"E6",x"07", -- 0x0CF8
    x"DD",x"86",x"03",x"DD",x"4E",x"04",x"C3",x"09", -- 0x0D00
    x"0D",x"11",x"E0",x"FF",x"18",x"03",x"11",x"01", -- 0x0D08
    x"00",x"77",x"CB",x"D4",x"71",x"CB",x"94",x"19", -- 0x0D10
    x"10",x"F7",x"C9",x"6F",x"26",x"00",x"29",x"11", -- 0x0D18
    x"84",x"17",x"19",x"5E",x"23",x"56",x"D5",x"DD", -- 0x0D20
    x"E1",x"DD",x"7E",x"00",x"DD",x"23",x"CD",x"5C", -- 0x0D28
    x"0C",x"DD",x"5E",x"00",x"DD",x"56",x"01",x"CD", -- 0x0D30
    x"6D",x"0B",x"DD",x"7E",x"02",x"B7",x"28",x"1C", -- 0x0D38
    x"47",x"CB",x"B8",x"E6",x"80",x"DD",x"7E",x"03", -- 0x0D40
    x"DD",x"4E",x"04",x"11",x"05",x"00",x"DD",x"19", -- 0x0D48
    x"28",x"05",x"CD",x"0E",x"0D",x"18",x"DA",x"CD", -- 0x0D50
    x"09",x"0D",x"18",x"D5",x"22",x"3F",x"4C",x"36", -- 0x0D58
    x"DE",x"2C",x"36",x"FE",x"CB",x"D4",x"36",x"09", -- 0x0D60
    x"2D",x"36",x"09",x"CB",x"94",x"11",x"E0",x"FF", -- 0x0D68
    x"19",x"36",x"DF",x"2C",x"36",x"FF",x"CB",x"D4", -- 0x0D70
    x"36",x"09",x"2D",x"36",x"09",x"DD",x"7E",x"03", -- 0x0D78
    x"DD",x"4E",x"04",x"DD",x"46",x"05",x"11",x"06", -- 0x0D80
    x"00",x"DD",x"19",x"B7",x"28",x"16",x"F5",x"DD", -- 0x0D88
    x"5E",x"00",x"DD",x"56",x"01",x"DD",x"23",x"DD", -- 0x0D90
    x"23",x"CD",x"6D",x"0B",x"71",x"CB",x"D4",x"70", -- 0x0D98
    x"F1",x"3D",x"20",x"EA",x"DD",x"7E",x"00",x"DD", -- 0x0DA0
    x"4E",x"01",x"DD",x"46",x"02",x"11",x"03",x"00", -- 0x0DA8
    x"DD",x"19",x"B7",x"28",x"16",x"F5",x"DD",x"5E", -- 0x0DB0
    x"00",x"DD",x"56",x"01",x"DD",x"23",x"DD",x"23", -- 0x0DB8
    x"CD",x"6D",x"0B",x"71",x"CB",x"D4",x"70",x"F1", -- 0x0DC0
    x"3D",x"20",x"EA",x"21",x"B0",x"43",x"11",x"E0", -- 0x0DC8
    x"FF",x"06",x"1C",x"36",x"A0",x"CB",x"D4",x"36", -- 0x0DD0
    x"09",x"CB",x"94",x"19",x"10",x"F5",x"DD",x"5E", -- 0x0DD8
    x"00",x"DD",x"23",x"16",x"10",x"CD",x"6D",x"0B", -- 0x0DE0
    x"EB",x"DD",x"E5",x"E1",x"0E",x"09",x"CD",x"93", -- 0x0DE8
    x"0B",x"22",x"37",x"4C",x"11",x"06",x"00",x"19", -- 0x0DF0
    x"7E",x"32",x"1D",x"4C",x"FE",x"10",x"07",x"17", -- 0x0DF8
    x"E6",x"02",x"32",x"1F",x"4C",x"23",x"7E",x"87", -- 0x0E00
    x"87",x"87",x"32",x"1E",x"4C",x"23",x"3E",x"01", -- 0x0E08
    x"32",x"20",x"4C",x"AF",x"32",x"24",x"4C",x"32", -- 0x0E10
    x"22",x"4C",x"3E",x"FF",x"32",x"25",x"4C",x"22", -- 0x0E18
    x"3D",x"4C",x"7E",x"47",x"32",x"3C",x"4C",x"23", -- 0x0E20
    x"7E",x"32",x"3A",x"4C",x"23",x"7E",x"32",x"3B", -- 0x0E28
    x"4C",x"23",x"5E",x"23",x"56",x"23",x"E5",x"CD", -- 0x0E30
    x"6D",x"0B",x"3A",x"3A",x"4C",x"77",x"CB",x"D4", -- 0x0E38
    x"3A",x"3B",x"4C",x"77",x"E1",x"10",x"EB",x"7E", -- 0x0E40
    x"23",x"47",x"1F",x"1F",x"1F",x"1F",x"E6",x"07", -- 0x0E48
    x"32",x"41",x"4C",x"78",x"E6",x"07",x"32",x"42", -- 0x0E50
    x"4C",x"3A",x"41",x"4C",x"06",x"00",x"4F",x"87", -- 0x0E58
    x"81",x"87",x"81",x"4F",x"28",x"04",x"11",x"71", -- 0x0E60
    x"4C",x"EF",x"3A",x"42",x"4C",x"06",x"00",x"4F", -- 0x0E68
    x"87",x"81",x"87",x"81",x"4F",x"28",x"04",x"11", -- 0x0E70
    x"8D",x"4C",x"EF",x"21",x"1F",x"28",x"11",x"B1", -- 0x0E78
    x"43",x"0E",x"01",x"CD",x"93",x"0B",x"0E",x"05", -- 0x0E80
    x"CD",x"93",x"0B",x"3E",x"BF",x"32",x"39",x"4C", -- 0x0E88
    x"11",x"00",x"14",x"CD",x"6D",x"0B",x"3A",x"27", -- 0x0E90
    x"4C",x"47",x"11",x"C0",x"FF",x"36",x"DB",x"CB", -- 0x0E98
    x"D4",x"36",x"01",x"2C",x"36",x"01",x"CB",x"94", -- 0x0EA0
    x"36",x"FB",x"2D",x"19",x"10",x"EF",x"21",x"3D", -- 0x0EA8
    x"28",x"11",x"B3",x"43",x"0E",x"19",x"CD",x"93", -- 0x0EB0
    x"0B",x"21",x"14",x"4C",x"CD",x"93",x"0B",x"21", -- 0x0EB8
    x"46",x"28",x"CD",x"93",x"0B",x"21",x"0D",x"4C", -- 0x0EC0
    x"C3",x"93",x"0B",x"06",x"08",x"11",x"F0",x"F0", -- 0x0EC8
    x"3E",x"08",x"90",x"CD",x"D5",x"0B",x"10",x"F5", -- 0x0ED0
    x"C9",x"E5",x"CD",x"6D",x"0B",x"EB",x"E1",x"E5", -- 0x0ED8
    x"D5",x"C5",x"7D",x"2C",x"12",x"CB",x"D2",x"7C", -- 0x0EE0
    x"12",x"CB",x"92",x"3E",x"E0",x"83",x"5F",x"7A", -- 0x0EE8
    x"CE",x"FF",x"57",x"0D",x"20",x"EC",x"C1",x"D1", -- 0x0EF0
    x"E1",x"13",x"7D",x"C6",x"20",x"6F",x"10",x"DF", -- 0x0EF8
    x"C9",x"E5",x"CD",x"6D",x"0B",x"EB",x"E1",x"E5", -- 0x0F00
    x"D5",x"C5",x"7D",x"12",x"CB",x"D2",x"7C",x"12", -- 0x0F08
    x"CB",x"92",x"3E",x"E0",x"83",x"5F",x"7A",x"CE", -- 0x0F10
    x"FF",x"57",x"0D",x"20",x"ED",x"C1",x"D1",x"E1", -- 0x0F18
    x"13",x"10",x"E4",x"C9",x"AF",x"CD",x"5C",x"0C", -- 0x0F20
    x"21",x"50",x"0F",x"16",x"04",x"0E",x"17",x"1E", -- 0x0F28
    x"00",x"06",x"1B",x"7E",x"23",x"E6",x"01",x"28", -- 0x0F30
    x"0D",x"E5",x"D5",x"CD",x"6D",x"0B",x"36",x"A0", -- 0x0F38
    x"CB",x"D4",x"36",x"09",x"D1",x"E1",x"1C",x"10", -- 0x0F40
    x"EA",x"14",x"0D",x"20",x"E2",x"C3",x"CB",x"0E", -- 0x0F48
    x"30",x"30",x"30",x"30",x"30",x"31",x"31",x"31", -- 0x0F50
    x"31",x"30",x"30",x"30",x"31",x"31",x"31",x"30", -- 0x0F58
    x"30",x"30",x"31",x"31",x"31",x"30",x"30",x"30", -- 0x0F60
    x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0F68
    x"31",x"30",x"30",x"30",x"31",x"30",x"31",x"30", -- 0x0F70
    x"30",x"30",x"31",x"30",x"31",x"30",x"30",x"30", -- 0x0F78
    x"31",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0F80
    x"30",x"30",x"30",x"31",x"31",x"31",x"31",x"30", -- 0x0F88
    x"30",x"31",x"31",x"31",x"31",x"31",x"30",x"31", -- 0x0F90
    x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0F98
    x"30",x"30",x"30",x"30",x"30",x"30",x"31",x"30", -- 0x0FA0
    x"30",x"30",x"30",x"30",x"31",x"30",x"30",x"30", -- 0x0FA8
    x"31",x"30",x"31",x"30",x"30",x"30",x"31",x"30", -- 0x0FB0
    x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0FB8
    x"30",x"31",x"30",x"30",x"30",x"30",x"30",x"31", -- 0x0FC0
    x"30",x"30",x"30",x"31",x"30",x"30",x"31",x"31", -- 0x0FC8
    x"31",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0FD0
    x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0FD8
    x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0FE0
    x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0FE8
    x"30",x"30",x"31",x"30",x"30",x"30",x"31",x"30", -- 0x0FF0
    x"30",x"31",x"31",x"31",x"30",x"30",x"31",x"30", -- 0x0FF8
    x"30",x"30",x"31",x"30",x"31",x"31",x"31",x"30", -- 0x1000
    x"30",x"31",x"31",x"31",x"30",x"31",x"31",x"30", -- 0x1008
    x"31",x"31",x"30",x"31",x"30",x"30",x"30",x"31", -- 0x1010
    x"30",x"31",x"31",x"30",x"30",x"31",x"30",x"30", -- 0x1018
    x"31",x"30",x"30",x"31",x"30",x"30",x"30",x"31", -- 0x1020
    x"31",x"30",x"31",x"30",x"31",x"30",x"31",x"31", -- 0x1028
    x"31",x"31",x"31",x"30",x"31",x"30",x"31",x"30", -- 0x1030
    x"31",x"30",x"30",x"31",x"30",x"30",x"31",x"30", -- 0x1038
    x"30",x"30",x"30",x"31",x"30",x"30",x"30",x"31", -- 0x1040
    x"30",x"31",x"30",x"30",x"30",x"31",x"30",x"31", -- 0x1048
    x"30",x"30",x"31",x"31",x"30",x"30",x"31",x"30", -- 0x1050
    x"30",x"31",x"30",x"30",x"30",x"31",x"31",x"30", -- 0x1058
    x"30",x"30",x"31",x"30",x"31",x"30",x"30",x"30", -- 0x1060
    x"31",x"30",x"31",x"30",x"30",x"30",x"31",x"30", -- 0x1068
    x"31",x"31",x"31",x"30",x"30",x"31",x"31",x"31", -- 0x1070
    x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x1078
    x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x1080
    x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x1088
    x"30",x"30",x"30",x"30",x"31",x"30",x"30",x"30", -- 0x1090
    x"31",x"30",x"31",x"31",x"31",x"30",x"31",x"30", -- 0x1098
    x"30",x"30",x"31",x"30",x"31",x"31",x"31",x"31", -- 0x10A0
    x"31",x"30",x"31",x"31",x"31",x"31",x"30",x"31", -- 0x10A8
    x"31",x"30",x"31",x"31",x"30",x"30",x"31",x"30", -- 0x10B0
    x"30",x"31",x"31",x"30",x"30",x"31",x"30",x"31", -- 0x10B8
    x"30",x"30",x"30",x"30",x"30",x"31",x"30",x"30", -- 0x10C0
    x"30",x"31",x"31",x"30",x"31",x"30",x"31",x"30", -- 0x10C8
    x"30",x"31",x"30",x"30",x"31",x"30",x"31",x"30", -- 0x10D0
    x"31",x"30",x"31",x"31",x"30",x"30",x"30",x"30", -- 0x10D8
    x"31",x"31",x"31",x"31",x"30",x"31",x"30",x"30", -- 0x10E0
    x"30",x"31",x"30",x"30",x"31",x"30",x"30",x"31", -- 0x10E8
    x"30",x"30",x"31",x"31",x"30",x"31",x"30",x"30", -- 0x10F0
    x"30",x"30",x"30",x"31",x"30",x"30",x"31",x"30", -- 0x10F8
    x"31",x"30",x"30",x"30",x"31",x"30",x"31",x"31", -- 0x1100
    x"31",x"30",x"31",x"30",x"30",x"30",x"31",x"30", -- 0x1108
    x"31",x"31",x"31",x"31",x"31",x"30",x"31",x"30", -- 0x1110
    x"30",x"30",x"31",x"30",x"30",x"30",x"30",x"30", -- 0x1118
    x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x1120
    x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x1128
    x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x1130
    x"30",x"30",x"30",x"31",x"30",x"30",x"30",x"31", -- 0x1138
    x"30",x"30",x"31",x"31",x"31",x"30",x"30",x"31", -- 0x1140
    x"30",x"30",x"30",x"31",x"30",x"30",x"30",x"30", -- 0x1148
    x"30",x"30",x"30",x"30",x"30",x"30",x"31",x"31", -- 0x1150
    x"30",x"31",x"31",x"30",x"31",x"30",x"30",x"30", -- 0x1158
    x"31",x"30",x"31",x"31",x"30",x"30",x"31",x"30", -- 0x1160
    x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x1168
    x"30",x"31",x"30",x"31",x"30",x"31",x"30",x"31", -- 0x1170
    x"31",x"31",x"31",x"31",x"30",x"31",x"30",x"31", -- 0x1178
    x"30",x"31",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x1180
    x"30",x"30",x"30",x"30",x"31",x"30",x"30",x"30", -- 0x1188
    x"31",x"30",x"31",x"30",x"30",x"30",x"31",x"30", -- 0x1190
    x"31",x"30",x"30",x"31",x"31",x"30",x"30",x"30", -- 0x1198
    x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"31", -- 0x11A0
    x"30",x"30",x"30",x"31",x"30",x"31",x"30",x"30", -- 0x11A8
    x"30",x"31",x"30",x"31",x"30",x"30",x"30",x"31", -- 0x11B0
    x"30",x"30",x"30",x"30",x"30",x"20",x"20",x"20", -- 0x11B8
    x"20",x"50",x"72",x"65",x"73",x"73",x"20",x"53", -- 0x11C0
    x"74",x"61",x"72",x"74",x"20",x"54",x"6F",x"20", -- 0x11C8
    x"50",x"6C",x"61",x"79",x"20",x"20",x"20",x"20", -- 0x11D0
    x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20", -- 0x11D8
    x"20",x"49",x"6E",x"73",x"65",x"72",x"74",x"20", -- 0x11E0
    x"43",x"6F",x"69",x"6E",x"20",x"20",x"20",x"20", -- 0x11E8
    x"20",x"20",x"20",x"20",x"00",x"1E",x"00",x"D6", -- 0x11F0
    x"0A",x"38",x"03",x"1C",x"18",x"F9",x"C6",x"0A", -- 0x11F8
    x"C9",x"3A",x"0A",x"4C",x"B7",x"C0",x"3A",x"00", -- 0x1200
    x"50",x"32",x"04",x"4C",x"2F",x"5F",x"3A",x"06", -- 0x1208
    x"4C",x"57",x"2F",x"A3",x"32",x"07",x"4C",x"7B", -- 0x1210
    x"32",x"06",x"4C",x"3A",x"40",x"50",x"32",x"05", -- 0x1218
    x"4C",x"2F",x"5F",x"3A",x"08",x"4C",x"57",x"2F", -- 0x1220
    x"A3",x"32",x"09",x"4C",x"7B",x"32",x"08",x"4C", -- 0x1228
    x"3A",x"09",x"4C",x"E6",x"01",x"28",x"08",x"3A", -- 0x1230
    x"4C",x"4C",x"EE",x"0F",x"32",x"4C",x"4C",x"3A", -- 0x1238
    x"09",x"4C",x"E6",x"08",x"28",x"08",x"3A",x"4D", -- 0x1240
    x"4C",x"EE",x"0F",x"32",x"4D",x"4C",x"3A",x"07", -- 0x1248
    x"4C",x"E6",x"20",x"28",x"13",x"3A",x"0B",x"4C", -- 0x1250
    x"FE",x"63",x"28",x"0C",x"3C",x"32",x"0B",x"4C", -- 0x1258
    x"CD",x"69",x"12",x"3E",x"01",x"32",x"0C",x"4C", -- 0x1260
    x"C9",x"11",x"99",x"12",x"21",x"FD",x"43",x"1A", -- 0x1268
    x"13",x"B7",x"28",x"0C",x"C6",x"80",x"77",x"CB", -- 0x1270
    x"D4",x"36",x"19",x"CB",x"94",x"2D",x"18",x"EF", -- 0x1278
    x"3A",x"0B",x"4C",x"CD",x"F5",x"11",x"57",x"7B", -- 0x1280
    x"C6",x"B0",x"77",x"CB",x"D4",x"36",x"19",x"2D", -- 0x1288
    x"36",x"19",x"CB",x"94",x"7A",x"C6",x"B0",x"77", -- 0x1290
    x"C9",x"43",x"72",x"65",x"64",x"69",x"74",x"73", -- 0x1298
    x"20",x"00",x"32",x"47",x"4C",x"AF",x"32",x"46", -- 0x12A0
    x"4C",x"3E",x"01",x"32",x"4B",x"4C",x"C9",x"CD", -- 0x12A8
    x"01",x"12",x"3A",x"47",x"4C",x"B7",x"CA",x"A1", -- 0x12B0
    x"13",x"3A",x"4B",x"4C",x"D6",x"04",x"32",x"4B", -- 0x12B8
    x"4C",x"D2",x"10",x"13",x"3A",x"47",x"4C",x"87", -- 0x12C0
    x"5F",x"16",x"00",x"21",x"4F",x"14",x"19",x"5E", -- 0x12C8
    x"23",x"56",x"EB",x"3A",x"46",x"4C",x"5F",x"3C", -- 0x12D0
    x"32",x"46",x"4C",x"16",x"00",x"19",x"19",x"19", -- 0x12D8
    x"7E",x"FE",x"FF",x"CA",x"A1",x"13",x"B7",x"20", -- 0x12E0
    x"14",x"3C",x"32",x"46",x"4C",x"3A",x"47",x"4C", -- 0x12E8
    x"87",x"5F",x"16",x"00",x"21",x"4F",x"14",x"19", -- 0x12F0
    x"5E",x"23",x"56",x"EB",x"7E",x"32",x"4B",x"4C", -- 0x12F8
    x"23",x"7E",x"CD",x"FD",x"13",x"32",x"48",x"4C", -- 0x1300
    x"23",x"7E",x"CD",x"FD",x"13",x"32",x"49",x"4C", -- 0x1308
    x"3A",x"24",x"4C",x"B7",x"28",x"16",x"3A",x"2A", -- 0x1310
    x"4C",x"3C",x"32",x"2A",x"4C",x"1F",x"1F",x"E6", -- 0x1318
    x"3F",x"5F",x"16",x"00",x"21",x"AE",x"13",x"19", -- 0x1320
    x"7E",x"32",x"4A",x"4C",x"3A",x"4F",x"4C",x"B7", -- 0x1328
    x"28",x"10",x"C6",x"02",x"32",x"4F",x"4C",x"32", -- 0x1330
    x"4A",x"4C",x"FE",x"40",x"38",x"04",x"AF",x"32", -- 0x1338
    x"4F",x"4C",x"3A",x"0C",x"4C",x"B7",x"28",x"10", -- 0x1340
    x"C6",x"01",x"32",x"0C",x"4C",x"32",x"4A",x"4C", -- 0x1348
    x"FE",x"20",x"38",x"04",x"AF",x"32",x"0C",x"4C", -- 0x1350
    x"3A",x"4E",x"4C",x"B7",x"28",x"08",x"D6",x"04", -- 0x1358
    x"32",x"4E",x"4C",x"32",x"4A",x"4C",x"DD",x"21", -- 0x1360
    x"45",x"50",x"DD",x"36",x"00",x"01",x"ED",x"4B", -- 0x1368
    x"4C",x"4C",x"3A",x"48",x"4C",x"CD",x"16",x"14", -- 0x1370
    x"DD",x"21",x"4A",x"50",x"DD",x"36",x"00",x"03", -- 0x1378
    x"ED",x"4B",x"4C",x"4C",x"3A",x"49",x"4C",x"CD", -- 0x1380
    x"16",x"14",x"DD",x"21",x"4F",x"50",x"DD",x"36", -- 0x1388
    x"00",x"01",x"ED",x"4B",x"4D",x"4C",x"3A",x"4A", -- 0x1390
    x"4C",x"CD",x"16",x"14",x"AF",x"32",x"4A",x"4C", -- 0x1398
    x"C9",x"AF",x"32",x"48",x"4C",x"32",x"49",x"4C", -- 0x13A0
    x"32",x"47",x"4C",x"C3",x"10",x"13",x"04",x"09", -- 0x13A8
    x"0B",x"0D",x"0F",x"11",x"13",x"15",x"16",x"15", -- 0x13B0
    x"13",x"11",x"0F",x"0D",x"0B",x"09",x"09",x"08", -- 0x13B8
    x"08",x"07",x"07",x"06",x"06",x"05",x"05",x"04", -- 0x13C0
    x"04",x"04",x"03",x"03",x"03",x"03",x"02",x"02", -- 0x13C8
    x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01", -- 0x13D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x13D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x13E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x13E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x13F0
    x"00",x"00",x"00",x"00",x"00",x"FE",x"FF",x"C8", -- 0x13F8
    x"B7",x"C8",x"E5",x"D5",x"5F",x"21",x"44",x"16", -- 0x1400
    x"16",x"00",x"BE",x"28",x"05",x"23",x"23",x"14", -- 0x1408
    x"18",x"F8",x"7A",x"D1",x"E1",x"C9",x"E5",x"D5", -- 0x1410
    x"B7",x"28",x"2D",x"87",x"5F",x"16",x"00",x"21", -- 0x1418
    x"AC",x"16",x"19",x"5E",x"23",x"56",x"7B",x"DD", -- 0x1420
    x"77",x"0C",x"1F",x"1F",x"1F",x"1F",x"DD",x"77", -- 0x1428
    x"0D",x"7A",x"DD",x"77",x"0E",x"1F",x"1F",x"1F", -- 0x1430
    x"1F",x"DD",x"77",x"0F",x"79",x"DD",x"77",x"10", -- 0x1438
    x"3E",x"01",x"32",x"01",x"50",x"D1",x"E1",x"C9", -- 0x1440
    x"DD",x"36",x"10",x"00",x"D1",x"E1",x"C9",x"00", -- 0x1448
    x"00",x"55",x"14",x"81",x"15",x"50",x"80",x"80", -- 0x1450
    x"50",x"66",x"66",x"50",x"56",x"56",x"32",x"56", -- 0x1458
    x"56",x"32",x"AB",x"CB",x"32",x"2B",x"33",x"32", -- 0x1460
    x"2B",x"33",x"32",x"AB",x"CB",x"32",x"33",x"40", -- 0x1468
    x"32",x"33",x"40",x"32",x"AB",x"CB",x"32",x"80", -- 0x1470
    x"80",x"32",x"80",x"80",x"32",x"66",x"66",x"32", -- 0x1478
    x"56",x"56",x"32",x"60",x"56",x"32",x"AB",x"C0", -- 0x1480
    x"32",x"2B",x"30",x"32",x"2B",x"30",x"32",x"AB", -- 0x1488
    x"C0",x"32",x"30",x"44",x"32",x"30",x"44",x"32", -- 0x1490
    x"AB",x"C0",x"32",x"88",x"88",x"32",x"88",x"88", -- 0x1498
    x"32",x"72",x"72",x"32",x"4C",x"4C",x"32",x"4C", -- 0x14A0
    x"4C",x"32",x"AB",x"C0",x"32",x"26",x"30",x"32", -- 0x14A8
    x"26",x"30",x"32",x"AB",x"C0",x"32",x"30",x"44", -- 0x14B0
    x"32",x"30",x"44",x"32",x"AB",x"C0",x"32",x"88", -- 0x14B8
    x"88",x"32",x"88",x"88",x"32",x"72",x"72",x"32", -- 0x14C0
    x"4C",x"4C",x"32",x"4C",x"4C",x"32",x"AB",x"CB", -- 0x14C8
    x"32",x"26",x"33",x"32",x"26",x"33",x"32",x"AB", -- 0x14D0
    x"CB",x"32",x"33",x"40",x"32",x"33",x"40",x"32", -- 0x14D8
    x"AB",x"CB",x"32",x"80",x"80",x"32",x"80",x"80", -- 0x14E0
    x"32",x"66",x"66",x"32",x"56",x"56",x"32",x"40", -- 0x14E8
    x"40",x"32",x"80",x"AB",x"32",x"20",x"2B",x"32", -- 0x14F0
    x"20",x"2B",x"32",x"80",x"AB",x"32",x"2B",x"33", -- 0x14F8
    x"32",x"2B",x"33",x"32",x"80",x"AB",x"32",x"80", -- 0x1500
    x"80",x"32",x"80",x"80",x"32",x"66",x"66",x"32", -- 0x1508
    x"56",x"56",x"32",x"40",x"40",x"32",x"80",x"98", -- 0x1510
    x"32",x"20",x"26",x"32",x"20",x"26",x"32",x"80", -- 0x1518
    x"98",x"32",x"26",x"30",x"32",x"26",x"30",x"32", -- 0x1520
    x"00",x"00",x"32",x"72",x"72",x"32",x"72",x"72", -- 0x1528
    x"32",x"60",x"60",x"32",x"4C",x"4C",x"32",x"4C", -- 0x1530
    x"98",x"32",x"4C",x"4C",x"32",x"4C",x"4C",x"32", -- 0x1538
    x"4C",x"98",x"32",x"5B",x"5B",x"32",x"56",x"56", -- 0x1540
    x"32",x"33",x"CB",x"32",x"33",x"33",x"32",x"33", -- 0x1548
    x"33",x"32",x"33",x"CB",x"32",x"40",x"40",x"32", -- 0x1550
    x"66",x"66",x"64",x"66",x"66",x"32",x"72",x"72", -- 0x1558
    x"64",x"4C",x"4C",x"32",x"56",x"56",x"32",x"80", -- 0x1560
    x"CB",x"19",x"80",x"00",x"19",x"80",x"80",x"32", -- 0x1568
    x"80",x"CB",x"FA",x"00",x"00",x"FA",x"00",x"00", -- 0x1570
    x"FA",x"00",x"00",x"FA",x"00",x"00",x"00",x"00", -- 0x1578
    x"00",x"32",x"80",x"80",x"32",x"72",x"72",x"32", -- 0x1580
    x"66",x"66",x"32",x"60",x"60",x"32",x"56",x"56", -- 0x1588
    x"32",x"66",x"66",x"32",x"56",x"56",x"32",x"56", -- 0x1590
    x"56",x"32",x"51",x"51",x"32",x"60",x"60",x"32", -- 0x1598
    x"51",x"51",x"32",x"51",x"51",x"32",x"56",x"56", -- 0x15A0
    x"32",x"66",x"66",x"32",x"56",x"56",x"32",x"56", -- 0x15A8
    x"56",x"32",x"80",x"80",x"32",x"72",x"72",x"32", -- 0x15B0
    x"66",x"66",x"32",x"60",x"60",x"32",x"56",x"56", -- 0x15B8
    x"32",x"66",x"66",x"32",x"56",x"56",x"32",x"56", -- 0x15C0
    x"56",x"32",x"51",x"51",x"32",x"60",x"60",x"32", -- 0x15C8
    x"51",x"51",x"32",x"51",x"51",x"32",x"56",x"56", -- 0x15D0
    x"32",x"56",x"56",x"32",x"56",x"56",x"32",x"56", -- 0x15D8
    x"56",x"32",x"80",x"80",x"32",x"72",x"72",x"32", -- 0x15E0
    x"66",x"66",x"32",x"60",x"60",x"32",x"56",x"56", -- 0x15E8
    x"32",x"66",x"66",x"32",x"56",x"56",x"32",x"56", -- 0x15F0
    x"56",x"32",x"51",x"51",x"32",x"60",x"60",x"32", -- 0x15F8
    x"51",x"51",x"32",x"51",x"51",x"32",x"56",x"56", -- 0x1600
    x"32",x"66",x"66",x"32",x"56",x"56",x"32",x"56", -- 0x1608
    x"56",x"32",x"80",x"80",x"32",x"72",x"72",x"32", -- 0x1610
    x"66",x"66",x"32",x"60",x"60",x"32",x"56",x"56", -- 0x1618
    x"32",x"66",x"66",x"32",x"56",x"56",x"32",x"40", -- 0x1620
    x"40",x"32",x"56",x"56",x"32",x"66",x"66",x"32", -- 0x1628
    x"80",x"80",x"32",x"66",x"66",x"32",x"56",x"56", -- 0x1630
    x"32",x"56",x"56",x"32",x"56",x"56",x"32",x"56", -- 0x1638
    x"56",x"00",x"00",x"00",x"00",x"24",x"FF",x"24", -- 0x1640
    x"F2",x"04",x"E6",x"25",x"D8",x"05",x"CB",x"26", -- 0x1648
    x"C0",x"27",x"B4",x"07",x"AB",x"28",x"A2",x"08", -- 0x1650
    x"98",x"29",x"90",x"09",x"88",x"2A",x"80",x"2B", -- 0x1658
    x"79",x"0B",x"72",x"2C",x"6C",x"0C",x"66",x"2D", -- 0x1660
    x"60",x"2E",x"5B",x"0E",x"56",x"2F",x"51",x"0F", -- 0x1668
    x"4C",x"30",x"48",x"10",x"44",x"31",x"40",x"32", -- 0x1670
    x"3C",x"12",x"39",x"33",x"36",x"13",x"33",x"34", -- 0x1678
    x"30",x"35",x"2D",x"15",x"2B",x"36",x"28",x"16", -- 0x1680
    x"26",x"37",x"24",x"17",x"22",x"38",x"20",x"39", -- 0x1688
    x"1F",x"19",x"1D",x"3A",x"1B",x"1A",x"19",x"3B", -- 0x1690
    x"18",x"3C",x"17",x"1C",x"16",x"3D",x"14",x"1D", -- 0x1698
    x"13",x"3E",x"12",x"1E",x"11",x"3F",x"10",x"2B", -- 0x16A0
    x"01",x"01",x"01",x"01",x"57",x"00",x"5C",x"00", -- 0x16A8
    x"62",x"00",x"6A",x"00",x"6F",x"00",x"75",x"00", -- 0x16B0
    x"7D",x"00",x"85",x"00",x"8E",x"00",x"96",x"00", -- 0x16B8
    x"9E",x"00",x"A6",x"00",x"AE",x"00",x"B9",x"00", -- 0x16C0
    x"C4",x"00",x"D5",x"00",x"DF",x"00",x"EA",x"00", -- 0x16C8
    x"FB",x"00",x"0B",x"01",x"1C",x"01",x"2C",x"01", -- 0x16D0
    x"3C",x"01",x"4D",x"01",x"5D",x"01",x"73",x"01", -- 0x16D8
    x"89",x"01",x"AA",x"01",x"BF",x"01",x"D5",x"01", -- 0x16E0
    x"F6",x"01",x"17",x"02",x"38",x"02",x"58",x"02", -- 0x16E8
    x"79",x"02",x"9A",x"02",x"BA",x"02",x"E6",x"02", -- 0x16F0
    x"12",x"03",x"54",x"03",x"7E",x"03",x"AA",x"03", -- 0x16F8
    x"EC",x"03",x"2E",x"04",x"70",x"04",x"B0",x"04", -- 0x1700
    x"F2",x"04",x"34",x"05",x"74",x"05",x"CC",x"05", -- 0x1708
    x"24",x"06",x"A8",x"06",x"FC",x"06",x"54",x"07", -- 0x1710
    x"D8",x"07",x"5C",x"08",x"E0",x"08",x"60",x"09", -- 0x1718
    x"E4",x"09",x"68",x"0A",x"E8",x"0A",x"98",x"0B", -- 0x1720
    x"48",x"0C",x"50",x"0D",x"F8",x"0D",x"A8",x"0E", -- 0x1728
    x"B0",x"0F",x"B8",x"10",x"C0",x"11",x"C0",x"12", -- 0x1730
    x"C8",x"13",x"D0",x"14",x"E8",x"0A",x"98",x"0B", -- 0x1738
    x"48",x"0C",x"50",x"0D",x"F8",x"0D",x"A8",x"0E", -- 0x1740
    x"B0",x"0F",x"B8",x"10",x"C0",x"11",x"C0",x"12", -- 0x1748
    x"C8",x"13",x"D0",x"14",x"E8",x"0A",x"98",x"0B", -- 0x1750
    x"48",x"0C",x"50",x"0D",x"F8",x"0D",x"A8",x"0E", -- 0x1758
    x"B0",x"0F",x"B8",x"10",x"C0",x"11",x"C0",x"12", -- 0x1760
    x"C8",x"13",x"D0",x"14",x"E8",x"0A",x"98",x"0B", -- 0x1768
    x"48",x"0C",x"50",x"0D",x"F8",x"0D",x"A8",x"0E", -- 0x1770
    x"B0",x"0F",x"B8",x"10",x"C0",x"11",x"C0",x"12", -- 0x1778
    x"C8",x"13",x"D0",x"14",x"AC",x"17",x"30",x"18", -- 0x1780
    x"D3",x"18",x"67",x"19",x"1F",x"1A",x"C9",x"1A", -- 0x1788
    x"71",x"1B",x"2F",x"1C",x"13",x"1D",x"CC",x"1D", -- 0x1790
    x"A0",x"1E",x"77",x"1F",x"59",x"20",x"13",x"21", -- 0x1798
    x"FA",x"21",x"AF",x"22",x"68",x"23",x"3E",x"24", -- 0x17A0
    x"F2",x"24",x"A6",x"25",x"00",x"00",x"05",x"1C", -- 0x17A8
    x"08",x"01",x"0C",x"05",x"04",x"80",x"01",x"11", -- 0x17B0
    x"05",x"04",x"80",x"01",x"00",x"07",x"03",x"08", -- 0x17B8
    x"01",x"11",x"08",x"03",x"20",x"09",x"00",x"09", -- 0x17C0
    x"04",x"08",x"01",x"08",x"09",x"10",x"58",x"0F", -- 0x17C8
    x"1A",x"0A",x"02",x"08",x"01",x"14",x"0C",x"03", -- 0x17D0
    x"20",x"09",x"17",x"0C",x"03",x"80",x"01",x"1A", -- 0x17D8
    x"0C",x"02",x"08",x"01",x"04",x"0D",x"10",x"08", -- 0x17E0
    x"01",x"00",x"0F",x"1C",x"08",x"01",x"1A",x"0D", -- 0x17E8
    x"00",x"04",x"30",x"0F",x"17",x"04",x"1B",x"04", -- 0x17F0
    x"15",x"08",x"0C",x"0C",x"02",x"38",x"05",x"0B", -- 0x17F8
    x"00",x"10",x"00",x"07",x"43",x"45",x"4E",x"54", -- 0x1800
    x"52",x"41",x"4C",x"20",x"43",x"41",x"56",x"45", -- 0x1808
    x"52",x"4E",x"00",x"08",x"09",x"10",x"58",x"0F", -- 0x1810
    x"00",x"01",x"0D",x"05",x"45",x"07",x"09",x"00", -- 0x1818
    x"10",x"01",x"19",x"00",x"18",x"04",x"1B",x"06", -- 0x1820
    x"10",x"28",x"08",x"38",x"40",x"40",x"7E",x"01", -- 0x1828
    x"01",x"10",x"00",x"0C",x"20",x"09",x"12",x"03", -- 0x1830
    x"03",x"88",x"01",x"15",x"03",x"01",x"09",x"01", -- 0x1838
    x"00",x"05",x"12",x"09",x"01",x"12",x"06",x"02", -- 0x1840
    x"09",x"01",x"00",x"07",x"01",x"09",x"01",x"01", -- 0x1848
    x"07",x"04",x"88",x"01",x"08",x"09",x"07",x"09", -- 0x1850
    x"01",x"11",x"0A",x"04",x"88",x"01",x"0D",x"0C", -- 0x1858
    x"03",x"09",x"01",x"07",x"0D",x"03",x"88",x"01", -- 0x1860
    x"00",x"0F",x"1C",x"09",x"01",x"16",x"06",x"87", -- 0x1868
    x"20",x"09",x"19",x"05",x"88",x"20",x"09",x"17", -- 0x1870
    x"06",x"02",x"88",x"01",x"17",x"08",x"02",x"88", -- 0x1878
    x"01",x"17",x"09",x"02",x"88",x"01",x"17",x"0A", -- 0x1880
    x"02",x"88",x"01",x"17",x"0B",x"02",x"88",x"01", -- 0x1888
    x"17",x"0C",x"02",x"88",x"01",x"1A",x"0D",x"00", -- 0x1890
    x"00",x"31",x"07",x"01",x"39",x"05",x"1B",x"01", -- 0x1898
    x"08",x"54",x"48",x"45",x"20",x"43",x"4F",x"4C", -- 0x18A0
    x"44",x"20",x"52",x"4F",x"4F",x"4D",x"00",x"02", -- 0x18A8
    x"0B",x"04",x"58",x"14",x"01",x"01",x"0D",x"05", -- 0x18B0
    x"44",x"07",x"02",x"09",x"07",x"01",x"15",x"01", -- 0x18B8
    x"18",x"07",x"11",x"0C",x"20",x"30",x"10",x"18", -- 0x18C0
    x"80",x"08",x"80",x"FF",x"30",x"13",x"68",x"98", -- 0x18C8
    x"58",x"D4",x"FF",x"00",x"09",x"00",x"01",x"1C", -- 0x18D0
    x"03",x"11",x"00",x"01",x"1B",x"03",x"11",x"01", -- 0x18D8
    x"01",x"1C",x"03",x"1A",x"00",x"01",x"1C",x"03", -- 0x18E0
    x"00",x"05",x"04",x"0A",x"05",x"04",x"05",x"18", -- 0x18E8
    x"98",x"05",x"00",x"07",x"05",x"0A",x"05",x"19", -- 0x18F0
    x"07",x"03",x"0A",x"05",x"00",x"08",x"83",x"1B", -- 0x18F8
    x"03",x"00",x"0B",x"01",x"1C",x"03",x"05",x"09", -- 0x1900
    x"06",x"48",x"01",x"17",x"0A",x"05",x"0A",x"05", -- 0x1908
    x"0C",x"0B",x"05",x"0A",x"05",x"04",x"0C",x"06", -- 0x1910
    x"0A",x"05",x"13",x"0D",x"09",x"0A",x"05",x"00", -- 0x1918
    x"0F",x"1C",x"0A",x"05",x"1A",x"08",x"00",x"00", -- 0x1920
    x"1B",x"07",x"00",x"1C",x"05",x"08",x"54",x"48", -- 0x1928
    x"45",x"20",x"4D",x"45",x"4E",x"41",x"47",x"45", -- 0x1930
    x"52",x"49",x"45",x"00",x"05",x"09",x"06",x"48", -- 0x1938
    x"01",x"00",x"01",x"0D",x"05",x"45",x"1B",x"05", -- 0x1940
    x"00",x"0D",x"00",x"15",x"00",x"12",x"06",x"19", -- 0x1948
    x"06",x"30",x"40",x"13",x"68",x"A0",x"08",x"D0", -- 0x1950
    x"FF",x"40",x"10",x"18",x"50",x"08",x"68",x"FF", -- 0x1958
    x"40",x"12",x"18",x"90",x"78",x"D0",x"01",x"00", -- 0x1960
    x"06",x"00",x"01",x"1C",x"03",x"0D",x"00",x"0F", -- 0x1968
    x"20",x"05",x"12",x"03",x"05",x"0A",x"07",x"19", -- 0x1970
    x"04",x"03",x"0A",x"07",x"00",x"05",x"01",x"0A", -- 0x1978
    x"07",x"06",x"05",x"01",x"0A",x"07",x"10",x"05", -- 0x1980
    x"01",x"0A",x"07",x"0B",x"06",x"02",x"0A",x"07", -- 0x1988
    x"14",x"06",x"03",x"0A",x"07",x"00",x"07",x"03", -- 0x1990
    x"98",x"14",x"06",x"08",x"02",x"0A",x"07",x"18", -- 0x1998
    x"08",x"04",x"0A",x"07",x"11",x"09",x"03",x"0A", -- 0x19A0
    x"07",x"00",x"0A",x"03",x"48",x"05",x"1B",x"0A", -- 0x19A8
    x"01",x"0A",x"07",x"0B",x"0B",x"03",x"0A",x"07", -- 0x19B0
    x"15",x"0B",x"03",x"0A",x"07",x"05",x"0C",x"02", -- 0x19B8
    x"0A",x"07",x"16",x"0C",x"01",x"1C",x"03",x"19", -- 0x19C0
    x"0C",x"03",x"0A",x"07",x"11",x"0D",x"02",x"0A", -- 0x19C8
    x"07",x"00",x"0F",x"1C",x"0A",x"07",x"1A",x"01", -- 0x19D0
    x"00",x"00",x"1B",x"07",x"00",x"1C",x"05",x"01", -- 0x19D8
    x"41",x"42",x"41",x"4E",x"44",x"4F",x"4E",x"45", -- 0x19E0
    x"44",x"20",x"55",x"52",x"41",x"4E",x"49",x"55", -- 0x19E8
    x"4D",x"20",x"57",x"4F",x"52",x"4B",x"49",x"4E", -- 0x19F0
    x"47",x"53",x"00",x"00",x"0A",x"03",x"48",x"05", -- 0x19F8
    x"01",x"1A",x"0D",x"05",x"45",x"1B",x"00",x"00", -- 0x1A00
    x"0B",x"01",x"16",x"01",x"0F",x"07",x"19",x"07", -- 0x1A08
    x"20",x"50",x"08",x"68",x"08",x"08",x"60",x"01", -- 0x1A10
    x"50",x"28",x"68",x"28",x"20",x"78",x"01",x"09", -- 0x1A18
    x"12",x"00",x"01",x"3A",x"01",x"00",x"05",x"0C", -- 0x1A20
    x"0C",x"0F",x"10",x"05",x"04",x"68",x"0F",x"14", -- 0x1A28
    x"05",x"05",x"0C",x"0F",x"1A",x"06",x"02",x"0C", -- 0x1A30
    x"0F",x"10",x"08",x"09",x"48",x"01",x"03",x"09", -- 0x1A38
    x"09",x"0C",x"0F",x"00",x"0B",x"02",x"68",x"0F", -- 0x1A40
    x"02",x"0B",x"0A",x"0C",x"0F",x"10",x"0B",x"06", -- 0x1A48
    x"0C",x"0F",x"1B",x"0B",x"01",x"0C",x"0F",x"00", -- 0x1A50
    x"0D",x"02",x"0C",x"0F",x"00",x"0F",x"1C",x"0C", -- 0x1A58
    x"0F",x"07",x"0C",x"83",x"23",x"0F",x"0C",x"0D", -- 0x1A60
    x"82",x"23",x"0F",x"0F",x"0D",x"82",x"23",x"0F", -- 0x1A68
    x"10",x"0E",x"06",x"23",x"0F",x"07",x"0F",x"0F", -- 0x1A70
    x"23",x"0F",x"0D",x"0D",x"00",x"05",x"33",x"09", -- 0x1A78
    x"14",x"07",x"17",x"04",x"04",x"0E",x"16",x"0E", -- 0x1A80
    x"17",x"0E",x"01",x"3A",x"01",x"12",x"00",x"08", -- 0x1A88
    x"45",x"55",x"47",x"45",x"4E",x"45",x"27",x"53", -- 0x1A90
    x"20",x"4C",x"41",x"49",x"52",x"00",x"10",x"08", -- 0x1A98
    x"09",x"48",x"01",x"00",x"00",x"03",x"05",x"44", -- 0x1AA0
    x"09",x"1B",x"01",x"1A",x"07",x"09",x"06",x"08", -- 0x1AA8
    x"0C",x"06",x"0C",x"21",x"60",x"50",x"18",x"50", -- 0x1AB0
    x"08",x"50",x"FF",x"60",x"20",x"38",x"20",x"20", -- 0x1AB8
    x"50",x"01",x"1C",x"0D",x"08",x"68",x"08",x"58", -- 0x1AC0
    x"01",x"00",x"14",x"04",x"01",x"3B",x"07",x"07", -- 0x1AC8
    x"05",x"03",x"0D",x"0F",x"0E",x"05",x"02",x"0D", -- 0x1AD0
    x"0F",x"14",x"05",x"05",x"0D",x"0F",x"02",x"06", -- 0x1AD8
    x"02",x"0D",x"0F",x"0F",x"06",x"82",x"24",x"09", -- 0x1AE0
    x"1A",x"06",x"02",x"0D",x"0F",x"15",x"08",x"04", -- 0x1AE8
    x"0D",x"0F",x"00",x"09",x"02",x"0D",x"0F",x"06", -- 0x1AF0
    x"0A",x"09",x"0D",x"0F",x"0F",x"0A",x"83",x"24", -- 0x1AF8
    x"09",x"10",x"0A",x"08",x"0D",x"0F",x"10",x"0B", -- 0x1B00
    x"01",x"3B",x"07",x"02",x"0C",x"01",x"34",x"03", -- 0x1B08
    x"1A",x"0C",x"02",x"0D",x"0F",x"02",x"0D",x"04", -- 0x1B10
    x"58",x"0F",x"15",x"0D",x"02",x"0D",x"0F",x"00", -- 0x1B18
    x"0F",x"1C",x"0D",x"0F",x"1A",x"00",x"00",x"00", -- 0x1B20
    x"33",x"01",x"00",x"3A",x"01",x"06",x"50",x"52", -- 0x1B28
    x"4F",x"43",x"45",x"53",x"53",x"49",x"4E",x"47", -- 0x1B30
    x"20",x"50",x"4C",x"41",x"4E",x"54",x"00",x"02", -- 0x1B38
    x"0D",x"04",x"58",x"0F",x"00",x"0F",x"03",x"05", -- 0x1B40
    x"45",x"1B",x"00",x"0A",x"0B",x"0B",x"0E",x"06", -- 0x1B48
    x"10",x"06",x"1B",x"07",x"40",x"70",x"30",x"40", -- 0x1B50
    x"30",x"30",x"60",x"01",x"70",x"70",x"40",x"70", -- 0x1B58
    x"70",x"A0",x"01",x"70",x"38",x"68",x"38",x"38", -- 0x1B60
    x"98",x"01",x"70",x"B8",x"68",x"B8",x"B8",x"D8", -- 0x1B68
    x"01",x"00",x"0D",x"00",x"0F",x"25",x"05",x"0E", -- 0x1B70
    x"03",x"02",x"0B",x"09",x"10",x"03",x"8A",x"25", -- 0x1B78
    x"05",x"11",x"03",x"0B",x"90",x"01",x"11",x"04", -- 0x1B80
    x"0B",x"90",x"01",x"06",x"05",x"04",x"58",x"0F", -- 0x1B88
    x"0D",x"05",x"03",x"0B",x"09",x"11",x"05",x"0B", -- 0x1B90
    x"90",x"01",x"00",x"06",x"03",x"0B",x"09",x"11", -- 0x1B98
    x"06",x"0B",x"90",x"01",x"11",x"07",x"0B",x"90", -- 0x1BA0
    x"01",x"00",x"08",x"01",x"0B",x"09",x"11",x"08", -- 0x1BA8
    x"0B",x"90",x"01",x"0D",x"09",x"03",x"0B",x"09", -- 0x1BB0
    x"11",x"09",x"0B",x"90",x"01",x"01",x"0A",x"0A", -- 0x1BB8
    x"0B",x"09",x"11",x"0A",x"0B",x"90",x"01",x"11", -- 0x1BC0
    x"0B",x"0B",x"90",x"01",x"0D",x"0C",x"03",x"25", -- 0x1BC8
    x"05",x"11",x"0C",x"0B",x"90",x"01",x"08",x"0D", -- 0x1BD0
    x"03",x"0B",x"09",x"0D",x"0D",x"82",x"25",x"05", -- 0x1BD8
    x"00",x"0F",x"1C",x"0B",x"09",x"0D",x"0F",x"0F", -- 0x1BE0
    x"25",x"05",x"0E",x"0D",x"00",x"00",x"34",x"01", -- 0x1BE8
    x"04",x"18",x"09",x"19",x"05",x"16",x"08",x"19", -- 0x1BF0
    x"0A",x"16",x"0C",x"0B",x"54",x"48",x"45",x"20", -- 0x1BF8
    x"56",x"41",x"54",x"00",x"06",x"05",x"04",x"58", -- 0x1C00
    x"0F",x"01",x"00",x"0D",x"05",x"45",x"1B",x"1B", -- 0x1C08
    x"03",x"13",x"06",x"18",x"07",x"12",x"0A",x"1B", -- 0x1C10
    x"0B",x"30",x"80",x"70",x"08",x"70",x"70",x"D0", -- 0x1C18
    x"01",x"80",x"08",x"40",x"08",x"08",x"50",x"01", -- 0x1C20
    x"80",x"80",x"68",x"80",x"80",x"D0",x"01",x"00", -- 0x1C28
    x"01",x"00",x"01",x"3C",x"09",x"09",x"00",x"01", -- 0x1C30
    x"3C",x"09",x"13",x"00",x"82",x"26",x"09",x"10", -- 0x1C38
    x"00",x"8F",x"26",x"09",x"0E",x"02",x"02",x"08", -- 0x1C40
    x"01",x"1A",x"02",x"02",x"08",x"01",x"00",x"05", -- 0x1C48
    x"03",x"08",x"01",x"08",x"05",x"06",x"08",x"01", -- 0x1C50
    x"11",x"05",x"02",x"08",x"01",x"14",x"06",x"02", -- 0x1C58
    x"08",x"01",x"1B",x"06",x"01",x"08",x"01",x"01", -- 0x1C60
    x"07",x"03",x"08",x"01",x"18",x"07",x"01",x"08", -- 0x1C68
    x"01",x"07",x"08",x"03",x"08",x"01",x"11",x"09", -- 0x1C70
    x"03",x"08",x"01",x"00",x"0A",x"01",x"08",x"01", -- 0x1C78
    x"0B",x"0A",x"03",x"08",x"01",x"18",x"0A",x"03", -- 0x1C80
    x"08",x"01",x"08",x"0B",x"02",x"08",x"01",x"03", -- 0x1C88
    x"0C",x"02",x"08",x"01",x"15",x"0C",x"04",x"08", -- 0x1C90
    x"01",x"0A",x"0D",x"02",x"58",x"0F",x"0D",x"0D", -- 0x1C98
    x"82",x"26",x"09",x"11",x"0D",x"02",x"08",x"01", -- 0x1CA0
    x"15",x"0E",x"01",x"30",x"0F",x"00",x"0F",x"1C", -- 0x1CA8
    x"08",x"01",x"05",x"00",x"01",x"46",x"0F",x"11", -- 0x1CB0
    x"00",x"01",x"46",x"0F",x"0E",x"0D",x"00",x"00", -- 0x1CB8
    x"33",x"01",x"00",x"3A",x"01",x"00",x"4D",x"49", -- 0x1CC0
    x"4E",x"45",x"52",x"20",x"57",x"49",x"4C",x"4C", -- 0x1CC8
    x"59",x"20",x"4D",x"45",x"45",x"54",x"53",x"20", -- 0x1CD0
    x"4B",x"4F",x"4E",x"47",x"20",x"42",x"45",x"41", -- 0x1CD8
    x"53",x"54",x"00",x"0A",x"0D",x"03",x"58",x"0F", -- 0x1CE0
    x"00",x"00",x"0D",x"04",x"45",x"1B",x"0C",x"02", -- 0x1CE8
    x"0D",x"06",x"01",x"08",x"1A",x"0D",x"31",x"A0", -- 0x1CF0
    x"44",x"68",x"44",x"00",x"48",x"FF",x"A0",x"68", -- 0x1CF8
    x"58",x"68",x"54",x"74",x"01",x"A0",x"88",x"38", -- 0x1D00
    x"88",x"88",x"98",x"01",x"90",x"0E",x"00",x"70", -- 0x1D08
    x"00",x"68",x"00",x"00",x"02",x"00",x"01",x"27", -- 0x1D10
    x"09",x"00",x"05",x"04",x"0B",x"09",x"06",x"05", -- 0x1D18
    x"02",x"0B",x"09",x"0A",x"05",x"08",x"0B",x"09", -- 0x1D20
    x"14",x"05",x"02",x"0B",x"09",x"18",x"05",x"02", -- 0x1D28
    x"0B",x"09",x"1A",x"07",x"02",x"0B",x"09",x"02", -- 0x1D30
    x"08",x"02",x"0B",x"09",x"06",x"08",x"02",x"0B", -- 0x1D38
    x"09",x"0A",x"08",x"08",x"58",x"0F",x"14",x"09", -- 0x1D40
    x"02",x"0B",x"09",x"18",x"09",x"02",x"0B",x"09", -- 0x1D48
    x"00",x"0A",x"02",x"0B",x"09",x"02",x"0C",x"02", -- 0x1D50
    x"0B",x"09",x"06",x"0C",x"02",x"0B",x"09",x"0A", -- 0x1D58
    x"0C",x"08",x"0B",x"09",x"14",x"0C",x"02",x"0B", -- 0x1D60
    x"09",x"18",x"0C",x"02",x"0B",x"09",x"1A",x"0D", -- 0x1D68
    x"02",x"0B",x"09",x"00",x"0F",x"1C",x"0B",x"09", -- 0x1D70
    x"00",x"00",x"00",x"00",x"33",x"01",x"00",x"3A", -- 0x1D78
    x"01",x"06",x"57",x"41",x"43",x"4B",x"59",x"20", -- 0x1D80
    x"41",x"4D",x"4F",x"45",x"42",x"41",x"54",x"52", -- 0x1D88
    x"4F",x"4E",x"53",x"00",x"0A",x"08",x"08",x"58", -- 0x1D90
    x"0F",x"01",x"00",x"0D",x"01",x"45",x"1B",x"10", -- 0x1D98
    x"01",x"24",x"C0",x"58",x"18",x"58",x"58",x"80", -- 0x1DA0
    x"01",x"C0",x"58",x"50",x"58",x"58",x"80",x"01", -- 0x1DA8
    x"B0",x"04",x"08",x"20",x"04",x"68",x"01",x"B0", -- 0x1DB0
    x"08",x"08",x"40",x"04",x"68",x"02",x"B0",x"12", -- 0x1DB8
    x"08",x"90",x"04",x"68",x"01",x"B0",x"16",x"08", -- 0x1DC0
    x"B0",x"04",x"68",x"02",x"00",x"0C",x"00",x"03", -- 0x1DC8
    x"0E",x"0F",x"0F",x"00",x"8C",x"28",x"09",x"14", -- 0x1DD0
    x"00",x"08",x"0E",x"0F",x"00",x"02",x"06",x"0E", -- 0x1DD8
    x"0F",x"1A",x"02",x"02",x"0E",x"0F",x"10",x"04", -- 0x1DE0
    x"04",x"0E",x"0F",x"07",x"05",x"01",x"0E",x"0F", -- 0x1DE8
    x"08",x"05",x"07",x"78",x"01",x"16",x"05",x"06", -- 0x1DF0
    x"0E",x"0F",x"00",x"06",x"04",x"0E",x"0F",x"10", -- 0x1DF8
    x"07",x"07",x"0E",x"0F",x"17",x"07",x"03",x"78", -- 0x1E00
    x"01",x"00",x"08",x"05",x"0E",x"0F",x"08",x"09", -- 0x1E08
    x"07",x"0E",x"0F",x"1A",x"09",x"02",x"0E",x"0F", -- 0x1E10
    x"00",x"0A",x"04",x"0E",x"0F",x"04",x"0A",x"02", -- 0x1E18
    x"78",x"01",x"10",x"0A",x"07",x"0E",x"0F",x"17", -- 0x1E20
    x"0B",x"03",x"78",x"01",x"07",x"0C",x"0A",x"13", -- 0x1E28
    x"05",x"00",x"0D",x"03",x"0E",x"0F",x"19",x"0D", -- 0x1E30
    x"03",x"0E",x"0F",x"00",x"0F",x"1C",x"13",x"05", -- 0x1E38
    x"0B",x"0D",x"00",x"08",x"37",x"0F",x"0A",x"00", -- 0x1E40
    x"11",x"00",x"13",x"00",x"14",x"01",x"02",x"03", -- 0x1E48
    x"00",x"09",x"1B",x"0A",x"16",x"0B",x"00",x"3B", -- 0x1E50
    x"01",x"05",x"54",x"48",x"45",x"20",x"45",x"4E", -- 0x1E58
    x"44",x"4F",x"52",x"49",x"41",x"4E",x"20",x"46", -- 0x1E60
    x"4F",x"52",x"45",x"53",x"54",x"00",x"02",x"0D", -- 0x1E68
    x"00",x"58",x"0F",x"00",x"00",x"04",x"05",x"45", -- 0x1E70
    x"1B",x"0D",x"01",x"1B",x"01",x"14",x"02",x"0B", -- 0x1E78
    x"06",x"11",x"08",x"40",x"D0",x"40",x"38",x"40", -- 0x1E80
    x"40",x"68",x"01",x"D0",x"38",x"50",x"38",x"38", -- 0x1E88
    x"68",x"01",x"D0",x"18",x"68",x"18",x"18",x"B8", -- 0x1E90
    x"01",x"D0",x"80",x"28",x"80",x"80",x"A0",x"01", -- 0x1E98
    x"00",x"00",x"00",x"06",x"2A",x"07",x"00",x"03", -- 0x1EA0
    x"04",x"0F",x"01",x"04",x"05",x"06",x"0F",x"01", -- 0x1EA8
    x"0E",x"05",x"02",x"0F",x"01",x"10",x"05",x"05", -- 0x1EB0
    x"14",x"05",x"15",x"05",x"02",x"0F",x"01",x"1A", -- 0x1EB8
    x"06",x"02",x"0F",x"01",x"00",x"08",x"02",x"0F", -- 0x1EC0
    x"01",x"04",x"08",x"02",x"80",x"09",x"1A",x"08", -- 0x1EC8
    x"02",x"0F",x"01",x"0A",x"09",x"07",x"0F",x"01", -- 0x1ED0
    x"19",x"0A",x"01",x"0F",x"01",x"05",x"0B",x"03", -- 0x1ED8
    x"80",x"10",x"08",x"0B",x"01",x"0F",x"01",x"19", -- 0x1EE0
    x"0C",x"03",x"0F",x"01",x"00",x"0D",x"02",x"0F", -- 0x1EE8
    x"01",x"14",x"0D",x"03",x"0F",x"01",x"00",x"0F", -- 0x1EF0
    x"1C",x"0F",x"0F",x"00",x"01",x"00",x"04",x"1A", -- 0x1EF8
    x"09",x"10",x"01",x"15",x"09",x"10",x"0B",x"0B", -- 0x1F00
    x"0C",x"07",x"1B",x"01",x"10",x"00",x"15",x"06", -- 0x1F08
    x"15",x"07",x"15",x"08",x"0B",x"0A",x"0B",x"0B", -- 0x1F10
    x"10",x"0A",x"01",x"41",x"54",x"54",x"41",x"43", -- 0x1F18
    x"4B",x"20",x"4F",x"46",x"20",x"54",x"48",x"45", -- 0x1F20
    x"20",x"4D",x"55",x"54",x"41",x"4E",x"54",x"20", -- 0x1F28
    x"50",x"48",x"4F",x"4E",x"45",x"53",x"00",x"04", -- 0x1F30
    x"08",x"02",x"50",x"09",x"00",x"02",x"01",x"05", -- 0x1F38
    x"45",x"1B",x"15",x"00",x"1B",x"01",x"00",x"04", -- 0x1F40
    x"11",x"06",x"1B",x"0D",x"24",x"F0",x"70",x"18", -- 0x1F48
    x"70",x"70",x"A8",x"01",x"F0",x"20",x"68",x"20", -- 0x1F50
    x"20",x"90",x"01",x"E0",x"02",x"20",x"10",x"20", -- 0x1F58
    x"68",x"02",x"E0",x"0B",x"02",x"58",x"02",x"38", -- 0x1F60
    x"01",x"E0",x"12",x"30",x"90",x"30",x"68",x"01", -- 0x1F68
    x"E0",x"17",x"02",x"B8",x"02",x"68",x"FD",x"00", -- 0x1F70
    x"05",x"00",x"01",x"46",x"07",x"10",x"00",x"01", -- 0x1F78
    x"25",x"07",x"11",x"00",x"01",x"46",x"07",x"14", -- 0x1F80
    x"00",x"01",x"25",x"07",x"0E",x"02",x"02",x"80", -- 0x1F88
    x"01",x"00",x"05",x"03",x"08",x"01",x"08",x"05", -- 0x1F90
    x"05",x"80",x"01",x"0D",x"05",x"85",x"25",x"07", -- 0x1F98
    x"10",x"05",x"8B",x"25",x"07",x"11",x"05",x"04", -- 0x1FA0
    x"80",x"01",x"15",x"05",x"02",x"08",x"01",x"1B", -- 0x1FA8
    x"06",x"01",x"08",x"01",x"05",x"07",x"02",x"08", -- 0x1FB0
    x"01",x"02",x"08",x"01",x"08",x"01",x"16",x"08", -- 0x1FB8
    x"06",x"08",x"0F",x"09",x"09",x"04",x"08",x"01", -- 0x1FC0
    x"05",x"0A",x"01",x"08",x"01",x"11",x"0A",x"03", -- 0x1FC8
    x"08",x"01",x"16",x"0B",x"02",x"08",x"01",x"00", -- 0x1FD0
    x"0C",x"06",x"08",x"01",x"0A",x"0D",x"03",x"08", -- 0x1FD8
    x"01",x"0D",x"0D",x"83",x"25",x"07",x"11",x"0D", -- 0x1FE0
    x"08",x"50",x"09",x"00",x"0F",x"0D",x"08",x"01", -- 0x1FE8
    x"0D",x"0F",x"03",x"08",x"01",x"11",x"0F",x"0B", -- 0x1FF0
    x"08",x"01",x"0E",x"0D",x"00",x"02",x"30",x"0F", -- 0x1FF8
    x"14",x"0C",x"19",x"0C",x"02",x"3C",x"05",x"01", -- 0x2000
    x"00",x"09",x"00",x"00",x"52",x"45",x"54",x"55", -- 0x2008
    x"52",x"4E",x"20",x"4F",x"46",x"20",x"41",x"4C", -- 0x2010
    x"49",x"45",x"4E",x"20",x"4B",x"4F",x"4E",x"47", -- 0x2018
    x"20",x"42",x"45",x"41",x"53",x"54",x"00",x"11", -- 0x2020
    x"0D",x"09",x"50",x"09",x"01",x"00",x"0D",x"05", -- 0x2028
    x"45",x"1B",x"0E",x"03",x"17",x"05",x"01",x"06", -- 0x2030
    x"0F",x"07",x"1A",x"0D",x"31",x"A0",x"40",x"68", -- 0x2038
    x"40",x"00",x"40",x"FF",x"A0",x"50",x"58",x"50", -- 0x2040
    x"50",x"70",x"01",x"A0",x"B0",x"30",x"B0",x"B0", -- 0x2048
    x"C8",x"01",x"90",x"0E",x"00",x"70",x"00",x"70", -- 0x2050
    x"00",x"00",x"00",x"00",x"1C",x"27",x"09",x"02", -- 0x2058
    x"01",x"8E",x"16",x"09",x"06",x"03",x"12",x"05", -- 0x2060
    x"05",x"1A",x"03",x"02",x"05",x"05",x"06",x"06", -- 0x2068
    x"02",x"05",x"05",x"0A",x"06",x"04",x"05",x"05", -- 0x2070
    x"10",x"06",x"05",x"05",x"05",x"17",x"06",x"02", -- 0x2078
    x"05",x"05",x"1B",x"06",x"01",x"05",x"05",x"06", -- 0x2080
    x"09",x"05",x"05",x"05",x"0D",x"09",x"03",x"05", -- 0x2088
    x"05",x"13",x"09",x"03",x"05",x"05",x"18",x"09", -- 0x2090
    x"04",x"05",x"05",x"06",x"0C",x"03",x"05",x"05", -- 0x2098
    x"0B",x"0C",x"03",x"05",x"05",x"10",x"0C",x"04", -- 0x20A0
    x"05",x"05",x"16",x"0C",x"02",x"05",x"05",x"1A", -- 0x20A8
    x"0C",x"02",x"05",x"05",x"00",x"0F",x"02",x"05", -- 0x20B0
    x"05",x"02",x"0F",x"18",x"58",x"0F",x"1A",x"0F", -- 0x20B8
    x"02",x"05",x"05",x"00",x"0D",x"00",x"00",x"33", -- 0x20C0
    x"01",x"00",x"3A",x"01",x"08",x"4F",x"52",x"45", -- 0x20C8
    x"20",x"52",x"45",x"46",x"49",x"4E",x"45",x"52", -- 0x20D0
    x"59",x"00",x"02",x"0F",x"18",x"58",x"0F",x"01", -- 0x20D8
    x"1A",x"0D",x"05",x"45",x"1B",x"18",x"03",x"09", -- 0x20E0
    x"06",x"12",x"09",x"17",x"09",x"0A",x"0C",x"41", -- 0x20E8
    x"C0",x"30",x"08",x"30",x"30",x"D0",x"02",x"C0", -- 0x20F0
    x"80",x"20",x"80",x"30",x"D0",x"01",x"C0",x"88", -- 0x20F8
    x"38",x"88",x"30",x"D0",x"FE",x"C0",x"98",x"50", -- 0x2100
    x"98",x"30",x"D0",x"01",x"B0",x"04",x"38",x"20", -- 0x2108
    x"08",x"68",x"02",x"01",x"0E",x"05",x"01",x"06", -- 0x2110
    x"05",x"0F",x"05",x"01",x"07",x"05",x"02",x"06", -- 0x2118
    x"01",x"06",x"05",x"03",x"06",x"01",x"07",x"05", -- 0x2120
    x"0A",x"06",x"01",x"06",x"05",x"0B",x"06",x"01", -- 0x2128
    x"07",x"05",x"12",x"06",x"01",x"06",x"05",x"13", -- 0x2130
    x"06",x"01",x"07",x"05",x"1A",x"06",x"01",x"06", -- 0x2138
    x"05",x"1B",x"06",x"01",x"07",x"05",x"06",x"07", -- 0x2140
    x"01",x"06",x"05",x"07",x"07",x"01",x"07",x"05", -- 0x2148
    x"16",x"07",x"01",x"06",x"05",x"17",x"07",x"01", -- 0x2150
    x"07",x"05",x"04",x"09",x"01",x"06",x"05",x"05", -- 0x2158
    x"09",x"01",x"07",x"05",x"0C",x"09",x"01",x"06", -- 0x2160
    x"05",x"0D",x"09",x"01",x"07",x"05",x"14",x"09", -- 0x2168
    x"01",x"06",x"05",x"15",x"09",x"01",x"07",x"05", -- 0x2170
    x"1A",x"09",x"01",x"06",x"05",x"1B",x"09",x"01", -- 0x2178
    x"07",x"05",x"00",x"0B",x"01",x"06",x"05",x"01", -- 0x2180
    x"0B",x"01",x"07",x"05",x"08",x"0B",x"01",x"06", -- 0x2188
    x"05",x"09",x"0B",x"01",x"07",x"05",x"0E",x"0B", -- 0x2190
    x"06",x"58",x"0F",x"18",x"0B",x"01",x"06",x"05", -- 0x2198
    x"19",x"0B",x"01",x"07",x"05",x"06",x"0D",x"01", -- 0x21A0
    x"06",x"05",x"07",x"0D",x"01",x"07",x"05",x"00", -- 0x21A8
    x"0F",x"1C",x"29",x"05",x"0E",x"00",x"00",x"00", -- 0x21B0
    x"33",x"01",x"00",x"3A",x"01",x"05",x"53",x"4B", -- 0x21B8
    x"59",x"4C",x"41",x"42",x"20",x"4C",x"41",x"4E", -- 0x21C0
    x"44",x"49",x"4E",x"47",x"20",x"42",x"41",x"59", -- 0x21C8
    x"00",x"0E",x"0B",x"06",x"58",x"0F",x"00",x"1A", -- 0x21D0
    x"0D",x"04",x"44",x"01",x"16",x"02",x"0F",x"07", -- 0x21D8
    x"1A",x"07",x"02",x"08",x"03",x"E0",x"00",x"20", -- 0x21E0
    x"00",x"00",x"48",x"04",x"E0",x"0A",x"00",x"50", -- 0x21E8
    x"00",x"20",x"01",x"E0",x"14",x"10",x"A0",x"00", -- 0x21F0
    x"38",x"03",x"00",x"04",x"00",x"18",x"2A",x"07", -- 0x21F8
    x"1A",x"01",x"8E",x"15",x"07",x"1B",x"01",x"8E", -- 0x2200
    x"15",x"07",x"06",x"03",x"0F",x"50",x"05",x"15", -- 0x2208
    x"03",x"05",x"0F",x"01",x"06",x"04",x"01",x"1B", -- 0x2210
    x"01",x"06",x"05",x"01",x"1A",x"09",x"19",x"04", -- 0x2218
    x"86",x"1B",x"01",x"19",x"0A",x"01",x"1A",x"09", -- 0x2220
    x"00",x"05",x"04",x"0F",x"01",x"15",x"06",x"02", -- 0x2228
    x"0F",x"01",x"05",x"07",x"01",x"80",x"10",x"0A", -- 0x2230
    x"07",x"02",x"0F",x"01",x"02",x"08",x"02",x"0F", -- 0x2238
    x"01",x"10",x"08",x"02",x"0F",x"01",x"16",x"09", -- 0x2240
    x"02",x"0F",x"01",x"00",x"0A",x"02",x"0F",x"01", -- 0x2248
    x"0A",x"0A",x"02",x"0F",x"01",x"10",x"0B",x"02", -- 0x2250
    x"0F",x"01",x"04",x"0C",x"02",x"0F",x"01",x"15", -- 0x2258
    x"0C",x"02",x"0F",x"01",x"0A",x"0D",x"02",x"0F", -- 0x2260
    x"01",x"00",x"0F",x"1C",x"0F",x"01",x"00",x"03", -- 0x2268
    x"00",x"00",x"33",x"01",x"00",x"3A",x"01",x"0A", -- 0x2270
    x"54",x"48",x"45",x"20",x"42",x"41",x"4E",x"4B", -- 0x2278
    x"00",x"06",x"03",x"0F",x"50",x"05",x"00",x"01", -- 0x2280
    x"0D",x"03",x"45",x"1B",x"16",x"02",x"0A",x"06", -- 0x2288
    x"18",x"0E",x"13",x"C0",x"78",x"68",x"78",x"78", -- 0x2290
    x"88",x"01",x"E0",x"07",x"28",x"38",x"24",x"68", -- 0x2298
    x"02",x"E0",x"0D",x"40",x"68",x"24",x"68",x"01", -- 0x22A0
    x"E0",x"12",x"50",x"90",x"20",x"68",x"FD",x"00", -- 0x22A8
    x"00",x"05",x"01",x"08",x"01",x"05",x"05",x"01", -- 0x22B0
    x"08",x"01",x"14",x"05",x"02",x"08",x"01",x"03", -- 0x22B8
    x"07",x"01",x"08",x"01",x"16",x"07",x"06",x"08", -- 0x22C0
    x"01",x"0A",x"05",x"84",x"2B",x"17",x"0D",x"05", -- 0x22C8
    x"84",x"2B",x"17",x"0E",x"06",x"83",x"2B",x"17", -- 0x22D0
    x"0F",x"07",x"82",x"2B",x"17",x"10",x"08",x"81", -- 0x22D8
    x"2B",x"17",x"00",x"09",x"02",x"80",x"01",x"02", -- 0x22E0
    x"09",x"18",x"50",x"09",x"09",x"0B",x"02",x"2B", -- 0x22E8
    x"17",x"0B",x"0B",x"02",x"08",x"01",x"0B",x"0B", -- 0x22F0
    x"02",x"08",x"01",x"19",x"0B",x"01",x"08",x"01", -- 0x22F8
    x"00",x"0C",x"09",x"08",x"01",x"13",x"0D",x"01", -- 0x2300
    x"08",x"01",x"19",x"0D",x"01",x"08",x"01",x"16", -- 0x2308
    x"0E",x"03",x"36",x"0F",x"00",x"0F",x"1C",x"08", -- 0x2310
    x"01",x"0B",x"05",x"00",x"00",x"33",x"01",x"00", -- 0x2318
    x"3A",x"01",x"04",x"54",x"48",x"45",x"20",x"53", -- 0x2320
    x"49",x"58",x"54",x"45",x"45",x"4E",x"54",x"48", -- 0x2328
    x"20",x"43",x"41",x"56",x"45",x"52",x"4E",x"00", -- 0x2330
    x"02",x"09",x"18",x"50",x"09",x"00",x"01",x"0D", -- 0x2338
    x"04",x"45",x"1B",x"00",x"00",x"1B",x"02",x"0C", -- 0x2340
    x"07",x"10",x"0A",x"40",x"20",x"B0",x"28",x"B0", -- 0x2348
    x"B0",x"D0",x"01",x"20",x"88",x"38",x"88",x"88", -- 0x2350
    x"A0",x"01",x"20",x"10",x"50",x"10",x"02",x"38", -- 0x2358
    x"01",x"20",x"50",x"68",x"50",x"02",x"88",x"01", -- 0x2360
    x"00",x"00",x"05",x"1C",x"90",x"05",x"00",x"06", -- 0x2368
    x"1C",x"90",x"05",x"00",x"07",x"1C",x"90",x"05", -- 0x2370
    x"00",x"08",x"1C",x"90",x"05",x"00",x"09",x"1C", -- 0x2378
    x"90",x"05",x"00",x"0A",x"1C",x"90",x"05",x"00", -- 0x2380
    x"0B",x"1C",x"90",x"05",x"00",x"0C",x"1C",x"90", -- 0x2388
    x"05",x"02",x"08",x"85",x"00",x"00",x"03",x"08", -- 0x2390
    x"85",x"00",x"00",x"08",x"05",x"88",x"00",x"00", -- 0x2398
    x"09",x"05",x"88",x"00",x"00",x"11",x"05",x"85", -- 0x23A0
    x"00",x"00",x"12",x"05",x"85",x"00",x"00",x"18", -- 0x23A8
    x"05",x"88",x"00",x"00",x"19",x"05",x"88",x"00", -- 0x23B0
    x"00",x"0C",x"08",x"05",x"58",x"0F",x"00",x"05", -- 0x23B8
    x"02",x"11",x"05",x"1A",x"05",x"02",x"11",x"05", -- 0x23C0
    x"18",x"0E",x"04",x"11",x"05",x"00",x"0F",x"1C", -- 0x23C8
    x"11",x"05",x"1A",x"01",x"00",x"06",x"32",x"07", -- 0x23D0
    x"05",x"04",x"07",x"04",x"0B",x"04",x"0E",x"04", -- 0x23D8
    x"14",x"04",x"16",x"04",x"04",x"3E",x"05",x"02", -- 0x23E0
    x"06",x"17",x"07",x"14",x"0A",x"07",x"0B",x"08", -- 0x23E8
    x"54",x"48",x"45",x"20",x"57",x"41",x"52",x"45", -- 0x23F0
    x"48",x"4F",x"55",x"53",x"45",x"00",x"0C",x"08", -- 0x23F8
    x"05",x"58",x"0F",x"01",x"00",x"03",x"05",x"45", -- 0x2400
    x"1B",x"16",x"05",x"0D",x"07",x"00",x"09",x"11", -- 0x2408
    x"0A",x"17",x"0B",x"24",x"70",x"20",x"68",x"20", -- 0x2410
    x"20",x"30",x"01",x"70",x"50",x"68",x"50",x"50", -- 0x2418
    x"B0",x"01",x"40",x"02",x"40",x"10",x"40",x"68", -- 0x2420
    x"02",x"40",x"08",x"40",x"40",x"00",x"68",x"FD", -- 0x2428
    x"40",x"11",x"30",x"88",x"00",x"40",x"01",x"40", -- 0x2430
    x"18",x"00",x"C0",x"00",x"60",x"04",x"00",x"19", -- 0x2438
    x"00",x"01",x"2D",x"09",x"02",x"05",x"1A",x"08", -- 0x2440
    x"01",x"00",x"07",x"02",x"08",x"01",x"0B",x"08", -- 0x2448
    x"11",x"08",x"01",x"02",x"09",x"07",x"08",x"01", -- 0x2450
    x"1B",x"0A",x"01",x"08",x"01",x"02",x"0C",x"1A", -- 0x2458
    x"08",x"01",x"00",x"0D",x"02",x"08",x"01",x"04", -- 0x2460
    x"05",x"88",x"00",x"00",x"05",x"05",x"88",x"00", -- 0x2468
    x"00",x"09",x"05",x"88",x"00",x"00",x"0A",x"05", -- 0x2470
    x"88",x"00",x"00",x"13",x"05",x"88",x"00",x"00", -- 0x2478
    x"14",x"05",x"88",x"00",x"00",x"18",x"05",x"88", -- 0x2480
    x"00",x"00",x"19",x"05",x"88",x"00",x"00",x"00", -- 0x2488
    x"0F",x"1C",x"08",x"01",x"1A",x"00",x"00",x"00", -- 0x2490
    x"34",x"01",x"00",x"3B",x"01",x"04",x"4F",x"4D", -- 0x2498
    x"4F",x"45",x"42",x"41",x"54",x"52",x"4F",x"4E", -- 0x24A0
    x"53",x"27",x"20",x"52",x"45",x"56",x"45",x"4E", -- 0x24A8
    x"47",x"45",x"00",x"02",x"0D",x"00",x"58",x"0F", -- 0x24B0
    x"00",x"1A",x"0D",x"01",x"45",x"1B",x"0F",x"01", -- 0x24B8
    x"34",x"C0",x"58",x"30",x"58",x"58",x"88",x"02", -- 0x24C0
    x"C0",x"78",x"50",x"78",x"58",x"88",x"01",x"C0", -- 0x24C8
    x"70",x"68",x"70",x"58",x"88",x"FE",x"B0",x"04", -- 0x24D0
    x"68",x"20",x"05",x"68",x"FC",x"B0",x"09",x"48", -- 0x24D8
    x"48",x"05",x"68",x"02",x"B0",x"13",x"48",x"98", -- 0x24E0
    x"05",x"68",x"04",x"B0",x"18",x"28",x"C0",x"05", -- 0x24E8
    x"68",x"01",x"0F",x"00",x"00",x"02",x"20",x"09", -- 0x24F0
    x"02",x"05",x"01",x"12",x"15",x"07",x"05",x"06", -- 0x24F8
    x"12",x"15",x"15",x"05",x"07",x"12",x"15",x"11", -- 0x2500
    x"07",x"02",x"12",x"15",x"00",x"08",x"01",x"12", -- 0x2508
    x"15",x"0B",x"08",x"03",x"12",x"15",x"15",x"08", -- 0x2510
    x"07",x"12",x"15",x"11",x"0A",x"01",x"12",x"15", -- 0x2518
    x"00",x"0B",x"03",x"12",x"15",x"0C",x"0C",x"05", -- 0x2520
    x"12",x"15",x"15",x"0B",x"07",x"12",x"15",x"00", -- 0x2528
    x"0E",x"02",x"20",x"09",x"00",x"0F",x"02",x"20", -- 0x2530
    x"09",x"02",x"0F",x"1A",x"12",x"15",x"14",x"0F", -- 0x2538
    x"01",x"20",x"09",x"00",x"01",x"00",x"00",x"33", -- 0x2540
    x"01",x"00",x"3A",x"01",x"04",x"53",x"4F",x"4C", -- 0x2548
    x"41",x"52",x"20",x"50",x"4F",x"57",x"45",x"52", -- 0x2550
    x"20",x"47",x"45",x"4E",x"45",x"52",x"41",x"54", -- 0x2558
    x"4F",x"52",x"00",x"05",x"0C",x"04",x"58",x"0F", -- 0x2560
    x"00",x"0C",x"0A",x"03",x"44",x"0F",x"1B",x"01", -- 0x2568
    x"00",x"05",x"1B",x"0C",x"43",x"70",x"B8",x"18", -- 0x2570
    x"B8",x"A0",x"D0",x"02",x"70",x"D0",x"30",x"D0", -- 0x2578
    x"98",x"D0",x"FE",x"70",x"C8",x"48",x"C8",x"98", -- 0x2580
    x"D0",x"FF",x"70",x"78",x"68",x"78",x"60",x"D0", -- 0x2588
    x"02",x"E0",x"03",x"58",x"18",x"04",x"68",x"03", -- 0x2590
    x"E0",x"09",x"38",x"48",x"30",x"68",x"FE",x"E0", -- 0x2598
    x"0E",x"48",x"70",x"02",x"50",x"FF",x"00",x"00", -- 0x25A0
    x"00",x"05",x"03",x"0F",x"00",x"01",x"05",x"03", -- 0x25A8
    x"0F",x"00",x"02",x"04",x"03",x"0F",x"02",x"02", -- 0x25B0
    x"84",x"28",x"09",x"05",x"00",x"17",x"01",x"01", -- 0x25B8
    x"05",x"01",x"17",x"01",x"01",x"04",x"02",x"18", -- 0x25C0
    x"01",x"01",x"17",x"02",x"05",x"04",x"01",x"17", -- 0x25C8
    x"03",x"05",x"04",x"01",x"00",x"03",x"83",x"01", -- 0x25D0
    x"01",x"01",x"03",x"83",x"01",x"01",x"03",x"03", -- 0x25D8
    x"0C",x"01",x"01",x"03",x"04",x"03",x"01",x"01", -- 0x25E0
    x"06",x"04",x"01",x"3F",x"09",x"05",x"05",x"01", -- 0x25E8
    x"3F",x"09",x"07",x"04",x"02",x"2E",x"09",x"06", -- 0x25F0
    x"05",x"04",x"2E",x"09",x"09",x"04",x"01",x"1F", -- 0x25F8
    x"09",x"0A",x"05",x"01",x"1F",x"09",x"13",x"00", -- 0x2600
    x"01",x"3F",x"09",x"14",x"00",x"02",x"2E",x"09", -- 0x2608
    x"16",x"00",x"01",x"1F",x"09",x"13",x"01",x"82", -- 0x2610
    x"2E",x"0F",x"14",x"01",x"82",x"1E",x"01",x"15", -- 0x2618
    x"01",x"82",x"1E",x"01",x"16",x"01",x"82",x"2E", -- 0x2620
    x"0F",x"13",x"03",x"04",x"2E",x"0F",x"0A",x"04", -- 0x2628
    x"03",x"01",x"01",x"03",x"05",x"02",x"01",x"01", -- 0x2630
    x"0B",x"05",x"01",x"01",x"01",x"1A",x"08",x"02", -- 0x2638
    x"08",x"01",x"18",x"0A",x"01",x"80",x"01",x"19", -- 0x2640
    x"0B",x"01",x"08",x"01",x"00",x"0C",x"01",x"08", -- 0x2648
    x"01",x"03",x"0D",x"01",x"08",x"01",x"00",x"0F", -- 0x2650
    x"1C",x"08",x"01",x"0F",x"04",x"0D",x"24",x"15", -- 0x2658
    x"0D",x"05",x"03",x"24",x"15",x"12",x"05",x"83", -- 0x2660
    x"24",x"15",x"0D",x"06",x"03",x"24",x"15",x"00", -- 0x2668
    x"06",x"04",x"24",x"15",x"00",x"07",x"10",x"24", -- 0x2670
    x"15",x"04",x"06",x"03",x"03",x"0F",x"07",x"06", -- 0x2678
    x"02",x"01",x"01",x"09",x"06",x"04",x"03",x"0F", -- 0x2680
    x"0C",x"05",x"01",x"03",x"0F",x"10",x"05",x"00", -- 0x2688
    x"06",x"31",x"05",x"0D",x"04",x"0E",x"04",x"0F", -- 0x2690
    x"03",x"10",x"03",x"11",x"03",x"12",x"03",x"04", -- 0x2698
    x"1A",x"05",x"06",x"0B",x"09",x"0B",x"0E",x"0B", -- 0x26A0
    x"12",x"0B",x"06",x"54",x"48",x"45",x"20",x"46", -- 0x26A8
    x"49",x"4E",x"41",x"4C",x"20",x"42",x"41",x"52", -- 0x26B0
    x"52",x"49",x"45",x"52",x"00",x"00",x"0A",x"14", -- 0x26B8
    x"58",x"0F",x"01",x"19",x"0D",x"05",x"45",x"1B", -- 0x26C0
    x"14",x"05",x"1B",x"06",x"07",x"0B",x"0B",x"0B", -- 0x26C8
    x"10",x"0B",x"11",x"70",x"38",x"68",x"38",x"20", -- 0x26D0
    x"98",x"02",x"E0",x"15",x"30",x"A8",x"28",x"68", -- 0x26D8
    x"01",x"00",x"21",x"07",x"27",x"16",x"16",x"0E", -- 0x26E0
    x"0A",x"1E",x"00",x"06",x"1C",x"7E",x"23",x"E5", -- 0x26E8
    x"D5",x"F5",x"CD",x"6D",x"0B",x"F1",x"C6",x"80", -- 0x26F0
    x"77",x"CB",x"D4",x"36",x"1B",x"D1",x"E1",x"1C", -- 0x26F8
    x"10",x"EB",x"14",x"0D",x"20",x"E3",x"C9",x"20", -- 0x2700
    x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20", -- 0x2708
    x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20", -- 0x2710
    x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20", -- 0x2718
    x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"50", -- 0x2720
    x"41",x"43",x"2D",x"4D",x"41",x"4E",x"49",x"43", -- 0x2728
    x"2D",x"4D",x"49",x"4E",x"45",x"52",x"2D",x"4D", -- 0x2730
    x"41",x"4E",x"20",x"20",x"20",x"20",x"20",x"20", -- 0x2738
    x"57",x"52",x"49",x"54",x"54",x"45",x"4E",x"20", -- 0x2740
    x"42",x"59",x"20",x"4A",x"49",x"4D",x"20",x"42", -- 0x2748
    x"41",x"47",x"4C",x"45",x"59",x"20",x"46",x"4F", -- 0x2750
    x"52",x"20",x"20",x"20",x"20",x"50",x"41",x"43", -- 0x2758
    x"4D",x"41",x"4E",x"20",x"41",x"52",x"43",x"41", -- 0x2760
    x"44",x"45",x"20",x"48",x"41",x"52",x"44",x"57", -- 0x2768
    x"41",x"52",x"45",x"2E",x"20",x"20",x"20",x"20", -- 0x2770
    x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20", -- 0x2778
    x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20", -- 0x2780
    x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20", -- 0x2788
    x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20", -- 0x2790
    x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20", -- 0x2798
    x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20", -- 0x27A0
    x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20", -- 0x27A8
    x"20",x"20",x"4A",x"55",x"4D",x"50",x"20",x"3D", -- 0x27B0
    x"20",x"4A",x"4F",x"59",x"20",x"32",x"20",x"2D", -- 0x27B8
    x"3E",x"20",x"52",x"49",x"47",x"48",x"54",x"20", -- 0x27C0
    x"20",x"20",x"20",x"20",x"4D",x"55",x"53",x"49", -- 0x27C8
    x"43",x"20",x"4F",x"4E",x"2F",x"4F",x"46",x"46", -- 0x27D0
    x"20",x"3D",x"20",x"4A",x"4F",x"59",x"20",x"32", -- 0x27D8
    x"20",x"2D",x"3E",x"20",x"55",x"50",x"20",x"20", -- 0x27E0
    x"46",x"58",x"20",x"4F",x"4E",x"2F",x"4F",x"46", -- 0x27E8
    x"46",x"20",x"3D",x"20",x"4A",x"4F",x"59",x"20", -- 0x27F0
    x"32",x"20",x"2D",x"3E",x"20",x"44",x"4F",x"57", -- 0x27F8
    x"4E",x"2E",x"20",x"20",x"20",x"20",x"20",x"20", -- 0x2800
    x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20", -- 0x2808
    x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20", -- 0x2810
    x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"41", -- 0x2818
    x"49",x"52",x"20",x"E7",x"E7",x"E7",x"E7",x"E7", -- 0x2820
    x"E7",x"00",x"E7",x"E7",x"E7",x"E7",x"E7",x"E7", -- 0x2828
    x"E7",x"E7",x"E7",x"E7",x"E7",x"E7",x"E7",x"E7", -- 0x2830
    x"E7",x"E7",x"E7",x"E7",x"00",x"48",x"49",x"53", -- 0x2838
    x"43",x"4F",x"52",x"45",x"20",x"00",x"20",x"20", -- 0x2840
    x"53",x"43",x"4F",x"52",x"45",x"20",x"00",x"00", -- 0x2848
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2850
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2858
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2860
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2868
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2870
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2878
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2880
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2888
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2890
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2898
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x28A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x28A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x28B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x28B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x28C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x28C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x28D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x28D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x28E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x28E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x28F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x28F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2900
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2908
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2910
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2918
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2920
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2928
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2930
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2938
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2940
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2948
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2950
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2958
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2960
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2968
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2970
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2978
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2980
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2988
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2990
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2998
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x29A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x29A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x29B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x29B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x29C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x29C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x29D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x29D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x29E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x29E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x29F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x29F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A08
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A10
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A18
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A28
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A30
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A38
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A40
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A48
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A50
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A58
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A60
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A68
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A78
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A80
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A88
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A90
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2AA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2AA8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2AB0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2AB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2AC0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2AC8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2AD0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2AD8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2AE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2AE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2AF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2AF8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B08
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B10
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B18
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B28
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B30
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B38
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B40
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B48
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B50
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B58
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B60
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B68
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B78
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B80
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B88
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B90
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2BA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2BA8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2BB0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2BB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2BC0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2BC8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2BD0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2BD8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2BE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2BE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2BF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2BF8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C08
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C10
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C18
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C28
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C30
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C38
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C40
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C48
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C50
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C58
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C60
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C68
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C78
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C80
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C88
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C90
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2CA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2CA8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2CB0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2CB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2CC0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2CC8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2CD0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2CD8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2CE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2CE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2CF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2CF8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D08
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D10
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D18
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D28
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D30
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D38
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D40
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D48
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D50
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D58
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D60
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D68
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D78
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D80
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D88
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D90
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2DA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2DA8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2DB0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2DB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2DC0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2DC8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2DD0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2DD8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2DE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2DE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2DF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2DF8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E08
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E10
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E18
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E28
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E30
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E38
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E40
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E48
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E50
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E58
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E60
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E68
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E78
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E80
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E88
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E90
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2EA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2EA8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2EB0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2EB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2EC0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2EC8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2ED0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2ED8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2EE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2EE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2EF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2EF8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F08
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F10
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F18
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F28
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F30
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F38
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F40
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F48
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F50
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F58
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F60
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F68
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F78
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F80
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F88
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F90
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2FA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2FA8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2FB0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2FB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2FC0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2FC8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2FD0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2FD8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2FE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2FE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2FF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2FF8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3000
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3008
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3010
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3018
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3020
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3028
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3030
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3038
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3040
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3048
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3050
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3058
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3060
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3068
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3070
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3078
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3080
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3088
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3090
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3098
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x30A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x30A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x30B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x30B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x30C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x30C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x30D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x30D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x30E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x30E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x30F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x30F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3100
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3108
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3110
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3118
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3120
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3128
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3130
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3138
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3140
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3148
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3150
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3158
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3160
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3168
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3170
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3178
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3180
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3188
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3190
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3198
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3200
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3208
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3210
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3218
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3220
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3228
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3230
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3238
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3240
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3248
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3250
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3258
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3260
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3268
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3270
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3278
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3280
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3288
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3290
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3298
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x32A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x32A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x32B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x32B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x32C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x32C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x32D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x32D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x32E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x32E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x32F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x32F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3300
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3308
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3310
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3318
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3320
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3328
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3330
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3338
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3340
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3348
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3350
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3358
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3360
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3368
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3370
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3378
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3380
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3388
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3390
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3398
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x33A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x33A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x33B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x33B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x33C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x33C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x33D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x33D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x33E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x33E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x33F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x33F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3400
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3408
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3410
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3418
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3420
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3428
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3430
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3438
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3440
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3448
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3450
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3458
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3460
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3468
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3470
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3478
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3480
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3488
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3490
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3498
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3500
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3508
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3510
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3518
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3520
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3528
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3530
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3538
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3540
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3548
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3550
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3558
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3560
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3568
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3570
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3578
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3580
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3588
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3590
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3598
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3600
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3608
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3610
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3618
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3620
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3628
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3630
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3638
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3640
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3648
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3650
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3658
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3660
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3668
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3670
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3678
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3680
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3688
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3690
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3698
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3700
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3708
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3710
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3718
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3720
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3728
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3730
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3738
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3740
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3748
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3750
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3758
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3760
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3768
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3770
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3778
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3780
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3788
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3790
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3798
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3800
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3808
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3810
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3818
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3820
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3828
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3830
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3838
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3840
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3848
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3850
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3858
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3860
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3868
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3870
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3878
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3880
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3888
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3890
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3898
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x38A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x38A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x38B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x38B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x38C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x38C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x38D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x38D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x38E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x38E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x38F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x38F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3900
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3908
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3910
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3918
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3920
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3928
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3930
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3938
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3940
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3948
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3950
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3958
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3960
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3968
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3970
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3978
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3980
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3988
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3990
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3998
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A08
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A10
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A18
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A28
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A30
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A38
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A40
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A48
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A50
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A58
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A60
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A68
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A78
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A80
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A88
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A90
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3AA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3AA8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3AB0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3AB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3AC0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3AC8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3AD0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3AD8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3AE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3AE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3AF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3AF8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B08
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B10
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B18
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B28
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B30
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B38
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B40
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B48
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B50
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B58
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B60
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B68
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B78
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B80
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B88
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B90
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3BA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3BA8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3BB0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3BB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3BC0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3BC8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3BD0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3BD8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3BE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3BE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3BF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3BF8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C08
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C10
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C18
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C28
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C30
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C38
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C40
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C48
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C50
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C58
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C60
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C68
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C78
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C80
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C88
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C90
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3CA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3CA8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3CB0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3CB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3CC0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3CC8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3CD0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3CD8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3CE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3CE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3CF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3CF8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D08
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D10
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D18
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D28
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D30
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D38
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D40
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D48
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D50
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D58
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D60
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D68
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D78
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D80
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D88
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D90
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3DA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3DA8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3DB0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3DB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3DC0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3DC8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3DD0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3DD8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3DE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3DE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3DF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3DF8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E08
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E10
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E18
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E28
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E30
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E38
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E40
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E48
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E50
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E58
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E60
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E68
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E78
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E80
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E88
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E90
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3EA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3EA8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3EB0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3EB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3EC0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3EC8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3ED0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3ED8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3EE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3EE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3EF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3EF8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F08
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F10
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F18
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F28
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F30
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F38
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F40
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F48
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F50
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F58
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F60
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F68
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F78
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F80
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F88
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F90
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3FA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3FA8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3FB0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3FB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3FC0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3FC8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3FD0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3FD8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3FE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3FE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3FF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"  -- 0x3FF8
  );

begin

  p_rom : process
  begin
    wait until rising_edge(CLK);
       DATA <= ROM(to_integer(unsigned(ADDR)));
  end process;
end RTL;
