library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity timber_bg_bits_1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of timber_bg_bits_1 is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"55",X"84",X"15",X"4A",X"A5",X"46",X"91",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"A9",X"AA",X"A9",X"AA",X"A9",X"AA",X"A9",X"AA",X"A9",X"AA",X"A9",
		X"97",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"56",X"55",X"56",X"55",X"56",X"55",X"56",X"57",X"56",X"55",X"56",X"55",X"56",X"55",X"56",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AB",
		X"AB",X"FD",X"AD",X"55",X"AD",X"45",X"B5",X"55",X"B5",X"55",X"D4",X"55",X"D5",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"7F",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AB",X"AA",X"AD",X"AA",X"AD",X"AA",X"B5",X"AA",X"B5",X"AA",X"D4",X"AA",X"D5",X"AB",X"55",
		X"55",X"55",X"45",X"55",X"5D",X"55",X"5F",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"75",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AB",X"55",X"AD",X"45",X"AD",X"55",X"B5",X"55",X"B5",X"55",X"D4",X"55",X"D5",X"55",X"D5",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"D5",X"55",X"54",X"55",X"55",X"55",X"55",
		X"57",X"55",X"17",X"15",X"5D",X"5D",X"5D",X"55",X"75",X"55",X"74",X"55",X"D5",X"55",X"D5",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"D5",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0B",X"80",X"02",X"C0",X"A2",X"28",X"2E",X"E0",X"0A",X"B0",X"3E",X"FC",X"FF",X"FF",X"3F",X"F0",
		X"00",X"00",X"00",X"00",X"02",X"00",X"22",X"EA",X"0A",X"AF",X"3F",X"BF",X"03",X"FC",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AB",X"AA",X"AB",X"AA",X"AD",X"AA",X"AD",
		X"BF",X"FF",X"D5",X"55",X"D4",X"55",X"D5",X"55",X"55",X"55",X"51",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"75",X"55",X"74",X"55",X"D5",X"55",X"D5",X"55",X"51",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"55",X"55",X"55",X"51",X"7D",X"55",X"55",X"55",X"55",X"47",X"55",X"57",X"55",X"55",
		X"FF",X"FF",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"75",X"55",X"75",X"15",X"D5",X"55",X"D5",X"55",X"55",X"55",X"45",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"51",X"55",X"55",X"55",X"55",X"55",X"57",X"55",X"17",X"55",X"5D",X"55",X"55",
		X"55",X"55",X"15",X"55",X"55",X"55",X"55",X"F5",X"55",X"F5",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AD",X"AA",X"B5",X"AA",X"B5",X"AA",X"D5",X"AA",X"D4",X"AA",X"D5",X"AB",X"55",X"AB",X"55",
		X"AD",X"55",X"AD",X"45",X"AD",X"55",X"B5",X"55",X"B5",X"15",X"D5",X"55",X"D5",X"55",X"D5",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"40",X"80",X"00",X"06",X"90",X"01",X"40",X"01",X"40",X"04",X"10",X"14",X"14",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"D5",X"51",X"D5",X"57",X"51",X"57",X"55",X"5D",X"55",X"5D",X"15",X"35",X"55",X"75",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"57",X"55",X"47",X"55",X"57",X"55",X"57",X"55",X"57",X"55",X"47",X"55",X"57",X"55",X"57",
		X"55",X"55",X"55",X"55",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"55",X"55",X"55",X"55",
		X"55",X"55",X"FF",X"FF",X"FF",X"FF",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"FF",X"FF",X"FF",X"FF",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"7D",X"55",X"55",
		X"55",X"55",X"FF",X"FF",X"FF",X"FF",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"D5",X"55",
		X"55",X"55",X"FF",X"FF",X"FF",X"FF",X"55",X"55",X"75",X"55",X"55",X"55",X"55",X"75",X"55",X"55",
		X"55",X"55",X"7F",X"FD",X"FF",X"FF",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"AA",X"BF",X"AA",X"FF",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"95",
		X"AA",X"95",X"AA",X"95",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"F6",X"55",X"00",X"15",
		X"55",X"55",X"55",X"55",X"55",X"7F",X"55",X"7D",X"55",X"7F",X"55",X"55",X"55",X"5F",X"55",X"5F",
		X"55",X"55",X"55",X"55",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"A9",X"55",X"69",X"55",X"A9",X"55",X"F5",X"55",X"A5",X"55",X"A5",X"55",
		X"55",X"55",X"55",X"55",X"56",X"AA",X"56",X"AA",X"56",X"9A",X"56",X"AA",X"54",X"01",X"55",X"A9",
		X"55",X"A9",X"55",X"A9",X"55",X"A9",X"55",X"A9",X"55",X"A9",X"55",X"A9",X"55",X"A9",X"55",X"A9",
		X"A5",X"55",X"A5",X"55",X"A5",X"55",X"A5",X"D5",X"A5",X"55",X"A5",X"55",X"A5",X"55",X"A5",X"55",
		X"55",X"5F",X"55",X"5F",X"55",X"5F",X"55",X"5F",X"55",X"5F",X"55",X"5F",X"55",X"5F",X"55",X"5F",
		X"00",X"15",X"00",X"15",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"15",
		X"00",X"15",X"00",X"15",X"00",X"55",X"00",X"55",X"80",X"55",X"20",X"55",X"E4",X"55",X"A8",X"15",
		X"55",X"A9",X"55",X"A9",X"55",X"A9",X"5D",X"A9",X"55",X"A1",X"55",X"80",X"55",X"91",X"55",X"95",
		X"55",X"95",X"55",X"95",X"55",X"B9",X"57",X"A9",X"7A",X"81",X"A8",X"05",X"80",X"94",X"05",X"94",
		X"55",X"55",X"57",X"55",X"57",X"55",X"57",X"55",X"FF",X"55",X"AA",X"55",X"AA",X"55",X"00",X"55",
		X"55",X"95",X"55",X"95",X"55",X"95",X"55",X"95",X"55",X"95",X"55",X"95",X"55",X"B9",X"5F",X"A9",
		X"57",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",X"00",X"00",
		X"55",X"41",X"55",X"00",X"75",X"41",X"55",X"55",X"FF",X"55",X"AA",X"55",X"AA",X"55",X"00",X"55",
		X"55",X"55",X"55",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"5F",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",X"00",X"00",
		X"88",X"01",X"C8",X"00",X"24",X"41",X"84",X"55",X"84",X"55",X"AA",X"55",X"AA",X"55",X"00",X"55",
		X"EB",X"55",X"89",X"55",X"28",X"55",X"B0",X"55",X"2A",X"55",X"8A",X"55",X"82",X"55",X"AA",X"55",
		X"62",X"AA",X"63",X"8F",X"E6",X"AA",X"88",X"8A",X"89",X"2E",X"98",X"6A",X"82",X"A3",X"8A",X"FA",
		X"28",X"AA",X"A8",X"AE",X"A2",X"8A",X"AA",X"48",X"69",X"E9",X"AA",X"AA",X"AA",X"AA",X"00",X"00",
		X"A7",X"20",X"92",X"A8",X"68",X"8A",X"AA",X"A0",X"4A",X"9A",X"20",X"8E",X"A9",X"A8",X"AC",X"69",
		X"02",X"00",X"82",X"00",X"08",X"20",X"28",X"80",X"B6",X"C0",X"A0",X"88",X"2A",X"A8",X"A8",X"AC",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FA",X"AA",X"0F",X"EA",X"00",X"0F",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"7B",X"55",X"0A",X"55",X"8A",X"55",X"A4",X"55",X"2B",X"55",X"10",X"55",X"82",X"55",X"88",X"55",
		X"A2",X"82",X"A6",X"00",X"2A",X"41",X"6A",X"55",X"FF",X"55",X"AA",X"55",X"AA",X"55",X"00",X"55",
		X"AA",X"A6",X"2A",X"2A",X"82",X"02",X"A1",X"28",X"85",X"A8",X"9A",X"AA",X"BC",X"94",X"AA",X"2A",
		X"08",X"33",X"08",X"B0",X"02",X"26",X"20",X"24",X"09",X"1A",X"2A",X"28",X"A2",X"8A",X"0A",X"8A",
		X"AA",X"AA",X"AA",X"AA",X"FE",X"AA",X"03",X"FE",X"00",X"03",X"00",X"00",X"00",X"20",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"00",X"F0",X"00",X"F0",X"02",X"FC",X"0A",X"FF",X"02",X"FF",X"C2",X"FF",X"8A",X"FE",X"0A",
		X"FF",X"A6",X"FF",X"C9",X"EA",X"08",X"82",X"A3",X"9A",X"94",X"26",X"6A",X"91",X"88",X"69",X"2A",
		X"B2",X"CA",X"A2",X"29",X"AB",X"89",X"8A",X"AC",X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",X"00",X"00",
		X"D0",X"A9",X"B8",X"82",X"26",X"0B",X"08",X"A2",X"A2",X"A6",X"8A",X"02",X"B9",X"25",X"82",X"6B",
		X"E8",X"55",X"AE",X"55",X"22",X"55",X"FC",X"55",X"B1",X"55",X"B4",X"55",X"82",X"55",X"8A",X"55",
		X"3E",X"82",X"FE",X"00",X"FC",X"41",X"FA",X"55",X"FF",X"55",X"AA",X"55",X"AA",X"55",X"00",X"55",
		X"00",X"3F",X"00",X"3F",X"00",X"FF",X"00",X"FA",X"03",X"E2",X"0F",X"FA",X"0F",X"F8",X"0F",X"82",
		X"0F",X"FF",X"03",X"FF",X"00",X"FF",X"00",X"3F",X"00",X"3F",X"00",X"0F",X"00",X"0F",X"00",X"0F",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"BF",X"FF",X"C0",X"00",X"00",X"FF",X"00",X"FF",X"F0",X"FF",X"FC",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AF",X"7F",X"F0",X"FF",X"FF",X"00",X"3F",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"55",X"AA",X"55",X"55",X"55",X"7F",X"7F",X"C0",X"C0",X"00",
		X"55",X"55",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",X"00",X"00",
		X"00",X"FF",X"03",X"FF",X"0F",X"FF",X"3F",X"FE",X"FF",X"FF",X"FF",X"FE",X"FF",X"FA",X"FF",X"FE",
		X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",
		X"00",X"00",X"00",X"00",X"00",X"41",X"00",X"55",X"FF",X"55",X"AA",X"55",X"AA",X"55",X"00",X"55",
		X"AA",X"AA",X"5A",X"AA",X"55",X"56",X"55",X"55",X"55",X"55",X"D5",X"55",X"FF",X"55",X"FF",X"FF",
		X"F5",X"6A",X"7F",X"55",X"57",X"D5",X"55",X"F5",X"55",X"7D",X"95",X"5F",X"55",X"57",X"55",X"55",
		X"55",X"55",X"55",X"57",X"95",X"FC",X"BF",X"00",X"A0",X"00",X"A0",X"00",X"20",X"00",X"00",X"00",
		X"7F",X"F0",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",X"00",X"00",
		X"28",X"00",X"8A",X"00",X"A2",X"41",X"88",X"55",X"FF",X"55",X"AA",X"55",X"AA",X"55",X"00",X"55",
		X"A0",X"55",X"88",X"55",X"8A",X"55",X"AA",X"55",X"28",X"55",X"8A",X"55",X"94",X"55",X"8A",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A2",X"AA",X"2C",X"28",X"80",X"8B",X"5A",X"82",X"02",X"2A",X"48",X"88",X"A8",X"A2",X"2A",X"2A",
		X"9A",X"22",X"8A",X"B0",X"08",X"82",X"AA",X"A8",X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",X"00",X"00",
		X"A9",X"AA",X"8A",X"22",X"05",X"8A",X"AA",X"AA",X"BC",X"9A",X"A2",X"A2",X"22",X"8A",X"A8",X"2A",
		X"80",X"00",X"A0",X"00",X"28",X"00",X"88",X"00",X"02",X"00",X"2B",X"00",X"80",X"00",X"A8",X"00",
		X"B3",X"21",X"AF",X"88",X"AA",X"A2",X"AA",X"28",X"A2",X"E2",X"68",X"0A",X"04",X"8A",X"A6",X"A0",
		X"AC",X"89",X"20",X"A5",X"80",X"25",X"28",X"99",X"2B",X"0A",X"8A",X"AA",X"22",X"05",X"82",X"85",
		X"88",X"AA",X"29",X"AA",X"02",X"2A",X"A8",X"AA",X"02",X"2A",X"AA",X"AA",X"EA",X"2A",X"8B",X"0A",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"0A",X"AA",X"A2",X"AA",X"2A",X"AA",
		X"55",X"55",X"56",X"95",X"56",X"95",X"55",X"55",X"55",X"55",X"56",X"95",X"56",X"95",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"55",X"55",X"56",X"A6",X"55",X"96",X"55",X"96",X"55",X"96",X"55",X"96",X"55",X"55",
		X"AA",X"AA",X"55",X"55",X"96",X"9A",X"66",X"59",X"96",X"9A",X"66",X"59",X"66",X"9A",X"55",X"55",
		X"AA",X"AA",X"55",X"55",X"5A",X"55",X"65",X"55",X"59",X"55",X"56",X"55",X"6A",X"55",X"55",X"55",
		X"AA",X"AA",X"55",X"55",X"65",X"A6",X"65",X"96",X"65",X"A6",X"65",X"96",X"69",X"A6",X"55",X"55",
		X"AA",X"AA",X"55",X"55",X"9A",X"95",X"56",X"55",X"96",X"55",X"56",X"55",X"56",X"55",X"55",X"55",
		X"AA",X"AA",X"55",X"55",X"55",X"6A",X"55",X"59",X"55",X"59",X"55",X"59",X"55",X"59",X"55",X"55",
		X"AA",X"AA",X"55",X"55",X"66",X"9A",X"66",X"AA",X"66",X"66",X"66",X"56",X"66",X"56",X"55",X"55",
		X"AA",X"AA",X"55",X"55",X"69",X"55",X"65",X"55",X"69",X"55",X"65",X"55",X"69",X"55",X"55",X"55",
		X"AA",X"AA",X"55",X"55",X"96",X"9A",X"96",X"59",X"96",X"9A",X"96",X"59",X"A6",X"99",X"55",X"55",
		X"AA",X"AA",X"55",X"55",X"6A",X"55",X"59",X"55",X"59",X"55",X"59",X"55",X"59",X"55",X"55",X"55",
		X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"8C",X"A2",X"7B",X"AB",X"3F",X"FF",X"FF",X"FF",
		X"FE",X"55",X"AA",X"55",X"AA",X"55",X"00",X"55",X"88",X"55",X"A2",X"55",X"EB",X"55",X"FF",X"D7",
		X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"55",X"AA",X"55",X"AA",X"55",X"00",X"55",X"3F",X"55",X"FF",X"55",X"FF",X"55",X"FF",X"D7",
		X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"55",X"AA",X"55",X"AA",X"55",X"00",X"55",X"AA",X"55",X"FA",X"55",X"FF",X"55",X"FF",X"D7",
		X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"2A",X"AA",X"AA",X"6A",X"FF",X"AB",X"FF",X"FF",
		X"FF",X"55",X"AA",X"55",X"AA",X"55",X"00",X"55",X"AB",X"55",X"FF",X"55",X"FF",X"55",X"FF",X"D7",
		X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"A6",X"EA",X"EB",X"FA",X"FF",X"0F",X"FF",X"FF",
		X"F5",X"55",X"AA",X"55",X"AA",X"55",X"00",X"55",X"AB",X"55",X"AF",X"55",X"FF",X"55",X"FF",X"D7",
		X"55",X"55",X"45",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"45",X"55",X"55",X"55",
		X"55",X"55",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"55",X"AA",X"55",X"AA",X"55",X"00",X"55",X"00",X"55",X"FF",X"55",X"FF",X"55",X"FF",X"D7",
		X"55",X"55",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"55",X"AA",X"55",X"AA",X"55",X"00",X"55",X"00",X"55",X"FF",X"55",X"FF",X"55",X"FF",X"D7",
		X"7A",X"81",X"A8",X"05",X"80",X"F7",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",
		X"55",X"41",X"55",X"01",X"55",X"45",X"55",X"55",X"7F",X"55",X"AA",X"55",X"AA",X"55",X"00",X"55",
		X"55",X"55",X"AA",X"57",X"AA",X"57",X"00",X"57",X"00",X"57",X"FF",X"57",X"FF",X"57",X"FF",X"DF",
		X"55",X"55",X"55",X"55",X"55",X"44",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"A9",X"55",X"A9",X"55",X"A9",X"55",X"A9",X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",X"00",X"00",
		X"55",X"01",X"55",X"A9",X"55",X"A9",X"55",X"A9",X"55",X"A9",X"55",X"A9",X"55",X"A9",X"55",X"55",
		X"55",X"55",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"A9",X"55",X"A9",X"55",X"A9",X"5D",X"A9",X"55",X"A9",X"55",X"A9",X"55",X"A9",X"55",X"A9",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"0F",X"00",X"3F",X"00",X"FF",
		X"FF",X"FF",X"00",X"FF",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FC",X"FF",X"F0",X"FF",X"F0",X"FF",X"C0",X"FF",X"C0",X"FF",X"C0",X"FF",X"00",X"FF",X"C0",
		X"FF",X"00",X"FC",X"00",X"FC",X"00",X"FC",X"00",X"F0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"03",X"FF",X"0F",X"FF",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"3F",X"00",X"FF",X"03",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FF",X"F0",X"FF",X"F0",X"FF",X"F0",X"FF",X"C0",
		X"55",X"5F",X"55",X"5F",X"55",X"55",X"55",X"7F",X"55",X"7D",X"55",X"7F",X"55",X"5F",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"55",X"55",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FC",X"00",X"FC",X"00",X"FC",X"00",X"F0",X"00",X"C0",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FF",X"FF",X"55",X"55",
		X"A5",X"55",X"A5",X"55",X"F5",X"55",X"A9",X"55",X"69",X"55",X"A9",X"55",X"F5",X"55",X"55",X"55",
		X"F5",X"55",X"FD",X"55",X"FD",X"55",X"FD",X"55",X"FD",X"55",X"FD",X"55",X"FD",X"69",X"FD",X"AA",
		X"00",X"03",X"00",X"0F",X"00",X"37",X"00",X"D7",X"03",X"57",X"03",X"57",X"03",X"57",X"0D",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",
		X"C0",X"00",X"70",X"00",X"70",X"00",X"5C",X"00",X"57",X"00",X"55",X"C0",X"55",X"70",X"55",X"5C",
		X"C0",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0D",X"55",X"0D",X"55",X"0D",X"55",X"03",X"55",X"03",X"55",X"03",X"55",X"03",X"55",X"00",X"D5",
		X"00",X"00",X"00",X"3F",X"03",X"F5",X"0F",X"55",X"0D",X"55",X"3D",X"55",X"35",X"55",X"35",X"55",
		X"FF",X"FF",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"D5",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FF",X"FC",X"FF",X"F0",X"FF",X"F0",X"FF",X"00",
		X"FC",X"00",X"FC",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"F0",X"FF",X"F0",X"FF",X"C0",X"FF",X"C0",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FC",X"00",
		X"F5",X"69",X"FD",X"55",X"5F",X"55",X"FF",X"55",X"7F",X"55",X"FF",X"55",X"FD",X"55",X"57",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",
		X"F0",X"00",X"F0",X"00",X"F0",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"FF",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"57",X"55",X"57",X"55",X"57",X"55",X"57",X"55",X"57",X"55",X"57",X"55",X"57",X"55",X"57",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"57",X"55",X"57",X"55",X"57",X"55",X"57",X"55",X"57",X"55",X"57",X"55",X"57",X"55",X"57",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"2A",X"80",X"A0",X"AA",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"0A",
		X"00",X"00",X"00",X"00",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"02",
		X"00",X"00",X"0A",X"A0",X"A8",X"28",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"02",
		X"00",X"00",X"2A",X"AA",X"A0",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",
		X"00",X"00",X"0A",X"AA",X"A0",X"00",X"00",X"00",X"00",X"00",X"2A",X"00",X"02",X"00",X"02",X"00",
		X"00",X"00",X"AA",X"80",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0A",X"AA",X"28",X"00",X"20",X"00",X"20",X"00",X"28",X"00",X"0A",X"00",X"02",X"00",
		X"00",X"00",X"A8",X"0A",X"0A",X"28",X"02",X"A0",X"00",X"00",X"02",X"80",X"00",X"A0",X"00",X"28",
		X"00",X"00",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",
		X"00",X"00",X"A0",X"00",X"2A",X"00",X"02",X"80",X"00",X"A0",X"00",X"28",X"80",X"08",X"A0",X"0A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"2A",X"AA",X"A0",X"00",X"80",X"00",X"80",X"00",X"80",X"00",
		X"00",X"00",X"00",X"02",X"00",X"02",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"A0",X"2A",X"28",X"A0",X"08",X"00",X"00",X"00",X"02",X"00",X"02",X"00",X"02",X"00",
		X"00",X"00",X"A8",X"00",X"0A",X"A8",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"00",X"25",X"00",X"25",X"00",X"25",X"00",X"25",X"00",X"25",X"00",X"25",
		X"02",X"15",X"02",X"55",X"02",X"55",X"02",X"55",X"02",X"15",X"82",X"85",X"80",X"81",X"80",X"80",
		X"00",X"00",X"0A",X"A0",X"09",X"58",X"09",X"58",X"09",X"56",X"09",X"55",X"09",X"55",X"09",X"55",
		X"00",X"00",X"00",X"00",X"94",X"00",X"94",X"00",X"94",X"00",X"94",X"00",X"94",X"00",X"84",X"00",
		X"60",X"02",X"68",X"02",X"58",X"02",X"58",X"00",X"58",X"00",X"58",X"00",X"58",X"00",X"18",X"00",
		X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"10",X"00",X"00",
		X"04",X"08",X"05",X"18",X"05",X"58",X"05",X"58",X"05",X"58",X"04",X"58",X"00",X"18",X"00",X"08",
		X"06",X"00",X"16",X"00",X"16",X"00",X"1A",X"00",X"18",X"00",X"08",X"00",X"08",X"00",X"28",X"00",
		X"00",X"40",X"00",X"50",X"00",X"50",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"80",X"05",X"80",X"55",X"80",X"55",X"80",X"55",X"80",X"41",X"80",X"42",X"80",X"02",X"00",
		X"80",X"00",X"A0",X"00",X"60",X"01",X"60",X"01",X"60",X"01",X"60",X"01",X"60",X"01",X"60",X"01",
		X"28",X"00",X"58",X"00",X"5A",X"01",X"56",X"01",X"56",X"81",X"55",X"81",X"55",X"A1",X"55",X"61",
		X"80",X"00",X"80",X"01",X"80",X"01",X"80",X"01",X"80",X"01",X"80",X"01",X"80",X"01",X"80",X"01",
		X"80",X"00",X"80",X"15",X"80",X"15",X"80",X"55",X"80",X"55",X"81",X"55",X"81",X"55",X"85",X"55",
		X"55",X"40",X"55",X"00",X"55",X"00",X"54",X"00",X"54",X"00",X"50",X"00",X"50",X"00",X"40",X"00",
		X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",
		X"15",X"54",X"05",X"54",X"05",X"54",X"01",X"54",X"01",X"54",X"00",X"54",X"00",X"54",X"00",X"14",
		X"60",X"01",X"20",X"00",X"20",X"00",X"20",X"00",X"20",X"00",X"20",X"00",X"20",X"00",X"20",X"00",
		X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"0A",X"00",X"08",X"00",X"08",X"00",X"08",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",
		X"20",X"00",X"20",X"00",X"20",X"00",X"A0",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"00",X"00",
		X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"08",
		X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",
		X"18",X"00",X"28",X"00",X"20",X"00",X"A0",X"00",X"80",X"00",X"00",X"00",X"00",X"02",X"00",X"02",
		X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"00",X"00",
		X"09",X"55",X"08",X"05",X"08",X"05",X"08",X"01",X"08",X"28",X"08",X"2A",X"08",X"22",X"08",X"22",
		X"60",X"80",X"60",X"80",X"58",X"80",X"55",X"00",X"55",X"40",X"55",X"40",X"55",X"40",X"15",X"40",
		X"00",X"25",X"00",X"20",X"00",X"20",X"00",X"20",X"00",X"20",X"00",X"20",X"00",X"20",X"00",X"20",
		X"00",X"20",X"00",X"20",X"00",X"20",X"00",X"20",X"00",X"20",X"00",X"20",X"00",X"20",X"00",X"08",
		X"95",X"40",X"85",X"40",X"80",X"00",X"A0",X"00",X"20",X"00",X"20",X"00",X"28",X"00",X"08",X"00",
		X"08",X"A2",X"02",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"80",X"00",X"A0",X"00",X"20",X"00",
		X"00",X"0A",X"00",X"08",X"80",X"08",X"A0",X"0A",X"60",X"02",X"68",X"00",X"58",X"00",X"5A",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",
		X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",
		X"08",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"28",X"00",X"20",X"00",
		X"20",X"00",X"20",X"00",X"20",X"00",X"20",X"00",X"20",X"00",X"20",X"00",X"20",X"00",X"20",X"00",
		X"20",X"00",X"20",X"00",X"20",X"00",X"A0",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",
		X"60",X"00",X"60",X"00",X"68",X"00",X"58",X"00",X"5A",X"00",X"56",X"00",X"56",X"00",X"16",X"80",
		X"00",X"60",X"00",X"60",X"00",X"60",X"01",X"60",X"01",X"60",X"05",X"60",X"05",X"60",X"05",X"20",
		X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"08",
		X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",
		X"56",X"00",X"56",X"00",X"56",X"00",X"56",X"00",X"56",X"00",X"16",X"00",X"1A",X"00",X"08",X"00",
		X"20",X"00",X"28",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"09",X"50",X"09",X"55",X"09",X"55",X"09",X"55",X"09",X"55",X"08",X"15",X"08",X"05",X"08",X"00",
		X"08",X"00",X"0A",X"00",X"42",X"00",X"50",X"00",X"50",X"00",X"54",X"00",X"54",X"A0",X"54",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"28",X"00",X"24",
		X"00",X"25",X"00",X"25",X"00",X"25",X"00",X"25",X"00",X"25",X"00",X"25",X"00",X"21",X"00",X"20",
		X"16",X"88",X"02",X"08",X"02",X"08",X"02",X"08",X"0A",X"08",X"08",X"08",X"A8",X"08",X"00",X"08",
		X"08",X"00",X"08",X"00",X"08",X"00",X"0A",X"00",X"02",X"A0",X"00",X"2A",X"00",X"02",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"50",X"00",X"40",X"00",X"54",X"00",X"55",X"40",
		X"A8",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"05",X"01",X"55",X"05",X"55",X"55",X"55",
		X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"50",X"55",X"50",X"55",X"54",X"55",X"55",
		X"00",X"28",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"05",X"05",X"45",X"55",X"45",X"55",X"55",
		X"15",X"20",X"15",X"20",X"14",X"A0",X"52",X"80",X"52",X"00",X"5A",X"00",X"68",X"15",X"40",X"15",
		X"15",X"80",X"15",X"80",X"05",X"A0",X"05",X"60",X"01",X"68",X"01",X"59",X"01",X"55",X"00",X"55",
		X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"02",
		X"20",X"00",X"20",X"00",X"A0",X"00",X"80",X"02",X"80",X"00",X"80",X"00",X"80",X"00",X"00",X"00",
		X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"00",X"05",X"00",X"15",X"41",X"55",X"55",X"55",
		X"00",X"55",X"00",X"55",X"00",X"15",X"00",X"15",X"00",X"04",X"00",X"00",X"00",X"00",X"40",X"00",
		X"40",X"15",X"40",X"55",X"01",X"55",X"01",X"55",X"05",X"55",X"15",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"51",X"55",X"50",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"54",X"15",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"54",X"55",X"55",X"05",X"55",X"05",X"55",X"15",X"55",X"01",X"55",X"00",X"15",X"00",X"01",
		X"00",X"00",X"40",X"00",X"55",X"00",X"55",X"50",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"08",X"50",X"04",X"54",X"00",X"55",X"40",
		X"00",X"20",X"00",X"20",X"00",X"20",X"00",X"28",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"08",
		X"00",X"0A",X"00",X"02",X"00",X"02",X"40",X"02",X"50",X"02",X"54",X"02",X"55",X"02",X"55",X"50",
		X"55",X"50",X"55",X"54",X"55",X"54",X"55",X"54",X"05",X"50",X"01",X"54",X"00",X"15",X"00",X"05",
		X"15",X"55",X"00",X"55",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"54",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"50",X"55",X"40",X"14",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"00",X"14",X"00",X"55",X"01",X"55",X"15",X"55",X"55",X"55",X"55",X"55",X"55",X"50",
		X"00",X"0A",X"00",X"08",X"00",X"28",X"00",X"20",X"00",X"A0",X"00",X"80",X"00",X"81",X"00",X"85",
		X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",
		X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"01",
		X"A8",X"05",X"00",X"15",X"00",X"15",X"00",X"55",X"00",X"55",X"00",X"54",X"00",X"50",X"54",X"00",
		X"55",X"40",X"55",X"00",X"54",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"54",X"55",X"55",X"15",X"55",X"05",X"55",X"01",X"55",X"00",X"55",X"00",X"05",X"00",X"01",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"54",X"00",X"50",X"00",X"40",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"05",X"00",X"05",X"00",X"15",X"00",X"15",X"00",X"55",X"01",X"54",X"01",X"54",X"05",X"50",
		X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"0A",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"28",
		X"00",X"20",X"00",X"20",X"00",X"20",X"00",X"20",X"00",X"20",X"00",X"21",X"00",X"15",X"00",X"15",
		X"05",X"50",X"15",X"40",X"15",X"40",X"55",X"00",X"54",X"00",X"54",X"00",X"50",X"00",X"50",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"40",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"14",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"50",X"00",X"50",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"50",X"15",X"54",X"05",X"55",X"01",X"55",X"00",X"55",X"00",X"15",X"00",X"15",X"00",X"05",
		X"80",X"00",X"20",X"00",X"20",X"00",X"20",X"00",X"00",X"00",X"40",X"00",X"40",X"00",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"04",X"00",X"01",X"00",X"01",X"00",X"55",X"00",X"55",X"00",X"15",X"00",X"05",X"00",X"01",
		X"00",X"08",X"00",X"08",X"40",X"0A",X"50",X"02",X"54",X"02",X"55",X"02",X"55",X"40",X"55",X"50",
		X"00",X"80",X"00",X"A0",X"00",X"20",X"00",X"20",X"00",X"20",X"00",X"28",X"00",X"08",X"00",X"08",
		X"80",X"40",X"80",X"50",X"00",X"54",X"00",X"54",X"00",X"00",X"40",X"00",X"40",X"00",X"40",X"10",
		X"08",X"00",X"0A",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"80",X"00",X"80",X"00",X"80",
		X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"40",X"81",X"40",X"81",X"40",
		X"14",X"00",X"14",X"00",X"14",X"00",X"14",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"00",X"00",
		X"80",X"00",X"A0",X"00",X"20",X"00",X"20",X"00",X"20",X"00",X"20",X"00",X"28",X"00",X"08",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"80",X"00",
		X"40",X"29",X"40",X"09",X"40",X"0A",X"40",X"02",X"40",X"02",X"50",X"02",X"50",X"02",X"10",X"00",
		X"00",X"02",X"00",X"02",X"00",X"0A",X"00",X"29",X"00",X"25",X"00",X"25",X"00",X"25",X"00",X"25",
		X"94",X"00",X"54",X"00",X"54",X"00",X"54",X"00",X"50",X"00",X"50",X"00",X"40",X"00",X"40",X"00",
		X"08",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"28",X"00",X"24",X"00",X"A4",X"00",X"94",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"54",X"00",X"54",X"00",X"14",X"00",X"04",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"08",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"80",X"00",X"A0",X"00",X"20",X"00",X"28",X"00",
		X"00",X"0A",X"00",X"02",X"00",X"02",X"40",X"02",X"50",X"00",X"50",X"00",X"50",X"00",X"54",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"A8",X"00",X"0A",X"80",X"00",X"A8",X"00",X"08",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"8A",X"AA",X"4A",X"AA",X"4A",X"AA",X"42",X"A9",X"00",X"A9",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A5",X"AA",X"95",X"62",X"95",X"82",X"5E",X"62",X"97",X"58",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"2A",X"9A",X"2A",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"8A",X"28",X"88",X"08",X"80",X"00",X"A0",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"2A",X"AA",X"2A",X"AA",X"0A",X"AA",X"02",X"AA",X"00",X"A2",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"82",X"AA",X"80",X"AA",X"02",X"AA",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"22",X"2A",X"88",X"9E",X"22",X"6A",X"8A",X"62",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"BA",X"AA",
		X"AA",X"00",X"A9",X"00",X"6A",X"41",X"6A",X"92",X"AA",X"A5",X"A6",X"A5",X"AA",X"A9",X"A9",X"A9",
		X"A5",X"58",X"65",X"56",X"95",X"68",X"65",X"58",X"55",X"56",X"57",X"56",X"55",X"95",X"D5",X"56",
		X"0A",X"AA",X"02",X"6A",X"02",X"AA",X"0A",X"96",X"09",X"AA",X"06",X"AA",X"8A",X"A9",X"4A",X"AA",
		X"A0",X"00",X"A0",X"00",X"A8",X"00",X"88",X"00",X"A8",X"00",X"AA",X"00",X"AA",X"80",X"2A",X"00",
		X"00",X"2A",X"00",X"2A",X"00",X"28",X"00",X"0A",X"00",X"02",X"00",X"0A",X"00",X"0A",X"00",X"08",
		X"28",X"00",X"A8",X"02",X"A0",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"AA",X"20",X"2B",X"80",X"6A",X"81",X"A8",X"0A",X"AB",X"26",X"8A",X"0A",X"AE",X"0A",X"8B",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"AA",X"A0",X"BA",X"80",X"A8",X"00",X"2A",X"00",X"AA",X"80",
		X"AA",X"AA",X"A9",X"6A",X"29",X"AA",X"02",X"A8",X"02",X"AA",X"00",X"A2",X"00",X"2A",X"00",X"9A",
		X"AA",X"AA",X"AA",X"AA",X"8A",X"88",X"2A",X"00",X"A8",X"80",X"A8",X"A0",X"AA",X"A0",X"2A",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"2A",X"AA",X"2A",X"A9",X"0A",X"AA",X"02",X"A2",X"02",X"2A",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A2",X"AA",X"6A",X"A2",X"6A",X"2A",X"6A",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"98",X"A0",X"A4",X"00",X"A4",X"00",X"24",X"00",
		X"AA",X"AA",X"AA",X"AA",X"2A",X"AA",X"0A",X"AA",X"00",X"99",X"00",X"25",X"00",X"25",X"00",X"24",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"6A",X"AA",X"60",X"2A",X"60",X"28",X"18",X"08",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"8A",X"2A",X"09",X"08",X"02",X"00",X"02",X"00",X"02",
		X"00",X"01",X"00",X"26",X"00",X"0A",X"00",X"0A",X"00",X"2A",X"00",X"28",X"00",X"2A",X"00",X"1A",
		X"56",X"00",X"41",X"80",X"54",X"60",X"55",X"18",X"45",X"24",X"55",X"90",X"41",X"A0",X"51",X"60",
		X"00",X"67",X"00",X"91",X"02",X"55",X"09",X"35",X"06",X"75",X"01",X"95",X"02",X"51",X"02",X"55",
		X"A8",X"00",X"A9",X"00",X"29",X"00",X"A4",X"00",X"A8",X"00",X"A8",X"00",X"A4",X"00",X"A9",X"00",
		X"6A",X"22",X"AA",X"0A",X"9A",X"AA",X"9A",X"AA",X"A2",X"62",X"A9",X"AA",X"A1",X"A8",X"AA",X"6A",
		X"0A",X"AA",X"02",X"2A",X"00",X"AA",X"00",X"22",X"00",X"2A",X"00",X"28",X"00",X"0A",X"00",X"02",
		X"8A",X"A0",X"A2",X"A8",X"2A",X"A8",X"AA",X"A0",X"A2",X"80",X"AA",X"A0",X"68",X"A8",X"AA",X"A8",
		X"00",X"2A",X"00",X"1A",X"00",X"26",X"00",X"0A",X"00",X"02",X"00",X"01",X"00",X"02",X"00",X"00",
		X"A2",X"80",X"BA",X"60",X"AA",X"A8",X"BA",X"A0",X"A2",X"E0",X"AA",X"A8",X"2A",X"AA",X"AB",X"AC",
		X"0A",X"EA",X"A2",X"AE",X"AA",X"EA",X"BE",X"2A",X"2A",X"AF",X"AA",X"AA",X"BA",X"BE",X"AA",X"E2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"0A",X"00",X"0A",X"00",X"02",X"00",X"02",
		X"00",X"A8",X"0A",X"80",X"2A",X"00",X"2A",X"00",X"22",X"80",X"AA",X"A0",X"8A",X"A0",X"AA",X"A0",
		X"A8",X"00",X"A8",X"00",X"AA",X"00",X"8A",X"80",X"AA",X"00",X"AA",X"00",X"A8",X"82",X"AA",X"A2",
		X"0A",X"6A",X"29",X"A8",X"AA",X"AA",X"6A",X"2A",X"9A",X"9A",X"62",X"AA",X"AA",X"AA",X"6A",X"A6",
		X"55",X"68",X"59",X"56",X"95",X"55",X"65",X"55",X"57",X"55",X"96",X"56",X"5D",X"55",X"55",X"55",
		X"AA",X"A9",X"A9",X"A5",X"AA",X"A5",X"AA",X"96",X"6A",X"A5",X"AA",X"A9",X"6A",X"A5",X"AA",X"95",
		X"A6",X"A5",X"AA",X"A9",X"9A",X"A5",X"6A",X"A5",X"AA",X"A5",X"A6",X"A9",X"A9",X"A9",X"AA",X"A5",
		X"7F",X"FF",X"1F",X"FF",X"07",X"FF",X"55",X"FF",X"55",X"FF",X"FF",X"7F",X"FF",X"7F",X"FF",X"DF",
		X"5A",X"A6",X"5A",X"9A",X"56",X"9A",X"56",X"AA",X"56",X"A9",X"55",X"AA",X"55",X"AA",X"D5",X"6A",
		X"AA",X"A9",X"A6",X"A2",X"6A",X"AA",X"9A",X"A2",X"A9",X"AA",X"AA",X"AA",X"AA",X"2A",X"6A",X"AA",
		X"AA",X"A9",X"6A",X"2A",X"6A",X"AA",X"9A",X"A9",X"A6",X"A0",X"AA",X"A9",X"9A",X"AA",X"6A",X"8A",
		X"00",X"0A",X"40",X"09",X"40",X"0A",X"00",X"0A",X"00",X"02",X"00",X"02",X"40",X"02",X"40",X"0A",
		X"6A",X"AA",X"AE",X"AA",X"AB",X"6A",X"6A",X"AB",X"9E",X"A2",X"6A",X"BA",X"A2",X"AB",X"AB",X"3A",
		X"AA",X"AA",X"E8",X"AA",X"A2",X"8A",X"AA",X"AE",X"B8",X"AA",X"A2",X"A2",X"AB",X"AA",X"2A",X"EA",
		X"00",X"00",X"00",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"00",X"00",X"80",X"00",X"80",X"00",
		X"AA",X"26",X"2A",X"89",X"AA",X"AA",X"AA",X"AA",X"2A",X"AA",X"0A",X"2A",X"2A",X"AA",X"AA",X"AA",
		X"00",X"0A",X"00",X"2A",X"00",X"0A",X"80",X"2A",X"80",X"2A",X"00",X"0A",X"80",X"0A",X"80",X"0A",
		X"2A",X"9A",X"AA",X"6A",X"A1",X"AA",X"AA",X"6A",X"8A",X"98",X"AA",X"66",X"8A",X"9A",X"AA",X"AA",
		X"8A",X"40",X"AA",X"40",X"2A",X"90",X"AA",X"90",X"AA",X"64",X"A2",X"98",X"8A",X"A9",X"AA",X"A6",
		X"01",X"5D",X"01",X"D5",X"00",X"D5",X"00",X"55",X"02",X"7D",X"01",X"5D",X"05",X"D4",X"09",X"75",
		X"55",X"50",X"44",X"90",X"15",X"58",X"50",X"94",X"55",X"49",X"59",X"46",X"55",X"15",X"45",X"15",
		X"00",X"28",X"00",X"6A",X"00",X"92",X"00",X"6A",X"01",X"A8",X"06",X"AA",X"99",X"A2",X"62",X"AA",
		X"80",X"A2",X"82",X"AA",X"8A",X"28",X"6A",X"AA",X"5A",X"A2",X"5A",X"2A",X"6A",X"AA",X"AA",X"A2",
		X"55",X"51",X"55",X"61",X"46",X"54",X"65",X"51",X"55",X"59",X"44",X"45",X"55",X"55",X"11",X"54",
		X"A7",X"56",X"A7",X"45",X"97",X"61",X"95",X"55",X"A5",X"D5",X"9D",X"54",X"95",X"56",X"B5",X"15",
		X"A8",X"AA",X"AA",X"2A",X"AA",X"AA",X"A8",X"A2",X"AA",X"AA",X"6A",X"A2",X"6A",X"2A",X"6A",X"AA",
		X"AA",X"A6",X"A8",X"9A",X"AA",X"9A",X"AA",X"A6",X"8A",X"A9",X"AA",X"AA",X"AA",X"AA",X"8A",X"2A",
		X"00",X"22",X"80",X"2A",X"80",X"22",X"A0",X"0A",X"A8",X"02",X"2A",X"0A",X"AA",X"8A",X"A2",X"8A",
		X"2A",X"A8",X"2A",X"AA",X"0A",X"A2",X"0A",X"A2",X"08",X"AA",X"02",X"AA",X"0A",X"8A",X"0A",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"80",X"00",X"A0",X"00",X"80",X"00",X"80",X"00",
		X"AA",X"2A",X"AA",X"A8",X"A2",X"AA",X"B2",X"8E",X"AA",X"AA",X"2A",X"AA",X"8B",X"A2",X"AA",X"8A",
		X"00",X"1F",X"00",X"1F",X"00",X"07",X"55",X"57",X"55",X"57",X"55",X"57",X"55",X"57",X"FF",X"FD",
		X"40",X"2A",X"90",X"2A",X"24",X"AB",X"A4",X"AA",X"29",X"AA",X"8A",X"6A",X"AA",X"AE",X"8A",X"A8",
		X"AA",X"2A",X"5A",X"AA",X"9A",X"AA",X"6A",X"2A",X"9A",X"AA",X"9A",X"A2",X"A6",X"AA",X"A9",X"AA",
		X"6A",X"A9",X"AA",X"4A",X"AA",X"AA",X"A9",X"AA",X"AA",X"8A",X"9A",X"AA",X"AA",X"26",X"AA",X"AA",
		X"AA",X"99",X"A9",X"A5",X"AA",X"96",X"9A",X"95",X"AA",X"95",X"AA",X"65",X"AA",X"65",X"AA",X"56",
		X"95",X"D9",X"55",X"5D",X"55",X"55",X"57",X"5D",X"55",X"55",X"55",X"DD",X"67",X"55",X"59",X"59",
		X"55",X"5A",X"55",X"5A",X"75",X"56",X"65",X"56",X"65",X"56",X"5D",X"5A",X"55",X"5A",X"D7",X"5A",
		X"AA",X"96",X"AA",X"95",X"AA",X"99",X"F9",X"A5",X"DF",X"D9",X"77",X"7F",X"FF",X"FF",X"AA",X"AE",
		X"55",X"57",X"55",X"5D",X"55",X"55",X"69",X"96",X"65",X"55",X"DA",X"A5",X"FF",X"FF",X"FE",X"AE",
		X"59",X"5A",X"55",X"56",X"65",X"D5",X"57",X"55",X"55",X"55",X"55",X"5A",X"FF",X"F5",X"BF",X"AB",
		X"A6",X"A8",X"AA",X"8A",X"AA",X"AA",X"AA",X"9A",X"A9",X"AA",X"AA",X"BF",X"AF",X"F7",X"AF",X"AA",
		X"6A",X"6A",X"AA",X"9A",X"8A",X"9A",X"AA",X"9A",X"FF",X"FF",X"75",X"FD",X"DF",X"77",X"AA",X"AF",
		X"AA",X"AB",X"A8",X"AA",X"AA",X"22",X"AA",X"8A",X"FF",X"FA",X"F7",X"EA",X"5D",X"7F",X"AF",X"BA",
		X"AB",X"AE",X"AA",X"AA",X"BA",X"8A",X"AA",X"AA",X"AA",X"A8",X"AA",X"AA",X"EE",X"AE",X"FE",X"FE",
		X"AA",X"AA",X"A8",X"AA",X"A8",X"EA",X"2A",X"2A",X"AE",X"A2",X"AA",X"AA",X"AA",X"AE",X"AA",X"FF",
		X"80",X"00",X"80",X"00",X"A0",X"00",X"88",X"00",X"AA",X"00",X"AA",X"03",X"BF",X"FF",X"AA",X"AA",
		X"02",X"A8",X"00",X"AA",X"00",X"8A",X"00",X"2A",X"03",X"FF",X"F7",X"FD",X"DD",X"DF",X"AE",X"BB",
		X"AA",X"6A",X"22",X"AA",X"AA",X"9A",X"AA",X"6A",X"FF",X"D6",X"DF",X"7D",X"DD",X"F7",X"FE",X"AB",
		X"AA",X"8A",X"A8",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"EA",X"AA",X"FA",X"BF",
		X"9A",X"8A",X"9A",X"A9",X"9A",X"AA",X"A6",X"AA",X"9A",X"BF",X"9A",X"FF",X"AF",X"FD",X"AE",X"FE",
		X"55",X"55",X"57",X"55",X"55",X"55",X"B5",X"D4",X"D5",X"55",X"5D",X"75",X"55",X"5D",X"EF",X"FB",
		X"55",X"55",X"59",X"52",X"56",X"65",X"55",X"15",X"54",X"64",X"55",X"59",X"45",X"45",X"FB",X"FA",
		X"68",X"AA",X"6A",X"8A",X"9A",X"AA",X"56",X"AA",X"5A",X"AA",X"1F",X"DE",X"57",X"7F",X"FA",X"FB",
		X"BF",X"FF",X"FF",X"FF",X"FF",X"BF",X"FF",X"FF",X"AA",X"03",X"FF",X"AA",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"AA",X"FF",X"FF",X"AA",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FB",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"AF",X"FF",X"FA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F3",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"AF",
		X"FF",X"FF",X"FF",X"FF",X"FA",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"AF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EB",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"F3",X"FF",X"FF",X"FF",X"FF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FB",X"FE",X"AF",X"FB",X"FF",X"EF",X"FF",X"BF",X"EB",X"BF",X"FF",X"AF",X"FF",X"FA",X"BF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"AF",X"AE",X"BF",X"AA",X"BF",X"AE",X"BF",X"EA",X"AF",
		X"FF",X"FF",X"FF",X"FF",X"AA",X"AF",X"AA",X"AA",X"AA",X"EA",X"EA",X"AE",X"AA",X"AA",X"AB",X"AE",
		X"FF",X"FF",X"AA",X"FF",X"AA",X"AA",X"BA",X"AA",X"AA",X"AB",X"AA",X"EA",X"AA",X"AA",X"BA",X"AE",
		X"AA",X"FF",X"AA",X"AA",X"AA",X"AA",X"AE",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AE",X"BA",X"EA",
		X"AA",X"AA",X"AA",X"EE",X"BA",X"AA",X"AE",X"BA",X"BA",X"EB",X"AA",X"AA",X"BE",X"EE",X"AA",X"AA",
		X"FF",X"FF",X"40",X"00",X"D4",X"00",X"F1",X"55",X"F0",X"55",X"50",X"5F",X"C4",X"1F",X"C1",X"07",
		X"FF",X"FF",X"FD",X"55",X"34",X"57",X"F4",X"57",X"D0",X"55",X"D1",X"17",X"71",X"17",X"74",X"15",
		X"FF",X"EA",X"FF",X"FF",X"AB",X"FF",X"AB",X"FF",X"AE",X"AF",X"AB",X"AA",X"EA",X"BA",X"AA",X"BB",
		X"BF",X"FF",X"EF",X"FF",X"FA",X"BF",X"FF",X"EA",X"FF",X"FF",X"BA",X"BF",X"AA",X"AB",X"AE",X"AA",
		X"FF",X"FF",X"EA",X"FA",X"FF",X"FF",X"AB",X"FF",X"FE",X"AB",X"FF",X"FE",X"FF",X"FF",X"AB",X"FA",
		X"FF",X"FF",X"FF",X"FF",X"FB",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"FF",X"FF",X"FF",
		X"41",X"04",X"10",X"44",X"11",X"55",X"15",X"55",X"55",X"55",X"55",X"55",X"75",X"55",X"77",X"55",
		X"77",X"47",X"F7",X"47",X"DF",X"75",X"5D",X"D5",X"55",X"D5",X"55",X"55",X"55",X"15",X"54",X"15",
		X"AF",X"AF",X"AF",X"EA",X"AB",X"FF",X"EB",X"BF",X"AB",X"AA",X"AA",X"EA",X"AB",X"AB",X"EA",X"AA",
		X"FB",X"3F",X"FF",X"FF",X"AB",X"FF",X"FE",X"BF",X"FF",X"EF",X"AB",X"FB",X"EF",X"AB",X"AB",X"BF",
		X"AF",X"EA",X"AB",X"FF",X"BB",X"AF",X"AA",X"EA",X"AA",X"AB",X"AE",X"AB",X"AA",X"AA",X"AA",X"BA",
		X"AB",X"FF",X"FE",X"BF",X"FF",X"EF",X"AF",X"EB",X"AB",X"FE",X"AE",X"FF",X"BA",X"FF",X"BA",X"AF",
		X"FF",X"FF",X"BF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"BF",X"FF",X"EF",X"FB",X"FB",X"FF",
		X"3F",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",X"EF",X"FF",X"BC",X"FE",X"F3",X"FB",X"CF",X"FB",X"F3",
		X"FE",X"FC",X"FF",X"BF",X"FF",X"EF",X"FF",X"FB",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"7F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AF",X"FF",X"FF",X"FF",X"FF",X"FF",X"5F",
		X"FF",X"57",X"DD",X"55",X"D5",X"55",X"55",X"95",X"55",X"99",X"56",X"25",X"65",X"41",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"F3",X"FF",X"FD",X"FF",X"3F",X"FF",X"FF",X"FF",X"F5",
		X"FF",X"D5",X"FF",X"D6",X"D7",X"56",X"75",X"65",X"75",X"95",X"D6",X"55",X"F5",X"A4",X"D5",X"68",
		X"FA",X"FF",X"AF",X"01",X"F0",X"FD",X"0F",X"FD",X"FF",X"A9",X"FA",X"F5",X"EF",X"F5",X"FA",X"FD",
		X"FF",X"AF",X"3F",X"FA",X"C3",X"FF",X"FC",X"3F",X"FF",X"C3",X"AF",X"FC",X"FA",X"FF",X"FF",X"AF",
		X"F7",X"56",X"FD",X"55",X"D6",X"55",X"D6",X"A9",X"55",X"55",X"D5",X"5A",X"F4",X"55",X"D5",X"59",
		X"FF",X"FF",X"FF",X"FF",X"30",X"CC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",
		X"51",X"15",X"55",X"54",X"55",X"55",X"56",X"45",X"12",X"59",X"54",X"94",X"5A",X"55",X"64",X"55",
		X"FF",X"FF",X"FA",X"FF",X"BE",X"BA",X"FB",X"AA",X"FE",X"AA",X"FA",X"89",X"EA",X"29",X"EA",X"A9",
		X"15",X"05",X"25",X"80",X"89",X"AA",X"A2",X"A2",X"2A",X"A2",X"68",X"AA",X"88",X"A8",X"A2",X"82",
		X"65",X"14",X"56",X"02",X"45",X"6A",X"95",X"6A",X"05",X"2A",X"50",X"0A",X"12",X"AA",X"AE",X"6A",
		X"FA",X"85",X"A0",X"25",X"A2",X"2A",X"8A",X"82",X"8A",X"AA",X"A0",X"8A",X"AA",X"AA",X"8A",X"8A",
		X"FF",X"FE",X"FF",X"EA",X"FF",X"BA",X"FE",X"AA",X"FA",X"A8",X"FE",X"AA",X"FE",X"EA",X"A5",X"5A",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F3",X"FF",X"3F",X"FF",X"FF",X"F3",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"EC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F3",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FE",X"BF",X"FF",X"F3",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"CF",X"FA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"BA",X"E5",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FB",X"FF",X"FF",X"FF",X"FF",X"FA",X"AA",X"A5",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AE",X"BA",X"55",X"55",X"55",X"55",X"55",X"57",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FA",X"AA",X"E5",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"FF",X"FF",
		X"FF",X"FE",X"EB",X"A5",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"7F",X"FF",X"FF",X"FF",
		X"EA",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"57",X"55",X"55",X"FF",X"FF",X"FF",X"AA",
		X"55",X"68",X"55",X"AA",X"7D",X"6A",X"FF",X"D9",X"FE",X"F7",X"FA",X"AF",X"FE",X"AB",X"AA",X"AA",
		X"28",X"26",X"AA",X"AD",X"5A",X"AF",X"F6",X"9F",X"F5",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"9D",X"82",X"7D",X"A0",X"F6",X"A8",X"F6",X"AA",X"F6",X"5A",X"FF",X"F5",X"FF",X"FF",X"EA",X"BF",
		X"2A",X"AA",X"2A",X"6A",X"2A",X"8A",X"A8",X"8A",X"56",X"0A",X"FD",X"66",X"FD",X"AA",X"FD",X"AA",
		X"FF",X"6A",X"FF",X"D9",X"FF",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AF",X"AA",X"AF",X"AA",X"AB",X"AA",X"AF",X"AF",X"BF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"EA",X"FF",X"EA",X"FB",X"EA",X"FE",X"AA",X"AA",X"AA",X"AA",X"AF",X"AA",X"FE",X"BF",X"FF",
		X"AA",X"AA",X"AA",X"AB",X"EF",X"FF",X"FF",X"FF",X"FB",X"FF",X"EA",X"FE",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"FE",X"AA",X"FA",X"AA",
		X"AB",X"FF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AF",X"FF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FA",X"AA",X"FF",X"EA",X"FF",X"FA",X"FF",X"FF",
		X"5F",X"FB",X"FA",X"AA",X"EA",X"AA",X"AA",X"AA",X"AA",X"AB",X"AB",X"EF",X"EF",X"FF",X"FF",X"FF",
		X"55",X"55",X"5F",X"FF",X"7F",X"EA",X"FF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AB",X"AA",X"BF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"7F",X"55",X"FF",X"FF",X"FE",X"FF",X"AA",X"EA",X"AA",
		X"AA",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"57",X"55",X"5F",
		X"FF",X"FF",X"EB",X"A9",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FE",X"BA",X"A9",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"3F",X"FF",X"FF",X"FF",X"FF",X"EA",X"BA",X"95",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"EB",X"E9",X"95",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"EF",X"FF",X"FF",X"FF",X"FF",X"BF",X"FF",X"FF",X"FE",X"BE",X"F9",X"55",
		X"FF",X"F7",X"FF",X"D5",X"FF",X"D7",X"FF",X"57",X"FF",X"45",X"FD",X"05",X"FD",X"D5",X"A9",X"D5",
		X"FF",X"FF",X"55",X"00",X"C1",X"40",X"55",X"55",X"55",X"55",X"55",X"DF",X"55",X"F7",X"55",X"07",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F3",X"FF",X"3F",X"F3",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"33",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",
		X"FF",X"FD",X"FF",X"FD",X"00",X"01",X"00",X"01",X"00",X"01",X"55",X"55",X"55",X"55",X"FF",X"FD",
		X"55",X"41",X"55",X"55",X"55",X"55",X"55",X"7D",X"55",X"7D",X"55",X"41",X"55",X"41",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FE",X"FF",X"E8",X"FF",X"AC",X"FF",X"BF",X"FF",X"EB",X"FF",X"FE",X"FF",X"FF",
		X"FA",X"00",X"A0",X"3F",X"03",X"FE",X"FF",X"FA",X"0F",X"FF",X"F3",X"FF",X"BC",X"3F",X"EF",X"C0",
		X"01",X"15",X"FD",X"15",X"A9",X"D5",X"FF",X"D5",X"AF",X"D5",X"FA",X"FD",X"FF",X"AF",X"FF",X"FA",
		X"C4",X"75",X"FC",X"7D",X"AF",X"FD",X"FA",X"FD",X"FF",X"AF",X"3F",X"FA",X"C3",X"FF",X"FC",X"3F",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"FF",X"FF",
		X"FF",X"FF",X"AF",X"AA",X"FF",X"FF",X"FF",X"FF",X"03",X"00",X"FF",X"FF",X"AE",X"AA",X"FF",X"FF",
		X"EB",X"FF",X"FE",X"AA",X"FF",X"FF",X"3F",X"FF",X"C0",X"00",X"FF",X"FF",X"AA",X"AA",X"FF",X"FF",
		X"0F",X"FF",X"F0",X"FF",X"BF",X"03",X"EB",X"FC",X"FE",X"AF",X"FF",X"FA",X"FF",X"FF",X"FF",X"FF",
		X"FA",X"FF",X"FF",X"AB",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"FF",X"F3",X"3F",
		X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"F3",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"AA",X"AA",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"AA",X"AA",X"FF",X"FF",
		X"FF",X"FF",X"AA",X"AA",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"EA",X"AA",X"FF",X"FF",
		X"FF",X"FF",X"AA",X"AA",X"FF",X"FF",X"FF",X"FF",X"0C",X"00",X"FF",X"FF",X"BA",X"AA",X"FF",X"FF",
		X"FF",X"FF",X"AA",X"AE",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"EA",X"AA",X"FF",X"FF",
		X"FF",X"FF",X"AA",X"AA",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"AA",X"AA",X"FF",X"FF",
		X"FF",X"FF",X"AA",X"AA",X"FF",X"FF",X"FF",X"FF",X"00",X"C0",X"FF",X"FF",X"AB",X"FA",X"FF",X"FF",
		X"FF",X"FF",X"AA",X"FA",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"AA",X"AA",X"FF",X"FF",
		X"FF",X"FF",X"AA",X"AA",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"AA",X"BA",X"FF",X"FF",
		X"FF",X"FF",X"AA",X"BE",X"FF",X"FF",X"FF",X"FF",X"C0",X"00",X"FF",X"FF",X"AA",X"AA",X"FF",X"FF",
		X"FF",X"FE",X"AA",X"AB",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FE",X"AA",X"AB",X"FF",X"FF",
		X"BC",X"2F",X"FF",X"0B",X"F0",X"EF",X"0E",X"BF",X"EB",X"FF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FC",
		X"FF",X"FF",X"33",X"FF",X"FF",X"3F",X"FF",X"CF",X"FF",X"FF",X"BF",X"FF",X"2B",X"FF",X"C2",X"BF",
		X"FF",X"FF",X"BF",X"FF",X"2B",X"FF",X"C2",X"BF",X"BC",X"2B",X"EB",X"C2",X"FE",X"BC",X"FF",X"EB",
		X"4D",X"D5",X"51",X"DF",X"51",X"FF",X"51",X"1F",X"D1",X"1F",X"FD",X"13",X"AF",X"D0",X"FA",X"FC",
		X"00",X"01",X"00",X"01",X"00",X"01",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"FF",X"FD",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"FF",X"FF",X"FF",X"F3",
		X"F7",X"FF",X"01",X"FF",X"00",X"7F",X"55",X"7F",X"55",X"5F",X"FF",X"DF",X"FF",X"F7",X"FF",X"F7",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"03",X"F0",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FB",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"FF",X"7F",X"FF",X"40",X"00",X"40",X"00",X"40",X"00",X"55",X"55",X"55",X"55",X"7F",X"FF",
		X"3F",X"FF",X"CF",X"FF",X"F3",X"FF",X"FC",X"FF",X"FF",X"C3",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"FF",X"C3",X"3F",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"C3",X"AF",X"FC",X"FA",X"FF",X"FF",X"AF",X"FF",X"FA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"AF",X"3F",X"FA",X"C3",X"FF",X"FC",X"3F",X"FF",X"C0",X"AF",X"FF",X"FA",X"AA",X"FF",X"FF",
		X"FF",X"FF",X"AA",X"AA",X"FF",X"FF",X"FF",X"FF",X"03",X"00",X"FF",X"FF",X"AE",X"AA",X"FF",X"FF",
		X"00",X"00",X"15",X"40",X"7F",X"D4",X"1F",X"FD",X"1F",X"7F",X"1F",X"5F",X"1F",X"5F",X"1F",X"5F",
		X"00",X"00",X"15",X"40",X"7F",X"D0",X"1F",X"40",X"5F",X"40",X"5F",X"41",X"DF",X"41",X"DF",X"41",
		X"00",X"00",X"10",X"15",X"74",X"7F",X"7D",X"1F",X"7D",X"1F",X"FF",X"47",X"FF",X"47",X"FF",X"41",
		X"00",X"00",X"40",X"55",X"D1",X"FF",X"40",X"77",X"D1",X"F7",X"D1",X"D7",X"F7",X"D7",X"F7",X"47",
		X"00",X"00",X"55",X"05",X"FF",X"5F",X"FF",X"57",X"DF",X"D7",X"D7",X"D7",X"D1",X"D7",X"D0",X"47",
		X"00",X"00",X"55",X"40",X"FF",X"D0",X"DF",X"F4",X"D7",X"F4",X"D7",X"FD",X"D5",X"FD",X"D1",X"FD",
		X"1F",X"5F",X"1F",X"5F",X"1A",X"5A",X"1A",X"5A",X"1A",X"5A",X"1A",X"5A",X"1A",X"9A",X"1A",X"AA",
		X"DF",X"41",X"DF",X"47",X"9A",X"46",X"9A",X"46",X"9A",X"46",X"9A",X"46",X"9A",X"46",X"5A",X"46",
		X"F7",X"D1",X"F7",X"D0",X"A6",X"90",X"96",X"90",X"91",X"A4",X"96",X"A4",X"9A",X"A4",X"A9",X"A4",
		X"FF",X"47",X"7D",X"07",X"69",X"06",X"69",X"06",X"69",X"06",X"69",X"06",X"69",X"06",X"69",X"06",
		X"D4",X"07",X"DD",X"07",X"AA",X"46",X"AA",X"46",X"9A",X"46",X"96",X"46",X"91",X"06",X"90",X"46",
		X"D1",X"FD",X"D1",X"FD",X"A6",X"A4",X"AA",X"90",X"9A",X"90",X"9A",X"90",X"9A",X"90",X"96",X"A4",
		X"1F",X"FD",X"1F",X"54",X"1F",X"40",X"1F",X"40",X"1F",X"40",X"1F",X"40",X"1F",X"40",X"1F",X"40",
		X"1F",X"47",X"1F",X"5F",X"1F",X"5F",X"1F",X"5F",X"1F",X"7D",X"1F",X"F4",X"1F",X"D0",X"1F",X"40",
		X"F5",X"FD",X"D1",X"FD",X"D0",X"7D",X"F5",X"FF",X"50",X"55",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7D",X"07",X"7D",X"07",X"7D",X"07",X"FF",X"5F",X"55",X"05",X"00",X"00",X"00",X"00",X"00",X"00",
		X"D1",X"D7",X"F7",X"D7",X"FF",X"D7",X"FF",X"D7",X"FF",X"D7",X"5F",X"D7",X"05",X"7F",X"00",X"17",
		X"D7",X"F4",X"D7",X"F4",X"D1",X"F4",X"D1",X"FD",X"D1",X"FD",X"D1",X"FD",X"F4",X"7D",X"F4",X"7D",
		X"1F",X"40",X"1F",X"40",X"1F",X"40",X"1F",X"40",X"1F",X"50",X"1F",X"74",X"1F",X"F4",X"1F",X"D0",
		X"7D",X"00",X"14",X"55",X"01",X"FF",X"07",X"F5",X"07",X"D0",X"1F",X"D0",X"1A",X"90",X"1A",X"90",
		X"00",X"00",X"50",X"55",X"F5",X"FF",X"FD",X"7F",X"7D",X"7F",X"7F",X"7F",X"6A",X"69",X"6A",X"69",
		X"00",X"00",X"01",X"55",X"47",X"FF",X"D1",X"D7",X"F5",X"D7",X"FD",X"D7",X"A9",X"96",X"AA",X"96",
		X"00",X"41",X"55",X"D0",X"FF",X"D0",X"FF",X"F4",X"D5",X"74",X"D7",X"50",X"AA",X"40",X"AA",X"40",
		X"FD",X"7F",X"7D",X"7F",X"15",X"FF",X"01",X"FF",X"00",X"7F",X"00",X"1F",X"00",X"1F",X"00",X"07",
		X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"D0",X"00",X"D0",X"00",X"F4",X"00",
		X"7F",X"40",X"FD",X"00",X"F4",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1A",X"90",X"1F",X"D0",X"1F",X"D0",X"07",X"F5",X"01",X"FF",X"00",X"55",X"00",X"00",X"00",X"00",
		X"6A",X"69",X"7F",X"7D",X"7D",X"7D",X"FD",X"7D",X"F5",X"FF",X"50",X"55",X"00",X"00",X"00",X"00",
		X"6A",X"96",X"1F",X"D7",X"1F",X"D7",X"07",X"D7",X"47",X"DF",X"01",X"45",X"00",X"00",X"00",X"00",
		X"96",X"40",X"D1",X"04",X"F5",X"5D",X"FF",X"FD",X"FF",X"F4",X"55",X"50",X"00",X"00",X"00",X"00",
		X"F4",X"00",X"7D",X"00",X"1D",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"15",X"40",X"6A",X"94",X"1A",X"A9",X"1A",X"6A",X"1A",X"5A",X"1A",X"5A",X"1A",X"5A",
		X"00",X"00",X"15",X"40",X"6A",X"90",X"1A",X"40",X"5A",X"40",X"5A",X"41",X"9A",X"41",X"9A",X"41",
		X"00",X"00",X"10",X"15",X"64",X"6A",X"69",X"1A",X"69",X"1A",X"AA",X"46",X"AA",X"46",X"AA",X"41",
		X"00",X"00",X"40",X"55",X"91",X"AA",X"40",X"66",X"91",X"A6",X"91",X"96",X"A6",X"96",X"A6",X"46",
		X"00",X"00",X"55",X"05",X"AA",X"5A",X"AA",X"56",X"9A",X"96",X"96",X"96",X"91",X"96",X"90",X"46",
		X"00",X"00",X"55",X"40",X"AA",X"90",X"9A",X"A4",X"96",X"A4",X"96",X"A9",X"95",X"A9",X"91",X"A9",
		X"1A",X"5A",X"1A",X"5A",X"1A",X"5A",X"1A",X"5A",X"1A",X"5A",X"1A",X"5A",X"1A",X"9A",X"1A",X"AA",
		X"9A",X"41",X"9A",X"46",X"9A",X"46",X"9A",X"46",X"9A",X"46",X"9A",X"46",X"9A",X"46",X"5A",X"46",
		X"A6",X"91",X"A6",X"90",X"A6",X"90",X"96",X"90",X"91",X"A4",X"96",X"A4",X"9A",X"A4",X"A9",X"A4",
		X"AA",X"46",X"69",X"06",X"69",X"06",X"69",X"06",X"69",X"06",X"69",X"06",X"69",X"06",X"69",X"06",
		X"94",X"06",X"99",X"06",X"AA",X"46",X"AA",X"46",X"9A",X"46",X"96",X"46",X"91",X"06",X"90",X"46",
		X"91",X"A9",X"91",X"A9",X"A6",X"A4",X"AA",X"90",X"9A",X"90",X"9A",X"90",X"9A",X"90",X"96",X"A4",
		X"1A",X"A9",X"1A",X"54",X"1A",X"40",X"1A",X"40",X"1A",X"40",X"1A",X"40",X"1A",X"40",X"1A",X"40",
		X"1A",X"46",X"1A",X"5A",X"1A",X"5A",X"1A",X"5A",X"1A",X"69",X"1A",X"A4",X"1A",X"90",X"1A",X"40",
		X"A5",X"A9",X"91",X"A9",X"90",X"69",X"A5",X"AA",X"50",X"55",X"00",X"00",X"00",X"00",X"00",X"00",
		X"69",X"06",X"69",X"06",X"69",X"06",X"AA",X"5A",X"55",X"05",X"00",X"00",X"00",X"00",X"00",X"00",
		X"91",X"96",X"A6",X"96",X"AA",X"96",X"AA",X"96",X"AA",X"96",X"5A",X"96",X"05",X"6A",X"00",X"16",
		X"96",X"A4",X"96",X"A4",X"91",X"A4",X"91",X"A9",X"91",X"A9",X"91",X"A9",X"A4",X"69",X"A4",X"69",
		X"1A",X"40",X"1A",X"40",X"1A",X"41",X"1A",X"41",X"1A",X"51",X"1A",X"64",X"1A",X"A4",X"1A",X"90",
		X"69",X"00",X"65",X"55",X"AA",X"AA",X"AA",X"AA",X"A5",X"A5",X"51",X"A4",X"01",X"A4",X"01",X"A4",
		X"40",X"00",X"95",X"50",X"AA",X"A4",X"A6",X"91",X"A6",X"96",X"56",X"91",X"06",X"A5",X"01",X"A6",
		X"00",X"00",X"01",X"54",X"06",X"A9",X"51",X"A5",X"A5",X"A5",X"91",X"A6",X"96",X"A6",X"A6",X"96",
		X"00",X"01",X"15",X"54",X"6A",X"A9",X"A9",X"6A",X"A4",X"1A",X"A4",X"1A",X"A4",X"1A",X"A4",X"1A",
		X"A9",X"6A",X"69",X"6A",X"15",X"AA",X"41",X"AA",X"40",X"6A",X"90",X"1A",X"90",X"1A",X"90",X"06",
		X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"90",X"00",X"90",X"00",X"A4",X"00",
		X"A4",X"00",X"69",X"00",X"19",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A4",X"1A",X"A4",X"1A",X"A4",X"1A",X"A9",X"6A",X"6A",X"A9",X"15",X"54",X"00",X"00",X"00",X"00",
		X"90",X"01",X"90",X"00",X"40",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"96",X"6A",X"96",X"1A",X"91",X"1A",X"41",X"06",X"40",X"01",X"00",X"00",X"00",X"00",X"00",
		X"01",X"A6",X"01",X"AA",X"01",X"A9",X"00",X"69",X"00",X"64",X"00",X"10",X"00",X"00",X"00",X"00",
		X"01",X"A4",X"01",X"A4",X"01",X"A4",X"01",X"A4",X"06",X"A9",X"01",X"54",X"00",X"00",X"00",X"00",
		X"6A",X"40",X"A9",X"00",X"A4",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"D5",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"57",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"80",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AB",X"55",X"AB",X"55",X"AD",X"55",X"AD",X"55",X"B5",X"55",X"B5",X"55",X"D5",X"55",X"D5",X"55",
		X"AA",X"AB",X"AA",X"AB",X"AA",X"AD",X"AA",X"AD",X"AA",X"B5",X"AA",X"B5",X"AA",X"D5",X"AA",X"D5",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FF",X"FF",
		X"FF",X"FF",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
