library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_8K is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_8K is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"02",X"03",X"0F",X"00",X"00",X"30",X"70",X"E0",X"ED",X"6F",X"6F",
		X"07",X"0F",X"03",X"02",X"00",X"00",X"00",X"00",X"7C",X"6F",X"6F",X"ED",X"E0",X"70",X"30",X"00",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CF",X"CF",X"CF",X"CF",X"C0",X"C0",X"FF",X"FF",
		X"CC",X"CC",X"CF",X"CF",X"C0",X"C0",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"F3",X"F3",X"F3",X"F3",X"03",X"03",X"FF",X"FF",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"33",X"33",X"F3",X"F3",X"03",X"03",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"03",X"03",X"F3",X"F3",X"33",X"33",
		X"FF",X"FF",X"03",X"03",X"F3",X"F3",X"F3",X"F3",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"FF",X"FF",X"C0",X"C0",X"CF",X"CF",X"CC",X"CC",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"FF",X"FF",X"C0",X"C0",X"CF",X"CF",X"CF",X"CF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"82",X"C6",X"7C",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"7C",X"C6",X"82",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"38",X"7C",X"C2",X"82",X"86",X"7C",X"38",X"00",X"00",X"02",X"02",X"FE",X"FE",X"42",X"02",X"00",
		X"62",X"F2",X"BA",X"9A",X"9E",X"CE",X"46",X"00",X"8C",X"DE",X"F2",X"B2",X"92",X"86",X"04",X"00",
		X"08",X"FE",X"FE",X"C8",X"68",X"38",X"18",X"00",X"9C",X"BE",X"A2",X"A2",X"A2",X"E6",X"E4",X"00",
		X"0C",X"9E",X"92",X"92",X"D2",X"7E",X"3C",X"00",X"C0",X"E0",X"B0",X"9E",X"8E",X"C0",X"C0",X"00",
		X"6C",X"FE",X"92",X"92",X"92",X"FE",X"6C",X"00",X"78",X"FC",X"96",X"92",X"92",X"F2",X"60",X"00",
		X"7C",X"82",X"AA",X"AA",X"BA",X"82",X"7C",X"00",X"7C",X"82",X"BA",X"AA",X"BE",X"82",X"7C",X"00",
		X"2E",X"2E",X"3A",X"3A",X"00",X"20",X"7E",X"7E",X"00",X"00",X"00",X"E0",X"C0",X"00",X"00",X"00",
		X"20",X"00",X"70",X"50",X"50",X"7E",X"7E",X"00",X"00",X"00",X"00",X"F0",X"FA",X"FA",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"7E",X"C8",X"88",X"C8",X"7E",X"3E",X"00",
		X"6C",X"FE",X"92",X"92",X"92",X"FE",X"FE",X"00",X"44",X"C6",X"82",X"82",X"C6",X"7C",X"38",X"00",
		X"38",X"7C",X"C6",X"82",X"82",X"FE",X"FE",X"00",X"00",X"82",X"92",X"92",X"92",X"FE",X"FE",X"00",
		X"80",X"90",X"90",X"90",X"90",X"FE",X"FE",X"00",X"9E",X"9E",X"92",X"82",X"C6",X"7C",X"38",X"00",
		X"FE",X"FE",X"10",X"10",X"10",X"FE",X"FE",X"00",X"00",X"82",X"82",X"FE",X"FE",X"82",X"82",X"00",
		X"FC",X"FE",X"02",X"02",X"02",X"06",X"04",X"00",X"82",X"C6",X"6E",X"3C",X"18",X"FE",X"FE",X"00",
		X"00",X"02",X"02",X"02",X"02",X"FE",X"FE",X"00",X"FE",X"FE",X"70",X"38",X"70",X"FE",X"FE",X"00",
		X"FE",X"FE",X"1C",X"38",X"70",X"FE",X"FE",X"00",X"7C",X"FE",X"82",X"82",X"82",X"FE",X"7C",X"00",
		X"70",X"88",X"88",X"88",X"88",X"FE",X"FE",X"00",X"7A",X"FC",X"8E",X"8A",X"82",X"FE",X"7C",X"00",
		X"72",X"F6",X"9E",X"8C",X"88",X"FE",X"FE",X"00",X"4C",X"DE",X"92",X"92",X"92",X"F6",X"64",X"00",
		X"00",X"80",X"80",X"FE",X"FE",X"80",X"80",X"00",X"FC",X"FE",X"02",X"02",X"02",X"FE",X"FC",X"00",
		X"F0",X"F8",X"1C",X"0E",X"1C",X"F8",X"F0",X"00",X"FC",X"FE",X"1C",X"38",X"1C",X"FE",X"FC",X"00",
		X"C6",X"EE",X"7C",X"38",X"7C",X"EE",X"C6",X"00",X"00",X"C0",X"F0",X"1E",X"1E",X"F0",X"C0",X"00",
		X"C2",X"E2",X"F2",X"BA",X"9E",X"8E",X"86",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"FF",
		X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"14",X"14",X"95",X"95",X"95",X"95",X"95",X"95",X"95",
		X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",
		X"7F",X"00",X"FF",X"00",X"FF",X"00",X"00",X"7F",X"FE",X"00",X"FF",X"00",X"FF",X"00",X"00",X"FE",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"00",X"FF",
		X"95",X"94",X"97",X"90",X"9F",X"80",X"80",X"FF",X"FF",X"80",X"9F",X"90",X"97",X"94",X"94",X"95",
		X"95",X"15",X"F5",X"05",X"FD",X"01",X"01",X"FF",X"FF",X"01",X"FD",X"05",X"F5",X"15",X"15",X"95",
		X"95",X"14",X"D7",X"00",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"FF",X"00",X"FF",X"14",X"14",X"95",
		X"95",X"94",X"97",X"90",X"97",X"90",X"94",X"95",X"95",X"15",X"F5",X"15",X"F5",X"15",X"15",X"95",
		X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"14",X"14",X"95",X"95",X"95",X"95",X"95",X"95",X"95",
		X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",
		X"7F",X"00",X"FF",X"00",X"FF",X"00",X"00",X"7F",X"FE",X"00",X"FF",X"00",X"FF",X"00",X"00",X"FE",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"00",X"FF",
		X"95",X"94",X"97",X"90",X"9F",X"80",X"80",X"FF",X"FF",X"80",X"9F",X"90",X"97",X"94",X"94",X"95",
		X"95",X"15",X"F5",X"05",X"FD",X"01",X"01",X"FF",X"FF",X"01",X"FD",X"05",X"F5",X"15",X"15",X"95",
		X"95",X"14",X"D7",X"00",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"FF",X"00",X"FF",X"14",X"14",X"95",
		X"95",X"94",X"97",X"90",X"97",X"90",X"94",X"95",X"95",X"15",X"F5",X"15",X"F5",X"15",X"15",X"95",
		X"00",X"00",X"00",X"00",X"00",X"02",X"01",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"38",
		X"0C",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"18",X"C0",X"E0",X"20",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",X"E0",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"04",X"08",X"10",X"20",X"20",X"00",X"00",X"C0",X"20",X"10",X"08",X"04",X"04",
		X"20",X"20",X"10",X"08",X"04",X"03",X"00",X"00",X"04",X"04",X"08",X"10",X"20",X"C0",X"00",X"00",
		X"07",X"08",X"10",X"20",X"40",X"80",X"80",X"80",X"E0",X"10",X"08",X"04",X"02",X"01",X"01",X"01",
		X"80",X"80",X"80",X"40",X"20",X"10",X"08",X"07",X"01",X"01",X"01",X"02",X"04",X"08",X"10",X"E0",
		X"20",X"00",X"00",X"80",X"28",X"A8",X"5C",X"24",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"5F",X"2F",X"AF",X"08",X"00",X"24",X"00",X"20",X"FF",X"FF",X"FE",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"08",X"81",X"03",X"50",X"00",X"27",X"00",X"00",X"40",X"E0",X"F8",X"3C",X"0E",X"86",
		X"07",X"57",X"03",X"83",X"09",X"00",X"00",X"00",X"E3",X"F3",X"F0",X"F8",X"F8",X"70",X"00",X"00",
		X"00",X"00",X"40",X"09",X"03",X"50",X"A8",X"43",X"00",X"00",X"40",X"E0",X"F8",X"3C",X"0E",X"86",
		X"27",X"17",X"27",X"83",X"21",X"14",X"00",X"20",X"E3",X"F3",X"F0",X"F8",X"F8",X"70",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"14",X"14",X"95",X"95",X"95",X"95",X"95",X"95",X"95",
		X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",
		X"7F",X"00",X"FF",X"00",X"FF",X"00",X"00",X"7F",X"FE",X"00",X"FF",X"00",X"FF",X"00",X"00",X"FE",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"00",X"FF",
		X"95",X"94",X"97",X"90",X"9F",X"80",X"80",X"FF",X"FF",X"80",X"9F",X"90",X"97",X"94",X"94",X"95",
		X"95",X"15",X"F5",X"05",X"FD",X"01",X"01",X"FF",X"FF",X"01",X"FD",X"05",X"F5",X"15",X"15",X"95",
		X"95",X"14",X"D7",X"00",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"FF",X"00",X"FF",X"14",X"14",X"95",
		X"95",X"94",X"97",X"90",X"97",X"90",X"94",X"95",X"95",X"15",X"F5",X"15",X"F5",X"15",X"15",X"95",
		X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"14",X"14",X"95",X"95",X"95",X"95",X"95",X"95",X"95",
		X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",
		X"7F",X"00",X"FF",X"00",X"FF",X"00",X"00",X"7F",X"FE",X"00",X"FF",X"00",X"FF",X"00",X"00",X"FE",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"00",X"FF",
		X"95",X"94",X"97",X"90",X"9F",X"80",X"80",X"FF",X"FF",X"80",X"9F",X"90",X"97",X"94",X"94",X"95",
		X"95",X"15",X"F5",X"05",X"FD",X"01",X"01",X"FF",X"FF",X"01",X"FD",X"05",X"F5",X"15",X"15",X"95",
		X"95",X"14",X"D7",X"00",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"FF",X"00",X"FF",X"14",X"14",X"95",
		X"95",X"94",X"97",X"90",X"97",X"90",X"94",X"95",X"95",X"15",X"F5",X"15",X"F5",X"15",X"15",X"95",
		X"C0",X"C2",X"C1",X"C0",X"C0",X"C0",X"C1",X"C2",X"03",X"0B",X"13",X"A3",X"43",X"A3",X"13",X"0B",
		X"C0",X"C0",X"C0",X"C0",X"FF",X"FF",X"FF",X"FF",X"03",X"03",X"03",X"03",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"C0",X"C0",X"C0",X"C0",X"FF",X"FF",X"FF",X"FF",X"03",X"03",X"03",X"1B",
		X"C0",X"DF",X"DF",X"C6",X"C6",X"C0",X"C0",X"C0",X"1B",X"FB",X"FB",X"1B",X"1B",X"03",X"03",X"03",
		X"FF",X"FF",X"FF",X"FF",X"C0",X"CF",X"DF",X"DD",X"FF",X"FF",X"FF",X"FF",X"03",X"1B",X"9B",X"9B",
		X"D9",X"D8",X"D8",X"DC",X"DE",X"CE",X"C0",X"C0",X"DB",X"FB",X"FB",X"7B",X"3B",X"1B",X"03",X"03",
		X"FF",X"FF",X"FF",X"FF",X"C0",X"DC",X"DF",X"DF",X"FF",X"FF",X"FF",X"FF",X"03",X"F3",X"FB",X"FB",
		X"DB",X"DB",X"DB",X"D8",X"D8",X"D8",X"C0",X"C0",X"3B",X"1B",X"1B",X"3B",X"7B",X"73",X"03",X"03",
		X"FF",X"FF",X"FF",X"FF",X"C0",X"C0",X"DF",X"DF",X"FF",X"FF",X"FF",X"FF",X"03",X"63",X"FB",X"FB",
		X"DC",X"CE",X"C7",X"C3",X"C1",X"C0",X"C0",X"C0",X"63",X"63",X"63",X"E3",X"E3",X"E3",X"03",X"03",
		X"FF",X"FF",X"FF",X"FF",X"C0",X"C1",X"DB",X"DB",X"FF",X"FF",X"FF",X"FF",X"03",X"F3",X"FB",X"BB",
		X"DB",X"DB",X"DB",X"DB",X"DF",X"DF",X"C0",X"C0",X"1B",X"1B",X"1B",X"3B",X"7B",X"73",X"03",X"03",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"2B",X"14",X"0B",X"04",X"03",X"00",X"00",X"00",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",
		X"00",X"00",X"03",X"04",X"0B",X"14",X"2B",X"2A",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"A8",X"50",X"A0",X"40",X"80",X"00",X"00",X"00",
		X"A8",X"A8",X"A8",X"A8",X"A8",X"A8",X"A8",X"A8",X"00",X"00",X"80",X"40",X"A0",X"50",X"A8",X"A8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"18",X"10",X"00",X"20",X"20",
		X"06",X"07",X"03",X"03",X"03",X"03",X"02",X"02",X"58",X"DE",X"C3",X"01",X"03",X"1F",X"D8",X"00",
		X"00",X"0F",X"24",X"C0",X"C0",X"63",X"3F",X"1E",X"00",X"00",X"01",X"00",X"C0",X"E3",X"15",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CF",X"CF",X"CF",X"CF",X"CF",X"CF",X"CF",X"CF",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CF",X"CF",X"CF",X"CF",X"CF",X"CF",X"CF",X"CF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"F3",X"F3",X"F3",X"F3",X"F3",X"F3",X"F3",X"F3",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"F3",X"F3",X"F3",X"F3",X"F3",X"F3",X"F3",X"F3",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"C0",X"C0",X"C0",X"E0",X"E0",X"E0",X"E0",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"F0",X"F0",X"F0",X"F0",X"F8",X"00",X"00",X"FF",X"01",X"01",X"01",X"03",X"02",X"06",X"1C",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F9",X"79",X"79",X"79",X"39",X"39",X"19",X"19",
		X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"19",X"09",X"09",X"01",X"01",X"01",X"01",X"01",
		X"3F",X"3F",X"1F",X"1F",X"1F",X"0F",X"0F",X"07",X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",
		X"07",X"07",X"03",X"03",X"01",X"01",X"01",X"00",X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"81",X"C1",X"E1",X"E1",X"F1",X"F9",X"F9",X"F9",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",
		X"3E",X"1C",X"09",X"03",X"03",X"01",X"00",X"C0",X"79",X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",X"79",
		X"E0",X"F0",X"F0",X"F8",X"FC",X"FE",X"FF",X"FF",X"39",X"19",X"09",X"01",X"01",X"01",X"01",X"81",
		X"1F",X"83",X"80",X"80",X"20",X"78",X"7E",X"3F",X"E1",X"E1",X"61",X"01",X"01",X"01",X"01",X"81",
		X"0F",X"07",X"01",X"80",X"E0",X"F0",X"F8",X"7C",X"E1",X"E1",X"C1",X"C1",X"01",X"01",X"19",X"39",
		X"00",X"00",X"01",X"00",X"00",X"E0",X"80",X"00",X"01",X"81",X"81",X"81",X"39",X"79",X"39",X"19",
		X"00",X"FE",X"FF",X"FF",X"00",X"00",X"00",X"7F",X"09",X"09",X"01",X"81",X"01",X"01",X"01",X"E1",
		X"7F",X"F8",X"F8",X"F8",X"38",X"F0",X"E0",X"C0",X"81",X"01",X"01",X"01",X"19",X"39",X"09",X"09",
		X"80",X"07",X"1F",X"3F",X"FF",X"FE",X"F8",X"60",X"09",X"89",X"89",X"89",X"89",X"09",X"09",X"01",
		X"0C",X"38",X"F8",X"F0",X"F0",X"E0",X"E0",X"C0",X"01",X"01",X"01",X"09",X"09",X"09",X"09",X"09",
		X"C0",X"81",X"03",X"07",X"0F",X"0F",X"1F",X"3F",X"89",X"89",X"89",X"89",X"89",X"81",X"81",X"81",
		X"00",X"0F",X"0F",X"1F",X"1F",X"1F",X"30",X"00",X"01",X"01",X"C1",X"C1",X"C1",X"C1",X"C1",X"41",
		X"0C",X"3E",X"7F",X"FF",X"FF",X"7F",X"3E",X"1C",X"19",X"09",X"09",X"01",X"01",X"01",X"01",X"01",
		X"C7",X"84",X"04",X"04",X"00",X"00",X"00",X"00",X"E1",X"01",X"01",X"01",X"41",X"41",X"41",X"C1",
		X"00",X"00",X"00",X"06",X"1C",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"1C",X"06",X"C2",X"E3",X"F1",X"F9",X"F9",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"F4",X"F9",X"F9",X"F9",X"E1",X"01",X"01",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"14",X"14",X"95",X"95",X"95",X"95",X"95",X"95",X"95",
		X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",
		X"7F",X"00",X"FF",X"00",X"FF",X"00",X"00",X"7F",X"FE",X"00",X"FF",X"00",X"FF",X"00",X"00",X"FE",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"00",X"FF",
		X"95",X"94",X"97",X"90",X"9F",X"80",X"80",X"FF",X"FF",X"80",X"9F",X"90",X"97",X"94",X"94",X"95",
		X"95",X"15",X"F5",X"05",X"FD",X"01",X"01",X"FF",X"FF",X"01",X"FD",X"05",X"F5",X"15",X"15",X"95",
		X"95",X"14",X"D7",X"00",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"FF",X"00",X"FF",X"14",X"14",X"95",
		X"95",X"94",X"97",X"90",X"97",X"90",X"94",X"95",X"95",X"15",X"F5",X"15",X"F5",X"15",X"15",X"95",
		X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"14",X"14",X"95",X"95",X"95",X"95",X"95",X"95",X"95",
		X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",
		X"7F",X"00",X"FF",X"00",X"FF",X"00",X"00",X"7F",X"FE",X"00",X"FF",X"00",X"FF",X"00",X"00",X"FE",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"00",X"FF",
		X"95",X"94",X"97",X"90",X"9F",X"80",X"80",X"FF",X"FF",X"80",X"9F",X"90",X"97",X"94",X"94",X"95",
		X"95",X"15",X"F5",X"05",X"FD",X"01",X"01",X"FF",X"FF",X"01",X"FD",X"05",X"F5",X"15",X"15",X"95",
		X"95",X"14",X"D7",X"00",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"FF",X"00",X"FF",X"14",X"14",X"95",
		X"95",X"94",X"97",X"90",X"97",X"90",X"94",X"95",X"95",X"15",X"F5",X"15",X"F5",X"15",X"15",X"95",
		X"00",X"00",X"00",X"07",X"04",X"07",X"00",X"07",X"00",X"00",X"00",X"C0",X"40",X"C0",X"00",X"C0",
		X"04",X"07",X"00",X"07",X"05",X"05",X"00",X"00",X"40",X"C0",X"00",X"40",X"40",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"06",X"0C",X"08",X"00",X"00",X"00",X"00",X"C0",X"60",X"30",X"10",
		X"08",X"0C",X"06",X"03",X"00",X"00",X"00",X"00",X"10",X"30",X"60",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"04",X"08",X"10",X"20",X"20",X"00",X"00",X"C0",X"20",X"10",X"08",X"04",X"04",
		X"20",X"20",X"10",X"08",X"04",X"03",X"00",X"00",X"04",X"04",X"08",X"10",X"20",X"C0",X"00",X"00",
		X"07",X"08",X"10",X"20",X"40",X"80",X"80",X"80",X"E0",X"10",X"08",X"04",X"02",X"01",X"01",X"01",
		X"80",X"80",X"80",X"40",X"20",X"10",X"08",X"07",X"01",X"01",X"01",X"02",X"04",X"08",X"10",X"E0",
		X"00",X"00",X"00",X"3E",X"22",X"3E",X"00",X"3E",X"00",X"00",X"00",X"00",X"74",X"54",X"5C",X"00",
		X"22",X"3E",X"00",X"3A",X"2A",X"2E",X"00",X"00",X"00",X"14",X"08",X"14",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"3E",X"22",X"3E",X"00",X"3E",X"00",X"00",X"00",X"00",X"7C",X"54",X"54",X"00",
		X"22",X"3E",X"00",X"3A",X"2A",X"2E",X"00",X"00",X"00",X"14",X"08",X"14",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"3E",X"22",X"3E",X"00",X"3E",X"00",X"00",X"00",X"00",X"7C",X"10",X"70",X"00",
		X"22",X"3E",X"00",X"3A",X"2A",X"2E",X"00",X"00",X"00",X"14",X"08",X"14",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"3E",X"22",X"3E",X"00",X"3E",X"00",X"00",X"00",X"00",X"5C",X"54",X"74",X"00",
		X"22",X"3E",X"00",X"3A",X"2A",X"2E",X"00",X"00",X"00",X"14",X"08",X"14",X"00",X"00",X"00",X"00",
		X"C3",X"C3",X"C3",X"C3",X"C3",X"C3",X"FF",X"FF",X"FF",X"FF",X"C3",X"C3",X"C3",X"C3",X"C3",X"C3",
		X"C3",X"C3",X"C3",X"C3",X"C3",X"C3",X"C3",X"C3",X"C3",X"C3",X"C3",X"C3",X"C3",X"C3",X"C3",X"C3",
		X"FF",X"81",X"85",X"9F",X"85",X"FD",X"81",X"FF",X"FF",X"81",X"DF",X"D3",X"D3",X"F3",X"81",X"FF",
		X"FF",X"81",X"DF",X"D3",X"D3",X"FF",X"81",X"FF",X"FF",X"81",X"FF",X"C1",X"C1",X"C1",X"81",X"FF",
		X"FF",X"81",X"FF",X"D3",X"D3",X"FF",X"81",X"FF",X"FF",X"81",X"FF",X"D3",X"D3",X"F3",X"81",X"FF",
		X"FF",X"81",X"FF",X"D1",X"D1",X"FF",X"81",X"FF",X"FF",X"81",X"9F",X"93",X"93",X"FF",X"81",X"FF",
		X"FF",X"81",X"E7",X"C3",X"C3",X"FF",X"81",X"FF",X"FF",X"81",X"FF",X"93",X"93",X"9F",X"81",X"FF",
		X"FF",X"81",X"C3",X"D3",X"D3",X"FF",X"81",X"FF",X"FF",X"81",X"C1",X"D1",X"D1",X"FF",X"81",X"FF",
		X"FF",X"81",X"FF",X"C3",X"C3",X"FF",X"81",X"FF",X"FF",X"81",X"83",X"FF",X"A3",X"81",X"81",X"FF",
		X"FF",X"81",X"FB",X"CB",X"CB",X"EF",X"81",X"FF",X"FF",X"81",X"FF",X"D3",X"C3",X"E7",X"81",X"FF",
		X"FF",X"81",X"85",X"9F",X"85",X"FD",X"81",X"FF",X"FF",X"81",X"DF",X"D3",X"D3",X"F3",X"81",X"FF",
		X"FF",X"81",X"DF",X"D3",X"D3",X"FF",X"81",X"FF",X"FF",X"81",X"FF",X"C1",X"C1",X"C1",X"81",X"FF",
		X"FF",X"81",X"FF",X"D3",X"D3",X"FF",X"81",X"FF",X"FF",X"81",X"FF",X"D3",X"D3",X"F3",X"81",X"FF",
		X"FF",X"81",X"FF",X"D1",X"D1",X"FF",X"81",X"FF",X"FF",X"81",X"9F",X"93",X"93",X"FF",X"81",X"FF",
		X"FF",X"81",X"E7",X"C3",X"C3",X"FF",X"81",X"FF",X"FF",X"81",X"FF",X"93",X"93",X"9F",X"81",X"FF",
		X"FF",X"81",X"C3",X"D3",X"D3",X"FF",X"81",X"FF",X"FF",X"81",X"C1",X"D1",X"D1",X"FF",X"81",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"08",X"1C",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"1F",X"0F",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FE",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"2F",X"00",X"00",X"00",X"00",X"E0",X"70",X"38",X"8C",
		X"57",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"C4",X"E0",X"F0",X"F0",X"60",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"03",X"00",X"00",X"13",X"00",X"00",X"40",X"E0",X"F8",X"3C",X"0E",X"86",
		X"2F",X"07",X"03",X"03",X"01",X"00",X"00",X"00",X"E3",X"F3",X"F0",X"F8",X"F8",X"70",X"00",X"00",
		X"00",X"00",X"00",X"01",X"03",X"00",X"00",X"07",X"00",X"00",X"40",X"E0",X"F8",X"3C",X"0E",X"86",
		X"07",X"07",X"03",X"03",X"01",X"00",X"00",X"00",X"E3",X"F3",X"F0",X"F8",X"F8",X"70",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"04",X"01",X"03",X"00",X"00",X"00",X"50",X"FC",X"50",X"FE",X"FE",
		X"03",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"00",X"00",X"00",X"30",X"FC",X"FE",X"FE",X"FF",
		X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FE",X"FE",X"FC",X"30",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"00",X"00",X"00",X"30",X"FC",X"FE",X"FE",X"FF",
		X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FE",X"FE",X"FC",X"30",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"00",X"00",X"00",X"30",X"FC",X"FE",X"FE",X"FF",
		X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FE",X"FE",X"FC",X"30",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
