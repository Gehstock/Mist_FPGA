library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_PGM is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_PGM is
	type rom is array(0 to  24575) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"3E",X"00",X"32",X"01",X"A8",X"C3",X"45",X"0E",X"77",X"23",X"10",X"FC",X"0D",X"20",X"F9",X"C9",
		X"85",X"6F",X"3E",X"00",X"8C",X"67",X"7E",X"C9",X"77",X"3C",X"23",X"77",X"3C",X"19",X"C9",X"FF",
		X"77",X"23",X"10",X"FC",X"C9",X"FF",X"FF",X"FF",X"87",X"5F",X"16",X"00",X"E1",X"19",X"5E",X"23",
		X"56",X"EB",X"E9",X"FF",X"FF",X"FF",X"FF",X"FF",X"3A",X"A0",X"80",X"E5",X"26",X"80",X"6F",X"CB",
		X"7E",X"28",X"0E",X"72",X"2C",X"73",X"2C",X"7D",X"FE",X"C0",X"30",X"02",X"3E",X"C0",X"32",X"A0",
		X"80",X"E1",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C3",X"69",X"00",X"F5",X"C5",X"D5",X"E5",X"08",X"D9",X"F5",
		X"C5",X"D5",X"E5",X"DD",X"E5",X"FD",X"E5",X"AF",X"32",X"01",X"A8",X"21",X"20",X"80",X"11",X"00",
		X"90",X"01",X"80",X"00",X"ED",X"B0",X"3A",X"00",X"B0",X"3A",X"15",X"80",X"32",X"16",X"80",X"3A",
		X"13",X"80",X"32",X"15",X"80",X"2A",X"10",X"80",X"22",X"13",X"80",X"21",X"12",X"80",X"3A",X"02",
		X"98",X"2F",X"77",X"2B",X"3A",X"01",X"98",X"2F",X"77",X"2B",X"3A",X"00",X"98",X"2F",X"77",X"21",
		X"5F",X"82",X"35",X"CD",X"DF",X"00",X"CD",X"5F",X"36",X"21",X"CB",X"00",X"E5",X"3A",X"05",X"80",
		X"EF",X"8E",X"01",X"8F",X"02",X"6E",X"07",X"AB",X"02",X"C5",X"02",X"FD",X"E1",X"DD",X"E1",X"E1",
		X"D1",X"C1",X"F1",X"D9",X"08",X"E1",X"D1",X"C1",X"3E",X"01",X"32",X"01",X"A8",X"F1",X"C9",X"21",
		X"18",X"80",X"7E",X"A7",X"28",X"03",X"35",X"3E",X"01",X"32",X"02",X"A8",X"21",X"10",X"80",X"7E",
		X"2C",X"2C",X"2C",X"B6",X"2C",X"2C",X"2F",X"A6",X"E6",X"C4",X"28",X"21",X"47",X"E6",X"C0",X"28",
		X"05",X"3E",X"06",X"32",X"18",X"80",X"CD",X"7D",X"03",X"21",X"02",X"80",X"7E",X"FE",X"63",X"38",
		X"02",X"36",X"63",X"3A",X"06",X"80",X"0F",X"38",X"04",X"11",X"01",X"07",X"FF",X"21",X"03",X"80",
		X"5E",X"16",X"06",X"1A",X"1C",X"73",X"23",X"86",X"3D",X"77",X"3A",X"B0",X"80",X"0F",X"D0",X"2A",
		X"B1",X"80",X"7E",X"E6",X"07",X"20",X"1B",X"EB",X"2A",X"B3",X"80",X"7E",X"FE",X"3F",X"28",X"11",
		X"23",X"22",X"B3",X"80",X"D6",X"30",X"2A",X"B5",X"80",X"77",X"01",X"E0",X"FF",X"09",X"22",X"B5",
		X"80",X"EB",X"35",X"C0",X"AF",X"32",X"B0",X"80",X"C9",X"21",X"C0",X"85",X"36",X"00",X"21",X"02",
		X"80",X"78",X"E6",X"84",X"3A",X"00",X"80",X"20",X"13",X"B7",X"28",X"16",X"3D",X"28",X"05",X"3D",
		X"28",X"04",X"18",X"05",X"34",X"34",X"34",X"34",X"34",X"34",X"34",X"C9",X"B7",X"20",X"FB",X"36",
		X"63",X"C9",X"2D",X"34",X"7E",X"FE",X"02",X"D8",X"36",X"00",X"2C",X"C3",X"7A",X"01",X"2A",X"0B",
		X"80",X"06",X"20",X"3E",X"10",X"E7",X"22",X"0B",X"80",X"21",X"08",X"80",X"35",X"C0",X"2D",X"2D",
		X"36",X"00",X"2D",X"36",X"01",X"AF",X"32",X"0A",X"80",X"21",X"CF",X"01",X"CD",X"BF",X"01",X"11",
		X"04",X"06",X"FF",X"11",X"00",X"05",X"FF",X"1E",X"02",X"FF",X"AF",X"32",X"14",X"85",X"C9",X"11",
		X"20",X"80",X"06",X"20",X"EB",X"36",X"00",X"2C",X"1A",X"77",X"2C",X"13",X"10",X"F7",X"C9",X"00",
		X"05",X"00",X"04",X"04",X"01",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",
		X"05",X"00",X"00",X"01",X"01",X"06",X"03",X"03",X"04",X"04",X"04",X"04",X"00",X"00",X"00",X"02",
		X"02",X"02",X"00",X"00",X"00",X"04",X"04",X"04",X"04",X"04",X"06",X"06",X"06",X"06",X"06",X"00",
		X"05",X"02",X"02",X"02",X"02",X"02",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"04",
		X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"06",X"06",X"00",X"06",X"06",X"06",X"00",
		X"05",X"06",X"06",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"06",X"00",
		X"05",X"04",X"04",X"04",X"04",X"04",X"02",X"02",X"02",X"02",X"02",X"02",X"06",X"06",X"06",X"06",
		X"06",X"06",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"06",X"06",X"06",X"06",X"06",X"00",
		X"05",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"02",X"03",X"03",X"04",X"04",X"05",X"05",X"06",
		X"06",X"07",X"07",X"01",X"01",X"02",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"06",X"21",
		X"60",X"07",X"E5",X"3A",X"41",X"85",X"EF",X"B2",X"03",X"E3",X"03",X"18",X"05",X"48",X"05",X"5D",
		X"05",X"83",X"06",X"83",X"06",X"83",X"06",X"9E",X"06",X"DA",X"06",X"3A",X"0A",X"80",X"EF",X"DF",
		X"02",X"8E",X"08",X"A6",X"08",X"30",X"09",X"6C",X"09",X"01",X"03",X"FA",X"09",X"B4",X"0A",X"39",
		X"03",X"F6",X"0B",X"5E",X"0D",X"3A",X"0A",X"80",X"EF",X"DF",X"02",X"8E",X"08",X"EB",X"08",X"30",
		X"09",X"6C",X"09",X"01",X"03",X"00",X"0B",X"1A",X"0B",X"39",X"03",X"F6",X"0B",X"5E",X"0D",X"AF",
		X"32",X"19",X"80",X"21",X"60",X"80",X"06",X"40",X"E7",X"21",X"0A",X"80",X"34",X"2D",X"36",X"20",
		X"21",X"00",X"88",X"22",X"0B",X"80",X"CD",X"8C",X"0A",X"3E",X"01",X"32",X"06",X"80",X"C3",X"7F",
		X"08",X"CD",X"EF",X"18",X"CD",X"A1",X"28",X"CD",X"A2",X"29",X"CD",X"A7",X"30",X"CD",X"97",X"35",
		X"CD",X"28",X"0D",X"CD",X"DA",X"37",X"CD",X"33",X"0D",X"21",X"80",X"83",X"7E",X"0F",X"D8",X"2C",
		X"7E",X"0F",X"D8",X"21",X"80",X"83",X"11",X"81",X"83",X"36",X"00",X"01",X"A0",X"01",X"ED",X"B0",
		X"21",X"0A",X"80",X"36",X"06",X"2D",X"36",X"64",X"C9",X"3A",X"81",X"85",X"EF",X"43",X"03",X"6E",
		X"0B",X"91",X"0B",X"CD",X"EF",X"18",X"CD",X"A1",X"28",X"CD",X"A2",X"29",X"CD",X"C9",X"30",X"CD",
		X"7D",X"0D",X"3A",X"23",X"81",X"3C",X"C0",X"3A",X"12",X"81",X"0F",X"38",X"06",X"3E",X"0A",X"32",
		X"0A",X"80",X"C9",X"32",X"23",X"81",X"21",X"80",X"85",X"36",X"01",X"2C",X"34",X"3E",X"01",X"32",
		X"04",X"A8",X"AF",X"32",X"03",X"A8",X"32",X"19",X"80",X"CD",X"36",X"37",X"C9",X"21",X"C0",X"85",
		X"36",X"00",X"21",X"02",X"80",X"78",X"E6",X"84",X"28",X"15",X"3A",X"00",X"80",X"B7",X"28",X"13",
		X"3D",X"28",X"0E",X"3D",X"28",X"10",X"2D",X"34",X"7E",X"FE",X"04",X"D8",X"36",X"00",X"2C",X"34",
		X"34",X"34",X"C9",X"36",X"63",X"C9",X"2D",X"34",X"7E",X"FE",X"02",X"D8",X"36",X"00",X"2C",X"C3",
		X"A1",X"03",X"3E",X"01",X"32",X"04",X"A8",X"3D",X"32",X"03",X"A8",X"AF",X"32",X"19",X"80",X"21",
		X"20",X"80",X"11",X"21",X"80",X"01",X"7F",X"00",X"36",X"00",X"ED",X"B0",X"21",X"02",X"88",X"22",
		X"0B",X"80",X"21",X"09",X"80",X"36",X"20",X"21",X"41",X"85",X"34",X"AF",X"32",X"06",X"80",X"32",
		X"48",X"85",X"C9",X"3A",X"48",X"85",X"EF",X"F1",X"03",X"4D",X"04",X"6C",X"04",X"A6",X"04",X"C4",
		X"04",X"2A",X"0B",X"80",X"06",X"1E",X"3E",X"10",X"E7",X"11",X"02",X"00",X"19",X"22",X"0B",X"80",
		X"21",X"09",X"80",X"35",X"C0",X"21",X"CF",X"01",X"CD",X"BF",X"01",X"AF",X"32",X"06",X"A8",X"32",
		X"07",X"A8",X"11",X"01",X"07",X"FF",X"11",X"06",X"06",X"FF",X"1E",X"12",X"FF",X"1D",X"FF",X"1E",
		X"0C",X"FF",X"AF",X"21",X"00",X"81",X"06",X"40",X"E7",X"21",X"80",X"83",X"01",X"02",X"A0",X"CF",
		X"21",X"40",X"80",X"06",X"60",X"E7",X"CD",X"B5",X"06",X"CD",X"E5",X"35",X"3E",X"BC",X"DD",X"21",
		X"60",X"82",X"21",X"17",X"88",X"CD",X"AE",X"16",X"21",X"48",X"85",X"34",X"C9",X"CD",X"CC",X"1D",
		X"CD",X"8C",X"1E",X"3A",X"5F",X"82",X"E6",X"03",X"CC",X"DF",X"1E",X"CD",X"A4",X"28",X"CD",X"0B",
		X"05",X"3A",X"83",X"83",X"FE",X"B8",X"D8",X"21",X"48",X"85",X"34",X"C9",X"CD",X"CC",X"1D",X"CD",
		X"DF",X"1E",X"CD",X"A4",X"28",X"CD",X"0B",X"05",X"3A",X"84",X"83",X"FE",X"8E",X"D0",X"21",X"01",
		X"00",X"22",X"C0",X"83",X"7D",X"32",X"C2",X"83",X"21",X"28",X"21",X"7D",X"32",X"CC",X"83",X"7C",
		X"32",X"CD",X"83",X"AF",X"32",X"CE",X"83",X"21",X"17",X"88",X"DD",X"21",X"60",X"82",X"CD",X"87",
		X"20",X"21",X"48",X"85",X"34",X"C9",X"CD",X"CC",X"1D",X"CD",X"74",X"1E",X"CD",X"6C",X"21",X"CD",
		X"A4",X"28",X"CD",X"0B",X"05",X"3A",X"83",X"83",X"FE",X"60",X"D0",X"11",X"0B",X"06",X"FF",X"21",
		X"48",X"85",X"34",X"C9",X"CD",X"CC",X"1D",X"CD",X"A4",X"28",X"CD",X"0B",X"05",X"21",X"40",X"85",
		X"35",X"7E",X"E6",X"1F",X"C0",X"7E",X"B7",X"28",X"10",X"CB",X"BF",X"FE",X"20",X"20",X"05",X"11",
		X"8B",X"06",X"FF",X"C9",X"11",X"0B",X"06",X"FF",X"C9",X"11",X"11",X"06",X"FF",X"AF",X"21",X"40",
		X"80",X"06",X"60",X"E7",X"21",X"41",X"85",X"34",X"21",X"02",X"88",X"11",X"04",X"00",X"3E",X"10",
		X"0E",X"20",X"06",X"1C",X"E7",X"19",X"0D",X"C8",X"18",X"F8",X"C9",X"21",X"4A",X"80",X"06",X"08",
		X"11",X"02",X"00",X"35",X"19",X"10",X"FC",X"C9",X"21",X"4F",X"02",X"CD",X"BF",X"01",X"11",X"86",
		X"06",X"FF",X"11",X"92",X"06",X"FF",X"11",X"8B",X"06",X"FF",X"11",X"8C",X"06",X"FF",X"21",X"50",
		X"85",X"34",X"7E",X"E6",X"03",X"21",X"41",X"85",X"20",X"09",X"34",X"2B",X"36",X"80",X"11",X"00",
		X"02",X"FF",X"C9",X"36",X"07",X"2B",X"34",X"C9",X"21",X"40",X"85",X"35",X"C0",X"21",X"02",X"88",
		X"22",X"0B",X"80",X"21",X"09",X"80",X"36",X"20",X"21",X"41",X"85",X"34",X"C9",X"2A",X"0B",X"80",
		X"06",X"1E",X"3E",X"10",X"E7",X"11",X"02",X"00",X"19",X"22",X"0B",X"80",X"21",X"09",X"80",X"35",
		X"C0",X"21",X"2F",X"02",X"CD",X"BF",X"01",X"11",X"0D",X"06",X"FF",X"11",X"37",X"06",X"FF",X"21",
		X"ED",X"05",X"11",X"60",X"80",X"01",X"20",X"00",X"ED",X"B0",X"3E",X"D3",X"32",X"AA",X"8A",X"3E",
		X"CE",X"32",X"38",X"8B",X"3E",X"CF",X"32",X"39",X"8B",X"3E",X"CD",X"32",X"19",X"8B",X"3E",X"A2",
		X"32",X"3B",X"8B",X"3E",X"A3",X"32",X"3C",X"8B",X"3E",X"A1",X"32",X"1C",X"8B",X"21",X"0D",X"06",
		X"22",X"44",X"85",X"21",X"47",X"8A",X"22",X"46",X"85",X"06",X"08",X"CD",X"CA",X"05",X"10",X"FB",
		X"21",X"40",X"85",X"36",X"78",X"2C",X"3E",X"07",X"77",X"C9",X"C5",X"DD",X"2A",X"44",X"85",X"2A",
		X"46",X"85",X"11",X"E0",X"FF",X"06",X"0D",X"DD",X"7E",X"00",X"77",X"19",X"DD",X"23",X"10",X"F7",
		X"DD",X"22",X"44",X"85",X"11",X"A3",X"01",X"19",X"22",X"46",X"85",X"C1",X"C9",X"30",X"1C",X"06",
		X"32",X"30",X"1E",X"04",X"4A",X"33",X"35",X"02",X"62",X"30",X"1F",X"00",X"7C",X"30",X"13",X"02",
		X"94",X"30",X"10",X"03",X"AA",X"4C",X"1B",X"03",X"32",X"4C",X"3F",X"05",X"93",X"0C",X"0C",X"0C",
		X"0C",X"0C",X"10",X"10",X"03",X"00",X"10",X"20",X"24",X"23",X"0C",X"0C",X"0C",X"0C",X"0C",X"10",
		X"10",X"05",X"00",X"10",X"20",X"24",X"23",X"0C",X"0C",X"0C",X"0C",X"0C",X"10",X"01",X"05",X"00",
		X"10",X"20",X"24",X"23",X"0C",X"0C",X"0C",X"0C",X"0C",X"10",X"10",X"05",X"00",X"10",X"20",X"24",
		X"23",X"0C",X"0C",X"0C",X"0C",X"0C",X"10",X"01",X"00",X"00",X"10",X"20",X"24",X"23",X"0C",X"0C",
		X"0C",X"0C",X"0C",X"10",X"10",X"05",X"00",X"10",X"20",X"24",X"23",X"0C",X"0C",X"0C",X"0C",X"0C",
		X"10",X"01",X"00",X"00",X"10",X"20",X"24",X"23",X"0C",X"0C",X"0C",X"0C",X"0C",X"10",X"1D",X"29",
		X"23",X"24",X"15",X"22",X"29",X"3E",X"10",X"1B",X"1F",X"1E",X"11",X"1D",X"19",X"10",X"10",X"01",
		X"09",X"08",X"01",X"21",X"40",X"85",X"35",X"C0",X"2C",X"34",X"21",X"60",X"80",X"3E",X"10",X"06",
		X"18",X"E7",X"CD",X"6B",X"0A",X"CD",X"8C",X"0A",X"21",X"CF",X"01",X"C3",X"BF",X"01",X"AF",X"21",
		X"00",X"81",X"06",X"40",X"E7",X"21",X"41",X"85",X"34",X"3E",X"01",X"32",X"19",X"80",X"11",X"07",
		X"06",X"FF",X"CD",X"E1",X"35",X"CD",X"7F",X"08",X"CD",X"53",X"09",X"21",X"01",X"00",X"22",X"80",
		X"83",X"22",X"A0",X"83",X"AF",X"32",X"82",X"83",X"3E",X"20",X"32",X"15",X"81",X"21",X"05",X"81",
		X"36",X"FF",X"2C",X"36",X"05",X"11",X"05",X"06",X"FF",X"C9",X"CD",X"EF",X"18",X"3A",X"80",X"83",
		X"B7",X"28",X"63",X"DD",X"21",X"80",X"83",X"3A",X"5F",X"82",X"E6",X"7F",X"20",X"07",X"ED",X"5F",
		X"E6",X"01",X"32",X"50",X"84",X"3A",X"50",X"84",X"B7",X"F5",X"CC",X"DF",X"1E",X"F1",X"C4",X"C7",
		X"1E",X"3A",X"16",X"81",X"47",X"3A",X"84",X"83",X"D6",X"04",X"90",X"E6",X"F8",X"0F",X"0F",X"C6",
		X"C0",X"6F",X"26",X"81",X"2C",X"7E",X"2D",X"86",X"1F",X"47",X"3E",X"C0",X"BD",X"20",X"02",X"2E",
		X"00",X"2D",X"7E",X"2D",X"86",X"1F",X"80",X"1F",X"47",X"3E",X"C0",X"BD",X"20",X"02",X"2E",X"00",
		X"2D",X"7E",X"2D",X"86",X"1F",X"80",X"1F",X"47",X"3A",X"83",X"83",X"B8",X"28",X"08",X"F5",X"D4",
		X"74",X"1E",X"F1",X"DC",X"8C",X"1E",X"CD",X"A1",X"28",X"CD",X"A2",X"29",X"CD",X"A7",X"30",X"CD",
		X"97",X"35",X"21",X"80",X"83",X"7E",X"2C",X"B6",X"0F",X"D8",X"21",X"41",X"85",X"36",X"00",X"C9",
		X"3A",X"02",X"80",X"A7",X"C8",X"21",X"05",X"80",X"34",X"AF",X"32",X"0A",X"80",X"C9",X"21",X"FE",
		X"07",X"E5",X"3A",X"0A",X"80",X"EF",X"7C",X"07",X"AA",X"07",X"F0",X"07",X"AF",X"32",X"19",X"80",
		X"3E",X"01",X"32",X"04",X"A8",X"3D",X"32",X"03",X"A8",X"21",X"EF",X"01",X"CD",X"BF",X"01",X"21",
		X"60",X"80",X"06",X"40",X"AF",X"E7",X"32",X"B0",X"80",X"32",X"06",X"80",X"21",X"02",X"88",X"22",
		X"0B",X"80",X"21",X"09",X"80",X"36",X"10",X"2C",X"34",X"C9",X"2A",X"0B",X"80",X"06",X"1D",X"3E",
		X"10",X"E7",X"11",X"03",X"00",X"19",X"06",X"1D",X"E7",X"19",X"22",X"0B",X"80",X"21",X"09",X"80",
		X"35",X"C0",X"2C",X"34",X"AF",X"32",X"06",X"A8",X"32",X"07",X"A8",X"32",X"0D",X"80",X"11",X"01",
		X"07",X"FF",X"11",X"01",X"06",X"FF",X"1E",X"16",X"FF",X"1C",X"FF",X"3A",X"17",X"80",X"47",X"E6",
		X"0F",X"32",X"58",X"89",X"78",X"E6",X"F0",X"C8",X"0F",X"0F",X"0F",X"0F",X"32",X"78",X"89",X"C9",
		X"3A",X"02",X"80",X"A7",X"C8",X"3D",X"11",X"18",X"06",X"28",X"01",X"1C",X"FF",X"C9",X"3A",X"11",
		X"80",X"CB",X"7F",X"C2",X"3E",X"08",X"CB",X"77",X"C8",X"3A",X"02",X"80",X"FE",X"02",X"D8",X"D6",
		X"02",X"32",X"02",X"80",X"21",X"00",X"01",X"22",X"0D",X"80",X"AF",X"32",X"0A",X"80",X"3E",X"03",
		X"32",X"05",X"80",X"3E",X"01",X"32",X"06",X"80",X"11",X"04",X"06",X"FF",X"CD",X"4D",X"08",X"CD",
		X"1D",X"37",X"11",X"00",X"04",X"FF",X"3A",X"0E",X"80",X"0F",X"D0",X"1C",X"FF",X"C9",X"3A",X"02",
		X"80",X"A7",X"C8",X"3D",X"32",X"02",X"80",X"21",X"00",X"00",X"C3",X"17",X"08",X"AF",X"21",X"00",
		X"81",X"47",X"E7",X"21",X"30",X"82",X"06",X"10",X"E7",X"21",X"60",X"80",X"06",X"40",X"E7",X"21",
		X"60",X"82",X"01",X"02",X"B0",X"CF",X"32",X"19",X"80",X"21",X"00",X"81",X"11",X"01",X"81",X"01",
		X"C0",X"00",X"36",X"00",X"ED",X"B0",X"3A",X"07",X"80",X"32",X"48",X"81",X"32",X"88",X"81",X"21",
		X"C0",X"81",X"11",X"28",X"C8",X"06",X"20",X"72",X"2C",X"73",X"2C",X"10",X"FA",X"C9",X"2A",X"0B",
		X"80",X"06",X"20",X"3E",X"10",X"E7",X"22",X"0B",X"80",X"21",X"09",X"80",X"35",X"C0",X"2C",X"34",
		X"21",X"CF",X"01",X"C3",X"BF",X"01",X"AF",X"32",X"5F",X"82",X"32",X"06",X"A8",X"32",X"07",X"A8",
		X"32",X"0D",X"80",X"21",X"0A",X"80",X"34",X"2D",X"36",X"96",X"3A",X"0E",X"80",X"0F",X"38",X"25",
		X"11",X"00",X"05",X"FF",X"1E",X"02",X"FF",X"14",X"FF",X"1E",X"04",X"FF",X"11",X"03",X"07",X"FF",
		X"1E",X"00",X"FF",X"21",X"40",X"81",X"11",X"00",X"81",X"01",X"40",X"00",X"ED",X"B0",X"2A",X"1D",
		X"81",X"22",X"18",X"81",X"C9",X"11",X"01",X"05",X"FF",X"18",X"D5",X"AF",X"32",X"5F",X"82",X"3A",
		X"0F",X"80",X"0F",X"30",X"08",X"3E",X"01",X"32",X"06",X"A8",X"32",X"07",X"A8",X"3E",X"01",X"32",
		X"0D",X"80",X"21",X"0A",X"80",X"34",X"2D",X"36",X"96",X"11",X"00",X"05",X"FF",X"1C",X"FF",X"1C",
		X"FF",X"11",X"03",X"06",X"FF",X"1C",X"FF",X"11",X"03",X"07",X"FF",X"1E",X"00",X"FF",X"21",X"80",
		X"81",X"11",X"00",X"81",X"01",X"40",X"00",X"ED",X"B0",X"2A",X"1D",X"81",X"22",X"18",X"81",X"C9",
		X"21",X"09",X"80",X"35",X"C0",X"36",X"20",X"2C",X"34",X"11",X"82",X"06",X"FF",X"1E",X"07",X"FF",
		X"CD",X"6B",X"0A",X"CD",X"8C",X"0A",X"CD",X"7F",X"08",X"AF",X"32",X"19",X"80",X"21",X"60",X"80",
		X"06",X"40",X"E7",X"21",X"19",X"88",X"11",X"1C",X"00",X"06",X"20",X"3E",X"36",X"0E",X"39",X"77",
		X"2C",X"71",X"2C",X"71",X"2C",X"71",X"2C",X"71",X"19",X"10",X"F4",X"C9",X"21",X"09",X"80",X"35",
		X"C0",X"36",X"0A",X"2C",X"34",X"3E",X"01",X"32",X"19",X"80",X"21",X"01",X"00",X"22",X"80",X"83",
		X"22",X"A0",X"83",X"AF",X"32",X"82",X"83",X"21",X"08",X"81",X"35",X"11",X"03",X"07",X"FF",X"21",
		X"10",X"81",X"11",X"11",X"81",X"01",X"0C",X"00",X"36",X"00",X"ED",X"B0",X"21",X"24",X"81",X"7E",
		X"B7",X"36",X"00",X"20",X"06",X"CD",X"E1",X"35",X"C3",X"D1",X"09",X"2A",X"20",X"81",X"3A",X"26",
		X"81",X"FE",X"08",X"30",X"0D",X"2B",X"2B",X"2B",X"2B",X"7E",X"3C",X"20",X"07",X"23",X"23",X"C3",
		X"C4",X"09",X"2B",X"2B",X"22",X"20",X"81",X"3E",X"FF",X"CD",X"A5",X"35",X"3E",X"10",X"32",X"26",
		X"81",X"3A",X"1E",X"81",X"D6",X"0A",X"20",X"0A",X"3A",X"25",X"81",X"B7",X"20",X"01",X"3C",X"32",
		X"12",X"81",X"11",X"02",X"07",X"FF",X"3E",X"08",X"32",X"15",X"81",X"3E",X"FF",X"32",X"05",X"81",
		X"3E",X"05",X"32",X"06",X"81",X"11",X"00",X"07",X"FF",X"C9",X"3A",X"08",X"81",X"A7",X"20",X"49",
		X"CD",X"6B",X"0A",X"CD",X"8C",X"0A",X"11",X"02",X"06",X"3A",X"0D",X"80",X"0F",X"30",X"01",X"1C",
		X"FF",X"1E",X"00",X"FF",X"3A",X"1F",X"80",X"47",X"3A",X"3F",X"81",X"B8",X"30",X"0F",X"1E",X"33",
		X"FF",X"1C",X"3A",X"02",X"80",X"B7",X"20",X"01",X"FF",X"1C",X"FF",X"1C",X"FF",X"3E",X"01",X"32",
		X"04",X"A8",X"3D",X"32",X"03",X"A8",X"32",X"C0",X"85",X"32",X"C1",X"85",X"3E",X"09",X"32",X"0A",
		X"80",X"AF",X"32",X"19",X"80",X"CD",X"99",X"37",X"C9",X"21",X"24",X"81",X"3E",X"01",X"77",X"23",
		X"3A",X"12",X"81",X"77",X"3A",X"0E",X"80",X"0F",X"38",X"09",X"21",X"0A",X"80",X"36",X"03",X"2D",
		X"36",X"32",X"C9",X"21",X"0A",X"80",X"34",X"2D",X"36",X"32",X"C9",X"21",X"03",X"88",X"11",X"05",
		X"00",X"0E",X"20",X"3E",X"10",X"06",X"1B",X"77",X"23",X"10",X"FC",X"19",X"0D",X"20",X"F6",X"21",
		X"2A",X"80",X"06",X"19",X"AF",X"77",X"2C",X"77",X"2C",X"10",X"FA",X"C9",X"21",X"60",X"80",X"11",
		X"61",X"80",X"01",X"3F",X"00",X"36",X"00",X"ED",X"B0",X"21",X"80",X"82",X"11",X"81",X"82",X"01",
		X"A0",X"02",X"36",X"00",X"ED",X"B0",X"21",X"60",X"82",X"11",X"61",X"82",X"01",X"1F",X"00",X"36",
		X"00",X"ED",X"B0",X"C9",X"21",X"53",X"0B",X"E5",X"21",X"09",X"80",X"35",X"C0",X"3A",X"08",X"81",
		X"A7",X"20",X"13",X"3A",X"0E",X"80",X"0F",X"38",X"1C",X"3E",X"01",X"32",X"05",X"80",X"AF",X"32",
		X"41",X"85",X"32",X"0D",X"80",X"C9",X"3A",X"88",X"81",X"A7",X"20",X"0F",X"21",X"0A",X"80",X"36",
		X"03",X"2D",X"36",X"01",X"C9",X"3A",X"88",X"81",X"A7",X"28",X"DE",X"21",X"00",X"81",X"11",X"40",
		X"81",X"01",X"40",X"00",X"ED",X"B0",X"AF",X"32",X"0A",X"80",X"3E",X"04",X"32",X"05",X"80",X"C9",
		X"3A",X"08",X"81",X"A7",X"CA",X"00",X"0A",X"21",X"24",X"81",X"3E",X"01",X"77",X"23",X"3A",X"12",
		X"81",X"77",X"21",X"0A",X"80",X"34",X"2D",X"36",X"64",X"C9",X"21",X"53",X"0B",X"E5",X"21",X"09",
		X"80",X"35",X"C0",X"3A",X"08",X"81",X"A7",X"20",X"06",X"3A",X"48",X"81",X"A7",X"28",X"9A",X"3A",
		X"48",X"81",X"A7",X"20",X"09",X"21",X"0A",X"80",X"36",X"03",X"2D",X"36",X"01",X"C9",X"21",X"00",
		X"81",X"11",X"80",X"81",X"01",X"40",X"00",X"ED",X"B0",X"AF",X"32",X"0A",X"80",X"3E",X"03",X"32",
		X"05",X"80",X"C9",X"3A",X"0E",X"80",X"0F",X"D2",X"FE",X"07",X"21",X"48",X"81",X"3A",X"0D",X"80",
		X"0F",X"38",X"03",X"21",X"88",X"81",X"3A",X"08",X"81",X"B6",X"CA",X"FE",X"07",X"C9",X"21",X"06",
		X"81",X"34",X"21",X"80",X"85",X"35",X"C0",X"36",X"AA",X"2C",X"34",X"CD",X"7F",X"0A",X"11",X"08",
		X"06",X"FF",X"1C",X"FF",X"1C",X"FF",X"C9",X"21",X"6F",X"02",X"CD",X"BF",X"01",X"CD",X"7F",X"08",
		X"C9",X"21",X"06",X"81",X"34",X"CD",X"EF",X"18",X"CD",X"A4",X"28",X"CD",X"A2",X"29",X"CD",X"0B",
		X"05",X"11",X"58",X"0D",X"21",X"18",X"81",X"73",X"23",X"72",X"3A",X"5F",X"82",X"E6",X"03",X"C0",
		X"3A",X"80",X"85",X"FE",X"40",X"CC",X"1D",X"37",X"21",X"80",X"85",X"35",X"C0",X"21",X"08",X"81",
		X"34",X"21",X"00",X"81",X"34",X"11",X"00",X"07",X"FF",X"AF",X"32",X"5F",X"82",X"21",X"0A",X"80",
		X"36",X"03",X"2D",X"36",X"32",X"AF",X"32",X"1E",X"81",X"21",X"CF",X"01",X"CD",X"BF",X"01",X"21",
		X"08",X"81",X"34",X"CD",X"1C",X"38",X"AF",X"32",X"23",X"81",X"21",X"6C",X"80",X"11",X"6D",X"80",
		X"01",X"33",X"00",X"C3",X"95",X"0A",X"21",X"53",X"0B",X"E5",X"3A",X"C1",X"85",X"EF",X"04",X"0C",
		X"A5",X"0C",X"C4",X"0C",X"3A",X"1F",X"80",X"47",X"3A",X"3F",X"81",X"B8",X"30",X"4D",X"3A",X"02",
		X"80",X"B7",X"28",X"2F",X"11",X"B4",X"06",X"FF",X"3A",X"0D",X"80",X"B7",X"20",X"1C",X"3A",X"10",
		X"80",X"E6",X"0A",X"20",X"53",X"3A",X"C0",X"85",X"47",X"E6",X"07",X"20",X"29",X"78",X"11",X"35",
		X"06",X"E6",X"1F",X"20",X"02",X"CB",X"FB",X"FF",X"18",X"1C",X"3A",X"11",X"80",X"E6",X"0C",X"20",
		X"37",X"18",X"E2",X"3A",X"C0",X"85",X"47",X"E6",X"07",X"20",X"0B",X"78",X"11",X"34",X"06",X"E6",
		X"1F",X"20",X"02",X"CB",X"FB",X"FF",X"3A",X"5F",X"82",X"0F",X"D8",X"21",X"C0",X"85",X"35",X"C0",
		X"2C",X"34",X"11",X"80",X"06",X"FF",X"1E",X"82",X"FF",X"1E",X"B3",X"FF",X"1C",X"FF",X"1C",X"FF",
		X"1C",X"FF",X"21",X"4F",X"02",X"C3",X"BF",X"01",X"CD",X"D2",X"0C",X"3A",X"07",X"80",X"32",X"08",
		X"81",X"3E",X"06",X"32",X"0A",X"80",X"21",X"A2",X"80",X"3A",X"0D",X"80",X"B7",X"28",X"03",X"23",
		X"23",X"23",X"AF",X"32",X"07",X"81",X"06",X"03",X"77",X"23",X"10",X"FC",X"21",X"02",X"80",X"35",
		X"21",X"3F",X"81",X"34",X"C9",X"CD",X"D2",X"0C",X"7D",X"FE",X"0A",X"28",X"0B",X"87",X"87",X"5F",
		X"16",X"00",X"21",X"2F",X"80",X"19",X"36",X"00",X"11",X"00",X"02",X"FF",X"21",X"C0",X"85",X"36",
		X"80",X"2C",X"34",X"C9",X"21",X"C0",X"85",X"35",X"C0",X"21",X"0A",X"80",X"36",X"07",X"2D",X"36",
		X"64",X"C9",X"01",X"1E",X"00",X"11",X"03",X"00",X"6A",X"DD",X"21",X"A2",X"80",X"3A",X"0D",X"80",
		X"0F",X"30",X"02",X"DD",X"19",X"FD",X"21",X"00",X"82",X"DD",X"7E",X"02",X"FD",X"BE",X"02",X"20",
		X"0F",X"DD",X"7E",X"01",X"FD",X"BE",X"01",X"20",X"07",X"DD",X"7E",X"00",X"FD",X"BE",X"00",X"C8",
		X"30",X"09",X"FD",X"19",X"2C",X"0D",X"0D",X"0D",X"C8",X"18",X"DE",X"7D",X"21",X"1D",X"82",X"11",
		X"20",X"82",X"ED",X"B8",X"6F",X"DD",X"7E",X"00",X"FD",X"77",X"00",X"DD",X"7E",X"01",X"FD",X"77",
		X"01",X"DD",X"7E",X"02",X"FD",X"77",X"02",X"C9",X"3A",X"5F",X"82",X"E6",X"3F",X"C0",X"11",X"0C",
		X"03",X"FF",X"C9",X"3A",X"07",X"81",X"A7",X"C0",X"21",X"A4",X"80",X"3A",X"0D",X"80",X"0F",X"30",
		X"03",X"21",X"A7",X"80",X"7E",X"A7",X"C8",X"CD",X"1C",X"38",X"21",X"08",X"81",X"34",X"11",X"03",
		X"07",X"FF",X"3E",X"01",X"32",X"07",X"81",X"C9",X"C8",X"36",X"C8",X"36",X"00",X"00",X"21",X"06",
		X"81",X"34",X"3A",X"23",X"81",X"B7",X"20",X"76",X"CD",X"EF",X"18",X"CD",X"A1",X"28",X"CD",X"A2",
		X"29",X"CD",X"E1",X"30",X"CD",X"28",X"0D",X"CD",X"0B",X"38",X"CD",X"33",X"0D",X"11",X"58",X"0D",
		X"21",X"18",X"81",X"73",X"23",X"72",X"21",X"80",X"83",X"7E",X"0F",X"D2",X"1F",X"03",X"21",X"22",
		X"81",X"35",X"CA",X"9D",X"0D",X"3A",X"5F",X"82",X"CB",X"47",X"C0",X"34",X"C9",X"34",X"23",X"35",
		X"3A",X"16",X"81",X"E6",X"07",X"28",X"02",X"34",X"C9",X"3A",X"12",X"81",X"FE",X"41",X"C8",X"AF",
		X"32",X"16",X"81",X"06",X"19",X"21",X"2A",X"80",X"77",X"2C",X"2C",X"10",X"FB",X"3A",X"1E",X"81",
		X"FE",X"0A",X"28",X"11",X"11",X"25",X"06",X"FF",X"CD",X"27",X"37",X"3A",X"1E",X"81",X"C6",X"26",
		X"16",X"06",X"5F",X"FF",X"C9",X"11",X"31",X"06",X"FF",X"1C",X"FF",X"C3",X"CB",X"0D",X"CD",X"F2",
		X"18",X"CD",X"A4",X"28",X"CD",X"A2",X"29",X"CD",X"E1",X"30",X"CD",X"28",X"0D",X"CD",X"0B",X"38",
		X"CD",X"33",X"0D",X"CD",X"0B",X"05",X"11",X"58",X"0D",X"21",X"18",X"81",X"73",X"23",X"72",X"21",
		X"80",X"83",X"7E",X"0F",X"D2",X"1F",X"03",X"16",X"06",X"21",X"23",X"81",X"35",X"28",X"12",X"3E",
		X"1F",X"A6",X"C0",X"3A",X"1E",X"81",X"C6",X"26",X"5F",X"CB",X"6E",X"20",X"02",X"CB",X"FB",X"FF",
		X"C9",X"21",X"05",X"81",X"3E",X"30",X"86",X"30",X"02",X"3E",X"FF",X"77",X"21",X"1E",X"81",X"34",
		X"7E",X"FE",X"0A",X"38",X"07",X"3E",X"01",X"32",X"12",X"81",X"36",X"0A",X"CD",X"E1",X"35",X"3E",
		X"05",X"32",X"0A",X"80",X"C9",X"3A",X"00",X"60",X"FE",X"55",X"CA",X"01",X"60",X"21",X"00",X"80",
		X"11",X"01",X"80",X"01",X"00",X"08",X"36",X"00",X"ED",X"B0",X"3E",X"9B",X"32",X"03",X"98",X"3E",
		X"88",X"32",X"03",X"A0",X"3E",X"08",X"32",X"42",X"82",X"32",X"01",X"A0",X"31",X"00",X"88",X"21",
		X"C0",X"80",X"06",X"40",X"3E",X"FF",X"E7",X"21",X"43",X"82",X"06",X"1C",X"E7",X"21",X"43",X"43",
		X"22",X"40",X"82",X"3A",X"00",X"B0",X"AF",X"32",X"01",X"A8",X"32",X"05",X"B0",X"32",X"06",X"A8",
		X"32",X"07",X"A8",X"21",X"C0",X"C0",X"22",X"A0",X"80",X"3C",X"32",X"04",X"A8",X"21",X"00",X"88",
		X"22",X"0B",X"80",X"3E",X"20",X"32",X"08",X"80",X"3E",X"10",X"32",X"17",X"80",X"3A",X"02",X"98",
		X"0F",X"47",X"E6",X"03",X"32",X"00",X"80",X"78",X"0F",X"0F",X"E6",X"01",X"32",X"0F",X"80",X"3A",
		X"01",X"98",X"47",X"CB",X"48",X"3E",X"03",X"28",X"02",X"3E",X"04",X"32",X"07",X"80",X"3E",X"00",
		X"CB",X"40",X"28",X"02",X"3E",X"04",X"32",X"1F",X"80",X"CD",X"9D",X"36",X"AF",X"3D",X"20",X"FD",
		X"CD",X"AC",X"36",X"21",X"00",X"90",X"01",X"00",X"01",X"16",X"00",X"72",X"23",X"0B",X"78",X"B1",
		X"20",X"F9",X"16",X"3F",X"21",X"00",X"88",X"01",X"00",X"08",X"72",X"3A",X"00",X"B0",X"23",X"0B",
		X"78",X"B1",X"20",X"F6",X"CD",X"30",X"0F",X"30",X"22",X"CD",X"30",X"0F",X"30",X"1D",X"3E",X"01",
		X"32",X"01",X"A8",X"21",X"00",X"82",X"06",X"0A",X"36",X"00",X"2C",X"36",X"00",X"2C",X"36",X"01",
		X"2C",X"10",X"F5",X"21",X"AA",X"80",X"36",X"01",X"C3",X"3F",X"0F",X"3A",X"00",X"B0",X"18",X"FB",
		X"0B",X"3A",X"00",X"B0",X"3A",X"01",X"98",X"07",X"D0",X"78",X"B1",X"20",X"F3",X"37",X"C9",X"26",
		X"80",X"3A",X"A1",X"80",X"6F",X"7E",X"87",X"30",X"05",X"CD",X"82",X"0F",X"18",X"F1",X"E6",X"1F",
		X"4F",X"06",X"00",X"36",X"FF",X"23",X"5E",X"36",X"FF",X"2C",X"7D",X"FE",X"C0",X"30",X"02",X"3E",
		X"C0",X"32",X"A1",X"80",X"7B",X"21",X"72",X"0F",X"09",X"5E",X"23",X"56",X"21",X"3F",X"0F",X"E5",
		X"EB",X"E9",X"E8",X"0F",X"E9",X"0F",X"EA",X"0F",X"48",X"10",X"DE",X"10",X"FA",X"10",X"41",X"11",
		X"85",X"15",X"3A",X"5F",X"82",X"47",X"E6",X"0F",X"CA",X"A1",X"0F",X"21",X"19",X"80",X"CB",X"46",
		X"C8",X"E6",X"03",X"CA",X"DB",X"16",X"3D",X"CA",X"89",X"16",X"3D",X"CA",X"D2",X"15",X"C3",X"89",
		X"16",X"11",X"E0",X"FF",X"21",X"E0",X"88",X"3A",X"0E",X"80",X"A7",X"28",X"22",X"36",X"02",X"CD",
		X"D9",X"0F",X"21",X"40",X"8B",X"CD",X"D7",X"0F",X"3A",X"0D",X"80",X"A7",X"21",X"40",X"8B",X"28",
		X"03",X"21",X"E0",X"88",X"CB",X"60",X"C8",X"3A",X"06",X"80",X"0F",X"D0",X"C3",X"E0",X"0F",X"21",
		X"E0",X"88",X"CD",X"E0",X"0F",X"18",X"DB",X"36",X"01",X"19",X"36",X"25",X"19",X"36",X"20",X"C9",
		X"3E",X"10",X"77",X"19",X"77",X"19",X"77",X"C9",X"C9",X"C9",X"3E",X"1A",X"06",X"0B",X"F5",X"C5",
		X"CD",X"41",X"11",X"C1",X"F1",X"3C",X"10",X"F6",X"21",X"87",X"89",X"11",X"20",X"00",X"06",X"0A",
		X"DD",X"21",X"00",X"82",X"DD",X"7E",X"00",X"4F",X"E6",X"0F",X"77",X"19",X"79",X"0F",X"0F",X"0F",
		X"0F",X"E6",X"0F",X"77",X"19",X"DD",X"23",X"DD",X"7E",X"00",X"4F",X"E6",X"0F",X"77",X"19",X"79",
		X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"77",X"19",X"DD",X"23",X"DD",X"7E",X"00",X"4F",X"E6",X"0F",
		X"77",X"19",X"79",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"28",X"01",X"77",X"11",X"62",X"FF",X"19",
		X"11",X"20",X"00",X"DD",X"23",X"10",X"BD",X"C9",X"4F",X"3A",X"06",X"80",X"0F",X"D0",X"79",X"A7",
		X"28",X"48",X"4F",X"CD",X"A5",X"10",X"87",X"81",X"4F",X"06",X"00",X"21",X"B4",X"10",X"09",X"A7",
		X"06",X"03",X"1A",X"8E",X"27",X"12",X"13",X"23",X"10",X"F8",X"D5",X"3A",X"0D",X"80",X"0F",X"30",
		X"02",X"3E",X"01",X"CD",X"FA",X"10",X"D1",X"1B",X"21",X"AA",X"80",X"06",X"03",X"1A",X"BE",X"D8",
		X"20",X"05",X"1B",X"2B",X"10",X"F7",X"C9",X"CD",X"A5",X"10",X"21",X"A8",X"80",X"06",X"03",X"1A",
		X"77",X"13",X"23",X"10",X"FA",X"3E",X"02",X"C3",X"FA",X"10",X"CD",X"A5",X"10",X"21",X"AB",X"80",
		X"A7",X"06",X"03",X"18",X"BD",X"F5",X"3A",X"0D",X"80",X"11",X"A2",X"80",X"0F",X"30",X"03",X"11",
		X"A5",X"80",X"F1",X"C9",X"00",X"00",X"00",X"30",X"00",X"00",X"50",X"01",X"00",X"50",X"00",X"00",
		X"50",X"00",X"00",X"00",X"01",X"00",X"00",X"02",X"00",X"00",X"03",X"00",X"00",X"01",X"00",X"00",
		X"02",X"00",X"50",X"00",X"00",X"00",X"02",X"00",X"10",X"00",X"00",X"00",X"08",X"00",X"F5",X"21",
		X"A2",X"80",X"A7",X"28",X"09",X"21",X"A5",X"80",X"3D",X"28",X"03",X"21",X"A8",X"80",X"36",X"00",
		X"23",X"36",X"00",X"23",X"36",X"00",X"F1",X"C3",X"FA",X"10",X"21",X"A4",X"80",X"DD",X"21",X"81",
		X"8B",X"A7",X"28",X"11",X"21",X"A7",X"80",X"DD",X"21",X"21",X"89",X"3D",X"28",X"07",X"21",X"AA",
		X"80",X"DD",X"21",X"41",X"8A",X"11",X"E0",X"FF",X"06",X"03",X"0E",X"04",X"7E",X"0F",X"0F",X"0F",
		X"0F",X"CD",X"2C",X"11",X"7E",X"CD",X"2C",X"11",X"2B",X"10",X"F1",X"C9",X"E6",X"0F",X"28",X"08",
		X"0E",X"00",X"DD",X"77",X"00",X"DD",X"19",X"C9",X"79",X"A7",X"28",X"F6",X"3E",X"10",X"0D",X"18",
		X"F1",X"87",X"F5",X"21",X"AE",X"11",X"E6",X"7F",X"5F",X"16",X"00",X"19",X"5E",X"23",X"56",X"EB",
		X"5E",X"23",X"56",X"23",X"EB",X"01",X"E0",X"FF",X"F1",X"38",X"0E",X"FA",X"73",X"11",X"1A",X"FE",
		X"3F",X"C8",X"D6",X"30",X"77",X"13",X"09",X"18",X"F5",X"1A",X"FE",X"3F",X"C8",X"36",X"10",X"13",
		X"09",X"18",X"F6",X"22",X"B5",X"80",X"ED",X"53",X"B3",X"80",X"EB",X"7B",X"E6",X"1F",X"47",X"87",
		X"C6",X"20",X"6F",X"26",X"80",X"22",X"B1",X"80",X"CB",X"3B",X"CB",X"3B",X"7A",X"E6",X"03",X"0F",
		X"0F",X"B3",X"E6",X"F8",X"4F",X"21",X"00",X"88",X"78",X"85",X"6F",X"11",X"20",X"00",X"43",X"36",
		X"10",X"19",X"10",X"FB",X"2A",X"B1",X"80",X"71",X"3E",X"01",X"32",X"B0",X"80",X"C9",X"1E",X"12",
		X"2B",X"12",X"3F",X"12",X"4C",X"12",X"59",X"12",X"66",X"12",X"7E",X"12",X"94",X"12",X"9B",X"12",
		X"AF",X"12",X"CC",X"12",X"E9",X"12",X"FC",X"12",X"0E",X"13",X"20",X"13",X"20",X"13",X"20",X"13",
		X"20",X"13",X"33",X"13",X"47",X"13",X"58",X"13",X"69",X"13",X"7A",X"13",X"8E",X"13",X"98",X"13",
		X"AA",X"13",X"BF",X"13",X"D3",X"13",X"E6",X"13",X"F9",X"13",X"0C",X"14",X"1F",X"14",X"32",X"14",
		X"45",X"14",X"58",X"14",X"6B",X"14",X"7E",X"14",X"92",X"14",X"A2",X"14",X"A9",X"14",X"B0",X"14",
		X"B7",X"14",X"BE",X"14",X"C5",X"14",X"CC",X"14",X"D3",X"14",X"DA",X"14",X"E1",X"14",X"E9",X"14",
		X"F6",X"14",X"FE",X"14",X"12",X"15",X"23",X"15",X"40",X"15",X"5C",X"15",X"72",X"15",X"89",X"8A",
		X"47",X"41",X"4D",X"45",X"40",X"40",X"4F",X"56",X"45",X"52",X"3F",X"F1",X"8A",X"50",X"55",X"53",
		X"48",X"40",X"53",X"54",X"41",X"52",X"54",X"40",X"42",X"55",X"54",X"54",X"4F",X"4E",X"3F",X"87",
		X"8A",X"50",X"4C",X"41",X"59",X"45",X"52",X"40",X"4F",X"4E",X"45",X"3F",X"87",X"8A",X"50",X"4C",
		X"41",X"59",X"45",X"52",X"40",X"54",X"57",X"4F",X"3F",X"80",X"8A",X"48",X"49",X"47",X"48",X"40",
		X"53",X"43",X"4F",X"52",X"45",X"3F",X"9F",X"8B",X"40",X"43",X"52",X"45",X"44",X"49",X"54",X"40",
		X"40",X"30",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"3F",X"07",X"8B",
		X"49",X"4E",X"56",X"41",X"44",X"45",X"40",X"54",X"48",X"45",X"40",X"42",X"41",X"53",X"45",X"40",
		X"41",X"4E",X"44",X"3F",X"5E",X"8B",X"46",X"55",X"45",X"4C",X"3F",X"CC",X"8A",X"43",X"4F",X"4E",
		X"47",X"52",X"41",X"54",X"55",X"4C",X"41",X"54",X"49",X"4F",X"4E",X"53",X"40",X"02",X"3F",X"6E",
		X"8B",X"59",X"4F",X"55",X"40",X"43",X"4F",X"4D",X"50",X"4C",X"45",X"54",X"45",X"44",X"40",X"59",
		X"4F",X"55",X"52",X"40",X"44",X"55",X"54",X"49",X"45",X"53",X"C0",X"3F",X"70",X"8B",X"47",X"4F",
		X"4F",X"44",X"40",X"4C",X"55",X"43",X"4B",X"40",X"4E",X"45",X"58",X"54",X"40",X"54",X"49",X"4D",
		X"45",X"40",X"41",X"47",X"41",X"49",X"4E",X"C0",X"3F",X"D3",X"8A",X"42",X"4F",X"4E",X"55",X"53",
		X"40",X"43",X"48",X"4F",X"50",X"50",X"45",X"52",X"40",X"3F",X"02",X"3F",X"C4",X"8A",X"5B",X"40",
		X"53",X"55",X"50",X"45",X"52",X"40",X"43",X"4F",X"42",X"52",X"41",X"40",X"5B",X"3F",X"C4",X"8A",
		X"5B",X"40",X"53",X"43",X"4F",X"52",X"45",X"40",X"54",X"41",X"42",X"4C",X"45",X"40",X"5B",X"3F",
		X"BD",X"8A",X"40",X"6E",X"40",X"4B",X"4F",X"4E",X"41",X"4D",X"49",X"40",X"40",X"31",X"39",X"38",
		X"31",X"40",X"3F",X"E9",X"8A",X"43",X"41",X"52",X"52",X"59",X"40",X"41",X"57",X"41",X"59",X"40",
		X"42",X"4F",X"4F",X"54",X"59",X"C0",X"3F",X"D5",X"8A",X"32",X"40",X"43",X"4F",X"49",X"4E",X"53",
		X"40",X"31",X"40",X"50",X"4C",X"41",X"59",X"3F",X"D5",X"8A",X"33",X"40",X"43",X"4F",X"49",X"4E",
		X"53",X"40",X"31",X"40",X"50",X"4C",X"41",X"59",X"3F",X"D5",X"8A",X"31",X"40",X"43",X"4F",X"49",
		X"4E",X"40",X"40",X"32",X"40",X"50",X"4C",X"41",X"59",X"3F",X"B8",X"8B",X"42",X"4F",X"4E",X"55",
		X"53",X"40",X"43",X"48",X"4F",X"50",X"50",X"45",X"52",X"40",X"46",X"4F",X"52",X"3F",X"38",X"89",
		X"30",X"30",X"30",X"40",X"50",X"54",X"53",X"3F",X"D4",X"8A",X"4F",X"4E",X"45",X"40",X"50",X"4C",
		X"41",X"59",X"45",X"52",X"40",X"4F",X"4E",X"4C",X"59",X"3F",X"F4",X"8A",X"4F",X"4E",X"45",X"40",
		X"4F",X"52",X"40",X"54",X"57",X"4F",X"40",X"50",X"4C",X"41",X"59",X"45",X"52",X"53",X"3F",X"04",
		X"8B",X"5B",X"40",X"53",X"43",X"4F",X"52",X"45",X"40",X"52",X"41",X"4E",X"4B",X"49",X"4E",X"47",
		X"40",X"5B",X"3F",X"E7",X"8A",X"31",X"53",X"54",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",
		X"40",X"40",X"50",X"54",X"53",X"3F",X"E9",X"8A",X"32",X"4E",X"44",X"40",X"40",X"40",X"40",X"40",
		X"40",X"40",X"40",X"40",X"40",X"50",X"54",X"53",X"3F",X"EB",X"8A",X"33",X"52",X"44",X"40",X"40",
		X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"50",X"54",X"53",X"3F",X"ED",X"8A",X"34",X"54",
		X"48",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"50",X"54",X"53",X"3F",X"EF",
		X"8A",X"35",X"54",X"48",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"50",X"54",
		X"53",X"3F",X"F1",X"8A",X"36",X"54",X"48",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",
		X"40",X"50",X"54",X"53",X"3F",X"F3",X"8A",X"37",X"54",X"48",X"40",X"40",X"40",X"40",X"40",X"40",
		X"40",X"40",X"40",X"40",X"50",X"54",X"53",X"3F",X"F5",X"8A",X"38",X"54",X"48",X"40",X"40",X"40",
		X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"50",X"54",X"53",X"3F",X"F7",X"8A",X"39",X"54",X"48",
		X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"50",X"54",X"53",X"3F",X"19",X"8B",
		X"31",X"30",X"54",X"48",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"50",X"54",
		X"53",X"3F",X"74",X"8A",X"4D",X"49",X"4C",X"45",X"53",X"40",X"43",X"4C",X"45",X"41",X"52",X"45",
		X"44",X"3F",X"14",X"8B",X"31",X"30",X"30",X"30",X"3F",X"14",X"8B",X"32",X"30",X"30",X"30",X"3F",
		X"14",X"8B",X"33",X"30",X"30",X"30",X"3F",X"14",X"8B",X"34",X"30",X"30",X"30",X"3F",X"14",X"8B",
		X"35",X"30",X"30",X"30",X"3F",X"14",X"8B",X"36",X"30",X"30",X"30",X"3F",X"14",X"8B",X"37",X"30",
		X"30",X"30",X"3F",X"14",X"8B",X"38",X"30",X"30",X"30",X"3F",X"14",X"8B",X"39",X"30",X"30",X"30",
		X"3F",X"34",X"8B",X"31",X"30",X"30",X"30",X"30",X"3F",X"2F",X"8A",X"44",X"45",X"53",X"54",X"52",
		X"4F",X"59",X"45",X"44",X"C0",X"3F",X"0F",X"8B",X"42",X"4F",X"4F",X"54",X"59",X"3F",X"12",X"8B",
		X"43",X"48",X"41",X"4C",X"4C",X"45",X"4E",X"47",X"45",X"40",X"41",X"47",X"41",X"49",X"4E",X"40",
		X"02",X"3F",X"55",X"8B",X"49",X"46",X"40",X"59",X"4F",X"55",X"40",X"57",X"49",X"53",X"48",X"40",
		X"54",X"4F",X"3F",X"6E",X"8B",X"49",X"4E",X"53",X"45",X"52",X"54",X"40",X"41",X"44",X"44",X"49",
		X"54",X"49",X"4F",X"4E",X"41",X"4C",X"40",X"43",X"4F",X"49",X"4E",X"40",X"41",X"4E",X"44",X"3F",
		X"71",X"8B",X"50",X"55",X"53",X"48",X"40",X"54",X"48",X"45",X"40",X"44",X"49",X"53",X"43",X"48",
		X"41",X"52",X"47",X"45",X"40",X"42",X"55",X"54",X"54",X"4F",X"4E",X"3F",X"17",X"8B",X"43",X"4F",
		X"4E",X"54",X"49",X"4E",X"55",X"45",X"40",X"59",X"4F",X"55",X"52",X"40",X"47",X"41",X"4D",X"45",
		X"C0",X"3F",X"BF",X"8A",X"40",X"6E",X"40",X"4B",X"4F",X"4E",X"41",X"4D",X"49",X"40",X"40",X"31",
		X"39",X"38",X"31",X"40",X"3F",X"A7",X"CA",X"7B",X"17",X"3D",X"CA",X"94",X"15",X"3D",X"CA",X"99",
		X"17",X"C3",X"56",X"17",X"3E",X"05",X"CD",X"41",X"11",X"3A",X"02",X"80",X"FE",X"63",X"38",X"02",
		X"3E",X"63",X"CD",X"B8",X"15",X"47",X"E6",X"F0",X"28",X"07",X"0F",X"0F",X"0F",X"0F",X"32",X"9F",
		X"8A",X"78",X"E6",X"0F",X"32",X"7F",X"8A",X"C9",X"47",X"E6",X"0F",X"C6",X"00",X"27",X"4F",X"78",
		X"E6",X"F0",X"28",X"0B",X"0F",X"0F",X"0F",X"0F",X"47",X"AF",X"C6",X"16",X"27",X"10",X"FB",X"81",
		X"27",X"C9",X"3A",X"10",X"81",X"0F",X"D0",X"3A",X"30",X"82",X"0F",X"D0",X"2A",X"35",X"82",X"7D",
		X"E6",X"E0",X"6F",X"11",X"05",X"00",X"19",X"3E",X"10",X"06",X"19",X"E7",X"11",X"07",X"00",X"19",
		X"06",X"19",X"E7",X"DD",X"21",X"30",X"82",X"DD",X"7E",X"01",X"DD",X"6E",X"02",X"DD",X"66",X"03",
		X"77",X"57",X"7D",X"E6",X"1F",X"47",X"3E",X"1D",X"90",X"28",X"0E",X"47",X"0E",X"39",X"7A",X"FE",
		X"2B",X"30",X"02",X"0E",X"3D",X"23",X"71",X"10",X"FC",X"DD",X"7E",X"04",X"DD",X"6E",X"05",X"DD",
		X"66",X"06",X"77",X"57",X"7D",X"E6",X"1F",X"47",X"3E",X"1D",X"90",X"28",X"0E",X"47",X"0E",X"39",
		X"7A",X"FE",X"2B",X"30",X"02",X"0E",X"D0",X"23",X"71",X"10",X"FC",X"DD",X"36",X"00",X"00",X"DD",
		X"CB",X"08",X"46",X"C8",X"DD",X"7E",X"09",X"DD",X"6E",X"0A",X"DD",X"66",X"0B",X"77",X"57",X"7D",
		X"E6",X"1F",X"D6",X"05",X"28",X"0E",X"47",X"0E",X"39",X"7A",X"FE",X"2B",X"30",X"02",X"0E",X"D0",
		X"2B",X"71",X"10",X"FC",X"DD",X"7E",X"0C",X"DD",X"6E",X"0D",X"DD",X"66",X"0E",X"77",X"57",X"7D",
		X"E6",X"1F",X"D6",X"05",X"28",X"0E",X"47",X"0E",X"39",X"7A",X"FE",X"2B",X"30",X"02",X"0E",X"3D",
		X"2B",X"71",X"10",X"FC",X"DD",X"36",X"08",X"00",X"C9",X"11",X"04",X"00",X"06",X"08",X"DD",X"21",
		X"60",X"82",X"D9",X"CD",X"9C",X"16",X"D9",X"DD",X"19",X"10",X"F7",X"C9",X"DD",X"CB",X"00",X"46",
		X"C8",X"DD",X"7E",X"01",X"87",X"87",X"38",X"18",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"77",X"3C",
		X"23",X"77",X"3C",X"11",X"1F",X"00",X"19",X"77",X"3C",X"23",X"77",X"DD",X"36",X"00",X"00",X"C9",
		X"DD",X"6E",X"02",X"DD",X"66",X"03",X"36",X"10",X"23",X"36",X"44",X"11",X"1F",X"00",X"19",X"36",
		X"10",X"23",X"DD",X"7E",X"01",X"77",X"DD",X"36",X"00",X"00",X"C9",X"3A",X"05",X"81",X"0F",X"4F",
		X"E6",X"78",X"0F",X"0F",X"0F",X"47",X"3E",X"0F",X"90",X"21",X"BE",X"8A",X"11",X"E0",X"FF",X"04",
		X"05",X"28",X"05",X"36",X"CB",X"19",X"10",X"FB",X"47",X"79",X"E6",X"07",X"D9",X"21",X"10",X"17",
		X"5F",X"16",X"00",X"19",X"7E",X"D9",X"77",X"04",X"05",X"C8",X"19",X"36",X"3C",X"10",X"FB",X"C9",
		X"3C",X"C4",X"C5",X"C6",X"C7",X"C8",X"C9",X"CA",X"CD",X"DB",X"16",X"3A",X"01",X"81",X"21",X"64",
		X"8B",X"11",X"E0",X"FF",X"47",X"3E",X"18",X"90",X"04",X"05",X"28",X"05",X"36",X"0C",X"19",X"10",
		X"FB",X"47",X"A7",X"28",X"05",X"36",X"10",X"19",X"10",X"FB",X"3A",X"02",X"81",X"21",X"63",X"8B",
		X"47",X"3E",X"18",X"90",X"04",X"05",X"28",X"05",X"36",X"0D",X"19",X"10",X"FB",X"47",X"A7",X"C8",
		X"36",X"10",X"19",X"10",X"FB",X"C9",X"21",X"BF",X"8B",X"11",X"E0",X"FF",X"06",X"0C",X"36",X"10",
		X"19",X"10",X"FB",X"21",X"BF",X"8B",X"3A",X"08",X"81",X"A7",X"C8",X"FE",X"07",X"38",X"02",X"3E",
		X"06",X"47",X"36",X"0A",X"19",X"36",X"0B",X"19",X"10",X"F8",X"C9",X"3A",X"00",X"81",X"E6",X"0F",
		X"3C",X"47",X"3E",X"10",X"90",X"21",X"5F",X"88",X"11",X"20",X"00",X"36",X"D1",X"19",X"10",X"FB",
		X"A7",X"C8",X"36",X"10",X"19",X"3D",X"20",X"FA",X"C9",X"DD",X"21",X"63",X"8B",X"11",X"E0",X"FF",
		X"21",X"E6",X"17",X"06",X"18",X"7E",X"DD",X"77",X"00",X"23",X"DD",X"19",X"10",X"F7",X"21",X"64",
		X"8B",X"11",X"E0",X"FF",X"DD",X"21",X"FE",X"17",X"06",X"18",X"DD",X"7E",X"00",X"77",X"DD",X"23",
		X"19",X"10",X"F7",X"3A",X"1E",X"81",X"3C",X"47",X"21",X"64",X"8B",X"36",X"81",X"19",X"36",X"83",
		X"19",X"10",X"F8",X"C6",X"F5",X"C0",X"01",X"40",X"00",X"09",X"36",X"81",X"19",X"36",X"82",X"19",
		X"36",X"82",X"19",X"36",X"83",X"C9",X"67",X"52",X"67",X"53",X"67",X"54",X"67",X"55",X"67",X"56",
		X"67",X"57",X"67",X"58",X"67",X"59",X"67",X"5A",X"50",X"5B",X"64",X"65",X"51",X"66",X"0F",X"80",
		X"0F",X"80",X"0F",X"80",X"0F",X"80",X"0F",X"80",X"0F",X"80",X"0F",X"80",X"0F",X"80",X"0F",X"80",
		X"0F",X"80",X"0F",X"3B",X"3B",X"80",X"DD",X"35",X"06",X"20",X"20",X"DD",X"6E",X"13",X"DD",X"66",
		X"14",X"7E",X"FE",X"80",X"20",X"06",X"23",X"5E",X"23",X"56",X"EB",X"7E",X"DD",X"77",X"05",X"23",
		X"7E",X"DD",X"77",X"06",X"23",X"DD",X"75",X"13",X"DD",X"74",X"14",X"DD",X"7E",X"05",X"DD",X"86",
		X"03",X"DD",X"77",X"03",X"ED",X"5F",X"E6",X"03",X"20",X"03",X"DD",X"34",X"04",X"DD",X"34",X"04",
		X"C9",X"21",X"BE",X"25",X"DD",X"75",X"0C",X"DD",X"74",X"0D",X"DD",X"36",X"0E",X"00",X"DD",X"36",
		X"06",X"01",X"21",X"85",X"18",X"DD",X"75",X"13",X"DD",X"74",X"14",X"DD",X"34",X"02",X"CD",X"82",
		X"1A",X"CD",X"C4",X"18",X"CD",X"16",X"18",X"DD",X"7E",X"04",X"FE",X"F0",X"D8",X"AF",X"DD",X"77",
		X"00",X"DD",X"77",X"01",X"C9",X"00",X"04",X"00",X"04",X"FF",X"30",X"FF",X"04",X"00",X"04",X"00",
		X"04",X"01",X"30",X"02",X"04",X"01",X"04",X"00",X"04",X"00",X"04",X"FF",X"04",X"FE",X"04",X"00",
		X"04",X"00",X"04",X"FF",X"04",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"04",X"00",
		X"04",X"00",X"04",X"01",X"04",X"FF",X"04",X"FF",X"04",X"01",X"04",X"00",X"04",X"00",X"04",X"00",
		X"04",X"80",X"85",X"18",X"3A",X"16",X"81",X"47",X"DD",X"7E",X"04",X"90",X"E6",X"F8",X"0F",X"0F",
		X"C6",X"C0",X"6F",X"26",X"81",X"7E",X"D6",X"1A",X"DD",X"BE",X"03",X"38",X"0C",X"2C",X"7E",X"C6",
		X"0C",X"DD",X"BE",X"03",X"D8",X"3E",X"01",X"18",X"02",X"3E",X"FF",X"DD",X"77",X"05",X"C9",X"CD",
		X"43",X"1C",X"CD",X"D4",X"1F",X"CD",X"CC",X"1D",X"CD",X"52",X"21",X"CD",X"2C",X"23",X"CD",X"14",
		X"25",X"CD",X"DB",X"24",X"CD",X"9D",X"26",X"CD",X"7D",X"27",X"CD",X"13",X"19",X"CD",X"A6",X"1D",
		X"C3",X"4A",X"1D",X"3A",X"1D",X"81",X"B7",X"F0",X"DD",X"21",X"00",X"84",X"11",X"20",X"00",X"06",
		X"04",X"D9",X"CD",X"2B",X"19",X"D9",X"DD",X"19",X"10",X"F7",X"C9",X"DD",X"7E",X"00",X"DD",X"B6",
		X"01",X"0F",X"D0",X"DD",X"7E",X"02",X"EF",X"4B",X"19",X"5C",X"19",X"29",X"1A",X"41",X"1A",X"42",
		X"1A",X"43",X"1A",X"44",X"1A",X"58",X"1A",X"70",X"1A",X"71",X"1A",X"21",X"22",X"21",X"DD",X"75",
		X"0C",X"DD",X"74",X"0D",X"DD",X"36",X"0E",X"00",X"DD",X"36",X"02",X"02",X"CD",X"82",X"1A",X"3A",
		X"22",X"81",X"D6",X"03",X"FE",X"60",X"DA",X"06",X"1A",X"DD",X"CB",X"0B",X"46",X"C2",X"06",X"1A",
		X"3A",X"16",X"81",X"47",X"DD",X"7E",X"04",X"4F",X"D6",X"06",X"90",X"E6",X"F8",X"0F",X"0F",X"C6",
		X"C0",X"6F",X"26",X"81",X"7E",X"D6",X"08",X"DD",X"BE",X"03",X"28",X"0A",X"38",X"05",X"DD",X"34",
		X"03",X"18",X"03",X"DD",X"35",X"03",X"FD",X"21",X"80",X"82",X"06",X"08",X"11",X"20",X"00",X"FD",
		X"CB",X"00",X"46",X"28",X"0B",X"FD",X"7E",X"04",X"B9",X"30",X"05",X"C6",X"10",X"B9",X"30",X"52",
		X"FD",X"19",X"10",X"EB",X"21",X"08",X"84",X"36",X"20",X"2C",X"36",X"40",X"2C",X"36",X"60",X"2E",
		X"28",X"36",X"40",X"2C",X"36",X"60",X"2C",X"36",X"00",X"2E",X"48",X"36",X"60",X"2C",X"36",X"00",
		X"2C",X"36",X"20",X"2E",X"68",X"36",X"00",X"2C",X"36",X"20",X"2C",X"36",X"40",X"DD",X"6E",X"08",
		X"CD",X"72",X"1A",X"38",X"1D",X"DD",X"6E",X"09",X"CD",X"72",X"1A",X"38",X"15",X"DD",X"6E",X"0A",
		X"CD",X"72",X"1A",X"38",X"0D",X"3A",X"84",X"83",X"91",X"D6",X"70",X"30",X"05",X"DD",X"35",X"04",
		X"18",X"04",X"DD",X"36",X"0B",X"01",X"3A",X"15",X"81",X"A7",X"20",X"03",X"DD",X"34",X"04",X"DD",
		X"7E",X"04",X"FE",X"F0",X"38",X"0B",X"AF",X"DD",X"77",X"00",X"DD",X"77",X"01",X"DD",X"77",X"0B",
		X"C9",X"DD",X"7E",X"03",X"FE",X"28",X"D0",X"18",X"ED",X"DD",X"35",X"02",X"D9",X"CB",X"40",X"D9",
		X"C8",X"DD",X"35",X"0E",X"C8",X"DD",X"34",X"02",X"3A",X"15",X"81",X"B7",X"C0",X"DD",X"34",X"04",
		X"C9",X"C9",X"C9",X"C9",X"21",X"1A",X"24",X"DD",X"75",X"0C",X"DD",X"74",X"0D",X"DD",X"36",X"0E",
		X"00",X"DD",X"36",X"0F",X"3F",X"DD",X"34",X"02",X"CD",X"82",X"1A",X"DD",X"35",X"0F",X"20",X"05",
		X"AF",X"DD",X"77",X"01",X"C9",X"3A",X"15",X"81",X"A7",X"C0",X"DD",X"34",X"04",X"C0",X"18",X"F0",
		X"C9",X"C9",X"7E",X"2C",X"B6",X"0F",X"D0",X"2C",X"2C",X"2C",X"7E",X"B9",X"D0",X"C6",X"10",X"B9",
		X"3F",X"C9",X"DD",X"7E",X"0E",X"A7",X"28",X"05",X"3D",X"DD",X"77",X"0E",X"C9",X"DD",X"6E",X"0C",
		X"DD",X"66",X"0D",X"7E",X"FE",X"FF",X"28",X"15",X"DD",X"77",X"16",X"23",X"7E",X"DD",X"77",X"12",
		X"23",X"7E",X"DD",X"77",X"0E",X"23",X"DD",X"75",X"0C",X"DD",X"74",X"0D",X"C9",X"23",X"7E",X"DD",
		X"77",X"0C",X"23",X"7E",X"DD",X"77",X"0D",X"18",X"C9",X"DD",X"E5",X"E1",X"3E",X"07",X"85",X"6F",
		X"DD",X"36",X"0A",X"00",X"DD",X"7E",X"05",X"DD",X"BE",X"03",X"28",X"04",X"38",X"1E",X"18",X"56",
		X"DD",X"7E",X"06",X"DD",X"BE",X"04",X"28",X"0E",X"38",X"06",X"36",X"00",X"2C",X"36",X"01",X"C9",
		X"36",X"00",X"2C",X"36",X"FF",X"C9",X"36",X"00",X"2C",X"36",X"00",X"C9",X"DD",X"7E",X"06",X"DD",
		X"BE",X"04",X"28",X"2C",X"38",X"15",X"36",X"FF",X"2C",X"36",X"01",X"DD",X"7E",X"03",X"DD",X"96",
		X"05",X"47",X"DD",X"7E",X"06",X"DD",X"96",X"04",X"4F",X"18",X"55",X"36",X"FF",X"2C",X"36",X"FF",
		X"DD",X"7E",X"03",X"DD",X"96",X"05",X"47",X"DD",X"7E",X"04",X"DD",X"96",X"06",X"4F",X"18",X"40",
		X"36",X"FF",X"2C",X"36",X"00",X"C9",X"DD",X"7E",X"06",X"DD",X"BE",X"04",X"28",X"2C",X"38",X"15",
		X"36",X"01",X"2C",X"36",X"01",X"DD",X"7E",X"05",X"DD",X"96",X"03",X"47",X"DD",X"7E",X"06",X"DD",
		X"96",X"04",X"4F",X"18",X"1B",X"36",X"01",X"2C",X"36",X"FF",X"DD",X"7E",X"05",X"DD",X"96",X"03",
		X"47",X"DD",X"7E",X"04",X"DD",X"96",X"06",X"4F",X"18",X"06",X"36",X"01",X"2C",X"36",X"00",X"C9",
		X"79",X"B8",X"28",X"16",X"38",X"0B",X"DD",X"36",X"09",X"00",X"CD",X"83",X"1B",X"DD",X"77",X"0B",
		X"C9",X"DD",X"36",X"09",X"01",X"78",X"41",X"4F",X"18",X"F0",X"DD",X"36",X"09",X"01",X"DD",X"36",
		X"0B",X"FF",X"C9",X"AF",X"67",X"68",X"57",X"59",X"06",X"08",X"CB",X"FF",X"07",X"29",X"A7",X"ED",
		X"52",X"38",X"03",X"10",X"F5",X"C9",X"19",X"CB",X"87",X"10",X"EF",X"C9",X"DD",X"7E",X"04",X"DD",
		X"BE",X"06",X"28",X"4A",X"DD",X"7E",X"03",X"DD",X"BE",X"05",X"28",X"58",X"DD",X"CB",X"09",X"46",
		X"28",X"1E",X"DD",X"7E",X"07",X"DD",X"86",X"03",X"DD",X"77",X"03",X"DD",X"7E",X"0B",X"DD",X"86",
		X"0A",X"DD",X"77",X"0A",X"D0",X"DD",X"7E",X"08",X"DD",X"86",X"04",X"DD",X"77",X"04",X"A7",X"C9",
		X"DD",X"7E",X"08",X"DD",X"86",X"04",X"DD",X"77",X"04",X"DD",X"7E",X"0B",X"DD",X"86",X"0A",X"DD",
		X"77",X"0A",X"D0",X"DD",X"7E",X"07",X"DD",X"86",X"03",X"DD",X"77",X"03",X"A7",X"C9",X"DD",X"7E",
		X"03",X"DD",X"BE",X"05",X"28",X"0C",X"30",X"05",X"DD",X"34",X"03",X"A7",X"C9",X"DD",X"35",X"03",
		X"A7",X"C9",X"37",X"C9",X"DD",X"7E",X"04",X"DD",X"BE",X"06",X"30",X"05",X"DD",X"34",X"04",X"A7",
		X"C9",X"DD",X"35",X"04",X"A7",X"C9",X"DD",X"6E",X"13",X"DD",X"66",X"14",X"7E",X"FE",X"80",X"20",
		X"0C",X"23",X"7E",X"DD",X"77",X"13",X"23",X"7E",X"DD",X"77",X"14",X"18",X"E9",X"DD",X"86",X"03",
		X"DD",X"77",X"03",X"23",X"7E",X"DD",X"86",X"04",X"DD",X"77",X"04",X"23",X"DD",X"75",X"13",X"DD",
		X"74",X"14",X"C9",X"DD",X"21",X"10",X"81",X"DD",X"7E",X"05",X"A7",X"20",X"12",X"DD",X"7E",X"04",
		X"DD",X"77",X"05",X"DD",X"7E",X"06",X"E6",X"0F",X"CC",X"63",X"1C",X"DD",X"34",X"06",X"C9",X"DD",
		X"35",X"05",X"C9",X"21",X"26",X"81",X"34",X"CD",X"6D",X"1C",X"C3",X"F9",X"1C",X"FD",X"2A",X"18",
		X"81",X"3E",X"01",X"32",X"10",X"81",X"32",X"30",X"82",X"DD",X"7E",X"06",X"2F",X"E6",X"F0",X"47",
		X"6F",X"26",X"22",X"29",X"29",X"E5",X"FD",X"7E",X"02",X"E6",X"F8",X"0F",X"0F",X"0F",X"5F",X"16",
		X"00",X"19",X"22",X"35",X"82",X"FD",X"7E",X"03",X"32",X"34",X"82",X"E1",X"1E",X"20",X"19",X"FD",
		X"7E",X"00",X"E6",X"F8",X"0F",X"0F",X"0F",X"5F",X"19",X"22",X"32",X"82",X"FD",X"7E",X"01",X"32",
		X"31",X"82",X"78",X"0F",X"0F",X"5F",X"21",X"C0",X"81",X"19",X"FD",X"7E",X"02",X"77",X"2C",X"36",
		X"28",X"2C",X"FD",X"7E",X"00",X"77",X"2C",X"36",X"28",X"AF",X"32",X"38",X"82",X"32",X"11",X"81",
		X"2A",X"18",X"81",X"1E",X"09",X"FD",X"7E",X"04",X"A7",X"20",X"02",X"1E",X"06",X"19",X"22",X"18",
		X"81",X"FD",X"7E",X"04",X"A7",X"FD",X"7E",X"08",X"20",X"03",X"FD",X"7E",X"05",X"32",X"1A",X"81",
		X"2A",X"35",X"82",X"2B",X"2B",X"22",X"1B",X"81",X"C9",X"FD",X"7E",X"04",X"A7",X"C8",X"68",X"26",
		X"22",X"29",X"29",X"E5",X"FD",X"7E",X"06",X"E6",X"F8",X"0F",X"0F",X"0F",X"5F",X"19",X"22",X"3D",
		X"82",X"FD",X"7E",X"07",X"32",X"3C",X"82",X"E1",X"1E",X"20",X"19",X"FD",X"7E",X"04",X"E6",X"F8",
		X"0F",X"0F",X"0F",X"5F",X"19",X"22",X"3A",X"82",X"FD",X"7E",X"05",X"32",X"39",X"82",X"78",X"0F",
		X"0F",X"5F",X"21",X"C0",X"81",X"19",X"2C",X"FD",X"7E",X"06",X"77",X"2C",X"2C",X"FD",X"7E",X"04",
		X"77",X"3E",X"01",X"32",X"11",X"81",X"32",X"38",X"82",X"C9",X"3A",X"1D",X"81",X"E6",X"10",X"20",
		X"32",X"DD",X"21",X"0C",X"85",X"11",X"03",X"00",X"06",X"03",X"CD",X"62",X"1D",X"DD",X"19",X"10",
		X"F9",X"C9",X"DD",X"CB",X"00",X"46",X"C8",X"DD",X"7E",X"02",X"C6",X"02",X"FE",X"F0",X"30",X"0E",
		X"DD",X"77",X"02",X"DD",X"7E",X"01",X"D6",X"03",X"DD",X"77",X"01",X"FE",X"1F",X"D0",X"DD",X"CB",
		X"00",X"86",X"C9",X"DD",X"21",X"0C",X"85",X"11",X"03",X"00",X"06",X"03",X"CD",X"94",X"1D",X"DD",
		X"19",X"10",X"F9",X"C9",X"DD",X"CB",X"00",X"46",X"C8",X"DD",X"7E",X"02",X"C6",X"03",X"FE",X"F0",
		X"30",X"DC",X"DD",X"77",X"02",X"C9",X"DD",X"21",X"00",X"85",X"11",X"03",X"00",X"06",X"04",X"CD",
		X"B7",X"1D",X"DD",X"19",X"10",X"F9",X"C9",X"DD",X"CB",X"00",X"46",X"C8",X"DD",X"7E",X"02",X"D6",
		X"03",X"DD",X"77",X"02",X"FE",X"1F",X"D0",X"DD",X"CB",X"00",X"86",X"C9",X"DD",X"21",X"80",X"83",
		X"DD",X"7E",X"00",X"DD",X"B6",X"01",X"0F",X"D0",X"DD",X"7E",X"02",X"EF",X"F0",X"1D",X"17",X"1E",
		X"F2",X"1E",X"30",X"1F",X"31",X"1F",X"32",X"1F",X"33",X"1F",X"51",X"1F",X"8A",X"1F",X"8B",X"1F",
		X"DD",X"36",X"03",X"58",X"DD",X"36",X"23",X"58",X"DD",X"36",X"04",X"D0",X"DD",X"36",X"24",X"E0",
		X"21",X"8C",X"1F",X"22",X"8C",X"83",X"21",X"98",X"1F",X"22",X"AC",X"83",X"DD",X"36",X"0E",X"00",
		X"DD",X"36",X"2E",X"00",X"DD",X"34",X"02",X"21",X"06",X"81",X"35",X"20",X"1B",X"3A",X"00",X"81",
		X"A7",X"28",X"07",X"3D",X"28",X"08",X"36",X"05",X"18",X"06",X"36",X"08",X"18",X"02",X"36",X"06",
		X"2D",X"35",X"20",X"04",X"DD",X"34",X"02",X"C9",X"DD",X"21",X"A0",X"83",X"CD",X"82",X"1A",X"DD",
		X"21",X"80",X"83",X"CD",X"82",X"1A",X"3A",X"06",X"80",X"0F",X"D0",X"CD",X"51",X"1E",X"C3",X"B1",
		X"1E",X"3A",X"0D",X"80",X"0F",X"38",X"43",X"3A",X"12",X"80",X"06",X"00",X"CB",X"67",X"28",X"02",
		X"CB",X"C0",X"CB",X"77",X"28",X"02",X"CB",X"C8",X"78",X"0F",X"30",X"16",X"3A",X"5F",X"82",X"E6",
		X"3F",X"CC",X"6C",X"37",X"DD",X"7E",X"03",X"3D",X"FE",X"38",X"D8",X"DD",X"77",X"03",X"DD",X"35",
		X"23",X"C9",X"0F",X"D0",X"3A",X"5F",X"82",X"E6",X"3F",X"CC",X"6C",X"37",X"DD",X"7E",X"03",X"3C",
		X"FE",X"D8",X"D0",X"DD",X"77",X"03",X"DD",X"34",X"23",X"C9",X"3A",X"12",X"80",X"06",X"00",X"CB",
		X"47",X"28",X"02",X"CB",X"C8",X"3A",X"10",X"80",X"CB",X"47",X"28",X"02",X"CB",X"C0",X"78",X"18",
		X"B8",X"3A",X"0D",X"80",X"0F",X"38",X"36",X"3A",X"10",X"80",X"07",X"07",X"07",X"30",X"16",X"3A",
		X"5F",X"82",X"E6",X"3F",X"CC",X"6C",X"37",X"DD",X"7E",X"04",X"3C",X"FE",X"D0",X"D0",X"DD",X"77",
		X"04",X"DD",X"34",X"24",X"C9",X"07",X"D0",X"3A",X"5F",X"82",X"E6",X"3F",X"CC",X"6C",X"37",X"DD",
		X"7E",X"04",X"3D",X"FE",X"80",X"D8",X"DD",X"77",X"04",X"DD",X"35",X"24",X"C9",X"3A",X"11",X"80",
		X"18",X"C8",X"DD",X"21",X"A0",X"83",X"CD",X"82",X"1A",X"DD",X"21",X"80",X"83",X"CD",X"82",X"1A",
		X"3A",X"05",X"81",X"B7",X"20",X"25",X"DD",X"34",X"03",X"DD",X"34",X"23",X"DD",X"7E",X"03",X"FE",
		X"F0",X"D8",X"DD",X"36",X"00",X"00",X"DD",X"36",X"01",X"01",X"DD",X"36",X"02",X"06",X"DD",X"36",
		X"20",X"00",X"DD",X"36",X"21",X"01",X"DD",X"36",X"22",X"06",X"C9",X"DD",X"36",X"02",X"01",X"C9",
		X"C9",X"C9",X"C9",X"CD",X"99",X"37",X"21",X"A4",X"1F",X"22",X"8C",X"83",X"DD",X"36",X"0E",X"00",
		X"DD",X"36",X"0F",X"6F",X"21",X"BC",X"1F",X"22",X"AC",X"83",X"DD",X"36",X"2E",X"00",X"DD",X"34",
		X"02",X"3A",X"5F",X"82",X"E6",X"03",X"CC",X"80",X"1F",X"DD",X"21",X"A0",X"83",X"CD",X"82",X"1A",
		X"DD",X"21",X"80",X"83",X"CD",X"82",X"1A",X"3A",X"15",X"81",X"A7",X"20",X"06",X"DD",X"34",X"04",
		X"DD",X"34",X"24",X"DD",X"35",X"0F",X"C0",X"DD",X"36",X"01",X"00",X"DD",X"36",X"21",X"00",X"C9",
		X"3A",X"17",X"81",X"3C",X"E6",X"07",X"32",X"17",X"81",X"C9",X"C9",X"C9",X"00",X"2A",X"01",X"00",
		X"2C",X"01",X"00",X"2E",X"01",X"FF",X"8C",X"1F",X"00",X"29",X"01",X"00",X"2B",X"01",X"00",X"2D",
		X"01",X"FF",X"98",X"1F",X"02",X"3C",X"07",X"02",X"3D",X"07",X"02",X"3C",X"07",X"02",X"3D",X"07",
		X"02",X"3C",X"07",X"02",X"3D",X"07",X"02",X"3E",X"07",X"FF",X"A4",X"1F",X"02",X"BC",X"07",X"02",
		X"BD",X"07",X"02",X"BC",X"07",X"02",X"BD",X"07",X"02",X"BC",X"07",X"02",X"BD",X"07",X"02",X"BE",
		X"07",X"FF",X"BC",X"1F",X"DD",X"21",X"80",X"82",X"11",X"20",X"00",X"06",X"08",X"D9",X"CD",X"E7",
		X"1F",X"D9",X"DD",X"19",X"10",X"F7",X"C9",X"DD",X"7E",X"00",X"DD",X"B6",X"01",X"0F",X"D0",X"DD",
		X"7E",X"02",X"EF",X"07",X"20",X"68",X"20",X"80",X"20",X"81",X"20",X"9B",X"20",X"9C",X"20",X"9D",
		X"20",X"EB",X"20",X"08",X"21",X"09",X"21",X"2A",X"1B",X"81",X"DD",X"75",X"18",X"DD",X"74",X"19",
		X"3A",X"16",X"81",X"E6",X"0F",X"C6",X"F8",X"DD",X"77",X"04",X"7D",X"E6",X"1F",X"07",X"07",X"07",
		X"C6",X"08",X"DD",X"77",X"03",X"DD",X"7E",X"17",X"A7",X"28",X"1D",X"3D",X"28",X"10",X"3D",X"28",
		X"12",X"3D",X"28",X"05",X"21",X"22",X"21",X"18",X"22",X"21",X"28",X"21",X"18",X"1D",X"21",X"0A",
		X"21",X"18",X"18",X"21",X"2E",X"21",X"18",X"13",X"21",X"0A",X"21",X"3A",X"1D",X"81",X"E6",X"06",
		X"20",X"02",X"3E",X"04",X"47",X"07",X"80",X"4F",X"06",X"00",X"09",X"DD",X"75",X"0C",X"DD",X"74",
		X"0D",X"DD",X"36",X"0E",X"00",X"DD",X"34",X"02",X"CD",X"82",X"1A",X"3A",X"15",X"81",X"A7",X"C0",
		X"DD",X"34",X"04",X"DD",X"7E",X"04",X"C6",X"0D",X"FE",X"08",X"D0",X"DD",X"36",X"02",X"03",X"C9",
		X"C9",X"DD",X"6E",X"18",X"DD",X"66",X"19",X"3E",X"10",X"77",X"23",X"77",X"11",X"1F",X"00",X"19",
		X"77",X"23",X"77",X"AF",X"DD",X"77",X"00",X"DD",X"77",X"01",X"C9",X"C9",X"C9",X"DD",X"7E",X"17",
		X"3D",X"28",X"05",X"3D",X"28",X"09",X"18",X"2E",X"21",X"43",X"21",X"3E",X"3F",X"18",X"2C",X"DD",
		X"36",X"0E",X"50",X"DD",X"36",X"0F",X"3F",X"DD",X"34",X"02",X"DD",X"46",X"1A",X"3E",X"4F",X"05",
		X"28",X"05",X"05",X"28",X"07",X"18",X"0A",X"DD",X"36",X"12",X"46",X"C9",X"DD",X"36",X"12",X"47",
		X"C9",X"DD",X"36",X"12",X"45",X"C9",X"21",X"34",X"21",X"3E",X"3F",X"DD",X"75",X"0C",X"DD",X"74",
		X"0D",X"DD",X"36",X"0E",X"00",X"DD",X"77",X"0F",X"DD",X"34",X"02",X"CD",X"82",X"1A",X"DD",X"35",
		X"0F",X"28",X"10",X"3A",X"15",X"81",X"A7",X"C0",X"DD",X"34",X"04",X"DD",X"7E",X"04",X"C6",X"14",
		X"FE",X"08",X"D0",X"DD",X"36",X"02",X"03",X"C9",X"C9",X"C9",X"02",X"10",X"10",X"FF",X"0A",X"21",
		X"00",X"1B",X"10",X"FF",X"10",X"21",X"02",X"1C",X"10",X"FF",X"16",X"21",X"00",X"1F",X"10",X"FF",
		X"1C",X"21",X"02",X"33",X"10",X"FF",X"22",X"21",X"00",X"2F",X"FF",X"FF",X"28",X"21",X"00",X"28",
		X"FF",X"FF",X"2E",X"21",X"07",X"38",X"10",X"07",X"39",X"10",X"07",X"3A",X"10",X"07",X"3B",X"10",
		X"FF",X"34",X"21",X"07",X"38",X"10",X"07",X"39",X"10",X"07",X"3A",X"10",X"07",X"3B",X"10",X"FF",
		X"43",X"21",X"3A",X"12",X"81",X"FE",X"41",X"28",X"13",X"DD",X"21",X"C0",X"83",X"11",X"20",X"00",
		X"06",X"02",X"D9",X"CD",X"BC",X"21",X"D9",X"DD",X"19",X"10",X"F7",X"C9",X"DD",X"21",X"C0",X"83",
		X"DD",X"7E",X"02",X"EF",X"DC",X"21",X"99",X"21",X"19",X"22",X"1A",X"22",X"1B",X"22",X"1C",X"22",
		X"88",X"21",X"31",X"22",X"47",X"22",X"48",X"22",X"3E",X"0A",X"32",X"12",X"81",X"21",X"BA",X"22",
		X"DD",X"75",X"13",X"DD",X"74",X"14",X"C3",X"1D",X"22",X"CD",X"82",X"1A",X"21",X"84",X"83",X"11",
		X"C4",X"83",X"7E",X"C6",X"03",X"12",X"2B",X"1B",X"7E",X"C6",X"06",X"12",X"2B",X"3E",X"06",X"BE",
		X"30",X"06",X"1B",X"EB",X"BE",X"38",X"01",X"77",X"DD",X"21",X"E0",X"83",X"DD",X"7E",X"00",X"DD",
		X"B6",X"01",X"0F",X"D0",X"DD",X"7E",X"02",X"EF",X"DC",X"21",X"05",X"22",X"19",X"22",X"1A",X"22",
		X"1B",X"22",X"1C",X"22",X"1D",X"22",X"31",X"22",X"47",X"22",X"48",X"22",X"3A",X"83",X"83",X"C6",
		X"04",X"DD",X"77",X"03",X"3A",X"84",X"83",X"C6",X"08",X"DD",X"77",X"04",X"21",X"49",X"22",X"DD",
		X"75",X"0C",X"DD",X"74",X"0D",X"DD",X"36",X"0E",X"00",X"21",X"64",X"22",X"DD",X"75",X"13",X"DD",
		X"74",X"14",X"DD",X"34",X"02",X"CD",X"82",X"1A",X"CD",X"16",X"1C",X"DD",X"7E",X"03",X"FE",X"F0",
		X"D8",X"AF",X"DD",X"77",X"00",X"DD",X"77",X"01",X"C9",X"C9",X"C9",X"C9",X"C9",X"21",X"55",X"22",
		X"DD",X"75",X"0C",X"DD",X"74",X"0D",X"DD",X"36",X"0E",X"00",X"DD",X"36",X"0F",X"23",X"DD",X"34",
		X"02",X"CD",X"82",X"1A",X"DD",X"35",X"0F",X"20",X"05",X"AF",X"DD",X"77",X"01",X"C9",X"3A",X"15",
		X"81",X"A7",X"C0",X"DD",X"34",X"04",X"C9",X"C9",X"C9",X"00",X"21",X"10",X"00",X"22",X"16",X"00",
		X"23",X"FE",X"FF",X"49",X"22",X"07",X"38",X"09",X"07",X"39",X"09",X"07",X"3A",X"09",X"07",X"3B",
		X"09",X"FF",X"55",X"22",X"00",X"00",X"01",X"00",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"01",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"01",X"FF",
		X"00",X"FF",X"00",X"FF",X"01",X"FF",X"00",X"FF",X"01",X"FF",X"01",X"FF",X"00",X"FF",X"01",X"FF",
		X"01",X"FF",X"01",X"FF",X"01",X"00",X"01",X"00",X"01",X"FF",X"01",X"FF",X"01",X"00",X"01",X"FF",
		X"01",X"00",X"01",X"FF",X"01",X"00",X"01",X"00",X"01",X"FF",X"01",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"80",X"BA",X"22",X"DD",X"21",X"00",X"84",X"11",X"20",X"00",X"06",X"04",X"D9",X"CD",
		X"D8",X"22",X"D9",X"DD",X"19",X"10",X"F7",X"C9",X"DD",X"7E",X"00",X"DD",X"B6",X"01",X"0F",X"D0",
		X"DD",X"7E",X"02",X"EF",X"F8",X"22",X"12",X"23",X"C1",X"23",X"D9",X"23",X"DA",X"23",X"DB",X"23",
		X"DC",X"23",X"F7",X"23",X"0F",X"24",X"10",X"24",X"21",X"26",X"23",X"DD",X"75",X"0C",X"DD",X"74",
		X"0D",X"DD",X"36",X"0E",X"00",X"21",X"2E",X"24",X"DD",X"75",X"13",X"DD",X"74",X"14",X"DD",X"36",
		X"02",X"02",X"CD",X"82",X"1A",X"CD",X"16",X"1C",X"3A",X"15",X"81",X"A7",X"C0",X"DD",X"34",X"04",
		X"C0",X"DD",X"36",X"00",X"00",X"C9",X"07",X"1F",X"10",X"FF",X"26",X"23",X"3A",X"1D",X"81",X"E6",
		X"06",X"C8",X"0F",X"3D",X"EF",X"33",X"24",X"3B",X"23",X"C5",X"22",X"DD",X"21",X"00",X"84",X"11",
		X"20",X"00",X"06",X"04",X"D9",X"CD",X"4E",X"23",X"D9",X"DD",X"19",X"10",X"F7",X"C9",X"DD",X"7E",
		X"00",X"DD",X"B6",X"01",X"0F",X"D0",X"DD",X"7E",X"02",X"EF",X"6E",X"23",X"8E",X"23",X"C1",X"23",
		X"D9",X"23",X"DA",X"23",X"DB",X"23",X"DC",X"23",X"F7",X"23",X"0F",X"24",X"10",X"24",X"DD",X"34",
		X"03",X"DD",X"34",X"03",X"21",X"11",X"24",X"DD",X"75",X"0C",X"DD",X"74",X"0D",X"DD",X"36",X"0E",
		X"00",X"21",X"29",X"24",X"DD",X"75",X"13",X"DD",X"74",X"14",X"DD",X"36",X"02",X"02",X"CD",X"82",
		X"1A",X"CD",X"16",X"1C",X"D9",X"CB",X"40",X"D9",X"28",X"07",X"DD",X"35",X"03",X"DD",X"36",X"16",
		X"06",X"3A",X"15",X"81",X"A7",X"20",X"03",X"DD",X"34",X"04",X"DD",X"7E",X"04",X"FE",X"F0",X"38",
		X"08",X"AF",X"DD",X"77",X"00",X"DD",X"77",X"01",X"C9",X"DD",X"7E",X"03",X"FE",X"28",X"D0",X"18",
		X"F0",X"DD",X"35",X"02",X"D9",X"CB",X"40",X"D9",X"C8",X"DD",X"35",X"0E",X"C8",X"DD",X"34",X"02",
		X"3A",X"15",X"81",X"B7",X"C0",X"DD",X"34",X"04",X"C9",X"C9",X"C9",X"C9",X"DD",X"7E",X"04",X"FE",
		X"0C",X"38",X"1C",X"21",X"1A",X"24",X"DD",X"75",X"0C",X"DD",X"74",X"0D",X"DD",X"36",X"0E",X"00",
		X"DD",X"36",X"0F",X"3F",X"DD",X"34",X"02",X"CD",X"82",X"1A",X"DD",X"35",X"0F",X"20",X"05",X"AF",
		X"DD",X"77",X"01",X"C9",X"3A",X"15",X"81",X"A7",X"C0",X"DD",X"34",X"04",X"C0",X"18",X"F0",X"C9",
		X"C9",X"04",X"1D",X"10",X"04",X"1E",X"10",X"FF",X"11",X"24",X"07",X"38",X"05",X"07",X"39",X"05",
		X"07",X"3A",X"05",X"07",X"3B",X"05",X"FF",X"1A",X"24",X"FF",X"00",X"80",X"29",X"24",X"01",X"00",
		X"80",X"2E",X"24",X"DD",X"21",X"00",X"84",X"11",X"20",X"00",X"06",X"04",X"D9",X"CD",X"46",X"24",
		X"D9",X"DD",X"19",X"10",X"F7",X"C9",X"DD",X"7E",X"00",X"DD",X"B6",X"01",X"0F",X"D0",X"DD",X"7E",
		X"02",X"EF",X"66",X"24",X"7D",X"24",X"7D",X"25",X"7E",X"25",X"7F",X"25",X"80",X"25",X"81",X"25",
		X"95",X"25",X"B0",X"25",X"B1",X"25",X"CD",X"C1",X"37",X"DD",X"7E",X"03",X"DD",X"77",X"05",X"DD",
		X"36",X"07",X"FD",X"DD",X"77",X"08",X"DD",X"34",X"02",X"DD",X"36",X"16",X"03",X"11",X"08",X"00",
		X"DD",X"66",X"07",X"DD",X"6E",X"08",X"19",X"DC",X"C6",X"37",X"DD",X"74",X"07",X"DD",X"75",X"08",
		X"E5",X"DD",X"56",X"03",X"DD",X"5E",X"06",X"19",X"3E",X"24",X"BC",X"30",X"01",X"7C",X"DD",X"77",
		X"03",X"DD",X"75",X"06",X"DD",X"7E",X"04",X"C6",X"02",X"D9",X"CB",X"40",X"D9",X"28",X"02",X"D6",
		X"03",X"DD",X"77",X"04",X"DC",X"14",X"33",X"C1",X"CB",X"11",X"CB",X"10",X"78",X"0E",X"00",X"30",
		X"03",X"0E",X"40",X"2F",X"CB",X"3F",X"FE",X"03",X"38",X"02",X"3E",X"02",X"C6",X"A5",X"81",X"D9",
		X"CB",X"40",X"D9",X"28",X"02",X"EE",X"80",X"DD",X"77",X"12",X"C9",X"3A",X"1D",X"81",X"E6",X"10",
		X"C8",X"DD",X"21",X"00",X"84",X"11",X"20",X"00",X"06",X"04",X"D9",X"CD",X"F4",X"24",X"D9",X"DD",
		X"19",X"10",X"F7",X"C9",X"DD",X"7E",X"00",X"DD",X"B6",X"01",X"0F",X"D0",X"DD",X"7E",X"02",X"EF",
		X"51",X"18",X"6E",X"18",X"7D",X"25",X"7E",X"25",X"7F",X"25",X"80",X"25",X"81",X"25",X"95",X"25",
		X"B0",X"25",X"B1",X"25",X"3A",X"1D",X"81",X"E6",X"08",X"C8",X"DD",X"21",X"00",X"84",X"11",X"20",
		X"00",X"06",X"04",X"D9",X"CD",X"2D",X"25",X"D9",X"DD",X"19",X"10",X"F7",X"C9",X"DD",X"7E",X"00",
		X"DD",X"B6",X"01",X"0F",X"D0",X"DD",X"7E",X"02",X"EF",X"4D",X"25",X"66",X"25",X"7D",X"25",X"7E",
		X"25",X"7F",X"25",X"80",X"25",X"81",X"25",X"95",X"25",X"B0",X"25",X"B1",X"25",X"21",X"B2",X"25",
		X"DD",X"75",X"0C",X"DD",X"74",X"0D",X"DD",X"36",X"0E",X"00",X"21",X"D6",X"25",X"DD",X"75",X"13",
		X"DD",X"74",X"14",X"DD",X"34",X"02",X"CD",X"82",X"1A",X"CD",X"6D",X"26",X"CD",X"16",X"1C",X"DD",
		X"7E",X"04",X"FE",X"F0",X"D8",X"AF",X"DD",X"77",X"00",X"DD",X"77",X"01",X"C9",X"C9",X"C9",X"C9",
		X"C9",X"21",X"C7",X"25",X"DD",X"75",X"0C",X"DD",X"74",X"0D",X"DD",X"36",X"0E",X"00",X"DD",X"36",
		X"0F",X"2B",X"DD",X"34",X"02",X"CD",X"82",X"1A",X"DD",X"35",X"0F",X"20",X"05",X"AF",X"DD",X"77",
		X"01",X"C9",X"3A",X"15",X"81",X"A7",X"C0",X"DD",X"34",X"04",X"C0",X"DD",X"36",X"01",X"00",X"C9",
		X"C9",X"C9",X"02",X"D2",X"01",X"02",X"D3",X"01",X"02",X"DA",X"01",X"FF",X"B2",X"25",X"05",X"3F",
		X"10",X"05",X"3F",X"10",X"FF",X"BE",X"25",X"05",X"38",X"0B",X"05",X"39",X"0B",X"05",X"3A",X"0B",
		X"05",X"3B",X"0B",X"FF",X"C7",X"25",X"FF",X"00",X"FE",X"00",X"FE",X"00",X"FE",X"00",X"FE",X"00",
		X"FE",X"00",X"FE",X"00",X"FE",X"00",X"FE",X"00",X"FE",X"02",X"FE",X"00",X"FE",X"02",X"FE",X"00",
		X"FE",X"02",X"FE",X"02",X"FE",X"02",X"FE",X"02",X"00",X"02",X"00",X"02",X"01",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"00",X"02",X"02",X"02",X"00",X"02",X"02",
		X"02",X"00",X"02",X"02",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"02",
		X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"02",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",
		X"02",X"02",X"02",X"00",X"02",X"02",X"02",X"00",X"02",X"00",X"02",X"02",X"02",X"02",X"02",X"02",
		X"00",X"02",X"00",X"02",X"00",X"02",X"FF",X"02",X"FE",X"02",X"FE",X"02",X"FE",X"02",X"FE",X"00",
		X"FE",X"02",X"FE",X"00",X"FE",X"02",X"FE",X"00",X"FE",X"02",X"FE",X"00",X"FE",X"02",X"FE",X"00",
		X"FE",X"00",X"FE",X"00",X"FE",X"00",X"FE",X"00",X"FE",X"00",X"80",X"D6",X"25",X"3A",X"16",X"81",
		X"47",X"DD",X"7E",X"04",X"90",X"E6",X"F8",X"0F",X"0F",X"C6",X"C0",X"6F",X"26",X"81",X"7E",X"D6",
		X"1A",X"DD",X"BE",X"03",X"38",X"0D",X"2C",X"7E",X"C6",X"0C",X"DD",X"BE",X"03",X"D8",X"21",X"FC",
		X"25",X"18",X"03",X"21",X"46",X"26",X"DD",X"75",X"13",X"DD",X"74",X"14",X"C9",X"3A",X"1D",X"81",
		X"E6",X"20",X"C8",X"DD",X"21",X"00",X"84",X"11",X"20",X"00",X"06",X"04",X"D9",X"CD",X"B6",X"26",
		X"D9",X"DD",X"19",X"10",X"F7",X"C9",X"DD",X"7E",X"00",X"DD",X"B6",X"01",X"0F",X"D0",X"DD",X"7E",
		X"02",X"EF",X"D6",X"26",X"FC",X"26",X"7D",X"25",X"7E",X"25",X"7F",X"25",X"80",X"25",X"81",X"25",
		X"95",X"25",X"B0",X"25",X"B1",X"25",X"11",X"49",X"27",X"21",X"73",X"27",X"D9",X"78",X"FE",X"01",
		X"D9",X"20",X"06",X"11",X"5E",X"27",X"21",X"78",X"27",X"DD",X"73",X"0C",X"DD",X"72",X"0D",X"DD",
		X"36",X"0E",X"00",X"DD",X"75",X"13",X"DD",X"74",X"14",X"DD",X"34",X"02",X"CD",X"82",X"1A",X"D9",
		X"78",X"FE",X"01",X"D9",X"28",X"1E",X"CD",X"16",X"1C",X"3E",X"AF",X"DD",X"BE",X"03",X"30",X"03",
		X"DD",X"77",X"03",X"DD",X"7E",X"04",X"FE",X"F0",X"D8",X"AF",X"DD",X"77",X"00",X"DD",X"77",X"01",
		X"DD",X"77",X"05",X"C9",X"DD",X"7E",X"05",X"C6",X"03",X"DD",X"77",X"16",X"21",X"09",X"27",X"E5",
		X"ED",X"5F",X"E6",X"03",X"C8",X"3A",X"83",X"83",X"DD",X"34",X"04",X"DD",X"BE",X"03",X"C8",X"38",
		X"04",X"DD",X"34",X"03",X"C9",X"DD",X"35",X"03",X"C9",X"02",X"35",X"05",X"02",X"36",X"05",X"02",
		X"37",X"05",X"02",X"30",X"05",X"02",X"37",X"05",X"02",X"36",X"05",X"FF",X"49",X"27",X"04",X"35",
		X"05",X"00",X"36",X"05",X"02",X"37",X"05",X"00",X"30",X"05",X"02",X"37",X"05",X"00",X"36",X"05",
		X"FF",X"5E",X"27",X"00",X"04",X"80",X"73",X"27",X"01",X"04",X"80",X"78",X"27",X"3A",X"1D",X"81",
		X"E6",X"40",X"C8",X"DD",X"21",X"00",X"84",X"11",X"20",X"00",X"06",X"04",X"D9",X"CD",X"96",X"27",
		X"D9",X"DD",X"19",X"10",X"F7",X"C9",X"DD",X"7E",X"00",X"DD",X"B6",X"01",X"0F",X"D0",X"DD",X"7E",
		X"02",X"EF",X"B6",X"27",X"C2",X"27",X"21",X"28",X"5D",X"28",X"7E",X"28",X"80",X"25",X"81",X"25",
		X"95",X"25",X"B0",X"25",X"B1",X"25",X"11",X"B2",X"25",X"DD",X"73",X"0C",X"DD",X"72",X"0D",X"DD",
		X"34",X"02",X"CD",X"82",X"1A",X"3A",X"5F",X"82",X"07",X"38",X"06",X"DD",X"34",X"03",X"C3",X"D4",
		X"27",X"DD",X"35",X"03",X"DD",X"34",X"04",X"ED",X"5B",X"83",X"83",X"ED",X"5F",X"E6",X"1F",X"DD",
		X"86",X"04",X"92",X"2F",X"47",X"DD",X"7E",X"03",X"FE",X"30",X"30",X"04",X"DD",X"36",X"03",X"30",
		X"FE",X"B0",X"38",X"04",X"DD",X"36",X"03",X"B0",X"93",X"30",X"01",X"2F",X"07",X"B8",X"D8",X"21",
		X"02",X"84",X"01",X"01",X"04",X"11",X"20",X"00",X"79",X"BE",X"28",X"07",X"19",X"10",X"FA",X"DD",
		X"34",X"02",X"C9",X"2C",X"2C",X"7E",X"3D",X"2D",X"2D",X"DD",X"BE",X"04",X"D0",X"79",X"C3",X"0C",
		X"28",X"CD",X"82",X"1A",X"DD",X"34",X"04",X"DD",X"34",X"04",X"DD",X"34",X"04",X"DD",X"7E",X"04",
		X"FE",X"F0",X"30",X"21",X"3A",X"83",X"83",X"DD",X"BE",X"03",X"CA",X"70",X"30",X"30",X"0B",X"DD",
		X"35",X"03",X"DD",X"36",X"02",X"03",X"CD",X"D5",X"37",X"C9",X"DD",X"34",X"03",X"DD",X"36",X"02",
		X"04",X"CD",X"D5",X"37",X"C9",X"AF",X"DD",X"77",X"00",X"DD",X"77",X"01",X"C9",X"CD",X"82",X"1A",
		X"DD",X"34",X"04",X"DD",X"34",X"04",X"DD",X"34",X"04",X"DD",X"7E",X"04",X"FE",X"F0",X"30",X"E5",
		X"DD",X"35",X"03",X"DD",X"7E",X"03",X"FE",X"30",X"D0",X"DD",X"36",X"02",X"02",X"C9",X"CD",X"82",
		X"1A",X"DD",X"34",X"04",X"DD",X"34",X"04",X"DD",X"34",X"04",X"DD",X"7E",X"04",X"FE",X"F0",X"30",
		X"C4",X"DD",X"34",X"03",X"DD",X"7E",X"03",X"FE",X"B0",X"D8",X"DD",X"36",X"02",X"02",X"C3",X"70",
		X"30",X"CD",X"B0",X"28",X"CD",X"C5",X"28",X"CD",X"F6",X"28",X"CD",X"00",X"29",X"C3",X"4F",X"29",
		X"21",X"2A",X"80",X"06",X"19",X"3A",X"16",X"81",X"ED",X"44",X"4F",X"3A",X"17",X"81",X"71",X"2C",
		X"77",X"2C",X"10",X"FA",X"C9",X"21",X"60",X"82",X"DD",X"21",X"80",X"82",X"11",X"20",X"00",X"06",
		X"08",X"CD",X"D9",X"28",X"DD",X"19",X"10",X"F9",X"C9",X"DD",X"7E",X"00",X"DD",X"B6",X"01",X"0F",
		X"36",X"00",X"D0",X"36",X"01",X"2C",X"DD",X"7E",X"12",X"77",X"2C",X"DD",X"7E",X"18",X"77",X"2C",
		X"DD",X"7E",X"19",X"77",X"2C",X"C9",X"DD",X"21",X"80",X"83",X"FD",X"21",X"60",X"80",X"18",X"12",
		X"DD",X"21",X"00",X"84",X"FD",X"21",X"70",X"80",X"18",X"08",X"DD",X"21",X"80",X"84",X"FD",X"21",
		X"70",X"80",X"01",X"08",X"04",X"DD",X"7E",X"00",X"DD",X"B6",X"01",X"0F",X"30",X"27",X"DD",X"7E",
		X"16",X"FD",X"77",X"02",X"DD",X"7E",X"03",X"91",X"FD",X"77",X"03",X"DD",X"7E",X"04",X"2F",X"91",
		X"FD",X"77",X"00",X"DD",X"7E",X"12",X"FD",X"77",X"01",X"11",X"20",X"00",X"DD",X"19",X"1E",X"04",
		X"FD",X"19",X"10",X"D1",X"C9",X"FD",X"36",X"00",X"F8",X"FD",X"36",X"03",X"F8",X"18",X"EA",X"DD",
		X"21",X"80",X"80",X"FD",X"21",X"00",X"85",X"06",X"07",X"CD",X"67",X"29",X"11",X"04",X"00",X"DD",
		X"19",X"1D",X"FD",X"19",X"10",X"F3",X"C9",X"FD",X"CB",X"00",X"46",X"28",X"23",X"FD",X"7E",X"02",
		X"2F",X"DD",X"77",X"01",X"FD",X"7E",X"01",X"C6",X"05",X"DD",X"77",X"03",X"3A",X"0F",X"80",X"0F",
		X"30",X"06",X"3A",X"0D",X"80",X"0F",X"38",X"11",X"DD",X"7E",X"03",X"2F",X"DD",X"77",X"03",X"C9",
		X"DD",X"36",X"01",X"00",X"DD",X"36",X"03",X"00",X"C9",X"DD",X"7E",X"03",X"D6",X"0D",X"DD",X"77",
		X"03",X"C9",X"CD",X"D9",X"29",X"CD",X"3D",X"2A",X"CD",X"EA",X"2A",X"CD",X"06",X"2B",X"CD",X"2B",
		X"2C",X"CD",X"CD",X"2A",X"CD",X"65",X"2B",X"CD",X"D5",X"2C",X"CD",X"A9",X"2D",X"CD",X"0D",X"2E",
		X"CD",X"47",X"2E",X"CD",X"B6",X"2E",X"CD",X"16",X"2F",X"CD",X"A7",X"2F",X"CD",X"12",X"30",X"CD",
		X"57",X"30",X"CD",X"C9",X"2B",X"CD",X"64",X"2C",X"C9",X"3A",X"80",X"83",X"0F",X"D0",X"3A",X"1D",
		X"81",X"E6",X"D8",X"C8",X"DD",X"21",X"00",X"84",X"11",X"20",X"00",X"06",X"04",X"CD",X"F5",X"29",
		X"DD",X"19",X"10",X"F9",X"C9",X"DD",X"CB",X"00",X"46",X"C8",X"21",X"83",X"83",X"7E",X"DD",X"96",
		X"03",X"C6",X"0A",X"FE",X"0F",X"D0",X"2C",X"7E",X"C6",X"04",X"DD",X"96",X"04",X"C6",X"0D",X"FE",
		X"19",X"D0",X"DD",X"CB",X"00",X"86",X"DD",X"CB",X"01",X"C6",X"DD",X"36",X"02",X"06",X"2D",X"2D",
		X"36",X"06",X"2D",X"36",X"01",X"2D",X"36",X"00",X"21",X"A0",X"83",X"36",X"00",X"2C",X"36",X"01",
		X"DD",X"36",X"17",X"00",X"3E",X"FF",X"32",X"15",X"81",X"CD",X"FD",X"36",X"C9",X"3A",X"80",X"83",
		X"0F",X"D0",X"3A",X"1D",X"81",X"E6",X"20",X"C8",X"DD",X"21",X"00",X"84",X"11",X"20",X"00",X"06",
		X"04",X"CD",X"F5",X"29",X"DD",X"19",X"10",X"F9",X"C9",X"DD",X"21",X"80",X"82",X"11",X"20",X"00",
		X"06",X"08",X"DD",X"7E",X"17",X"FE",X"03",X"28",X"08",X"CD",X"F5",X"29",X"DD",X"19",X"10",X"F2",
		X"C9",X"21",X"6C",X"2A",X"E5",X"DD",X"CB",X"00",X"46",X"C8",X"21",X"83",X"83",X"7E",X"DD",X"96",
		X"03",X"C6",X"0B",X"FE",X"06",X"D0",X"2C",X"7E",X"C6",X"04",X"DD",X"96",X"04",X"C6",X"0D",X"FE",
		X"19",X"D0",X"DD",X"36",X"02",X"03",X"11",X"C4",X"83",X"01",X"05",X"00",X"ED",X"B8",X"21",X"80",
		X"85",X"36",X"96",X"2C",X"36",X"00",X"21",X"0A",X"80",X"36",X"08",X"2D",X"36",X"64",X"3E",X"41",
		X"32",X"12",X"81",X"3E",X"82",X"32",X"22",X"81",X"3E",X"01",X"32",X"CE",X"83",X"2A",X"20",X"81",
		X"23",X"23",X"22",X"20",X"81",X"21",X"28",X"21",X"22",X"CC",X"83",X"E1",X"C9",X"3A",X"80",X"83",
		X"0F",X"D0",X"3A",X"1E",X"81",X"FE",X"0A",X"28",X"80",X"DD",X"21",X"80",X"82",X"11",X"20",X"00",
		X"06",X"08",X"CD",X"F5",X"29",X"DD",X"19",X"10",X"F9",X"C9",X"3A",X"80",X"83",X"0F",X"D0",X"3A",
		X"1D",X"81",X"E6",X"06",X"C8",X"DD",X"21",X"00",X"84",X"11",X"20",X"00",X"06",X"04",X"CD",X"F5",
		X"29",X"DD",X"19",X"10",X"F9",X"C9",X"3A",X"80",X"83",X"0F",X"D0",X"3A",X"16",X"81",X"47",X"3A",
		X"84",X"83",X"D6",X"04",X"90",X"E6",X"F8",X"0F",X"0F",X"C6",X"C0",X"6F",X"26",X"81",X"01",X"04",
		X"04",X"3A",X"83",X"83",X"C6",X"03",X"5F",X"D6",X"06",X"57",X"7E",X"81",X"BB",X"38",X"1A",X"2C",
		X"7E",X"91",X"BA",X"30",X"14",X"0E",X"00",X"78",X"FE",X"02",X"20",X"02",X"0E",X"04",X"2C",X"28",
		X"03",X"10",X"E7",X"C9",X"2E",X"C0",X"10",X"E2",X"C9",X"21",X"80",X"83",X"36",X"00",X"2C",X"36",
		X"01",X"2C",X"36",X"06",X"21",X"A0",X"83",X"36",X"00",X"2C",X"36",X"01",X"3E",X"FF",X"32",X"15",
		X"81",X"CD",X"FD",X"36",X"C9",X"3A",X"1D",X"81",X"E6",X"58",X"C8",X"FD",X"21",X"00",X"85",X"06",
		X"04",X"11",X"20",X"00",X"CD",X"80",X"2B",X"FD",X"23",X"FD",X"23",X"FD",X"23",X"10",X"F5",X"C9",
		X"FD",X"CB",X"00",X"46",X"C8",X"DD",X"21",X"00",X"84",X"0E",X"04",X"D9",X"CD",X"96",X"2B",X"D9",
		X"DD",X"19",X"0D",X"20",X"F6",X"C9",X"DD",X"CB",X"00",X"46",X"C8",X"FD",X"7E",X"01",X"DD",X"96",
		X"03",X"C6",X"04",X"FE",X"09",X"D0",X"FD",X"7E",X"02",X"DD",X"96",X"04",X"C6",X"04",X"FE",X"09",
		X"D0",X"DD",X"36",X"00",X"00",X"DD",X"36",X"01",X"01",X"DD",X"36",X"02",X"06",X"FD",X"36",X"00",
		X"00",X"11",X"08",X"03",X"FF",X"CD",X"F5",X"36",X"C9",X"3A",X"1D",X"81",X"E6",X"80",X"C8",X"FD",
		X"21",X"00",X"85",X"06",X"04",X"11",X"20",X"00",X"CD",X"E4",X"2B",X"FD",X"23",X"FD",X"23",X"FD",
		X"23",X"10",X"F5",X"C9",X"FD",X"CB",X"00",X"46",X"C8",X"DD",X"21",X"00",X"84",X"0E",X"04",X"D9",
		X"CD",X"FA",X"2B",X"D9",X"DD",X"19",X"0D",X"20",X"F6",X"C9",X"DD",X"CB",X"00",X"46",X"C8",X"FD",
		X"7E",X"01",X"DD",X"96",X"03",X"FE",X"09",X"D0",X"FD",X"7E",X"02",X"DD",X"96",X"04",X"C6",X"04",
		X"FE",X"09",X"D0",X"DD",X"36",X"00",X"00",X"DD",X"36",X"01",X"01",X"DD",X"36",X"02",X"06",X"FD",
		X"36",X"00",X"00",X"11",X"08",X"03",X"FF",X"CD",X"F5",X"36",X"C9",X"FD",X"21",X"0C",X"85",X"06",
		X"03",X"CD",X"3D",X"2C",X"FD",X"23",X"FD",X"23",X"FD",X"23",X"10",X"F5",X"C9",X"FD",X"CB",X"00",
		X"46",X"C8",X"DD",X"21",X"80",X"83",X"DD",X"CB",X"00",X"46",X"C8",X"FD",X"7E",X"01",X"DD",X"96",
		X"03",X"C6",X"03",X"FE",X"07",X"D0",X"FD",X"7E",X"02",X"DD",X"96",X"04",X"C6",X"04",X"FE",X"14",
		X"D0",X"C3",X"49",X"2B",X"3A",X"1D",X"81",X"E6",X"20",X"C8",X"FD",X"21",X"00",X"85",X"06",X"04",
		X"11",X"20",X"00",X"CD",X"7F",X"2C",X"FD",X"23",X"FD",X"23",X"FD",X"23",X"10",X"F5",X"C9",X"FD",
		X"CB",X"00",X"46",X"C8",X"DD",X"21",X"00",X"84",X"0E",X"04",X"D9",X"CD",X"95",X"2C",X"D9",X"DD",
		X"19",X"0D",X"20",X"F6",X"C9",X"DD",X"CB",X"00",X"46",X"C8",X"FD",X"7E",X"01",X"DD",X"96",X"03",
		X"C6",X"04",X"FE",X"0A",X"D0",X"FD",X"7E",X"02",X"DD",X"96",X"04",X"C6",X"04",X"FE",X"09",X"D0",
		X"FD",X"36",X"00",X"00",X"DD",X"34",X"05",X"3E",X"05",X"DD",X"96",X"05",X"C0",X"DD",X"36",X"05",
		X"00",X"DD",X"36",X"00",X"00",X"DD",X"36",X"01",X"01",X"DD",X"36",X"02",X"06",X"11",X"02",X"03",
		X"FF",X"CD",X"F5",X"36",X"C9",X"FD",X"21",X"00",X"85",X"06",X"04",X"11",X"20",X"00",X"CD",X"EA",
		X"2C",X"FD",X"23",X"FD",X"23",X"FD",X"23",X"10",X"F5",X"C9",X"FD",X"CB",X"00",X"46",X"C8",X"DD",
		X"21",X"80",X"82",X"0E",X"08",X"D9",X"CD",X"00",X"2D",X"D9",X"DD",X"19",X"0D",X"20",X"F6",X"C9",
		X"DD",X"CB",X"00",X"46",X"C8",X"FD",X"7E",X"01",X"DD",X"96",X"03",X"C6",X"08",X"FE",X"0E",X"D0",
		X"FD",X"7E",X"02",X"DD",X"96",X"04",X"C6",X"04",X"FE",X"09",X"D0",X"DD",X"36",X"00",X"00",X"DD",
		X"36",X"01",X"01",X"DD",X"36",X"02",X"06",X"FD",X"36",X"00",X"00",X"DD",X"7E",X"17",X"A7",X"28",
		X"0B",X"3D",X"28",X"10",X"3D",X"28",X"26",X"3D",X"28",X"56",X"18",X"65",X"11",X"01",X"03",X"FF",
		X"CD",X"05",X"37",X"C9",X"3A",X"80",X"83",X"0F",X"30",X"0B",X"21",X"05",X"81",X"7E",X"C6",X"30",
		X"30",X"02",X"3E",X"FF",X"77",X"11",X"03",X"03",X"FF",X"CD",X"D8",X"36",X"C9",X"ED",X"5F",X"E6",
		X"03",X"A7",X"28",X"08",X"3D",X"28",X"05",X"3D",X"28",X"0E",X"18",X"18",X"DD",X"36",X"1A",X"00",
		X"11",X"05",X"03",X"FF",X"CD",X"E0",X"36",X"C9",X"DD",X"36",X"1A",X"01",X"11",X"06",X"03",X"FF",
		X"CD",X"E0",X"36",X"C9",X"DD",X"36",X"1A",X"02",X"11",X"07",X"03",X"FF",X"CD",X"E0",X"36",X"C9",
		X"CD",X"E0",X"36",X"3E",X"0A",X"32",X"0A",X"80",X"32",X"12",X"81",X"3E",X"82",X"32",X"22",X"81",
		X"C9",X"11",X"08",X"03",X"FF",X"CD",X"05",X"37",X"C9",X"3A",X"1D",X"81",X"E6",X"06",X"C8",X"FD",
		X"21",X"00",X"85",X"06",X"04",X"11",X"20",X"00",X"CD",X"C4",X"2D",X"FD",X"23",X"FD",X"23",X"FD",
		X"23",X"10",X"F5",X"C9",X"FD",X"CB",X"00",X"46",X"C8",X"DD",X"21",X"00",X"84",X"0E",X"04",X"D9",
		X"CD",X"DA",X"2D",X"D9",X"DD",X"19",X"0D",X"20",X"F6",X"C9",X"DD",X"CB",X"00",X"46",X"C8",X"FD",
		X"7E",X"01",X"DD",X"96",X"03",X"C6",X"05",X"FE",X"0B",X"D0",X"FD",X"7E",X"02",X"DD",X"96",X"04",
		X"C6",X"03",X"FE",X"07",X"D0",X"DD",X"36",X"00",X"00",X"DD",X"36",X"01",X"01",X"DD",X"36",X"02",
		X"06",X"FD",X"36",X"00",X"00",X"11",X"0A",X"03",X"FF",X"CD",X"05",X"37",X"C9",X"DD",X"21",X"00",
		X"85",X"11",X"03",X"00",X"06",X"07",X"D9",X"CD",X"20",X"2E",X"D9",X"DD",X"19",X"10",X"F7",X"C9",
		X"DD",X"CB",X"00",X"46",X"C8",X"3A",X"16",X"81",X"47",X"DD",X"7E",X"02",X"90",X"E6",X"F8",X"0F",
		X"0F",X"C6",X"C0",X"6F",X"26",X"81",X"7E",X"DD",X"BE",X"01",X"38",X"06",X"2C",X"7E",X"DD",X"BE",
		X"01",X"D8",X"DD",X"36",X"00",X"00",X"C9",X"3A",X"1D",X"81",X"E6",X"F8",X"C8",X"FD",X"21",X"C0",
		X"83",X"06",X"02",X"11",X"20",X"00",X"CD",X"5E",X"2E",X"FD",X"19",X"10",X"F9",X"C9",X"FD",X"CB",
		X"00",X"46",X"C8",X"DD",X"21",X"00",X"84",X"0E",X"04",X"D9",X"CD",X"74",X"2E",X"D9",X"DD",X"19",
		X"0D",X"20",X"F6",X"C9",X"DD",X"CB",X"00",X"46",X"C8",X"FD",X"7E",X"03",X"DD",X"96",X"03",X"C6",
		X"05",X"FE",X"0B",X"D0",X"FD",X"7E",X"04",X"DD",X"96",X"04",X"C6",X"06",X"FE",X"0D",X"D0",X"DD",
		X"36",X"00",X"00",X"DD",X"36",X"01",X"01",X"DD",X"36",X"02",X"06",X"DD",X"36",X"05",X"00",X"FD",
		X"36",X"00",X"00",X"FD",X"36",X"01",X"01",X"FD",X"36",X"02",X"06",X"11",X"08",X"03",X"FF",X"CD",
		X"E8",X"36",X"CD",X"F5",X"36",X"C9",X"FD",X"21",X"C0",X"83",X"06",X"02",X"11",X"20",X"00",X"CD",
		X"C7",X"2E",X"FD",X"19",X"10",X"F9",X"C9",X"FD",X"CB",X"00",X"46",X"C8",X"DD",X"21",X"80",X"82",
		X"0E",X"08",X"D9",X"CD",X"DD",X"2E",X"D9",X"DD",X"19",X"0D",X"20",X"F6",X"C9",X"DD",X"CB",X"00",
		X"46",X"C8",X"FD",X"7E",X"03",X"DD",X"96",X"03",X"C6",X"07",X"FE",X"0E",X"D0",X"FD",X"7E",X"04",
		X"DD",X"96",X"04",X"C6",X"07",X"FE",X"0E",X"D0",X"DD",X"36",X"00",X"00",X"DD",X"36",X"01",X"01",
		X"DD",X"36",X"02",X"06",X"FD",X"36",X"00",X"00",X"FD",X"36",X"01",X"01",X"FD",X"36",X"02",X"06",
		X"CD",X"E8",X"36",X"C3",X"2B",X"2D",X"3A",X"1D",X"81",X"E6",X"02",X"C8",X"FD",X"21",X"00",X"84",
		X"06",X"04",X"11",X"20",X"00",X"CD",X"2D",X"2F",X"FD",X"19",X"10",X"F9",X"C9",X"FD",X"CB",X"00",
		X"46",X"C8",X"DD",X"21",X"80",X"82",X"0E",X"08",X"D9",X"CD",X"43",X"2F",X"D9",X"DD",X"19",X"0D",
		X"20",X"F6",X"C9",X"DD",X"CB",X"00",X"46",X"C8",X"FD",X"7E",X"03",X"DD",X"96",X"03",X"C6",X"07",
		X"FE",X"0E",X"D0",X"FD",X"7E",X"04",X"DD",X"96",X"04",X"C6",X"07",X"FE",X"0E",X"D0",X"DD",X"36",
		X"00",X"00",X"DD",X"36",X"01",X"01",X"DD",X"36",X"02",X"06",X"FD",X"36",X"00",X"00",X"FD",X"36",
		X"01",X"01",X"FD",X"36",X"02",X"06",X"CD",X"E8",X"36",X"DD",X"7E",X"17",X"A7",X"28",X"08",X"3D",
		X"28",X"09",X"3D",X"28",X"0A",X"18",X"0F",X"CD",X"05",X"37",X"C9",X"CD",X"D8",X"36",X"C9",X"DD",
		X"35",X"17",X"CD",X"E0",X"36",X"C9",X"CD",X"E0",X"36",X"3E",X"0A",X"32",X"0A",X"80",X"32",X"12",
		X"81",X"3E",X"82",X"32",X"22",X"81",X"C9",X"3A",X"1D",X"81",X"E6",X"06",X"C8",X"FD",X"21",X"C0",
		X"83",X"06",X"02",X"11",X"20",X"00",X"CD",X"BE",X"2F",X"FD",X"19",X"10",X"F9",X"C9",X"FD",X"CB",
		X"00",X"46",X"C8",X"DD",X"21",X"00",X"84",X"0E",X"04",X"D9",X"CD",X"D4",X"2F",X"D9",X"DD",X"19",
		X"0D",X"20",X"F6",X"C9",X"DD",X"CB",X"00",X"46",X"C8",X"FD",X"7E",X"03",X"DD",X"96",X"03",X"C6",
		X"06",X"FE",X"0D",X"D0",X"FD",X"7E",X"04",X"DD",X"96",X"04",X"C6",X"04",X"FE",X"09",X"D0",X"DD",
		X"36",X"00",X"00",X"DD",X"36",X"01",X"01",X"DD",X"36",X"02",X"06",X"FD",X"36",X"00",X"00",X"FD",
		X"36",X"01",X"01",X"FD",X"36",X"02",X"06",X"11",X"0A",X"03",X"FF",X"CD",X"E8",X"36",X"CD",X"05",
		X"37",X"C9",X"DD",X"21",X"C0",X"83",X"06",X"02",X"11",X"20",X"00",X"D9",X"CD",X"25",X"30",X"D9",
		X"DD",X"19",X"10",X"F7",X"C9",X"DD",X"CB",X"00",X"46",X"C8",X"3A",X"16",X"81",X"47",X"DD",X"7E",
		X"04",X"90",X"E6",X"F8",X"0F",X"0F",X"C6",X"C0",X"6F",X"26",X"81",X"7E",X"DD",X"BE",X"03",X"38",
		X"06",X"2C",X"7E",X"DD",X"BE",X"03",X"D8",X"DD",X"36",X"00",X"00",X"DD",X"36",X"01",X"01",X"DD",
		X"36",X"02",X"06",X"CD",X"E8",X"36",X"C9",X"3A",X"1D",X"81",X"E6",X"06",X"C8",X"DD",X"21",X"00",
		X"84",X"06",X"04",X"11",X"20",X"00",X"D9",X"CD",X"70",X"30",X"D9",X"DD",X"19",X"10",X"F7",X"C9",
		X"DD",X"CB",X"00",X"46",X"C8",X"3A",X"16",X"81",X"47",X"DD",X"7E",X"04",X"90",X"E6",X"F8",X"0F",
		X"0F",X"C6",X"C0",X"6F",X"26",X"81",X"7E",X"DD",X"BE",X"03",X"38",X"0B",X"2C",X"7E",X"FE",X"29",
		X"D8",X"C6",X"04",X"DD",X"BE",X"03",X"D8",X"DD",X"36",X"00",X"00",X"DD",X"36",X"01",X"01",X"DD",
		X"36",X"02",X"06",X"CD",X"05",X"37",X"C9",X"3A",X"06",X"80",X"0F",X"38",X"19",X"3A",X"80",X"83",
		X"0F",X"30",X"19",X"3A",X"5F",X"82",X"E6",X"67",X"CC",X"3C",X"31",X"3A",X"5F",X"82",X"E6",X"3F",
		X"CC",X"7F",X"34",X"C3",X"CC",X"30",X"CD",X"55",X"34",X"CD",X"12",X"31",X"CD",X"6E",X"32",X"CD",
		X"4C",X"33",X"CD",X"B3",X"33",X"CD",X"FB",X"33",X"CD",X"AA",X"32",X"CD",X"5F",X"31",X"C3",X"EA",
		X"30",X"CD",X"55",X"34",X"CD",X"12",X"31",X"C3",X"EA",X"30",X"3A",X"1A",X"81",X"47",X"E6",X"07",
		X"C8",X"B8",X"28",X"12",X"32",X"1A",X"81",X"4F",X"78",X"E6",X"F8",X"0F",X"0F",X"0F",X"ED",X"44",
		X"21",X"1B",X"81",X"86",X"77",X"79",X"3D",X"EF",X"D6",X"34",X"A4",X"34",X"08",X"35",X"3A",X"35",
		X"6B",X"35",X"3A",X"06",X"80",X"0F",X"D0",X"3A",X"80",X"83",X"0F",X"D0",X"3A",X"0D",X"80",X"0F",
		X"38",X"0E",X"3A",X"10",X"80",X"CB",X"5F",X"C8",X"3A",X"13",X"80",X"CB",X"5F",X"C0",X"18",X"0C",
		X"3A",X"11",X"80",X"CB",X"5F",X"C8",X"3A",X"14",X"80",X"CB",X"5F",X"C0",X"21",X"00",X"85",X"06",
		X"04",X"CB",X"46",X"20",X"14",X"CB",X"C6",X"2C",X"3A",X"83",X"83",X"C6",X"02",X"77",X"2C",X"3A",
		X"84",X"83",X"D6",X"07",X"77",X"CD",X"0D",X"37",X"C9",X"2C",X"2C",X"2C",X"10",X"E3",X"C9",X"3A",
		X"1D",X"81",X"E6",X"90",X"20",X"6F",X"3A",X"5F",X"82",X"E6",X"27",X"C0",X"3A",X"1D",X"81",X"0F",
		X"38",X"13",X"21",X"27",X"81",X"34",X"7E",X"47",X"E6",X"3C",X"C0",X"78",X"2F",X"E6",X"03",X"20",
		X"04",X"3E",X"10",X"80",X"77",X"3A",X"80",X"83",X"0F",X"D0",X"DD",X"21",X"80",X"82",X"11",X"20",
		X"00",X"06",X"08",X"DD",X"CB",X"00",X"46",X"20",X"05",X"DD",X"19",X"10",X"F6",X"C9",X"DD",X"7E",
		X"17",X"CB",X"47",X"20",X"F4",X"B7",X"28",X"F1",X"3A",X"A4",X"83",X"DD",X"96",X"04",X"FE",X"80",
		X"30",X"E7",X"21",X"0C",X"85",X"06",X"04",X"CB",X"46",X"20",X"14",X"CB",X"C6",X"2C",X"DD",X"7E",
		X"03",X"C6",X"FD",X"77",X"2C",X"DD",X"7E",X"04",X"C6",X"03",X"77",X"CD",X"CB",X"37",X"C9",X"2C",
		X"2C",X"2C",X"10",X"E3",X"C9",X"FA",X"20",X"32",X"3A",X"80",X"83",X"0F",X"D0",X"3A",X"5F",X"82",
		X"E6",X"2F",X"C0",X"DD",X"21",X"00",X"84",X"11",X"20",X"00",X"06",X"04",X"DD",X"CB",X"00",X"46",
		X"20",X"05",X"DD",X"19",X"10",X"F6",X"C9",X"3A",X"A4",X"83",X"DD",X"96",X"04",X"38",X"F3",X"21",
		X"0C",X"85",X"06",X"04",X"CB",X"46",X"20",X"12",X"CB",X"C6",X"2C",X"DD",X"7E",X"03",X"77",X"2C",
		X"DD",X"7E",X"04",X"C6",X"08",X"77",X"CD",X"0D",X"37",X"C9",X"2C",X"2C",X"2C",X"10",X"E5",X"C9",
		X"3A",X"80",X"83",X"0F",X"D0",X"3A",X"5F",X"82",X"E6",X"27",X"C0",X"DD",X"21",X"00",X"84",X"11",
		X"20",X"00",X"06",X"04",X"DD",X"CB",X"00",X"46",X"20",X"07",X"DD",X"19",X"10",X"F6",X"C3",X"8A",
		X"31",X"3A",X"A4",X"83",X"DD",X"96",X"04",X"FE",X"80",X"30",X"EF",X"21",X"0C",X"85",X"06",X"04",
		X"CB",X"46",X"20",X"14",X"CB",X"C6",X"2C",X"DD",X"7E",X"03",X"C6",X"FD",X"77",X"2C",X"DD",X"7E",
		X"04",X"C6",X"03",X"77",X"CD",X"CB",X"37",X"C9",X"2C",X"2C",X"2C",X"10",X"E3",X"C9",X"3A",X"1D",
		X"81",X"E6",X"18",X"C8",X"3A",X"5F",X"82",X"E6",X"3F",X"C0",X"DD",X"21",X"00",X"84",X"11",X"20",
		X"00",X"06",X"04",X"DD",X"7E",X"00",X"DD",X"B6",X"01",X"0F",X"30",X"05",X"DD",X"19",X"10",X"F3",
		X"C9",X"DD",X"36",X"00",X"01",X"DD",X"36",X"01",X"00",X"DD",X"36",X"02",X"00",X"ED",X"5F",X"E6",
		X"0F",X"C6",X"09",X"DD",X"77",X"04",X"CD",X"14",X"33",X"C9",X"3A",X"1D",X"81",X"B7",X"F0",X"3A",
		X"5F",X"82",X"E6",X"1F",X"C0",X"ED",X"5F",X"0F",X"D8",X"DD",X"21",X"80",X"82",X"11",X"20",X"00",
		X"06",X"08",X"DD",X"CB",X"00",X"46",X"20",X"05",X"DD",X"19",X"10",X"F6",X"C9",X"DD",X"7E",X"17",
		X"FE",X"04",X"20",X"F4",X"3A",X"84",X"83",X"DD",X"96",X"04",X"FE",X"50",X"30",X"EA",X"FD",X"21",
		X"00",X"84",X"06",X"04",X"FD",X"7E",X"00",X"FD",X"B6",X"01",X"0F",X"30",X"05",X"FD",X"19",X"10",
		X"F3",X"C9",X"DD",X"36",X"02",X"03",X"DD",X"7E",X"03",X"FD",X"77",X"03",X"DD",X"7E",X"04",X"FD",
		X"77",X"04",X"AF",X"FD",X"77",X"01",X"FD",X"77",X"02",X"FD",X"77",X"0B",X"3C",X"FD",X"77",X"00",
		X"DD",X"77",X"00",X"C9",X"3A",X"16",X"81",X"47",X"DD",X"7E",X"04",X"90",X"E6",X"F8",X"0F",X"0F",
		X"C6",X"C0",X"6F",X"26",X"81",X"ED",X"5F",X"CB",X"47",X"28",X"08",X"7E",X"2C",X"86",X"1F",X"DD",
		X"77",X"03",X"C9",X"CB",X"4F",X"28",X"0B",X"7E",X"47",X"2C",X"86",X"1F",X"80",X"1F",X"DD",X"77",
		X"03",X"C9",X"7E",X"2C",X"86",X"1F",X"86",X"1F",X"DD",X"77",X"03",X"C9",X"3A",X"1D",X"81",X"E6",
		X"06",X"C8",X"3A",X"5F",X"82",X"E6",X"1F",X"C0",X"ED",X"5F",X"0F",X"D8",X"DD",X"21",X"80",X"82",
		X"11",X"20",X"00",X"06",X"08",X"DD",X"CB",X"00",X"46",X"20",X"05",X"DD",X"19",X"10",X"F6",X"C9",
		X"DD",X"7E",X"17",X"A7",X"20",X"F5",X"3A",X"A4",X"83",X"C6",X"10",X"DD",X"96",X"04",X"FE",X"90",
		X"30",X"E9",X"FD",X"21",X"00",X"84",X"06",X"04",X"FD",X"7E",X"00",X"FD",X"B6",X"01",X"0F",X"30",
		X"05",X"FD",X"19",X"10",X"F3",X"C9",X"DD",X"36",X"02",X"03",X"DD",X"7E",X"03",X"FD",X"77",X"03",
		X"DD",X"7E",X"04",X"FD",X"77",X"04",X"FD",X"36",X"00",X"01",X"FD",X"36",X"01",X"00",X"FD",X"36",
		X"02",X"00",X"C9",X"3A",X"1D",X"81",X"E6",X"20",X"C8",X"3A",X"5F",X"82",X"E6",X"0F",X"C0",X"DD",
		X"21",X"00",X"84",X"11",X"20",X"00",X"06",X"04",X"DD",X"7E",X"00",X"DD",X"B6",X"01",X"0F",X"30",
		X"05",X"DD",X"19",X"10",X"F3",X"C9",X"DD",X"36",X"00",X"01",X"DD",X"36",X"01",X"00",X"DD",X"36",
		X"02",X"00",X"ED",X"5F",X"E6",X"7F",X"C6",X"30",X"21",X"83",X"83",X"86",X"1F",X"FE",X"B0",X"38",
		X"02",X"3E",X"B0",X"DD",X"77",X"03",X"DD",X"36",X"04",X"08",X"C9",X"3A",X"1D",X"81",X"E6",X"40",
		X"C8",X"3A",X"5F",X"82",X"67",X"E6",X"4F",X"C0",X"DD",X"21",X"00",X"84",X"11",X"20",X"00",X"06",
		X"04",X"DD",X"7E",X"00",X"DD",X"B6",X"01",X"0F",X"30",X"05",X"DD",X"19",X"10",X"F3",X"C9",X"DD",
		X"36",X"00",X"01",X"AF",X"DD",X"77",X"01",X"DD",X"77",X"02",X"DD",X"36",X"04",X"08",X"DD",X"77",
		X"0E",X"3E",X"30",X"A4",X"0F",X"0F",X"0F",X"0F",X"21",X"51",X"34",X"5F",X"19",X"3A",X"83",X"83",
		X"FE",X"9C",X"38",X"02",X"3E",X"9C",X"FE",X"44",X"30",X"02",X"3E",X"44",X"86",X"DD",X"77",X"03",
		X"C9",X"FC",X"EC",X"14",X"04",X"3A",X"06",X"80",X"0F",X"D0",X"3A",X"80",X"83",X"0F",X"D0",X"3A",
		X"0D",X"80",X"0F",X"38",X"0E",X"3A",X"10",X"80",X"CB",X"4F",X"C8",X"3A",X"13",X"80",X"CB",X"4F",
		X"C0",X"18",X"0C",X"3A",X"11",X"80",X"CB",X"57",X"C8",X"3A",X"14",X"80",X"CB",X"57",X"C0",X"21",
		X"C0",X"83",X"11",X"1F",X"00",X"06",X"02",X"7E",X"2C",X"B6",X"0F",X"30",X"04",X"19",X"10",X"F7",
		X"C9",X"2D",X"36",X"01",X"2C",X"36",X"00",X"2C",X"36",X"00",X"CD",X"12",X"37",X"C9",X"3A",X"1A",
		X"81",X"E6",X"02",X"C8",X"DD",X"21",X"80",X"82",X"11",X"20",X"00",X"06",X"08",X"DD",X"7E",X"00",
		X"DD",X"B6",X"01",X"0F",X"30",X"05",X"DD",X"19",X"10",X"F3",X"C9",X"DD",X"36",X"00",X"01",X"DD",
		X"36",X"01",X"00",X"DD",X"36",X"02",X"00",X"DD",X"36",X"17",X"01",X"AF",X"32",X"1A",X"81",X"C9",
		X"3A",X"1A",X"81",X"E6",X"01",X"C8",X"DD",X"21",X"80",X"82",X"11",X"20",X"00",X"06",X"08",X"DD",
		X"7E",X"00",X"DD",X"B6",X"01",X"0F",X"30",X"05",X"DD",X"19",X"10",X"F3",X"C9",X"DD",X"36",X"00",
		X"01",X"DD",X"36",X"01",X"00",X"DD",X"36",X"02",X"00",X"DD",X"36",X"17",X"00",X"AF",X"32",X"1A",
		X"81",X"C9",X"3A",X"1A",X"81",X"E6",X"04",X"C8",X"DD",X"21",X"80",X"82",X"11",X"20",X"00",X"06",
		X"08",X"DD",X"7E",X"00",X"DD",X"B6",X"01",X"0F",X"30",X"05",X"DD",X"19",X"10",X"F3",X"C9",X"DD",
		X"36",X"00",X"01",X"DD",X"36",X"01",X"00",X"DD",X"36",X"02",X"00",X"DD",X"36",X"17",X"02",X"AF",
		X"32",X"1A",X"81",X"C9",X"3A",X"1A",X"81",X"E6",X"08",X"C8",X"3A",X"12",X"81",X"0F",X"D0",X"DD",
		X"21",X"80",X"82",X"11",X"20",X"00",X"06",X"08",X"DD",X"7E",X"00",X"DD",X"B6",X"01",X"0F",X"30",
		X"05",X"DD",X"19",X"10",X"F3",X"C9",X"DD",X"36",X"00",X"01",X"DD",X"36",X"01",X"00",X"DD",X"36",
		X"02",X"00",X"DD",X"36",X"17",X"03",X"AF",X"32",X"1A",X"81",X"C9",X"DD",X"21",X"80",X"82",X"11",
		X"20",X"00",X"06",X"08",X"DD",X"7E",X"00",X"DD",X"B6",X"01",X"0F",X"30",X"05",X"DD",X"19",X"10",
		X"F3",X"C9",X"DD",X"36",X"00",X"01",X"DD",X"36",X"01",X"00",X"DD",X"36",X"02",X"00",X"DD",X"36",
		X"17",X"04",X"AF",X"32",X"1A",X"81",X"C9",X"CD",X"9E",X"35",X"CD",X"11",X"36",X"C9",X"2A",X"18",
		X"81",X"7E",X"FE",X"FF",X"C0",X"21",X"26",X"81",X"36",X"00",X"2A",X"20",X"81",X"5E",X"23",X"56",
		X"23",X"22",X"20",X"81",X"ED",X"53",X"18",X"81",X"BA",X"C0",X"3A",X"12",X"81",X"0F",X"38",X"0E",
		X"3E",X"0A",X"32",X"0A",X"80",X"32",X"26",X"81",X"3E",X"82",X"32",X"22",X"81",X"C9",X"21",X"D0",
		X"38",X"11",X"B7",X"5B",X"22",X"20",X"81",X"ED",X"53",X"18",X"81",X"3E",X"10",X"32",X"26",X"81",
		X"C9",X"11",X"02",X"07",X"FF",X"21",X"21",X"38",X"3A",X"1E",X"81",X"47",X"87",X"80",X"5F",X"16",
		X"00",X"19",X"5E",X"23",X"56",X"23",X"3A",X"00",X"81",X"B7",X"7E",X"28",X"02",X"CB",X"C7",X"32",
		X"1D",X"81",X"EB",X"7E",X"32",X"18",X"81",X"23",X"7E",X"32",X"19",X"81",X"23",X"22",X"20",X"81",
		X"C9",X"3A",X"5F",X"82",X"A7",X"C0",X"21",X"1B",X"80",X"34",X"7E",X"0F",X"D8",X"21",X"17",X"81",
		X"7E",X"3C",X"E6",X"07",X"FE",X"01",X"28",X"03",X"77",X"18",X"02",X"3C",X"77",X"47",X"3A",X"11",
		X"81",X"0F",X"38",X"13",X"78",X"21",X"4F",X"36",X"16",X"00",X"87",X"5F",X"19",X"7E",X"32",X"04",
		X"A8",X"23",X"7E",X"32",X"03",X"A8",X"C9",X"AF",X"32",X"04",X"A8",X"32",X"03",X"A8",X"C9",X"01",
		X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"01",X"01",X"01",X"01",X"00",X"01",X"00",X"11",
		X"41",X"82",X"1A",X"6F",X"26",X"82",X"7E",X"FE",X"FF",X"C8",X"47",X"3A",X"06",X"80",X"A7",X"78",
		X"C4",X"BC",X"36",X"36",X"FF",X"7D",X"FE",X"5E",X"28",X"03",X"3C",X"12",X"C9",X"3E",X"43",X"12",
		X"C9",X"C5",X"D5",X"E5",X"47",X"11",X"40",X"82",X"1A",X"6F",X"26",X"82",X"70",X"7D",X"FE",X"5E",
		X"28",X"04",X"3C",X"12",X"18",X"03",X"3E",X"43",X"12",X"E1",X"D1",X"C1",X"C9",X"3A",X"42",X"82",
		X"F6",X"10",X"32",X"42",X"82",X"32",X"01",X"A0",X"AF",X"C3",X"BC",X"36",X"AF",X"CD",X"BC",X"36",
		X"3A",X"42",X"82",X"E6",X"EF",X"32",X"42",X"82",X"32",X"01",X"A0",X"C9",X"32",X"00",X"A0",X"3A",
		X"42",X"82",X"E6",X"F7",X"32",X"01",X"A0",X"00",X"00",X"00",X"00",X"3A",X"42",X"82",X"F6",X"08",
		X"32",X"01",X"A0",X"C9",X"3E",X"08",X"18",X"E4",X"3E",X"01",X"CD",X"81",X"36",X"C3",X"40",X"37",
		X"3E",X"01",X"CD",X"81",X"36",X"C3",X"40",X"37",X"3E",X"30",X"CD",X"81",X"36",X"3E",X"02",X"CD",
		X"81",X"36",X"C3",X"40",X"37",X"3E",X"04",X"CD",X"81",X"36",X"C3",X"40",X"37",X"3E",X"05",X"CD",
		X"81",X"36",X"C3",X"40",X"37",X"3E",X"03",X"CD",X"81",X"36",X"C3",X"40",X"37",X"3E",X"06",X"C3",
		X"81",X"36",X"3E",X"20",X"C3",X"81",X"36",X"C9",X"3E",X"0A",X"C3",X"81",X"36",X"3E",X"09",X"CD",
		X"81",X"36",X"3E",X"0A",X"C3",X"81",X"36",X"3E",X"0C",X"CD",X"81",X"36",X"3E",X"0D",X"CD",X"81",
		X"36",X"3E",X"0E",X"C3",X"81",X"36",X"3E",X"0F",X"CD",X"81",X"36",X"3E",X"10",X"C3",X"81",X"36",
		X"3E",X"13",X"CD",X"81",X"36",X"3E",X"14",X"CD",X"81",X"36",X"3E",X"15",X"C3",X"81",X"36",X"3A",
		X"42",X"82",X"F6",X"40",X"B0",X"32",X"42",X"82",X"32",X"01",X"A0",X"C9",X"3A",X"42",X"82",X"E6",
		X"BF",X"32",X"42",X"82",X"32",X"01",X"A0",X"AF",X"32",X"1C",X"80",X"C9",X"3E",X"32",X"CD",X"81",
		X"36",X"3E",X"38",X"CD",X"81",X"36",X"3E",X"29",X"C3",X"81",X"36",X"3E",X"39",X"CD",X"81",X"36",
		X"3E",X"38",X"CD",X"81",X"36",X"3E",X"22",X"C3",X"81",X"36",X"3E",X"32",X"CD",X"81",X"36",X"3E",
		X"39",X"CD",X"81",X"36",X"3E",X"28",X"C3",X"81",X"36",X"3E",X"32",X"CD",X"81",X"36",X"3E",X"38",
		X"CD",X"81",X"36",X"3E",X"39",X"C3",X"81",X"36",X"3E",X"21",X"C3",X"81",X"36",X"3E",X"07",X"C3",
		X"81",X"36",X"3E",X"23",X"C3",X"81",X"36",X"00",X"00",X"00",X"00",X"00",X"3E",X"24",X"C3",X"81",
		X"36",X"3E",X"11",X"C3",X"81",X"36",X"3E",X"25",X"C3",X"81",X"36",X"3E",X"16",X"C3",X"81",X"36",
		X"3E",X"26",X"C3",X"81",X"36",X"3E",X"27",X"C3",X"81",X"36",X"3A",X"80",X"83",X"0F",X"D0",X"3A",
		X"5F",X"82",X"E6",X"3F",X"C0",X"3A",X"05",X"81",X"FE",X"50",X"DC",X"AD",X"37",X"3A",X"1D",X"81",
		X"CB",X"6F",X"C4",X"B2",X"37",X"3A",X"1D",X"81",X"E6",X"58",X"CA",X"6C",X"37",X"CB",X"67",X"C2",
		X"D0",X"37",X"3A",X"5F",X"82",X"E6",X"7F",X"CA",X"A8",X"37",X"C9",X"3A",X"5F",X"82",X"E6",X"3F",
		X"C0",X"3A",X"05",X"81",X"FE",X"50",X"DC",X"AD",X"37",X"C3",X"6C",X"37",X"3E",X"08",X"C3",X"81",
		X"36",X"44",X"38",X"04",X"52",X"38",X"02",X"6E",X"38",X"40",X"60",X"38",X"08",X"7C",X"38",X"06",
		X"8C",X"38",X"81",X"9A",X"38",X"20",X"A4",X"38",X"11",X"B2",X"38",X"02",X"C2",X"38",X"04",X"CC",
		X"38",X"03",X"FF",X"FF",X"A1",X"43",X"A8",X"4E",X"A3",X"49",X"09",X"54",X"53",X"42",X"85",X"50",
		X"FF",X"FF",X"DC",X"51",X"11",X"4E",X"A3",X"49",X"05",X"41",X"C9",X"3F",X"D6",X"4F",X"FF",X"FF",
		X"D6",X"4F",X"85",X"50",X"C9",X"3F",X"C4",X"48",X"7A",X"4D",X"6D",X"4B",X"FF",X"FF",X"4C",X"4C",
		X"E3",X"4C",X"7A",X"4D",X"11",X"4E",X"A8",X"4E",X"3F",X"4F",X"FF",X"FF",X"2D",X"55",X"E0",X"44",
		X"2D",X"55",X"2E",X"46",X"2D",X"55",X"7C",X"47",X"2D",X"55",X"FF",X"FF",X"D2",X"38",X"2A",X"53",
		X"B1",X"39",X"2A",X"53",X"DB",X"3A",X"1D",X"3C",X"FF",X"FF",X"7A",X"4D",X"4C",X"4C",X"3F",X"4F",
		X"E3",X"4C",X"FF",X"FF",X"8E",X"4A",X"6D",X"4B",X"53",X"42",X"C9",X"3F",X"7A",X"4D",X"C4",X"48",
		X"FF",X"FF",X"A3",X"49",X"2C",X"3D",X"0B",X"3E",X"EA",X"3E",X"0B",X"3E",X"EA",X"3E",X"2C",X"3D",
		X"FF",X"FF",X"2A",X"56",X"66",X"57",X"63",X"58",X"72",X"59",X"FF",X"FF",X"E4",X"5A",X"B7",X"5B",
		X"FF",X"FF",X"C8",X"36",X"C8",X"36",X"00",X"00",X"C8",X"36",X"C0",X"30",X"00",X"00",X"B8",X"33",
		X"B0",X"32",X"00",X"00",X"A8",X"31",X"A0",X"33",X"00",X"00",X"98",X"30",X"90",X"33",X"00",X"00",
		X"88",X"30",X"80",X"32",X"00",X"00",X"80",X"36",X"80",X"36",X"00",X"01",X"80",X"36",X"78",X"31",
		X"00",X"00",X"70",X"33",X"68",X"30",X"00",X"00",X"60",X"34",X"68",X"2C",X"00",X"00",X"70",X"2C",
		X"78",X"2D",X"00",X"00",X"80",X"2E",X"88",X"2C",X"00",X"00",X"90",X"36",X"90",X"36",X"00",X"02",
		X"90",X"36",X"90",X"36",X"00",X"02",X"90",X"36",X"90",X"36",X"00",X"01",X"90",X"36",X"90",X"36",
		X"00",X"05",X"88",X"31",X"80",X"30",X"00",X"00",X"78",X"33",X"70",X"32",X"00",X"00",X"70",X"2E",
		X"78",X"2D",X"00",X"00",X"80",X"2C",X"88",X"2D",X"00",X"00",X"90",X"2F",X"98",X"2D",X"00",X"00",
		X"A0",X"2E",X"A8",X"2C",X"00",X"00",X"B0",X"2F",X"B8",X"2C",X"00",X"00",X"C0",X"36",X"C0",X"36",
		X"00",X"05",X"C0",X"36",X"C0",X"36",X"00",X"02",X"B8",X"31",X"B0",X"30",X"00",X"00",X"A8",X"33",
		X"A0",X"32",X"00",X"00",X"A0",X"2E",X"A8",X"2C",X"00",X"00",X"B0",X"2E",X"B8",X"2C",X"00",X"00",
		X"C0",X"2D",X"C8",X"2F",X"00",X"00",X"D0",X"2F",X"D8",X"2C",X"00",X"00",X"E0",X"36",X"E0",X"36",
		X"00",X"01",X"E0",X"36",X"E0",X"36",X"00",X"05",X"E0",X"36",X"D8",X"31",X"00",X"00",X"D0",X"33",
		X"C8",X"32",X"00",X"00",X"C8",X"36",X"C8",X"36",X"00",X"00",X"C8",X"36",X"C8",X"36",X"00",X"00",
		X"FF",X"C8",X"36",X"C8",X"36",X"00",X"00",X"C8",X"36",X"C8",X"36",X"00",X"00",X"C8",X"36",X"C8",
		X"36",X"00",X"00",X"C8",X"36",X"C8",X"36",X"00",X"00",X"C0",X"31",X"B8",X"31",X"00",X"00",X"B0",
		X"33",X"A8",X"30",X"00",X"00",X"A0",X"30",X"98",X"31",X"28",X"5F",X"28",X"62",X"00",X"90",X"33",
		X"88",X"30",X"30",X"63",X"38",X"62",X"00",X"80",X"32",X"80",X"2E",X"40",X"63",X"48",X"63",X"00",
		X"88",X"2F",X"90",X"2D",X"50",X"62",X"58",X"63",X"00",X"98",X"2C",X"A0",X"2D",X"60",X"62",X"68",
		X"63",X"00",X"A8",X"36",X"A8",X"36",X"70",X"5C",X"68",X"61",X"02",X"A8",X"36",X"A8",X"36",X"60",
		X"60",X"58",X"60",X"01",X"A0",X"31",X"98",X"30",X"50",X"61",X"50",X"63",X"00",X"90",X"30",X"90",
		X"2C",X"58",X"63",X"60",X"63",X"00",X"98",X"2D",X"A0",X"36",X"60",X"61",X"60",X"62",X"00",X"A0",
		X"36",X"A0",X"36",X"68",X"62",X"70",X"5C",X"01",X"98",X"33",X"90",X"31",X"68",X"61",X"60",X"60",
		X"00",X"88",X"34",X"90",X"36",X"58",X"5D",X"60",X"62",X"00",X"90",X"36",X"90",X"36",X"68",X"63",
		X"68",X"60",X"02",X"90",X"36",X"90",X"36",X"60",X"60",X"58",X"60",X"05",X"88",X"31",X"80",X"30",
		X"50",X"61",X"48",X"61",X"00",X"78",X"32",X"78",X"2E",X"40",X"60",X"38",X"60",X"00",X"80",X"2F",
		X"88",X"2D",X"30",X"61",X"30",X"5F",X"00",X"90",X"2C",X"90",X"37",X"30",X"62",X"38",X"63",X"00",
		X"98",X"36",X"98",X"36",X"40",X"63",X"48",X"62",X"01",X"98",X"36",X"90",X"30",X"50",X"63",X"58",
		X"62",X"00",X"90",X"36",X"90",X"36",X"58",X"60",X"50",X"61",X"02",X"88",X"30",X"80",X"33",X"48",
		X"61",X"40",X"61",X"00",X"78",X"31",X"70",X"32",X"38",X"60",X"30",X"60",X"00",X"70",X"2E",X"78",
		X"2C",X"28",X"61",X"28",X"5F",X"00",X"80",X"2D",X"88",X"2E",X"00",X"00",X"90",X"2F",X"98",X"2C",
		X"00",X"00",X"A0",X"2C",X"A8",X"2D",X"00",X"00",X"B0",X"2E",X"B8",X"2C",X"00",X"00",X"C0",X"2C",
		X"C8",X"36",X"00",X"00",X"C8",X"36",X"C8",X"36",X"00",X"00",X"FF",X"C8",X"36",X"C8",X"36",X"00",
		X"00",X"C8",X"36",X"C8",X"36",X"28",X"5F",X"28",X"62",X"02",X"C0",X"30",X"B8",X"30",X"30",X"62",
		X"38",X"63",X"00",X"B0",X"33",X"A8",X"31",X"40",X"63",X"48",X"62",X"00",X"A0",X"32",X"A0",X"2E",
		X"50",X"62",X"58",X"62",X"00",X"A8",X"2C",X"B0",X"2F",X"60",X"62",X"68",X"63",X"00",X"B8",X"2D",
		X"C0",X"2F",X"70",X"63",X"78",X"62",X"00",X"C8",X"2F",X"D0",X"2D",X"80",X"62",X"88",X"63",X"00",
		X"D8",X"36",X"D8",X"36",X"90",X"63",X"98",X"62",X"05",X"D8",X"36",X"D8",X"36",X"A0",X"62",X"A8",
		X"5C",X"05",X"D8",X"36",X"D8",X"36",X"A0",X"60",X"98",X"61",X"02",X"D8",X"36",X"D8",X"36",X"90",
		X"60",X"88",X"60",X"01",X"D0",X"31",X"C8",X"30",X"80",X"61",X"78",X"61",X"00",X"C0",X"32",X"B8",
		X"31",X"70",X"60",X"68",X"60",X"00",X"B0",X"33",X"A8",X"33",X"60",X"61",X"58",X"5D",X"00",X"A0",
		X"30",X"98",X"32",X"60",X"62",X"68",X"63",X"00",X"98",X"2E",X"A0",X"2F",X"68",X"61",X"60",X"60",
		X"00",X"A8",X"2D",X"A8",X"37",X"58",X"60",X"50",X"61",X"00",X"B0",X"36",X"B0",X"36",X"48",X"60",
		X"40",X"61",X"02",X"B0",X"36",X"B0",X"36",X"38",X"61",X"38",X"63",X"05",X"A8",X"37",X"A8",X"31",
		X"40",X"62",X"48",X"63",X"00",X"A0",X"31",X"98",X"30",X"50",X"62",X"58",X"5C",X"00",X"90",X"31",
		X"88",X"33",X"50",X"60",X"48",X"61",X"00",X"80",X"30",X"78",X"30",X"40",X"61",X"38",X"61",X"00",
		X"70",X"31",X"68",X"33",X"30",X"60",X"28",X"60",X"00",X"60",X"32",X"60",X"2E",X"28",X"5F",X"28",
		X"5F",X"00",X"68",X"2F",X"70",X"2D",X"28",X"5F",X"28",X"5F",X"00",X"78",X"2F",X"80",X"2D",X"28",
		X"5F",X"28",X"5F",X"00",X"88",X"2D",X"90",X"2F",X"28",X"62",X"30",X"63",X"00",X"98",X"2F",X"A0",
		X"2C",X"38",X"63",X"40",X"63",X"00",X"A8",X"2C",X"B0",X"2F",X"48",X"62",X"50",X"63",X"00",X"B8",
		X"2F",X"C0",X"2D",X"50",X"60",X"48",X"61",X"00",X"C8",X"2D",X"D0",X"2C",X"40",X"61",X"38",X"60",
		X"00",X"D8",X"36",X"D8",X"36",X"30",X"61",X"28",X"61",X"00",X"D8",X"36",X"D8",X"36",X"00",X"05",
		X"D0",X"31",X"C8",X"32",X"00",X"00",X"C8",X"36",X"C8",X"36",X"00",X"00",X"FF",X"C8",X"36",X"C8",
		X"36",X"00",X"00",X"C8",X"36",X"C0",X"31",X"00",X"00",X"B8",X"33",X"B0",X"30",X"00",X"00",X"A8",
		X"30",X"A0",X"30",X"00",X"00",X"98",X"33",X"90",X"32",X"00",X"00",X"90",X"2E",X"98",X"2F",X"00",
		X"00",X"A0",X"2D",X"A8",X"36",X"28",X"62",X"30",X"62",X"00",X"A8",X"36",X"A8",X"36",X"38",X"63",
		X"40",X"62",X"01",X"A8",X"36",X"A8",X"36",X"48",X"62",X"50",X"63",X"02",X"A8",X"36",X"A8",X"2F",
		X"58",X"63",X"60",X"62",X"00",X"B0",X"2D",X"B8",X"2C",X"68",X"63",X"70",X"63",X"00",X"C0",X"2C",
		X"C0",X"37",X"78",X"63",X"80",X"5C",X"00",X"C8",X"36",X"C8",X"36",X"78",X"60",X"70",X"61",X"05",
		X"C0",X"32",X"C0",X"2E",X"70",X"62",X"78",X"62",X"00",X"C8",X"2F",X"D0",X"2F",X"80",X"63",X"88",
		X"62",X"00",X"D8",X"36",X"D8",X"36",X"90",X"5C",X"88",X"60",X"05",X"D8",X"36",X"D8",X"36",X"80",
		X"60",X"78",X"61",X"02",X"D0",X"37",X"D0",X"33",X"70",X"61",X"68",X"60",X"00",X"C8",X"33",X"C0",
		X"31",X"60",X"60",X"58",X"60",X"00",X"B8",X"31",X"B0",X"30",X"50",X"61",X"48",X"60",X"00",X"A8",
		X"30",X"A0",X"30",X"40",X"60",X"38",X"60",X"00",X"98",X"33",X"90",X"31",X"30",X"61",X"28",X"60",
		X"00",X"88",X"31",X"80",X"31",X"00",X"00",X"78",X"32",X"78",X"2E",X"00",X"00",X"80",X"2C",X"88",
		X"2D",X"00",X"00",X"90",X"2D",X"90",X"37",X"00",X"00",X"98",X"36",X"98",X"36",X"00",X"01",X"98",
		X"36",X"98",X"36",X"00",X"01",X"98",X"36",X"98",X"36",X"00",X"05",X"90",X"31",X"88",X"33",X"00",
		X"00",X"80",X"32",X"80",X"2E",X"00",X"00",X"88",X"2C",X"90",X"2D",X"00",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"60",X"00",X"C0",X"36",X"C0",X"36",X"4F",X"62",X"4C",X"60",X"02",X"C0",X"36",X"C4",X"2C",X"44",
		X"61",X"3C",X"61",X"00",X"C8",X"36",X"C8",X"36",X"3A",X"5F",X"3A",X"5F",X"03",X"C8",X"36",X"C8",
		X"36",X"3A",X"5F",X"3A",X"5F",X"02",X"C8",X"36",X"C4",X"30",X"3C",X"62",X"44",X"62",X"00",X"BC",
		X"33",X"B4",X"31",X"4C",X"63",X"54",X"62",X"00",X"AC",X"30",X"A0",X"34",X"5C",X"62",X"64",X"62",
		X"00",X"AC",X"2D",X"B0",X"36",X"6C",X"63",X"74",X"62",X"00",X"B0",X"36",X"B0",X"36",X"7F",X"63",
		X"7C",X"60",X"01",X"B0",X"36",X"B0",X"36",X"74",X"60",X"77",X"5C",X"01",X"B0",X"36",X"B0",X"36",
		X"6F",X"3A",X"6F",X"3A",X"01",X"B0",X"36",X"B0",X"36",X"6C",X"60",X"64",X"60",X"01",X"B4",X"2C",
		X"BC",X"2D",X"5C",X"61",X"54",X"60",X"00",X"C4",X"2E",X"CC",X"2F",X"52",X"5F",X"52",X"5F",X"00",
		X"D2",X"35",X"CE",X"37",X"4C",X"60",X"44",X"60",X"00",X"C8",X"34",X"D0",X"36",X"3C",X"60",X"34",
		X"61",X"00",X"D0",X"36",X"D0",X"36",X"2C",X"60",X"28",X"10",X"02",X"D0",X"36",X"D0",X"36",X"00",
		X"03",X"D0",X"36",X"D0",X"36",X"00",X"02",X"CC",X"33",X"C4",X"30",X"00",X"00",X"BC",X"31",X"B6",
		X"37",X"00",X"00",X"B8",X"36",X"B8",X"36",X"28",X"10",X"2C",X"62",X"00",X"B8",X"36",X"BC",X"2C",
		X"34",X"62",X"3C",X"63",X"00",X"C4",X"2D",X"C8",X"36",X"44",X"62",X"4F",X"5C",X"00",X"C8",X"36",
		X"C8",X"36",X"44",X"61",X"44",X"63",X"01",X"C8",X"36",X"C4",X"31",X"4F",X"5C",X"44",X"60",X"00",
		X"B8",X"34",X"C4",X"2F",X"44",X"62",X"4F",X"5C",X"00",X"CC",X"2D",X"D0",X"36",X"47",X"3A",X"47",
		X"3A",X"00",X"D0",X"36",X"D0",X"36",X"44",X"61",X"3C",X"60",X"03",X"D0",X"36",X"CC",X"30",X"34",
		X"61",X"2C",X"60",X"00",X"FF",X"C0",X"34",X"CC",X"2C",X"2F",X"5C",X"2F",X"5C",X"00",X"D4",X"2D",
		X"D8",X"36",X"2A",X"5F",X"2C",X"62",X"00",X"D8",X"36",X"D8",X"36",X"34",X"62",X"3C",X"63",X"01",
		X"D8",X"36",X"D8",X"36",X"44",X"63",X"4C",X"62",X"01",X"D8",X"36",X"D8",X"36",X"54",X"63",X"5F",
		X"62",X"01",X"D8",X"36",X"D8",X"36",X"5C",X"61",X"57",X"5E",X"02",X"D4",X"33",X"CC",X"32",X"55",
		X"5D",X"5C",X"63",X"00",X"C4",X"31",X"BC",X"30",X"64",X"62",X"6C",X"63",X"00",X"B4",X"31",X"AC",
		X"33",X"74",X"62",X"7A",X"5F",X"00",X"A4",X"30",X"9C",X"31",X"74",X"60",X"6C",X"61",X"00",X"90",
		X"30",X"92",X"2C",X"64",X"60",X"5C",X"60",X"00",X"94",X"33",X"8C",X"32",X"54",X"61",X"4C",X"60",
		X"00",X"84",X"30",X"7C",X"31",X"44",X"61",X"3E",X"5D",X"00",X"74",X"32",X"68",X"30",X"3C",X"60",
		X"34",X"61",X"00",X"6A",X"2D",X"74",X"2E",X"2E",X"5E",X"32",X"5F",X"00",X"7C",X"2F",X"84",X"2C",
		X"37",X"5C",X"2E",X"5E",X"00",X"88",X"36",X"88",X"36",X"34",X"62",X"3F",X"62",X"01",X"88",X"36",
		X"88",X"36",X"3C",X"61",X"3A",X"5F",X"03",X"88",X"36",X"88",X"36",X"3A",X"5F",X"3A",X"5F",X"02",
		X"88",X"36",X"88",X"36",X"3A",X"5F",X"3C",X"63",X"01",X"8C",X"2C",X"94",X"2D",X"44",X"62",X"47",
		X"3A",X"00",X"90",X"34",X"9A",X"35",X"47",X"3A",X"47",X"3A",X"00",X"9C",X"2C",X"A4",X"2D",X"47",
		X"3A",X"47",X"3A",X"00",X"AC",X"2F",X"B4",X"2E",X"47",X"3A",X"47",X"3A",X"00",X"B8",X"36",X"B8",
		X"36",X"47",X"3A",X"47",X"3A",X"01",X"B8",X"36",X"B8",X"36",X"44",X"60",X"3C",X"61",X"03",X"B8",
		X"36",X"B8",X"36",X"34",X"60",X"2E",X"5E",X"01",X"BA",X"35",X"B0",X"34",X"2E",X"5E",X"2E",X"5E",
		X"00",X"B8",X"36",X"B8",X"36",X"2E",X"5E",X"34",X"62",X"02",X"B4",X"33",X"AC",X"30",X"3C",X"62",
		X"47",X"63",X"00",X"A8",X"36",X"A8",X"36",X"45",X"60",X"3C",X"61",X"01",X"A8",X"36",X"A8",X"36",
		X"34",X"60",X"34",X"62",X"01",X"A8",X"36",X"A8",X"36",X"3F",X"5C",X"37",X"3A",X"01",X"A0",X"34",
		X"A0",X"34",X"37",X"3A",X"34",X"60",X"00",X"A8",X"36",X"A8",X"36",X"2C",X"60",X"2F",X"5C",X"03",
		X"AC",X"2C",X"B4",X"2F",X"2A",X"5F",X"2F",X"62",X"00",X"BC",X"2C",X"C4",X"2F",X"2F",X"61",X"2F",
		X"5C",X"00",X"FF",X"C4",X"30",X"B8",X"30",X"2F",X"62",X"2C",X"60",X"00",X"BA",X"2F",X"C4",X"2E",
		X"2C",X"62",X"34",X"63",X"00",X"CC",X"2C",X"D4",X"2D",X"3F",X"62",X"3C",X"61",X"00",X"D8",X"36",
		X"D8",X"36",X"37",X"5E",X"3C",X"62",X"01",X"D8",X"36",X"D8",X"36",X"44",X"62",X"4C",X"62",X"01",
		X"D4",X"30",X"C8",X"34",X"4C",X"60",X"46",X"5D",X"00",X"D0",X"36",X"D0",X"36",X"4C",X"62",X"54",
		X"62",X"03",X"D0",X"36",X"D0",X"36",X"5C",X"62",X"67",X"5C",X"03",X"CC",X"33",X"C0",X"34",X"5C",
		X"60",X"5C",X"62",X"00",X"C8",X"36",X"C8",X"36",X"5F",X"3A",X"5F",X"3A",X"01",X"C8",X"36",X"C8",
		X"36",X"5F",X"3A",X"5F",X"3A",X"01",X"C4",X"33",X"B8",X"34",X"5F",X"3A",X"5F",X"3A",X"00",X"C0",
		X"36",X"C0",X"36",X"5F",X"3A",X"67",X"5C",X"02",X"C0",X"36",X"C0",X"36",X"5E",X"5D",X"62",X"5F",
		X"02",X"BC",X"30",X"B4",X"31",X"5C",X"60",X"54",X"61",X"00",X"AC",X"33",X"A6",X"37",X"4C",X"60",
		X"44",X"60",X"00",X"AA",X"38",X"A0",X"34",X"3F",X"5E",X"3F",X"5E",X"00",X"AA",X"35",X"A6",X"37",
		X"3F",X"5E",X"3F",X"5E",X"00",X"AC",X"2E",X"B0",X"36",X"3F",X"5E",X"3F",X"5E",X"00",X"B0",X"36",
		X"B0",X"36",X"3F",X"5E",X"3F",X"5E",X"01",X"B0",X"36",X"B0",X"36",X"3F",X"5E",X"3F",X"5E",X"01",
		X"B4",X"2C",X"B8",X"36",X"3F",X"5E",X"3F",X"5E",X"00",X"B8",X"36",X"B8",X"36",X"3F",X"5E",X"3F",
		X"5E",X"03",X"B8",X"36",X"B8",X"36",X"3F",X"5E",X"3F",X"5E",X"03",X"BC",X"2C",X"C0",X"36",X"3F",
		X"5E",X"3F",X"5E",X"00",X"C0",X"36",X"C0",X"36",X"3F",X"5E",X"3F",X"5E",X"01",X"C0",X"36",X"C0",
		X"36",X"44",X"62",X"4F",X"62",X"01",X"B8",X"34",X"C2",X"38",X"4C",X"60",X"47",X"5E",X"00",X"C0",
		X"36",X"C0",X"36",X"44",X"61",X"3C",X"60",X"02",X"C4",X"2E",X"CC",X"2F",X"37",X"5E",X"37",X"5E",
		X"00",X"D4",X"2C",X"DA",X"35",X"37",X"3A",X"37",X"5E",X"00",X"D8",X"36",X"D8",X"36",X"3F",X"62",
		X"3C",X"60",X"01",X"D4",X"31",X"CC",X"30",X"34",X"60",X"2F",X"5E",X"00",X"C4",X"33",X"BC",X"32",
		X"2F",X"5E",X"2F",X"5E",X"00",X"B0",X"30",X"B2",X"2F",X"37",X"5C",X"2E",X"5E",X"00",X"BC",X"2C",
		X"C4",X"2D",X"32",X"5F",X"2C",X"60",X"00",X"CC",X"2F",X"CC",X"33",X"2A",X"5F",X"2A",X"5F",X"00",
		X"FF",X"C4",X"30",X"BC",X"31",X"00",X"00",X"B4",X"32",X"AC",X"33",X"00",X"00",X"A6",X"37",X"AC",
		X"2C",X"28",X"10",X"2C",X"63",X"00",X"B0",X"36",X"B0",X"36",X"34",X"62",X"3F",X"5C",X"01",X"B0",
		X"36",X"B4",X"2C",X"36",X"5E",X"3A",X"5F",X"00",X"B8",X"36",X"B8",X"36",X"3C",X"63",X"44",X"62",
		X"01",X"B8",X"36",X"BC",X"2C",X"4F",X"62",X"4C",X"60",X"00",X"C0",X"36",X"C0",X"36",X"4F",X"62",
		X"4C",X"60",X"02",X"C0",X"36",X"C4",X"2C",X"44",X"61",X"3C",X"61",X"00",X"C8",X"36",X"C8",X"36",
		X"3A",X"5F",X"3A",X"5F",X"03",X"C8",X"36",X"C8",X"36",X"3A",X"5F",X"3A",X"5F",X"02",X"78",X"0E",
		X"78",X"0E",X"3C",X"62",X"44",X"62",X"00",X"88",X"0E",X"88",X"0E",X"4C",X"63",X"57",X"0E",X"00",
		X"88",X"0E",X"88",X"0E",X"4F",X"0E",X"57",X"0E",X"01",X"88",X"0E",X"88",X"0E",X"4F",X"0E",X"57",
		X"0E",X"01",X"88",X"0E",X"88",X"0E",X"4F",X"0E",X"57",X"0E",X"01",X"88",X"0E",X"88",X"0E",X"4F",
		X"0E",X"57",X"0E",X"02",X"88",X"0E",X"80",X"0E",X"4F",X"0E",X"57",X"0E",X"00",X"80",X"0E",X"A0",
		X"0E",X"4F",X"0E",X"57",X"0E",X"00",X"A0",X"0E",X"A0",X"0E",X"4F",X"0E",X"57",X"0E",X"02",X"A0",
		X"0E",X"A0",X"0E",X"4F",X"0E",X"57",X"0E",X"03",X"A0",X"0E",X"A0",X"0E",X"4F",X"0E",X"57",X"0E",
		X"03",X"A0",X"0E",X"A0",X"0E",X"4F",X"0E",X"57",X"0E",X"01",X"BC",X"2C",X"C0",X"36",X"3F",X"5E",
		X"3F",X"5E",X"00",X"C0",X"36",X"C0",X"36",X"3F",X"5E",X"3F",X"5E",X"01",X"C0",X"36",X"C0",X"36",
		X"44",X"62",X"4F",X"62",X"01",X"B8",X"34",X"C2",X"38",X"4C",X"60",X"47",X"5E",X"00",X"C0",X"36",
		X"C0",X"36",X"44",X"61",X"3C",X"60",X"02",X"C4",X"2E",X"CC",X"2F",X"37",X"5E",X"37",X"5E",X"00",
		X"D4",X"2C",X"DA",X"35",X"37",X"3A",X"37",X"5E",X"00",X"D8",X"36",X"D8",X"36",X"3F",X"62",X"3C",
		X"60",X"01",X"D4",X"31",X"CC",X"30",X"34",X"60",X"2F",X"5E",X"00",X"C4",X"33",X"BC",X"32",X"2F",
		X"5E",X"2F",X"5E",X"00",X"B0",X"30",X"B2",X"2F",X"37",X"5C",X"2E",X"5E",X"00",X"BC",X"2C",X"C4",
		X"2D",X"32",X"5F",X"2C",X"60",X"00",X"CC",X"2F",X"CC",X"33",X"2A",X"5F",X"2A",X"5F",X"00",X"FF",
		X"C4",X"30",X"BC",X"31",X"2C",X"62",X"34",X"62",X"00",X"B4",X"32",X"AC",X"33",X"3C",X"63",X"44",
		X"62",X"00",X"A0",X"34",X"AA",X"38",X"4C",X"63",X"54",X"63",X"00",X"A6",X"37",X"AC",X"2C",X"5C",
		X"62",X"64",X"62",X"00",X"B0",X"36",X"B0",X"36",X"6C",X"62",X"77",X"5C",X"02",X"B0",X"36",X"B0",
		X"36",X"6F",X"5E",X"6F",X"5E",X"03",X"B0",X"36",X"B0",X"36",X"6F",X"3A",X"6F",X"3A",X"31",X"B0",
		X"36",X"B0",X"36",X"74",X"62",X"77",X"5E",X"02",X"A8",X"34",X"AE",X"37",X"77",X"5E",X"77",X"5E",
		X"21",X"AC",X"31",X"A4",X"32",X"74",X"60",X"6C",X"61",X"00",X"9C",X"31",X"94",X"33",X"67",X"5E",
		X"67",X"5E",X"19",X"8C",X"30",X"86",X"37",X"67",X"5E",X"67",X"5E",X"09",X"8A",X"35",X"87",X"37",
		X"6C",X"62",X"76",X"5C",X"00",X"86",X"37",X"88",X"38",X"6C",X"61",X"64",X"60",X"00",X"8C",X"2E",
		X"90",X"36",X"61",X"5F",X"5E",X"3A",X"00",X"90",X"38",X"90",X"38",X"61",X"5F",X"5E",X"5E",X"00",
		X"88",X"34",X"92",X"38",X"5C",X"60",X"57",X"5E",X"00",X"92",X"35",X"88",X"34",X"57",X"5E",X"57",
		X"5E",X"21",X"90",X"36",X"90",X"36",X"57",X"5E",X"57",X"5E",X"29",X"90",X"36",X"90",X"36",X"5C",
		X"62",X"64",X"63",X"00",X"90",X"36",X"90",X"36",X"6F",X"5C",X"67",X"5E",X"00",X"90",X"36",X"90",
		X"36",X"67",X"5E",X"67",X"5E",X"19",X"90",X"36",X"90",X"36",X"67",X"5E",X"67",X"5E",X"19",X"90",
		X"36",X"90",X"36",X"64",X"61",X"5C",X"60",X"03",X"88",X"34",X"94",X"2C",X"54",X"60",X"4E",X"3A",
		X"00",X"98",X"38",X"98",X"38",X"51",X"5F",X"4E",X"5D",X"00",X"98",X"38",X"98",X"38",X"4F",X"5E",
		X"4F",X"5E",X"39",X"98",X"38",X"90",X"34",X"4F",X"5E",X"4F",X"5E",X"31",X"98",X"36",X"98",X"36",
		X"4C",X"60",X"44",X"60",X"02",X"9C",X"2C",X"A4",X"2D",X"3F",X"5E",X"3F",X"5E",X"51",X"A8",X"36",
		X"A8",X"36",X"3F",X"5E",X"3F",X"5E",X"59",X"A8",X"36",X"A0",X"34",X"3F",X"5E",X"3F",X"5E",X"51",
		X"A8",X"36",X"A8",X"36",X"3C",X"61",X"34",X"61",X"02",X"A4",X"31",X"98",X"33",X"2F",X"5E",X"2F",
		X"5E",X"59",X"9A",X"2C",X"A4",X"2D",X"2F",X"5E",X"2F",X"5E",X"61",X"AC",X"2E",X"B4",X"2F",X"2C",
		X"60",X"2C",X"63",X"00",X"BC",X"2C",X"C4",X"2D",X"2C",X"60",X"2A",X"5F",X"00",X"FF",X"C4",X"30",
		X"BC",X"32",X"2C",X"62",X"34",X"63",X"00",X"B0",X"31",X"B2",X"2E",X"3C",X"62",X"3F",X"5E",X"00",
		X"BC",X"2D",X"C4",X"2C",X"3F",X"3A",X"3F",X"3A",X"71",X"CC",X"2F",X"D0",X"36",X"3F",X"3A",X"3F",
		X"3A",X"81",X"D0",X"36",X"D0",X"36",X"44",X"62",X"4C",X"63",X"03",X"D0",X"36",X"D0",X"36",X"54",
		X"62",X"5C",X"63",X"00",X"D0",X"36",X"D0",X"36",X"67",X"5C",X"5F",X"3A",X"02",X"D0",X"36",X"D0",
		X"36",X"5F",X"3A",X"5F",X"3A",X"61",X"D0",X"36",X"C8",X"34",X"5F",X"3A",X"5F",X"3A",X"59",X"CC",
		X"31",X"C4",X"30",X"5F",X"3A",X"5F",X"3A",X"51",X"B8",X"33",X"BA",X"2F",X"64",X"62",X"6C",X"62",
		X"00",X"C4",X"2C",X"C0",X"34",X"74",X"63",X"7C",X"63",X"00",X"CA",X"35",X"C8",X"36",X"84",X"62",
		X"8F",X"5C",X"00",X"C8",X"36",X"C8",X"36",X"84",X"60",X"7F",X"3A",X"02",X"C8",X"36",X"C8",X"36",
		X"7F",X"3A",X"7F",X"3A",X"39",X"C8",X"36",X"C8",X"36",X"7F",X"3A",X"7F",X"3A",X"39",X"C8",X"36",
		X"C8",X"36",X"7F",X"3A",X"7F",X"3A",X"39",X"C8",X"36",X"C8",X"36",X"84",X"63",X"8C",X"62",X"03",
		X"C8",X"36",X"C8",X"36",X"97",X"63",X"95",X"60",X"00",X"C8",X"36",X"C8",X"36",X"8F",X"3A",X"8F",
		X"3A",X"29",X"C8",X"36",X"C8",X"36",X"8F",X"3A",X"8F",X"3A",X"29",X"C8",X"36",X"C8",X"36",X"8F",
		X"3A",X"8F",X"3A",X"29",X"CC",X"2C",X"D4",X"2C",X"8C",X"60",X"87",X"3A",X"00",X"D8",X"36",X"D8",
		X"36",X"87",X"3A",X"87",X"3A",X"41",X"D8",X"36",X"D8",X"36",X"87",X"3A",X"87",X"3A",X"41",X"D8",
		X"36",X"D8",X"36",X"87",X"3A",X"8C",X"63",X"03",X"D8",X"36",X"D8",X"36",X"94",X"62",X"9F",X"5C",
		X"03",X"D8",X"36",X"D8",X"36",X"97",X"3A",X"97",X"3A",X"31",X"D8",X"36",X"D8",X"36",X"97",X"3A",
		X"97",X"3A",X"31",X"D4",X"31",X"CC",X"30",X"97",X"3A",X"97",X"3A",X"21",X"C4",X"33",X"BC",X"30",
		X"94",X"60",X"8C",X"60",X"00",X"B0",X"34",X"B8",X"36",X"84",X"61",X"7C",X"60",X"00",X"B8",X"36",
		X"B8",X"36",X"74",X"60",X"6C",X"60",X"03",X"B8",X"36",X"BC",X"2D",X"64",X"61",X"5C",X"61",X"00",
		X"C0",X"36",X"C0",X"36",X"54",X"60",X"4C",X"61",X"02",X"C0",X"36",X"C0",X"36",X"44",X"60",X"3C",
		X"60",X"02",X"C4",X"2C",X"CA",X"35",X"34",X"61",X"2C",X"60",X"00",X"FF",X"C4",X"30",X"BC",X"31",
		X"00",X"00",X"B4",X"32",X"A8",X"33",X"2C",X"62",X"34",X"62",X"00",X"AA",X"2C",X"B4",X"2D",X"3C",
		X"63",X"77",X"0E",X"00",X"BC",X"2F",X"BC",X"31",X"77",X"0E",X"77",X"0E",X"31",X"B0",X"30",X"B2",
		X"2C",X"4F",X"0E",X"4F",X"0E",X"00",X"BA",X"38",X"B0",X"34",X"4F",X"0E",X"4F",X"0E",X"00",X"B6",
		X"37",X"BA",X"35",X"3C",X"60",X"3C",X"62",X"00",X"70",X"0E",X"70",X"0E",X"44",X"62",X"4F",X"5C",
		X"00",X"70",X"0E",X"70",X"0E",X"44",X"61",X"47",X"0E",X"03",X"B8",X"0E",X"B8",X"0E",X"47",X"0E",
		X"47",X"0E",X"61",X"B8",X"0E",X"B8",X"0E",X"47",X"0E",X"47",X"0E",X"61",X"B8",X"0E",X"B8",X"0E",
		X"47",X"0E",X"47",X"0E",X"02",X"B8",X"0E",X"B8",X"0E",X"47",X"0E",X"47",X"0E",X"61",X"B8",X"0E",
		X"B8",X"0E",X"47",X"0E",X"47",X"0E",X"02",X"B8",X"0E",X"B8",X"0E",X"47",X"0E",X"47",X"0E",X"61",
		X"B8",X"0E",X"B8",X"0E",X"47",X"0E",X"47",X"0E",X"02",X"B8",X"0E",X"B8",X"0E",X"47",X"0E",X"47",
		X"0E",X"61",X"B8",X"0E",X"B8",X"0E",X"47",X"0E",X"47",X"0E",X"02",X"B8",X"0E",X"B8",X"0E",X"47",
		X"0E",X"47",X"0E",X"61",X"70",X"0E",X"70",X"0E",X"36",X"5D",X"34",X"60",X"03",X"70",X"0E",X"9C",
		X"2C",X"2C",X"61",X"28",X"10",X"00",X"A4",X"2D",X"AC",X"2F",X"00",X"00",X"B4",X"2C",X"B4",X"33",
		X"28",X"10",X"2C",X"62",X"00",X"AC",X"30",X"A0",X"34",X"34",X"62",X"3C",X"63",X"00",X"A8",X"36",
		X"A8",X"36",X"44",X"62",X"4C",X"63",X"03",X"AC",X"2C",X"AE",X"37",X"54",X"62",X"57",X"3A",X"00",
		X"B2",X"38",X"B4",X"2C",X"57",X"3A",X"57",X"3A",X"49",X"BC",X"2D",X"C4",X"2F",X"57",X"3A",X"57",
		X"3A",X"59",X"C4",X"31",X"B8",X"34",X"57",X"3A",X"5F",X"5C",X"00",X"C4",X"2C",X"CC",X"2D",X"54",
		X"61",X"4C",X"60",X"00",X"D0",X"36",X"D0",X"36",X"4C",X"62",X"54",X"62",X"02",X"D0",X"36",X"D0",
		X"36",X"57",X"3A",X"57",X"3A",X"69",X"D0",X"36",X"D0",X"36",X"57",X"3A",X"57",X"3A",X"69",X"D0",
		X"36",X"CC",X"31",X"57",X"3A",X"57",X"3A",X"61",X"C4",X"30",X"BC",X"33",X"54",X"61",X"4C",X"60",
		X"00",X"B0",X"31",X"B2",X"2C",X"44",X"60",X"3C",X"61",X"00",X"BC",X"2D",X"C4",X"2F",X"34",X"60",
		X"2C",X"61",X"00",X"FF",X"C4",X"31",X"BC",X"30",X"00",X"00",X"B4",X"33",X"AC",X"32",X"00",X"00",
		X"A4",X"33",X"9C",X"31",X"00",X"00",X"94",X"31",X"8C",X"30",X"00",X"00",X"84",X"32",X"7C",X"30",
		X"00",X"00",X"74",X"33",X"6C",X"31",X"00",X"00",X"60",X"34",X"6C",X"2C",X"00",X"00",X"6C",X"30",
		X"64",X"32",X"00",X"00",X"5C",X"33",X"54",X"31",X"00",X"00",X"4C",X"30",X"40",X"34",X"00",X"00",
		X"4C",X"2D",X"54",X"2C",X"00",X"00",X"58",X"36",X"58",X"36",X"00",X"01",X"5C",X"2F",X"62",X"38",
		X"00",X"00",X"60",X"36",X"60",X"36",X"00",X"03",X"62",X"38",X"64",X"2E",X"00",X"00",X"68",X"36",
		X"68",X"36",X"00",X"02",X"6A",X"38",X"64",X"31",X"00",X"00",X"5C",X"30",X"50",X"32",X"00",X"00",
		X"52",X"2E",X"5C",X"2C",X"00",X"00",X"64",X"2D",X"6C",X"2C",X"00",X"00",X"74",X"2E",X"7C",X"2F",
		X"00",X"00",X"84",X"2D",X"8C",X"2F",X"00",X"00",X"90",X"36",X"90",X"36",X"00",X"01",X"90",X"36",
		X"90",X"36",X"00",X"01",X"90",X"36",X"90",X"36",X"00",X"03",X"88",X"34",X"92",X"36",X"00",X"00",
		X"90",X"36",X"90",X"36",X"00",X"02",X"90",X"36",X"90",X"36",X"00",X"01",X"90",X"36",X"90",X"36",
		X"00",X"01",X"94",X"2E",X"9C",X"2C",X"00",X"00",X"A4",X"2F",X"AC",X"2D",X"00",X"00",X"B4",X"2C",
		X"BC",X"2E",X"00",X"00",X"C4",X"2F",X"CC",X"2E",X"00",X"00",X"D0",X"36",X"D0",X"36",X"00",X"03",
		X"D0",X"36",X"D0",X"36",X"00",X"01",X"D0",X"36",X"D0",X"36",X"00",X"03",X"D0",X"36",X"CC",X"31",
		X"00",X"00",X"FF",X"CC",X"2E",X"D4",X"2D",X"00",X"00",X"D8",X"36",X"D8",X"36",X"00",X"03",X"DC",
		X"2F",X"D8",X"34",X"00",X"00",X"50",X"0E",X"40",X"0E",X"00",X"00",X"60",X"0E",X"60",X"0E",X"00",
		X"00",X"E0",X"36",X"E0",X"36",X"00",X"00",X"DC",X"31",X"D4",X"33",X"00",X"00",X"CC",X"30",X"C4",
		X"33",X"00",X"00",X"BC",X"31",X"B4",X"30",X"00",X"00",X"AC",X"30",X"A0",X"32",X"00",X"00",X"A2",
		X"2F",X"AC",X"2C",X"00",X"00",X"B0",X"36",X"B0",X"36",X"00",X"01",X"B0",X"36",X"B0",X"36",X"00",
		X"02",X"B4",X"2F",X"BC",X"2E",X"00",X"00",X"C0",X"36",X"C0",X"36",X"00",X"01",X"C0",X"36",X"C0",
		X"36",X"00",X"02",X"BC",X"30",X"B4",X"33",X"00",X"00",X"AC",X"31",X"A4",X"32",X"00",X"00",X"9C",
		X"31",X"94",X"30",X"00",X"00",X"88",X"34",X"92",X"38",X"00",X"00",X"90",X"36",X"90",X"36",X"00",
		X"00",X"8E",X"37",X"8C",X"30",X"00",X"00",X"88",X"36",X"88",X"36",X"00",X"01",X"88",X"36",X"88",
		X"36",X"00",X"02",X"84",X"32",X"78",X"31",X"00",X"00",X"7A",X"2D",X"84",X"2E",X"00",X"00",X"88",
		X"36",X"88",X"36",X"00",X"01",X"88",X"36",X"88",X"36",X"00",X"01",X"86",X"37",X"8A",X"35",X"00",
		X"00",X"80",X"34",X"8A",X"35",X"00",X"00",X"88",X"36",X"88",X"36",X"00",X"03",X"88",X"36",X"88",
		X"36",X"00",X"03",X"8C",X"2C",X"94",X"2D",X"00",X"00",X"9C",X"2D",X"A4",X"2C",X"00",X"00",X"AC",
		X"2C",X"B4",X"2F",X"00",X"00",X"B8",X"36",X"B8",X"36",X"00",X"03",X"B8",X"36",X"B8",X"36",X"00",
		X"02",X"BC",X"2D",X"C4",X"2C",X"00",X"00",X"CA",X"35",X"C0",X"34",X"00",X"00",X"FF",X"C4",X"31",
		X"BC",X"32",X"00",X"00",X"B4",X"30",X"AC",X"33",X"00",X"00",X"A4",X"31",X"9C",X"30",X"00",X"00",
		X"90",X"30",X"92",X"2E",X"00",X"00",X"98",X"36",X"98",X"36",X"00",X"01",X"98",X"36",X"98",X"36",
		X"00",X"01",X"98",X"36",X"98",X"36",X"00",X"01",X"98",X"36",X"98",X"36",X"00",X"02",X"9C",X"2C",
		X"A4",X"2E",X"00",X"00",X"A8",X"36",X"A8",X"36",X"00",X"03",X"A8",X"36",X"A8",X"36",X"00",X"03",
		X"A8",X"36",X"A8",X"36",X"00",X"03",X"A8",X"36",X"A8",X"36",X"00",X"02",X"A4",X"31",X"9C",X"33",
		X"00",X"00",X"94",X"30",X"8C",X"33",X"00",X"00",X"84",X"30",X"7C",X"31",X"00",X"00",X"74",X"33",
		X"6C",X"30",X"00",X"00",X"64",X"33",X"5C",X"31",X"00",X"00",X"54",X"30",X"4E",X"37",X"00",X"00",
		X"54",X"2E",X"5C",X"2D",X"00",X"00",X"60",X"36",X"60",X"36",X"00",X"03",X"60",X"36",X"60",X"36",
		X"00",X"01",X"60",X"36",X"60",X"36",X"00",X"01",X"5E",X"37",X"5C",X"31",X"00",X"00",X"50",X"34",
		X"5C",X"2F",X"00",X"00",X"60",X"36",X"60",X"36",X"00",X"02",X"60",X"36",X"60",X"36",X"00",X"03",
		X"60",X"36",X"60",X"36",X"00",X"01",X"60",X"36",X"60",X"36",X"00",X"01",X"58",X"34",X"64",X"2C",
		X"00",X"00",X"6C",X"2D",X"74",X"2F",X"00",X"00",X"7C",X"2C",X"84",X"2D",X"00",X"00",X"8C",X"2F",
		X"94",X"2C",X"00",X"00",X"9C",X"2D",X"A4",X"2F",X"00",X"00",X"A8",X"36",X"A8",X"36",X"00",X"01",
		X"AC",X"2E",X"B4",X"2F",X"00",X"00",X"BC",X"2C",X"C4",X"2D",X"00",X"00",X"FF",X"C4",X"31",X"BC",
		X"33",X"00",X"00",X"B0",X"34",X"BC",X"2C",X"00",X"00",X"C4",X"2D",X"C8",X"36",X"00",X"00",X"C8",
		X"36",X"C8",X"36",X"00",X"01",X"C8",X"36",X"CC",X"2E",X"00",X"00",X"D0",X"36",X"D0",X"36",X"00",
		X"01",X"D0",X"36",X"D0",X"36",X"00",X"02",X"CC",X"30",X"C4",X"31",X"00",X"00",X"BC",X"33",X"B4",
		X"31",X"00",X"00",X"AC",X"30",X"A4",X"31",X"00",X"00",X"9C",X"32",X"94",X"33",X"00",X"00",X"8C",
		X"31",X"84",X"30",X"00",X"00",X"7E",X"37",X"82",X"38",X"00",X"00",X"78",X"34",X"7E",X"37",X"00",
		X"00",X"82",X"35",X"84",X"2E",X"00",X"00",X"88",X"36",X"88",X"36",X"00",X"03",X"88",X"36",X"88",
		X"36",X"00",X"01",X"8C",X"2F",X"88",X"34",X"00",X"00",X"90",X"36",X"90",X"36",X"00",X"03",X"8C",
		X"30",X"84",X"31",X"00",X"00",X"7C",X"33",X"74",X"32",X"00",X"00",X"68",X"34",X"74",X"2D",X"00",
		X"00",X"7C",X"2F",X"84",X"2C",X"00",X"00",X"8C",X"2D",X"92",X"38",X"00",X"00",X"90",X"36",X"90",
		X"36",X"00",X"01",X"88",X"34",X"90",X"36",X"00",X"00",X"90",X"36",X"90",X"36",X"00",X"02",X"90",
		X"36",X"8C",X"31",X"00",X"00",X"80",X"33",X"82",X"2F",X"00",X"00",X"8C",X"2D",X"8E",X"37",X"00",
		X"00",X"90",X"36",X"90",X"36",X"00",X"01",X"90",X"36",X"90",X"36",X"00",X"02",X"90",X"36",X"90",
		X"36",X"00",X"03",X"94",X"2D",X"9C",X"2E",X"00",X"00",X"9E",X"37",X"A4",X"2E",X"00",X"00",X"AC",
		X"2F",X"B4",X"2D",X"00",X"00",X"BC",X"2C",X"C4",X"2C",X"00",X"00",X"FF",X"C0",X"34",X"C0",X"34",
		X"00",X"00",X"C4",X"30",X"BC",X"32",X"00",X"00",X"B6",X"37",X"BA",X"35",X"00",X"00",X"BA",X"38",
		X"BA",X"38",X"00",X"00",X"BC",X"2C",X"C4",X"2D",X"00",X"00",X"CC",X"2E",X"D4",X"2C",X"00",X"00",
		X"DC",X"2F",X"E0",X"36",X"00",X"00",X"E0",X"36",X"E0",X"36",X"00",X"01",X"E0",X"36",X"E0",X"36",
		X"00",X"02",X"E0",X"36",X"E2",X"35",X"00",X"00",X"E0",X"36",X"E0",X"36",X"00",X"01",X"D8",X"34",
		X"DC",X"31",X"00",X"00",X"D0",X"34",X"DC",X"2F",X"00",X"00",X"E0",X"36",X"E0",X"36",X"00",X"03",
		X"E0",X"36",X"E0",X"36",X"00",X"02",X"E0",X"36",X"DC",X"33",X"00",X"00",X"D4",X"31",X"CE",X"37",
		X"00",X"00",X"D2",X"38",X"C8",X"34",X"00",X"00",X"D0",X"36",X"D0",X"36",X"00",X"02",X"D0",X"36",
		X"D0",X"36",X"00",X"01",X"CC",X"31",X"C4",X"30",X"00",X"00",X"BC",X"33",X"B6",X"37",X"00",X"00",
		X"B8",X"38",X"B8",X"36",X"00",X"00",X"B8",X"36",X"B8",X"38",X"00",X"00",X"BC",X"2C",X"C4",X"2F",
		X"00",X"00",X"FF",X"CC",X"2C",X"D0",X"36",X"00",X"00",X"D0",X"36",X"D0",X"36",X"00",X"03",X"D4",
		X"2C",X"DC",X"2D",X"00",X"00",X"E0",X"36",X"E0",X"36",X"00",X"01",X"E0",X"36",X"E0",X"36",X"00",
		X"02",X"E0",X"36",X"E0",X"36",X"00",X"01",X"E0",X"36",X"E0",X"36",X"00",X"02",X"DC",X"30",X"D4",
		X"31",X"00",X"00",X"CC",X"33",X"C4",X"30",X"00",X"00",X"B8",X"34",X"BE",X"37",X"00",X"00",X"BE",
		X"37",X"C2",X"35",X"00",X"00",X"C3",X"2E",X"C3",X"31",X"00",X"00",X"B8",X"34",X"C4",X"2C",X"00",
		X"00",X"CC",X"2D",X"D0",X"36",X"00",X"00",X"D0",X"36",X"D0",X"36",X"00",X"03",X"D0",X"36",X"D0",
		X"36",X"00",X"02",X"CC",X"30",X"C8",X"36",X"00",X"00",X"C8",X"36",X"C8",X"36",X"00",X"01",X"C8",
		X"36",X"C8",X"36",X"00",X"03",X"C0",X"34",X"C8",X"36",X"00",X"00",X"C8",X"36",X"C8",X"36",X"00",
		X"02",X"C8",X"36",X"C8",X"36",X"00",X"01",X"C4",X"30",X"BC",X"31",X"00",X"00",X"B7",X"37",X"B7",
		X"37",X"00",X"00",X"BC",X"2F",X"C4",X"2E",X"00",X"00",X"FF",X"C6",X"37",X"C6",X"37",X"00",X"00",
		X"CA",X"35",X"C0",X"34",X"00",X"00",X"C8",X"36",X"C8",X"36",X"00",X"01",X"C8",X"36",X"C8",X"36",
		X"00",X"01",X"C8",X"36",X"CC",X"2C",X"00",X"00",X"D4",X"2D",X"D8",X"36",X"00",X"00",X"D8",X"36",
		X"D8",X"36",X"00",X"01",X"D8",X"36",X"D8",X"36",X"00",X"02",X"D8",X"36",X"D8",X"36",X"00",X"02",
		X"D4",X"33",X"CC",X"31",X"00",X"00",X"C4",X"33",X"B8",X"31",X"00",X"00",X"BA",X"2E",X"C4",X"2F",
		X"00",X"00",X"CC",X"2D",X"C8",X"34",X"00",X"00",X"D0",X"36",X"D0",X"36",X"00",X"02",X"D0",X"36",
		X"D0",X"36",X"00",X"03",X"D0",X"36",X"D0",X"36",X"00",X"02",X"CC",X"31",X"C0",X"34",X"00",X"00",
		X"C8",X"36",X"C8",X"36",X"00",X"03",X"C8",X"36",X"C8",X"36",X"00",X"01",X"C8",X"36",X"C8",X"36",
		X"00",X"01",X"C8",X"36",X"C8",X"36",X"00",X"01",X"CC",X"2C",X"D4",X"2D",X"00",X"00",X"D8",X"36",
		X"D8",X"36",X"00",X"02",X"D4",X"33",X"CC",X"31",X"00",X"00",X"C0",X"30",X"C2",X"2D",X"00",X"00",
		X"FF",X"CC",X"2C",X"D4",X"2D",X"00",X"00",X"D0",X"34",X"D0",X"34",X"00",X"00",X"D8",X"36",X"D8",
		X"36",X"00",X"03",X"D4",X"32",X"CC",X"31",X"00",X"00",X"C4",X"30",X"BC",X"33",X"00",X"00",X"B6",
		X"37",X"B7",X"37",X"00",X"00",X"BC",X"2C",X"C4",X"2D",X"00",X"00",X"CC",X"2F",X"D4",X"2E",X"00",
		X"00",X"D8",X"36",X"D8",X"36",X"00",X"01",X"D8",X"36",X"D8",X"36",X"00",X"01",X"D8",X"36",X"DC",
		X"2E",X"00",X"00",X"E0",X"36",X"E0",X"36",X"00",X"02",X"E0",X"36",X"E0",X"36",X"00",X"02",X"DC",
		X"30",X"D4",X"33",X"00",X"00",X"C8",X"34",X"D0",X"35",X"00",X"00",X"D0",X"36",X"D0",X"36",X"00",
		X"03",X"D0",X"36",X"D0",X"36",X"00",X"01",X"CC",X"31",X"C4",X"30",X"00",X"00",X"B8",X"33",X"BA",
		X"2E",X"00",X"00",X"C4",X"2F",X"CC",X"2C",X"00",X"00",X"D0",X"36",X"D0",X"36",X"00",X"01",X"D0",
		X"36",X"D0",X"36",X"00",X"02",X"D0",X"36",X"CC",X"30",X"00",X"00",X"C0",X"34",X"C8",X"36",X"00",
		X"00",X"C8",X"36",X"C8",X"36",X"00",X"02",X"FF",X"CC",X"2E",X"D4",X"2D",X"00",X"00",X"D8",X"36",
		X"D8",X"36",X"00",X"00",X"DC",X"2C",X"E4",X"2C",X"00",X"00",X"E6",X"37",X"E0",X"34",X"00",X"00",
		X"E4",X"33",X"DC",X"30",X"00",X"00",X"D0",X"34",X"DC",X"2F",X"00",X"00",X"E0",X"36",X"E0",X"36",
		X"00",X"02",X"E0",X"36",X"E0",X"36",X"00",X"03",X"E0",X"36",X"E0",X"36",X"00",X"02",X"DC",X"30",
		X"D4",X"33",X"00",X"00",X"CC",X"31",X"C4",X"33",X"00",X"00",X"B8",X"34",X"C0",X"36",X"00",X"00",
		X"C4",X"2E",X"C8",X"36",X"00",X"00",X"C8",X"36",X"C8",X"36",X"00",X"01",X"C8",X"36",X"C8",X"36",
		X"00",X"02",X"C8",X"36",X"C4",X"33",X"00",X"00",X"B8",X"30",X"BA",X"2D",X"00",X"00",X"C4",X"2C",
		X"CC",X"2F",X"00",X"00",X"D4",X"2E",X"DC",X"2D",X"00",X"00",X"E0",X"36",X"E0",X"36",X"00",X"01",
		X"E0",X"36",X"E0",X"36",X"00",X"03",X"D8",X"34",X"E2",X"35",X"00",X"00",X"E0",X"36",X"E0",X"36",
		X"00",X"02",X"DC",X"31",X"D0",X"34",X"00",X"00",X"D4",X"33",X"CC",X"30",X"00",X"00",X"FF",X"C4",
		X"33",X"B8",X"34",X"00",X"00",X"C4",X"2C",X"C8",X"36",X"00",X"00",X"C8",X"36",X"C8",X"36",X"00",
		X"03",X"C8",X"36",X"C8",X"36",X"00",X"01",X"C8",X"36",X"CC",X"2D",X"00",X"00",X"D4",X"2E",X"DC",
		X"2C",X"00",X"00",X"E0",X"36",X"E0",X"36",X"00",X"01",X"E0",X"36",X"E0",X"36",X"00",X"01",X"E0",
		X"36",X"E0",X"36",X"00",X"01",X"E0",X"36",X"E0",X"36",X"00",X"02",X"DC",X"32",X"D0",X"31",X"00",
		X"00",X"D2",X"2F",X"D0",X"34",X"00",X"00",X"DC",X"2D",X"E0",X"36",X"00",X"00",X"E0",X"36",X"E0",
		X"36",X"00",X"03",X"E0",X"36",X"E0",X"36",X"00",X"02",X"E0",X"36",X"DC",X"33",X"00",X"00",X"D4",
		X"31",X"CC",X"33",X"00",X"00",X"C0",X"33",X"C2",X"2E",X"00",X"00",X"C8",X"36",X"C8",X"36",X"00",
		X"01",X"C8",X"36",X"C8",X"36",X"00",X"02",X"C4",X"30",X"BC",X"31",X"00",X"00",X"B8",X"38",X"B8",
		X"38",X"00",X"00",X"BC",X"2E",X"C4",X"2D",X"00",X"00",X"CC",X"2F",X"D2",X"35",X"00",X"00",X"CE",
		X"37",X"CC",X"30",X"00",X"00",X"FF",X"C4",X"30",X"BC",X"31",X"00",X"00",X"B4",X"33",X"AC",X"30",
		X"00",X"00",X"A4",X"30",X"9C",X"31",X"00",X"00",X"94",X"33",X"8E",X"37",X"00",X"00",X"88",X"34",
		X"94",X"2E",X"00",X"00",X"98",X"36",X"98",X"36",X"00",X"01",X"9C",X"2F",X"A4",X"2C",X"00",X"00",
		X"A9",X"36",X"A9",X"36",X"00",X"03",X"A9",X"36",X"A9",X"36",X"00",X"02",X"AC",X"2E",X"B4",X"2D",
		X"00",X"00",X"BC",X"2C",X"C4",X"2C",X"00",X"00",X"C9",X"36",X"C9",X"36",X"00",X"01",X"C9",X"36",
		X"C9",X"36",X"00",X"02",X"C0",X"34",X"C0",X"34",X"00",X"00",X"CC",X"2F",X"CC",X"33",X"00",X"00",
		X"C8",X"36",X"C8",X"36",X"00",X"01",X"C4",X"33",X"BC",X"30",X"00",X"00",X"B0",X"34",X"B6",X"37",
		X"00",X"00",X"BC",X"2E",X"C4",X"2F",X"00",X"00",X"C8",X"36",X"C8",X"36",X"00",X"03",X"C4",X"33",
		X"BC",X"32",X"00",X"00",X"B4",X"30",X"AC",X"30",X"00",X"00",X"A4",X"31",X"9C",X"33",X"00",X"00",
		X"90",X"34",X"9C",X"2D",X"00",X"00",X"A4",X"2F",X"A8",X"36",X"00",X"00",X"A8",X"36",X"A8",X"36",
		X"00",X"01",X"A8",X"36",X"A8",X"36",X"00",X"01",X"AC",X"2C",X"B4",X"2E",X"00",X"00",X"BA",X"2D",
		X"C4",X"2C",X"00",X"00",X"FF",X"C4",X"37",X"C4",X"31",X"00",X"00",X"BC",X"30",X"B4",X"30",X"00",
		X"00",X"AC",X"31",X"A4",X"31",X"00",X"00",X"9C",X"30",X"94",X"30",X"28",X"63",X"34",X"63",X"00",
		X"8C",X"32",X"84",X"30",X"37",X"5E",X"37",X"5E",X"00",X"7C",X"30",X"74",X"33",X"37",X"5E",X"3C",
		X"62",X"00",X"6C",X"33",X"66",X"37",X"3F",X"5E",X"3F",X"5E",X"00",X"6C",X"2C",X"74",X"2D",X"3F",
		X"5E",X"44",X"63",X"00",X"7C",X"2F",X"84",X"2F",X"4C",X"63",X"54",X"62",X"00",X"8C",X"2C",X"8E",
		X"37",X"5A",X"5F",X"5C",X"62",X"00",X"90",X"36",X"90",X"36",X"64",X"62",X"6A",X"5F",X"01",X"90",
		X"36",X"90",X"36",X"6A",X"5F",X"6A",X"5F",X"01",X"90",X"36",X"90",X"36",X"64",X"61",X"5C",X"61",
		X"03",X"90",X"36",X"90",X"36",X"57",X"5E",X"57",X"5E",X"02",X"8C",X"30",X"88",X"38",X"57",X"5E",
		X"57",X"5E",X"00",X"80",X"34",X"8C",X"2F",X"54",X"61",X"4C",X"61",X"00",X"90",X"36",X"90",X"36",
		X"47",X"5E",X"47",X"5E",X"01",X"94",X"2C",X"9C",X"2C",X"47",X"5E",X"47",X"5E",X"00",X"A4",X"2F",
		X"AC",X"2D",X"47",X"5E",X"44",X"61",X"00",X"B0",X"36",X"B0",X"36",X"3C",X"61",X"3C",X"62",X"01",
		X"B0",X"2F",X"B8",X"35",X"44",X"63",X"4C",X"62",X"00",X"BC",X"2F",X"C4",X"2F",X"4F",X"5E",X"4F",
		X"5E",X"00",X"CC",X"2C",X"C8",X"34",X"54",X"63",X"5C",X"63",X"00",X"D0",X"36",X"D0",X"36",X"64",
		X"62",X"6C",X"62",X"01",X"D0",X"36",X"D0",X"36",X"6F",X"5E",X"6F",X"5E",X"02",X"D4",X"2C",X"DC",
		X"2D",X"6F",X"5E",X"6F",X"5E",X"00",X"E4",X"2F",X"E8",X"36",X"6F",X"5E",X"6C",X"60",X"00",X"E8",
		X"36",X"E8",X"36",X"64",X"60",X"5C",X"61",X"03",X"E8",X"36",X"E4",X"31",X"54",X"60",X"4C",X"61",
		X"00",X"DC",X"30",X"D4",X"31",X"44",X"60",X"3C",X"61",X"00",X"D0",X"36",X"D0",X"36",X"3C",X"62",
		X"44",X"62",X"01",X"D0",X"36",X"D0",X"36",X"4C",X"63",X"54",X"63",X"01",X"D0",X"36",X"D0",X"36",
		X"5C",X"62",X"64",X"63",X"02",X"D0",X"36",X"D0",X"36",X"6C",X"62",X"74",X"63",X"03",X"CC",X"30",
		X"C4",X"33",X"74",X"60",X"6C",X"60",X"00",X"BC",X"31",X"B4",X"31",X"64",X"60",X"5C",X"61",X"00",
		X"AC",X"30",X"AC",X"2D",X"54",X"61",X"4C",X"60",X"00",X"B4",X"2C",X"BC",X"2C",X"44",X"61",X"3C",
		X"60",X"00",X"C4",X"2F",X"C4",X"37",X"34",X"60",X"2C",X"60",X"00",X"FF",X"C4",X"30",X"B8",X"34",
		X"2C",X"62",X"37",X"5C",X"00",X"C4",X"2D",X"C0",X"34",X"34",X"63",X"3E",X"62",X"00",X"C8",X"36",
		X"C8",X"36",X"44",X"62",X"4C",X"63",X"02",X"C8",X"36",X"C8",X"36",X"54",X"62",X"5C",X"63",X"01",
		X"C8",X"36",X"C8",X"36",X"64",X"62",X"6C",X"63",X"01",X"C4",X"30",X"BC",X"30",X"74",X"62",X"7A",
		X"5F",X"00",X"B4",X"33",X"AC",X"31",X"7A",X"5F",X"7A",X"5F",X"00",X"A4",X"31",X"98",X"34",X"7C",
		X"62",X"7F",X"5E",X"00",X"A4",X"2C",X"AC",X"2F",X"87",X"5C",X"7F",X"5E",X"00",X"B0",X"36",X"B0",
		X"36",X"7F",X"5D",X"80",X"5C",X"03",X"B0",X"36",X"B0",X"36",X"80",X"5F",X"80",X"5F",X"03",X"B0",
		X"36",X"B0",X"36",X"80",X"5F",X"7C",X"60",X"02",X"B0",X"36",X"B0",X"36",X"74",X"60",X"6C",X"61",
		X"01",X"B0",X"36",X"B0",X"36",X"64",X"60",X"5C",X"60",X"01",X"B0",X"36",X"B0",X"36",X"54",X"61",
		X"4C",X"61",X"01",X"B4",X"2C",X"BC",X"2C",X"44",X"61",X"3C",X"61",X"00",X"C4",X"2F",X"C4",X"37",
		X"34",X"61",X"2C",X"61",X"00",X"C4",X"37",X"C4",X"33",X"2C",X"63",X"34",X"63",X"00",X"BC",X"30",
		X"B4",X"32",X"3C",X"63",X"40",X"5F",X"00",X"AC",X"30",X"A4",X"31",X"40",X"5F",X"40",X"5F",X"00",
		X"9C",X"30",X"94",X"30",X"40",X"5F",X"39",X"5D",X"00",X"94",X"2C",X"94",X"37",X"40",X"5C",X"3F",
		X"5D",X"00",X"9C",X"2D",X"A4",X"2F",X"40",X"5C",X"40",X"5F",X"00",X"AC",X"36",X"AC",X"2D",X"44",
		X"62",X"4C",X"63",X"00",X"B4",X"2F",X"BC",X"2C",X"54",X"63",X"5C",X"62",X"00",X"C4",X"2D",X"CC",
		X"2F",X"64",X"62",X"6C",X"62",X"00",X"D0",X"36",X"D0",X"36",X"6F",X"5D",X"6F",X"5D",X"01",X"D0",
		X"36",X"D0",X"36",X"70",X"5C",X"6F",X"5D",X"01",X"D0",X"36",X"D0",X"36",X"70",X"5C",X"6F",X"5D",
		X"01",X"D0",X"36",X"D0",X"36",X"6C",X"60",X"64",X"60",X"03",X"D0",X"36",X"D0",X"36",X"5C",X"61",
		X"54",X"60",X"02",X"D0",X"36",X"D0",X"36",X"4C",X"60",X"44",X"60",X"02",X"D4",X"2D",X"DC",X"2F",
		X"40",X"5F",X"3F",X"5E",X"00",X"E0",X"36",X"E0",X"36",X"40",X"5C",X"40",X"5F",X"01",X"E0",X"36",
		X"E0",X"36",X"40",X"5C",X"3F",X"5D",X"01",X"E0",X"36",X"D8",X"30",X"3C",X"61",X"34",X"60",X"00",
		X"D4",X"33",X"CC",X"31",X"2C",X"61",X"2A",X"5F",X"00",X"FF",X"C4",X"33",X"BC",X"31",X"00",X"00",
		X"B4",X"33",X"AC",X"30",X"00",X"00",X"A4",X"30",X"A4",X"2F",X"00",X"00",X"AC",X"2C",X"AF",X"37",
		X"00",X"00",X"AF",X"37",X"B0",X"35",X"00",X"00",X"B4",X"2F",X"BC",X"2C",X"00",X"00",X"C0",X"36",
		X"C0",X"36",X"00",X"02",X"C0",X"36",X"C0",X"36",X"00",X"05",X"C0",X"36",X"C0",X"36",X"00",X"00",
		X"C0",X"36",X"C0",X"36",X"00",X"00",X"C4",X"2F",X"CC",X"2C",X"00",X"00",X"D4",X"2F",X"DC",X"2C",
		X"00",X"00",X"E0",X"35",X"E0",X"35",X"00",X"00",X"E0",X"36",X"E0",X"36",X"00",X"02",X"E0",X"36",
		X"E0",X"36",X"00",X"02",X"E0",X"36",X"E0",X"36",X"00",X"05",X"E0",X"36",X"E0",X"36",X"00",X"00",
		X"E0",X"36",X"E0",X"36",X"00",X"00",X"E0",X"36",X"E0",X"36",X"00",X"00",X"DC",X"33",X"D4",X"31",
		X"00",X"00",X"CC",X"31",X"C4",X"33",X"00",X"00",X"BC",X"32",X"B4",X"30",X"00",X"00",X"B0",X"36",
		X"B0",X"36",X"00",X"00",X"AC",X"33",X"A4",X"30",X"00",X"00",X"9C",X"30",X"94",X"31",X"00",X"00",
		X"8C",X"33",X"84",X"32",X"00",X"00",X"84",X"2F",X"8C",X"2C",X"00",X"00",X"90",X"36",X"90",X"36",
		X"00",X"00",X"94",X"2F",X"9C",X"2C",X"00",X"00",X"A0",X"36",X"A0",X"36",X"00",X"02",X"A0",X"36",
		X"A0",X"36",X"00",X"05",X"A0",X"36",X"A0",X"36",X"00",X"05",X"A0",X"36",X"A0",X"36",X"00",X"00",
		X"A0",X"36",X"A0",X"36",X"00",X"00",X"A0",X"36",X"A4",X"2D",X"00",X"00",X"AC",X"2D",X"B4",X"2F",
		X"00",X"00",X"BC",X"2C",X"C4",X"2C",X"00",X"00",X"FF",X"C4",X"33",X"BC",X"31",X"2C",X"62",X"34",
		X"63",X"00",X"B4",X"30",X"AC",X"32",X"3C",X"62",X"42",X"5C",X"00",X"A4",X"30",X"9C",X"30",X"3E",
		X"5D",X"44",X"62",X"00",X"94",X"33",X"88",X"32",X"4C",X"62",X"54",X"63",X"00",X"8A",X"2F",X"94",
		X"2D",X"5C",X"62",X"64",X"63",X"00",X"9C",X"2C",X"9E",X"37",X"6C",X"63",X"74",X"62",X"00",X"A0",
		X"36",X"A3",X"2D",X"7C",X"63",X"84",X"62",X"00",X"AA",X"36",X"AA",X"35",X"87",X"60",X"86",X"5F",
		X"00",X"AA",X"36",X"AA",X"36",X"87",X"63",X"84",X"61",X"02",X"A7",X"37",X"A5",X"34",X"7C",X"61",
		X"74",X"61",X"00",X"AC",X"2F",X"B4",X"2C",X"6C",X"60",X"64",X"60",X"00",X"B8",X"36",X"B8",X"36",
		X"5F",X"5D",X"64",X"5C",X"01",X"B8",X"36",X"B8",X"36",X"5F",X"5D",X"5C",X"61",X"01",X"B0",X"34",
		X"B0",X"34",X"54",X"60",X"4C",X"61",X"00",X"B8",X"36",X"B8",X"36",X"47",X"5E",X"47",X"5E",X"02",
		X"B4",X"31",X"AC",X"30",X"4A",X"5C",X"47",X"5E",X"00",X"A4",X"33",X"98",X"34",X"4A",X"5F",X"4A",
		X"5F",X"00",X"9E",X"37",X"9C",X"30",X"47",X"5D",X"4F",X"5C",X"00",X"94",X"31",X"8C",X"33",X"47",
		X"5E",X"47",X"3A",X"00",X"84",X"30",X"78",X"32",X"4F",X"5C",X"47",X"3A",X"00",X"7A",X"2C",X"84",
		X"2F",X"44",X"60",X"3C",X"61",X"00",X"88",X"36",X"88",X"38",X"34",X"60",X"2C",X"61",X"03",X"84",
		X"30",X"7C",X"31",X"2F",X"5C",X"2A",X"5F",X"00",X"74",X"33",X"6C",X"31",X"00",X"00",X"60",X"34",
		X"6C",X"2C",X"00",X"00",X"74",X"2D",X"76",X"37",X"00",X"00",X"78",X"36",X"78",X"36",X"00",X"01",
		X"78",X"36",X"78",X"36",X"00",X"01",X"78",X"36",X"78",X"36",X"00",X"03",X"74",X"33",X"6C",X"31",
		X"00",X"00",X"60",X"34",X"60",X"34",X"00",X"00",X"6C",X"2C",X"74",X"2D",X"00",X"00",X"7C",X"2D",
		X"84",X"2F",X"00",X"00",X"8C",X"2F",X"94",X"2C",X"00",X"00",X"9C",X"2D",X"A4",X"2F",X"00",X"00",
		X"AC",X"2C",X"B4",X"2F",X"00",X"00",X"BC",X"2C",X"C4",X"2D",X"00",X"00",X"FF",X"C0",X"31",X"B8",
		X"30",X"28",X"62",X"30",X"62",X"00",X"B0",X"32",X"B0",X"36",X"38",X"62",X"40",X"62",X"00",X"B0",
		X"2E",X"B8",X"2D",X"48",X"62",X"50",X"62",X"00",X"C0",X"2E",X"C8",X"2D",X"5F",X"62",X"5F",X"3A",
		X"00",X"D0",X"36",X"D0",X"36",X"5F",X"3A",X"5F",X"60",X"02",X"D0",X"36",X"D0",X"36",X"50",X"3A",
		X"50",X"3A",X"68",X"D0",X"36",X"D0",X"36",X"5F",X"62",X"5F",X"3A",X"02",X"D0",X"36",X"D0",X"36",
		X"5F",X"3A",X"5F",X"3A",X"61",X"D0",X"36",X"D0",X"2E",X"5F",X"3A",X"5F",X"3A",X"61",X"D8",X"36",
		X"D8",X"36",X"5F",X"3A",X"5F",X"60",X"03",X"D8",X"36",X"D8",X"36",X"50",X"60",X"48",X"60",X"03",
		X"D0",X"32",X"D0",X"36",X"40",X"60",X"38",X"60",X"00",X"D0",X"36",X"D0",X"36",X"30",X"3A",X"30",
		X"3A",X"89",X"C8",X"31",X"C0",X"32",X"30",X"3A",X"30",X"3A",X"79",X"C0",X"36",X"C0",X"36",X"30",
		X"3A",X"30",X"3A",X"79",X"B8",X"31",X"B0",X"32",X"30",X"3A",X"30",X"60",X"00",X"B0",X"36",X"B0",
		X"36",X"28",X"3A",X"28",X"3A",X"71",X"B0",X"36",X"B0",X"36",X"28",X"3A",X"28",X"3A",X"71",X"B0",
		X"2E",X"B8",X"2D",X"30",X"62",X"30",X"3A",X"00",X"C0",X"36",X"C0",X"2E",X"30",X"3A",X"30",X"3A",
		X"79",X"C8",X"36",X"C8",X"36",X"38",X"62",X"40",X"62",X"03",X"C8",X"36",X"C8",X"36",X"48",X"62",
		X"48",X"3A",X"02",X"C8",X"2E",X"D0",X"36",X"48",X"3A",X"50",X"62",X"00",X"D0",X"36",X"D0",X"36",
		X"5F",X"62",X"5F",X"3A",X"03",X"D0",X"36",X"D0",X"2D",X"5F",X"3A",X"5F",X"60",X"00",X"D8",X"36",
		X"D8",X"36",X"50",X"60",X"48",X"60",X"03",X"D8",X"36",X"D8",X"36",X"40",X"60",X"38",X"60",X"02",
		X"D0",X"31",X"C8",X"32",X"30",X"60",X"28",X"60",X"00",X"FF",X"60",X"0E",X"60",X"0E",X"47",X"0E",
		X"47",X"0E",X"02",X"60",X"0E",X"60",X"0E",X"47",X"0E",X"47",X"0E",X"02",X"60",X"0E",X"60",X"0E",
		X"37",X"0E",X"37",X"0E",X"00",X"60",X"0E",X"60",X"0E",X"37",X"0E",X"37",X"0E",X"00",X"60",X"0E",
		X"60",X"0E",X"37",X"0E",X"37",X"0E",X"00",X"50",X"0E",X"50",X"0E",X"37",X"0E",X"37",X"0E",X"02",
		X"50",X"0E",X"50",X"0E",X"37",X"0E",X"37",X"0E",X"00",X"60",X"0E",X"60",X"0E",X"37",X"0E",X"37",
		X"0E",X"00",X"60",X"0E",X"60",X"0E",X"37",X"0E",X"37",X"0E",X"00",X"60",X"0E",X"60",X"0E",X"37",
		X"0E",X"47",X"0E",X"00",X"60",X"0E",X"60",X"0E",X"47",X"0E",X"47",X"0E",X"00",X"60",X"0E",X"60",
		X"0E",X"47",X"0E",X"47",X"0E",X"00",X"60",X"0E",X"60",X"0E",X"47",X"0E",X"47",X"0E",X"02",X"60",
		X"0E",X"60",X"0E",X"47",X"0E",X"47",X"0E",X"02",X"60",X"0E",X"60",X"0E",X"47",X"0E",X"47",X"0E",
		X"02",X"60",X"0E",X"60",X"0E",X"2F",X"0E",X"2F",X"0E",X"02",X"60",X"0E",X"60",X"0E",X"2F",X"0E",
		X"2F",X"0E",X"00",X"60",X"0E",X"60",X"0E",X"2F",X"0E",X"2F",X"0E",X"00",X"40",X"0E",X"40",X"0E",
		X"2F",X"0E",X"2F",X"0E",X"00",X"40",X"0E",X"40",X"0E",X"2F",X"0E",X"2F",X"0E",X"00",X"40",X"0E",
		X"40",X"0E",X"2F",X"0E",X"2F",X"0E",X"00",X"40",X"0E",X"40",X"0E",X"2F",X"0E",X"2F",X"0E",X"00",
		X"40",X"0E",X"40",X"0E",X"2F",X"0E",X"2F",X"0E",X"00",X"A0",X"0E",X"A0",X"0E",X"2F",X"0E",X"2F",
		X"0E",X"01",X"A0",X"0E",X"A0",X"0E",X"2F",X"0E",X"2F",X"0E",X"01",X"A0",X"0E",X"A0",X"0E",X"2F",
		X"0E",X"2F",X"0E",X"03",X"A0",X"0E",X"A0",X"0E",X"2F",X"0E",X"2F",X"0E",X"00",X"A0",X"0E",X"A0",
		X"0E",X"2F",X"0E",X"2F",X"0E",X"00",X"A0",X"0E",X"A0",X"0E",X"2F",X"0E",X"2F",X"0E",X"02",X"A0",
		X"0E",X"A0",X"0E",X"37",X"0E",X"37",X"0E",X"02",X"A0",X"0E",X"A0",X"0E",X"8F",X"0E",X"8F",X"0E",
		X"02",X"A0",X"0E",X"A0",X"0E",X"8F",X"0E",X"8F",X"0E",X"02",X"A0",X"0E",X"A0",X"0E",X"8F",X"0E",
		X"8F",X"0E",X"02",X"A0",X"0E",X"A0",X"0E",X"8F",X"0E",X"8F",X"0E",X"00",X"A0",X"0E",X"A0",X"0E",
		X"8F",X"0E",X"8F",X"0E",X"00",X"FF",X"A0",X"0E",X"A0",X"0E",X"8F",X"0E",X"8F",X"0E",X"00",X"D8",
		X"0E",X"D8",X"0E",X"8F",X"0E",X"8F",X"0E",X"00",X"D8",X"0E",X"D8",X"0E",X"8F",X"0E",X"8F",X"0E",
		X"00",X"D8",X"0E",X"D8",X"0E",X"8F",X"0E",X"8F",X"0E",X"00",X"D8",X"0E",X"D8",X"0E",X"C7",X"0E",
		X"C7",X"0E",X"00",X"D8",X"0E",X"D8",X"0E",X"C7",X"0E",X"C7",X"0E",X"02",X"D8",X"0E",X"D8",X"0E",
		X"C7",X"0E",X"C7",X"0E",X"02",X"D8",X"0E",X"D8",X"0E",X"C7",X"0E",X"C7",X"0E",X"02",X"D8",X"0E",
		X"D8",X"0E",X"C7",X"0E",X"C7",X"0E",X"02",X"D8",X"0E",X"D8",X"0E",X"C7",X"0E",X"C7",X"0E",X"00",
		X"D8",X"0E",X"D8",X"0E",X"3F",X"0E",X"3F",X"0E",X"01",X"D8",X"0E",X"D8",X"0E",X"3F",X"0E",X"3F",
		X"0E",X"01",X"D8",X"0E",X"D8",X"0E",X"3F",X"0E",X"3F",X"0E",X"01",X"D8",X"0E",X"D8",X"0E",X"3F",
		X"0E",X"3F",X"0E",X"01",X"D8",X"0E",X"D8",X"0E",X"3F",X"0E",X"3F",X"0E",X"01",X"D8",X"0E",X"D8",
		X"0E",X"3F",X"0E",X"3F",X"0E",X"03",X"50",X"0E",X"50",X"0E",X"3F",X"0E",X"3F",X"0E",X"00",X"50",
		X"0E",X"50",X"0E",X"3F",X"0E",X"3F",X"0E",X"00",X"50",X"0E",X"50",X"0E",X"3F",X"0E",X"3F",X"0E",
		X"00",X"50",X"0E",X"50",X"0E",X"3F",X"0E",X"3F",X"0E",X"00",X"50",X"0E",X"50",X"0E",X"3F",X"0E",
		X"3F",X"0E",X"00",X"D8",X"0E",X"D8",X"0E",X"3F",X"0E",X"3F",X"0E",X"01",X"D8",X"0E",X"D8",X"0E",
		X"3F",X"0E",X"3F",X"0E",X"00",X"D8",X"0E",X"D8",X"0E",X"3F",X"0E",X"3F",X"0E",X"00",X"D8",X"0E",
		X"D8",X"0E",X"3F",X"0E",X"3F",X"0E",X"01",X"D8",X"0E",X"D8",X"0E",X"3F",X"0E",X"3F",X"0E",X"01",
		X"D8",X"0E",X"D8",X"0E",X"3F",X"0E",X"3F",X"0E",X"00",X"D8",X"0E",X"D8",X"0E",X"3F",X"0E",X"3F",
		X"0E",X"00",X"FF",X"C8",X"0E",X"C8",X"0E",X"AF",X"0E",X"AF",X"0E",X"00",X"E0",X"0E",X"E0",X"0E",
		X"AF",X"0E",X"AF",X"0E",X"00",X"E0",X"0E",X"E0",X"0E",X"AF",X"0E",X"AF",X"0E",X"00",X"E0",X"0E",
		X"E0",X"0E",X"B7",X"0E",X"CF",X"0E",X"00",X"E0",X"0E",X"E0",X"0E",X"CF",X"0E",X"C7",X"0E",X"00",
		X"E0",X"0E",X"E0",X"0E",X"BF",X"0E",X"BF",X"0E",X"00",X"E0",X"0E",X"E0",X"0E",X"BF",X"0E",X"BF",
		X"0E",X"00",X"D8",X"0E",X"D8",X"0E",X"4F",X"0E",X"4F",X"0E",X"01",X"D8",X"0E",X"D8",X"0E",X"4F",
		X"0E",X"4F",X"0E",X"01",X"D8",X"0E",X"D8",X"0E",X"4F",X"0E",X"4F",X"0E",X"01",X"D8",X"0E",X"D8",
		X"0E",X"4F",X"0E",X"4F",X"0E",X"01",X"D8",X"0E",X"D8",X"0E",X"4F",X"0E",X"4F",X"0E",X"03",X"60",
		X"0E",X"60",X"0E",X"4F",X"0E",X"4F",X"0E",X"00",X"60",X"0E",X"60",X"0E",X"4F",X"0E",X"4F",X"0E",
		X"00",X"60",X"0E",X"60",X"0E",X"4F",X"0E",X"37",X"0E",X"00",X"60",X"0E",X"60",X"0E",X"37",X"0E",
		X"37",X"0E",X"00",X"60",X"0E",X"60",X"0E",X"37",X"0E",X"37",X"0E",X"00",X"48",X"0E",X"48",X"0E",
		X"37",X"0E",X"37",X"0E",X"00",X"48",X"0E",X"48",X"0E",X"37",X"0E",X"37",X"0E",X"00",X"48",X"0E",
		X"48",X"0E",X"37",X"0E",X"37",X"0E",X"00",X"48",X"0E",X"58",X"0E",X"37",X"0E",X"37",X"0E",X"00",
		X"60",X"0E",X"60",X"0E",X"37",X"0E",X"37",X"0E",X"00",X"60",X"0E",X"60",X"0E",X"37",X"0E",X"37",
		X"0E",X"00",X"60",X"0E",X"60",X"0E",X"47",X"0E",X"47",X"0E",X"00",X"60",X"0E",X"60",X"0E",X"47",
		X"0E",X"4F",X"0E",X"00",X"60",X"0E",X"60",X"0E",X"4F",X"0E",X"4F",X"0E",X"00",X"60",X"0E",X"60",
		X"0E",X"4F",X"0E",X"4F",X"0E",X"00",X"60",X"0E",X"60",X"0E",X"4F",X"0E",X"4F",X"0E",X"00",X"60",
		X"0E",X"60",X"0E",X"4F",X"0E",X"4F",X"0E",X"00",X"60",X"0E",X"60",X"0E",X"4F",X"0E",X"4F",X"0E",
		X"00",X"FF",X"60",X"0E",X"60",X"0E",X"47",X"0E",X"47",X"0E",X"00",X"70",X"0E",X"70",X"0E",X"47",
		X"0E",X"47",X"0E",X"00",X"70",X"0E",X"70",X"0E",X"47",X"0E",X"47",X"0E",X"00",X"70",X"0E",X"70",
		X"0E",X"47",X"0E",X"47",X"0E",X"00",X"70",X"0E",X"70",X"0E",X"5F",X"0E",X"5F",X"0E",X"00",X"70",
		X"0E",X"70",X"0E",X"5F",X"0E",X"5F",X"0E",X"00",X"70",X"0E",X"70",X"0E",X"5F",X"0E",X"5F",X"0E",
		X"00",X"70",X"0E",X"70",X"0E",X"57",X"0E",X"57",X"0E",X"00",X"70",X"0E",X"70",X"0E",X"57",X"0E",
		X"57",X"0E",X"00",X"70",X"0E",X"68",X"0E",X"57",X"0E",X"4F",X"0E",X"00",X"68",X"0E",X"68",X"0E",
		X"4F",X"0E",X"4F",X"0E",X"00",X"68",X"0E",X"68",X"0E",X"4F",X"0E",X"47",X"0E",X"00",X"68",X"0E",
		X"60",X"0E",X"47",X"0E",X"47",X"0E",X"00",X"60",X"0E",X"60",X"0E",X"47",X"0E",X"47",X"0E",X"00",
		X"58",X"0E",X"58",X"0E",X"47",X"0E",X"47",X"0E",X"00",X"58",X"0E",X"D8",X"0E",X"47",X"0E",X"47",
		X"0E",X"00",X"D8",X"0E",X"D8",X"0E",X"47",X"0E",X"47",X"0E",X"00",X"D8",X"0E",X"D8",X"0E",X"47",
		X"0E",X"47",X"0E",X"01",X"D8",X"0E",X"D8",X"0E",X"47",X"0E",X"47",X"0E",X"00",X"D8",X"0E",X"D8",
		X"0E",X"47",X"0E",X"47",X"0E",X"00",X"D8",X"0E",X"D8",X"0E",X"47",X"0E",X"47",X"0E",X"00",X"D8",
		X"0E",X"D8",X"0E",X"C7",X"0E",X"C7",X"0E",X"00",X"D8",X"0E",X"D8",X"0E",X"C7",X"0E",X"C7",X"0E",
		X"00",X"D8",X"0E",X"D8",X"0E",X"C7",X"0E",X"C7",X"0E",X"00",X"D8",X"0E",X"D8",X"0E",X"C7",X"0E",
		X"C7",X"0E",X"00",X"D8",X"0E",X"D8",X"0E",X"C7",X"0E",X"C7",X"0E",X"00",X"D8",X"0E",X"D8",X"0E",
		X"C7",X"0E",X"C7",X"0E",X"00",X"D8",X"0E",X"D8",X"0E",X"C7",X"0E",X"C7",X"0E",X"00",X"D8",X"0E",
		X"D8",X"0E",X"C7",X"0E",X"C7",X"0E",X"00",X"D8",X"0E",X"D8",X"0E",X"3F",X"0E",X"3F",X"0E",X"01",
		X"D8",X"0E",X"D8",X"0E",X"3F",X"0E",X"3F",X"0E",X"01",X"D8",X"0E",X"D8",X"0E",X"3F",X"0E",X"3F",
		X"0E",X"01",X"D8",X"0E",X"D8",X"0E",X"3F",X"0E",X"3F",X"0E",X"01",X"D8",X"0E",X"D8",X"0E",X"3F",
		X"0E",X"3F",X"0E",X"01",X"D8",X"0E",X"D8",X"0E",X"3F",X"0E",X"3F",X"0E",X"03",X"50",X"0E",X"50",
		X"0E",X"3F",X"0E",X"3F",X"0E",X"00",X"50",X"0E",X"50",X"0E",X"3F",X"0E",X"3F",X"0E",X"00",X"50",
		X"0E",X"50",X"0E",X"3F",X"0E",X"3F",X"0E",X"00",X"60",X"0E",X"60",X"0E",X"3F",X"0E",X"3F",X"0E",
		X"01",X"60",X"0E",X"60",X"0E",X"3F",X"0E",X"3F",X"0E",X"02",X"60",X"0E",X"60",X"0E",X"3F",X"0E",
		X"3F",X"0E",X"03",X"FF",X"C8",X"0E",X"C8",X"0E",X"00",X"00",X"80",X"0E",X"80",X"0E",X"00",X"01",
		X"80",X"0E",X"80",X"0E",X"00",X"01",X"80",X"0E",X"C8",X"0E",X"00",X"00",X"C8",X"0E",X"C8",X"0E",
		X"00",X"00",X"C8",X"0E",X"C8",X"0E",X"00",X"03",X"50",X"0E",X"50",X"0E",X"00",X"03",X"50",X"0E",
		X"50",X"0E",X"00",X"01",X"50",X"0E",X"50",X"0E",X"00",X"00",X"60",X"0E",X"60",X"0E",X"00",X"00",
		X"60",X"0E",X"60",X"0E",X"00",X"01",X"60",X"0E",X"60",X"0E",X"00",X"01",X"C8",X"0E",X"C8",X"0E",
		X"00",X"00",X"C8",X"0E",X"C8",X"0E",X"00",X"00",X"C8",X"0E",X"C8",X"0E",X"00",X"00",X"88",X"0E",
		X"88",X"0E",X"00",X"03",X"88",X"0E",X"88",X"0E",X"00",X"01",X"88",X"0E",X"78",X"0E",X"00",X"00",
		X"78",X"0E",X"78",X"0E",X"00",X"01",X"78",X"0E",X"C8",X"0E",X"00",X"00",X"C8",X"0E",X"C8",X"0E",
		X"00",X"00",X"48",X"0E",X"49",X"1F",X"00",X"00",X"49",X"23",X"49",X"11",X"00",X"00",X"49",X"1B",
		X"49",X"11",X"00",X"00",X"48",X"0E",X"C8",X"0E",X"00",X"00",X"C8",X"0E",X"C8",X"0E",X"00",X"00",
		X"C8",X"0E",X"C8",X"0E",X"00",X"00",X"C8",X"0E",X"C8",X"0E",X"00",X"03",X"C8",X"0E",X"C8",X"0E",
		X"00",X"00",X"C8",X"0E",X"C8",X"0E",X"00",X"01",X"C8",X"0E",X"C8",X"0E",X"00",X"02",X"C8",X"0E",
		X"C8",X"0E",X"00",X"00",X"80",X"0E",X"80",X"0E",X"00",X"03",X"80",X"0E",X"80",X"0E",X"00",X"00",
		X"C8",X"0E",X"C8",X"0E",X"00",X"00",X"FF",X"C8",X"0E",X"C8",X"0E",X"00",X"00",X"C8",X"0E",X"C8",
		X"0E",X"00",X"03",X"90",X"0E",X"90",X"0E",X"00",X"00",X"50",X"0E",X"50",X"0E",X"00",X"03",X"90",
		X"0E",X"90",X"0E",X"00",X"00",X"C8",X"0E",X"C8",X"0E",X"00",X"00",X"C8",X"0E",X"C8",X"0E",X"00",
		X"03",X"98",X"0E",X"98",X"0E",X"00",X"01",X"98",X"0E",X"98",X"0E",X"00",X"01",X"98",X"0E",X"98",
		X"0E",X"00",X"00",X"C8",X"0E",X"C8",X"0E",X"00",X"00",X"48",X"1B",X"48",X"1F",X"00",X"00",X"48",
		X"1E",X"48",X"11",X"00",X"00",X"48",X"1D",X"48",X"19",X"00",X"00",X"C8",X"0E",X"C8",X"0E",X"00",
		X"00",X"C8",X"0E",X"C8",X"0E",X"00",X"00",X"98",X"0E",X"98",X"0E",X"00",X"00",X"98",X"0E",X"98",
		X"0E",X"00",X"00",X"98",X"0E",X"98",X"0E",X"00",X"03",X"C8",X"0E",X"C8",X"0E",X"00",X"00",X"C8",
		X"0E",X"C8",X"0E",X"00",X"00",X"C8",X"0E",X"C8",X"0E",X"00",X"04",X"C8",X"0E",X"C8",X"0E",X"00",
		X"00",X"C8",X"0E",X"C8",X"0E",X"00",X"01",X"C8",X"0E",X"C8",X"0E",X"00",X"00",X"C8",X"0E",X"C8",
		X"0E",X"00",X"00",X"78",X"0E",X"78",X"0E",X"00",X"03",X"78",X"0E",X"78",X"0E",X"00",X"03",X"C8",
		X"0E",X"C8",X"0E",X"00",X"00",X"C8",X"0E",X"C8",X"0E",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
