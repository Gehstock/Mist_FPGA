library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity fg2_rom is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of fg2_rom is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"99",X"99",X"AA",X"AA",X"99",X"99",X"AA",X"AA",X"99",X"99",X"AA",X"AA",X"99",X"99",
		X"55",X"55",X"EE",X"E5",X"88",X"88",X"BB",X"BB",X"99",X"BB",X"77",X"99",X"9A",X"AA",X"AA",X"AA",
		X"55",X"55",X"EE",X"5E",X"88",X"55",X"99",X"88",X"BB",X"B9",X"AA",X"AA",X"AA",X"99",X"99",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"11",X"11",X"11",X"11",X"12",X"12",
		X"21",X"22",X"22",X"22",X"22",X"22",X"23",X"23",X"32",X"32",X"33",X"33",X"33",X"33",X"34",X"34",
		X"43",X"43",X"34",X"34",X"44",X"44",X"45",X"45",X"54",X"54",X"55",X"55",X"55",X"55",X"56",X"56",
		X"65",X"65",X"66",X"66",X"66",X"66",X"67",X"67",X"76",X"76",X"77",X"77",X"77",X"77",X"78",X"78",
		X"87",X"87",X"88",X"88",X"88",X"88",X"89",X"89",X"98",X"98",X"99",X"99",X"99",X"99",X"9A",X"9A",
		X"A9",X"A9",X"AA",X"AA",X"AA",X"AA",X"AB",X"AB",X"BA",X"BA",X"BB",X"BB",X"BB",X"BB",X"BC",X"BC",
		X"CB",X"CB",X"CC",X"CC",X"CC",X"CC",X"CD",X"CD",X"DC",X"DC",X"DD",X"DD",X"DD",X"DD",X"DE",X"DE",
		X"ED",X"ED",X"EE",X"EE",X"EE",X"EE",X"EF",X"EF",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"4A",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"4A",X"04",X"AA",X"4A",X"AA",X"AA",X"AA",X"4A",X"DA",
		X"4A",X"00",X"AA",X"40",X"DA",X"A4",X"AA",X"AA",X"AA",X"A4",X"DA",X"AA",X"AA",X"AA",X"AA",X"DA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"A4",X"40",X"A4",X"A4",X"AA",X"AA",X"AA",X"A4",
		X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"11",X"00",X"11",X"04",X"11",X"41",X"11",X"11",X"11",
		X"00",X"04",X"00",X"41",X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"11",
		X"44",X"44",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"44",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"44",X"44",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"44",X"44",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"44",X"44",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"14",X"00",X"11",X"40",X"11",X"14",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"AA",X"AA",X"AA",X"A4",X"AA",X"AA",X"AA",X"44",X"AA",X"AA",X"AA",X"AA",X"DA",X"44",X"AA",X"A4",
		X"41",X"11",X"A4",X"33",X"43",X"33",X"44",X"43",X"A4",X"33",X"43",X"33",X"33",X"33",X"44",X"44",
		X"AA",X"A4",X"AA",X"4F",X"AA",X"FF",X"AA",X"FF",X"AA",X"44",X"AA",X"84",X"44",X"84",X"40",X"84",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"44",X"44",X"4D",X"DD",X"4D",X"DD",X"4D",X"DD",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"44",X"44",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"44",X"44",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"44",X"44",X"DD",X"DD",X"D4",X"DD",X"D4",X"DD",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"44",X"44",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"44",X"44",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"44",X"44",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"44",X"44",X"DD",X"44",X"DD",X"44",X"DD",X"44",
		X"4C",X"56",X"4C",X"56",X"4C",X"56",X"45",X"66",X"45",X"66",X"85",X"66",X"5E",X"66",X"5E",X"66",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"44",X"44",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"44",X"44",
		X"55",X"88",X"66",X"77",X"66",X"88",X"65",X"55",X"65",X"22",X"59",X"99",X"5B",X"B9",X"99",X"99",
		X"88",X"88",X"77",X"77",X"88",X"85",X"55",X"53",X"22",X"23",X"99",X"93",X"BB",X"93",X"99",X"93",
		X"40",X"84",X"E4",X"84",X"E4",X"84",X"E4",X"84",X"5E",X"84",X"5E",X"84",X"5E",X"84",X"44",X"84",
		X"4D",X"DD",X"4D",X"DD",X"45",X"44",X"48",X"44",X"48",X"44",X"48",X"44",X"48",X"44",X"48",X"44",
		X"04",X"84",X"04",X"84",X"00",X"84",X"00",X"84",X"00",X"84",X"00",X"E4",X"00",X"E4",X"00",X"E4",
		X"48",X"44",X"48",X"44",X"48",X"44",X"44",X"44",X"99",X"99",X"4B",X"44",X"4A",X"44",X"4A",X"44",
		X"D4",X"DD",X"D4",X"DD",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"DD",X"DD",X"DD",X"DD",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"46",X"44",X"88",X"88",X"99",X"99",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"34",X"44",X"34",X"44",X"99",X"99",X"44",X"44",X"44",X"44",X"44",X"44",
		X"DD",X"45",X"DD",X"45",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"45",
		X"5E",X"66",X"E5",X"66",X"E5",X"66",X"E5",X"66",X"56",X"65",X"56",X"65",X"56",X"65",X"55",X"65",
		X"44",X"45",X"44",X"45",X"44",X"4E",X"44",X"4E",X"99",X"4E",X"BB",X"E5",X"4A",X"E5",X"4A",X"E5",
		X"39",X"59",X"39",X"B9",X"39",X"B9",X"39",X"B9",X"39",X"B9",X"32",X"22",X"35",X"55",X"35",X"88",
		X"9B",X"9B",X"9B",X"9B",X"9B",X"9B",X"9B",X"9B",X"9B",X"9B",X"9B",X"9B",X"9B",X"9B",X"9B",X"9B",
		X"B9",X"B3",X"B9",X"B3",X"B9",X"B3",X"B9",X"B3",X"B9",X"B3",X"B9",X"B3",X"B9",X"B3",X"B9",X"B3",
		X"9B",X"9B",X"9B",X"9B",X"9B",X"9B",X"9B",X"9B",X"9B",X"9B",X"22",X"22",X"55",X"55",X"58",X"85",
		X"B9",X"B3",X"B9",X"B3",X"B9",X"B3",X"B9",X"B3",X"B9",X"B3",X"22",X"23",X"55",X"53",X"88",X"53",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",
		X"00",X"00",X"00",X"00",X"99",X"99",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"D9",X"00",X"D9",X"00",X"DD",X"00",
		X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"99",X"99",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"99",X"99",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"9B",X"BB",X"09",X"BB",X"00",X"99",
		X"9D",X"DD",X"9D",X"DD",X"9D",X"DD",X"9D",X"DD",X"99",X"DD",X"BB",X"99",X"BB",X"BB",X"BB",X"BB",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"D9",X"99",X"99",X"BB",X"BB",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"9D",X"00",X"9D",X"00",X"9D",X"00",X"9D",X"00",X"9D",X"00",X"9D",X"00",X"9D",X"00",X"9D",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"99",X"00",X"BB",X"90",X"BB",X"B9",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"00",X"9D",X"00",X"9D",X"00",X"9D",X"00",X"9D",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",
		X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"D9",X"00",X"D9",X"00",X"D9",X"00",X"D9",X"00",
		X"00",X"09",X"00",X"9D",X"00",X"DD",X"00",X"DD",X"09",X"DD",X"09",X"DD",X"09",X"DD",X"09",X"DD",
		X"99",X"90",X"DD",X"D9",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"BB",X"BB",X"99",X"BB",X"DD",X"99",X"DD",X"DD",X"DD",X"DD",X"9D",X"DD",X"09",X"99",X"00",X"DD",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"99",X"9B",X"DD",X"09",X"D9",X"00",X"99",X"90",X"DD",X"D9",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"B9",X"BB",X"99",X"99",X"9D",X"00",X"DD",X"00",X"DD",X"00",X"DD",
		X"00",X"DD",X"99",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"D9",
		X"D9",X"00",X"D9",X"00",X"90",X"00",X"90",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"99",X"00",
		X"09",X"DD",X"09",X"DD",X"09",X"DD",X"09",X"DD",X"09",X"DD",X"09",X"DD",X"9D",X"DD",X"9D",X"DD",
		X"09",X"DD",X"9D",X"DD",X"9D",X"DD",X"9D",X"DD",X"9D",X"DD",X"9D",X"DD",X"9D",X"DD",X"9D",X"DD",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"D9",X"DD",X"9B",X"DD",X"BB",X"DD",X"BB",X"DD",X"BB",X"DD",X"BB",
		X"00",X"9D",X"00",X"09",X"99",X"00",X"BB",X"09",X"BB",X"9B",X"BB",X"B9",X"BB",X"B9",X"BB",X"BB",
		X"DD",X"DD",X"DD",X"DD",X"99",X"DD",X"BB",X"99",X"BB",X"B9",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"DD",X"9D",X"99",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"9D",X"DD",
		X"DD",X"00",X"DD",X"90",X"DD",X"D9",X"DD",X"D9",X"DD",X"D9",X"DD",X"D9",X"DD",X"D9",X"DD",X"D9",
		X"9D",X"DD",X"9D",X"DD",X"9D",X"DD",X"9D",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"9D",X"DD",X"9D",X"DD",X"9D",X"DD",X"9D",X"DD",X"9D",X"DD",X"9D",X"DD",X"9D",X"DD",X"9D",X"DD",
		X"DD",X"BB",X"DD",X"BB",X"DD",X"BB",X"DD",X"BB",X"DD",X"BB",X"DD",X"9B",X"DD",X"D9",X"DD",X"DD",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"9B",X"99",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"99",X"BB",
		X"9D",X"DD",X"B9",X"DD",X"B9",X"DD",X"B9",X"DD",X"B9",X"DD",X"B9",X"DD",X"9D",X"DD",X"DD",X"DD",
		X"DD",X"D9",X"DD",X"D9",X"DD",X"D9",X"DD",X"D9",X"DD",X"D9",X"DD",X"D9",X"DD",X"D9",X"DD",X"D9",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"9D",X"DD",X"9D",X"DD",X"09",X"DD",X"00",X"99",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"D9",X"DD",X"D9",X"DD",X"90",X"DD",X"00",X"99",X"00",
		X"9D",X"DD",X"09",X"DD",X"09",X"DD",X"00",X"DD",X"00",X"9D",X"00",X"09",X"00",X"00",X"00",X"00",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"9D",X"DD",X"09",X"99",
		X"D9",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"99",X"99",
		X"DD",X"99",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"99",X"99",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"99",X"99",
		X"DD",X"D9",X"DD",X"D9",X"DD",X"90",X"DD",X"90",X"DD",X"00",X"DD",X"00",X"99",X"00",X"00",X"00",
		X"09",X"99",X"9D",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"99",X"00",X"DD",X"90",X"DD",X"90",X"DD",X"D9",X"DD",X"D9",X"DD",X"D9",X"DD",X"D9",X"DD",X"D9",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"09",X"00",X"09",
		X"00",X"00",X"09",X"99",X"9D",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"00",X"00",X"99",X"99",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"DD",X"D9",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"D9",X"DD",X"9B",X"D9",X"BB",
		X"00",X"00",X"99",X"99",X"DD",X"9B",X"D9",X"BB",X"9B",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"00",X"00",X"99",X"00",X"BB",X"99",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"90",X"00",
		X"00",X"09",X"00",X"09",X"00",X"09",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"9D",X"DD",X"09",X"99",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"D9",X"DD",X"9B",X"99",X"BB",
		X"DD",X"DD",X"DD",X"D9",X"DD",X"9B",X"D9",X"BB",X"9B",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"9B",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"B9",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"B9",X"BB",X"90",X"B9",X"00",X"90",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"09",X"DD",X"9D",X"DD",X"9D",X"DD",X"DD",X"DD",X"DD",X"D9",X"DD",X"9B",X"D9",X"BB",
		X"99",X"99",X"DD",X"D9",X"DD",X"9B",X"D9",X"BB",X"9B",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"9B",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"B9",X"BB",X"9D",X"B9",X"DD",X"9D",X"DD",X"DD",X"DD",
		X"BB",X"99",X"B9",X"DD",X"9D",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"99",X"99",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"90",X"00",X"D9",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"90",X"DD",X"90",X"DD",X"90",X"DD",X"90",
		X"D9",X"BB",X"9B",X"BB",X"9B",X"BB",X"9B",X"BB",X"9B",X"BB",X"9B",X"BB",X"09",X"BB",X"09",X"BB",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"B9",X"BB",X"9D",X"B9",X"DD",X"9D",X"DD",X"99",X"99",
		X"BB",X"9D",X"B9",X"DD",X"9D",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"99",X"99",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"99",X"99",
		X"DD",X"90",X"DD",X"90",X"DD",X"90",X"DD",X"90",X"DD",X"00",X"DD",X"00",X"D9",X"00",X"90",X"00",
		X"00",X"BB",X"00",X"BB",X"00",X"99",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",
		X"BB",X"9D",X"B9",X"DD",X"9D",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"99",X"D9",X"BB",X"9B",X"BB",X"BB",X"BB",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"9D",X"DD",X"B9",X"DD",X"BB",X"DD",X"BB",X"9D",
		X"DD",X"D9",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"00",X"00",X"00",X"00",X"90",X"00",X"90",X"00",X"D9",X"00",X"D9",X"00",X"D9",X"00",X"D9",X"00",
		X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"D9",X"DD",X"D9",X"99",X"99",X"DD",X"D9",X"DD",X"DD",X"DD",X"DD",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"BB",X"B9",X"BB",X"B9",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"B9",X"BB",X"B9",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"99",X"9D",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"D9",X"00",X"D9",X"00",X"D9",X"00",X"D9",X"00",X"D9",X"00",X"D9",X"00",X"D9",X"00",X"D9",X"00",
		X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"9D",X"00",X"09",X"00",X"00",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"99",X"99",
		X"BB",X"BB",X"9B",X"BB",X"D9",X"BB",X"DD",X"99",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"99",X"99",
		X"D9",X"00",X"D9",X"00",X"D9",X"00",X"90",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",
		X"BB",X"9D",X"BB",X"DD",X"B9",X"DD",X"9D",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"99",X"99",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"D9",X"99",X"90",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"DD",X"09",X"DD",X"9D",X"DD",X"DD",X"DD",
		X"00",X"00",X"00",X"00",X"90",X"00",X"D9",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"90",X"DD",X"90",
		X"00",X"00",X"00",X"09",X"00",X"9D",X"00",X"DD",X"00",X"DD",X"09",X"DD",X"09",X"DD",X"9D",X"DD",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"DD",X"90",X"DD",X"90",X"DD",X"90",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"D9",X"00",X"90",X"00",
		X"9D",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"D9",X"DD",X"D9",X"DD",X"D9",X"DD",X"D9",X"DD",X"DD",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DD",X"DD",X"9D",X"DD",X"9D",X"DD",X"9D",X"DD",X"09",X"DD",X"09",X"DD",X"09",X"DD",X"00",X"DD",
		X"00",X"00",X"00",X"00",X"90",X"00",X"D9",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"90",
		X"00",X"DD",X"00",X"9D",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"9D",
		X"DD",X"DD",X"DD",X"99",X"D9",X"DD",X"9D",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"DD",X"90",X"DD",X"90",X"9D",X"90",X"D9",X"90",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",
		X"00",X"9D",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"09",X"DD",X"09",X"DD",X"09",X"DD",
		X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"D9",X"00",X"90",X"90",X"99",X"D9",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"9D",X"DD",X"9D",X"DD",X"9D",X"DD",X"9D",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"D9",X"DD",X"9D",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"00",X"00",X"90",X"00",X"D9",X"00",X"D9",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",X"DD",X"00",
		X"DD",X"DD",X"9D",X"DD",X"9D",X"DD",X"9D",X"DD",X"09",X"DD",X"09",X"DD",X"00",X"DD",X"00",X"99",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"9D",X"DD",X"9D",X"DD",X"09",X"99",
		X"DD",X"90",X"DD",X"90",X"DD",X"90",X"DD",X"90",X"DD",X"90",X"DD",X"00",X"DD",X"00",X"99",X"00",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"99",X"DD",
		X"89",X"98",X"88",X"88",X"89",X"89",X"88",X"88",X"89",X"88",X"88",X"88",X"89",X"89",X"98",X"88",
		X"99",X"89",X"88",X"88",X"98",X"99",X"88",X"89",X"88",X"99",X"88",X"89",X"98",X"88",X"88",X"89",
		X"98",X"99",X"98",X"88",X"98",X"99",X"98",X"88",X"99",X"88",X"99",X"89",X"98",X"99",X"88",X"90",
		X"99",X"88",X"88",X"88",X"99",X"89",X"88",X"89",X"89",X"99",X"89",X"99",X"89",X"89",X"88",X"88",
		X"99",X"00",X"89",X"99",X"89",X"89",X"89",X"88",X"89",X"89",X"88",X"89",X"89",X"88",X"89",X"89",
		X"88",X"88",X"88",X"89",X"88",X"89",X"88",X"88",X"98",X"99",X"98",X"90",X"88",X"89",X"88",X"89",
		X"89",X"89",X"89",X"89",X"89",X"89",X"88",X"88",X"88",X"89",X"89",X"99",X"99",X"00",X"98",X"00",
		X"88",X"89",X"89",X"98",X"89",X"98",X"89",X"88",X"89",X"88",X"88",X"88",X"89",X"89",X"90",X"90",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"D9",X"09",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"D9",X"00",X"D0",X"00",
		X"09",X"09",X"09",X"09",X"09",X"99",X"00",X"DD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"D0",X"00",X"D0",X"09",X"00",X"99",X"00",X"DD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"99",X"55",X"55",X"55",X"99",X"55",X"99",X"55",X"55",X"55",X"99",X"55",X"99",X"55",X"55",
		X"99",X"99",X"55",X"59",X"99",X"59",X"99",X"59",X"55",X"59",X"99",X"59",X"99",X"59",X"55",X"59",
		X"99",X"99",X"55",X"55",X"55",X"99",X"55",X"55",X"55",X"99",X"55",X"55",X"55",X"99",X"55",X"55",
		X"99",X"90",X"55",X"90",X"95",X"90",X"55",X"90",X"95",X"90",X"55",X"90",X"95",X"90",X"55",X"90",
		X"99",X"09",X"55",X"95",X"95",X"55",X"95",X"59",X"59",X"55",X"55",X"99",X"95",X"55",X"95",X"99",
		X"59",X"00",X"55",X"00",X"55",X"00",X"99",X"90",X"55",X"59",X"99",X"95",X"55",X"59",X"99",X"59",
		X"55",X"99",X"99",X"55",X"90",X"95",X"90",X"95",X"90",X"55",X"90",X"55",X"99",X"59",X"95",X"99",
		X"99",X"59",X"55",X"59",X"99",X"99",X"59",X"00",X"55",X"00",X"55",X"99",X"95",X"55",X"99",X"99",
		X"00",X"09",X"00",X"09",X"00",X"09",X"00",X"09",X"00",X"09",X"00",X"09",X"00",X"09",X"00",X"09",
		X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"50",X"99",X"95",X"55",X"55",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"00",X"00",
		X"00",X"50",X"50",X"95",X"95",X"95",X"59",X"95",X"05",X"95",X"00",X"95",X"00",X"95",X"00",X"50",
		X"AA",X"AA",X"44",X"AA",X"4A",X"AA",X"04",X"AA",X"4A",X"AA",X"AD",X"AD",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"DA",X"AD",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AD",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AD",X"DA",X"AA",X"AD",X"AA",X"AA",
		X"AA",X"AA",X"AD",X"AA",X"AA",X"AD",X"AA",X"AA",X"AD",X"55",X"AA",X"66",X"AA",X"66",X"AA",X"66",
		X"AA",X"AA",X"AD",X"AA",X"AA",X"AA",X"4A",X"DA",X"4A",X"AA",X"04",X"44",X"00",X"00",X"00",X"00",
		X"AA",X"66",X"A5",X"66",X"58",X"56",X"A5",X"56",X"4A",X"85",X"04",X"85",X"00",X"88",X"00",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"88",X"00",X"88",X"00",X"88",X"00",X"88",X"00",X"88",X"00",X"88",X"00",X"88",X"04",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"14",X"00",X"11",X"00",X"11",X"44",X"11",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"44",X"44",
		X"00",X"00",X"40",X"00",X"14",X"00",X"14",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"88",X"77",X"77",X"88",X"85",X"55",X"53",X"22",X"23",X"99",X"93",X"BB",X"93",X"99",X"93",
		X"40",X"00",X"74",X"00",X"40",X"04",X"44",X"43",X"22",X"23",X"99",X"93",X"BB",X"93",X"99",X"93",
		X"B9",X"B3",X"B9",X"B3",X"B9",X"B3",X"B9",X"B3",X"B9",X"B3",X"B9",X"B3",X"B9",X"B3",X"B9",X"B3",
		X"B9",X"B3",X"B9",X"B3",X"B9",X"B3",X"B9",X"B3",X"B9",X"B3",X"B9",X"B3",X"B9",X"B3",X"B9",X"B3",
		X"B9",X"B3",X"B9",X"B3",X"B9",X"B3",X"B9",X"B3",X"B9",X"B3",X"22",X"23",X"54",X"43",X"80",X"43",
		X"B9",X"B3",X"B9",X"B3",X"B9",X"B3",X"B9",X"B3",X"B9",X"B3",X"22",X"23",X"44",X"43",X"00",X"43",
		X"44",X"44",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"44",X"44",
		X"44",X"00",X"66",X"00",X"66",X"40",X"66",X"64",X"66",X"64",X"66",X"40",X"66",X"00",X"44",X"00",
		X"00",X"44",X"44",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"44",X"66",X"00",X"44",
		X"44",X"66",X"00",X"66",X"00",X"46",X"00",X"04",X"00",X"04",X"00",X"46",X"00",X"66",X"44",X"66",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",
		X"66",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"66",X"00",
		X"44",X"44",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"44",X"44",
		X"AA",X"AA",X"99",X"AA",X"AA",X"AA",X"99",X"AA",X"44",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"4A",
		X"47",X"4A",X"47",X"99",X"47",X"AA",X"47",X"44",X"77",X"99",X"74",X"94",X"49",X"4A",X"49",X"99",
		X"4A",X"4A",X"94",X"4A",X"AA",X"4A",X"99",X"4A",X"AA",X"4A",X"99",X"4A",X"AA",X"4A",X"99",X"4A",
		X"49",X"AA",X"49",X"99",X"49",X"AA",X"49",X"99",X"44",X"AA",X"44",X"99",X"44",X"AA",X"44",X"99",
		X"AA",X"AA",X"49",X"99",X"A4",X"AA",X"4A",X"99",X"4A",X"AA",X"94",X"49",X"A4",X"4A",X"94",X"A4",
		X"AA",X"AA",X"99",X"99",X"AA",X"AA",X"99",X"94",X"AA",X"4A",X"99",X"AA",X"AA",X"44",X"99",X"B4",
		X"AA",X"44",X"99",X"74",X"AA",X"74",X"99",X"74",X"AA",X"74",X"94",X"74",X"A4",X"4A",X"94",X"49",
		X"AA",X"B4",X"99",X"49",X"AA",X"4A",X"99",X"99",X"AA",X"AA",X"99",X"99",X"AA",X"AA",X"99",X"99",
		X"AA",X"AA",X"99",X"99",X"AA",X"AA",X"99",X"99",X"4A",X"AA",X"B4",X"99",X"BB",X"AA",X"BB",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"4B",X"AA",X"4B",X"99",X"A4",X"AA",X"94",X"99",X"AA",X"AA",X"99",X"99",X"AA",X"AA",X"99",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"66",X"66",X"99",X"99",X"77",X"77",X"22",X"22",X"66",X"66",X"11",X"11",X"00",X"00",X"00",
		X"66",X"00",X"7C",X"00",X"2C",X"00",X"6C",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"73",X"01",X"73",X"01",X"73",X"01",X"73",X"01",X"73",X"01",X"73",X"01",X"73",X"01",X"73",
		X"95",X"BD",X"95",X"BD",X"95",X"BD",X"95",X"BD",X"95",X"BD",X"95",X"BD",X"95",X"BD",X"95",X"BD",
		X"01",X"73",X"01",X"73",X"01",X"73",X"01",X"73",X"01",X"73",X"01",X"73",X"01",X"73",X"01",X"73",
		X"95",X"BD",X"95",X"BD",X"95",X"BD",X"95",X"BD",X"95",X"BD",X"95",X"BD",X"95",X"BD",X"95",X"BD",
		X"CA",X"48",X"CA",X"48",X"CA",X"48",X"CA",X"48",X"CA",X"48",X"CA",X"48",X"CA",X"48",X"CA",X"48",
		X"26",X"00",X"26",X"00",X"26",X"00",X"26",X"00",X"26",X"00",X"26",X"00",X"26",X"00",X"26",X"00",
		X"CA",X"48",X"CA",X"48",X"CA",X"48",X"CA",X"48",X"CA",X"C4",X"C5",X"CC",X"C5",X"1C",X"51",X"11",
		X"26",X"00",X"26",X"00",X"26",X"00",X"7C",X"11",X"77",X"66",X"33",X"11",X"11",X"33",X"C1",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"12",X"00",X"21",X"00",X"12",X"00",X"21",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"02",X"00",X"21",X"00",X"12",X"00",X"21",
		X"10",X"12",X"20",X"21",X"10",X"12",X"20",X"21",X"12",X"12",X"21",X"21",X"12",X"00",X"21",X"21",
		X"00",X"12",X"00",X"21",X"02",X"12",X"01",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",
		X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",
		X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",
		X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",
		X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"20",
		X"12",X"12",X"21",X"20",X"12",X"06",X"21",X"66",X"10",X"66",X"06",X"66",X"66",X"66",X"66",X"66",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"21",X"44",X"12",X"44",X"21",X"44",X"12",X"44",X"21",X"40",X"12",X"40",X"21",X"40",X"12",
		X"44",X"44",X"00",X"04",X"66",X"60",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",
		X"40",X"21",X"40",X"12",X"40",X"21",X"02",X"12",X"01",X"21",X"02",X"12",X"21",X"21",X"12",X"12",
		X"44",X"40",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"44",X"00",X"44",X"00",X"44",X"00",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"00",X"44",X"00",X"44",X"20",X"44",X"10",X"44",X"20",X"44",X"10",X"44",X"21",X"44",X"12",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"00",X"44",X"33",X"40",X"33",
		X"44",X"44",X"44",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"33",X"03",X"33",X"03",X"33",X"03",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"03",X"00",X"03",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"40",X"44",X"00",X"40",X"00",X"00",X"00",
		X"44",X"44",X"44",X"00",X"44",X"00",X"44",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"30",X"33",X"30",X"33",X"30",X"33",X"00",
		X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"44",X"00",X"44",X"00",X"44",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"40",X"00",X"40",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"40",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"00",X"00",X"00",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"11",X"11",X"44",X"41",X"14",X"41",X"41",X"41",X"44",X"41",X"44",X"41",X"44",X"11",X"11",X"11",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"00",X"44",X"33",X"44",X"33",X"00",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"00",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"77",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"74",X"44",
		X"44",X"44",X"44",X"44",X"44",X"77",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"34",X"44",X"34",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"33",X"34",X"33",X"44",X"44",X"34",X"44",X"43",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"34",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"40",X"44",X"40",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"40",X"00",X"40",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"30",X"00",X"30",X"00",X"30",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"44",X"00",X"44",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"04",X"44",X"00",X"44",
		X"11",X"11",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",
		X"00",X"44",X"00",X"24",X"00",X"99",X"02",X"99",X"29",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"11",X"11",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"11",X"11",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"00",X"40",X"CC",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"22",X"44",X"22",X"44",X"22",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"24",X"44",X"24",X"44",X"24",X"44",X"44",X"44",X"24",X"44",X"42",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"29",X"00",X"29",X"00",X"29",
		X"99",X"29",X"92",X"20",X"92",X"05",X"29",X"55",X"29",X"CC",X"00",X"55",X"CC",X"55",X"CC",X"CC",
		X"00",X"20",X"00",X"0C",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"CC",X"CC",X"CC",X"C5",X"C5",X"55",X"5C",X"55",X"55",X"CC",X"55",X"C5",X"50",X"00",X"00",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"55",X"CC",X"50",X"CC",X"0F",X"CC",X"FF",X"CC",X"FF",
		X"C0",X"44",X"0F",X"04",X"FF",X"F0",X"FF",X"F0",X"FF",X"00",X"00",X"00",X"FF",X"00",X"F0",X"00",
		X"C0",X"FF",X"C0",X"FF",X"0F",X"FF",X"0F",X"F0",X"FF",X"F0",X"FF",X"0F",X"FF",X"0F",X"FF",X"FF",
		X"0F",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"F0",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"00",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"11",X"11",
		X"00",X"44",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"04",X"44",X"00",X"44",X"00",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"FF",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"F0",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"44",X"00",X"44",X"04",X"44",X"04",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"00",X"44",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"04",X"44",
		X"00",X"00",X"00",X"03",X"00",X"33",X"00",X"33",X"03",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"30",X"44",X"33",X"44",X"33",X"04",X"33",X"30",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"66",X"00",X"60",X"11",X"00",X"00",X"11",X"33",X"00",X"33",X"33",X"30",X"33",X"00",X"33",X"00",
		X"03",X"33",X"33",X"00",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"60",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"00",X"60",X"11",X"01",X"10",X"11",X"03",
		X"66",X"01",X"60",X"11",X"00",X"11",X"11",X"10",X"11",X"03",X"11",X"33",X"11",X"33",X"10",X"33",
		X"10",X"33",X"03",X"33",X"33",X"33",X"33",X"33",X"33",X"30",X"33",X"00",X"33",X"00",X"33",X"00",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"60",X"60",X"60",X"66",X"00",X"66",X"60",X"66",X"66",
		X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"02",X"12",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",
		X"60",X"21",X"66",X"12",X"66",X"01",X"66",X"60",X"66",X"60",X"66",X"60",X"66",X"06",X"66",X"06",
		X"21",X"06",X"12",X"66",X"21",X"66",X"10",X"66",X"20",X"66",X"06",X"66",X"06",X"66",X"66",X"66",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"60",X"66",X"01",X"66",X"11",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"40",X"44",X"06",X"44",X"66",X"44",X"66",X"40",X"66",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"00",X"00",X"30",X"00",X"30",
		X"40",X"66",X"06",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"06",X"66",
		X"00",X"03",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"66",X"10",X"66",X"11",X"66",X"01",X"66",X"30",X"06",X"33",X"10",X"33",X"11",X"03",X"01",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"40",X"44",X"03",X"44",X"33",X"44",X"33",X"40",X"33",X"40",X"33",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"03",X"33",X"03",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"44",X"40",X"44",X"40",X"44",X"40",X"44",X"40",X"44",X"03",X"44",X"03",X"44",X"03",X"44",X"03",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"30",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"30",X"33",X"30",
		X"03",X"30",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"03",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"30",X"00",X"33",X"00",X"33",X"00",
		X"06",X"66",X"11",X"66",X"11",X"66",X"01",X"06",X"30",X"10",X"33",X"11",X"33",X"11",X"33",X"00",
		X"66",X"06",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"00",X"66",X"11",X"66",
		X"33",X"33",X"33",X"33",X"03",X"33",X"00",X"33",X"00",X"33",X"00",X"33",X"00",X"00",X"00",X"00",
		X"11",X"00",X"11",X"11",X"00",X"11",X"01",X"11",X"11",X"10",X"11",X"03",X"11",X"33",X"10",X"33",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"60",X"66",X"00",X"66",X"11",X"00",X"11",X"11",X"11",
		X"66",X"11",X"60",X"11",X"01",X"10",X"11",X"03",X"11",X"33",X"11",X"33",X"10",X"33",X"03",X"33",
		X"11",X"10",X"11",X"03",X"10",X"33",X"03",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"30",X"33",X"00",X"33",X"00",X"33",X"00",
		X"03",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"30",X"33",X"00",X"33",X"00",X"33",X"00",
		X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"04",X"44",X"30",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"00",X"33",X"00",X"33",X"00",X"33",X"03",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"33",X"00",X"33",X"00",X"33",X"03",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"30",X"44",X"33",X"44",X"33",X"44",X"33",X"44",X"33",X"44",X"33",X"44",X"33",X"04",X"33",X"04",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"33",X"04",X"33",X"30",X"33",X"30",X"33",X"30",X"33",X"30",X"33",X"33",X"33",X"33",X"33",X"33",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"12",X"00",X"21",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"12",X"00",X"21",X"00",X"12",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"12",X"21",X"21",
		X"00",X"12",X"00",X"21",X"02",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"17",X"21",X"21",
		X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"77",X"88",X"21",X"21",
		X"00",X"00",X"00",X"00",X"00",X"12",X"00",X"20",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",
		X"00",X"00",X"00",X"00",X"02",X"00",X"01",X"00",X"10",X"00",X"21",X"04",X"12",X"04",X"21",X"04",
		X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"88",X"21",
		X"12",X"04",X"21",X"04",X"12",X"44",X"21",X"44",X"12",X"44",X"21",X"44",X"12",X"44",X"21",X"44",
		X"00",X"00",X"00",X"04",X"00",X"44",X"00",X"44",X"44",X"44",X"44",X"44",X"04",X"44",X"40",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"12",X"00",X"21",X"00",X"12",X"00",X"21",X"00",X"12",X"00",X"21",X"00",X"12",X"00",X"21",X"01",
		X"02",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",
		X"12",X"02",X"21",X"01",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",
		X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",
		X"12",X"12",X"21",X"21",X"1A",X"12",X"28",X"A7",X"12",X"88",X"21",X"71",X"12",X"17",X"21",X"21",
		X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"A1",X"7A",X"12",X"80",X"21",X"10",X"88",X"80",X"21",
		X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",
		X"A8",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",
		X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"10",X"21",X"04",
		X"10",X"44",X"20",X"44",X"04",X"44",X"04",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"12",X"44",X"21",X"44",X"12",X"44",X"20",X"44",X"10",X"44",X"20",X"44",X"10",X"44",X"20",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"22",X"44",X"22",X"44",X"22",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"24",X"44",X"24",X"44",X"24",X"44",X"44",X"44",X"24",X"44",X"42",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",
		X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",
		X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"02",X"12",X"20",X"21",
		X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",
		X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",
		X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",
		X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"44",X"12",X"4F",X"21",X"24",
		X"12",X"12",X"21",X"21",X"12",X"00",X"21",X"44",X"12",X"44",X"40",X"44",X"40",X"44",X"04",X"44",
		X"10",X"44",X"20",X"44",X"10",X"44",X"20",X"44",X"10",X"44",X"20",X"44",X"10",X"44",X"20",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"10",X"44",X"04",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"10",X"12",X"20",X"21",X"10",X"02",X"20",X"40",X"10",X"44",X"20",X"40",X"10",X"06",X"20",X"66",
		X"12",X"12",X"21",X"21",X"12",X"12",X"21",X"21",X"12",X"12",X"01",X"21",X"60",X"12",X"66",X"00",
		X"06",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",
		X"12",X"00",X"21",X"44",X"12",X"44",X"21",X"00",X"12",X"66",X"20",X"66",X"06",X"66",X"66",X"66",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"00",X"44",X"66",X"44",X"66",X"44",X"66",X"04",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",
		X"66",X"04",X"66",X"04",X"66",X"00",X"66",X"01",X"66",X"10",X"66",X"03",X"60",X"33",X"11",X"33",
		X"44",X"44",X"44",X"42",X"44",X"44",X"44",X"22",X"44",X"22",X"44",X"22",X"44",X"44",X"44",X"44",
		X"24",X"44",X"24",X"44",X"22",X"44",X"22",X"44",X"24",X"44",X"44",X"44",X"44",X"44",X"24",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"04",X"44",X"00",X"44",
		X"22",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"00",X"40",X"21",X"44",X"00",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"00",X"00",X"00",X"02",X"20",X"21",X"12",X"00",X"01",X"21",X"40",X"12",
		X"44",X"00",X"44",X"12",X"44",X"01",X"44",X"00",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"21",X"04",X"02",X"20",X"40",X"12",X"00",X"01",X"21",X"00",X"12",X"40",X"21",X"44",X"02");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
