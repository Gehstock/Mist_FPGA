library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity dotron_bg_bits_2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of dotron_bg_bits_2 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"02",X"AA",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"0A",X"AA",X"02",X"AA",X"00",X"AA",X"00",X"2A",
		X"00",X"2A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"2A",X"00",X"2A",
		X"00",X"AA",X"00",X"AA",X"02",X"AA",X"0A",X"AA",X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"2A",X"2A",X"AA",
		X"02",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"2A",X"AA",X"02",X"AA",X"00",X"2A",X"00",X"02",X"00",X"00",
		X"0A",X"AA",X"02",X"AA",X"00",X"AA",X"00",X"2A",X"00",X"0A",X"00",X"02",X"00",X"00",X"00",X"00",
		X"2A",X"AA",X"0A",X"AA",X"0A",X"AA",X"02",X"AA",X"02",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",
		X"AA",X"AA",X"00",X"AA",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"2A",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"02",X"AA",
		X"A8",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A8",X"00",X"A8",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"AA",X"80",X"AA",X"00",X"A8",X"00",
		X"AA",X"AA",X"AA",X"80",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"15",X"54",X"14",X"04",X"14",X"04",X"10",X"04",X"10",X"04",X"10",X"04",X"15",X"54",
		X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",
		X"00",X"00",X"15",X"54",X"10",X"04",X"10",X"00",X"15",X"54",X"00",X"14",X"00",X"14",X"15",X"54",
		X"00",X"00",X"05",X"54",X"04",X"00",X"15",X"00",X"14",X"00",X"14",X"00",X"14",X"04",X"15",X"54",
		X"00",X"00",X"04",X"00",X"04",X"04",X"04",X"04",X"04",X"04",X"15",X"54",X"05",X"00",X"05",X"00",
		X"00",X"00",X"15",X"54",X"00",X"04",X"00",X"04",X"15",X"54",X"14",X"00",X"14",X"04",X"15",X"54",
		X"00",X"00",X"15",X"54",X"00",X"04",X"00",X"04",X"15",X"54",X"14",X"04",X"14",X"04",X"15",X"54",
		X"00",X"00",X"15",X"54",X"10",X"00",X"10",X"00",X"14",X"00",X"14",X"00",X"14",X"00",X"14",X"00",
		X"00",X"00",X"05",X"50",X"04",X"10",X"04",X"10",X"15",X"54",X"14",X"04",X"14",X"04",X"15",X"54",
		X"00",X"00",X"15",X"54",X"10",X"04",X"10",X"04",X"15",X"54",X"14",X"00",X"14",X"00",X"15",X"54",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",
		X"00",X"00",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"20",X"00",X"20",X"00",X"00",X"00",X"20",
		X"00",X"00",X"00",X"28",X"00",X"28",X"00",X"00",X"00",X"00",X"00",X"28",X"00",X"28",X"00",X"00",
		X"00",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",
		X"00",X"00",X"2A",X"A8",X"20",X"08",X"20",X"00",X"2A",X"A8",X"00",X"28",X"00",X"28",X"2A",X"A8",
		X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"FF",X"FF",
		X"00",X"00",X"0A",X"A0",X"08",X"20",X"08",X"20",X"2A",X"A8",X"20",X"28",X"20",X"28",X"20",X"28",
		X"00",X"00",X"0A",X"A8",X"08",X"08",X"08",X"08",X"2A",X"A8",X"20",X"28",X"20",X"28",X"2A",X"A8",
		X"00",X"00",X"2A",X"A8",X"20",X"08",X"00",X"08",X"00",X"28",X"00",X"28",X"20",X"28",X"2A",X"A8",
		X"00",X"00",X"0A",X"A8",X"28",X"08",X"20",X"08",X"20",X"28",X"20",X"28",X"28",X"28",X"0A",X"A8",
		X"00",X"00",X"2A",X"A8",X"00",X"08",X"00",X"08",X"2A",X"A8",X"00",X"28",X"00",X"28",X"2A",X"A8",
		X"00",X"00",X"2A",X"A8",X"00",X"08",X"00",X"08",X"2A",X"A8",X"00",X"28",X"00",X"28",X"00",X"28",
		X"00",X"00",X"2A",X"A8",X"20",X"08",X"00",X"08",X"2A",X"28",X"20",X"28",X"20",X"28",X"2A",X"A8",
		X"00",X"00",X"20",X"08",X"20",X"08",X"20",X"08",X"2A",X"A8",X"20",X"28",X"20",X"28",X"20",X"28",
		X"00",X"00",X"00",X"80",X"00",X"80",X"00",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",
		X"00",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"28",X"00",X"28",X"00",X"28",X"08",X"2A",X"A8",
		X"00",X"00",X"28",X"08",X"08",X"08",X"08",X"08",X"0A",X"A8",X"28",X"28",X"20",X"28",X"20",X"28",
		X"00",X"00",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"28",X"00",X"28",X"00",X"28",X"2A",X"A8",
		X"00",X"00",X"2A",X"A8",X"22",X"08",X"22",X"08",X"22",X"28",X"22",X"28",X"22",X"28",X"22",X"28",
		X"00",X"00",X"20",X"A8",X"22",X"88",X"22",X"08",X"22",X"28",X"2A",X"28",X"28",X"28",X"28",X"28",
		X"00",X"00",X"2A",X"A8",X"28",X"08",X"28",X"08",X"20",X"08",X"20",X"08",X"20",X"08",X"2A",X"A8",
		X"00",X"00",X"2A",X"A8",X"20",X"08",X"20",X"08",X"2A",X"A8",X"00",X"28",X"00",X"28",X"00",X"28",
		X"00",X"00",X"2A",X"A8",X"20",X"08",X"20",X"08",X"22",X"08",X"2A",X"08",X"28",X"08",X"2A",X"A8",
		X"00",X"00",X"0A",X"A8",X"08",X"08",X"08",X"08",X"2A",X"A8",X"20",X"28",X"20",X"28",X"20",X"28",
		X"00",X"00",X"2A",X"A8",X"20",X"08",X"00",X"08",X"2A",X"A8",X"28",X"00",X"28",X"08",X"2A",X"A8",
		X"00",X"00",X"2A",X"A8",X"00",X"80",X"00",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",
		X"00",X"00",X"20",X"08",X"20",X"08",X"20",X"08",X"20",X"28",X"20",X"28",X"20",X"28",X"2A",X"A8",
		X"00",X"00",X"20",X"28",X"20",X"28",X"20",X"28",X"08",X"28",X"08",X"20",X"08",X"20",X"0A",X"A0",
		X"00",X"00",X"22",X"08",X"22",X"08",X"22",X"08",X"22",X"28",X"22",X"28",X"22",X"28",X"2A",X"A8",
		X"00",X"00",X"20",X"08",X"20",X"08",X"20",X"20",X"0A",X"80",X"20",X"28",X"20",X"28",X"20",X"28",
		X"00",X"00",X"20",X"08",X"20",X"08",X"28",X"28",X"0A",X"A0",X"02",X"80",X"02",X"80",X"02",X"80",
		X"00",X"00",X"2A",X"A8",X"28",X"08",X"0A",X"00",X"02",X"80",X"00",X"A0",X"20",X"28",X"2A",X"A8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"A8",X"00",X"AA",X"A8",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"80",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",
		X"AA",X"A8",X"AA",X"A0",X"AA",X"A0",X"AA",X"80",X"AA",X"80",X"AA",X"00",X"AA",X"00",X"AA",X"00",
		X"AA",X"A0",X"AA",X"80",X"AA",X"00",X"A8",X"00",X"A0",X"00",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"AA",X"80",X"A8",X"00",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"00",X"AA",X"00",X"AA",X"80",X"AA",X"A0",X"AA",X"A8",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"01",X"55",X"01",X"55",X"01",X"55",X"01",X"55",X"01",X"55",X"01",X"55",X"01",X"55",
		X"01",X"55",X"01",X"55",X"01",X"55",X"01",X"55",X"01",X"55",X"01",X"55",X"01",X"55",X"A1",X"55",
		X"A1",X"55",X"01",X"55",X"01",X"55",X"01",X"55",X"01",X"55",X"01",X"11",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"05",
		X"00",X"05",X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"55",X"00",X"55",X"00",X"55",X"28",X"55",
		X"28",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"88",X"02",X"AA",X"02",X"AA",X"02",X"AA",X"02",X"AA",X"00",X"00",
		X"85",X"54",X"05",X"54",X"05",X"54",X"05",X"54",X"15",X"54",X"11",X"10",X"00",X"00",X"00",X"00",
		X"55",X"40",X"55",X"50",X"55",X"50",X"15",X"50",X"15",X"54",X"05",X"54",X"05",X"54",X"85",X"54",
		X"00",X"05",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",
		X"00",X"00",X"55",X"54",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"55",
		X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"00",
		X"00",X"00",X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"A0",X"00",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"10",X"00",X"00",X"00",X"00",X"22",X"22",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"22",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"00",X"2A",X"00",X"2A",X"00",X"2A",X"00",X"00",
		X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"40",X"00",X"50",X"00",X"54",X"00",X"55",X"00",X"55",X"00",X"55",X"40",
		X"00",X"00",X"00",X"55",X"05",X"55",X"15",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"54",
		X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"00",
		X"00",X"00",X"54",X"00",X"54",X"00",X"54",X"00",X"54",X"00",X"54",X"00",X"54",X"00",X"00",X"00",
		X"55",X"40",X"55",X"00",X"54",X"00",X"50",X"00",X"50",X"00",X"40",X"00",X"40",X"00",X"4A",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",
		X"0A",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",
		X"00",X"10",X"00",X"00",X"00",X"00",X"88",X"88",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"00",X"A0",X"00",X"80",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"05",X"54",X"05",X"54",X"05",X"54",X"15",X"50",X"04",X"40",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"88",X"A2",X"88",X"88",X"88",X"80",X"88",
		X"FF",X"FF",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"FF",X"FF",
		X"A1",X"55",X"01",X"55",X"01",X"55",X"01",X"55",X"00",X"55",X"00",X"44",X"00",X"00",X"00",X"00",
		X"00",X"15",X"00",X"55",X"00",X"55",X"00",X"55",X"01",X"55",X"01",X"55",X"01",X"55",X"A1",X"55",
		X"55",X"02",X"54",X"02",X"50",X"02",X"40",X"02",X"40",X"02",X"00",X"02",X"00",X"02",X"2A",X"AA",
		X"00",X"00",X"01",X"55",X"15",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"50",
		X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"22",X"AA",X"AA",X"2A",X"AA",X"02",X"AA",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"22",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",
		X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"FF",X"FF",
		X"2A",X"AA",X"00",X"02",X"00",X"02",X"40",X"02",X"40",X"02",X"40",X"02",X"00",X"02",X"00",X"02",
		X"AA",X"AA",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",
		X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"05",X"00",X"05",X"00",X"15",
		X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0A",X"00",X"2A",X"00",X"AA",X"00",X"A8",X"02",X"A2",X"02",X"82",X"02",X"82",
		X"02",X"82",X"02",X"82",X"02",X"A2",X"00",X"A8",X"00",X"AA",X"00",X"2A",X"00",X"0A",X"00",X"00",
		X"82",X"80",X"82",X"80",X"8A",X"80",X"2A",X"00",X"AA",X"00",X"A8",X"00",X"A0",X"00",X"00",X"00",
		X"00",X"00",X"A0",X"00",X"A8",X"00",X"AA",X"00",X"2A",X"00",X"8A",X"80",X"82",X"80",X"82",X"80",
		X"2A",X"AA",X"2A",X"AA",X"2A",X"00",X"2A",X"00",X"2A",X"00",X"2A",X"00",X"2A",X"00",X"00",X"00",
		X"00",X"00",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"00",X"2A",X"00",X"2A",X"00",X"2A",X"AA",
		X"00",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",
		X"A0",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"0A",X"A8",X"0A",X"A8",X"0A",X"A8",
		X"00",X"00",X"00",X"2A",X"00",X"2A",X"00",X"2A",X"00",X"2A",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"A8",X"0A",X"A8",X"0A",X"A8",X"8A",X"A8",X"8A",X"A8",X"0A",X"A8",X"0A",X"A8",X"0A",X"A8",
		X"0A",X"A8",X"0A",X"A8",X"0A",X"A8",X"0A",X"A8",X"0A",X"A8",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"A0",X"00",X"A8",X"00",X"AA",X"00",X"AA",X"00",X"2A",X"80",X"0A",X"80",
		X"0A",X"80",X"0A",X"A0",X"02",X"A0",X"A0",X"02",X"AA",X"AA",X"00",X"00",X"80",X"00",X"A0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"00",X"00",X"A0",X"AA",X"A0",X"2A",X"A0",X"0A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"A0",X"00",X"02",X"00",X"02",X"00",X"02",
		X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A0",X"02",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A8",X"00",X"AA",X"00",X"2A",X"80",X"0A",X"A0",X"02",X"A8",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"A2",X"02",X"A8",X"02",X"AA",X"00",X"AA",X"00",X"0A",X"00",X"00",X"00",X"02",X"00",X"02",
		X"8A",X"A0",X"2A",X"80",X"AA",X"80",X"AA",X"00",X"A0",X"00",X"00",X"00",X"80",X"00",X"80",X"00",
		X"2A",X"02",X"2A",X"02",X"28",X"02",X"28",X"AA",X"28",X"AA",X"2A",X"02",X"0A",X"02",X"0A",X"82",
		X"00",X"00",X"00",X"0A",X"00",X"AA",X"02",X"AA",X"02",X"AA",X"0A",X"A8",X"0A",X"A2",X"0A",X"82",
		X"00",X"00",X"A0",X"00",X"AA",X"00",X"AA",X"80",X"AA",X"80",X"2A",X"A0",X"8A",X"A0",X"82",X"A8",
		X"80",X"A8",X"80",X"A8",X"80",X"28",X"AA",X"28",X"AA",X"28",X"80",X"A8",X"80",X"A0",X"82",X"A0",
		X"0A",X"80",X"0A",X"80",X"0A",X"80",X"0A",X"80",X"0A",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"8A",X"80",X"8A",X"8A",X"0A",X"80",X"0A",X"80",X"0A",X"80",
		X"00",X"00",X"00",X"00",X"08",X"00",X"0A",X"00",X"0A",X"80",X"0A",X"A0",X"0A",X"A8",X"0A",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"20",X"20",X"80",X"20",X"80",X"28",X"80",
		X"80",X"00",X"A0",X"00",X"A8",X"00",X"00",X"2A",X"AA",X"80",X"00",X"02",X"00",X"00",X"00",X"00",
		X"02",X"A0",X"02",X"A0",X"02",X"A0",X"A2",X"A2",X"02",X"A2",X"AA",X"A0",X"AA",X"A0",X"2A",X"A0",
		X"0A",X"A0",X"02",X"A0",X"00",X"A0",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"A0",X"02",X"A0",X"02",X"A0",X"02",X"A0",X"02",X"A0",X"02",X"A0",X"02",X"A0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"08",X"08",X"88",X"8A",X"88",X"88",X"8A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2A",X"00",X"22",X"00",X"28",X"00",X"2A",
		X"0A",X"80",X"20",X"20",X"82",X"08",X"88",X"08",X"88",X"08",X"82",X"08",X"20",X"20",X"0A",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"00",X"02",X"00",X"02",X"AA",X"AA",X"AA",X"AA",X"00",X"02",X"00",X"02",X"00",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"A0",X"AA",X"A8",X"00",X"2A",X"00",X"0A",X"00",X"02",
		X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",
		X"00",X"00",X"22",X"A2",X"22",X"22",X"22",X"22",X"22",X"A2",X"20",X"22",X"20",X"22",X"00",X"00",
		X"00",X"00",X"A2",X"A0",X"20",X"20",X"A2",X"A0",X"20",X"20",X"20",X"20",X"A2",X"A0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"20",X"00",X"A0",X"00",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"28",X"00",X"22",X"00",X"22",X"00",X"2A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"08",X"22",X"88",X"22",X"28",X"22",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"28",X"A2",X"28",X"8A",X"20",X"82",X"28",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"80",X"88",X"A2",X"A0",X"88",X"88",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"08",X"88",X"8A",X"8A",X"88",X"88",X"88",
		X"0A",X"80",X"20",X"20",X"82",X"08",X"88",X"88",X"8A",X"88",X"88",X"88",X"20",X"20",X"0A",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"28",X"2A",X"22",X"20",X"2A",X"28",X"22",X"20",X"22",X"20",X"2A",X"20",X"00",X"00",
		X"00",X"00",X"0A",X"00",X"20",X"80",X"20",X"00",X"20",X"00",X"20",X"80",X"0A",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"80",X"88",X"88",X"88",X"22",X"A0",X"22",
		X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"AA",X"AA",
		X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"AA",X"2A",X"80",X"A8",X"00",X"A0",X"00",X"A0",X"00",X"80",X"00",X"80",X"00",X"80",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"08",X"88",X"82",X"0A",X"82",X"08",X"82",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"05",X"50",X"15",X"54",X"55",X"55",X"55",X"55",X"55",X"45",X"55",X"41",
		X"55",X"01",X"15",X"01",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"50",X"00",X"05",X"40",X"00",X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"54",X"00",X"01",X"50",X"00",X"05",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"15",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"54",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"50",X"00",X"05",X"55",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"04",X"00",X"00",
		X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",
		X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"04",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"04",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"10",X"00",X"04",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"10",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"40",X"00",X"00",X"00",X"00",X"04",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"40",X"04",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"0F",X"FF",X"F1",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"0C",X"00",X"F0",
		X"00",X"0C",X"00",X"F0",X"03",X"00",X"0C",X"00",X"F0",X"00",X"00",X"03",X"00",X"0C",X"00",X"30",
		X"01",X"00",X"01",X"00",X"03",X"FF",X"0D",X"00",X"F1",X"00",X"01",X"00",X"01",X"00",X"03",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"0C",X"00",X"F0",X"03",X"00",X"0C",X"00",
		X"03",X"00",X"0C",X"00",X"F0",X"00",X"00",X"00",X"00",X"0F",X"00",X"30",X"00",X"C0",X"03",X"00",
		X"03",X"C0",X"0C",X"00",X"30",X"00",X"C0",X"03",X"00",X"0C",X"00",X"30",X"00",X"C0",X"03",X"00",
		X"0D",X"00",X"31",X"00",X"C1",X"00",X"01",X"00",X"03",X"FF",X"0D",X"00",X"31",X"00",X"C1",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"00",X"00",X"00",X"03",X"00",X"0C",X"00",X"F0",X"03",X"00",X"0C",X"00",X"F0",X"00",X"00",X"00",
		X"F0",X"00",X"00",X"00",X"00",X"03",X"00",X"0C",X"00",X"F0",X"03",X"00",X"0C",X"00",X"30",X"00",
		X"3C",X"00",X"C0",X"00",X"00",X"03",X"00",X"0C",X"00",X"30",X"00",X"C0",X"03",X"00",X"0C",X"00",
		X"3C",X"03",X"C0",X"0C",X"00",X"30",X"00",X"C0",X"03",X"00",X"0C",X"02",X"30",X"08",X"C0",X"08",
		X"01",X"00",X"02",X"AA",X"09",X"00",X"21",X"00",X"81",X"00",X"01",X"00",X"02",X"AA",X"09",X"00",
		X"00",X"00",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"00",X"00",
		X"02",X"AA",X"00",X"0A",X"00",X"00",X"00",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"0C",X"00",X"F0",
		X"00",X"0C",X"00",X"F0",X"03",X"00",X"0C",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"00",X"03",X"00",X"0C",X"00",X"30",X"00",X"C0",X"0F",X"00",X"30",X"00",X"C0",X"00",X"00",X"00",
		X"C0",X"00",X"00",X"03",X"00",X"0C",X"00",X"30",X"00",X"C0",X"03",X"00",X"0C",X"00",X"30",X"00",
		X"30",X"03",X"C0",X"0C",X"00",X"30",X"00",X"C0",X"03",X"00",X"0C",X"00",X"30",X"00",X"C0",X"02",
		X"00",X"20",X"00",X"80",X"02",X"00",X"08",X"02",X"20",X"08",X"80",X"20",X"80",X"80",X"00",X"80",
		X"21",X"00",X"21",X"00",X"81",X"00",X"01",X"55",X"05",X"00",X"11",X"00",X"11",X"00",X"41",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"42",X"AA",X"40",X"0A",X"40",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"0C",X"00",X"F0",X"03",X"00",X"0C",X"00",
		X"03",X"00",X"0C",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"0C",X"00",X"30",
		X"00",X"3C",X"00",X"C0",X"03",X"00",X"0C",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"00",X"3C",X"00",X"C0",X"03",X"00",X"0C",X"00",X"30",X"00",X"C0",X"00",
		X"C0",X"03",X"00",X"0C",X"00",X"30",X"00",X"C0",X"03",X"00",X"0C",X"00",X"30",X"00",X"C0",X"02",
		X"00",X"08",X"00",X"20",X"00",X"80",X"02",X"00",X"08",X"02",X"20",X"02",X"80",X"08",X"00",X"20",
		X"02",X"01",X"08",X"04",X"20",X"04",X"80",X"10",X"00",X"40",X"01",X"00",X"01",X"00",X"04",X"00",
		X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"00",X"40",X"00",X"40",X"00",X"15",X"55",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",
		X"02",X"AA",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"40",X"00",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"00",X"00",X"00",X"03",X"00",X"0C",X"00",X"F0",X"03",X"00",X"0C",X"00",X"F0",X"00",X"00",X"00",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"30",X"00",X"C0",X"03",X"00",
		X"03",X"C0",X"0C",X"00",X"30",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"00",X"03",X"00",X"0C",X"00",X"F0",X"03",X"00",X"0C",X"00",X"30",X"00",X"C0",X"00",X"00",X"00",
		X"00",X"03",X"00",X"0C",X"00",X"30",X"00",X"C0",X"03",X"00",X"0C",X"00",X"30",X"00",X"C0",X"00",
		X"00",X"08",X"00",X"08",X"00",X"20",X"00",X"80",X"02",X"00",X"08",X"00",X"20",X"02",X"80",X"08",
		X"00",X"80",X"02",X"00",X"08",X"00",X"08",X"01",X"20",X"04",X"80",X"10",X"00",X"10",X"00",X"40",
		X"10",X"00",X"40",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"AA",X"40",X"00",X"40",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"42",X"AA",X"40",X"0A",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",
		X"00",X"0C",X"00",X"F0",X"03",X"00",X"0C",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"0C",X"00",X"F0",X"03",X"00",X"0C",X"00",X"30",X"00",
		X"3C",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"0C",
		X"00",X"0C",X"00",X"30",X"00",X"C0",X"0F",X"00",X"30",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"00",X"0C",X"00",X"30",X"00",X"C0",X"03",X"00",X"0C",X"00",X"30",X"00",X"C0",X"00",
		X"00",X"02",X"00",X"08",X"00",X"20",X"00",X"80",X"00",X"80",X"02",X"00",X"08",X"00",X"20",X"00",
		X"00",X"20",X"00",X"20",X"00",X"80",X"02",X"00",X"08",X"00",X"20",X"01",X"80",X"01",X"80",X"04",
		X"01",X"00",X"04",X"00",X"04",X"00",X"10",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",
		X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",
		X"00",X"03",X"00",X"0C",X"00",X"30",X"00",X"C0",X"0F",X"00",X"30",X"00",X"C0",X"00",X"00",X"00",
		X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"0C",X"00",X"30",
		X"00",X"30",X"00",X"C0",X"03",X"00",X"3C",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"00",X"0C",X"00",X"30",X"00",X"C0",X"03",X"00",X"0C",X"00",X"30",X"00",X"C0",X"00",
		X"00",X"00",X"00",X"02",X"00",X"08",X"00",X"20",X"00",X"80",X"02",X"00",X"08",X"00",X"08",X"00",
		X"80",X"02",X"00",X"08",X"00",X"20",X"00",X"80",X"02",X"00",X"02",X"00",X"08",X"00",X"20",X"00",
		X"00",X"10",X"00",X"40",X"00",X"40",X"01",X"00",X"04",X"00",X"10",X"00",X"10",X"00",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"00",X"40",X"00",X"40",X"00",X"55",X"55",X"6A",X"AA",X"6A",X"AA",X"6A",X"AA",X"6A",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"6A",X"A8",X"6A",X"AA",X"6A",X"AA",X"6A",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"15",X"55",X"6A",X"AA",X"6A",X"AA",X"6A",X"AA",X"6A",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"40",X"00",X"40",X"00",X"40",X"55",X"40",X"AA",X"40",X"AA",X"90",X"AA",X"90",X"AA",X"A4",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"0C",X"00",X"30",X"00",X"C0",
		X"00",X"C0",X"03",X"00",X"0C",X"00",X"30",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"00",X"0C",X"00",X"30",X"00",X"C0",X"03",X"00",X"0C",X"00",X"30",X"00",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"08",X"00",X"20",X"00",X"80",X"02",X"00",X"08",X"00",
		X"20",X"00",X"80",X"02",X"00",X"08",X"00",X"08",X"00",X"20",X"00",X"80",X"02",X"00",X"08",X"00",
		X"80",X"01",X"00",X"04",X"00",X"04",X"00",X"10",X"00",X"40",X"01",X"00",X"01",X"00",X"04",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"6A",X"AA",X"6A",X"AA",X"6A",X"AA",X"6A",X"AA",X"6A",X"AA",X"6A",X"AA",X"6A",X"AA",X"6A",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"6A",X"AA",X"6A",X"AA",X"6A",X"AA",X"6A",X"AA",
		X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"6A",X"AA",X"6A",X"AA",X"6A",X"AA",X"6A",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"A4",X"AA",X"A9",X"AA",X"A9",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"40",X"00",X"90",X"00",X"90",X"00",X"A4",X"00",
		X"03",X"00",X"0C",X"00",X"30",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"00",X"0C",X"00",X"30",X"00",X"C0",X"03",X"00",X"0C",X"00",X"30",X"00",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"08",X"00",X"20",X"00",X"80",X"02",X"00",
		X"20",X"00",X"80",X"00",X"80",X"00",X"00",X"02",X"00",X"08",X"00",X"20",X"00",X"80",X"00",X"80",
		X"20",X"00",X"20",X"00",X"80",X"00",X"00",X"01",X"00",X"04",X"00",X"10",X"00",X"10",X"00",X"40",
		X"10",X"00",X"40",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"80",X"A8",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"AA",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",
		X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"40",X"00",X"40",X"00",
		X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"40",X"00",X"40",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"AA",X"00",X"A0",X"00",X"80",X"00",X"00",X"00",X"00",X"00",
		X"A8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"AA",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"2A",X"AA",X"02",X"AA",X"00",X"2A",X"00",X"0A",X"00",X"02",X"00",X"00",
		X"A4",X"00",X"A9",X"00",X"A9",X"00",X"AA",X"40",X"AA",X"40",X"AA",X"90",X"AA",X"90",X"AA",X"A4",
		X"00",X"03",X"00",X"0C",X"00",X"30",X"00",X"C0",X"03",X"00",X"0C",X"00",X"30",X"00",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"08",X"00",X"08",X"00",X"20",X"00",X"80",
		X"08",X"00",X"20",X"00",X"80",X"00",X"00",X"00",X"00",X"02",X"00",X"02",X"00",X"08",X"00",X"20",
		X"02",X"00",X"08",X"00",X"20",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"04",
		X"01",X"00",X"04",X"00",X"04",X"00",X"10",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"A8",X"00",X"AA",X"80",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"00",
		X"00",X"00",X"80",X"00",X"A0",X"00",X"A8",X"00",X"AA",X"80",X"AA",X"A8",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"AA",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2A",
		X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"0A",X"00",X"AA",X"0A",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"A4",X"AA",X"A9",X"AA",X"A9",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"40",X"00",X"90",X"00",X"90",X"00",X"A4",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"08",X"00",X"20",X"00",X"80",
		X"02",X"00",X"08",X"00",X"20",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"08",
		X"00",X"80",X"02",X"00",X"08",X"00",X"08",X"00",X"20",X"00",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"10",X"00",X"40",X"00",X"40",X"01",X"00",X"04",X"00",X"10",X"00",X"10",X"00",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"A4",X"00",X"A9",X"00",X"A9",X"00",X"AA",X"40",X"AA",X"40",X"AA",X"90",X"AA",X"90",X"AA",X"A4",
		X"00",X"80",X"02",X"00",X"08",X"00",X"20",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"20",X"00",X"20",X"00",X"80",X"02",X"00",X"08",X"00",X"20",X"00",X"80",X"00",X"80",X"00",
		X"00",X"01",X"00",X"04",X"00",X"04",X"00",X"10",X"00",X"40",X"01",X"00",X"01",X"00",X"04",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"00",X"08",X"00",X"20",X"00",X"80",X"02",X"00",X"02",X"00",X"08",X"00",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"04",X"00",X"10",X"00",X"40",
		X"04",X"00",X"10",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"04",
		X"00",X"40",X"01",X"00",X"04",X"00",X"10",X"00",X"10",X"00",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"00",X"10",X"00",X"40",X"01",X"00",X"01",X"00",X"04",X"00",X"10",X"00",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",
		X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",
		X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"50",X"2A",
		X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"00",X"2A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"00",
		X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"5A",X"AA",X"50",X"2A",
		X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"00",X"2A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"AA",X"00",X"A8",X"00",X"A0",X"00",
		X"AA",X"A8",X"AA",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"AA",X"A0",X"AA",X"A0",X"AA",X"80",X"AA",X"80",X"AA",X"00",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1A",X"AA",X"6A",X"AA",X"6A",X"A8",X"AA",X"A0",X"AA",X"A0",X"AA",X"80",X"AA",X"80",X"AA",X"00",
		X"6A",X"AA",X"6A",X"AA",X"6A",X"AA",X"6A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"AA",
		X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",
		X"40",X"00",X"40",X"00",X"40",X"00",X"55",X"55",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",
		X"40",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"40",X"00",
		X"40",X"00",X"40",X"00",X"00",X"00",X"15",X"55",X"00",X"00",X"00",X"00",X"40",X"00",X"40",X"00",
		X"AA",X"AA",X"AA",X"AA",X"2A",X"AA",X"0A",X"AA",X"0A",X"AA",X"02",X"AA",X"02",X"AA",X"00",X"AA",
		X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"0A",X"AA",X"00",X"AA",X"00",X"2A",X"00",X"0A",
		X"2A",X"AA",X"00",X"AA",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1A",X"AA",X"6A",X"AA",X"6A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"01",X"00",X"15",X"40",X"01",X"10",X"01",X"00",X"01",X"00",X"04",X"40",X"04",X"40",X"04",X"10");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
