library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity crater_ch_bits is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of crater_ch_bits is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"C0",X"01",X"C0",X"01",X"C0",X"01",X"C0",X"01",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"C0",X"05",X"C0",X"05",X"C0",X"05",X"C0",X"05",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"C0",X"15",X"C0",X"15",X"C0",X"15",X"C0",X"15",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"C0",X"55",X"C0",X"55",X"C0",X"55",X"C0",X"55",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"C1",X"55",X"C1",X"55",X"C1",X"55",X"C1",X"55",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"C5",X"55",X"C5",X"55",X"C5",X"55",X"C5",X"55",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"D5",X"55",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"15",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"55",X"01",X"55",X"01",X"55",X"01",X"55",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"05",X"55",X"05",X"55",X"05",X"55",X"05",X"55",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"15",X"55",X"15",X"55",X"15",X"55",X"15",X"55",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"07",X"00",X"07",X"00",X"07",X"00",X"07",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"17",X"00",X"17",X"00",X"17",X"00",X"17",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"57",X"00",X"57",X"00",X"57",X"00",X"57",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"01",X"57",X"01",X"57",X"01",X"57",X"01",X"57",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"05",X"57",X"05",X"57",X"05",X"57",X"05",X"57",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"15",X"57",X"15",X"57",X"15",X"57",X"15",X"57",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"55",X"57",X"55",X"57",X"55",X"57",X"55",X"57",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"FF",X"FF",
		X"00",X"00",X"00",X"10",X"00",X"50",X"01",X"50",X"05",X"50",X"00",X"10",X"00",X"10",X"00",X"10",
		X"00",X"00",X"00",X"30",X"00",X"F0",X"03",X"F0",X"0F",X"F0",X"00",X"30",X"00",X"30",X"00",X"30",
		X"00",X"C0",X"30",X"C3",X"30",X"C3",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"33",X"F3",X"30",X"03",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"03",X"C0",X"03",X"C0",X"3F",X"FC",X"3F",X"FC",X"03",X"C0",X"03",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"3F",X"FC",X"00",X"00",X"00",X"00",X"3F",X"FC",X"00",X"00",X"00",X"00",
		X"00",X"00",X"30",X"0C",X"0C",X"30",X"03",X"C0",X"0C",X"30",X"30",X"0C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0C",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"0C",X"00",X"00",X"00",
		X"FF",X"FF",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"FF",X"FF",
		X"00",X"00",X"0F",X"C0",X"0F",X"C0",X"03",X"00",X"3F",X"F0",X"03",X"00",X"0C",X"C0",X"30",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"3F",X"FC",X"3C",X"0C",X"3C",X"0C",X"30",X"0C",X"30",X"0C",X"30",X"0C",X"3F",X"FC",
		X"00",X"00",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",
		X"00",X"00",X"3F",X"FC",X"30",X"0C",X"30",X"00",X"3F",X"FC",X"00",X"3C",X"00",X"3C",X"3F",X"FC",
		X"00",X"00",X"0F",X"FC",X"0C",X"00",X"3F",X"00",X"3C",X"00",X"3C",X"00",X"3C",X"0C",X"3F",X"FC",
		X"00",X"00",X"0C",X"00",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"3F",X"FC",X"0F",X"00",X"0F",X"00",
		X"00",X"00",X"3F",X"FC",X"00",X"0C",X"00",X"0C",X"3F",X"FC",X"3C",X"00",X"3C",X"0C",X"3F",X"FC",
		X"00",X"00",X"3F",X"FC",X"00",X"0C",X"00",X"0C",X"3F",X"FC",X"3C",X"0C",X"3C",X"0C",X"3F",X"FC",
		X"00",X"00",X"3F",X"FC",X"30",X"00",X"30",X"00",X"3C",X"00",X"3C",X"00",X"3C",X"00",X"3C",X"00",
		X"00",X"00",X"0F",X"F0",X"0C",X"30",X"0C",X"30",X"3F",X"FC",X"3C",X"0C",X"3C",X"0C",X"3F",X"FC",
		X"00",X"00",X"3F",X"FC",X"30",X"0C",X"30",X"0C",X"3F",X"FC",X"3C",X"00",X"3C",X"00",X"3F",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"F0",X"0C",X"30",X"0C",X"30",X"3F",X"FC",X"30",X"3C",X"30",X"3C",X"30",X"3C",
		X"00",X"00",X"0F",X"FC",X"0C",X"0C",X"0C",X"0C",X"3F",X"FC",X"30",X"3C",X"30",X"3C",X"3F",X"FC",
		X"00",X"00",X"3F",X"FC",X"30",X"0C",X"00",X"0C",X"00",X"3C",X"00",X"3C",X"30",X"3C",X"3F",X"FC",
		X"00",X"00",X"0F",X"FC",X"3C",X"0C",X"30",X"0C",X"30",X"3C",X"30",X"3C",X"3C",X"3C",X"0F",X"FC",
		X"00",X"00",X"3F",X"FC",X"00",X"0C",X"00",X"0C",X"3F",X"FC",X"00",X"3C",X"00",X"3C",X"3F",X"FC",
		X"00",X"00",X"3F",X"FC",X"00",X"0C",X"00",X"0C",X"3F",X"FC",X"00",X"3C",X"00",X"3C",X"00",X"3C",
		X"00",X"00",X"3F",X"FC",X"30",X"0C",X"00",X"0C",X"3F",X"3C",X"30",X"3C",X"30",X"3C",X"3F",X"FC",
		X"00",X"00",X"30",X"0C",X"30",X"0C",X"30",X"0C",X"3F",X"FC",X"30",X"3C",X"30",X"3C",X"30",X"3C",
		X"00",X"00",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",
		X"00",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"3C",X"00",X"3C",X"00",X"3C",X"0C",X"3F",X"FC",
		X"00",X"00",X"3C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0F",X"FC",X"3C",X"3C",X"30",X"3C",X"30",X"3C",
		X"00",X"00",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"3C",X"00",X"3C",X"00",X"3C",X"3F",X"FC",
		X"00",X"00",X"3F",X"FC",X"33",X"0C",X"33",X"0C",X"33",X"3C",X"33",X"3C",X"33",X"3C",X"33",X"3C",
		X"00",X"00",X"30",X"FC",X"33",X"CC",X"33",X"0C",X"33",X"3C",X"3F",X"3C",X"3C",X"3C",X"3C",X"3C",
		X"00",X"00",X"3F",X"FC",X"3C",X"0C",X"3C",X"0C",X"30",X"0C",X"30",X"0C",X"30",X"0C",X"3F",X"FC",
		X"00",X"00",X"3F",X"FC",X"30",X"0C",X"30",X"0C",X"3F",X"FC",X"00",X"3C",X"00",X"3C",X"00",X"3C",
		X"00",X"00",X"3F",X"FC",X"30",X"0C",X"30",X"0C",X"33",X"0C",X"3F",X"0C",X"3C",X"0C",X"3F",X"FC",
		X"00",X"00",X"0F",X"FC",X"0C",X"0C",X"0C",X"0C",X"3F",X"FC",X"30",X"3C",X"30",X"3C",X"30",X"3C",
		X"00",X"00",X"3F",X"FC",X"30",X"0C",X"00",X"0C",X"3F",X"FC",X"3C",X"00",X"3C",X"0C",X"3F",X"FC",
		X"00",X"00",X"3F",X"FC",X"00",X"C0",X"00",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",
		X"00",X"00",X"30",X"0C",X"30",X"0C",X"30",X"0C",X"30",X"3C",X"30",X"3C",X"30",X"3C",X"3F",X"FC",
		X"00",X"00",X"30",X"3C",X"30",X"3C",X"30",X"3C",X"0C",X"3C",X"0C",X"30",X"0C",X"30",X"0F",X"F0",
		X"00",X"00",X"33",X"0C",X"33",X"0C",X"33",X"0C",X"33",X"3C",X"33",X"3C",X"33",X"3C",X"3F",X"FC",
		X"00",X"00",X"30",X"0C",X"30",X"0C",X"30",X"30",X"0F",X"C0",X"30",X"3C",X"30",X"3C",X"30",X"3C",
		X"00",X"00",X"30",X"0C",X"30",X"0C",X"3C",X"3C",X"0F",X"F0",X"03",X"C0",X"03",X"C0",X"03",X"C0",
		X"00",X"00",X"3F",X"FC",X"3C",X"0C",X"0F",X"00",X"03",X"C0",X"00",X"F0",X"30",X"3C",X"3F",X"FC",
		X"00",X"00",X"15",X"54",X"14",X"04",X"14",X"04",X"10",X"04",X"10",X"04",X"10",X"04",X"15",X"54",
		X"00",X"00",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",
		X"00",X"00",X"15",X"54",X"10",X"04",X"10",X"00",X"15",X"54",X"00",X"14",X"00",X"14",X"15",X"54",
		X"00",X"00",X"05",X"54",X"04",X"00",X"15",X"00",X"14",X"00",X"14",X"00",X"14",X"04",X"15",X"54",
		X"00",X"00",X"04",X"00",X"04",X"04",X"04",X"04",X"04",X"04",X"15",X"54",X"05",X"00",X"05",X"00",
		X"00",X"00",X"15",X"54",X"00",X"04",X"00",X"04",X"15",X"54",X"14",X"00",X"14",X"04",X"15",X"54",
		X"00",X"00",X"15",X"54",X"00",X"04",X"00",X"04",X"15",X"54",X"14",X"04",X"14",X"04",X"15",X"54",
		X"00",X"00",X"15",X"54",X"10",X"00",X"10",X"00",X"14",X"00",X"14",X"00",X"14",X"00",X"14",X"00",
		X"00",X"00",X"05",X"50",X"04",X"10",X"04",X"10",X"15",X"54",X"14",X"04",X"14",X"04",X"15",X"54",
		X"00",X"00",X"15",X"54",X"10",X"04",X"10",X"04",X"15",X"54",X"14",X"00",X"14",X"00",X"15",X"54",
		X"00",X"00",X"05",X"50",X"04",X"10",X"04",X"10",X"15",X"54",X"10",X"14",X"10",X"14",X"10",X"14",
		X"00",X"00",X"05",X"54",X"04",X"04",X"04",X"04",X"15",X"54",X"10",X"14",X"10",X"14",X"15",X"54",
		X"00",X"00",X"15",X"54",X"10",X"04",X"00",X"04",X"00",X"14",X"00",X"14",X"10",X"14",X"15",X"54",
		X"00",X"00",X"05",X"54",X"14",X"04",X"10",X"04",X"10",X"14",X"10",X"14",X"14",X"14",X"05",X"54",
		X"00",X"00",X"15",X"54",X"00",X"04",X"00",X"04",X"15",X"54",X"00",X"14",X"00",X"14",X"15",X"54",
		X"00",X"00",X"15",X"54",X"00",X"04",X"00",X"04",X"15",X"54",X"00",X"14",X"00",X"14",X"00",X"14",
		X"00",X"00",X"15",X"54",X"10",X"04",X"00",X"04",X"15",X"14",X"10",X"14",X"10",X"14",X"15",X"54",
		X"00",X"00",X"10",X"04",X"10",X"04",X"10",X"04",X"15",X"54",X"10",X"14",X"10",X"14",X"10",X"14",
		X"00",X"00",X"00",X"40",X"00",X"40",X"00",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",
		X"00",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"14",X"00",X"14",X"00",X"14",X"04",X"15",X"54",
		X"00",X"00",X"14",X"04",X"04",X"04",X"04",X"04",X"05",X"54",X"14",X"14",X"10",X"14",X"10",X"14",
		X"00",X"00",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"14",X"00",X"14",X"00",X"14",X"15",X"54",
		X"00",X"00",X"15",X"54",X"11",X"04",X"11",X"04",X"11",X"14",X"11",X"14",X"11",X"14",X"11",X"14",
		X"00",X"00",X"10",X"54",X"11",X"44",X"11",X"04",X"11",X"14",X"15",X"14",X"14",X"14",X"14",X"14",
		X"00",X"00",X"15",X"54",X"14",X"04",X"14",X"04",X"10",X"04",X"10",X"04",X"10",X"04",X"15",X"54",
		X"00",X"00",X"15",X"54",X"10",X"04",X"10",X"04",X"15",X"54",X"00",X"14",X"00",X"14",X"00",X"14",
		X"00",X"00",X"15",X"54",X"10",X"04",X"10",X"04",X"11",X"04",X"15",X"04",X"14",X"04",X"15",X"54",
		X"00",X"00",X"05",X"54",X"04",X"04",X"04",X"04",X"15",X"54",X"10",X"14",X"10",X"14",X"10",X"14",
		X"00",X"00",X"15",X"54",X"10",X"04",X"00",X"04",X"15",X"54",X"14",X"00",X"14",X"04",X"15",X"54",
		X"00",X"00",X"15",X"54",X"00",X"40",X"00",X"40",X"01",X"40",X"01",X"40",X"01",X"40",X"01",X"40",
		X"00",X"00",X"10",X"04",X"10",X"04",X"10",X"04",X"10",X"14",X"10",X"14",X"10",X"14",X"15",X"54",
		X"00",X"00",X"10",X"14",X"10",X"14",X"10",X"14",X"04",X"14",X"04",X"10",X"04",X"10",X"05",X"50",
		X"00",X"00",X"11",X"04",X"11",X"04",X"11",X"04",X"11",X"14",X"11",X"14",X"11",X"14",X"15",X"54",
		X"00",X"00",X"10",X"04",X"10",X"04",X"10",X"10",X"05",X"40",X"10",X"14",X"10",X"14",X"10",X"14",
		X"00",X"00",X"10",X"04",X"10",X"04",X"14",X"14",X"05",X"50",X"01",X"40",X"01",X"40",X"01",X"40",
		X"00",X"00",X"15",X"54",X"14",X"04",X"05",X"00",X"01",X"40",X"00",X"50",X"10",X"14",X"15",X"54",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
