library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity fg_sp_graphx_3 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of fg_sp_graphx_3 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"90",X"10",X"FC",X"FE",X"FE",X"FE",X"FF",X"FF",X"FE",X"FE",X"FE",X"FC",X"D0",X"10",X"00",
		X"03",X"06",X"06",X"1F",X"9F",X"FF",X"FF",X"1F",X"1F",X"0F",X"7F",X"7F",X"5F",X"06",X"16",X"0C",
		X"00",X"10",X"10",X"FC",X"FE",X"FE",X"FE",X"FF",X"FF",X"FE",X"FE",X"FE",X"FC",X"D0",X"90",X"00",
		X"0C",X"16",X"06",X"1F",X"5F",X"7F",X"7F",X"1F",X"1F",X"0F",X"FF",X"FF",X"9F",X"06",X"06",X"03",
		X"00",X"10",X"10",X"FC",X"FE",X"FE",X"FE",X"FF",X"FF",X"FE",X"FE",X"FE",X"FC",X"10",X"90",X"00",
		X"0C",X"16",X"06",X"5F",X"7F",X"7F",X"1F",X"1F",X"1F",X"FF",X"FF",X"9F",X"1F",X"06",X"06",X"03",
		X"00",X"90",X"10",X"FC",X"FE",X"FE",X"FE",X"FF",X"FF",X"FE",X"FE",X"FE",X"FC",X"10",X"10",X"00",
		X"03",X"06",X"06",X"9F",X"FF",X"FF",X"1F",X"1F",X"1F",X"7F",X"7F",X"5F",X"1F",X"06",X"16",X"0C",
		X"00",X"E0",X"F8",X"FE",X"FE",X"FF",X"FF",X"FE",X"FE",X"FE",X"FC",X"D0",X"10",X"00",X"00",X"00",
		X"00",X"1F",X"9F",X"FF",X"FF",X"1F",X"1F",X"0F",X"7F",X"7F",X"5F",X"06",X"16",X"0C",X"00",X"00",
		X"00",X"C0",X"F8",X"FE",X"FF",X"FF",X"FF",X"FF",X"FE",X"68",X"48",X"80",X"00",X"00",X"00",X"00",
		X"00",X"3F",X"3F",X"0F",X"0F",X"07",X"7F",X"7F",X"4F",X"03",X"03",X"01",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"F8",X"FE",X"FF",X"FF",X"FF",X"B4",X"84",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"07",X"03",X"1F",X"1F",X"17",X"01",X"05",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"F8",X"FE",X"FF",X"DA",X"D2",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"1F",X"1F",X"13",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"D2",X"C2",X"FF",X"FE",X"F8",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"13",X"1F",X"1F",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"84",X"84",X"FF",X"FF",X"FF",X"FE",X"F8",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"05",X"01",X"17",X"1F",X"1F",X"07",X"07",X"07",X"00",
		X"00",X"00",X"00",X"00",X"80",X"48",X"08",X"FE",X"FF",X"FF",X"FF",X"FF",X"FE",X"F8",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"4F",X"7F",X"7F",X"0F",X"0F",X"0F",X"3F",X"3F",X"00",
		X"00",X"00",X"00",X"10",X"10",X"FC",X"FE",X"FE",X"FE",X"FF",X"FF",X"FE",X"FE",X"F8",X"C0",X"00",
		X"00",X"00",X"0C",X"16",X"06",X"5F",X"7F",X"7F",X"1F",X"1F",X"1F",X"FF",X"FF",X"9F",X"1F",X"00",
		X"C0",X"60",X"E1",X"FB",X"FE",X"FC",X"F8",X"F8",X"F8",X"F8",X"FC",X"FE",X"FB",X"E1",X"60",X"C0",
		X"20",X"A1",X"50",X"5F",X"BF",X"7F",X"3F",X"BF",X"7F",X"BF",X"3F",X"7F",X"BF",X"50",X"51",X"88",
		X"00",X"80",X"C0",X"F0",X"F1",X"FF",X"FF",X"F0",X"F0",X"FF",X"FF",X"F1",X"F0",X"C0",X"80",X"00",
		X"40",X"27",X"A1",X"7F",X"7F",X"7F",X"7F",X"FF",X"7F",X"7F",X"FF",X"7F",X"BF",X"21",X"47",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"F0",X"FC",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"F8",
		X"F0",X"DC",X"92",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"93",X"DF",X"F0",
		X"00",X"01",X"07",X"1F",X"9F",X"FF",X"FF",X"1F",X"1F",X"FF",X"FF",X"9F",X"1F",X"07",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"C0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"E0",X"C0",X"00",X"00",
		X"80",X"4F",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"4F",X"80",
		X"01",X"03",X"07",X"1F",X"9F",X"FF",X"FF",X"1F",X"1F",X"FF",X"FF",X"9F",X"1F",X"07",X"03",X"01",
		X"00",X"00",X"80",X"C0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"C0",X"00",X"00",X"00",
		X"00",X"0F",X"3F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"1F",X"00",
		X"00",X"E0",X"F8",X"F8",X"FC",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FC",X"FC",X"F8",X"E0",X"00",
		X"00",X"01",X"03",X"0F",X"0F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"0F",X"07",X"07",X"01",X"00",
		X"00",X"00",X"C1",X"08",X"80",X"A4",X"00",X"80",X"20",X"00",X"48",X"00",X"81",X"C8",X"00",X"00",
		X"00",X"00",X"00",X"1B",X"37",X"1C",X"4A",X"B0",X"C4",X"69",X"34",X"33",X"0B",X"04",X"00",X"00",
		X"78",X"8E",X"25",X"19",X"1A",X"30",X"00",X"00",X"00",X"00",X"28",X"16",X"06",X"35",X"02",X"58",
		X"04",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"90",X"44",X"88",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"A4",X"40",X"A2",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"01",X"02",X"02",X"02",X"05",X"10",X"04",X"42",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"00",X"00",X"40",X"00",X"00",X"54",X"02",X"4A",X"A6",X"8B",X"F3",X"EE",X"5A",
		X"00",X"08",X"00",X"01",X"10",X"00",X"00",X"09",X"00",X"06",X"03",X"00",X"05",X"00",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"08",X"00",X"A0",X"00",X"00",X"20",X"84",X"00",X"10",X"90",X"48",X"68",X"68",X"A0",X"28",
		X"F0",X"0C",X"82",X"71",X"C1",X"BD",X"41",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"0C",X"13",X"17",X"0E",X"2D",X"5B",X"56",X"4E",X"55",X"19",X"19",X"15",X"0D",X"55",X"59",
		X"F0",X"0C",X"82",X"71",X"C1",X"BD",X"41",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"0C",X"13",X"17",X"2E",X"2D",X"1B",X"16",X"0E",X"15",X"59",X"59",X"55",X"4D",X"15",X"19",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"59",X"55",X"0D",X"15",X"19",X"19",X"55",X"4D",X"4D",X"55",X"19",X"19",X"15",X"0D",X"55",X"59",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"19",X"15",X"4D",X"55",X"59",X"59",X"15",X"0D",X"0D",X"15",X"59",X"59",X"55",X"4D",X"15",X"19",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"42",X"5C",X"60",X"41",X"4E",X"70",X"40",X"40",X"70",X"4E",X"41",X"60",X"5C",X"42",X"01",
		X"00",X"00",X"03",X"0F",X"0E",X"0D",X"03",X"0F",X"0F",X"03",X"0D",X"0E",X"0F",X"03",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"40",X"F0",X"F8",X"F8",X"F8",X"FC",X"FC",X"F8",X"F8",X"F8",X"F0",X"40",X"40",X"00",
		X"0D",X"5A",X"5C",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"5C",X"5A",X"0D",
		X"00",X"00",X"03",X"0F",X"0E",X"0D",X"03",X"0F",X"0F",X"03",X"0D",X"0E",X"0F",X"03",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"44",X"7C",X"40",X"00",X"7C",X"44",X"7C",X"00",X"7C",X"44",X"7C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"48",X"64",X"54",X"48",X"00",X"7C",X"44",X"7C",X"00",X"7C",X"44",X"7C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"30",X"28",X"7C",X"20",X"00",X"7C",X"44",X"7C",X"00",X"7C",X"44",X"7C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"78",X"54",X"54",X"74",X"00",X"7C",X"44",X"7C",X"00",X"7C",X"44",X"7C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"6C",X"54",X"54",X"6C",X"00",X"7C",X"44",X"7C",X"00",X"7C",X"44",X"7C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"01",X"81",X"01",X"02",X"04",X"08",X"10",X"30",X"48",X"88",X"04",X"04",X"04",X"04",
		X"02",X"01",X"01",X"00",X"01",X"02",X"04",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"04",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"18",X"0C",X"05",X"03",X"07",X"07",X"07",X"07",X"03",X"05",X"0C",X"18",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"18",X"0C",X"02",X"04",X"0C",X"1C",X"18",X"18",X"1C",X"0C",X"04",X"02",X"0C",X"18",X"00",
		X"00",X"00",X"00",X"00",X"40",X"E0",X"F0",X"F0",X"F0",X"F0",X"E0",X"40",X"00",X"00",X"00",X"00",
		X"00",X"00",X"06",X"03",X"01",X"00",X"01",X"01",X"01",X"01",X"00",X"01",X"03",X"06",X"00",X"00",
		X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",
		X"00",X"06",X"03",X"00",X"01",X"03",X"07",X"06",X"06",X"07",X"03",X"01",X"00",X"03",X"06",X"00",
		X"00",X"00",X"80",X"04",X"06",X"02",X"82",X"96",X"6E",X"FE",X"92",X"04",X"00",X"50",X"00",X"00",
		X"00",X"82",X"80",X"80",X"80",X"81",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"10",X"0E",
		X"00",X"00",X"50",X"06",X"07",X"03",X"87",X"CF",X"7B",X"D2",X"84",X"00",X"00",X"80",X"00",X"00",
		X"0E",X"10",X"20",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"82",X"00",
		X"00",X"10",X"58",X"08",X"78",X"FC",X"FC",X"FC",X"FC",X"FC",X"7C",X"18",X"30",X"A0",X"60",X"00",
		X"0E",X"10",X"20",X"00",X"00",X"01",X"01",X"00",X"01",X"01",X"80",X"80",X"80",X"80",X"82",X"00",
		X"00",X"60",X"A0",X"30",X"7C",X"FE",X"FE",X"FE",X"FE",X"FE",X"7C",X"18",X"08",X"58",X"10",X"00",
		X"00",X"82",X"80",X"80",X"80",X"81",X"01",X"00",X"01",X"01",X"00",X"00",X"00",X"20",X"10",X"0E",
		X"0A",X"46",X"0F",X"07",X"03",X"80",X"80",X"00",X"80",X"81",X"01",X"01",X"01",X"01",X"00",X"00",
		X"00",X"06",X"05",X"0C",X"7E",X"FF",X"FF",X"FF",X"FF",X"FF",X"7E",X"18",X"10",X"90",X"20",X"80",
		X"00",X"00",X"01",X"01",X"01",X"01",X"81",X"80",X"00",X"80",X"80",X"03",X"07",X"0F",X"46",X"0A",
		X"80",X"20",X"90",X"10",X"18",X"7E",X"FF",X"FF",X"FF",X"FF",X"FF",X"7E",X"0C",X"05",X"06",X"00",
		X"00",X"00",X"08",X"04",X"04",X"2C",X"DC",X"FC",X"24",X"08",X"00",X"A0",X"00",X"00",X"00",X"00",
		X"00",X"80",X"80",X"82",X"03",X"01",X"00",X"01",X"01",X"00",X"00",X"40",X"20",X"1C",X"00",X"00",
		X"00",X"00",X"80",X"CE",X"7B",X"D2",X"84",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"82",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"30",X"7E",X"49",X"02",X"00",X"28",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"08",X"07",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"20",X"00",X"00",X"20",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"20",X"20",X"20",X"20",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"98",X"28",X"0C",X"1E",X"78",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"20",X"20",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"2C",X"04",X"3C",X"FE",X"FE",X"78",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"08",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"60",X"A0",X"30",X"7C",X"FE",X"FE",X"FE",X"FE",X"F8",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"82",X"80",X"80",X"80",X"81",X"01",X"00",X"01",X"01",X"00",X"00",
		X"00",X"00",X"00",X"20",X"B0",X"10",X"F0",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"30",X"40",X"00",
		X"00",X"00",X"1C",X"20",X"40",X"00",X"00",X"03",X"03",X"01",X"03",X"03",X"80",X"80",X"80",X"00",
		X"80",X"B4",X"E0",X"C8",X"D0",X"B1",X"C4",X"80",X"C0",X"80",X"CC",X"78",X"60",X"B0",X"02",X"90",
		X"09",X"AF",X"6B",X"3F",X"CF",X"D4",X"FF",X"F7",X"FB",X"DF",X"BF",X"17",X"F7",X"33",X"4F",X"0B",
		X"01",X"C0",X"E8",X"C0",X"64",X"F0",X"E8",X"E0",X"F0",X"E4",X"E0",X"C2",X"C0",X"14",X"E8",X"81",
		X"87",X"2E",X"4F",X"5F",X"1E",X"2B",X"B7",X"27",X"2F",X"EF",X"DB",X"BC",X"DE",X"8F",X"4F",X"15",
		X"00",X"D0",X"C2",X"60",X"F8",X"FC",X"FC",X"FC",X"FC",X"FC",X"F8",X"30",X"90",X"B0",X"21",X"90",
		X"08",X"A4",X"65",X"D0",X"E8",X"C3",X"F3",X"71",X"33",X"93",X"6A",X"D0",X"F4",X"B0",X"B2",X"10",
		X"C4",X"F0",X"F2",X"F8",X"F8",X"FC",X"FD",X"FC",X"FC",X"FE",X"FE",X"FC",X"F8",X"F9",X"F4",X"C0",
		X"47",X"1F",X"3F",X"3F",X"FF",X"7F",X"7F",X"7F",X"7F",X"FF",X"7F",X"3F",X"3F",X"1F",X"0F",X"27",
		X"90",X"E0",X"F0",X"F0",X"F8",X"FC",X"F8",X"F8",X"F8",X"F8",X"F8",X"F0",X"F8",X"E0",X"F0",X"80",
		X"0F",X"5F",X"3F",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"BF",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E4",X"F8",X"FC",X"FC",X"FE",X"F8",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"17",X"0F",X"3F",X"1F",X"3F",X"3F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E2",X"F8",X"F9",X"FC",X"FC",X"FE",X"F8",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"23",X"0F",X"1F",X"1F",X"7F",X"3F",X"3F",X"3F",X"00",
		X"00",X"00",X"00",X"00",X"90",X"E0",X"F0",X"F0",X"F8",X"FC",X"F8",X"F8",X"F8",X"F8",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"5F",X"3F",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"00",X"00",X"00",X"88",X"E0",X"E4",X"F0",X"F0",X"F8",X"FA",X"F8",X"F8",X"FC",X"F8",X"C0",X"00",
		X"00",X"00",X"00",X"8F",X"3F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"00",
		X"80",X"E8",X"E2",X"B0",X"F8",X"F0",X"FD",X"D8",X"F0",X"E2",X"F8",X"A1",X"F0",X"E4",X"C0",X"88",
		X"0F",X"1F",X"3F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"3F",X"0F",
		X"88",X"E0",X"E4",X"F0",X"A1",X"F8",X"E0",X"74",X"D8",X"FD",X"F0",X"C8",X"F0",X"E2",X"E8",X"80",
		X"0F",X"3F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"3F",X"1F",X"0F",
		X"04",X"30",X"72",X"78",X"78",X"B0",X"C1",X"EC",X"6C",X"8E",X"6E",X"24",X"A0",X"B9",X"B4",X"00",
		X"46",X"13",X"39",X"38",X"13",X"87",X"AD",X"1E",X"6F",X"F7",X"58",X"3D",X"37",X"1F",X"0F",X"27",
		X"00",X"80",X"80",X"10",X"30",X"00",X"00",X"82",X"00",X"10",X"30",X"20",X"80",X"00",X"90",X"00",
		X"02",X"13",X"57",X"3B",X"70",X"81",X"D0",X"B0",X"C8",X"70",X"50",X"A1",X"45",X"0F",X"0B",X"27",
		X"00",X"00",X"00",X"00",X"10",X"00",X"02",X"00",X"00",X"04",X"00",X"40",X"00",X"00",X"20",X"00",
		X"00",X"04",X"22",X"20",X"60",X"04",X"0E",X"B4",X"C0",X"E4",X"A0",X"40",X"14",X"08",X"11",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"20",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"60",X"F0",X"F0",X"F0",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"60",X"F0",X"F0",X"F0",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"0F",X"0F",X"0F",X"06",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"A0",X"A0",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"07",X"07",X"03",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"58",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"BC",X"BC",X"B8",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"78",X"78",X"78",X"30",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"F0",X"F0",X"F0",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"F0",X"F0",X"60",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"60",X"F0",X"F0",X"F0",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"F0",X"F0",X"60",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"78",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"07",X"03",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",X"E0",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"3C",X"3C",X"18",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"40",X"C0",X"E0",X"E0",X"C0",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"40",X"40",X"C0",X"C0",X"40",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"FC",X"FE",X"E1",X"C0",X"80",X"80",X"00",X"80",X"C0",X"E1",X"FE",X"FC",X"E0",X"00",X"00",
		X"3F",X"FF",X"07",X"0F",X"07",X"03",X"C3",X"38",X"03",X"07",X"0F",X"07",X"FF",X"3F",X"00",X"00",
		X"00",X"E0",X"FC",X"E3",X"C0",X"80",X"80",X"00",X"80",X"C0",X"E3",X"FC",X"E0",X"00",X"00",X"00",
		X"00",X"3F",X"FF",X"0F",X"07",X"03",X"33",X"C8",X"03",X"07",X"0F",X"FF",X"3F",X"00",X"00",X"00",
		X"60",X"1C",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"1C",X"E0",X"00",X"00",
		X"3F",X"C0",X"00",X"00",X"00",X"00",X"C0",X"38",X"00",X"00",X"00",X"00",X"C0",X"3F",X"00",X"00",
		X"00",X"E0",X"1C",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"1C",X"60",X"00",X"00",X"00",
		X"00",X"3F",X"C0",X"00",X"00",X"00",X"38",X"C0",X"00",X"00",X"00",X"C0",X"3F",X"00",X"00",X"00",
		X"F8",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"03",X"00",X"00",X"00",X"01",X"5C",X"00",
		X"00",X"0D",X"10",X"20",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"70",X"0F",X"00",
		X"00",X"5C",X"03",X"00",X"00",X"00",X"03",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"F8",
		X"00",X"0F",X"70",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"20",X"10",X"0D",X"00",
		X"00",X"C0",X"80",X"00",X"00",X"00",X"00",X"80",X"C2",X"FC",X"F8",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"1F",X"0F",X"07",X"87",X"70",X"07",X"0F",X"1F",X"0F",X"FF",X"7F",X"00",X"00",X"00",X"00",
		X"00",X"80",X"80",X"00",X"80",X"C0",X"E3",X"FC",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"33",X"C8",X"03",X"07",X"0F",X"FF",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"E0",X"F0",X"FF",X"FE",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"1C",X"01",X"03",X"07",X"03",X"7F",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"F8",X"FE",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"03",X"3F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"07",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"30",X"00",X"00",X"00",X"0E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"0E",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"60",X"00",X"00",X"00",X"00",X"60",X"1C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"1C",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"3F",X"C0",X"00",X"00",X"00",X"38",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"38",X"04",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",
		X"00",X"00",X"7E",X"80",X"00",X"00",X"00",X"00",X"80",X"70",X"00",X"00",X"00",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"E0",X"FC",X"FF",X"00",X"00",X"FF",X"FC",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"3F",X"FF",X"C0",X"38",X"FF",X"3F",X"07",X"00",X"00",X"00",X"00",
		X"00",X"00",X"E0",X"F8",X"1C",X"03",X"00",X"00",X"00",X"03",X"FE",X"FC",X"E0",X"00",X"00",X"00",
		X"00",X"00",X"3F",X"7F",X"C0",X"00",X"00",X"38",X"C0",X"00",X"FF",X"7F",X"1F",X"00",X"00",X"00",
		X"00",X"60",X"1C",X"02",X"01",X"00",X"00",X"00",X"00",X"01",X"02",X"1E",X"FC",X"E0",X"00",X"00",
		X"00",X"3F",X"C0",X"00",X"00",X"00",X"00",X"C0",X"38",X"00",X"00",X"C0",X"7F",X"3F",X"00",X"00",
		X"00",X"00",X"FC",X"F8",X"C6",X"1E",X"3C",X"F8",X"F0",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"07",X"0F",X"1F",X"3C",X"38",X"63",X"4F",X"7F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"E0",X"F0",X"F8",X"3C",X"1E",X"C6",X"F8",X"FC",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"7F",X"4F",X"63",X"38",X"3C",X"1F",X"0F",X"07",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"13",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"FE",X"F1",X"C7",X"0E",X"38",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"0F",X"0E",X"18",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"E0",X"F0",X"F8",X"38",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"4F",X"63",X"38",X"3C",X"1F",X"00",
		X"00",X"00",X"00",X"00",X"F8",X"F0",X"8C",X"3C",X"78",X"F0",X"E0",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"0F",X"1F",X"3E",X"78",X"71",X"C7",X"9F",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"F9",X"C7",X"3E",X"FE",X"FC",X"F8",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"07",X"1F",X"3C",X"70",X"9F",X"1F",X"2F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"C0",X"F8",X"FC",X"FE",X"3E",X"07",X"01",X"C0",X"F8",X"FE",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"2F",X"1F",X"80",X"60",X"30",X"3C",X"1F",X"07",X"01",X"00",X"00",X"00",
		X"40",X"C0",X"C0",X"80",X"0C",X"3C",X"38",X"C0",X"E0",X"C0",X"00",X"80",X"A0",X"70",X"F0",X"78",
		X"00",X"00",X"03",X"05",X"10",X"36",X"78",X"71",X"C7",X"99",X"FC",X"0F",X"07",X"02",X"00",X"00",
		X"C0",X"A0",X"00",X"04",X"08",X"40",X"F0",X"80",X"40",X"30",X"00",X"00",X"C0",X"88",X"20",X"10",
		X"00",X"91",X"25",X"49",X"28",X"60",X"70",X"C2",X"0B",X"B1",X"B0",X"5C",X"0C",X"02",X"40",X"00",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",
		X"00",X"01",X"10",X"40",X"20",X"80",X"80",X"48",X"10",X"45",X"00",X"00",X"40",X"28",X"0C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"0F",X"0F",X"09",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"0F",X"0F",X"09",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"06",X"06",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"06",X"0E",X"0F",X"0F",X"0E",X"06",X"02",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"06",X"06",X"00",X"00",X"00",X"00",X"06",X"06",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"06",X"0E",X"0F",X"0F",X"0E",X"06",X"02",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"D0",X"F0",X"D0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"20",X"00",X"00",X"00",X"01",X"01",X"00",X"10",X"00",X"10",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"D0",X"F0",X"D0",X"80",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"00",X"10",X"00",X"01",X"01",X"00",X"00",X"00",X"20",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"12",X"1E",X"1E",X"12",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"0F",X"0F",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"07",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"00",X"00",X"80",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"07",X"07",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"06",X"0E",X"0F",X"0F",X"0E",X"06",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"0C",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0C",X"1C",X"1E",X"1E",X"1C",X"0C",X"04",X"00",X"00",
		X"00",X"E0",X"50",X"80",X"1C",X"38",X"30",X"70",X"60",X"60",X"00",X"30",X"20",X"00",X"00",X"00",
		X"00",X"08",X"18",X"09",X"03",X"0C",X"08",X"1D",X"34",X"03",X"01",X"00",X"02",X"02",X"00",X"00",
		X"00",X"00",X"30",X"70",X"F2",X"64",X"23",X"19",X"30",X"00",X"B2",X"72",X"06",X"4C",X"98",X"80",
		X"06",X"0D",X"A0",X"00",X"50",X"82",X"D6",X"0E",X"16",X"37",X"53",X"58",X"00",X"08",X"44",X"01",
		X"00",X"00",X"00",X"00",X"0C",X"0C",X"00",X"00",X"00",X"00",X"0C",X"0C",X"00",X"00",X"40",X"00",
		X"22",X"60",X"08",X"40",X"84",X"44",X"1C",X"8E",X"DE",X"5C",X"0C",X"04",X"40",X"60",X"42",X"06",
		X"F0",X"C0",X"E4",X"EC",X"7C",X"38",X"30",X"70",X"E0",X"E0",X"F0",X"30",X"20",X"00",X"00",X"00",
		X"00",X"08",X"1D",X"1F",X"3F",X"0E",X"0C",X"1F",X"37",X"07",X"07",X"03",X"03",X"02",X"00",X"00",
		X"00",X"00",X"00",X"20",X"30",X"F0",X"E0",X"E0",X"70",X"30",X"38",X"7C",X"EC",X"E4",X"C0",X"F0",
		X"00",X"00",X"02",X"03",X"03",X"07",X"07",X"37",X"1F",X"0C",X"0E",X"3F",X"1F",X"1D",X"08",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"24",X"32",X"33",X"7C",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"3C",X"30",X"79",X"FB",X"DF",X"8E",X"0C",X"DC",X"F8",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"07",X"07",X"0F",X"03",X"03",X"07",X"0D",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"98",X"F8",X"F0",X"F0",X"B8",X"18",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"03",X"03",X"1B",X"0F",X"06",X"07",X"00",
		X"00",X"00",X"F0",X"C0",X"E4",X"EC",X"7C",X"38",X"30",X"70",X"E0",X"E0",X"F0",X"30",X"20",X"00",
		X"00",X"00",X"00",X"08",X"1D",X"1F",X"3F",X"0E",X"0C",X"1F",X"37",X"07",X"07",X"03",X"03",X"00",
		X"00",X"00",X"20",X"B8",X"EC",X"C6",X"E0",X"E0",X"E0",X"C0",X"82",X"82",X"C4",X"40",X"E0",X"E0",
		X"00",X"00",X"03",X"03",X"27",X"3D",X"7C",X"7C",X"66",X"67",X"23",X"37",X"1C",X"0C",X"03",X"00",
		X"E0",X"E0",X"40",X"C4",X"82",X"82",X"C0",X"E0",X"E0",X"E0",X"C6",X"EC",X"B8",X"20",X"00",X"00",
		X"00",X"03",X"0C",X"1C",X"37",X"23",X"67",X"66",X"7C",X"7C",X"3D",X"27",X"03",X"03",X"00",X"00",
		X"00",X"00",X"00",X"20",X"20",X"00",X"60",X"E0",X"70",X"30",X"78",X"1C",X"80",X"50",X"E0",X"00",
		X"00",X"00",X"02",X"02",X"00",X"01",X"03",X"35",X"1C",X"0A",X"0C",X"03",X"09",X"18",X"08",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"80",X"00",X"80",X"00",X"00",
		X"10",X"00",X"00",X"11",X"00",X"08",X"1B",X"2F",X"62",X"50",X"01",X"08",X"0C",X"82",X"07",X"20",
		X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"20",X"60",X"12",X"40",X"00",X"40",X"02",X"60",X"00",X"A1",X"30",X"40",X"60",X"08",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C4",X"F0",X"F2",X"F8",X"F8",X"FC",X"FD",X"FC",X"FC",X"FE",X"FE",X"FC",X"F8",X"F9",X"F4",X"C0",
		X"47",X"1F",X"3F",X"3F",X"FF",X"7F",X"7F",X"7F",X"7F",X"FF",X"7F",X"3F",X"3F",X"1F",X"0F",X"27",
		X"C4",X"F0",X"F2",X"F8",X"F8",X"FC",X"FC",X"FC",X"FC",X"FE",X"FE",X"FC",X"F8",X"F8",X"F4",X"C0",
		X"47",X"1F",X"3F",X"3F",X"FF",X"7F",X"7F",X"7F",X"7F",X"FF",X"7F",X"3F",X"3F",X"1F",X"0F",X"27",
		X"C4",X"F0",X"F0",X"F8",X"F8",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"F8",X"F8",X"F4",X"C0",
		X"47",X"1F",X"3F",X"3F",X"FF",X"7F",X"7F",X"7F",X"7F",X"FF",X"7F",X"3F",X"3F",X"1F",X"0F",X"27",
		X"C0",X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F0",X"C0",
		X"47",X"1F",X"3F",X"3F",X"FF",X"7F",X"7F",X"7F",X"7F",X"FF",X"7F",X"3F",X"3F",X"1F",X"0F",X"27",
		X"C0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"C0",
		X"47",X"1F",X"3F",X"3F",X"FF",X"7F",X"7F",X"7F",X"7F",X"FF",X"7F",X"3F",X"3F",X"1F",X"0F",X"27",
		X"C0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"C0",
		X"47",X"1F",X"3F",X"3F",X"FF",X"7F",X"7F",X"7F",X"7F",X"FF",X"7F",X"3F",X"3F",X"1F",X"0F",X"27",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"47",X"1F",X"3F",X"3F",X"FF",X"7F",X"7F",X"7F",X"7F",X"FF",X"7F",X"3F",X"3F",X"1F",X"0F",X"27",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"47",X"1F",X"3F",X"3F",X"FF",X"7F",X"7F",X"7F",X"7F",X"FF",X"7F",X"3F",X"3F",X"1F",X"0F",X"27",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"47",X"1F",X"3F",X"3F",X"FF",X"7F",X"7F",X"7F",X"7F",X"FF",X"7F",X"3F",X"3F",X"1F",X"0F",X"27",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"46",X"1E",X"3E",X"3E",X"FE",X"7E",X"7E",X"7E",X"7E",X"FE",X"7E",X"3E",X"3E",X"1E",X"0E",X"26",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"1C",X"3C",X"3C",X"FC",X"7C",X"7C",X"7C",X"7C",X"FC",X"7C",X"3C",X"3C",X"1C",X"0C",X"24",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"18",X"38",X"38",X"F8",X"78",X"78",X"78",X"78",X"F8",X"78",X"38",X"38",X"18",X"08",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"10",X"30",X"30",X"F0",X"70",X"70",X"70",X"70",X"F0",X"70",X"30",X"30",X"10",X"00",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"00",X"20",X"20",X"E0",X"60",X"60",X"60",X"60",X"E0",X"60",X"20",X"20",X"00",X"00",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"00",X"00",X"00",X"C0",X"40",X"40",X"40",X"40",X"C0",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"F0",X"F0",X"60",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"F0",X"F0",X"60",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"F0",X"F0",X"60",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"F0",X"F0",X"60",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"F0",X"F0",X"60",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"E0",X"E0",X"60",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"C0",X"C0",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FC",X"F8",X"C6",X"1E",X"3C",X"F8",X"F0",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"07",X"0F",X"1F",X"3C",X"38",X"63",X"4F",X"7F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FC",X"F8",X"C6",X"1E",X"3C",X"F8",X"F0",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"07",X"0F",X"1F",X"3C",X"38",X"63",X"4F",X"7F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FC",X"F8",X"C4",X"1C",X"3C",X"F8",X"F0",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"07",X"0F",X"1F",X"3C",X"38",X"63",X"4F",X"7F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"F8",X"F8",X"C0",X"18",X"38",X"F8",X"F0",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"07",X"0F",X"1F",X"3C",X"38",X"63",X"4F",X"7F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"F0",X"F0",X"C0",X"10",X"30",X"F0",X"F0",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"07",X"0F",X"1F",X"3C",X"38",X"63",X"4F",X"7F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"E0",X"E0",X"C0",X"00",X"20",X"E0",X"E0",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"07",X"0F",X"1F",X"3C",X"38",X"63",X"4F",X"7F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"C0",X"C0",X"00",X"00",X"C0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"07",X"0F",X"1F",X"3C",X"38",X"63",X"4F",X"7F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"80",X"80",X"00",X"00",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"07",X"0F",X"1F",X"3C",X"38",X"63",X"4F",X"7F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"07",X"0F",X"1F",X"3C",X"38",X"63",X"4F",X"7F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"06",X"0E",X"1E",X"3C",X"38",X"62",X"4E",X"7E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"04",X"0C",X"1C",X"3C",X"38",X"60",X"4C",X"7C",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"18",X"38",X"38",X"60",X"48",X"78",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"30",X"60",X"40",X"70",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"60",X"40",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"C0",X"E4",X"EC",X"7C",X"38",X"30",X"70",X"E0",X"E0",X"F0",X"30",X"20",X"00",X"00",X"00",
		X"00",X"08",X"1D",X"1F",X"3F",X"0E",X"0C",X"1F",X"37",X"07",X"07",X"03",X"03",X"02",X"00",X"00",
		X"F0",X"C0",X"E4",X"EC",X"7C",X"38",X"30",X"70",X"E0",X"E0",X"F0",X"30",X"20",X"00",X"00",X"00",
		X"00",X"08",X"1D",X"1F",X"3F",X"0E",X"0C",X"1F",X"37",X"07",X"07",X"03",X"03",X"02",X"00",X"00",
		X"F0",X"C0",X"E4",X"EC",X"7C",X"38",X"30",X"70",X"E0",X"E0",X"F0",X"30",X"20",X"00",X"00",X"00",
		X"00",X"08",X"1D",X"1F",X"3F",X"0E",X"0C",X"1F",X"37",X"07",X"07",X"03",X"03",X"02",X"00",X"00",
		X"F0",X"C0",X"E0",X"E8",X"78",X"38",X"30",X"70",X"E0",X"E0",X"F0",X"30",X"20",X"00",X"00",X"00",
		X"00",X"08",X"1D",X"1F",X"3F",X"0E",X"0C",X"1F",X"37",X"07",X"07",X"03",X"03",X"02",X"00",X"00",
		X"F0",X"C0",X"E0",X"E0",X"70",X"30",X"30",X"70",X"E0",X"E0",X"F0",X"30",X"20",X"00",X"00",X"00",
		X"00",X"08",X"1D",X"1F",X"3F",X"0E",X"0C",X"1F",X"37",X"07",X"07",X"03",X"03",X"02",X"00",X"00",
		X"E0",X"C0",X"E0",X"E0",X"60",X"20",X"20",X"60",X"E0",X"E0",X"E0",X"20",X"20",X"00",X"00",X"00",
		X"00",X"08",X"1D",X"1F",X"3F",X"0E",X"0C",X"1F",X"37",X"07",X"07",X"03",X"03",X"02",X"00",X"00",
		X"C0",X"C0",X"C0",X"C0",X"40",X"00",X"00",X"40",X"C0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"1D",X"1F",X"3F",X"0E",X"0C",X"1F",X"37",X"07",X"07",X"03",X"03",X"02",X"00",X"00",
		X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"1D",X"1F",X"3F",X"0E",X"0C",X"1F",X"37",X"07",X"07",X"03",X"03",X"02",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"1D",X"1F",X"3F",X"0E",X"0C",X"1F",X"37",X"07",X"07",X"03",X"03",X"02",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"1C",X"1E",X"3E",X"0E",X"0C",X"1E",X"36",X"06",X"06",X"02",X"02",X"02",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"1C",X"1C",X"3C",X"0C",X"0C",X"1C",X"34",X"04",X"04",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"18",X"18",X"38",X"08",X"08",X"18",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"10",X"30",X"00",X"00",X"10",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
