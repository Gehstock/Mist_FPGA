library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_OBJ_1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_OBJ_1 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"38",X"7C",X"C2",X"82",X"86",X"7C",X"38",X"00",X"02",X"02",X"FE",X"FE",X"42",X"02",X"00",X"00",
		X"62",X"F2",X"BA",X"9A",X"9E",X"CE",X"46",X"00",X"8C",X"DE",X"F2",X"B2",X"92",X"86",X"04",X"00",
		X"08",X"FE",X"FE",X"C8",X"68",X"38",X"18",X"00",X"1C",X"BE",X"A2",X"A2",X"A2",X"E6",X"E4",X"00",
		X"0C",X"9E",X"92",X"92",X"D2",X"7E",X"3C",X"00",X"C0",X"E0",X"B0",X"9E",X"8E",X"C0",X"C0",X"00",
		X"0C",X"6E",X"9A",X"9A",X"B2",X"F2",X"6C",X"00",X"78",X"FC",X"96",X"92",X"92",X"F2",X"60",X"00",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"3C",X"42",X"81",X"A5",X"A5",X"99",X"42",X"3C",
		X"00",X"00",X"00",X"06",X"06",X"00",X"00",X"00",X"00",X"70",X"F8",X"8D",X"85",X"C0",X"60",X"00",
		X"8E",X"4A",X"2E",X"10",X"E8",X"A4",X"E2",X"00",X"18",X"3C",X"7E",X"FF",X"3C",X"3C",X"3C",X"3C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"7E",X"C8",X"88",X"C8",X"7E",X"3E",X"00",
		X"6C",X"FE",X"92",X"92",X"92",X"FE",X"FE",X"00",X"44",X"C6",X"82",X"82",X"C6",X"7C",X"38",X"00",
		X"38",X"7C",X"C6",X"82",X"82",X"FE",X"FE",X"00",X"82",X"92",X"92",X"92",X"FE",X"FE",X"00",X"00",
		X"80",X"90",X"90",X"90",X"90",X"FE",X"FE",X"00",X"9E",X"9E",X"92",X"82",X"C6",X"7C",X"38",X"00",
		X"FE",X"FE",X"10",X"10",X"10",X"FE",X"FE",X"00",X"82",X"82",X"FE",X"FE",X"82",X"82",X"00",X"00",
		X"FC",X"FE",X"02",X"02",X"02",X"06",X"04",X"00",X"82",X"C6",X"6E",X"3C",X"18",X"FE",X"FE",X"00",
		X"02",X"02",X"02",X"02",X"FE",X"FE",X"00",X"00",X"FE",X"FE",X"70",X"38",X"70",X"FE",X"FE",X"00",
		X"FE",X"FE",X"1C",X"38",X"70",X"FE",X"FE",X"00",X"7C",X"FE",X"82",X"82",X"82",X"FE",X"7C",X"00",
		X"70",X"F8",X"88",X"88",X"88",X"FE",X"FE",X"00",X"7A",X"FC",X"8E",X"8A",X"82",X"FE",X"7C",X"00",
		X"72",X"F6",X"9E",X"8C",X"88",X"FE",X"FE",X"00",X"0C",X"5E",X"D2",X"92",X"92",X"F6",X"64",X"00",
		X"80",X"80",X"FE",X"FE",X"80",X"80",X"00",X"00",X"FC",X"FE",X"02",X"02",X"02",X"FE",X"FC",X"00",
		X"F0",X"F8",X"1C",X"0E",X"1C",X"F8",X"F0",X"00",X"F8",X"FE",X"1C",X"38",X"1C",X"FE",X"F8",X"00",
		X"C6",X"EE",X"7C",X"38",X"7C",X"EE",X"C6",X"00",X"C0",X"F0",X"1E",X"1E",X"F0",X"C0",X"00",X"00",
		X"C2",X"E2",X"F2",X"BA",X"9E",X"8E",X"86",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",
		X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"08",X"02",X"07",X"00",X"00",X"00",X"00",X"00",X"20",X"80",X"C0",
		X"02",X"07",X"02",X"08",X"00",X"00",X"00",X"00",X"80",X"C0",X"80",X"20",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"00",X"02",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"C0",
		X"02",X"07",X"12",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"80",X"00",X"40",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"00",X"02",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"D0",
		X"02",X"17",X"02",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"80",X"00",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"02",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",
		X"12",X"07",X"02",X"00",X"01",X"00",X"00",X"00",X"90",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",
		X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"60",X"80",
		X"01",X"06",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"38",X"10",X"20",X"C4",X"4F",
		X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"20",X"10",X"38",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"03",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"F8",
		X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"C8",X"5C",X"CE",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"05",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",
		X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"7C",X"C0",X"90",X"B8",X"98",X"84",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"05",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"01",X"01",X"01",X"03",X"03",X"00",X"00",X"00",X"58",X"78",X"80",X"20",X"30",X"20",X"10",X"00",
		X"00",X"00",X"00",X"00",X"02",X"02",X"02",X"02",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",
		X"02",X"03",X"14",X"18",X"13",X"01",X"01",X"00",X"80",X"80",X"50",X"30",X"90",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"38",X"10",X"20",X"C8",X"4E",
		X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C8",X"20",X"10",X"38",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"03",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"F8",
		X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"C8",X"5C",X"C8",X"C6",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"05",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",
		X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"7C",X"C0",X"90",X"B8",X"98",X"84",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"05",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"01",X"01",X"01",X"03",X"03",X"00",X"00",X"00",X"58",X"78",X"80",X"20",X"30",X"20",X"10",X"00",
		X"00",X"00",X"00",X"00",X"02",X"02",X"02",X"02",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",
		X"02",X"03",X"14",X"18",X"13",X"03",X"01",X"01",X"80",X"80",X"50",X"30",X"10",X"80",X"00",X"00",
		X"03",X"03",X"07",X"07",X"03",X"03",X"07",X"0F",X"80",X"80",X"C0",X"C0",X"80",X"80",X"C0",X"E0",
		X"AF",X"5F",X"AF",X"5F",X"0F",X"0F",X"08",X"1C",X"F4",X"EA",X"F4",X"EA",X"E0",X"E0",X"10",X"38",
		X"00",X"00",X"00",X"00",X"06",X"0F",X"19",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"EC",
		X"18",X"18",X"0E",X"06",X"00",X"00",X"00",X"00",X"6C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"60",X"60",X"80",
		X"01",X"06",X"06",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"F8",X"F0",X"E0",X"C0",X"C1",X"C0",X"FF",X"FF",X"3F",X"0F",X"03",X"63",X"E1",X"E1",
		X"C2",X"E7",X"E3",X"E0",X"F0",X"F8",X"FE",X"FF",X"61",X"21",X"81",X"01",X"03",X"03",X"0F",X"FF",
		X"FF",X"C1",X"80",X"8E",X"10",X"20",X"07",X"0F",X"FF",X"E7",X"5B",X"1B",X"A7",X"1F",X"1B",X"95",
		X"93",X"80",X"80",X"C0",X"C1",X"E0",X"F0",X"FF",X"CB",X"CF",X"CF",X"8F",X"1F",X"3F",X"7F",X"FF",
		X"DF",X"F8",X"76",X"EE",X"EE",X"EF",X"F7",X"F8",X"87",X"03",X"01",X"01",X"11",X"01",X"03",X"87",
		X"8F",X"07",X"03",X"03",X"83",X"83",X"C7",X"FF",X"FF",X"FF",X"FB",X"F0",X"F9",X"FF",X"7F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"F7",X"E3",X"F7",X"FF",X"E3",X"C5",X"9E",X"96",X"BA",X"DC",X"E1",X"F3",
		X"FF",X"FF",X"CF",X"97",X"B3",X"C7",X"CF",X"FF",X"FF",X"FF",X"C7",X"BB",X"AB",X"BB",X"C7",X"FD",
		X"FF",X"E3",X"C5",X"9E",X"9E",X"BE",X"DC",X"E1",X"FF",X"FF",X"F1",X"E2",X"E6",X"EE",X"F0",X"FD",
		X"FF",X"FF",X"FF",X"CE",X"B6",X"B6",X"CF",X"FF",X"FF",X"8F",X"77",X"FB",X"FB",X"FB",X"77",X"8F",
		X"FF",X"FB",X"F5",X"FB",X"C7",X"83",X"3D",X"3C",X"FF",X"FF",X"FF",X"C7",X"8B",X"3D",X"2D",X"74",
		X"7C",X"B9",X"C3",X"8B",X"9B",X"B9",X"C1",X"E3",X"B9",X"C3",X"F7",X"F3",X"ED",X"ED",X"F3",X"FF",
		X"FF",X"FF",X"FB",X"F1",X"FB",X"DF",X"FF",X"FF",X"FD",X"FA",X"FD",X"FF",X"DF",X"AF",X"DF",X"FF",
		X"FF",X"FF",X"FF",X"F9",X"F6",X"F6",X"F9",X"FF",X"FF",X"F7",X"E3",X"F3",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"F7",X"EB",X"F7",X"FF",X"C7",X"83",X"FF",X"9F",X"0F",X"07",X"87",X"CF",X"C7",X"83",
		X"99",X"99",X"C1",X"E3",X"FF",X"FF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"07",X"0F",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"06",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"03",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"04",X"01",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",
		X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"20",X"60",X"E0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"60",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"01",X"03",X"02",X"02",X"02",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",
		X"01",X"03",X"0B",X"0B",X"0B",X"1B",X"1B",X"16",X"00",X"80",X"A0",X"A0",X"A0",X"B0",X"B0",X"D0",
		X"00",X"00",X"01",X"01",X"03",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",
		X"0B",X"0D",X"08",X"00",X"00",X"00",X"00",X"00",X"A0",X"60",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"1F",X"00",X"00",X"00",X"00",X"A0",X"40",X"A0",X"00",
		X"03",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"01",X"03",X"02",X"02",X"02",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",
		X"01",X"03",X"0B",X"0A",X"08",X"18",X"10",X"00",X"00",X"80",X"A0",X"A0",X"20",X"30",X"10",X"00",
		X"00",X"00",X"01",X"01",X"03",X"02",X"02",X"02",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",
		X"00",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"18",X"20",X"40",X"40",X"80",X"81",X"FF",X"E0",X"98",X"84",X"82",X"82",X"81",X"81",X"C1",
		X"83",X"81",X"81",X"41",X"41",X"21",X"19",X"07",X"FF",X"81",X"01",X"02",X"02",X"04",X"18",X"E0",
		X"07",X"1C",X"24",X"44",X"42",X"82",X"83",X"83",X"E0",X"18",X"04",X"02",X"02",X"0F",X"F1",X"C1",
		X"83",X"8F",X"F0",X"40",X"40",X"20",X"18",X"07",X"C1",X"C1",X"41",X"42",X"22",X"24",X"38",X"E0",
		X"07",X"18",X"20",X"50",X"48",X"84",X"83",X"83",X"E0",X"18",X"04",X"0A",X"12",X"21",X"C1",X"C1",
		X"83",X"83",X"84",X"48",X"50",X"20",X"18",X"07",X"C1",X"41",X"21",X"12",X"0A",X"04",X"18",X"E0",
		X"00",X"00",X"00",X"02",X"00",X"84",X"10",X"00",X"00",X"40",X"04",X"00",X"00",X"50",X"00",X"22",
		X"8A",X"00",X"00",X"00",X"04",X"00",X"20",X"04",X"00",X"80",X"10",X"00",X"14",X"80",X"20",X"00",
		X"00",X"00",X"08",X"04",X"00",X"01",X"23",X"01",X"00",X"00",X"41",X"02",X"08",X"C0",X"B2",X"68",
		X"86",X"13",X"20",X"07",X"03",X"00",X"10",X"00",X"48",X"D4",X"B0",X"64",X"C0",X"08",X"01",X"10",
		X"00",X"00",X"00",X"00",X"0C",X"14",X"05",X"28",X"00",X"00",X"00",X"00",X"80",X"00",X"40",X"40",
		X"21",X"06",X"33",X"01",X"0B",X"04",X"00",X"00",X"40",X"00",X"00",X"40",X"00",X"00",X"00",X"00",
		X"07",X"18",X"23",X"4C",X"50",X"90",X"A1",X"A2",X"E0",X"18",X"C4",X"32",X"0A",X"09",X"85",X"45",
		X"A2",X"A1",X"90",X"50",X"4C",X"23",X"18",X"07",X"45",X"85",X"09",X"0A",X"32",X"C4",X"18",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"38",X"10",X"20",X"C0",X"40",
		X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"20",X"10",X"38",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"03",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"F8",
		X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"C0",X"40",X"C0",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"05",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",
		X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"7C",X"C0",X"80",X"80",X"80",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"05",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"01",X"01",X"01",X"03",X"03",X"00",X"00",X"00",X"58",X"78",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"02",X"02",X"02",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",
		X"02",X"03",X"14",X"18",X"10",X"00",X"00",X"00",X"80",X"80",X"50",X"30",X"10",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
