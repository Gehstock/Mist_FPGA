library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity bg2_rom is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of bg2_rom is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"0F",X"1E",X"3C",X"78",X"F0",X"E1",X"C3",X"87",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F0",X"E1",X"C3",X"87",X"0F",X"1E",X"3C",X"78",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"38",X"6C",X"C6",X"83",X"83",X"C6",X"6C",X"38",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3C",X"3C",X"78",X"F0",X"F0",X"F0",X"78",X"3C",X"C3",X"C3",X"87",X"0F",X"0F",X"0F",X"87",X"C3",
		X"3C",X"3C",X"78",X"F0",X"F0",X"F0",X"78",X"3C",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"F8",X"88",X"F8",X"00",X"F8",X"88",X"F8",
		X"00",X"48",X"F8",X"08",X"00",X"F8",X"88",X"F8",X"00",X"48",X"F8",X"08",X"00",X"E8",X"A8",X"B8",
		X"00",X"B8",X"A8",X"E8",X"00",X"F8",X"88",X"F8",X"00",X"B8",X"A8",X"E8",X"00",X"E8",X"A8",X"B8",
		X"00",X"88",X"A8",X"F8",X"00",X"F8",X"88",X"F8",X"00",X"88",X"A8",X"F8",X"00",X"E8",X"A8",X"B8",
		X"00",X"F0",X"10",X"F8",X"00",X"F8",X"88",X"F8",X"00",X"F0",X"10",X"F8",X"00",X"E8",X"A8",X"B8",
		X"00",X"E8",X"A8",X"B8",X"00",X"F8",X"88",X"F8",X"00",X"F8",X"A8",X"B8",X"00",X"F8",X"88",X"F8",
		X"00",X"80",X"80",X"F8",X"00",X"F8",X"88",X"F8",X"00",X"F8",X"A8",X"F8",X"00",X"F8",X"88",X"F8",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"FE",X"FE",X"FE",X"FC",X"FC",X"FC",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FC",X"FC",X"FC",X"F8",X"F8",X"F8",X"F8",X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"E0",X"E0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"E0",X"E0",X"E0",X"F0",X"F0",X"F0",X"F8",X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F8",X"FC",X"FC",X"FC",X"FE",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"FE",X"FC",X"FC",X"F8",X"F8",X"F8",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F0",X"E0",X"E0",X"F0",X"F8",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FC",X"F8",X"F8",X"F0",X"F0",X"E0",X"C0",X"C0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"C0",X"80",X"80",X"80",X"80",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FE",X"FC",X"FC",X"F8",X"F8",X"F8",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"E0",X"E0",X"E0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"F0",X"F8",X"FC",X"FC",X"FC",X"FC",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"C0",X"E0",X"E0",X"E0",X"F0",X"F0",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"C3",X"FF",X"FF",X"C7",X"03",X"00",X"00",X"60",X"A0",X"A3",X"FF",X"FF",X"F0",
		X"3C",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"80",X"80",X"80",X"00",X"80",X"C0",X"80",X"FF",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"E0",X"FF",X"FF",X"7F",X"00",X"00",X"00",X"00",X"C7",X"9F",X"7F",X"FC",X"C8",X"98",X"D0",X"DC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E6",X"E0",X"C0",X"80",X"C0",X"80",X"C0",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"C7",X"03",
		X"FF",X"7F",X"3F",X"7F",X"1F",X"3F",X"0F",X"9F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"7F",X"3F",X"BF",X"FF",X"FF",X"FF",X"01",X"00",X"00",X"08",X"0F",X"1F",X"07",X"01",
		X"FF",X"FF",X"3F",X"0F",X"1F",X"1F",X"1F",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"E0",X"F0",X"F0",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",X"F0",X"F8",X"FC",X"FC",
		X"00",X"FE",X"FF",X"7F",X"27",X"23",X"01",X"01",X"00",X"0F",X"38",X"F0",X"F0",X"F0",X"F8",X"F8",
		X"F8",X"F8",X"F8",X"F9",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"03",X"0F",X"01",X"00",X"00",X"00",X"01",X"63",
		X"F0",X"F0",X"C0",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"F8",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"01",X"07",X"FF",X"FF",X"FF",X"F9",X"F0",
		X"9C",X"0E",X"0F",X"9F",X"FF",X"FF",X"F9",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F3",X"E0",X"E0",X"E0",X"60",X"60",X"E0",X"F0",X"FF",X"FF",X"F9",X"F0",X"E0",X"E0",X"F0",X"F9",
		X"70",X"79",X"FF",X"FF",X"FF",X"FF",X"FF",X"F3",X"E0",X"E0",X"F0",X"F9",X"FF",X"07",X"03",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F8",X"FC",X"FC",X"F8",X"F8",X"F0",X"E0",
		X"FF",X"FF",X"FF",X"E3",X"C1",X"C1",X"C1",X"E3",X"E1",X"E1",X"73",X"7F",X"7F",X"7F",X"FF",X"E7",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FE",X"F8",X"00",X"00",X"00",X"00",
		X"C3",X"C3",X"E7",X"FF",X"FF",X"00",X"00",X"00",X"03",X"07",X"0F",X"1F",X"1F",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FF",X"FF",X"FF",X"9F",X"1F",X"13",X"33",X"00",X"03",X"0F",X"1F",X"3F",X"7E",X"FC",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"FF",X"FF",X"FF",X"F3",X"73",X"3F",X"1F",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"F8",X"F8",X"03",X"03",X"07",X"07",X"0F",X"0F",X"1F",X"1F",
		X"0F",X"1F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"1F",X"3F",X"3F",X"3F",X"7F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"3F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"E0",X"C0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",
		X"3F",X"1F",X"0F",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"FF",X"00",X"00",X"00",X"00",X"80",X"FC",X"FF",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"F8",X"F0",X"E0",X"E0",X"C0",X"80",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"F0",X"E0",X"80",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"E0",X"E0",X"E0",X"E0",X"F0",X"F8",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"80",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"82",X"C2",X"C7",X"C7",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"C0",X"E7",X"E3",X"F3",X"F1",X"F9",X"F9",X"FC",X"7C",
		X"C3",X"47",X"6E",X"B8",X"4F",X"FF",X"DF",X"D9",X"3C",X"1C",X"0E",X"07",X"00",X"71",X"FB",X"FF",
		X"00",X"80",X"C0",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"F8",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"F0",X"00",X"80",X"C0",X"F0",X"FC",X"FE",X"FF",X"FF",
		X"C0",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"0F",X"00",X"00",X"00",X"C0",X"FF",X"FF",
		X"FF",X"FC",X"FC",X"F8",X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"00",X"C0",X"FF",X"FF",
		X"FF",X"3F",X"00",X"00",X"00",X"3F",X"00",X"3F",X"FF",X"FC",X"F0",X"F8",X"F0",X"F8",X"FC",X"FE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"C0",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"F8",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FE",X"FC",X"FC",X"FC",X"78",X"30",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"1E",X"00",X"7F",X"FF",X"23",X"01",X"00",X"00",X"00",X"00",
		X"1F",X"0F",X"3F",X"1F",X"FF",X"7F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"8F",X"0F",X"07",X"0F",X"0F",X"0F",X"07",X"03",X"01",X"00",
		X"07",X"01",X"0F",X"3F",X"3F",X"1F",X"0B",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"F0",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"F8",X"F8",
		X"00",X"06",X"06",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"BF",X"3F",X"73",X"F3",X"00",X"03",X"0F",X"1F",X"3F",X"77",X"F2",X"FA",
		X"FF",X"FF",X"FF",X"F3",X"F3",X"FF",X"7F",X"7F",X"F8",X"FD",X"FD",X"FD",X"FC",X"F8",X"FA",X"FB",
		X"3F",X"9F",X"CF",X"EF",X"EF",X"FF",X"FF",X"FF",X"FB",X"F3",X"F7",X"F7",X"F7",X"F7",X"F7",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"07",X"0F",X"1F",X"1F",X"1F",X"1F",X"0F",X"8F",
		X"CF",X"DF",X"7F",X"7F",X"7F",X"7F",X"7F",X"40",X"40",X"78",X"78",X"78",X"78",X"78",X"F8",X"F8",
		X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"78",X"38",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"E0",X"60",X"30",X"98",X"CC",X"CC",X"00",X"00",X"02",X"02",X"03",X"07",X"0F",X"1F",
		X"98",X"B8",X"30",X"70",X"60",X"E0",X"00",X"00",X"0F",X"07",X"03",X"03",X"02",X"02",X"00",X"00",
		X"00",X"00",X"C0",X"E0",X"E0",X"00",X"FC",X"FE",X"00",X"00",X"0F",X"1F",X"1F",X"1E",X"1C",X"1D",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FC",X"00",X"00",X"1D",X"0D",X"01",X"01",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"E0",X"F0",X"F8",X"F0",X"E0",X"00",X"00",X"00",X"00",X"07",X"0F",X"1F",X"1F",
		X"E0",X"F0",X"F8",X"F0",X"E0",X"00",X"00",X"00",X"1F",X"1F",X"0F",X"07",X"00",X"00",X"00",X"00",
		X"00",X"00",X"40",X"60",X"30",X"32",X"36",X"7E",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"1C",
		X"FE",X"F6",X"B2",X"30",X"60",X"40",X"00",X"00",X"1C",X"09",X"03",X"07",X"0E",X"0C",X"00",X"00",
		X"00",X"00",X"00",X"98",X"AC",X"D6",X"D6",X"D6",X"00",X"00",X"00",X"07",X"0F",X"1F",X"1F",X"1F",
		X"D6",X"D6",X"D6",X"AC",X"98",X"00",X"00",X"00",X"1F",X"1F",X"1F",X"0F",X"07",X"00",X"00",X"00",
		X"00",X"00",X"F8",X"FC",X"FE",X"FE",X"FE",X"FE",X"00",X"00",X"01",X"03",X"07",X"07",X"0F",X"1F",
		X"FE",X"FE",X"FE",X"FE",X"FC",X"F8",X"00",X"00",X"1F",X"0F",X"07",X"07",X"03",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"1F",X"1F",X"1F",X"1F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"1F",X"1F",X"1F",X"1F",X"1F",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FE",X"FE",X"FE",X"7E",X"00",X"00",X"00",X"07",X"03",X"01",X"00",X"1E",
		X"3E",X"9E",X"C0",X"E0",X"F0",X"00",X"00",X"00",X"1F",X"1F",X"1F",X"1F",X"1F",X"00",X"00",X"00",
		X"00",X"C2",X"DE",X"E2",X"DE",X"E2",X"FE",X"42",X"00",X"44",X"6F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"FE",X"02",X"FE",X"02",X"E6",X"DA",X"DA",X"00",X"7F",X"7F",X"7F",X"7F",X"7F",X"6F",X"44",X"00",
		X"00",X"00",X"F0",X"F8",X"FC",X"FE",X"FE",X"FE",X"00",X"00",X"03",X"07",X"07",X"0F",X"1F",X"1F",
		X"FE",X"FC",X"FC",X"F0",X"E0",X"C0",X"00",X"00",X"1F",X"1F",X"1F",X"0F",X"0F",X"07",X"00",X"00",
		X"00",X"00",X"00",X"F0",X"F8",X"FC",X"FC",X"FC",X"00",X"00",X"00",X"07",X"0F",X"1F",X"1F",X"1F",
		X"FC",X"FC",X"FC",X"F8",X"F0",X"00",X"00",X"00",X"1F",X"1F",X"1F",X"0F",X"07",X"00",X"00",X"00",
		X"00",X"00",X"00",X"E0",X"31",X"19",X"0F",X"19",X"00",X"00",X"00",X"07",X"04",X"04",X"04",X"1C",
		X"31",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"34",X"27",X"21",X"33",X"1E",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"60",X"60",X"60",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"60",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"9E",X"9E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E7",X"E7",X"00",X"00",X"00",X"00",X"00",X"00",X"79",X"79",X"00",
		X"00",X"00",X"00",X"00",X"00",X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"06",
		X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"06",X"00",X"60",X"60",X"60",X"60",X"60",X"60",X"60",
		X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"00",
		X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"06",
		X"00",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"60",X"00",X"00",X"60",X"60",X"60",X"60",X"00",
		X"60",X"60",X"60",X"00",X"00",X"60",X"60",X"60",X"00",X"60",X"60",X"60",X"60",X"00",X"00",X"60",
		X"00",X"06",X"06",X"06",X"06",X"00",X"00",X"06",X"06",X"06",X"06",X"00",X"00",X"06",X"06",X"06",
		X"06",X"00",X"00",X"06",X"06",X"06",X"06",X"00",X"00",X"E0",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"60",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"60",X"60",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"79",X"79",X"00",X"00",X"00",X"00",X"00",X"00",X"E7",X"E7",X"00",X"00",X"00",X"00",X"00",
		X"00",X"9E",X"9E",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"06",X"00",X"00",X"00",X"00",X"00",
		X"06",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"07",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"F0",X"F8",X"FC",X"FE",X"FF",
		X"01",X"03",X"07",X"0F",X"1F",X"3F",X"7F",X"FF",X"80",X"C0",X"E0",X"F0",X"F8",X"FC",X"0E",X"00",
		X"FF",X"FF",X"FF",X"FF",X"0F",X"00",X"00",X"00",X"FF",X"3F",X"0F",X"03",X"03",X"0F",X"3F",X"FF",
		X"00",X"0E",X"FC",X"F8",X"F0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"0F",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FC",X"F0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FE",X"FC",X"F8",X"F0",X"E0",X"C0",X"80",X"C0",X"70",X"3C",X"1F",X"0F",X"07",X"03",X"01",
		X"00",X"00",X"00",X"00",X"00",X"03",X"0F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FC",X"F0",X"C0",X"00",
		X"00",X"C0",X"F0",X"FC",X"FF",X"FF",X"FF",X"FF",X"3F",X"0F",X"03",X"00",X"00",X"00",X"00",X"00",
		X"01",X"03",X"07",X"0F",X"1F",X"3C",X"70",X"C0",X"00",X"C0",X"F0",X"FC",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"3F",X"0F",X"03",X"03",X"0F",X"3F",X"FF",X"FF",X"7F",X"3F",X"1F",X"0F",X"07",X"03",X"01",
		X"00",X"00",X"00",X"00",X"1C",X"3C",X"7F",X"FF",X"00",X"00",X"00",X"00",X"00",X"0C",X"0E",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"70",X"F0",X"78",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"F0",X"F8",X"FC",X"FE",X"FF",X"F0",X"E0",X"01",X"00",X"00",X"00",X"00",X"81",X"C3",X"FF",
		X"00",X"00",X"01",X"03",X"03",X"07",X"07",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FC",X"FF",X"FF",X"FE",X"F0",X"38",X"18",X"39",X"F0",X"F0",X"F0",X"F9",X"FF",X"FF",X"FE",
		X"7C",X"3F",X"1F",X"FF",X"FF",X"7F",X"1F",X"7F",X"00",X"00",X"00",X"0F",X"3E",X"FC",X"F0",X"FC",
		X"02",X"03",X"06",X"0C",X"1E",X"FF",X"FF",X"FF",X"30",X"30",X"38",X"3C",X"7E",X"FF",X"FF",X"FF",
		X"C0",X"C0",X"C0",X"C0",X"E0",X"B0",X"3F",X"3F",X"FF",X"FF",X"FF",X"FF",X"0F",X"07",X"03",X"02",
		X"0F",X"1F",X"7F",X"FF",X"9F",X"1E",X"3C",X"FC",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"F8",X"F8",X"F8",X"F8",X"F0",X"E0",X"80",
		X"FF",X"FF",X"FF",X"7F",X"1F",X"7F",X"FF",X"FF",X"FE",X"FF",X"FE",X"FC",X"F0",X"FC",X"FE",X"EF",
		X"FF",X"FF",X"7F",X"3F",X"1F",X"1F",X"0F",X"0F",X"FF",X"E1",X"80",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"7F",X"FF",X"FF",X"FE",X"FE",X"FC",X"7C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FF",X"EE",X"CC",X"00",X"00",X"00",X"00",X"1F",X"1F",X"3F",X"3F",X"1F",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"C0",X"C0",X"C0",X"60",X"60",X"00",X"00",X"40",
		X"0F",X"0F",X"18",X"10",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"E0",X"FC",
		X"7C",X"3C",X"3E",X"1E",X"3F",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"EF",X"FF",X"FF",X"87",X"03",X"01",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"F8",X"F8",X"F8",X"F8",X"88",X"00",X"00",
		X"01",X"01",X"01",X"03",X"87",X"FF",X"FF",X"FE",X"00",X"00",X"00",X"01",X"03",X"03",X"03",X"03",
		X"80",X"C0",X"C0",X"C0",X"FC",X"FC",X"F8",X"C0",X"01",X"03",X"07",X"1F",X"1F",X"1F",X"1F",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"00",X"00",X"00",X"80",X"FE",X"E7",X"E1",X"E1",
		X"1E",X"0E",X"07",X"07",X"07",X"07",X"0F",X"1F",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"E0",X"60",X"00",X"00",X"00",X"00",X"00",X"3F",X"3F",X"3F",X"1B",X"00",X"00",X"00",X"00",
		X"F0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"7E",X"00",X"00",X"00",X"00",
		X"1F",X"3F",X"3F",X"3F",X"3E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"38",X"78",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"00",X"00",X"C0",X"F0",X"FC",X"FE",X"0F",X"03",
		X"00",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"1E",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F8",X"F8",X"78",X"78",X"78",X"78",X"78",X"40",X"01",X"00",X"00",X"FE",X"FE",X"B6",X"B6",X"B6",
		X"0E",X"0E",X"1C",X"3D",X"F9",X"F1",X"E1",X"F1",X"7E",X"7C",X"7C",X"3E",X"3F",X"3F",X"1F",X"0F",
		X"40",X"7F",X"7F",X"7F",X"7F",X"7F",X"DF",X"CF",X"B6",X"B6",X"B6",X"86",X"86",X"00",X"00",X"01",
		X"F1",X"E1",X"F1",X"F9",X"3D",X"1C",X"0E",X"0E",X"0F",X"1F",X"3F",X"3F",X"3E",X"7C",X"7C",X"7E",
		X"8F",X"0F",X"1F",X"1F",X"1F",X"1F",X"0F",X"07",X"03",X"0F",X"FE",X"FC",X"F0",X"C0",X"00",X"00",
		X"1E",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"60",X"E0",X"E0",X"E0",X"E0",X"E0",X"F0",X"70",X"10",X"30",X"71",X"F3",X"F7",X"F7",X"9F",X"1C",
		X"0C",X"3C",X"7C",X"FC",X"FD",X"FD",X"CF",X"9E",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"0F",
		X"10",X"00",X"00",X"06",X"0F",X"1F",X"1F",X"9F",X"30",X"22",X"07",X"07",X"02",X"80",X"80",X"30",
		X"18",X"10",X"00",X"00",X"03",X"07",X"07",X"03",X"1E",X"18",X"30",X"20",X"40",X"00",X"00",X"00",
		X"CF",X"87",X"07",X"07",X"0F",X"0F",X"07",X"03",X"31",X"00",X"0E",X"1F",X"3F",X"7F",X"7F",X"FE",
		X"30",X"F8",X"FB",X"FB",X"38",X"18",X"18",X"10",X"00",X"00",X"03",X"07",X"06",X"04",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FF",X"FF",X"FF",X"F9",X"FC",X"EC",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"80",X"80",X"C0",X"E0",X"C0",X"F0",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"1F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"03",X"07",X"0F",X"0F",X"0F",
		X"F0",X"F8",X"00",X"00",X"80",X"E0",X"F0",X"F0",X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1C",
		X"C0",X"00",X"C0",X"F0",X"E0",X"C0",X"80",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"10",X"07",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"20",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"FE",X"FC",X"FF",X"FF",X"FF",X"FE",X"F0",X"C0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"1F",X"0F",X"0F",X"0F",X"07",X"03",X"01",X"00",X"00",
		X"00",X"00",X"00",X"80",X"C8",X"E0",X"C0",X"C0",X"00",X"00",X"07",X"0F",X"1F",X"3F",X"3F",X"FF",
		X"00",X"00",X"00",X"00",X"F0",X"F8",X"7C",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"03",
		X"00",X"00",X"00",X"00",X"00",X"20",X"60",X"70",X"80",X"C0",X"E0",X"F0",X"F8",X"F8",X"F8",X"FA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"9D",X"CF",X"E3",X"F9",X"FD",X"1C",X"1E",X"1E",
		X"03",X"03",X"03",X"81",X"E0",X"F8",X"F8",X"E0",X"78",X"7C",X"7E",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"F0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"7F",X"3F",X"BF",X"9E",X"DC",X"D0",X"C0",X"C0",
		X"0F",X"8F",X"DF",X"FF",X"FF",X"FF",X"F7",X"F7",X"80",X"03",X"01",X"1F",X"3F",X"77",X"E3",X"80",
		X"7F",X"7F",X"3F",X"3E",X"3E",X"1E",X"1E",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"E0",X"E0",X"C0",X"C0",X"C0",X"C0",X"80",X"F7",X"F7",X"E7",X"83",X"01",X"07",X"3F",X"32",
		X"E3",X"F7",X"FF",X"1F",X"07",X"00",X"00",X"00",X"06",X"03",X"01",X"00",X"00",X"00",X"00",X"00",
		X"30",X"78",X"F8",X"F8",X"FC",X"7C",X"3E",X"9E",X"30",X"22",X"07",X"07",X"02",X"80",X"80",X"30",
		X"DF",X"8F",X"0F",X"0F",X"07",X"00",X"00",X"00",X"31",X"00",X"70",X"F8",X"FC",X"FE",X"7E",X"7F",
		X"C0",X"F8",X"F8",X"C0",X"E0",X"E0",X"00",X"80",X"7F",X"7F",X"3F",X"3F",X"1F",X"0F",X"07",X"03",
		X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"00",X"00",X"00",X"1D",X"3E",X"7F",X"7F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"F0",X"10",X"10",X"10",X"10",
		X"00",X"00",X"00",X"FF",X"10",X"10",X"10",X"10",X"00",X"00",X"00",X"1F",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"F0",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"FF",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"1F",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"F0",X"00",X"00",X"00",X"00",
		X"10",X"10",X"10",X"FF",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"1F",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
