library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity sbagman_tile_bit1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of sbagman_tile_bit1 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"3E",X"41",X"41",X"41",X"41",X"41",X"3E",X"00",X"00",X"00",X"7F",X"20",X"10",X"00",X"00",
		X"00",X"31",X"49",X"49",X"49",X"49",X"49",X"27",X"00",X"46",X"69",X"59",X"49",X"41",X"41",X"41",
		X"00",X"04",X"7F",X"44",X"44",X"24",X"14",X"0C",X"00",X"46",X"49",X"49",X"49",X"49",X"49",X"79",
		X"00",X"46",X"49",X"49",X"49",X"49",X"49",X"3E",X"00",X"60",X"50",X"48",X"47",X"40",X"40",X"40",
		X"00",X"36",X"49",X"49",X"49",X"49",X"49",X"36",X"00",X"3E",X"49",X"49",X"49",X"49",X"49",X"31",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"18",X"24",X"62",X"51",X"85",X"46",X"24",X"18",X"18",X"24",X"46",X"89",X"91",X"62",X"24",X"18",
		X"18",X"24",X"42",X"D5",X"AB",X"42",X"24",X"18",X"00",X"00",X"80",X"80",X"80",X"80",X"FF",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"48",X"48",X"48",X"48",X"48",X"3F",
		X"00",X"36",X"49",X"49",X"49",X"49",X"49",X"7F",X"00",X"41",X"41",X"41",X"41",X"41",X"41",X"3E",
		X"00",X"3E",X"41",X"41",X"41",X"41",X"41",X"7F",X"00",X"41",X"41",X"49",X"49",X"49",X"49",X"7F",
		X"00",X"40",X"40",X"48",X"48",X"48",X"48",X"7F",X"00",X"4F",X"49",X"49",X"41",X"41",X"41",X"3E",
		X"00",X"7F",X"08",X"08",X"08",X"08",X"08",X"7F",X"00",X"00",X"00",X"00",X"7F",X"00",X"00",X"00",
		X"00",X"7E",X"01",X"01",X"01",X"01",X"01",X"06",X"00",X"41",X"22",X"14",X"08",X"04",X"02",X"7F",
		X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"7F",X"00",X"7F",X"20",X"10",X"08",X"10",X"20",X"7F",
		X"00",X"7F",X"02",X"04",X"08",X"10",X"20",X"7F",X"00",X"3E",X"41",X"41",X"41",X"41",X"41",X"3E",
		X"00",X"30",X"48",X"48",X"48",X"48",X"48",X"7F",X"00",X"3D",X"42",X"45",X"41",X"41",X"41",X"3E",
		X"00",X"31",X"4A",X"4C",X"48",X"48",X"48",X"7F",X"00",X"46",X"49",X"49",X"49",X"49",X"49",X"31",
		X"00",X"40",X"40",X"40",X"7F",X"40",X"40",X"40",X"00",X"7E",X"01",X"01",X"01",X"01",X"01",X"7E",
		X"00",X"78",X"04",X"02",X"01",X"02",X"04",X"78",X"00",X"7C",X"02",X"01",X"06",X"01",X"02",X"7C",
		X"00",X"41",X"22",X"14",X"08",X"14",X"22",X"41",X"00",X"40",X"20",X"10",X"0F",X"10",X"20",X"40",
		X"00",X"41",X"61",X"51",X"49",X"45",X"43",X"41",X"00",X"00",X"00",X"00",X"06",X"06",X"00",X"00",
		X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"00",X"00",X"40",X"40",X"40",X"40",X"40",X"40",X"00",
		X"00",X"00",X"00",X"00",X"28",X"00",X"00",X"00",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",
		X"00",X"00",X"82",X"C6",X"6C",X"38",X"00",X"00",X"00",X"00",X"38",X"6C",X"C6",X"82",X"00",X"00",
		X"00",X"00",X"82",X"FE",X"FE",X"82",X"00",X"00",X"82",X"FE",X"FE",X"82",X"82",X"FE",X"FE",X"82",
		X"00",X"28",X"28",X"28",X"28",X"28",X"28",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"00",
		X"F6",X"F6",X"00",X"00",X"F6",X"F6",X"00",X"00",X"FA",X"FA",X"00",X"00",X"FA",X"FA",X"00",X"00",
		X"00",X"00",X"00",X"F6",X"F6",X"00",X"00",X"00",X"00",X"00",X"00",X"FA",X"FA",X"00",X"00",X"00",
		X"00",X"00",X"00",X"E0",X"C0",X"00",X"00",X"00",X"00",X"E0",X"C0",X"00",X"E0",X"C0",X"00",X"00",
		X"00",X"60",X"E0",X"00",X"60",X"E0",X"00",X"00",X"00",X"00",X"C0",X"00",X"C0",X"00",X"00",X"00",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"FF",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"1B",X"80",X"80",X"C0",X"C0",X"80",X"44",X"54",X"55",
		X"3F",X"35",X"31",X"23",X"00",X"00",X"00",X"00",X"55",X"51",X"51",X"50",X"40",X"40",X"00",X"00",
		X"00",X"00",X"C8",X"EA",X"02",X"42",X"62",X"60",X"00",X"00",X"00",X"20",X"A8",X"A8",X"A8",X"A0",
		X"60",X"62",X"42",X"02",X"02",X"00",X"00",X"00",X"A1",X"AB",X"AB",X"AA",X"A0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"36",X"7F",X"6B",X"00",X"00",X"00",X"09",X"3B",X"2B",X"AB",X"A8",
		X"62",X"46",X"01",X"07",X"07",X"03",X"00",X"00",X"A9",X"AB",X"AB",X"AB",X"80",X"80",X"00",X"00",
		X"00",X"10",X"38",X"10",X"00",X"40",X"02",X"07",X"D7",X"D0",X"D7",X"80",X"0F",X"20",X"3F",X"00",
		X"02",X"20",X"70",X"21",X"00",X"04",X"0E",X"04",X"07",X"0C",X"1F",X"39",X"2C",X"18",X"1F",X"0F",
		X"00",X"00",X"00",X"10",X"38",X"10",X"00",X"40",X"D7",X"D0",X"D7",X"80",X"0F",X"10",X"1F",X"00",
		X"04",X"0E",X"04",X"00",X"20",X"70",X"21",X"00",X"07",X"0C",X"1F",X"39",X"2C",X"18",X"1F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D7",X"D0",X"D7",X"80",X"0F",X"10",X"1F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"0C",X"1F",X"39",X"2C",X"18",X"1F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D7",X"D0",X"D7",X"80",X"0F",X"00",X"3F",X"D0",
		X"03",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"FF",X"A0",X"AE",X"12",X"0A",X"0A",X"02",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"06",X"1F",X"00",X"00",X"00",X"11",X"17",X"97",X"07",X"05",
		X"1D",X"1D",X"01",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"D5",X"54",X"54",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"36",X"FF",X"00",X"00",X"00",X"00",X"09",X"2B",X"2B",X"AB",
		X"EA",X"EA",X"46",X"00",X"00",X"00",X"00",X"00",X"A8",X"A9",X"AB",X"AB",X"2B",X"00",X"00",X"00",
		X"00",X"03",X"01",X"00",X"01",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"80",X"80",
		X"0C",X"36",X"7F",X"6B",X"62",X"46",X"00",X"00",X"00",X"E0",X"00",X"C0",X"00",X"00",X"00",X"00",
		X"0F",X"07",X"00",X"07",X"00",X"0F",X"80",X"EF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"E8",X"1F",X"68",X"FF",X"D4",X"C7",X"8C",X"00",X"00",X"80",X"00",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"40",X"70",X"75",X"00",X"F0",X"70",X"00",X"70",X"40",X"40",X"41",
		X"05",X"1D",X"6D",X"FF",X"D5",X"C5",X"8C",X"00",X"57",X"57",X"56",X"40",X"40",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"18",X"6C",X"FE",X"00",X"00",X"78",X"B8",X"90",X"D0",X"50",X"50",
		X"D7",X"C5",X"8D",X"01",X"00",X"00",X"01",X"00",X"50",X"50",X"50",X"50",X"50",X"90",X"B8",X"3C",
		X"00",X"00",X"00",X"00",X"06",X"1B",X"3F",X"35",X"00",X"00",X"00",X"30",X"20",X"35",X"97",X"D7",
		X"31",X"23",X"00",X"00",X"00",X"00",X"00",X"00",X"53",X"50",X"50",X"54",X"54",X"54",X"DC",X"1E",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"36",X"7F",X"00",X"00",X"3C",X"DC",X"88",X"88",X"88",X"A8",
		X"6B",X"62",X"46",X"00",X"00",X"00",X"00",X"00",X"A8",X"A8",X"A8",X"A9",X"2F",X"2F",X"66",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"36",X"7F",X"00",X"00",X"00",X"00",X"09",X"2B",X"3B",X"AB",
		X"6B",X"62",X"46",X"00",X"00",X"00",X"00",X"00",X"A8",X"A9",X"AB",X"AB",X"2B",X"00",X"00",X"00",
		X"00",X"10",X"38",X"10",X"00",X"40",X"02",X"07",X"C0",X"C0",X"C0",X"80",X"00",X"3F",X"3F",X"0F",
		X"02",X"20",X"70",X"21",X"00",X"04",X"0E",X"04",X"07",X"0F",X"1F",X"7F",X"2F",X"1F",X"00",X"00",
		X"00",X"00",X"00",X"10",X"38",X"10",X"00",X"40",X"C0",X"C0",X"C0",X"80",X"00",X"1F",X"1F",X"0F",
		X"04",X"0E",X"04",X"00",X"20",X"70",X"21",X"00",X"07",X"0F",X"1F",X"7F",X"2F",X"1F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"C0",X"80",X"00",X"1F",X"1F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"0F",X"1F",X"7F",X"2F",X"1F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"C0",X"80",X"00",X"10",X"38",X"5C",
		X"02",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"7C",X"FC",X"FE",X"FF",X"FF",X"3F",X"06",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"13",X"00",X"00",X"00",X"01",X"03",X"23",X"F3",X"F0",
		X"1F",X"1F",X"07",X"07",X"01",X"00",X"00",X"00",X"F0",X"F8",X"FC",X"FC",X"FC",X"5C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"0C",X"16",X"9F",X"00",X"00",X"00",X"00",X"01",X"23",X"63",X"E3",
		X"FF",X"FF",X"3F",X"3E",X"0E",X"02",X"00",X"00",X"E0",X"E1",X"E3",X"E3",X"63",X"00",X"00",X"00",
		X"00",X"00",X"DC",X"FF",X"1F",X"3D",X"1C",X"1E",X"00",X"00",X"00",X"00",X"08",X"88",X"88",X"00",
		X"1E",X"1C",X"3D",X"1B",X"03",X"01",X"00",X"00",X"01",X"83",X"83",X"82",X"C0",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"06",X"0B",X"80",X"80",X"C0",X"C0",X"80",X"C0",X"C0",X"C1",
		X"0F",X"0F",X"0F",X"1F",X"1F",X"07",X"01",X"00",X"C1",X"E1",X"E1",X"E0",X"E0",X"40",X"00",X"00",
		X"00",X"00",X"00",X"04",X"0C",X"16",X"1F",X"1F",X"00",X"00",X"10",X"11",X"13",X"73",X"F3",X"E0",
		X"10",X"3F",X"3E",X"0E",X"07",X"03",X"00",X"00",X"E1",X"F3",X"F3",X"E3",X"C0",X"80",X"00",X"00",
		X"08",X"04",X"02",X"01",X"04",X"0C",X"16",X"1F",X"00",X"00",X"00",X"80",X"C0",X"61",X"E3",X"E3",
		X"1F",X"1F",X"3F",X"3E",X"0E",X"02",X"00",X"00",X"C3",X"C0",X"E0",X"E1",X"67",X"07",X"06",X"00",
		X"00",X"00",X"00",X"1F",X"01",X"04",X"0C",X"16",X"00",X"00",X"00",X"80",X"80",X"C1",X"E3",X"E3",
		X"1F",X"1F",X"1F",X"3F",X"3E",X"0E",X"02",X"00",X"E3",X"C0",X"C0",X"E1",X"E7",X"67",X"06",X"00",
		X"08",X"04",X"02",X"01",X"00",X"04",X"0C",X"16",X"00",X"00",X"00",X"80",X"C0",X"41",X"63",X"E3",
		X"1F",X"1F",X"1F",X"3F",X"3E",X"0E",X"02",X"00",X"E3",X"C0",X"C0",X"E1",X"E7",X"67",X"06",X"00",
		X"00",X"00",X"00",X"00",X"04",X"0C",X"16",X"1F",X"20",X"20",X"20",X"60",X"60",X"41",X"E3",X"E3",
		X"1F",X"1F",X"3F",X"3E",X"0E",X"02",X"00",X"00",X"C3",X"C0",X"E0",X"E1",X"67",X"07",X"06",X"00",
		X"00",X"00",X"00",X"02",X"06",X"0B",X"0F",X"0F",X"10",X"10",X"10",X"30",X"30",X"21",X"B3",X"F3",
		X"0F",X"1F",X"1F",X"07",X"01",X"00",X"00",X"00",X"F3",X"E0",X"E0",X"60",X"60",X"40",X"DC",X"DE",
		X"00",X"00",X"00",X"00",X"04",X"0C",X"16",X"1F",X"00",X"80",X"BC",X"DC",X"C0",X"60",X"60",X"E0",
		X"1F",X"1F",X"3F",X"3E",X"0E",X"02",X"00",X"00",X"E0",X"E0",X"E0",X"60",X"40",X"DC",X"DE",X"DE",
		X"00",X"00",X"00",X"00",X"04",X"0C",X"16",X"1F",X"40",X"40",X"7C",X"DC",X"C0",X"80",X"C0",X"C0",
		X"1F",X"1F",X"3F",X"3E",X"0E",X"02",X"00",X"00",X"C0",X"C0",X"E0",X"E1",X"67",X"27",X"66",X"60",
		X"00",X"00",X"00",X"00",X"04",X"0C",X"16",X"1F",X"00",X"00",X"00",X"10",X"11",X"13",X"33",X"33",
		X"1F",X"1F",X"3F",X"3E",X"0E",X"02",X"00",X"00",X"E0",X"E1",X"F3",X"F3",X"63",X"00",X"00",X"00",
		X"07",X"08",X"08",X"07",X"00",X"07",X"08",X"08",X"C0",X"20",X"20",X"C0",X"00",X"C0",X"20",X"20",
		X"00",X"00",X"0E",X"8C",X"CC",X"EA",X"00",X"00",X"01",X"01",X"00",X"00",X"20",X"60",X"F0",X"F0",
		X"1F",X"20",X"40",X"80",X"80",X"80",X"80",X"80",X"FF",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"80",X"80",X"80",X"80",X"80",X"40",X"20",X"1F",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"5C",X"FE",X"54",X"FE",X"54",X"74",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"9C",X"C8",X"E8",X"F2",X"F3",X"F2",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F2",X"F3",X"F2",X"E8",X"C8",X"9C",
		X"01",X"01",X"00",X"00",X"3F",X"7F",X"FF",X"FF",X"01",X"01",X"00",X"00",X"E0",X"E0",X"F0",X"F0",
		X"01",X"01",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"01",X"00",X"00",X"01",X"01",X"00",X"00",
		X"07",X"02",X"02",X"02",X"02",X"02",X"02",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"F0",X"F0",
		X"01",X"01",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"07",X"07",X"03",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"C0",X"C0",X"E0",X"E0",X"F0",X"F0",X"F8",X"F8",X"FC",X"FC",X"FE",X"FE",X"FF",X"FF",
		X"7F",X"7F",X"3F",X"3F",X"1F",X"0F",X"0F",X"07",X"07",X"07",X"03",X"03",X"01",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",
		X"00",X"00",X"00",X"00",X"40",X"70",X"78",X"0C",X"00",X"F0",X"70",X"00",X"00",X"00",X"00",X"01",
		X"0F",X"1F",X"2F",X"3F",X"3F",X"3F",X"7E",X"7C",X"87",X"87",X"86",X"80",X"80",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FB",X"FB",X"FB",X"3B",X"BC",X"04",X"04",X"04",X"02",X"02",X"03",X"01",X"01",
		X"00",X"01",X"01",X"03",X"06",X"04",X"04",X"04",X"06",X"03",X"01",X"00",X"00",X"00",X"00",X"00",
		X"35",X"17",X"17",X"13",X"0B",X"09",X"0D",X"04",X"5F",X"4F",X"4F",X"6F",X"2F",X"2F",X"27",X"27",
		X"BF",X"BF",X"9F",X"DF",X"5F",X"5F",X"57",X"5F",X"FE",X"FF",X"FE",X"FF",X"7F",X"7F",X"3F",X"BF",
		X"DE",X"BC",X"7E",X"7D",X"7F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"01",X"07",X"0C",X"39",X"67",
		X"3F",X"00",X"80",X"E1",X"3F",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"7D",X"FF",X"FF",X"EE",X"FF",
		X"FF",X"FF",X"FF",X"DF",X"FF",X"FF",X"FF",X"7F",X"FB",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3F",X"1F",X"1F",X"8F",X"6F",X"D7",X"F7",X"F7",X"7D",X"73",X"7F",X"FF",X"FF",X"FF",X"FF",X"3E",
		X"3E",X"63",X"DC",X"DF",X"7B",X"7D",X"7B",X"76",X"1C",X"36",X"63",X"C1",X"00",X"00",X"00",X"00",
		X"FF",X"BF",X"FD",X"F9",X"F1",X"E1",X"C5",X"8C",X"FF",X"FF",X"FF",X"FF",X"BF",X"FF",X"FF",X"FF",
		X"FB",X"FB",X"FD",X"FD",X"FD",X"FD",X"FE",X"FE",X"9F",X"5F",X"EF",X"FF",X"FF",X"FB",X"FB",X"FB",
		X"FF",X"FF",X"FF",X"FB",X"FB",X"FB",X"3B",X"BC",X"BF",X"BE",X"60",X"C0",X"BF",X"BF",X"7F",X"FF",
		X"07",X"1C",X"11",X"37",X"2F",X"6F",X"5F",X"DF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"08",X"0C",X"06",X"03",X"01",X"00",X"00",X"00",X"47",X"67",X"27",X"23",X"33",X"13",X"11",X"19",
		X"04",X"06",X"06",X"C6",X"46",X"46",X"46",X"46",X"BF",X"7B",X"77",X"B3",X"F0",X"E0",X"E0",X"C0",
		X"7F",X"7F",X"BF",X"BB",X"DF",X"FF",X"FF",X"9F",X"67",X"6B",X"8D",X"BE",X"DF",X"CE",X"F0",X"FF",
		X"DE",X"9E",X"AC",X"B0",X"79",X"39",X"52",X"63",X"FD",X"FC",X"F9",X"C3",X"DB",X"83",X"AD",X"0E",
		X"03",X"33",X"73",X"F3",X"F3",X"FB",X"F9",X"F9",X"16",X"06",X"F2",X"F8",X"FC",X"FE",X"87",X"03",
		X"13",X"13",X"13",X"17",X"17",X"17",X"16",X"F6",X"03",X"02",X"06",X"04",X"04",X"0C",X"08",X"18",
		X"00",X"01",X"01",X"03",X"02",X"02",X"03",X"01",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",
		X"C0",X"43",X"43",X"03",X"80",X"E0",X"3F",X"00",X"0F",X"0F",X"8F",X"8F",X"8F",X"8F",X"87",X"83",
		X"3D",X"1F",X"1F",X"1F",X"1E",X"1D",X"1F",X"0F",X"BF",X"3E",X"39",X"3F",X"3F",X"3F",X"3F",X"3E",
		X"EF",X"FB",X"7E",X"FC",X"F3",X"EF",X"5F",X"9F",X"DF",X"DF",X"DE",X"BF",X"3F",X"37",X"7E",X"FF",
		X"6F",X"6D",X"2F",X"CF",X"D7",X"DF",X"5E",X"8D",X"FF",X"FB",X"7F",X"BF",X"BF",X"1E",X"6B",X"6F",
		X"FB",X"FF",X"FE",X"FF",X"BD",X"FF",X"EF",X"FD",X"03",X"03",X"07",X"07",X"0F",X"0F",X"1F",X"FF",
		X"83",X"87",X"06",X"06",X"05",X"0D",X"0D",X"0C",X"3F",X"3F",X"3F",X"3F",X"CF",X"C1",X"C2",X"83",
		X"B9",X"A7",X"7F",X"7F",X"FF",X"FF",X"7F",X"7E",X"DF",X"BF",X"DC",X"BB",X"77",X"6F",X"7F",X"3F",
		X"06",X"1D",X"33",X"67",X"5F",X"DC",X"BB",X"B7",X"0E",X"0C",X"03",X"0F",X"38",X"E0",X"80",X"00",
		X"FC",X"FC",X"C0",X"F8",X"18",X"1C",X"0C",X"0E",X"FE",X"FE",X"FE",X"04",X"F8",X"FC",X"FC",X"FC",
		X"80",X"7C",X"FC",X"FE",X"FE",X"82",X"7C",X"FE",X"B0",X"30",X"B0",X"C0",X"F0",X"F8",X"FC",X"FC",
		X"D0",X"D0",X"D0",X"D0",X"B0",X"B0",X"B0",X"B0",X"90",X"B0",X"90",X"D0",X"D0",X"D0",X"D0",X"D0",
		X"EC",X"F8",X"78",X"F0",X"F0",X"E0",X"E0",X"C0",X"FC",X"FC",X"F4",X"FC",X"FC",X"F4",X"BC",X"FC",
		X"90",X"90",X"E0",X"E0",X"B0",X"F0",X"F8",X"78",X"7C",X"7C",X"F8",X"F8",X"70",X"40",X"B0",X"10",
		X"E0",X"F0",X"F8",X"FC",X"FC",X"FC",X"FC",X"7C",X"E0",X"F8",X"FC",X"FC",X"F8",X"F8",X"00",X"C0",
		X"F8",X"F0",X"00",X"F0",X"FC",X"FC",X"FC",X"18",X"18",X"ED",X"F7",X"F0",X"30",X"C0",X"F0",X"F0",
		X"80",X"C0",X"60",X"BF",X"40",X"3F",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"83",X"83",X"83",X"83",X"80",X"80",X"80",X"80",X"80",X"80",X"C0",X"80",X"80",X"80",
		X"FF",X"FF",X"FF",X"E0",X"C0",X"80",X"80",X"80",X"80",X"80",X"80",X"C0",X"E0",X"FF",X"FF",X"FF",
		X"80",X"80",X"C0",X"E0",X"C0",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"C0",X"C0",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"C0",X"E0",X"F0",X"E0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"E0",X"C0",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"C0",X"E0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"D8",X"B0",X"60",X"C0",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"07",X"0C",X"1B",X"36",X"6C",
		X"07",X"0F",X"18",X"F7",X"0C",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",
		X"38",X"78",X"F0",X"E0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"3C",
		X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3C",X"3C",X"3C",X"1C",X"00",X"00",X"00",X"00",X"00",X"3F",X"3F",X"3F",X"3E",X"3C",X"3C",X"3C",
		X"3E",X"63",X"DC",X"BD",X"78",X"7A",X"79",X"76",X"00",X"00",X"00",X"18",X"3C",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"03",X"FC",X"07",X"01",
		X"F0",X"F0",X"10",X"D8",X"64",X"37",X"18",X"0F",X"1F",X"3F",X"7F",X"FF",X"FC",X"F8",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"1F",X"9F",X"9F",X"5F",X"DF",X"EF",X"F7",X"1F",X"1F",X"5F",X"AF",X"FF",X"FE",X"FE",X"FE",
		X"FE",X"FE",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"1F",X"1F",X"1F",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",
		X"07",X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"1F",X"0F",X"07",X"07",X"07",
		X"DF",X"DF",X"EF",X"F5",X"FF",X"FF",X"FF",X"9F",X"00",X"00",X"03",X"07",X"07",X"00",X"00",X"00",
		X"70",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"06",X"9D",X"F3",X"2E",X"D8",
		X"00",X"00",X"01",X"03",X"07",X"FE",X"01",X"FF",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"01",X"00",X"00",
		X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"00",X"00",X"00",X"01",X"03",X"01",X"00",X"00",X"FF",X"03",X"01",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"03",X"1F",X"FF",
		X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"7F",X"FF",X"FF",X"FF",X"FF",X"03",X"01",X"00",
		X"00",X"00",X"00",X"00",X"01",X"03",X"0F",X"1F",X"C7",X"BF",X"63",X"C1",X"80",X"00",X"00",X"00",
		X"05",X"05",X"05",X"05",X"05",X"05",X"0D",X"7B",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",
		X"05",X"05",X"05",X"05",X"04",X"07",X"03",X"06",X"00",X"01",X"03",X"06",X"05",X"05",X"05",X"05",
		X"00",X"00",X"00",X"80",X"C0",X"7F",X"80",X"FF",X"01",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"FC",X"FF",X"FF",X"FF",X"FF",X"F8",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"7F",X"7F",X"70",X"40",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"00",X"03",X"03",X"03",X"03",X"00",X"00",X"00",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",
		X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"7F",X"7F",X"7F",X"7F",X"7F",X"7E",X"78",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"F8",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"C0",X"F8",X"FF",X"FF",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"FF",X"FF",X"FF",X"FC",X"D7",X"D3",X"65",X"6E",X"77",X"72",X"BC",X"BF",
		X"00",X"00",X"00",X"80",X"C0",X"7F",X"3F",X"7C",X"FF",X"80",X"7F",X"C0",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"FF",X"80",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",X"E0",X"E0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"F0",X"F0",X"F9",X"FF",X"00",X"00",X"00",
		X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"E0",X"F8",X"E0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"F8",X"F6",X"E6",X"EC",X"E0",X"D9",X"DD",X"C2",X"D3",
		X"00",X"00",X"00",X"00",X"FF",X"FC",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"F0",X"80",X"00",X"FF",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"FD",X"FC",X"FA",X"C2",X"DD",X"9B",X"B9",X"32",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"1C",X"7F",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"E0",X"F0",X"F0",X"F0",X"E0",X"00",X"C0",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",
		X"FE",X"FC",X"00",X"F0",X"F8",X"F8",X"F0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"07",X"1F",X"00",X"00",X"00",X"18",X"ED",X"F7",X"F0",X"00",X"F0",X"FC",X"FE",
		X"00",X"00",X"00",X"1F",X"07",X"01",X"00",X"00",X"80",X"80",X"80",X"80",X"C0",X"C0",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"03",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"1C",X"1E",X"18",X"10",X"18",X"10",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"18",X"24",X"42",X"42",X"24",X"18",
		X"FE",X"FC",X"FC",X"F8",X"F8",X"F8",X"B0",X"B0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"BE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"80",X"C0",X"E0",X"F0",X"F8",X"F8",X"BC",X"BE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0E",X"1F",X"1F",X"0E",X"0C",X"10",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"20",X"A0",X"40",X"40",X"A0",X"90",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"52",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"C0",
		X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"52",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"07",X"06",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"04",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"20",X"20",X"20",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0E",X"1F",X"1F",X"0E",X"04",X"04",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"14",X"0C",X"0C",X"0A",X"18",X"10",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0E",X"0F",X"0F",X"0E",X"04",X"04",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"04",X"0C",X"0C",X"0A",X"09",X"08",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"D8",X"5C",X"76",X"74",X"2C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3C",X"9C",X"C4",X"70",X"98",X"8C",X"87",X"81",X"09",X"0C",X"0E",X"1E",X"1E",X"1E",X"3C",X"3C",
		X"C0",X"40",X"60",X"30",X"18",X"0C",X"06",X"03",X"79",X"33",X"06",X"0C",X"18",X"30",X"60",X"C0",
		X"03",X"41",X"E0",X"E0",X"F0",X"F0",X"F8",X"7C",X"86",X"85",X"85",X"8D",X"BB",X"E3",X"C7",X"83",
		X"AD",X"B1",X"96",X"9A",X"94",X"96",X"98",X"8E",X"7F",X"E1",X"9E",X"BF",X"BF",X"DF",X"E3",X"AD",
		X"FB",X"0D",X"06",X"03",X"00",X"00",X"00",X"00",X"1F",X"1F",X"3F",X"3F",X"3F",X"3F",X"0E",X"A7",
		X"83",X"C6",X"6D",X"1B",X"17",X"0F",X"1F",X"1F",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"01",
		X"80",X"00",X"00",X"01",X"03",X"02",X"02",X"02",X"FF",X"FE",X"E1",X"5F",X"30",X"10",X"30",X"E0",
		X"FB",X"FD",X"FE",X"FF",X"F7",X"FB",X"FB",X"FF",X"D8",X"E8",X"EC",X"F4",X"F4",X"F6",X"FA",X"FA",
		X"00",X"80",X"C0",X"60",X"A0",X"B0",X"D0",X"D0",X"F4",X"F4",X"6C",X"98",X"F0",X"00",X"00",X"00",
		X"FD",X"FD",X"FB",X"FA",X"BA",X"BA",X"76",X"F4",X"5D",X"C5",X"BD",X"DD",X"E5",X"DD",X"D9",X"E5",
		X"FD",X"FD",X"FD",X"FE",X"FE",X"EE",X"F6",X"F6",X"7A",X"8A",X"BA",X"BA",X"CA",X"BA",X"B2",X"CB",
		X"FA",X"7A",X"0A",X"FA",X"FA",X"3A",X"CA",X"FA",X"00",X"00",X"00",X"F0",X"18",X"EC",X"F6",X"FA",
		X"00",X"00",X"00",X"01",X"07",X"04",X"05",X"05",X"06",X"03",X"03",X"02",X"02",X"03",X"02",X"02",
		X"03",X"02",X"02",X"06",X"FD",X"0B",X"87",X"8F",X"7D",X"BD",X"C5",X"BD",X"BD",X"DD",X"A5",X"BD",
		X"00",X"00",X"00",X"F8",X"8C",X"76",X"FB",X"FD",X"A0",X"60",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"80",X"C0",X"60",X"A0",X"A0",X"A0",X"A0",X"AF",X"AF",X"AF",X"AF",X"B7",X"97",X"98",X"8F",
		X"0F",X"1F",X"9F",X"DF",X"DD",X"DD",X"DE",X"EF",X"F1",X"E0",X"C0",X"80",X"80",X"01",X"03",X"07",
		X"19",X"13",X"06",X"0C",X"0C",X"24",X"76",X"F2",X"3C",X"7C",X"FE",X"7E",X"7F",X"3F",X"3E",X"3C",
		X"80",X"83",X"86",X"8C",X"98",X"F0",X"C0",X"98",X"F9",X"F6",X"EF",X"D9",X"B0",X"60",X"C0",X"80",
		X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",X"FF",X"80",X"C0",X"40",X"60",X"B8",X"CE",X"F3",X"FD",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"1F",X"09",X"06",X"0F",X"18",X"70",X"C0",
		X"37",X"EF",X"9F",X"7F",X"7F",X"3F",X"3F",X"1F",X"35",X"36",X"2A",X"2D",X"36",X"1A",X"15",X"1B",
		X"1F",X"31",X"2E",X"2F",X"2F",X"37",X"2B",X"2D",X"FD",X"FD",X"7D",X"BD",X"DD",X"6B",X"36",X"1C",
		X"DD",X"5D",X"AD",X"CD",X"FD",X"FD",X"FD",X"FD",X"00",X"00",X"00",X"00",X"7C",X"C6",X"BA",X"BB",
		X"ED",X"FD",X"FD",X"7B",X"86",X"FC",X"00",X"00",X"FA",X"F5",X"FA",X"F5",X"FA",X"F5",X"FA",X"75",
		X"7A",X"35",X"3A",X"15",X"1A",X"05",X"0A",X"05",X"1A",X"15",X"1A",X"15",X"0A",X"05",X"0A",X"05",
		X"FA",X"F5",X"7A",X"75",X"7A",X"35",X"3A",X"35",X"FA",X"F5",X"FA",X"75",X"7A",X"35",X"3A",X"15",
		X"EA",X"E5",X"CA",X"C5",X"CA",X"C5",X"CA",X"C5",X"CA",X"C5",X"8A",X"85",X"8A",X"85",X"8A",X"85",
		X"8A",X"85",X"8A",X"C5",X"CA",X"C5",X"CA",X"C5",X"CA",X"C5",X"EA",X"E5",X"EA",X"E5",X"EA",X"E5",
		X"7A",X"75",X"7A",X"75",X"FA",X"F5",X"FA",X"F5",X"1A",X"15",X"3A",X"35",X"3A",X"35",X"7A",X"75",
		X"7A",X"75",X"7A",X"75",X"3A",X"35",X"3A",X"35",X"3A",X"35",X"3A",X"35",X"7A",X"75",X"7A",X"75",
		X"EA",X"C5",X"CA",X"85",X"8A",X"05",X"0A",X"05",X"FA",X"F5",X"FA",X"F5",X"FA",X"F5",X"FA",X"E5",
		X"0A",X"85",X"CA",X"E5",X"FA",X"F5",X"FA",X"F5",X"0A",X"05",X"0A",X"05",X"0A",X"05",X"0A",X"05",
		X"FA",X"F5",X"FA",X"E5",X"EA",X"E5",X"CA",X"C5",X"CA",X"C5",X"8A",X"85",X"8A",X"85",X"8A",X"85",
		X"8A",X"85",X"8A",X"85",X"8A",X"85",X"8A",X"C5",X"CA",X"C5",X"CA",X"C5",X"CA",X"C5",X"EA",X"E5",
		X"0A",X"05",X"0A",X"05",X"0A",X"05",X"0A",X"05",X"1A",X"15",X"1A",X"15",X"3A",X"75",X"7A",X"75",
		X"FA",X"F5",X"FA",X"F5",X"FA",X"F5",X"FA",X"F5",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"40",X"20",X"10",X"08",X"04",X"FF",X"04",X"08",X"10",X"20",X"40",X"80",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"50",X"A0",X"50",X"A0",X"50",X"A0",X"50",X"A0",X"50",X"A0",X"40",X"A0",X"50",
		X"A0",X"50",X"A0",X"50",X"A0",X"50",X"A0",X"50",X"A0",X"50",X"A0",X"50",X"A0",X"50",X"A0",X"50",
		X"A0",X"50",X"A0",X"40",X"A0",X"50",X"A0",X"50",X"A0",X"50",X"A0",X"50",X"A0",X"00",X"00",X"00",
		X"04",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"04",X"08",X"10",X"3E",X"00",X"1A",
		X"24",X"24",X"24",X"3E",X"00",X"3E",X"02",X"02",X"02",X"3E",X"00",X"20",X"20",X"3E",X"20",X"20",
		X"00",X"22",X"2A",X"2A",X"2A",X"3E",X"00",X"1A",X"24",X"24",X"24",X"3E",X"00",X"00",X"00",X"00",
		X"00",X"02",X"02",X"02",X"02",X"3E",X"00",X"3E",X"02",X"02",X"02",X"3E",X"00",X"22",X"22",X"22",
		X"22",X"3E",X"00",X"22",X"2A",X"2A",X"2A",X"3E",X"00",X"1A",X"24",X"24",X"24",X"3E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"22",X"2A",X"2A",X"2A",X"3E",X"00",X"2E",X"2A",X"2A",X"2A",X"3A",
		X"00",X"1E",X"24",X"24",X"24",X"1E",X"00",X"1A",X"24",X"24",X"24",X"3E",X"00",X"22",X"2A",X"2A",
		X"2A",X"3E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",
		X"20",X"3E",X"20",X"20",X"00",X"3E",X"04",X"08",X"10",X"3E",X"00",X"22",X"2A",X"2A",X"2A",X"3E",
		X"00",X"3E",X"10",X"08",X"10",X"3E",X"00",X"22",X"2A",X"2A",X"2A",X"3E",X"00",X"22",X"22",X"22",
		X"22",X"3E",X"20",X"1E",X"24",X"24",X"24",X"1E",X"00",X"20",X"28",X"28",X"28",X"3E",X"00",X"20",
		X"28",X"28",X"28",X"3E",X"00",X"22",X"2A",X"2A",X"2A",X"3E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"2A",X"2A",X"2A",X"3E",X"00",X"22",X"22",X"22",X"22",
		X"3E",X"00",X"3E",X"04",X"08",X"10",X"3E",X"00",X"1E",X"24",X"24",X"24",X"1E",X"00",X"38",X"04",
		X"02",X"04",X"38",X"00",X"1C",X"22",X"22",X"22",X"3E",X"00",X"1E",X"24",X"24",X"24",X"1E",X"00",
		X"00",X"00",X"00",X"00",X"22",X"2A",X"2A",X"2A",X"3E",X"00",X"22",X"22",X"22",X"22",X"3E",X"00",
		X"3E",X"04",X"08",X"10",X"3E",X"00",X"1E",X"24",X"24",X"24",X"1E",X"00",X"38",X"04",X"02",X"04",
		X"38",X"00",X"1E",X"24",X"24",X"24",X"1A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"2A",
		X"2A",X"2A",X"3E",X"00",X"1A",X"24",X"24",X"24",X"3E",X"00",X"3E",X"02",X"02",X"02",X"3E",X"00",
		X"20",X"20",X"3E",X"20",X"20",X"00",X"3E",X"00",X"00",X"1A",X"24",X"24",X"24",X"3E",X"00",X"22",
		X"22",X"22",X"22",X"3E",X"00",X"22",X"2A",X"2A",X"2A",X"3E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"2A",X"2A",X"2A",X"3E",X"00",X"20",X"20",X"3E",
		X"20",X"20",X"00",X"3E",X"00",X"1A",X"24",X"24",X"24",X"3E",X"00",X"38",X"04",X"02",X"3C",X"02",
		X"08",X"08",X"08",X"08",X"08",X"0C",X"06",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"08",X"08",X"08",X"08",X"08",X"18",X"30",X"E0",X"E0",X"30",X"18",X"08",X"08",X"08",X"08",X"08",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"06",X"0C",X"08",X"08",X"08",X"08",X"08",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"02",X"02",X"02",X"06",X"FD",X"03",X"FE",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"03",X"03",X"07",X"02",X"02",X"02",X"02",X"02",
		X"3C",X"38",X"38",X"3C",X"0E",X"06",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"06",X"0E",
		X"02",X"02",X"02",X"02",X"02",X"06",X"0E",X"06",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"06",X"0D",X"06",
		X"1D",X"7B",X"F6",X"F6",X"FB",X"05",X"05",X"06",X"06",X"06",X"02",X"02",X"02",X"02",X"06",X"0E",
		X"02",X"06",X"1D",X"FB",X"F6",X"FB",X"3D",X"0C",X"0D",X"0D",X"02",X"02",X"02",X"02",X"02",X"02",
		X"1D",X"05",X"06",X"02",X"02",X"02",X"02",X"06",X"02",X"02",X"06",X"0E",X"3D",X"3B",X"36",X"3B",
		X"02",X"02",X"06",X"0D",X"06",X"02",X"02",X"02",X"F6",X"FB",X"0D",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"05",X"0D",X"FB",X"F8",X"0C",X"F6",X"1B",X"0D",X"06",X"02",X"02",
		X"F4",X"F4",X"F4",X"F6",X"FB",X"FD",X"FD",X"DD",X"F4",X"F4",X"F4",X"F4",X"F4",X"F4",X"F4",X"F4",
		X"00",X"C0",X"60",X"B0",X"D8",X"E8",X"E8",X"E8",X"CD",X"86",X"83",X"81",X"80",X"80",X"80",X"80",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"CF",X"B7",X"7B",X"03",X"E1",X"3B",X"CE",X"F6",X"FB",X"FD",X"FE",
		X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"01",X"FE",X"C0",X"60",X"38",X"0F",X"01",X"06",X"07",X"07",
		X"EC",X"D8",X"30",X"E0",X"00",X"00",X"00",X"00",X"34",X"F4",X"F4",X"F4",X"F4",X"F4",X"F4",X"F4",
		X"C6",X"FF",X"19",X"E8",X"EC",X"74",X"74",X"B4",X"8F",X"8F",X"8F",X"8F",X"8E",X"8E",X"8E",X"01",
		X"00",X"00",X"01",X"03",X"FE",X"0D",X"83",X"8F",X"FD",X"7D",X"9B",X"E6",X"3C",X"00",X"00",X"00",
		X"FD",X"FD",X"FD",X"FB",X"FB",X"FD",X"ED",X"ED",X"DD",X"C5",X"BD",X"5D",X"E5",X"DD",X"D9",X"E5",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"02",X"02",X"02",
		X"30",X"60",X"C0",X"80",X"80",X"01",X"03",X"07",X"06",X"FF",X"41",X"60",X"B8",X"CE",X"F3",X"FD",
		X"7D",X"FD",X"9B",X"E6",X"7C",X"C6",X"BA",X"BB",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0A",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"00",
		X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"80",X"80",X"80",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",
		X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"04",X"04",X"04",X"0C",X"0C",X"0C",X"0C",X"0C",
		X"0C",X"0C",X"0C",X"0C",X"04",X"06",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"04",X"04",
		X"04",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"04",X"04",X"02",X"03",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"04",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"07",X"00",X"00",X"03",X"04",X"04",
		X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"06",X"01",X"00",X"00",X"00",X"01",X"02",X"02",X"04",
		X"04",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"04",X"04",X"02",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"02",X"04",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",
		X"0C",X"04",X"06",X"01",X"00",X"00",X"00",X"00",X"01",X"02",X"04",X"04",X"0C",X"0C",X"0C",X"0C",
		X"0C",X"0C",X"0C",X"0C",X"0C",X"04",X"03",X"00",X"00",X"00",X"00",X"01",X"06",X"04",X"04",X"0C",
		X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"04",X"04",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"04",X"04",X"04",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"04",X"03",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"20",X"E0",X"E0",X"E0",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"0F",X"3F",X"FF",X"FF",X"FF",X"E7",X"87",X"07",X"07",X"07",X"07",X"87",X"E7",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"03",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"E0",X"E0",X"20",X"00",X"00",X"00",
		X"3F",X"0F",X"07",X"07",X"07",X"07",X"07",X"07",X"00",X"E0",X"E0",X"E0",X"C0",X"C0",X"C0",X"80",
		X"07",X"3F",X"3F",X"3F",X"1F",X"1F",X"1F",X"0F",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"E0",
		X"0F",X"0F",X"07",X"07",X"07",X"07",X"07",X"3F",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"80",X"00",X"00",X"00",
		X"3F",X"07",X"07",X"07",X"07",X"C7",X"F7",X"FF",X"FF",X"7F",X"1F",X"07",X"01",X"00",X"00",X"00",
		X"00",X"01",X"07",X"1F",X"7F",X"FF",X"FC",X"F8",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"04",X"07",X"07",X"07",X"07",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"07",X"07",X"07",X"04",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"12",X"01",X"00",X"22",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"05",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"50",X"00",X"00",X"00",X"00",X"02",X"15",X"2A",X"55",
		X"00",X"00",X"00",X"00",X"80",X"40",X"A8",X"55",X"00",X"01",X"02",X"15",X"AA",X"55",X"AA",X"55",
		X"80",X"40",X"80",X"50",X"A8",X"55",X"AA",X"55",X"0A",X"15",X"2A",X"55",X"AA",X"55",X"AA",X"55",
		X"0A",X"50",X"A8",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",
		X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"FF",X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",X"FF",
		X"00",X"04",X"44",X"40",X"00",X"08",X"08",X"00",X"00",X"00",X"00",X"02",X"02",X"40",X"40",X"00",
		X"00",X"02",X"42",X"00",X"00",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"00",X"00",
		X"00",X"00",X"00",X"20",X"20",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"02",X"02",X"20",X"00",
		X"00",X"02",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",
		X"00",X"04",X"44",X"40",X"00",X"08",X"08",X"00",X"00",X"00",X"00",X"02",X"02",X"40",X"40",X"00",
		X"00",X"02",X"42",X"00",X"00",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"00",X"00",
		X"00",X"00",X"00",X"20",X"20",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"02",X"02",X"20",X"00",
		X"00",X"02",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",
		X"7F",X"3F",X"3F",X"1F",X"1F",X"0F",X"0F",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",
		X"80",X"C0",X"C0",X"C0",X"E0",X"E0",X"E0",X"F0",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",
		X"FF",X"FE",X"FE",X"FE",X"00",X"00",X"10",X"10",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",
		X"07",X"07",X"07",X"07",X"00",X"00",X"10",X"10",X"E0",X"C0",X"00",X"00",X"00",X"00",X"10",X"10",
		X"01",X"01",X"00",X"00",X"E0",X"E0",X"E0",X"E0",X"01",X"01",X"00",X"00",X"1F",X"1F",X"0F",X"0F",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"E0",X"E0",X"F0",X"F0",
		X"FE",X"FE",X"FC",X"FC",X"FC",X"F8",X"F8",X"F8",X"07",X"07",X"06",X"04",X"00",X"00",X"10",X"10",
		X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"F0",X"F0",X"E0",X"E0",X"C0",X"C0",X"80",X"00",
		X"80",X"80",X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"80",X"80",
		X"1F",X"0F",X"0F",X"0F",X"0F",X"07",X"07",X"07",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"E0",
		X"00",X"80",X"80",X"C0",X"C0",X"E0",X"E0",X"F0",X"F0",X"F8",X"F8",X"FC",X"FC",X"FE",X"FE",X"FE",
		X"7E",X"FF",X"F3",X"AD",X"AD",X"DD",X"FF",X"9F",X"FF",X"FF",X"81",X"F7",X"F7",X"81",X"FF",X"BF",
		X"81",X"BF",X"FF",X"81",X"FF",X"81",X"DF",X"EF",X"DF",X"81",X"FF",X"F3",X"AD",X"AD",X"DD",X"FF",
		X"81",X"F7",X"EF",X"81",X"FF",X"83",X"FD",X"FD",X"83",X"FF",X"B1",X"BD",X"BD",X"C3",X"FF",X"7E",
		X"7E",X"FF",X"FF",X"FF",X"B5",X"B5",X"81",X"FF",X"81",X"FF",X"CD",X"B3",X"B7",X"81",X"FF",X"B5",
		X"B5",X"81",X"FF",X"CD",X"B3",X"B7",X"81",X"FF",X"83",X"FD",X"FD",X"83",X"FF",X"81",X"DF",X"EF",
		X"DF",X"81",X"FF",X"CD",X"B3",X"B7",X"81",X"FF",X"C1",X"B7",X"B7",X"C1",X"FF",X"FF",X"FF",X"7E",
		X"00",X"1C",X"3C",X"38",X"38",X"1C",X"1C",X"00",X"00",X"06",X"0E",X"0E",X"06",X"06",X"02",X"00",
		X"00",X"3C",X"6A",X"56",X"6A",X"56",X"6A",X"56",X"6A",X"56",X"6A",X"56",X"6A",X"56",X"3C",X"00",
		X"00",X"00",X"00",X"10",X"38",X"3C",X"3E",X"3E",X"1E",X"1E",X"0E",X"0E",X"0C",X"08",X"10",X"00",
		X"0A",X"05",X"0A",X"05",X"0A",X"05",X"0A",X"05",X"00",X"00",X"30",X"38",X"7C",X"7C",X"7C",X"78",
		X"78",X"78",X"10",X"18",X"08",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"40",X"20",X"10",X"08",X"04",X"FF",X"04",X"08",X"10",X"20",X"40",X"80",X"00",
		X"FF",X"02",X"04",X"08",X"10",X"20",X"40",X"55",X"AA",X"40",X"20",X"10",X"08",X"04",X"02",X"FF",
		X"FF",X"40",X"20",X"10",X"08",X"04",X"02",X"55",X"AA",X"02",X"04",X"08",X"10",X"20",X"40",X"FF",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"10",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"40",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"3C",X"7E",X"7E",X"3E",
		X"3E",X"1C",X"1C",X"18",X"18",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"02",X"00",X"00",X"00",
		X"40",X"00",X"00",X"04",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3E",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"3E",X"00",
		X"00",X"3C",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"3C",X"00",
		X"A0",X"40",X"A0",X"40",X"00",X"00",X"00",X"00",X"A0",X"55",X"AA",X"40",X"A0",X"40",X"A0",X"40",
		X"A0",X"40",X"A0",X"40",X"A0",X"40",X"A0",X"40",X"40",X"40",X"20",X"20",X"10",X"10",X"28",X"28",
		X"24",X"24",X"22",X"26",X"25",X"25",X"24",X"66",X"44",X"78",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"40",X"20",X"20",X"10",X"10",X"08",X"08",X"14",X"14",X"12",X"12",X"11",X"13",X"12",X"12",
		X"12",X"33",X"22",X"3C",X"00",X"00",X"00",X"00",X"40",X"40",X"20",X"A0",X"10",X"10",X"08",X"08",
		X"04",X"04",X"0A",X"0A",X"09",X"09",X"08",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"20",X"40",X"44",X"C0",X"B0",X"A0",X"E0",X"C0",X"E0",X"80",X"C0",X"C0",X"E0",X"E0",X"B0",
		X"90",X"90",X"88",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"04",
		X"04",X"04",X"06",X"06",X"0B",X"07",X"1B",X"01",X"03",X"03",X"07",X"0F",X"33",X"06",X"04",X"18",
		X"10",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"20",X"40",X"40",X"D0",X"B0",X"E0",X"C0",X"C0",X"E0",X"80",X"C0",X"C0",X"E0",X"C0",X"80",
		X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",
		X"04",X"04",X"06",X"02",X"03",X"07",X"03",X"01",X"03",X"03",X"07",X"0F",X"13",X"02",X"04",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"40",
		X"00",X"D0",X"80",X"C0",X"C0",X"C0",X"C0",X"80",X"C0",X"80",X"80",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"02",
		X"00",X"01",X"05",X"02",X"00",X"00",X"00",X"01",X"07",X"01",X"02",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"00",X"00",X"01",X"01",X"00",X"00",X"05",X"02",X"04",X"88",X"50",X"20",X"40",X"88",
		X"00",X"00",X"AC",X"00",X"00",X"08",X"00",X"20",X"06",X"0D",X"0B",X"09",X"09",X"0B",X"0D",X"09",
		X"09",X"0D",X"0B",X"09",X"09",X"0B",X"0D",X"09",X"09",X"0D",X"0B",X"09",X"09",X"0B",X"0D",X"06",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"80",X"04",X"80",X"40",X"28",X"10",X"20",
		X"05",X"FA",X"04",X"88",X"50",X"20",X"50",X"A8",X"05",X"FA",X"04",X"8A",X"51",X"BF",X"40",X"80",
		X"01",X"02",X"05",X"08",X"10",X"2F",X"50",X"88",X"01",X"03",X"05",X"09",X"11",X"2F",X"51",X"89",
		X"05",X"FA",X"04",X"88",X"50",X"A0",X"40",X"80",X"FF",X"20",X"51",X"0A",X"04",X"FF",X"00",X"00",
		X"FF",X"82",X"44",X"28",X"10",X"FF",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"FF",X"21",X"11",X"09",X"05",X"03",X"01",X"01",X"01",X"03",X"05",X"09",X"11",X"21",X"FF",
		X"01",X"FF",X"03",X"05",X"09",X"11",X"21",X"41",X"81",X"41",X"21",X"11",X"09",X"05",X"03",X"FF",
		X"02",X"FF",X"22",X"12",X"0A",X"06",X"02",X"03",X"02",X"03",X"02",X"06",X"0A",X"12",X"22",X"FF",
		X"02",X"FF",X"02",X"06",X"0A",X"12",X"22",X"42",X"82",X"42",X"22",X"12",X"0A",X"06",X"02",X"FF",
		X"04",X"FF",X"24",X"14",X"0C",X"04",X"06",X"05",X"04",X"05",X"06",X"04",X"0C",X"14",X"24",X"FF",
		X"04",X"FF",X"06",X"04",X"0C",X"14",X"24",X"44",X"84",X"44",X"24",X"14",X"0C",X"04",X"06",X"FF",
		X"08",X"FF",X"28",X"18",X"08",X"0C",X"0A",X"09",X"08",X"09",X"0A",X"0C",X"08",X"18",X"28",X"FF",
		X"08",X"FF",X"0A",X"0C",X"08",X"18",X"28",X"48",X"88",X"48",X"28",X"18",X"08",X"0C",X"0A",X"FF",
		X"10",X"FF",X"30",X"10",X"18",X"14",X"12",X"11",X"10",X"11",X"12",X"14",X"18",X"10",X"30",X"FF",
		X"10",X"FF",X"12",X"14",X"18",X"10",X"30",X"50",X"90",X"50",X"30",X"10",X"18",X"14",X"12",X"FF",
		X"20",X"FF",X"20",X"30",X"28",X"24",X"22",X"21",X"20",X"21",X"22",X"24",X"28",X"30",X"20",X"FF",
		X"20",X"FF",X"22",X"24",X"28",X"30",X"20",X"60",X"A0",X"60",X"20",X"30",X"28",X"24",X"22",X"FF",
		X"40",X"FF",X"60",X"50",X"48",X"44",X"42",X"41",X"40",X"41",X"42",X"44",X"48",X"50",X"60",X"FF",
		X"40",X"FF",X"42",X"44",X"48",X"50",X"60",X"40",X"C0",X"40",X"60",X"50",X"48",X"44",X"42",X"FF",
		X"80",X"FF",X"A0",X"90",X"88",X"84",X"82",X"81",X"80",X"81",X"82",X"84",X"88",X"90",X"A0",X"FF",
		X"80",X"FF",X"82",X"84",X"88",X"90",X"A0",X"C0",X"80",X"C0",X"A0",X"90",X"88",X"84",X"82",X"FF",
		X"00",X"FF",X"20",X"10",X"08",X"04",X"02",X"01",X"00",X"01",X"02",X"04",X"08",X"10",X"20",X"FF",
		X"00",X"FF",X"02",X"04",X"08",X"10",X"20",X"40",X"80",X"40",X"20",X"10",X"08",X"04",X"02",X"FF",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"1C",X"1A",X"1A",X"1A",X"1E",X"1F",X"18",
		X"00",X"4F",X"5F",X"5F",X"5F",X"7F",X"7F",X"00",X"00",X"F9",X"FB",X"FB",X"FB",X"7F",X"7F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"09",X"09",X"19",X"11",X"1E",X"00",X"00",
		X"40",X"C0",X"A0",X"A0",X"90",X"D0",X"88",X"08",X"04",X"04",X"02",X"02",X"05",X"05",X"04",X"04",
		X"04",X"04",X"04",X"04",X"04",X"0C",X"08",X"0F",X"40",X"40",X"20",X"60",X"50",X"50",X"48",X"68",
		X"44",X"84",X"02",X"02",X"01",X"01",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"06",
		X"04",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"20",X"20",X"10",X"30",X"28",X"28",
		X"24",X"34",X"22",X"C2",X"01",X"01",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"03",X"02",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"00",
		X"40",X"40",X"A0",X"A0",X"90",X"90",X"88",X"98",X"94",X"94",X"92",X"9A",X"11",X"E1",X"00",X"00",
		X"40",X"40",X"20",X"20",X"50",X"50",X"48",X"48",X"44",X"4C",X"4A",X"4A",X"49",X"CD",X"88",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"01",X"01",X"01",X"01",X"01",X"01",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"11",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"F0",X"F0",
		X"01",X"01",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"07",X"07",X"03",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"C0",X"C0",X"E0",X"E0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"05",X"02",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"01",X"02",X"05",
		X"0B",X"05",X"0A",X"16",X"2C",X"14",X"28",X"58",X"B0",X"50",X"A0",X"60",X"C0",X"40",X"80",X"80",
		X"80",X"80",X"C0",X"40",X"A0",X"60",X"B0",X"50",X"28",X"58",X"2C",X"14",X"0A",X"16",X"0B",X"05",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"40",X"A0",X"50",X"28",X"14",X"0A",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"05",X"0A",X"14",X"28",X"50",X"A0",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"11",
		X"11",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"11",
		X"11",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
