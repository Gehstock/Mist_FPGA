library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity pooyan_sprite_grphx1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of pooyan_sprite_grphx1 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"30",X"10",X"00",X"00",X"00",X"00",
		X"E0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"88",X"E8",X"30",X"30",X"31",X"00",X"10",X"30",X"31",X"71",X"F2",X"F2",X"EE",
		X"88",X"00",X"88",X"FC",X"F8",X"F7",X"F7",X"F0",X"00",X"00",X"00",X"80",X"E0",X"F0",X"C0",X"80",
		X"31",X"30",X"30",X"E8",X"88",X"00",X"00",X"00",X"EE",X"F2",X"F2",X"71",X"31",X"30",X"10",X"00",
		X"F3",X"F7",X"F7",X"FB",X"FC",X"88",X"00",X"88",X"80",X"C8",X"F8",X"E0",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"77",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"88",X"CC",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"20",X"32",X"33",X"00",X"00",X"10",X"77",X"FF",X"F7",X"FF",X"FF",
		X"00",X"00",X"80",X"CC",X"EE",X"FE",X"FE",X"FF",X"00",X"00",X"00",X"00",X"51",X"79",X"68",X"E0",
		X"33",X"11",X"11",X"20",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"77",X"00",X"00",X"00",
		X"FF",X"FE",X"EE",X"CC",X"88",X"00",X"00",X"00",X"F1",X"F1",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"20",X"10",X"33",X"33",X"00",X"00",X"00",X"77",X"F7",X"FF",X"BF",X"FE",
		X"00",X"00",X"02",X"89",X"CC",X"DC",X"FE",X"F6",X"00",X"00",X"00",X"22",X"F3",X"F3",X"E2",X"E0",
		X"33",X"33",X"31",X"00",X"00",X"00",X"00",X"00",X"FE",X"BF",X"FF",X"FF",X"77",X"00",X"00",X"00",
		X"F6",X"FE",X"DC",X"CC",X"89",X"02",X"00",X"00",X"E0",X"E2",X"F3",X"F3",X"22",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"11",X"11",X"33",X"33",X"66",X"00",X"00",X"FF",X"FF",X"FE",X"FD",X"FC",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E2",X"F3",X"33",X"33",X"11",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"EE",X"FF",X"FF",X"30",X"30",
		X"00",X"10",X"FC",X"EC",X"10",X"70",X"F0",X"30",X"33",X"C0",X"F1",X"33",X"F1",X"F4",X"FE",X"FE",
		X"91",X"40",X"B8",X"DC",X"FC",X"FC",X"F6",X"F7",X"88",X"80",X"00",X"80",X"C0",X"80",X"C0",X"80",
		X"10",X"10",X"31",X"F1",X"70",X"10",X"00",X"00",X"F4",X"FC",X"FE",X"FE",X"FC",X"F1",X"33",X"11",
		X"77",X"77",X"F7",X"E6",X"CC",X"CC",X"CC",X"88",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"B0",X"10",X"33",X"77",X"33",X"10",X"30",X"70",X"00",X"80",X"C0",X"C8",X"EC",X"EE",X"E2",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"76",X"00",X"00",X"00",X"60",X"66",X"EE",X"F1",X"F1",
		X"30",X"10",X"33",X"77",X"33",X"10",X"B0",X"C0",X"E2",X"EE",X"EC",X"C8",X"C0",X"80",X"00",X"00",
		X"70",X"70",X"FC",X"FF",X"F3",X"F1",X"F1",X"F5",X"F2",X"F0",X"F0",X"F0",X"F1",X"E8",X"AA",X"99",
		X"F6",X"F6",X"D4",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F3",X"FF",X"FF",X"77",X"FF",X"EE",X"88",X"00",X"99",X"99",X"88",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"20",X"32",X"33",X"00",X"00",X"10",X"77",X"FF",X"F7",X"FF",X"FF",
		X"00",X"00",X"80",X"CC",X"EE",X"FE",X"FF",X"FF",X"00",X"00",X"00",X"00",X"C0",X"F1",X"F1",X"68",
		X"33",X"11",X"11",X"20",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"77",X"00",X"00",X"00",
		X"FE",X"FE",X"EE",X"CC",X"88",X"00",X"00",X"00",X"68",X"B1",X"D1",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"10",X"31",X"33",X"76",X"BC",X"60",X"E0",X"E6",X"FF",X"EE",X"E8",X"E0",X"F0",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"76",X"33",X"31",X"10",X"10",X"00",X"00",X"00",X"E0",X"E8",X"EE",X"FF",X"E6",X"E0",X"60",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FC",X"CC",X"10",X"70",X"F1",X"31",X"10",X"00",X"F0",X"73",X"F3",X"FD",X"FE",X"FE",X"FC",
		X"00",X"00",X"80",X"C8",X"EC",X"F4",X"F6",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C8",
		X"10",X"30",X"F0",X"70",X"10",X"00",X"00",X"00",X"F4",X"FE",X"FE",X"F5",X"F3",X"33",X"00",X"11",
		X"77",X"F6",X"F4",X"FC",X"98",X"30",X"40",X"99",X"88",X"C0",X"C0",X"C0",X"80",X"00",X"80",X"88",
		X"74",X"F8",X"F0",X"F1",X"B3",X"32",X"E1",X"71",X"C0",X"F1",X"F1",X"E8",X"BF",X"7E",X"FE",X"F7",
		X"00",X"00",X"00",X"00",X"EE",X"FF",X"FF",X"F2",X"00",X"00",X"00",X"00",X"00",X"50",X"F8",X"EC",
		X"76",X"DD",X"DD",X"11",X"11",X"11",X"00",X"00",X"F8",X"F8",X"F2",X"F1",X"F4",X"F2",X"FC",X"33",
		X"FD",X"F7",X"F3",X"F3",X"F3",X"F7",X"FF",X"EE",X"CC",X"CC",X"CC",X"CC",X"CC",X"E8",X"C0",X"00",
		X"99",X"FF",X"77",X"FF",X"FF",X"FF",X"FF",X"67",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"33",X"FF",X"FF",X"FB",X"FD",X"F9",X"00",X"00",X"88",X"CC",X"CC",X"EF",X"EF",X"EF",
		X"77",X"33",X"11",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"70",X"00",X"00",X"00",X"00",
		X"F3",X"B3",X"80",X"00",X"11",X"11",X"33",X"33",X"CC",X"88",X"CC",X"EE",X"EE",X"CC",X"88",X"00",
		X"00",X"76",X"74",X"70",X"71",X"71",X"70",X"74",X"00",X"D0",X"90",X"E6",X"DF",X"BE",X"7F",X"FF",
		X"00",X"00",X"88",X"88",X"F7",X"FC",X"F0",X"F2",X"00",X"00",X"00",X"00",X"CC",X"E2",X"EA",X"F5",
		X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FD",X"FE",X"FE",X"FF",X"76",X"33",X"71",X"30",
		X"F1",X"F8",X"FC",X"F7",X"FF",X"FF",X"FF",X"00",X"F1",X"F3",X"F7",X"FF",X"EE",X"EC",X"E8",X"40",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"B0",X"10",X"33",X"77",X"33",X"10",X"30",X"70",X"00",X"80",X"C0",X"C8",X"EC",X"EE",X"E2",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"10",X"33",X"77",X"33",X"10",X"30",X"00",X"E2",X"EE",X"EC",X"C8",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"11",X"30",X"70",X"70",X"70",
		X"00",X"88",X"CC",X"88",X"C0",X"E0",X"E0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"70",X"70",X"70",X"30",X"11",X"33",X"11",
		X"C0",X"E0",X"E0",X"E0",X"C0",X"88",X"CC",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"10",X"31",X"33",X"76",X"BC",X"60",X"E0",X"E6",X"EE",X"EE",X"E8",X"E0",X"E0",
		X"F0",X"00",X"60",X"51",X"33",X"77",X"77",X"77",X"F0",X"00",X"77",X"FF",X"FF",X"FF",X"FF",X"FD",
		X"76",X"33",X"31",X"10",X"10",X"00",X"00",X"00",X"E0",X"E8",X"EE",X"EE",X"E6",X"E0",X"60",X"00",
		X"77",X"77",X"77",X"33",X"33",X"00",X"00",X"00",X"FD",X"32",X"77",X"FF",X"FF",X"FE",X"30",X"00",
		X"F0",X"00",X"CC",X"EE",X"FF",X"FF",X"FF",X"FF",X"F0",X"88",X"CC",X"FC",X"74",X"7C",X"18",X"B0",
		X"B0",X"10",X"33",X"77",X"B3",X"90",X"B0",X"F0",X"00",X"80",X"C0",X"C8",X"EC",X"EE",X"E2",X"E0",
		X"FD",X"FD",X"F3",X"FE",X"EC",X"C0",X"80",X"00",X"7C",X"7C",X"F4",X"7C",X"7C",X"74",X"44",X"44",
		X"B0",X"90",X"B3",X"F7",X"B3",X"10",X"30",X"00",X"E2",X"EE",X"EC",X"C8",X"C0",X"80",X"00",X"00",
		X"80",X"60",X"10",X"00",X"00",X"00",X"00",X"00",X"44",X"44",X"F4",X"44",X"E4",X"40",X"00",X"00",
		X"20",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"88",X"88",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",
		X"88",X"88",X"88",X"88",X"88",X"88",X"C8",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"D1",X"F5",X"73",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",
		X"00",X"00",X"88",X"DD",X"DE",X"FE",X"DE",X"FC",X"00",X"00",X"00",X"D1",X"F1",X"F1",X"E0",X"E0",
		X"FF",X"77",X"77",X"33",X"11",X"00",X"00",X"00",X"FB",X"FC",X"FF",X"FF",X"FF",X"F0",X"00",X"00",
		X"DA",X"F5",X"DF",X"DD",X"BB",X"11",X"00",X"00",X"E0",X"E0",X"F9",X"F9",X"D9",X"00",X"00",X"00",
		X"F0",X"00",X"00",X"CC",X"EE",X"FF",X"FF",X"FE",X"F0",X"00",X"88",X"CC",X"FC",X"BC",X"BC",X"F8",
		X"B0",X"10",X"33",X"77",X"33",X"90",X"B0",X"F0",X"00",X"80",X"C0",X"C8",X"EC",X"EE",X"E2",X"E0",
		X"FD",X"F3",X"77",X"33",X"33",X"11",X"00",X"00",X"BC",X"BC",X"F8",X"BC",X"BC",X"34",X"74",X"44",
		X"B0",X"90",X"B3",X"F7",X"B3",X"90",X"30",X"00",X"E2",X"EE",X"EC",X"C8",X"C0",X"80",X"00",X"00",
		X"C0",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"60",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"60",X"10",X"00",X"00",X"00",X"00",X"22",X"00",X"30",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"30",X"C0",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"22",X"00",X"00",X"00",X"00",X"10",X"AA",X"FF",X"BB",
		X"77",X"10",X"32",X"F3",X"F1",X"FC",X"FE",X"FE",X"00",X"22",X"22",X"B1",X"D1",X"C0",X"C0",X"C0",
		X"00",X"00",X"00",X"00",X"55",X"70",X"10",X"00",X"22",X"00",X"00",X"10",X"74",X"F0",X"E0",X"80",
		X"FC",X"FE",X"F6",X"F6",X"F6",X"70",X"10",X"10",X"E0",X"F0",X"F0",X"E0",X"C8",X"C8",X"80",X"00",
		X"00",X"33",X"10",X"10",X"11",X"22",X"11",X"33",X"70",X"F0",X"F0",X"F0",X"A5",X"FF",X"F8",X"F4",
		X"E2",X"31",X"30",X"F0",X"B5",X"EE",X"FF",X"F7",X"00",X"88",X"00",X"00",X"00",X"88",X"00",X"88",
		X"77",X"77",X"77",X"77",X"22",X"33",X"31",X"30",X"F1",X"F8",X"FC",X"FF",X"FF",X"FF",X"DD",X"77",
		X"F3",X"F2",X"F5",X"FB",X"FB",X"FF",X"FF",X"DC",X"CC",X"C4",X"CC",X"CC",X"CC",X"88",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"20",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"2B",X"37",X"00",X"00",X"00",X"30",X"60",X"58",X"38",X"0C",X"FE",
		X"00",X"00",X"00",X"E0",X"90",X"70",X"E1",X"E1",X"00",X"00",X"00",X"00",X"00",X"80",X"0C",X"8C",
		X"11",X"23",X"22",X"00",X"00",X"00",X"00",X"00",X"0C",X"38",X"58",X"70",X"30",X"00",X"00",X"00",
		X"F0",X"70",X"90",X"E0",X"80",X"00",X"00",X"00",X"0C",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"70",X"F0",X"30",X"10",X"00",X"11",X"33",X"F1",X"F0",X"FE",X"FE",X"F0",
		X"33",X"A8",X"C8",X"C8",X"E4",X"F4",X"F7",X"77",X"00",X"00",X"11",X"31",X"51",X"C0",X"C0",X"C0",
		X"10",X"31",X"F1",X"70",X"10",X"00",X"00",X"00",X"FC",X"FE",X"FE",X"FC",X"F1",X"33",X"11",X"00",
		X"77",X"F7",X"F4",X"E4",X"C8",X"C8",X"A8",X"33",X"C0",X"C0",X"C0",X"51",X"31",X"11",X"00",X"00",
		X"00",X"00",X"71",X"D9",X"77",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"88",X"CC",X"DE",X"FC",X"DF",X"FD",X"00",X"00",X"00",X"C0",X"20",X"A8",X"F9",X"F9",
		X"FF",X"77",X"77",X"33",X"11",X"00",X"00",X"00",X"F7",X"FB",X"FC",X"FF",X"FF",X"F0",X"00",X"00",
		X"DF",X"F8",X"D6",X"D8",X"80",X"00",X"00",X"00",X"F1",X"F1",X"E0",X"E0",X"40",X"00",X"00",X"00",
		X"0F",X"00",X"00",X"00",X"00",X"10",X"F0",X"50",X"0E",X"01",X"00",X"00",X"11",X"F3",X"F1",X"FE",
		X"00",X"0E",X"45",X"40",X"40",X"C8",X"E8",X"F4",X"00",X"00",X"0C",X"03",X"22",X"E2",X"A2",X"80",
		X"30",X"10",X"10",X"30",X"50",X"F0",X"10",X"00",X"FE",X"F0",X"F0",X"FE",X"FE",X"F1",X"F3",X"11",
		X"F0",X"90",X"90",X"F0",X"F4",X"E8",X"C8",X"71",X"80",X"88",X"88",X"80",X"80",X"A2",X"E2",X"22",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0E",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"03",X"11",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"77",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DD",
		X"00",X"00",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"EE",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",
		X"00",X"22",X"33",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"BB",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DD",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"CC",X"22",X"00",X"00",X"00",X"00",
		X"00",X"00",X"44",X"88",X"00",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"DD",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"22",X"11",X"00",X"00",X"00",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"10",X"31",X"33",X"76",X"BC",X"60",X"E0",X"E6",X"EE",X"EE",X"E8",X"E0",X"E0",
		X"F0",X"00",X"30",X"20",X"11",X"33",X"33",X"77",X"F0",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FD",
		X"76",X"33",X"31",X"10",X"10",X"00",X"00",X"00",X"E0",X"E8",X"EE",X"EE",X"E6",X"E0",X"60",X"00",
		X"77",X"77",X"77",X"77",X"33",X"33",X"11",X"00",X"FD",X"FE",X"33",X"BB",X"FF",X"FF",X"FC",X"60",
		X"31",X"20",X"71",X"E0",X"71",X"70",X"30",X"10",X"00",X"00",X"00",X"00",X"00",X"11",X"80",X"F3",
		X"00",X"CC",X"66",X"EE",X"44",X"CC",X"CC",X"EE",X"00",X"00",X"00",X"00",X"CC",X"66",X"40",X"40",
		X"31",X"30",X"F0",X"73",X"30",X"00",X"00",X"00",X"FF",X"FC",X"F0",X"F0",X"F0",X"F0",X"30",X"00",
		X"FF",X"FF",X"F7",X"F0",X"F0",X"A0",X"20",X"22",X"C8",X"C8",X"C0",X"C0",X"A0",X"20",X"31",X"33",
		X"10",X"10",X"30",X"70",X"70",X"30",X"30",X"10",X"88",X"11",X"88",X"11",X"88",X"33",X"91",X"F3",
		X"00",X"88",X"CC",X"CC",X"88",X"88",X"88",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"31",X"31",X"30",X"71",X"F0",X"00",X"00",X"00",X"FF",X"FE",X"F0",X"F0",X"F0",X"F0",X"30",X"00",
		X"FF",X"CC",X"F0",X"C0",X"F0",X"80",X"00",X"00",X"99",X"55",X"F9",X"51",X"80",X"00",X"00",X"00",
		X"00",X"00",X"10",X"30",X"30",X"30",X"10",X"10",X"C4",X"91",X"C4",X"90",X"D5",X"91",X"D1",X"F3",
		X"00",X"88",X"CC",X"CC",X"88",X"AA",X"A8",X"EC",X"00",X"00",X"00",X"00",X"CC",X"66",X"40",X"40",
		X"30",X"31",X"F0",X"73",X"30",X"00",X"00",X"00",X"FD",X"FE",X"F0",X"F0",X"F0",X"F0",X"30",X"00",
		X"FD",X"FD",X"F0",X"F0",X"F0",X"80",X"00",X"00",X"88",X"CC",X"CC",X"E0",X"A0",X"20",X"31",X"33",
		X"00",X"0F",X"00",X"00",X"00",X"10",X"70",X"F2",X"00",X"0E",X"01",X"00",X"11",X"F3",X"F1",X"FE",
		X"00",X"00",X"0E",X"81",X"C0",X"E8",X"FC",X"F4",X"00",X"00",X"00",X"0C",X"03",X"71",X"51",X"C0",
		X"30",X"10",X"10",X"30",X"F2",X"70",X"10",X"00",X"FE",X"F0",X"F0",X"FE",X"FE",X"F1",X"F3",X"11",
		X"F0",X"90",X"90",X"F0",X"F4",X"EC",X"B8",X"00",X"C0",X"C4",X"C4",X"C0",X"C0",X"51",X"F9",X"11",
		X"31",X"20",X"71",X"E0",X"71",X"70",X"30",X"10",X"00",X"0F",X"00",X"00",X"00",X"11",X"80",X"F3",
		X"00",X"CC",X"67",X"EE",X"44",X"CC",X"CC",X"EE",X"00",X"00",X"08",X"07",X"CC",X"66",X"40",X"40",
		X"31",X"30",X"F0",X"73",X"30",X"00",X"00",X"00",X"FD",X"FC",X"F0",X"F0",X"F0",X"F0",X"30",X"00",
		X"FF",X"FF",X"F7",X"F0",X"F0",X"A0",X"20",X"22",X"C8",X"C8",X"C0",X"C0",X"A0",X"20",X"31",X"33",
		X"18",X"10",X"30",X"70",X"70",X"30",X"30",X"10",X"88",X"15",X"8B",X"11",X"88",X"33",X"91",X"F3",
		X"00",X"88",X"CC",X"CC",X"9E",X"A8",X"A8",X"EC",X"00",X"00",X"00",X"00",X"00",X"0C",X"03",X"00",
		X"31",X"31",X"30",X"71",X"F0",X"00",X"00",X"00",X"FF",X"FE",X"FC",X"E0",X"D0",X"E2",X"30",X"00",
		X"FF",X"FC",X"70",X"F0",X"70",X"80",X"00",X"00",X"99",X"D5",X"F1",X"D1",X"80",X"00",X"00",X"00",
		X"00",X"00",X"11",X"33",X"72",X"F2",X"74",X"FC",X"00",X"00",X"CC",X"FF",X"F1",X"FC",X"FC",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"DC",X"F2",X"90",X"00",X"00",X"00",X"D1",X"31",X"D1",X"C0",X"C0",
		X"FC",X"74",X"F2",X"72",X"33",X"11",X"00",X"00",X"F0",X"FC",X"FC",X"F1",X"FF",X"CC",X"00",X"00",
		X"90",X"F2",X"DC",X"00",X"00",X"00",X"00",X"00",X"C0",X"D1",X"71",X"11",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"11",X"00",X"30",X"73",X"F0",X"31",X"31",X"F0",X"20",X"F0",X"F0",X"F0",X"F0",X"FE",X"FF",
		X"80",X"C0",X"40",X"F0",X"F0",X"F0",X"F8",X"FC",X"00",X"22",X"E2",X"A2",X"80",X"80",X"11",X"B3",
		X"10",X"10",X"30",X"30",X"30",X"10",X"10",X"00",X"C0",X"91",X"C4",X"00",X"88",X"00",X"88",X"00",
		X"FC",X"FE",X"66",X"FF",X"33",X"66",X"00",X"00",X"EE",X"80",X"D1",X"31",X"11",X"00",X"00",X"00",
		X"73",X"F0",X"30",X"10",X"00",X"00",X"00",X"00",X"F0",X"F0",X"FF",X"FF",X"F1",X"E0",X"F1",X"E0",
		X"F0",X"F0",X"E6",X"EE",X"CC",X"CC",X"CC",X"66",X"D1",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F1",X"E2",X"51",X"62",X"00",X"00",X"00",X"00",
		X"EE",X"CC",X"CC",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"30",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"40",X"20",X"30",X"90",X"40",X"30",X"03",X"00",X"40",X"20",X"20",X"2C",X"4B",X"7A",X"78",
		X"40",X"90",X"E0",X"80",X"B0",X"E0",X"8F",X"C2",X"00",X"C0",X"40",X"80",X"20",X"40",X"80",X"00",
		X"80",X"50",X"21",X"40",X"10",X"20",X"40",X"80",X"3F",X"1A",X"38",X"0B",X"10",X"20",X"40",X"00",
		X"CB",X"E4",X"61",X"50",X"40",X"20",X"10",X"80",X"C0",X"20",X"90",X"08",X"C0",X"60",X"00",X"00",
		X"00",X"60",X"F0",X"70",X"40",X"40",X"00",X"00",X"00",X"00",X"80",X"E0",X"80",X"20",X"A0",X"43",
		X"00",X"10",X"30",X"40",X"00",X"40",X"80",X"08",X"00",X"00",X"00",X"80",X"40",X"E0",X"00",X"00",
		X"00",X"00",X"40",X"D0",X"F0",X"70",X"10",X"00",X"43",X"A1",X"20",X"00",X"20",X"E0",X"E0",X"00",
		X"48",X"20",X"00",X"20",X"30",X"00",X"00",X"00",X"00",X"20",X"60",X"E0",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"20",X"70",X"F0",X"60",X"20",X"00",X"00",
		X"00",X"00",X"80",X"00",X"80",X"40",X"00",X"00",X"00",X"00",X"00",X"40",X"C0",X"20",X"00",X"00",
		X"00",X"30",X"10",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"D0",X"F0",X"60",X"00",
		X"00",X"00",X"00",X"90",X"80",X"00",X"00",X"00",X"00",X"60",X"20",X"E0",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"60",X"60",X"00",
		X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"E0",X"70",X"00",X"00",X"00",
		X"10",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"0F",X"07",X"03",X"70",X"F0",
		X"99",X"FF",X"77",X"FF",X"FF",X"FF",X"FF",X"67",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"33",X"FF",X"FF",X"FB",X"F8",X"FC",X"00",X"00",X"88",X"EF",X"EF",X"88",X"CC",X"EF",
		X"77",X"33",X"11",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"70",X"00",X"00",X"00",X"00",
		X"F4",X"B8",X"10",X"10",X"11",X"11",X"33",X"33",X"EF",X"01",X"CC",X"EE",X"EE",X"CC",X"88",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"40",X"40",X"30",X"00",X"77",X"04",
		X"00",X"E0",X"10",X"10",X"E0",X"00",X"8E",X"89",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"47",X"00",X"00",X"34",X"20",X"00",X"00",
		X"89",X"7F",X"00",X"01",X"69",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"C3",X"E1",X"30",X"10",X"00",X"00",X"00",X"F0",X"F0",X"C3",X"5A",X"F0",X"F0",X"30",X"00",
		X"00",X"00",X"C0",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"08",X"08",X"07",X"00",X"07",X"08",
		X"00",X"0C",X"02",X"02",X"0C",X"00",X"0C",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"07",X"00",X"00",X"6F",X"44",X"02",X"11",
		X"02",X"0C",X"00",X"08",X"CE",X"88",X"08",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"88",X"77",X"00",X"77",X"88",X"77",X"00",
		X"CC",X"22",X"CC",X"00",X"CC",X"22",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"99",X"77",X"00",X"00",X"FF",X"44",X"00",
		X"CC",X"22",X"CC",X"00",X"22",X"EE",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"77",X"33",X"00",X"00",X"00",X"00",
		X"00",X"00",X"88",X"CC",X"EE",X"66",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"33",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"BB",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0C",X"78",X"34",
		X"00",X"00",X"00",X"0B",X"08",X"20",X"F0",X"F0",X"00",X"00",X"00",X"08",X"0C",X"06",X"02",X"83",
		X"00",X"00",X"08",X"08",X"0C",X"0E",X"87",X"E1",X"30",X"30",X"30",X"10",X"00",X"00",X"08",X"68",
		X"F0",X"F0",X"F0",X"F0",X"70",X"10",X"00",X"00",X"81",X"E1",X"F0",X"F0",X"E0",X"E0",X"E0",X"60");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
