library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_PGM_0 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_PGM_0 is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"F3",X"AF",X"06",X"08",X"21",X"00",X"50",X"77",X"23",X"10",X"FC",X"ED",X"56",X"31",X"F1",X"4F",
		X"C3",X"00",X"3F",X"3A",X"A6",X"4C",X"FE",X"00",X"C8",X"47",X"3E",X"18",X"21",X"1D",X"40",X"77",
		X"2B",X"10",X"FC",X"C9",X"3A",X"A7",X"4C",X"FE",X"00",X"C8",X"47",X"3E",X"18",X"21",X"02",X"40",
		X"77",X"23",X"10",X"FC",X"C9",X"D6",X"FF",X"00",X"08",X"D9",X"DD",X"E5",X"FD",X"E5",X"AF",X"32",
		X"00",X"50",X"2A",X"0C",X"4C",X"3A",X"0E",X"4C",X"77",X"2A",X"0F",X"4C",X"3A",X"11",X"4C",X"77",
		X"2A",X"14",X"4C",X"3A",X"16",X"4C",X"77",X"2A",X"17",X"4C",X"3A",X"19",X"4C",X"77",X"2A",X"1C",
		X"4C",X"3A",X"1E",X"4C",X"77",X"2A",X"1F",X"4C",X"3A",X"21",X"4C",X"77",X"2A",X"24",X"4C",X"3A",
		X"26",X"4C",X"77",X"2A",X"27",X"4C",X"3A",X"29",X"4C",X"77",X"2A",X"2C",X"4C",X"3A",X"2E",X"4C",
		X"77",X"2A",X"2F",X"4C",X"3A",X"31",X"4C",X"77",X"2A",X"34",X"4C",X"3A",X"36",X"4C",X"77",X"2A",
		X"37",X"4C",X"3A",X"39",X"4C",X"77",X"2A",X"3C",X"4C",X"3A",X"3E",X"4C",X"77",X"2A",X"3F",X"4C",
		X"3A",X"41",X"4C",X"77",X"2A",X"44",X"4C",X"3A",X"46",X"4C",X"77",X"2A",X"47",X"4C",X"3A",X"49",
		X"4C",X"77",X"2A",X"4C",X"4C",X"3A",X"4E",X"4C",X"77",X"2A",X"4F",X"4C",X"3A",X"51",X"4C",X"77",
		X"2A",X"54",X"4C",X"3A",X"56",X"4C",X"77",X"2A",X"57",X"4C",X"3A",X"59",X"4C",X"77",X"21",X"96",
		X"4C",X"CB",X"7E",X"28",X"31",X"CB",X"6E",X"20",X"2D",X"06",X"06",X"21",X"64",X"4C",X"11",X"62",
		X"50",X"3E",X"06",X"0E",X"02",X"ED",X"A0",X"ED",X"A0",X"CD",X"BA",X"15",X"10",X"F3",X"06",X"06",
		X"21",X"66",X"4C",X"11",X"F2",X"4F",X"3E",X"06",X"0E",X"02",X"ED",X"A0",X"ED",X"A0",X"CD",X"BA",
		X"15",X"10",X"F3",X"C3",X"7E",X"01",X"ED",X"5B",X"64",X"4C",X"CD",X"3D",X"0F",X"ED",X"53",X"62",
		X"50",X"ED",X"5B",X"6C",X"4C",X"CD",X"3D",X"0F",X"ED",X"53",X"64",X"50",X"ED",X"5B",X"74",X"4C",
		X"CD",X"3D",X"0F",X"ED",X"53",X"66",X"50",X"ED",X"5B",X"7C",X"4C",X"CD",X"3D",X"0F",X"ED",X"53",
		X"68",X"50",X"ED",X"5B",X"84",X"4C",X"CD",X"3D",X"0F",X"ED",X"53",X"6A",X"50",X"ED",X"5B",X"8C",
		X"4C",X"CD",X"3D",X"0F",X"ED",X"53",X"6C",X"50",X"2A",X"66",X"4C",X"CD",X"56",X"0F",X"22",X"F2",
		X"4F",X"2A",X"6E",X"4C",X"CD",X"56",X"0F",X"22",X"F4",X"4F",X"2A",X"76",X"4C",X"CD",X"56",X"0F",
		X"22",X"F6",X"4F",X"2A",X"7E",X"4C",X"CD",X"56",X"0F",X"22",X"F8",X"4F",X"2A",X"86",X"4C",X"CD",
		X"56",X"0F",X"22",X"FA",X"4F",X"2A",X"8E",X"4C",X"CD",X"56",X"0F",X"22",X"FC",X"4F",X"2A",X"93",
		X"4C",X"23",X"22",X"93",X"4C",X"7E",X"FE",X"FF",X"20",X"06",X"21",X"DB",X"3C",X"22",X"93",X"4C",
		X"21",X"95",X"4C",X"CB",X"46",X"20",X"56",X"3A",X"00",X"50",X"CB",X"6F",X"CA",X"2A",X"02",X"CB",
		X"8E",X"CB",X"56",X"20",X"3D",X"3A",X"00",X"50",X"CB",X"7F",X"CA",X"38",X"02",X"3A",X"98",X"4C",
		X"FE",X"06",X"28",X"07",X"3C",X"32",X"98",X"4C",X"C3",X"3D",X"02",X"AF",X"32",X"98",X"4C",X"CB",
		X"5E",X"20",X"0A",X"3A",X"99",X"4C",X"FE",X"00",X"20",X"0B",X"C3",X"3D",X"02",X"AF",X"32",X"07",
		X"50",X"CB",X"9E",X"18",X"68",X"3D",X"32",X"99",X"4C",X"3E",X"01",X"32",X"07",X"50",X"CB",X"DE",
		X"18",X"5B",X"3A",X"00",X"50",X"CB",X"7F",X"28",X"C4",X"CB",X"96",X"18",X"10",X"3A",X"00",X"50",
		X"CB",X"6F",X"28",X"AD",X"CB",X"86",X"3A",X"99",X"4C",X"3C",X"32",X"99",X"4C",X"3A",X"9A",X"4C",
		X"FE",X"14",X"30",X"1A",X"47",X"3A",X"9C",X"4C",X"80",X"32",X"9A",X"4C",X"CB",X"3F",X"06",X"00",
		X"80",X"27",X"32",X"9D",X"4C",X"CD",X"27",X"15",X"CB",X"66",X"20",X"02",X"CB",X"EE",X"3A",X"05",
		X"4D",X"CB",X"C7",X"32",X"05",X"4D",X"CB",X"F6",X"18",X"83",X"CB",X"4E",X"20",X"05",X"CB",X"CE",
		X"C3",X"A1",X"01",X"CB",X"C6",X"C3",X"9F",X"01",X"CB",X"D6",X"C3",X"AD",X"01",X"00",X"21",X"96",
		X"4C",X"CB",X"46",X"28",X"16",X"CD",X"49",X"16",X"21",X"96",X"4C",X"CB",X"7E",X"28",X"04",X"CB",
		X"6E",X"28",X"05",X"CD",X"29",X"16",X"18",X"03",X"CD",X"39",X"16",X"3A",X"9F",X"4C",X"3C",X"32",
		X"9F",X"4C",X"3A",X"9E",X"4C",X"3C",X"32",X"9E",X"4C",X"FE",X"3C",X"20",X"0B",X"AF",X"32",X"9E",
		X"4C",X"3A",X"A0",X"4C",X"3C",X"32",X"A0",X"4C",X"21",X"95",X"4C",X"CB",X"BE",X"3A",X"00",X"50",
		X"CB",X"77",X"20",X"35",X"AF",X"32",X"01",X"50",X"21",X"62",X"50",X"06",X"0C",X"36",X"00",X"23",
		X"10",X"FB",X"3E",X"40",X"CD",X"07",X"15",X"3E",X"09",X"CD",X"17",X"15",X"11",X"D0",X"41",X"21",
		X"9C",X"19",X"3E",X"01",X"06",X"04",X"CD",X"DF",X"15",X"06",X"FF",X"21",X"FF",X"FF",X"2B",X"7D",
		X"BC",X"32",X"C0",X"50",X"20",X"F8",X"10",X"F3",X"76",X"FB",X"3E",X"01",X"32",X"00",X"50",X"FD",
		X"E1",X"DD",X"E1",X"D9",X"08",X"ED",X"4D",X"3A",X"00",X"50",X"CB",X"67",X"C2",X"93",X"05",X"AF",
		X"06",X"08",X"21",X"00",X"50",X"77",X"23",X"10",X"FC",X"3E",X"00",X"32",X"03",X"50",X"31",X"F1",
		X"4F",X"CD",X"14",X"16",X"F3",X"08",X"AF",X"08",X"21",X"00",X"40",X"CD",X"16",X"05",X"08",X"CB",
		X"47",X"28",X"02",X"CB",X"D7",X"CB",X"4F",X"28",X"02",X"CB",X"DF",X"08",X"21",X"00",X"44",X"CD",
		X"16",X"05",X"08",X"CB",X"47",X"28",X"02",X"CB",X"E7",X"CB",X"4F",X"28",X"02",X"CB",X"EF",X"08",
		X"31",X"FD",X"43",X"21",X"00",X"4C",X"CD",X"16",X"05",X"08",X"CB",X"47",X"28",X"02",X"CB",X"F7",
		X"CB",X"4F",X"28",X"02",X"CB",X"FF",X"08",X"3E",X"01",X"CD",X"17",X"15",X"21",X"00",X"40",X"11",
		X"01",X"40",X"01",X"FE",X"03",X"36",X"40",X"ED",X"B0",X"11",X"66",X"41",X"21",X"60",X"1A",X"3E",
		X"01",X"06",X"0B",X"CD",X"DF",X"15",X"11",X"8A",X"40",X"21",X"6B",X"1A",X"3E",X"01",X"06",X"18",
		X"CD",X"DF",X"15",X"11",X"EC",X"40",X"21",X"83",X"1A",X"3E",X"01",X"06",X"14",X"CD",X"DF",X"15",
		X"11",X"ED",X"40",X"21",X"97",X"1A",X"3E",X"01",X"06",X"14",X"CD",X"DF",X"15",X"11",X"EE",X"40",
		X"21",X"AB",X"1A",X"3E",X"01",X"06",X"14",X"CD",X"DF",X"15",X"11",X"EF",X"40",X"21",X"BF",X"1A",
		X"3E",X"01",X"06",X"14",X"CD",X"DF",X"15",X"11",X"93",X"40",X"21",X"4F",X"1B",X"3E",X"01",X"06",
		X"18",X"CD",X"DF",X"15",X"11",X"F5",X"40",X"21",X"D3",X"1A",X"3E",X"01",X"06",X"14",X"CD",X"DF",
		X"15",X"11",X"F6",X"40",X"21",X"E7",X"1A",X"3E",X"01",X"06",X"14",X"CD",X"DF",X"15",X"11",X"F7",
		X"40",X"21",X"FB",X"1A",X"3E",X"01",X"06",X"14",X"CD",X"DF",X"15",X"11",X"F8",X"40",X"21",X"0F",
		X"1B",X"3E",X"01",X"06",X"14",X"CD",X"DF",X"15",X"11",X"F9",X"40",X"21",X"23",X"1B",X"3E",X"01",
		X"06",X"14",X"CD",X"DF",X"15",X"11",X"FA",X"40",X"21",X"37",X"1B",X"3E",X"01",X"06",X"14",X"CD",
		X"DF",X"15",X"08",X"32",X"FE",X"4C",X"08",X"3A",X"FE",X"4C",X"CB",X"57",X"28",X"0D",X"11",X"F5",
		X"40",X"21",X"4B",X"1B",X"3E",X"01",X"06",X"04",X"CD",X"DF",X"15",X"3A",X"FE",X"4C",X"CB",X"5F",
		X"28",X"0D",X"11",X"F6",X"40",X"21",X"4B",X"1B",X"3E",X"01",X"06",X"04",X"CD",X"DF",X"15",X"3A",
		X"FE",X"4C",X"CB",X"67",X"28",X"0D",X"11",X"F7",X"40",X"21",X"4B",X"1B",X"3E",X"01",X"06",X"04",
		X"CD",X"DF",X"15",X"3A",X"FE",X"4C",X"CB",X"6F",X"28",X"0D",X"11",X"F8",X"40",X"21",X"4B",X"1B",
		X"3E",X"01",X"06",X"04",X"CD",X"DF",X"15",X"3A",X"FE",X"4C",X"CB",X"77",X"28",X"0D",X"11",X"F9",
		X"40",X"21",X"4B",X"1B",X"3E",X"01",X"06",X"04",X"CD",X"DF",X"15",X"3A",X"FE",X"4C",X"CB",X"7F",
		X"28",X"0D",X"11",X"FA",X"40",X"21",X"4B",X"1B",X"3E",X"01",X"06",X"04",X"CD",X"DF",X"15",X"1E",
		X"00",X"21",X"00",X"00",X"CD",X"FD",X"04",X"30",X"02",X"CB",X"C3",X"21",X"00",X"10",X"CD",X"FD",
		X"04",X"30",X"02",X"CB",X"CB",X"21",X"00",X"20",X"CD",X"FD",X"04",X"30",X"02",X"CB",X"D3",X"21",
		X"00",X"30",X"CD",X"FD",X"04",X"30",X"02",X"CB",X"DB",X"3A",X"FE",X"4C",X"FE",X"00",X"28",X"02",
		X"3E",X"80",X"B3",X"32",X"FE",X"4C",X"CB",X"47",X"28",X"0D",X"11",X"EC",X"40",X"21",X"4B",X"1B",
		X"3E",X"01",X"06",X"04",X"CD",X"DF",X"15",X"3A",X"FE",X"4C",X"CB",X"4F",X"28",X"0D",X"11",X"ED",
		X"40",X"21",X"4B",X"1B",X"3E",X"01",X"06",X"04",X"CD",X"DF",X"15",X"3A",X"FE",X"4C",X"CB",X"57",
		X"28",X"0D",X"11",X"EE",X"40",X"21",X"4B",X"1B",X"3E",X"01",X"06",X"04",X"CD",X"DF",X"15",X"3A",
		X"FE",X"4C",X"CB",X"5F",X"28",X"0D",X"11",X"EF",X"40",X"21",X"4B",X"1B",X"3E",X"01",X"06",X"04",
		X"CD",X"DF",X"15",X"3A",X"FE",X"4C",X"FE",X"00",X"20",X"0E",X"FB",X"3E",X"01",X"32",X"00",X"50",
		X"3E",X"02",X"CD",X"59",X"15",X"C3",X"D9",X"02",X"32",X"C0",X"50",X"18",X"FB",X"01",X"00",X"10",
		X"AF",X"32",X"C0",X"50",X"86",X"23",X"57",X"0B",X"79",X"B0",X"7A",X"20",X"F7",X"FE",X"FF",X"28",
		X"02",X"37",X"C9",X"37",X"3F",X"C9",X"08",X"E6",X"FC",X"08",X"E5",X"3E",X"11",X"CD",X"35",X"05",
		X"E1",X"E5",X"3E",X"22",X"CD",X"35",X"05",X"E1",X"E5",X"3E",X"44",X"CD",X"35",X"05",X"E1",X"3E",
		X"88",X"CD",X"35",X"05",X"C9",X"32",X"C0",X"50",X"E5",X"E5",X"D1",X"13",X"01",X"FF",X"03",X"77",
		X"ED",X"B0",X"E1",X"01",X"00",X"04",X"BE",X"C4",X"53",X"05",X"23",X"5F",X"0B",X"79",X"B0",X"7B",
		X"20",X"F4",X"C9",X"5F",X"7E",X"E6",X"0F",X"57",X"7B",X"E6",X"0F",X"BA",X"28",X"04",X"08",X"CB",
		X"CF",X"08",X"7E",X"E6",X"F0",X"57",X"7B",X"E6",X"F0",X"BA",X"C8",X"08",X"CB",X"C7",X"08",X"7B",
		X"C9",X"47",X"4F",X"52",X"4B",X"41",X"4E",X"53",X"2C",X"43",X"4F",X"50",X"59",X"52",X"49",X"47",
		X"48",X"54",X"20",X"31",X"39",X"38",X"33",X"54",X"45",X"43",X"48",X"53",X"54",X"41",X"52",X"20",
		X"49",X"4E",X"43",X"32",X"C0",X"50",X"21",X"00",X"40",X"11",X"01",X"40",X"01",X"FE",X"07",X"36",
		X"40",X"ED",X"B0",X"32",X"C0",X"50",X"21",X"00",X"4C",X"11",X"01",X"4C",X"01",X"FE",X"03",X"36",
		X"00",X"ED",X"B0",X"32",X"C0",X"50",X"21",X"60",X"50",X"11",X"61",X"50",X"01",X"0F",X"00",X"36",
		X"00",X"ED",X"B0",X"32",X"C0",X"50",X"21",X"F0",X"4F",X"11",X"F1",X"4F",X"01",X"0F",X"00",X"36",
		X"00",X"ED",X"B0",X"32",X"C0",X"50",X"21",X"40",X"50",X"11",X"41",X"50",X"01",X"1F",X"00",X"36",
		X"00",X"ED",X"B0",X"21",X"0C",X"4C",X"11",X"0D",X"4C",X"01",X"4F",X"00",X"36",X"FF",X"ED",X"B0",
		X"21",X"DB",X"3C",X"22",X"93",X"4C",X"3A",X"80",X"50",X"47",X"E6",X"03",X"32",X"9B",X"4C",X"21",
		X"A5",X"1B",X"CD",X"BA",X"15",X"7E",X"32",X"9C",X"4C",X"78",X"E6",X"0C",X"CB",X"3F",X"CB",X"3F",
		X"21",X"D7",X"3C",X"CD",X"BA",X"15",X"7E",X"32",X"A2",X"4C",X"78",X"E6",X"30",X"21",X"97",X"3C",
		X"CD",X"BA",X"15",X"22",X"A3",X"4C",X"78",X"E6",X"30",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",
		X"3F",X"32",X"A5",X"4C",X"78",X"CB",X"77",X"20",X"05",X"21",X"96",X"4C",X"CB",X"FE",X"FB",X"3E",
		X"01",X"32",X"00",X"50",X"CD",X"9A",X"38",X"21",X"C2",X"43",X"11",X"C3",X"43",X"01",X"3C",X"00",
		X"36",X"40",X"ED",X"B0",X"21",X"C2",X"47",X"11",X"C3",X"47",X"01",X"1C",X"00",X"36",X"05",X"ED",
		X"B0",X"32",X"C0",X"50",X"21",X"E2",X"47",X"11",X"E3",X"47",X"01",X"1C",X"00",X"36",X"09",X"ED",
		X"B0",X"32",X"C0",X"50",X"21",X"95",X"18",X"11",X"C3",X"43",X"01",X"1A",X"00",X"ED",X"B0",X"AF",
		X"32",X"E4",X"43",X"32",X"ED",X"43",X"32",X"F6",X"43",X"21",X"F0",X"3C",X"11",X"B3",X"4C",X"01",
		X"3C",X"00",X"ED",X"B0",X"21",X"B8",X"4C",X"11",X"F2",X"43",X"CD",X"1B",X"10",X"21",X"02",X"40",
		X"11",X"03",X"40",X"01",X"3C",X"00",X"36",X"40",X"ED",X"B0",X"32",X"C0",X"50",X"21",X"02",X"44",
		X"11",X"03",X"44",X"01",X"1C",X"00",X"36",X"01",X"ED",X"B0",X"21",X"22",X"44",X"11",X"23",X"44",
		X"01",X"1C",X"00",X"36",X"11",X"ED",X"B0",X"32",X"C0",X"50",X"21",X"AF",X"18",X"11",X"0F",X"40",
		X"01",X"06",X"00",X"ED",X"B0",X"AF",X"32",X"0C",X"40",X"3A",X"9B",X"4C",X"FE",X"00",X"20",X"0B",
		X"21",X"B5",X"18",X"11",X"0C",X"40",X"01",X"09",X"00",X"ED",X"B0",X"32",X"C0",X"50",X"21",X"05",
		X"4D",X"11",X"06",X"4D",X"01",X"FF",X"00",X"36",X"00",X"ED",X"B0",X"21",X"FE",X"39",X"22",X"1E",
		X"4D",X"22",X"06",X"4D",X"21",X"1D",X"4D",X"22",X"0D",X"4D",X"21",X"2C",X"3A",X"22",X"39",X"4D",
		X"22",X"21",X"4D",X"21",X"38",X"4D",X"22",X"28",X"4D",X"21",X"43",X"3A",X"22",X"54",X"4D",X"22",
		X"3C",X"4D",X"21",X"53",X"4D",X"22",X"43",X"4D",X"21",X"66",X"3A",X"22",X"6F",X"4D",X"22",X"57",
		X"4D",X"21",X"6E",X"4D",X"22",X"5E",X"4D",X"21",X"92",X"3A",X"22",X"8A",X"4D",X"22",X"72",X"4D",
		X"21",X"89",X"4D",X"22",X"79",X"4D",X"21",X"AB",X"3A",X"22",X"A5",X"4D",X"22",X"8D",X"4D",X"21",
		X"A4",X"4D",X"22",X"94",X"4D",X"21",X"C4",X"3A",X"22",X"C0",X"4D",X"22",X"A8",X"4D",X"21",X"BF",
		X"4D",X"22",X"AF",X"4D",X"21",X"DD",X"3A",X"22",X"DB",X"4D",X"22",X"C3",X"4D",X"21",X"DA",X"4D",
		X"22",X"CA",X"4D",X"06",X"20",X"21",X"40",X"50",X"36",X"00",X"23",X"10",X"FB",X"3E",X"00",X"32",
		X"03",X"50",X"21",X"96",X"4C",X"CB",X"EE",X"3A",X"9B",X"4C",X"FE",X"00",X"CA",X"38",X"09",X"3A",
		X"9A",X"4C",X"FE",X"00",X"C2",X"38",X"09",X"21",X"95",X"4C",X"CB",X"A6",X"AF",X"32",X"01",X"50",
		X"21",X"96",X"4C",X"CB",X"86",X"CD",X"14",X"16",X"32",X"C0",X"50",X"CD",X"DC",X"35",X"21",X"95",
		X"4C",X"CB",X"6E",X"C2",X"38",X"09",X"CD",X"71",X"10",X"3E",X"07",X"CD",X"59",X"15",X"21",X"95",
		X"4C",X"CB",X"6E",X"C2",X"38",X"09",X"3E",X"40",X"CD",X"07",X"15",X"11",X"44",X"44",X"21",X"2C",
		X"3D",X"3E",X"01",X"06",X"1C",X"CD",X"F5",X"15",X"11",X"49",X"44",X"21",X"2E",X"3D",X"3E",X"03",
		X"06",X"1C",X"CD",X"F5",X"15",X"11",X"50",X"44",X"21",X"2D",X"3D",X"3E",X"03",X"06",X"1C",X"CD",
		X"F5",X"15",X"11",X"58",X"44",X"21",X"2E",X"3D",X"3E",X"03",X"06",X"1C",X"CD",X"F5",X"15",X"11",
		X"5B",X"44",X"21",X"2F",X"3D",X"3E",X"03",X"06",X"1C",X"CD",X"F5",X"15",X"11",X"C4",X"40",X"21",
		X"A0",X"19",X"3E",X"01",X"06",X"15",X"CD",X"DF",X"15",X"11",X"C9",X"40",X"21",X"B5",X"19",X"3E",
		X"01",X"06",X"14",X"CD",X"DF",X"15",X"11",X"AB",X"40",X"21",X"C9",X"19",X"3E",X"01",X"06",X"17",
		X"CD",X"DF",X"15",X"11",X"B0",X"40",X"21",X"E0",X"19",X"3E",X"01",X"06",X"16",X"CD",X"DF",X"15",
		X"11",X"52",X"41",X"21",X"F6",X"19",X"3E",X"01",X"06",X"0C",X"CD",X"DF",X"15",X"3A",X"9B",X"4C",
		X"FE",X"01",X"20",X"0F",X"11",X"19",X"41",X"21",X"02",X"1A",X"3E",X"01",X"06",X"0F",X"CD",X"DF",
		X"15",X"18",X"20",X"FE",X"02",X"20",X"0F",X"11",X"19",X"41",X"21",X"11",X"1A",X"3E",X"01",X"06",
		X"0F",X"CD",X"DF",X"15",X"18",X"0D",X"11",X"19",X"41",X"21",X"20",X"1A",X"3E",X"01",X"06",X"0F",
		X"CD",X"DF",X"15",X"11",X"9C",X"40",X"21",X"2F",X"1A",X"3E",X"01",X"06",X"19",X"CD",X"DF",X"15",
		X"3A",X"A5",X"4C",X"FE",X"00",X"20",X"0F",X"11",X"7C",X"41",X"21",X"48",X"1A",X"3E",X"01",X"06",
		X"06",X"CD",X"DF",X"15",X"18",X"33",X"FE",X"01",X"20",X"0F",X"11",X"7C",X"41",X"21",X"4E",X"1A",
		X"3E",X"01",X"06",X"06",X"CD",X"DF",X"15",X"18",X"20",X"FE",X"02",X"20",X"0F",X"11",X"7C",X"41",
		X"21",X"54",X"1A",X"3E",X"01",X"06",X"06",X"CD",X"DF",X"15",X"18",X"0D",X"11",X"7C",X"41",X"21",
		X"5A",X"1A",X"3E",X"01",X"06",X"06",X"CD",X"DF",X"15",X"3E",X"08",X"CD",X"59",X"15",X"21",X"95",
		X"4C",X"CB",X"6E",X"20",X"53",X"CD",X"9B",X"38",X"AF",X"32",X"FF",X"4C",X"32",X"01",X"4D",X"32",
		X"03",X"4D",X"32",X"00",X"4D",X"32",X"02",X"4D",X"32",X"04",X"4D",X"CD",X"BD",X"38",X"CD",X"EF",
		X"0E",X"CD",X"CA",X"38",X"CD",X"C5",X"1B",X"AF",X"32",X"20",X"4D",X"32",X"3B",X"4D",X"32",X"56",
		X"4D",X"32",X"71",X"4D",X"32",X"8C",X"4D",X"32",X"A7",X"4D",X"32",X"C2",X"4D",X"CD",X"1F",X"16",
		X"32",X"C0",X"50",X"21",X"95",X"4C",X"CB",X"6E",X"20",X"0E",X"21",X"96",X"4C",X"CB",X"4E",X"20",
		X"02",X"18",X"CE",X"CB",X"8E",X"C3",X"A5",X"07",X"CD",X"14",X"16",X"21",X"95",X"4C",X"CB",X"E6",
		X"CB",X"AE",X"21",X"96",X"4C",X"CB",X"8E",X"CB",X"96",X"CB",X"9E",X"21",X"97",X"4C",X"CB",X"96",
		X"21",X"96",X"4C",X"CB",X"C6",X"21",X"0C",X"4C",X"11",X"0D",X"4C",X"01",X"4F",X"00",X"36",X"FF",
		X"ED",X"B0",X"3E",X"FF",X"32",X"01",X"50",X"21",X"97",X"4C",X"CB",X"56",X"20",X"0F",X"3A",X"FD",
		X"4C",X"3C",X"32",X"FD",X"4C",X"FE",X"0A",X"20",X"04",X"CB",X"D6",X"CB",X"DE",X"00",X"32",X"C0",
		X"50",X"3E",X"40",X"CD",X"07",X"15",X"3E",X"03",X"CD",X"17",X"15",X"3A",X"9B",X"4C",X"FE",X"00",
		X"CA",X"13",X"0A",X"3A",X"9A",X"4C",X"FE",X"02",X"30",X"4C",X"11",X"70",X"41",X"21",X"BE",X"18",
		X"3E",X"01",X"06",X"0B",X"CD",X"DF",X"15",X"3A",X"40",X"50",X"CB",X"6F",X"20",X"74",X"3A",X"9B",
		X"4C",X"FE",X"00",X"28",X"15",X"3A",X"9A",X"4C",X"FE",X"02",X"38",X"66",X"D6",X"02",X"32",X"9A",
		X"4C",X"3A",X"9D",X"4C",X"D6",X"01",X"27",X"32",X"9D",X"4C",X"21",X"96",X"4C",X"CB",X"E6",X"3A",
		X"A2",X"4C",X"32",X"A6",X"4C",X"CD",X"13",X"00",X"3A",X"9B",X"4C",X"FE",X"00",X"CA",X"6E",X"0A",
		X"CD",X"27",X"15",X"C3",X"6E",X"0A",X"FE",X"04",X"30",X"29",X"11",X"0E",X"41",X"21",X"C9",X"18",
		X"3E",X"01",X"06",X"11",X"CD",X"DF",X"15",X"11",X"10",X"42",X"21",X"DA",X"18",X"3E",X"01",X"06",
		X"02",X"CD",X"DF",X"15",X"11",X"72",X"41",X"21",X"BE",X"18",X"3E",X"01",X"06",X"0B",X"CD",X"DF",
		X"15",X"18",X"94",X"11",X"90",X"40",X"21",X"DC",X"18",X"3E",X"01",X"06",X"19",X"CD",X"DF",X"15",
		X"18",X"85",X"3A",X"40",X"50",X"CB",X"77",X"20",X"33",X"3A",X"9B",X"4C",X"FE",X"00",X"28",X"15",
		X"3A",X"9A",X"4C",X"FE",X"04",X"38",X"25",X"D6",X"04",X"32",X"9A",X"4C",X"3A",X"9D",X"4C",X"D6",
		X"02",X"27",X"32",X"9D",X"4C",X"21",X"96",X"4C",X"CB",X"A6",X"3A",X"A2",X"4C",X"32",X"A6",X"4C",
		X"32",X"A7",X"4C",X"CD",X"13",X"00",X"CD",X"24",X"00",X"C3",X"D8",X"09",X"32",X"C0",X"50",X"21",
		X"95",X"4C",X"CB",X"76",X"20",X"03",X"C3",X"A7",X"09",X"CB",X"B6",X"C3",X"7E",X"09",X"AF",X"21",
		X"A8",X"4C",X"11",X"A9",X"4C",X"01",X"05",X"00",X"77",X"ED",X"B0",X"32",X"B1",X"4C",X"32",X"B2",
		X"4C",X"3E",X"40",X"21",X"E4",X"43",X"11",X"E5",X"43",X"01",X"05",X"00",X"77",X"ED",X"B0",X"21",
		X"F6",X"43",X"11",X"F7",X"43",X"01",X"05",X"00",X"77",X"ED",X"B0",X"AF",X"32",X"E4",X"43",X"32",
		X"F6",X"43",X"AF",X"32",X"FF",X"4C",X"32",X"01",X"4D",X"32",X"03",X"4D",X"32",X"00",X"4D",X"32",
		X"02",X"4D",X"32",X"04",X"4D",X"CD",X"AC",X"38",X"CD",X"C9",X"38",X"21",X"97",X"4C",X"CB",X"CE",
		X"21",X"96",X"4C",X"CB",X"66",X"28",X"02",X"18",X"1A",X"3E",X"00",X"32",X"03",X"50",X"CD",X"4E",
		X"15",X"11",X"50",X"41",X"21",X"F5",X"18",X"3E",X"01",X"06",X"0D",X"CD",X"DF",X"15",X"3E",X"03",
		X"CD",X"59",X"15",X"21",X"96",X"4C",X"CB",X"EE",X"3A",X"A6",X"4C",X"3D",X"32",X"A6",X"4C",X"3E",
		X"40",X"21",X"16",X"40",X"11",X"17",X"40",X"01",X"08",X"00",X"77",X"ED",X"B0",X"CD",X"13",X"00",
		X"3A",X"FF",X"4C",X"32",X"03",X"4D",X"3A",X"00",X"4D",X"32",X"04",X"4D",X"CD",X"09",X"39",X"C3",
		X"9A",X"0B",X"21",X"96",X"4C",X"CB",X"66",X"20",X"CA",X"CB",X"6E",X"28",X"AC",X"3A",X"96",X"4C",
		X"CB",X"7F",X"20",X"43",X"CD",X"4E",X"15",X"11",X"50",X"41",X"21",X"02",X"19",X"3E",X"01",X"06",
		X"0D",X"CD",X"DF",X"15",X"3E",X"03",X"CD",X"59",X"15",X"21",X"96",X"4C",X"CB",X"AE",X"3A",X"A7",
		X"4C",X"3D",X"32",X"A7",X"4C",X"3E",X"40",X"21",X"02",X"40",X"11",X"03",X"40",X"01",X"08",X"00",
		X"77",X"ED",X"B0",X"CD",X"24",X"00",X"3A",X"01",X"4D",X"32",X"03",X"4D",X"3A",X"02",X"4D",X"32",
		X"04",X"4D",X"CD",X"11",X"39",X"18",X"33",X"3E",X"01",X"32",X"03",X"50",X"18",X"B6",X"CD",X"4E",
		X"15",X"21",X"96",X"4C",X"CB",X"66",X"C2",X"E8",X"0A",X"11",X"10",X"41",X"21",X"0F",X"19",X"3E",
		X"01",X"06",X"11",X"CD",X"DF",X"15",X"21",X"20",X"4D",X"CB",X"C6",X"3E",X"01",X"CD",X"59",X"15",
		X"21",X"96",X"4C",X"CB",X"6E",X"28",X"A7",X"C3",X"E8",X"0A",X"CD",X"EF",X"0E",X"21",X"97",X"4C",
		X"CB",X"4E",X"28",X"13",X"CB",X"8E",X"21",X"C2",X"4D",X"CB",X"C6",X"32",X"C0",X"50",X"3A",X"C2",
		X"4D",X"FE",X"00",X"20",X"F6",X"18",X"05",X"3E",X"02",X"CD",X"59",X"15",X"CD",X"C5",X"1B",X"ED",
		X"5B",X"AE",X"4C",X"7B",X"B2",X"28",X"09",X"21",X"00",X"00",X"22",X"AE",X"4C",X"CD",X"5B",X"0F",
		X"32",X"C0",X"50",X"CD",X"1F",X"16",X"21",X"96",X"4C",X"CB",X"4E",X"28",X"DF",X"CB",X"8E",X"CD",
		X"14",X"16",X"21",X"96",X"4C",X"CB",X"56",X"20",X"0F",X"CD",X"1B",X"39",X"CD",X"14",X"16",X"21",
		X"96",X"4C",X"CB",X"5E",X"20",X"09",X"18",X"67",X"CB",X"96",X"CD",X"1A",X"39",X"18",X"EA",X"CB",
		X"9E",X"21",X"97",X"4C",X"CB",X"CE",X"21",X"96",X"4C",X"CB",X"6E",X"20",X"29",X"3A",X"01",X"4D",
		X"3C",X"FE",X"0C",X"20",X"02",X"3E",X"0B",X"32",X"01",X"4D",X"32",X"03",X"4D",X"3A",X"02",X"4D",
		X"3C",X"FE",X"19",X"20",X"02",X"3E",X"18",X"32",X"02",X"4D",X"32",X"04",X"4D",X"CD",X"1C",X"39",
		X"CD",X"19",X"39",X"C3",X"9A",X"0B",X"3A",X"FF",X"4C",X"3C",X"FE",X"0C",X"20",X"02",X"3E",X"0B",
		X"32",X"FF",X"4C",X"32",X"03",X"4D",X"3A",X"00",X"4D",X"3C",X"FE",X"19",X"20",X"02",X"3E",X"18",
		X"32",X"00",X"4D",X"32",X"04",X"4D",X"CD",X"1C",X"39",X"CD",X"18",X"39",X"C3",X"9A",X"0B",X"3A",
		X"B0",X"4C",X"FE",X"00",X"20",X"2E",X"21",X"96",X"4C",X"CB",X"6E",X"20",X"2F",X"3A",X"A7",X"4C",
		X"FE",X"00",X"20",X"4E",X"CD",X"4E",X"15",X"11",X"90",X"41",X"21",X"20",X"19",X"3E",X"01",X"06",
		X"09",X"CD",X"DF",X"15",X"3E",X"02",X"CD",X"59",X"15",X"CD",X"F8",X"11",X"21",X"95",X"4C",X"CB",
		X"F6",X"C3",X"7D",X"07",X"D6",X"01",X"32",X"B0",X"4C",X"C3",X"6E",X"0B",X"3A",X"A6",X"4C",X"FE",
		X"00",X"20",X"25",X"21",X"96",X"4C",X"CB",X"66",X"20",X"CA",X"CD",X"4E",X"15",X"11",X"F0",X"40",
		X"21",X"29",X"19",X"3E",X"01",X"06",X"14",X"CD",X"DF",X"15",X"3E",X"03",X"CD",X"59",X"15",X"C3",
		X"1D",X"0B",X"CD",X"10",X"39",X"C3",X"12",X"0B",X"CD",X"08",X"39",X"C3",X"12",X"0B",X"2A",X"91",
		X"4C",X"EB",X"DD",X"21",X"00",X"00",X"DD",X"19",X"DD",X"7E",X"01",X"DD",X"86",X"02",X"47",X"E6",
		X"0F",X"DD",X"77",X"02",X"CB",X"38",X"CB",X"38",X"CB",X"38",X"CB",X"38",X"DD",X"7E",X"00",X"21",
		X"FC",X"0C",X"CB",X"27",X"CD",X"BA",X"15",X"5E",X"23",X"56",X"EB",X"E9",X"08",X"0D",X"08",X"0D",
		X"09",X"0D",X"11",X"0D",X"19",X"0D",X"21",X"0D",X"C9",X"DD",X"7E",X"04",X"90",X"DD",X"77",X"04",
		X"C9",X"DD",X"7E",X"04",X"80",X"DD",X"77",X"04",X"C9",X"DD",X"7E",X"03",X"80",X"DD",X"77",X"03",
		X"C9",X"DD",X"7E",X"03",X"90",X"DD",X"77",X"03",X"C9",X"2A",X"5E",X"4C",X"EB",X"DD",X"21",X"00",
		X"00",X"DD",X"19",X"EB",X"01",X"00",X"4C",X"37",X"3F",X"ED",X"42",X"E5",X"DD",X"7E",X"00",X"21",
		X"4C",X"0D",X"CB",X"27",X"CD",X"BA",X"15",X"5E",X"23",X"56",X"EB",X"E9",X"1C",X"0E",X"58",X"0D",
		X"9B",X"0D",X"2B",X"0E",X"35",X"0E",X"48",X"0E",X"DD",X"7E",X"03",X"32",X"5C",X"4C",X"DD",X"7E",
		X"04",X"32",X"5D",X"4C",X"CD",X"B2",X"0E",X"DD",X"7E",X"06",X"12",X"3A",X"0A",X"4C",X"FE",X"00",
		X"20",X"17",X"3A",X"0B",X"4C",X"FE",X"00",X"20",X"17",X"C1",X"21",X"0C",X"4C",X"09",X"E5",X"D1",
		X"13",X"01",X"05",X"00",X"36",X"FF",X"ED",X"B0",X"C9",X"DD",X"7E",X"06",X"13",X"12",X"18",X"E9",
		X"DD",X"7E",X"06",X"21",X"20",X"00",X"19",X"EB",X"12",X"18",X"DE",X"CD",X"DA",X"0E",X"DD",X"7E",
		X"03",X"90",X"32",X"5C",X"4C",X"DD",X"7E",X"04",X"32",X"5D",X"4C",X"CD",X"B2",X"0E",X"3A",X"0A",
		X"4C",X"FE",X"00",X"28",X"32",X"3A",X"0A",X"4C",X"CB",X"27",X"DD",X"46",X"05",X"80",X"3D",X"C1",
		X"FD",X"21",X"0C",X"4C",X"FD",X"09",X"FD",X"73",X"00",X"FD",X"72",X"01",X"FD",X"77",X"02",X"3C",
		X"13",X"FD",X"73",X"03",X"FD",X"72",X"04",X"FD",X"77",X"05",X"3A",X"5C",X"4C",X"DD",X"77",X"03",
		X"3A",X"5D",X"4C",X"DD",X"77",X"04",X"C9",X"3A",X"0B",X"4C",X"FE",X"00",X"CA",X"51",X"0E",X"3A",
		X"0B",X"4C",X"CB",X"27",X"C6",X"0F",X"DD",X"46",X"05",X"80",X"C1",X"FD",X"21",X"0C",X"4C",X"FD",
		X"09",X"FD",X"73",X"00",X"FD",X"72",X"01",X"FD",X"77",X"02",X"3C",X"21",X"20",X"00",X"19",X"EB",
		X"FD",X"73",X"03",X"FD",X"72",X"04",X"FD",X"77",X"05",X"C3",X"DA",X"0D",X"DD",X"7E",X"03",X"32",
		X"5C",X"4C",X"DD",X"7E",X"04",X"32",X"5D",X"4C",X"C3",X"AB",X"0D",X"CD",X"DA",X"0E",X"DD",X"7E",
		X"03",X"80",X"C3",X"A2",X"0D",X"CD",X"DA",X"0E",X"DD",X"7E",X"04",X"90",X"32",X"5D",X"4C",X"DD",
		X"7E",X"03",X"32",X"5C",X"4C",X"C3",X"AB",X"0D",X"CD",X"DA",X"0E",X"DD",X"7E",X"04",X"80",X"18",
		X"EB",X"DD",X"7E",X"05",X"C1",X"FD",X"21",X"0C",X"4C",X"FD",X"09",X"FD",X"73",X"00",X"FD",X"72",
		X"01",X"FD",X"77",X"02",X"3A",X"5C",X"4C",X"DD",X"77",X"03",X"3A",X"5D",X"4C",X"DD",X"77",X"04",
		X"DD",X"7E",X"00",X"21",X"85",X"0E",X"CB",X"27",X"CD",X"BA",X"15",X"D5",X"5E",X"23",X"56",X"EB",
		X"D1",X"DD",X"7E",X"06",X"E9",X"91",X"0E",X"91",X"0E",X"92",X"0E",X"9D",X"0E",X"A0",X"0E",X"A7",
		X"0E",X"C9",X"13",X"FD",X"73",X"03",X"FD",X"72",X"04",X"FD",X"77",X"05",X"C9",X"1B",X"18",X"F3",
		X"21",X"20",X"00",X"19",X"EB",X"18",X"EC",X"EB",X"11",X"20",X"00",X"37",X"3F",X"ED",X"52",X"EB",
		X"18",X"E1",X"3A",X"5C",X"4C",X"E6",X"07",X"32",X"0A",X"4C",X"3A",X"5D",X"4C",X"E6",X"07",X"32",
		X"0B",X"4C",X"3A",X"5C",X"4C",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"57",X"3A",X"5D",X"4C",X"CB",
		X"3F",X"CB",X"3F",X"CB",X"3F",X"5F",X"CD",X"E9",X"14",X"C9",X"DD",X"7E",X"01",X"DD",X"86",X"02",
		X"47",X"E6",X"0F",X"DD",X"77",X"02",X"CB",X"38",X"CB",X"38",X"CB",X"38",X"CB",X"38",X"C9",X"3A",
		X"03",X"4D",X"21",X"FD",X"0E",X"CB",X"27",X"CB",X"27",X"CD",X"BA",X"15",X"E9",X"CD",X"CA",X"29",
		X"C9",X"CD",X"23",X"2A",X"C9",X"CD",X"7C",X"2A",X"C9",X"CD",X"D5",X"2A",X"C9",X"CD",X"2E",X"2B",
		X"C9",X"CD",X"87",X"2B",X"C9",X"CD",X"E0",X"2B",X"C9",X"CD",X"36",X"2C",X"C9",X"CD",X"8C",X"2C",
		X"C9",X"CD",X"E5",X"2C",X"C9",X"CD",X"3E",X"2D",X"C9",X"CD",X"8A",X"2D",X"C9",X"CD",X"D6",X"2D",
		X"C9",X"CD",X"D7",X"2D",X"C9",X"CD",X"D8",X"2D",X"C9",X"CD",X"D9",X"2D",X"C9",X"D5",X"37",X"3F",
		X"21",X"0E",X"01",X"16",X"00",X"ED",X"52",X"7D",X"37",X"3F",X"21",X"10",X"01",X"D1",X"5A",X"16",
		X"00",X"ED",X"52",X"55",X"5F",X"C9",X"7D",X"EE",X"03",X"6F",X"C9",X"21",X"96",X"4C",X"CB",X"46",
		X"C8",X"CB",X"6E",X"28",X"43",X"21",X"A8",X"4C",X"7B",X"86",X"27",X"77",X"23",X"7A",X"8E",X"27",
		X"77",X"23",X"3E",X"00",X"8E",X"27",X"77",X"38",X"02",X"18",X"32",X"21",X"96",X"4C",X"CB",X"6E",
		X"28",X"13",X"21",X"F6",X"43",X"11",X"F7",X"43",X"01",X"05",X"00",X"36",X"40",X"ED",X"B0",X"AF",
		X"32",X"F6",X"43",X"18",X"18",X"21",X"E4",X"43",X"11",X"E5",X"43",X"01",X"05",X"00",X"36",X"40",
		X"ED",X"B0",X"AF",X"32",X"E4",X"43",X"18",X"05",X"21",X"AB",X"4C",X"18",X"BB",X"21",X"96",X"4C",
		X"CB",X"6E",X"28",X"5C",X"21",X"AA",X"4C",X"11",X"FB",X"43",X"3A",X"B1",X"4C",X"F5",X"CD",X"1B",
		X"10",X"23",X"23",X"23",X"EB",X"2A",X"A3",X"4C",X"F1",X"FE",X"04",X"D0",X"CB",X"27",X"CB",X"27",
		X"3C",X"3C",X"CD",X"BA",X"15",X"CD",X"B0",X"11",X"D0",X"3A",X"B0",X"4C",X"3C",X"32",X"B0",X"4C",
		X"21",X"20",X"4D",X"CB",X"C6",X"21",X"96",X"4C",X"CB",X"6E",X"28",X"12",X"3A",X"B1",X"4C",X"3C",
		X"32",X"B1",X"4C",X"3A",X"A6",X"4C",X"3C",X"32",X"A6",X"4C",X"CD",X"13",X"00",X"C9",X"3A",X"B2",
		X"4C",X"3C",X"32",X"B2",X"4C",X"3A",X"A7",X"4C",X"3C",X"32",X"A7",X"4C",X"CD",X"24",X"00",X"C9",
		X"21",X"AD",X"4C",X"11",X"E9",X"43",X"3A",X"B2",X"4C",X"18",X"A2",X"3E",X"03",X"F5",X"7E",X"E6",
		X"F0",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"47",X"3A",X"96",X"4C",X"CB",X"77",X"28",
		X"22",X"78",X"12",X"1B",X"7E",X"E6",X"0F",X"47",X"3A",X"96",X"4C",X"CB",X"77",X"32",X"96",X"4C",
		X"28",X"20",X"78",X"12",X"2B",X"1B",X"F1",X"3D",X"20",X"D3",X"3A",X"96",X"4C",X"CB",X"B7",X"32",
		X"96",X"4C",X"C9",X"78",X"FE",X"00",X"28",X"DB",X"3A",X"96",X"4C",X"CB",X"F7",X"32",X"96",X"4C",
		X"18",X"CF",X"78",X"FE",X"00",X"28",X"DD",X"3A",X"96",X"4C",X"CB",X"F7",X"32",X"96",X"4C",X"18",
		X"D1",X"21",X"97",X"4C",X"CB",X"5E",X"28",X"3D",X"CB",X"9E",X"21",X"40",X"40",X"CD",X"A7",X"10",
		X"FE",X"DC",X"20",X"1C",X"21",X"40",X"44",X"CD",X"A7",X"10",X"FE",X"DD",X"20",X"12",X"47",X"E6",
		X"F0",X"32",X"51",X"4F",X"78",X"32",X"50",X"4F",X"3A",X"51",X"4F",X"B8",X"20",X"02",X"18",X"15",
		X"3E",X"40",X"CD",X"07",X"15",X"F3",X"C9",X"AF",X"11",X"80",X"03",X"86",X"23",X"1B",X"47",X"7A",
		X"B3",X"78",X"20",X"F7",X"C9",X"00",X"3E",X"40",X"CD",X"07",X"15",X"3E",X"09",X"CD",X"17",X"15",
		X"11",X"29",X"45",X"21",X"F4",X"10",X"3E",X"15",X"06",X"0B",X"CD",X"F5",X"15",X"11",X"45",X"41",
		X"21",X"3D",X"19",X"3E",X"01",X"06",X"0C",X"CD",X"DF",X"15",X"21",X"68",X"1B",X"11",X"CA",X"42",
		X"01",X"FF",X"09",X"ED",X"A0",X"13",X"10",X"FB",X"AF",X"12",X"CD",X"0C",X"16",X"3E",X"01",X"12",
		X"CD",X"F5",X"10",X"C9",X"03",X"21",X"B3",X"4C",X"11",X"6A",X"42",X"CD",X"35",X"11",X"11",X"6C",
		X"42",X"CD",X"35",X"11",X"11",X"6E",X"42",X"CD",X"35",X"11",X"11",X"70",X"42",X"CD",X"35",X"11",
		X"11",X"72",X"42",X"CD",X"35",X"11",X"11",X"74",X"42",X"CD",X"35",X"11",X"11",X"76",X"42",X"CD",
		X"35",X"11",X"11",X"78",X"42",X"CD",X"35",X"11",X"11",X"7A",X"42",X"CD",X"35",X"11",X"11",X"7C",
		X"42",X"CD",X"35",X"11",X"C9",X"06",X"03",X"0E",X"0F",X"3E",X"21",X"ED",X"A0",X"CD",X"D3",X"15",
		X"10",X"F7",X"23",X"23",X"3E",X"40",X"CD",X"D3",X"15",X"CD",X"52",X"11",X"3E",X"04",X"CD",X"BA",
		X"15",X"C9",X"3E",X"03",X"F5",X"7E",X"E6",X"F0",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",
		X"47",X"3A",X"96",X"4C",X"CB",X"77",X"28",X"2A",X"78",X"12",X"3E",X"20",X"CD",X"D3",X"15",X"7E",
		X"E6",X"0F",X"47",X"3A",X"96",X"4C",X"CB",X"77",X"32",X"96",X"4C",X"28",X"24",X"78",X"12",X"2B",
		X"3E",X"20",X"CD",X"D3",X"15",X"F1",X"3D",X"20",X"CB",X"3A",X"96",X"4C",X"CB",X"B7",X"32",X"96",
		X"4C",X"C9",X"78",X"FE",X"00",X"28",X"D3",X"3A",X"96",X"4C",X"CB",X"F7",X"32",X"96",X"4C",X"18",
		X"C7",X"78",X"FE",X"00",X"28",X"D9",X"3A",X"96",X"4C",X"CB",X"F7",X"32",X"96",X"4C",X"18",X"CD",
		X"06",X"03",X"1A",X"BE",X"38",X"08",X"20",X"0E",X"2B",X"1B",X"10",X"F6",X"18",X"06",X"CD",X"CB",
		X"11",X"37",X"3F",X"C9",X"37",X"C9",X"CD",X"CB",X"11",X"37",X"C9",X"78",X"FE",X"00",X"C8",X"2B",
		X"1B",X"3D",X"20",X"FB",X"C9",X"DE",X"47",X"4F",X"52",X"4B",X"41",X"4E",X"53",X"2C",X"43",X"4F",
		X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"20",X"31",X"39",X"38",X"33",X"54",X"45",X"43",X"48",
		X"53",X"54",X"41",X"52",X"20",X"49",X"4E",X"43",X"21",X"96",X"4C",X"CB",X"EE",X"21",X"A8",X"4C",
		X"11",X"F5",X"4C",X"01",X"03",X"00",X"ED",X"B0",X"CD",X"22",X"12",X"21",X"96",X"4C",X"CB",X"66",
		X"C0",X"CB",X"AE",X"21",X"AB",X"4C",X"11",X"F5",X"4C",X"01",X"03",X"00",X"ED",X"B0",X"CD",X"22",
		X"12",X"C9",X"01",X"00",X"0A",X"21",X"F1",X"4C",X"11",X"F7",X"4C",X"2B",X"2B",X"2B",X"C5",X"CD",
		X"B0",X"11",X"C1",X"30",X"0A",X"3E",X"06",X"81",X"4F",X"10",X"ED",X"2B",X"2B",X"18",X"08",X"79",
		X"FE",X"00",X"C8",X"23",X"23",X"23",X"23",X"C5",X"E5",X"06",X"00",X"21",X"EE",X"4C",X"11",X"F4",
		X"4C",X"ED",X"B8",X"3E",X"40",X"CD",X"07",X"15",X"21",X"96",X"4C",X"CB",X"6E",X"20",X"1B",X"11",
		X"62",X"41",X"21",X"05",X"19",X"3E",X"01",X"06",X"0A",X"CD",X"DF",X"15",X"21",X"96",X"4C",X"CB",
		X"7E",X"28",X"19",X"3E",X"01",X"32",X"03",X"50",X"18",X"12",X"11",X"62",X"41",X"21",X"F8",X"18",
		X"3E",X"01",X"06",X"0A",X"CD",X"DF",X"15",X"3E",X"00",X"32",X"03",X"50",X"11",X"40",X"44",X"21",
		X"E5",X"14",X"3E",X"0B",X"06",X"1C",X"CD",X"F5",X"15",X"11",X"4C",X"44",X"21",X"E6",X"14",X"3E",
		X"03",X"06",X"1C",X"CD",X"F5",X"15",X"11",X"51",X"44",X"21",X"E7",X"14",X"3E",X"10",X"06",X"1C",
		X"CD",X"F5",X"15",X"11",X"50",X"44",X"21",X"E8",X"14",X"3E",X"02",X"06",X"1C",X"CD",X"F5",X"15",
		X"D1",X"D5",X"3E",X"40",X"D5",X"E1",X"13",X"01",X"03",X"00",X"77",X"ED",X"B0",X"36",X"00",X"01",
		X"02",X"00",X"ED",X"B0",X"D1",X"C1",X"D5",X"78",X"21",X"A9",X"1B",X"CB",X"27",X"CD",X"BA",X"15",
		X"4E",X"23",X"46",X"C5",X"21",X"80",X"04",X"09",X"0E",X"01",X"06",X"0F",X"71",X"3E",X"20",X"CD",
		X"C9",X"15",X"10",X"F8",X"11",X"C3",X"40",X"21",X"49",X"19",X"3E",X"01",X"06",X"14",X"CD",X"DF",
		X"15",X"11",X"A5",X"41",X"21",X"5D",X"19",X"3E",X"01",X"06",X"07",X"CD",X"DF",X"15",X"11",X"A7",
		X"40",X"21",X"64",X"19",X"3E",X"01",X"06",X"16",X"CD",X"DF",X"15",X"11",X"88",X"40",X"21",X"7A",
		X"19",X"3E",X"01",X"06",X"17",X"CD",X"DF",X"15",X"11",X"69",X"42",X"21",X"91",X"19",X"3E",X"01",
		X"06",X"08",X"CD",X"DF",X"15",X"11",X"4C",X"40",X"21",X"99",X"19",X"3E",X"03",X"06",X"01",X"CD",
		X"DF",X"15",X"11",X"8D",X"40",X"21",X"8B",X"1B",X"3E",X"01",X"06",X"1A",X"CD",X"DF",X"15",X"3E",
		X"01",X"11",X"AD",X"47",X"12",X"AF",X"32",X"F9",X"4C",X"32",X"FA",X"4C",X"21",X"AD",X"47",X"22",
		X"FB",X"4C",X"11",X"71",X"41",X"21",X"3D",X"19",X"3E",X"01",X"06",X"0C",X"CD",X"DF",X"15",X"21",
		X"68",X"1B",X"11",X"F4",X"42",X"01",X"09",X"00",X"ED",X"B0",X"AF",X"12",X"CD",X"0C",X"16",X"3E",
		X"01",X"12",X"21",X"B3",X"4C",X"11",X"94",X"42",X"CD",X"35",X"11",X"11",X"95",X"42",X"CD",X"35",
		X"11",X"11",X"96",X"42",X"CD",X"35",X"11",X"11",X"97",X"42",X"CD",X"35",X"11",X"11",X"98",X"42",
		X"CD",X"35",X"11",X"11",X"99",X"42",X"CD",X"35",X"11",X"11",X"9A",X"42",X"CD",X"35",X"11",X"11",
		X"9B",X"42",X"CD",X"35",X"11",X"11",X"9C",X"42",X"CD",X"35",X"11",X"11",X"9D",X"42",X"CD",X"35",
		X"11",X"3A",X"F8",X"4C",X"CB",X"4F",X"CA",X"4D",X"14",X"CB",X"57",X"CA",X"85",X"14",X"3A",X"F8",
		X"4C",X"CB",X"67",X"C2",X"C6",X"14",X"3A",X"F9",X"4C",X"FE",X"1B",X"28",X"1F",X"21",X"71",X"1B",
		X"CD",X"BA",X"15",X"7E",X"E1",X"D1",X"12",X"13",X"77",X"3E",X"20",X"CD",X"C9",X"15",X"D5",X"E5",
		X"3A",X"FA",X"4C",X"3C",X"32",X"FA",X"4C",X"FE",X"03",X"C2",X"D9",X"14",X"21",X"BD",X"1B",X"3A",
		X"FA",X"4C",X"CD",X"BA",X"15",X"7E",X"E1",X"D1",X"E5",X"CD",X"BF",X"15",X"21",X"F5",X"4C",X"01",
		X"03",X"00",X"ED",X"B0",X"3A",X"FA",X"4C",X"FE",X"00",X"28",X"25",X"21",X"C1",X"1B",X"CD",X"BA",
		X"15",X"7E",X"D1",X"CD",X"D3",X"15",X"21",X"F7",X"4C",X"CD",X"52",X"11",X"21",X"B8",X"4C",X"11",
		X"F2",X"43",X"CD",X"1B",X"10",X"21",X"97",X"4C",X"CB",X"86",X"3E",X"01",X"CD",X"59",X"15",X"C9",
		X"D1",X"3E",X"80",X"CD",X"D3",X"15",X"3E",X"20",X"CD",X"D3",X"15",X"18",X"D9",X"3A",X"F9",X"4C",
		X"FE",X"00",X"CA",X"CE",X"13",X"3D",X"32",X"F9",X"4C",X"FE",X"1A",X"28",X"14",X"3E",X"05",X"2A",
		X"FB",X"4C",X"77",X"3E",X"20",X"CD",X"BA",X"15",X"22",X"FB",X"4C",X"3E",X"01",X"77",X"C3",X"CE",
		X"13",X"3D",X"32",X"F9",X"4C",X"3E",X"05",X"2A",X"FB",X"4C",X"2B",X"77",X"23",X"77",X"23",X"77",
		X"2B",X"3E",X"40",X"18",X"E0",X"3A",X"F9",X"4C",X"FE",X"1B",X"CA",X"CE",X"13",X"3C",X"32",X"F9",
		X"4C",X"FE",X"1A",X"28",X"14",X"3E",X"05",X"2A",X"FB",X"4C",X"77",X"3E",X"20",X"CD",X"C9",X"15",
		X"22",X"FB",X"4C",X"3E",X"01",X"77",X"C3",X"CE",X"13",X"3C",X"32",X"F9",X"4C",X"3E",X"05",X"2A",
		X"FB",X"4C",X"77",X"3E",X"40",X"CD",X"C9",X"15",X"22",X"FB",X"4C",X"3E",X"01",X"2B",X"77",X"23",
		X"77",X"23",X"77",X"C3",X"CE",X"13",X"3E",X"08",X"CD",X"A5",X"15",X"32",X"C0",X"50",X"06",X"14",
		X"CD",X"71",X"15",X"DA",X"FC",X"13",X"C3",X"C1",X"13",X"3A",X"F8",X"4C",X"CB",X"67",X"32",X"C0",
		X"50",X"28",X"F6",X"18",X"E6",X"09",X"05",X"10",X"01",X"D5",X"AF",X"CB",X"23",X"17",X"CB",X"23",
		X"17",X"CB",X"23",X"17",X"CB",X"23",X"17",X"CB",X"23",X"17",X"57",X"EB",X"01",X"40",X"40",X"09",
		X"06",X"00",X"D1",X"4A",X"09",X"EB",X"C9",X"21",X"40",X"40",X"11",X"41",X"40",X"01",X"7F",X"03",
		X"77",X"ED",X"B0",X"32",X"C0",X"50",X"C9",X"21",X"40",X"44",X"11",X"41",X"44",X"01",X"7F",X"03",
		X"77",X"ED",X"B0",X"32",X"C0",X"50",X"C9",X"3A",X"9B",X"4C",X"FE",X"00",X"C8",X"3A",X"9D",X"4C",
		X"E6",X"F0",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"FE",X"00",X"28",X"0C",X"32",X"0D",
		X"40",X"3A",X"9D",X"4C",X"E6",X"0F",X"32",X"0C",X"40",X"C9",X"3E",X"40",X"18",X"F0",X"3E",X"09",
		X"CD",X"17",X"15",X"3E",X"40",X"CD",X"07",X"15",X"C9",X"47",X"AF",X"32",X"9E",X"4C",X"32",X"A0",
		X"4C",X"3A",X"A0",X"4C",X"B8",X"C8",X"21",X"95",X"4C",X"CB",X"6E",X"C0",X"32",X"C0",X"50",X"18",
		X"F0",X"3A",X"97",X"4C",X"CB",X"47",X"28",X"0D",X"3A",X"A1",X"4C",X"47",X"3A",X"A0",X"4C",X"B8",
		X"30",X"19",X"37",X"3F",X"C9",X"78",X"32",X"A1",X"4C",X"3A",X"97",X"4C",X"CB",X"C7",X"32",X"97",
		X"4C",X"AF",X"32",X"A0",X"4C",X"32",X"9E",X"4C",X"37",X"3F",X"C9",X"3A",X"97",X"4C",X"CB",X"87",
		X"32",X"97",X"4C",X"37",X"C9",X"47",X"AF",X"32",X"9F",X"4C",X"3A",X"9F",X"4C",X"B8",X"C8",X"21",
		X"95",X"4C",X"CB",X"6E",X"C0",X"32",X"C0",X"50",X"18",X"F0",X"85",X"6F",X"D0",X"24",X"C9",X"83",
		X"5F",X"D0",X"14",X"C9",X"81",X"4F",X"D0",X"04",X"C9",X"D5",X"16",X"00",X"5F",X"37",X"3F",X"ED",
		X"52",X"D1",X"C9",X"E5",X"EB",X"16",X"00",X"5F",X"37",X"3F",X"ED",X"52",X"EB",X"E1",X"C9",X"32",
		X"60",X"4C",X"D5",X"3A",X"60",X"4C",X"4F",X"ED",X"A0",X"79",X"FE",X"00",X"20",X"F9",X"D1",X"CD",
		X"0C",X"16",X"10",X"EE",X"C9",X"32",X"60",X"4C",X"D5",X"3A",X"60",X"4C",X"4F",X"ED",X"A0",X"2B",
		X"79",X"FE",X"00",X"20",X"F8",X"D1",X"CD",X"0C",X"16",X"10",X"ED",X"C9",X"E5",X"21",X"20",X"00",
		X"19",X"EB",X"E1",X"C9",X"21",X"61",X"4C",X"06",X"2F",X"36",X"00",X"23",X"10",X"FB",X"C9",X"21",
		X"95",X"4C",X"CB",X"FE",X"CB",X"7E",X"C8",X"18",X"FB",X"3A",X"00",X"50",X"E6",X"0F",X"47",X"3A",
		X"40",X"50",X"E6",X"F0",X"B0",X"32",X"F8",X"4C",X"C9",X"3A",X"40",X"50",X"47",X"E6",X"0F",X"CB",
		X"78",X"28",X"02",X"CB",X"E7",X"32",X"F8",X"4C",X"C9",X"DD",X"21",X"05",X"4D",X"DD",X"CB",X"00",
		X"46",X"C4",X"7A",X"17",X"DD",X"CB",X"00",X"56",X"28",X"10",X"CD",X"82",X"17",X"FD",X"21",X"51",
		X"50",X"CD",X"51",X"17",X"DD",X"7E",X"06",X"32",X"45",X"50",X"DD",X"21",X"20",X"4D",X"DD",X"CB",
		X"00",X"46",X"C4",X"7A",X"17",X"DD",X"CB",X"00",X"56",X"28",X"10",X"CD",X"82",X"17",X"FD",X"21",
		X"51",X"50",X"CD",X"51",X"17",X"DD",X"7E",X"06",X"32",X"45",X"50",X"DD",X"21",X"3B",X"4D",X"DD",
		X"CB",X"00",X"46",X"C4",X"7A",X"17",X"DD",X"CB",X"00",X"56",X"28",X"10",X"CD",X"82",X"17",X"FD",
		X"21",X"51",X"50",X"CD",X"51",X"17",X"DD",X"7E",X"06",X"32",X"45",X"50",X"DD",X"21",X"56",X"4D",
		X"DD",X"CB",X"00",X"46",X"C4",X"7A",X"17",X"DD",X"CB",X"00",X"56",X"28",X"10",X"CD",X"82",X"17",
		X"FD",X"21",X"56",X"50",X"CD",X"51",X"17",X"DD",X"7E",X"06",X"32",X"4A",X"50",X"DD",X"21",X"71",
		X"4D",X"DD",X"CB",X"00",X"46",X"C4",X"7A",X"17",X"DD",X"CB",X"00",X"56",X"28",X"10",X"CD",X"82",
		X"17",X"FD",X"21",X"56",X"50",X"CD",X"51",X"17",X"DD",X"7E",X"06",X"32",X"4A",X"50",X"DD",X"21",
		X"8C",X"4D",X"DD",X"CB",X"00",X"46",X"C4",X"7A",X"17",X"DD",X"CB",X"00",X"56",X"28",X"10",X"CD",
		X"82",X"17",X"FD",X"21",X"56",X"50",X"CD",X"51",X"17",X"DD",X"7E",X"06",X"32",X"4A",X"50",X"DD",
		X"21",X"A7",X"4D",X"DD",X"CB",X"00",X"46",X"C4",X"7A",X"17",X"DD",X"CB",X"00",X"56",X"28",X"10",
		X"CD",X"82",X"17",X"FD",X"21",X"5B",X"50",X"CD",X"51",X"17",X"DD",X"7E",X"06",X"32",X"4F",X"50",
		X"DD",X"21",X"C2",X"4D",X"DD",X"CB",X"00",X"46",X"C4",X"7A",X"17",X"DD",X"CB",X"00",X"56",X"C8",
		X"CD",X"82",X"17",X"FD",X"21",X"5B",X"50",X"CD",X"51",X"17",X"DD",X"7E",X"06",X"32",X"4F",X"50",
		X"C9",X"DD",X"7E",X"03",X"FD",X"77",X"00",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"FD",
		X"77",X"01",X"DD",X"7E",X"04",X"FD",X"77",X"02",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",
		X"FD",X"77",X"03",X"DD",X"7E",X"05",X"FD",X"77",X"04",X"C9",X"CD",X"56",X"18",X"DD",X"CB",X"00",
		X"D6",X"C9",X"DD",X"CB",X"00",X"4E",X"C2",X"56",X"18",X"DD",X"6E",X"01",X"DD",X"66",X"02",X"7E",
		X"CB",X"27",X"11",X"A0",X"17",X"CD",X"BF",X"15",X"23",X"E5",X"1A",X"6F",X"13",X"1A",X"67",X"E9",
		X"BA",X"17",X"BE",X"17",X"CC",X"17",X"D5",X"17",X"EB",X"17",X"F8",X"17",X"12",X"18",X"2B",X"18",
		X"4D",X"18",X"55",X"18",X"74",X"18",X"80",X"18",X"8C",X"18",X"E1",X"C3",X"8F",X"17",X"E1",X"7E",
		X"DD",X"77",X"03",X"23",X"7E",X"23",X"DD",X"77",X"04",X"C3",X"8F",X"17",X"E1",X"7E",X"DD",X"77",
		X"05",X"23",X"C3",X"8F",X"17",X"E1",X"7E",X"DD",X"46",X"03",X"80",X"DD",X"77",X"03",X"23",X"7E",
		X"23",X"DD",X"46",X"04",X"88",X"DD",X"77",X"04",X"C3",X"8F",X"17",X"E1",X"7E",X"DD",X"46",X"05",
		X"80",X"DD",X"77",X"05",X"23",X"C3",X"8F",X"17",X"E1",X"DD",X"7E",X"07",X"BE",X"30",X"0B",X"DD",
		X"34",X"07",X"2B",X"DD",X"75",X"01",X"DD",X"74",X"02",X"C9",X"DD",X"36",X"07",X"00",X"23",X"C3",
		X"8F",X"17",X"DD",X"6E",X"08",X"DD",X"66",X"09",X"D1",X"D5",X"2B",X"72",X"2B",X"73",X"2B",X"36",
		X"00",X"DD",X"75",X"08",X"DD",X"74",X"09",X"E1",X"C3",X"8F",X"17",X"D1",X"1A",X"DD",X"6E",X"08",
		X"DD",X"66",X"09",X"BE",X"28",X"09",X"34",X"23",X"5E",X"23",X"56",X"EB",X"C3",X"8F",X"17",X"23",
		X"23",X"23",X"DD",X"75",X"08",X"DD",X"74",X"09",X"13",X"EB",X"C3",X"8F",X"17",X"E1",X"5E",X"23",
		X"56",X"EB",X"C3",X"8F",X"17",X"E1",X"DD",X"E5",X"DD",X"E5",X"E1",X"D1",X"13",X"36",X"00",X"01",
		X"18",X"00",X"ED",X"B0",X"1A",X"DD",X"77",X"01",X"13",X"1A",X"DD",X"77",X"02",X"DD",X"75",X"08",
		X"DD",X"74",X"09",X"C9",X"E1",X"DD",X"75",X"01",X"DD",X"74",X"02",X"DD",X"36",X"00",X"00",X"C9",
		X"E1",X"5E",X"23",X"56",X"EB",X"36",X"06",X"13",X"EB",X"C3",X"8F",X"17",X"E1",X"7E",X"DD",X"77",
		X"06",X"23",X"C3",X"8F",X"17",X"32",X"40",X"52",X"45",X"59",X"41",X"4C",X"50",X"40",X"45",X"52",
		X"4F",X"43",X"53",X"50",X"4F",X"54",X"40",X"31",X"40",X"52",X"45",X"59",X"41",X"4C",X"50",X"54",
		X"49",X"44",X"45",X"52",X"43",X"59",X"41",X"4C",X"50",X"45",X"45",X"52",X"46",X"40",X"4E",X"49",
		X"4F",X"43",X"40",X"54",X"52",X"45",X"53",X"4E",X"49",X"52",X"45",X"59",X"41",X"4C",X"50",X"40",
		X"45",X"4E",X"4F",X"40",X"54",X"43",X"45",X"4C",X"45",X"53",X"52",X"4F",X"53",X"52",X"45",X"59",
		X"41",X"4C",X"50",X"40",X"4F",X"57",X"54",X"40",X"52",X"4F",X"40",X"45",X"4E",X"4F",X"40",X"54",
		X"43",X"45",X"4C",X"45",X"53",X"50",X"55",X"40",X"45",X"4E",X"4F",X"40",X"52",X"45",X"59",X"41",
		X"4C",X"50",X"50",X"55",X"40",X"4F",X"57",X"54",X"40",X"52",X"45",X"59",X"41",X"4C",X"50",X"4E",
		X"49",X"41",X"47",X"41",X"40",X"52",X"45",X"59",X"41",X"4C",X"50",X"40",X"45",X"4D",X"41",X"53",
		X"52",X"45",X"56",X"4F",X"40",X"45",X"4D",X"41",X"47",X"52",X"45",X"56",X"4F",X"40",X"45",X"4D",
		X"41",X"47",X"40",X"45",X"4E",X"4F",X"40",X"52",X"45",X"59",X"41",X"4C",X"50",X"45",X"4D",X"41",
		X"46",X"40",X"46",X"4F",X"40",X"4C",X"4C",X"41",X"48",X"45",X"48",X"54",X"40",X"4E",X"49",X"40",
		X"53",X"49",X"40",X"45",X"52",X"4F",X"43",X"53",X"40",X"52",X"55",X"4F",X"59",X"4E",X"45",X"54",
		X"40",X"50",X"4F",X"54",X"54",X"43",X"45",X"4C",X"45",X"53",X"40",X"4F",X"54",X"40",X"4B",X"43",
		X"49",X"54",X"53",X"59",X"4F",X"4A",X"40",X"45",X"53",X"55",X"4E",X"4F",X"54",X"54",X"55",X"42",
		X"40",X"44",X"45",X"45",X"50",X"53",X"40",X"44",X"4E",X"41",X"40",X"52",X"45",X"54",X"54",X"45",
		X"4C",X"54",X"4E",X"49",X"52",X"50",X"40",X"4F",X"54",X"45",X"4E",X"44",X"4D",X"41",X"4C",X"53",
		X"45",X"43",X"4E",X"41",X"56",X"44",X"41",X"40",X"45",X"52",X"4F",X"43",X"53",X"40",X"53",X"4E",
		X"41",X"4B",X"52",X"4F",X"47",X"45",X"52",X"4F",X"43",X"53",X"40",X"40",X"53",X"4E",X"4F",X"49",
		X"54",X"43",X"45",X"53",X"52",X"45",X"54",X"4E",X"49",X"52",X"45",X"42",X"4D",X"55",X"4E",X"40",
		X"45",X"53",X"41",X"42",X"40",X"58",X"40",X"53",X"54",X"4E",X"49",X"4F",X"50",X"40",X"30",X"31",
		X"40",X"53",X"45",X"52",X"4F",X"43",X"40",X"52",X"41",X"45",X"4C",X"43",X"55",X"4E",X"40",X"4E",
		X"41",X"4B",X"52",X"4F",X"47",X"40",X"64",X"64",X"64",X"64",X"40",X"40",X"40",X"45",X"52",X"4F",
		X"43",X"53",X"40",X"59",X"41",X"4C",X"50",X"40",X"31",X"40",X"53",X"4E",X"49",X"4F",X"43",X"40",
		X"32",X"53",X"59",X"41",X"4C",X"50",X"40",X"32",X"40",X"40",X"4E",X"49",X"4F",X"43",X"40",X"31",
		X"40",X"59",X"41",X"4C",X"50",X"40",X"31",X"40",X"40",X"4E",X"49",X"4F",X"43",X"40",X"31",X"53",
		X"54",X"4E",X"49",X"4F",X"50",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"59",X"52",X"45",
		X"56",X"45",X"40",X"53",X"55",X"4E",X"4F",X"42",X"30",X"30",X"30",X"30",X"35",X"31",X"30",X"30",
		X"30",X"35",X"32",X"31",X"30",X"30",X"30",X"30",X"30",X"31",X"40",X"30",X"30",X"30",X"35",X"37",
		X"53",X"43",X"49",X"54",X"53",X"4F",X"4E",X"47",X"41",X"49",X"44",X"4E",X"4F",X"49",X"54",X"49",
		X"44",X"4E",X"4F",X"43",X"40",X"40",X"4E",X"4F",X"49",X"54",X"41",X"43",X"4F",X"4C",X"40",X"40",
		X"4D",X"4F",X"52",X"44",X"4F",X"4F",X"47",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"44",X"37",
		X"40",X"40",X"40",X"40",X"40",X"40",X"31",X"44",X"4F",X"4F",X"47",X"40",X"40",X"40",X"40",X"40",
		X"40",X"40",X"46",X"37",X"40",X"40",X"40",X"40",X"40",X"40",X"32",X"44",X"4F",X"4F",X"47",X"40",
		X"40",X"40",X"40",X"40",X"40",X"40",X"48",X"37",X"40",X"40",X"40",X"40",X"40",X"40",X"33",X"44",
		X"4F",X"4F",X"47",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"4A",X"37",X"40",X"40",X"40",X"40",
		X"40",X"40",X"34",X"44",X"4F",X"4F",X"47",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"48",X"34",
		X"40",X"40",X"40",X"40",X"40",X"40",X"31",X"44",X"4F",X"4F",X"47",X"40",X"40",X"40",X"40",X"40",
		X"40",X"40",X"4C",X"34",X"40",X"40",X"40",X"40",X"40",X"40",X"32",X"44",X"4F",X"4F",X"47",X"40",
		X"40",X"40",X"40",X"40",X"40",X"40",X"4A",X"34",X"40",X"40",X"40",X"40",X"40",X"40",X"33",X"44",
		X"4F",X"4F",X"47",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"4D",X"34",X"40",X"40",X"40",X"40",
		X"40",X"40",X"34",X"44",X"4F",X"4F",X"47",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"4B",X"34",
		X"40",X"40",X"40",X"40",X"40",X"40",X"35",X"44",X"4F",X"4F",X"47",X"40",X"40",X"40",X"40",X"40",
		X"40",X"40",X"4E",X"34",X"40",X"40",X"40",X"40",X"40",X"40",X"36",X"44",X"41",X"42",X"40",X"4E",
		X"4F",X"49",X"54",X"49",X"44",X"4E",X"4F",X"43",X"40",X"40",X"4E",X"4F",X"49",X"54",X"41",X"43",
		X"4F",X"4C",X"40",X"40",X"4D",X"41",X"52",X"00",X"01",X"02",X"03",X"04",X"05",X"06",X"07",X"08",
		X"09",X"41",X"42",X"43",X"44",X"45",X"46",X"47",X"48",X"49",X"4A",X"4B",X"4C",X"4D",X"4E",X"4F",
		X"50",X"51",X"52",X"53",X"54",X"55",X"56",X"57",X"58",X"59",X"5A",X"5A",X"59",X"58",X"57",X"56",
		X"55",X"54",X"53",X"52",X"51",X"50",X"4F",X"4E",X"4D",X"4C",X"4B",X"4A",X"49",X"48",X"47",X"46",
		X"45",X"44",X"43",X"42",X"41",X"00",X"01",X"04",X"02",X"94",X"42",X"95",X"42",X"96",X"42",X"97",
		X"42",X"98",X"42",X"99",X"42",X"9A",X"42",X"9B",X"42",X"9C",X"42",X"9D",X"42",X"03",X"02",X"01",
		X"00",X"00",X"80",X"60",X"40",X"21",X"DD",X"4D",X"CB",X"46",X"C2",X"5B",X"1C",X"CB",X"C6",X"11",
		X"CE",X"44",X"21",X"9B",X"4E",X"3E",X"05",X"06",X"14",X"CD",X"F5",X"15",X"06",X"14",X"21",X"37",
		X"4E",X"11",X"CE",X"40",X"C5",X"01",X"05",X"00",X"ED",X"B0",X"3E",X"1B",X"CD",X"BF",X"15",X"C1",
		X"10",X"F2",X"2A",X"9D",X"4E",X"23",X"7E",X"2B",X"FE",X"00",X"20",X"1F",X"2A",X"2F",X"4E",X"06",
		X"10",X"3A",X"34",X"4E",X"5E",X"23",X"56",X"12",X"CD",X"10",X"1C",X"23",X"10",X"F3",X"18",X"41",
		X"E5",X"21",X"00",X"04",X"19",X"3A",X"E2",X"4E",X"77",X"E1",X"C9",X"06",X"10",X"5E",X"23",X"56",
		X"7A",X"FE",X"00",X"28",X"11",X"3A",X"34",X"4E",X"12",X"CD",X"10",X"1C",X"3A",X"2A",X"4E",X"3C",
		X"32",X"2A",X"4E",X"23",X"10",X"E7",X"3A",X"2A",X"4E",X"47",X"3E",X"10",X"90",X"32",X"29",X"4E",
		X"AF",X"32",X"2A",X"4E",X"2A",X"9D",X"4E",X"E5",X"D1",X"13",X"01",X"1F",X"00",X"36",X"00",X"ED",
		X"B0",X"3E",X"3C",X"CD",X"A5",X"15",X"21",X"71",X"4D",X"CB",X"C6",X"00",X"3E",X"04",X"32",X"15",
		X"4E",X"3A",X"31",X"4E",X"32",X"16",X"4E",X"21",X"74",X"27",X"11",X"17",X"4E",X"01",X"04",X"00",
		X"ED",X"B0",X"FD",X"21",X"89",X"4C",X"FD",X"7E",X"07",X"E6",X"E0",X"47",X"3A",X"F8",X"4C",X"E6",
		X"1F",X"B0",X"FD",X"77",X"07",X"2A",X"11",X"4E",X"22",X"0F",X"4E",X"21",X"F8",X"4D",X"CD",X"A7",
		X"1F",X"3A",X"E4",X"4E",X"FD",X"BE",X"05",X"28",X"12",X"3A",X"90",X"4C",X"CB",X"77",X"28",X"0B",
		X"21",X"A7",X"4D",X"CB",X"C6",X"FD",X"7E",X"05",X"32",X"E4",X"4E",X"21",X"00",X"00",X"22",X"0F",
		X"4E",X"3A",X"13",X"4E",X"32",X"15",X"4E",X"3A",X"14",X"4E",X"32",X"16",X"4E",X"21",X"78",X"27",
		X"11",X"17",X"4E",X"01",X"04",X"00",X"ED",X"B0",X"3A",X"1B",X"4E",X"FE",X"B5",X"28",X"25",X"FE",
		X"3C",X"28",X"0A",X"FE",X"78",X"28",X"0D",X"FE",X"B4",X"28",X"10",X"18",X"13",X"21",X"70",X"4C",
		X"CB",X"F6",X"18",X"0C",X"21",X"78",X"4C",X"CB",X"F6",X"18",X"05",X"21",X"80",X"4C",X"CB",X"F6",
		X"3C",X"32",X"1B",X"4E",X"00",X"DD",X"21",X"89",X"4C",X"FD",X"21",X"61",X"4C",X"CD",X"CD",X"27",
		X"CD",X"7B",X"28",X"DD",X"21",X"89",X"4C",X"21",X"FB",X"4D",X"CD",X"A7",X"1F",X"DD",X"21",X"89",
		X"4C",X"FD",X"21",X"69",X"4C",X"CD",X"CD",X"27",X"CD",X"AB",X"28",X"DD",X"21",X"89",X"4C",X"21",
		X"FE",X"4D",X"CD",X"A7",X"1F",X"DD",X"21",X"89",X"4C",X"FD",X"21",X"71",X"4C",X"CD",X"CD",X"27",
		X"CD",X"CD",X"28",X"DD",X"21",X"89",X"4C",X"21",X"01",X"4E",X"CD",X"A7",X"1F",X"DD",X"21",X"89",
		X"4C",X"FD",X"21",X"79",X"4C",X"CD",X"CD",X"27",X"21",X"04",X"4E",X"CD",X"A7",X"1F",X"3A",X"33",
		X"4E",X"3C",X"32",X"33",X"4E",X"FE",X"04",X"20",X"2C",X"AF",X"32",X"33",X"4E",X"3A",X"32",X"4E",
		X"FE",X"02",X"28",X"1E",X"3C",X"32",X"32",X"4E",X"47",X"3A",X"34",X"4E",X"80",X"4F",X"2A",X"2F",
		X"4E",X"06",X"10",X"5E",X"23",X"56",X"23",X"1A",X"FE",X"66",X"38",X"02",X"79",X"12",X"10",X"F3",
		X"18",X"03",X"AF",X"18",X"E0",X"00",X"3A",X"84",X"4C",X"FE",X"00",X"28",X"51",X"3A",X"2B",X"4E",
		X"3C",X"32",X"2B",X"4E",X"FE",X"03",X"C2",X"DE",X"1D",X"AF",X"32",X"2B",X"4E",X"3A",X"2C",X"4E",
		X"3C",X"32",X"2C",X"4E",X"FE",X"07",X"30",X"19",X"3A",X"84",X"4C",X"FE",X"01",X"28",X"0A",X"32",
		X"2E",X"4E",X"3E",X"01",X"32",X"84",X"4C",X"18",X"25",X"3A",X"2E",X"4E",X"32",X"84",X"4C",X"18",
		X"1D",X"FE",X"14",X"28",X"0D",X"3A",X"2D",X"4E",X"32",X"86",X"4C",X"3E",X"07",X"32",X"87",X"4C",
		X"18",X"0C",X"AF",X"32",X"2C",X"4E",X"32",X"84",X"4C",X"3E",X"09",X"32",X"87",X"4C",X"3A",X"26",
		X"4E",X"FE",X"04",X"20",X"22",X"AF",X"32",X"26",X"4E",X"3A",X"30",X"40",X"47",X"3A",X"2F",X"40",
		X"4F",X"3A",X"27",X"4E",X"32",X"30",X"40",X"3A",X"28",X"4E",X"32",X"2F",X"40",X"78",X"32",X"27",
		X"4E",X"79",X"32",X"28",X"4E",X"18",X"04",X"3C",X"32",X"26",X"4E",X"3A",X"29",X"4E",X"FE",X"FF",
		X"CA",X"79",X"1E",X"FE",X"10",X"C2",X"9E",X"1E",X"21",X"A7",X"4D",X"CB",X"CE",X"21",X"8C",X"4D",
		X"CB",X"C6",X"3E",X"5A",X"CD",X"A5",X"15",X"CD",X"14",X"16",X"11",X"4E",X"40",X"21",X"4E",X"1F",
		X"3E",X"05",X"06",X"1C",X"CD",X"F5",X"15",X"11",X"4E",X"44",X"21",X"A6",X"1F",X"3E",X"05",X"06",
		X"1C",X"CD",X"F5",X"15",X"11",X"2F",X"41",X"21",X"6A",X"1F",X"3E",X"01",X"06",X"0F",X"CD",X"DF",
		X"15",X"11",X"71",X"40",X"21",X"4F",X"1F",X"3E",X"01",X"06",X"1B",X"CD",X"DF",X"15",X"3E",X"B4",
		X"CD",X"A5",X"15",X"AF",X"32",X"62",X"4C",X"32",X"6A",X"4C",X"32",X"72",X"4C",X"32",X"7A",X"4C",
		X"32",X"82",X"4C",X"32",X"8A",X"4C",X"C3",X"3A",X"1F",X"AF",X"32",X"62",X"4C",X"32",X"6A",X"4C",
		X"32",X"72",X"4C",X"32",X"7A",X"4C",X"32",X"82",X"4C",X"32",X"8A",X"4C",X"21",X"71",X"4D",X"CB",
		X"CE",X"21",X"A7",X"4D",X"CB",X"CE",X"21",X"3B",X"4D",X"CB",X"CE",X"C3",X"33",X"1F",X"3A",X"90",
		X"4C",X"CB",X"6F",X"C2",X"4D",X"1F",X"CB",X"77",X"20",X"10",X"21",X"96",X"4C",X"CB",X"CE",X"3E",
		X"40",X"32",X"2F",X"40",X"32",X"30",X"40",X"C3",X"4D",X"1F",X"3A",X"68",X"4C",X"47",X"3A",X"70",
		X"4C",X"B0",X"47",X"3A",X"78",X"4C",X"B0",X"47",X"3A",X"80",X"4C",X"B0",X"47",X"3A",X"88",X"4C",
		X"B0",X"CB",X"77",X"C2",X"4D",X"1F",X"47",X"AF",X"32",X"8A",X"4C",X"21",X"71",X"4D",X"CB",X"CE",
		X"21",X"A7",X"4D",X"CB",X"CE",X"CB",X"68",X"20",X"64",X"21",X"00",X"00",X"22",X"E0",X"4E",X"3E",
		X"5A",X"CD",X"A5",X"15",X"3A",X"34",X"4E",X"47",X"3A",X"32",X"4E",X"80",X"32",X"9F",X"4E",X"01",
		X"80",X"03",X"21",X"40",X"40",X"3A",X"9F",X"4E",X"ED",X"B1",X"78",X"B1",X"28",X"21",X"2B",X"36",
		X"0A",X"C5",X"E5",X"11",X"00",X"04",X"19",X"3A",X"40",X"44",X"77",X"11",X"00",X"10",X"CD",X"5B",
		X"0F",X"21",X"8C",X"4D",X"CB",X"C6",X"3E",X"0F",X"CD",X"A5",X"15",X"E1",X"C1",X"18",X"D6",X"AF",
		X"32",X"84",X"4C",X"3A",X"84",X"4C",X"FE",X"00",X"20",X"13",X"21",X"96",X"4C",X"CB",X"DE",X"CB",
		X"CE",X"AF",X"32",X"1B",X"4E",X"3E",X"40",X"32",X"2F",X"40",X"32",X"30",X"40",X"C9",X"40",X"44",
		X"45",X"59",X"4F",X"52",X"54",X"53",X"45",X"44",X"40",X"45",X"52",X"4F",X"43",X"40",X"52",X"41",
		X"45",X"4C",X"43",X"55",X"4E",X"40",X"54",X"53",X"41",X"4C",X"53",X"4E",X"4F",X"49",X"54",X"41",
		X"4C",X"55",X"54",X"41",X"52",X"47",X"4E",X"4F",X"43",X"45",X"48",X"54",X"40",X"48",X"54",X"49",
		X"57",X"40",X"44",X"45",X"44",X"49",X"4C",X"4C",X"4F",X"43",X"40",X"55",X"4F",X"59",X"4C",X"4C",
		X"41",X"57",X"40",X"54",X"4E",X"45",X"4D",X"4E",X"49",X"41",X"54",X"4E",X"4F",X"43",X"40",X"52",
		X"41",X"45",X"4C",X"43",X"55",X"4E",X"09",X"DD",X"2A",X"F6",X"4D",X"FD",X"CB",X"07",X"6E",X"C2",
		X"06",X"24",X"FD",X"CB",X"07",X"76",X"C8",X"7E",X"CB",X"BF",X"CB",X"B7",X"FE",X"03",X"CA",X"7B",
		X"23",X"3C",X"47",X"7E",X"E6",X"C0",X"B0",X"77",X"3E",X"F3",X"FD",X"46",X"03",X"90",X"32",X"5D",
		X"4C",X"FD",X"7E",X"04",X"D6",X"0C",X"32",X"5C",X"4C",X"E5",X"CD",X"B2",X"0E",X"E1",X"3A",X"0A",
		X"4C",X"FE",X"00",X"C2",X"5C",X"23",X"3A",X"0B",X"4C",X"FE",X"00",X"C2",X"5C",X"23",X"CB",X"76",
		X"C2",X"54",X"23",X"CB",X"F6",X"1A",X"32",X"0A",X"4E",X"D5",X"1B",X"1A",X"32",X"0B",X"4E",X"13",
		X"13",X"1A",X"32",X"0C",X"4E",X"3E",X"21",X"CD",X"D3",X"15",X"1A",X"32",X"0D",X"4E",X"3E",X"40",
		X"CD",X"BF",X"15",X"1A",X"32",X"0E",X"4E",X"D1",X"CB",X"7E",X"C2",X"F3",X"20",X"3A",X"9C",X"4E",
		X"FE",X"00",X"CA",X"F3",X"20",X"FE",X"01",X"28",X"02",X"18",X"56",X"3A",X"90",X"4C",X"CB",X"47",
		X"28",X"07",X"CB",X"5F",X"28",X"27",X"CB",X"B6",X"C9",X"FD",X"46",X"00",X"FD",X"36",X"00",X"02",
		X"3A",X"18",X"4E",X"FD",X"77",X"05",X"AF",X"32",X"9C",X"4E",X"78",X"FE",X"04",X"28",X"07",X"DD",
		X"7E",X"02",X"12",X"C3",X"BF",X"22",X"DD",X"7E",X"03",X"12",X"C3",X"BF",X"22",X"FD",X"46",X"00",
		X"FD",X"36",X"00",X"03",X"3A",X"17",X"4E",X"FD",X"77",X"05",X"AF",X"32",X"9C",X"4E",X"78",X"FE",
		X"04",X"28",X"07",X"DD",X"7E",X"04",X"12",X"C3",X"BF",X"22",X"DD",X"7E",X"05",X"12",X"C3",X"BF",
		X"22",X"3A",X"90",X"4C",X"CB",X"4F",X"28",X"07",X"CB",X"57",X"28",X"27",X"CB",X"B6",X"C9",X"FD",
		X"46",X"00",X"FD",X"36",X"00",X"05",X"3A",X"19",X"4E",X"FD",X"77",X"05",X"AF",X"32",X"9C",X"4E",
		X"78",X"FE",X"02",X"28",X"07",X"DD",X"7E",X"03",X"12",X"C3",X"95",X"21",X"DD",X"7E",X"05",X"12",
		X"C3",X"95",X"21",X"FD",X"46",X"00",X"FD",X"36",X"00",X"04",X"3A",X"1A",X"4E",X"FD",X"77",X"05",
		X"AF",X"32",X"9C",X"4E",X"78",X"FE",X"02",X"28",X"07",X"DD",X"7E",X"02",X"12",X"C3",X"95",X"21",
		X"DD",X"7E",X"04",X"12",X"C3",X"95",X"21",X"AF",X"32",X"9C",X"4E",X"C3",X"BF",X"22",X"AF",X"32",
		X"9C",X"4E",X"C3",X"BF",X"22",X"AF",X"32",X"9C",X"4E",X"C3",X"95",X"21",X"AF",X"32",X"9C",X"4E",
		X"C3",X"95",X"21",X"FD",X"7E",X"00",X"FE",X"02",X"CA",X"2A",X"22",X"FE",X"03",X"CA",X"2A",X"22",
		X"FD",X"CB",X"07",X"46",X"20",X"2F",X"3A",X"0A",X"4E",X"DD",X"BE",X"01",X"CA",X"17",X"21",X"FE",
		X"66",X"DA",X"A6",X"21",X"CD",X"45",X"29",X"CD",X"BA",X"29",X"FD",X"7E",X"00",X"FE",X"05",X"28",
		X"0A",X"DD",X"7E",X"03",X"32",X"0A",X"4E",X"12",X"C3",X"05",X"22",X"DD",X"7E",X"02",X"32",X"0A",
		X"4E",X"12",X"C3",X"05",X"22",X"FD",X"CB",X"07",X"5E",X"CA",X"5A",X"21",X"3A",X"0A",X"4E",X"DD",
		X"BE",X"01",X"CA",X"4D",X"21",X"FE",X"66",X"DA",X"A6",X"21",X"CD",X"45",X"29",X"CD",X"BA",X"29",
		X"DD",X"7E",X"07",X"32",X"0A",X"4E",X"12",X"C3",X"D7",X"21",X"3A",X"0A",X"4E",X"DD",X"BE",X"01",
		X"28",X"08",X"FE",X"66",X"DA",X"A6",X"21",X"CD",X"45",X"29",X"CD",X"BA",X"29",X"FD",X"7E",X"00",
		X"FE",X"05",X"28",X"29",X"DD",X"7E",X"05",X"32",X"0A",X"4E",X"12",X"3A",X"17",X"4E",X"FD",X"77",
		X"05",X"FD",X"36",X"00",X"03",X"3A",X"0C",X"4E",X"DD",X"BE",X"00",X"CA",X"AF",X"25",X"C3",X"FC",
		X"25",X"FD",X"CB",X"07",X"FE",X"FD",X"22",X"91",X"4C",X"CD",X"CE",X"0C",X"C9",X"DD",X"7E",X"04",
		X"32",X"0A",X"4E",X"12",X"18",X"D5",X"FD",X"7E",X"00",X"FE",X"05",X"28",X"11",X"3A",X"0A",X"4E",
		X"DD",X"BE",X"02",X"20",X"13",X"DD",X"7E",X"08",X"32",X"0A",X"4E",X"12",X"18",X"BD",X"3A",X"0A",
		X"4E",X"DD",X"BE",X"03",X"20",X"02",X"18",X"ED",X"3A",X"0A",X"4E",X"DD",X"BE",X"06",X"20",X"1F",
		X"DD",X"7E",X"08",X"32",X"0A",X"4E",X"12",X"FD",X"7E",X"00",X"FE",X"05",X"28",X"0C",X"3A",X"0D",
		X"4E",X"DD",X"BE",X"00",X"CA",X"99",X"25",X"C3",X"95",X"21",X"3A",X"0E",X"4E",X"18",X"F2",X"FD",
		X"7E",X"00",X"FE",X"05",X"28",X"25",X"3A",X"0A",X"4E",X"DD",X"BE",X"04",X"20",X"27",X"DD",X"7E",
		X"08",X"32",X"0A",X"4E",X"12",X"3A",X"18",X"4E",X"FD",X"77",X"05",X"FD",X"36",X"00",X"02",X"3A",
		X"0B",X"4E",X"DD",X"BE",X"00",X"CA",X"69",X"25",X"C3",X"DF",X"25",X"3A",X"0A",X"4E",X"DD",X"BE",
		X"05",X"20",X"02",X"18",X"D9",X"FD",X"CB",X"07",X"EE",X"C9",X"FD",X"CB",X"07",X"56",X"20",X"2F",
		X"3A",X"0A",X"4E",X"DD",X"BE",X"01",X"CA",X"41",X"22",X"FE",X"66",X"DA",X"D0",X"22",X"CD",X"45",
		X"29",X"CD",X"BA",X"29",X"FD",X"7E",X"00",X"FE",X"03",X"28",X"0A",X"DD",X"7E",X"04",X"32",X"0A",
		X"4E",X"12",X"C3",X"2F",X"23",X"DD",X"7E",X"02",X"32",X"0A",X"4E",X"12",X"C3",X"2F",X"23",X"FD",
		X"CB",X"07",X"4E",X"CA",X"84",X"22",X"3A",X"0A",X"4E",X"DD",X"BE",X"01",X"CA",X"77",X"22",X"FE",
		X"66",X"DA",X"D0",X"22",X"CD",X"45",X"29",X"CD",X"BA",X"29",X"DD",X"7E",X"06",X"32",X"0A",X"4E",
		X"12",X"C3",X"01",X"23",X"3A",X"0A",X"4E",X"DD",X"BE",X"01",X"28",X"08",X"FE",X"66",X"DA",X"D0",
		X"22",X"CD",X"45",X"29",X"CD",X"BA",X"29",X"FD",X"7E",X"00",X"FE",X"03",X"28",X"29",X"DD",X"7E",
		X"05",X"32",X"0A",X"4E",X"12",X"3A",X"19",X"4E",X"FD",X"77",X"05",X"FD",X"36",X"00",X"05",X"3A",
		X"0E",X"4E",X"DD",X"BE",X"00",X"CA",X"5F",X"26",X"C3",X"AC",X"26",X"FD",X"CB",X"07",X"FE",X"FD",
		X"22",X"91",X"4C",X"CD",X"CE",X"0C",X"C9",X"DD",X"7E",X"03",X"32",X"0A",X"4E",X"12",X"18",X"D5",
		X"FD",X"7E",X"00",X"FE",X"03",X"28",X"11",X"3A",X"0A",X"4E",X"DD",X"BE",X"02",X"20",X"13",X"DD",
		X"7E",X"08",X"32",X"0A",X"4E",X"12",X"18",X"BD",X"3A",X"0A",X"4E",X"DD",X"BE",X"04",X"20",X"02",
		X"18",X"ED",X"3A",X"0A",X"4E",X"DD",X"BE",X"07",X"20",X"1F",X"DD",X"7E",X"08",X"32",X"0A",X"4E",
		X"12",X"FD",X"7E",X"00",X"FE",X"03",X"28",X"0C",X"3A",X"0B",X"4E",X"DD",X"BE",X"00",X"CA",X"49",
		X"26",X"C3",X"BF",X"22",X"3A",X"0C",X"4E",X"18",X"F2",X"FD",X"7E",X"00",X"FE",X"03",X"28",X"25",
		X"3A",X"0A",X"4E",X"DD",X"BE",X"03",X"20",X"27",X"DD",X"7E",X"08",X"32",X"0A",X"4E",X"12",X"3A",
		X"1A",X"4E",X"FD",X"77",X"05",X"FD",X"36",X"00",X"04",X"3A",X"0D",X"4E",X"DD",X"BE",X"00",X"CA",
		X"19",X"26",X"C3",X"8F",X"26",X"3A",X"0A",X"4E",X"DD",X"BE",X"05",X"20",X"02",X"18",X"D9",X"FD",
		X"CB",X"07",X"EE",X"C9",X"FD",X"22",X"91",X"4C",X"CD",X"CE",X"0C",X"C9",X"CB",X"B6",X"CB",X"7E",
		X"20",X"F2",X"3A",X"9C",X"4E",X"FE",X"00",X"28",X"EB",X"FE",X"03",X"CA",X"D7",X"20",X"FE",X"04",
		X"CA",X"DE",X"20",X"FE",X"05",X"CA",X"E5",X"20",X"C3",X"EC",X"20",X"3E",X"C0",X"A6",X"77",X"CB",
		X"7F",X"20",X"2A",X"FD",X"7E",X"01",X"FE",X"00",X"C8",X"FD",X"CB",X"07",X"66",X"C2",X"C4",X"23",
		X"FD",X"7E",X"01",X"06",X"02",X"B8",X"CA",X"C8",X"1F",X"D6",X"02",X"FE",X"04",X"38",X"06",X"FD",
		X"77",X"01",X"C3",X"C8",X"1F",X"3E",X"02",X"FD",X"77",X"01",X"C3",X"C8",X"1F",X"FD",X"CB",X"07",
		X"7E",X"20",X"32",X"3A",X"16",X"4E",X"FD",X"46",X"01",X"B8",X"CA",X"C8",X"1F",X"04",X"FD",X"70",
		X"01",X"C3",X"C8",X"1F",X"3A",X"31",X"4E",X"FD",X"46",X"01",X"B8",X"CA",X"C8",X"1F",X"90",X"FE",
		X"02",X"38",X"09",X"78",X"C6",X"02",X"FD",X"77",X"01",X"C3",X"C8",X"1F",X"3A",X"31",X"4E",X"FD",
		X"77",X"01",X"C3",X"C8",X"1F",X"FD",X"CB",X"07",X"BE",X"FD",X"7E",X"01",X"FE",X"00",X"28",X"C3",
		X"3A",X"15",X"4E",X"FD",X"77",X"01",X"3A",X"8C",X"4D",X"FE",X"00",X"20",X"B6",X"E5",X"21",X"71",
		X"4D",X"CB",X"C6",X"E1",X"18",X"AD",X"23",X"7E",X"FE",X"02",X"20",X"1D",X"36",X"00",X"23",X"7E",
		X"FE",X"00",X"28",X"17",X"FE",X"28",X"CA",X"69",X"27",X"34",X"21",X"7C",X"27",X"CD",X"BA",X"15",
		X"7E",X"FD",X"77",X"05",X"FD",X"36",X"06",X"01",X"C9",X"34",X"C9",X"34",X"2B",X"2B",X"FD",X"CB",
		X"07",X"B6",X"CB",X"7E",X"28",X"35",X"3A",X"14",X"4E",X"FE",X"0D",X"D2",X"45",X"24",X"C6",X"04",
		X"32",X"14",X"4E",X"18",X"05",X"3E",X"10",X"32",X"14",X"4E",X"3A",X"13",X"4E",X"FE",X"0D",X"30",
		X"07",X"C6",X"04",X"32",X"13",X"4E",X"18",X"05",X"3E",X"10",X"32",X"13",X"4E",X"3A",X"20",X"4D",
		X"FE",X"00",X"20",X"B6",X"21",X"3B",X"4D",X"CB",X"C6",X"18",X"AF",X"21",X"56",X"4D",X"CB",X"C6",
		X"21",X"68",X"4C",X"CB",X"B6",X"21",X"70",X"4C",X"CB",X"B6",X"21",X"78",X"4C",X"CB",X"B6",X"21",
		X"80",X"4C",X"CB",X"B6",X"21",X"88",X"4C",X"CB",X"B6",X"21",X"90",X"4C",X"CB",X"AE",X"CB",X"B6",
		X"3E",X"B5",X"32",X"1B",X"4E",X"2A",X"9D",X"4E",X"E5",X"E5",X"D1",X"13",X"01",X"1F",X"00",X"36",
		X"00",X"ED",X"B0",X"D1",X"3A",X"34",X"4E",X"47",X"3A",X"32",X"4E",X"80",X"32",X"9F",X"4E",X"01",
		X"80",X"03",X"21",X"40",X"40",X"3A",X"9F",X"4E",X"ED",X"B1",X"78",X"B1",X"28",X"0A",X"2B",X"EB",
		X"73",X"23",X"72",X"23",X"EB",X"23",X"18",X"ED",X"3E",X"07",X"32",X"8F",X"4C",X"AF",X"32",X"64",
		X"4C",X"32",X"6C",X"4C",X"32",X"74",X"4C",X"32",X"7C",X"4C",X"32",X"84",X"4C",X"21",X"A4",X"27",
		X"7E",X"FE",X"FF",X"28",X"0D",X"32",X"8E",X"4C",X"23",X"E5",X"3E",X"02",X"CD",X"A5",X"15",X"E1",
		X"18",X"EE",X"AF",X"32",X"8C",X"4C",X"3A",X"E3",X"4E",X"CB",X"47",X"CA",X"39",X"25",X"AF",X"32",
		X"E3",X"4E",X"11",X"4E",X"40",X"21",X"4E",X"1F",X"3E",X"05",X"06",X"1C",X"CD",X"F5",X"15",X"11",
		X"4E",X"44",X"21",X"A6",X"1F",X"3E",X"05",X"06",X"1C",X"CD",X"F5",X"15",X"CD",X"14",X"16",X"11",
		X"CF",X"40",X"21",X"79",X"1F",X"3E",X"01",X"06",X"15",X"CD",X"DF",X"15",X"11",X"91",X"40",X"21",
		X"8E",X"1F",X"3E",X"01",X"06",X"18",X"CD",X"DF",X"15",X"3E",X"B4",X"CD",X"A5",X"15",X"21",X"90",
		X"4C",X"CB",X"AE",X"C9",X"21",X"61",X"4C",X"22",X"91",X"4C",X"CD",X"CE",X"0C",X"21",X"69",X"4C",
		X"22",X"91",X"4C",X"CD",X"CE",X"0C",X"21",X"71",X"4C",X"22",X"91",X"4C",X"CD",X"CE",X"0C",X"21",
		X"79",X"4C",X"22",X"91",X"4C",X"CD",X"CE",X"0C",X"C9",X"CB",X"7E",X"C2",X"25",X"22",X"3A",X"0A",
		X"4E",X"DD",X"BE",X"08",X"CA",X"FC",X"26",X"DD",X"BE",X"03",X"20",X"11",X"3A",X"1A",X"4E",X"FD",
		X"77",X"05",X"FD",X"36",X"00",X"04",X"DD",X"7E",X"07",X"12",X"C3",X"95",X"21",X"3A",X"19",X"4E",
		X"FD",X"77",X"05",X"FD",X"36",X"00",X"05",X"18",X"ED",X"CB",X"7E",X"C2",X"25",X"22",X"3A",X"0A",
		X"4E",X"DD",X"BE",X"08",X"CA",X"FC",X"26",X"3E",X"01",X"32",X"9C",X"4E",X"CB",X"B6",X"C9",X"CB",
		X"7E",X"C2",X"25",X"22",X"3A",X"0A",X"4E",X"DD",X"BE",X"08",X"CA",X"FC",X"26",X"DD",X"BE",X"05",
		X"20",X"11",X"3A",X"1A",X"4E",X"FD",X"77",X"05",X"FD",X"36",X"00",X"04",X"DD",X"7E",X"07",X"12",
		X"C3",X"95",X"21",X"3A",X"19",X"4E",X"FD",X"77",X"05",X"FD",X"36",X"00",X"05",X"18",X"ED",X"CB",
		X"7E",X"C2",X"91",X"21",X"3A",X"0A",X"4E",X"DD",X"BE",X"08",X"C2",X"95",X"21",X"FD",X"CB",X"07",
		X"46",X"CA",X"95",X"21",X"3E",X"03",X"32",X"9C",X"4E",X"C3",X"95",X"21",X"CB",X"7E",X"C2",X"91",
		X"21",X"3A",X"0A",X"4E",X"DD",X"BE",X"08",X"C2",X"95",X"21",X"FD",X"CB",X"07",X"5E",X"CA",X"95",
		X"21",X"3E",X"04",X"32",X"9C",X"4E",X"C3",X"95",X"21",X"CB",X"7E",X"C2",X"4F",X"23",X"3A",X"0A",
		X"4E",X"DD",X"BE",X"08",X"CA",X"FC",X"26",X"DD",X"BE",X"04",X"20",X"11",X"3A",X"18",X"4E",X"FD",
		X"77",X"05",X"FD",X"36",X"00",X"02",X"DD",X"7E",X"06",X"12",X"C3",X"BF",X"22",X"3A",X"17",X"4E",
		X"FD",X"77",X"05",X"FD",X"36",X"00",X"03",X"18",X"ED",X"CB",X"7E",X"C2",X"4F",X"23",X"3A",X"0A",
		X"4E",X"DD",X"BE",X"08",X"CA",X"FC",X"26",X"3E",X"02",X"32",X"9C",X"4E",X"CB",X"B6",X"C9",X"CB",
		X"7E",X"C2",X"4F",X"23",X"3A",X"0A",X"4E",X"DD",X"BE",X"08",X"CA",X"FC",X"26",X"DD",X"BE",X"05",
		X"20",X"11",X"3A",X"18",X"4E",X"FD",X"77",X"05",X"FD",X"36",X"00",X"02",X"DD",X"7E",X"06",X"12",
		X"C3",X"BF",X"22",X"3A",X"17",X"4E",X"FD",X"77",X"05",X"FD",X"36",X"00",X"03",X"18",X"ED",X"CB",
		X"7E",X"C2",X"BB",X"22",X"3A",X"0A",X"4E",X"DD",X"BE",X"08",X"C2",X"BF",X"22",X"FD",X"CB",X"07",
		X"56",X"CA",X"BF",X"22",X"3E",X"05",X"32",X"9C",X"4E",X"C3",X"BF",X"22",X"CB",X"7E",X"C2",X"BB",
		X"22",X"3A",X"0A",X"4E",X"DD",X"BE",X"08",X"C2",X"BF",X"22",X"FD",X"CB",X"07",X"4E",X"CA",X"BF",
		X"22",X"3E",X"06",X"32",X"9C",X"4E",X"C3",X"BF",X"22",X"FD",X"7E",X"07",X"47",X"FD",X"7E",X"00",
		X"FE",X"02",X"28",X"10",X"FE",X"03",X"28",X"14",X"FE",X"05",X"28",X"18",X"CB",X"48",X"CA",X"90",
		X"23",X"C3",X"B3",X"23",X"CB",X"58",X"CA",X"90",X"23",X"C3",X"B3",X"23",X"CB",X"40",X"CA",X"90",
		X"23",X"C3",X"B3",X"23",X"CB",X"50",X"CA",X"90",X"23",X"C3",X"B3",X"23",X"FD",X"CB",X"07",X"EE",
		X"CB",X"7E",X"C0",X"21",X"E3",X"4E",X"CB",X"C6",X"C9",X"05",X"20",X"00",X"E0",X"70",X"42",X"09",
		X"00",X"05",X"20",X"00",X"F0",X"70",X"3E",X"09",X"00",X"05",X"20",X"00",X"DF",X"60",X"3A",X"09",
		X"00",X"05",X"20",X"00",X"EF",X"60",X"36",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"20",X"00",X"02",X"70",X"2E",X"09",
		X"00",X"04",X"20",X"00",X"12",X"70",X"2A",X"09",X"00",X"04",X"20",X"00",X"01",X"60",X"26",X"09",
		X"00",X"04",X"20",X"00",X"11",X"60",X"22",X"09",X"00",X"04",X"20",X"00",X"FA",X"80",X"32",X"09",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"36",X"00",X"FD",X"CB",X"07",X"AE",X"FD",
		X"36",X"03",X"00",X"C9",X"5D",X"5C",X"60",X"62",X"5D",X"5C",X"60",X"62",X"04",X"08",X"0C",X"09",
		X"04",X"08",X"0C",X"09",X"10",X"14",X"18",X"15",X"10",X"14",X"18",X"15",X"1C",X"20",X"24",X"21",
		X"1C",X"20",X"24",X"21",X"28",X"2C",X"30",X"2D",X"28",X"2C",X"30",X"2D",X"34",X"38",X"3C",X"39",
		X"34",X"38",X"3C",X"39",X"04",X"08",X"0C",X"09",X"04",X"08",X"0C",X"09",X"10",X"14",X"18",X"15",
		X"10",X"14",X"18",X"15",X"1C",X"20",X"24",X"21",X"1C",X"20",X"24",X"21",X"28",X"2C",X"30",X"2D",
		X"28",X"2C",X"30",X"2D",X"34",X"38",X"3C",X"39",X"34",X"38",X"3C",X"39",X"FF",X"FD",X"CB",X"07",
		X"76",X"C8",X"FD",X"7E",X"00",X"FE",X"04",X"DA",X"3E",X"28",X"DD",X"7E",X"03",X"FD",X"BE",X"03",
		X"DA",X"2B",X"28",X"CA",X"3E",X"28",X"FD",X"7E",X"00",X"FE",X"05",X"CA",X"5D",X"28",X"FD",X"7E",
		X"07",X"F6",X"1F",X"E6",X"FB",X"FD",X"77",X"07",X"DD",X"7E",X"03",X"FD",X"46",X"03",X"90",X"FE",
		X"05",X"38",X"05",X"FE",X"FB",X"30",X"01",X"C9",X"DD",X"7E",X"04",X"FD",X"46",X"04",X"90",X"FE",
		X"05",X"38",X"05",X"FE",X"FB",X"30",X"01",X"C9",X"DD",X"CB",X"07",X"EE",X"FD",X"CB",X"07",X"EE",
		X"C9",X"FD",X"7E",X"03",X"DD",X"BE",X"03",X"38",X"C5",X"18",X"07",X"FD",X"7E",X"00",X"FE",X"04",
		X"28",X"2B",X"FD",X"7E",X"07",X"F6",X"1F",X"E6",X"FD",X"FD",X"77",X"07",X"18",X"BA",X"DD",X"7E",
		X"04",X"FD",X"BE",X"04",X"38",X"21",X"CA",X"DA",X"27",X"FD",X"7E",X"00",X"FE",X"02",X"28",X"D1",
		X"FD",X"7E",X"07",X"F6",X"1F",X"E6",X"F7",X"FD",X"77",X"07",X"C3",X"F8",X"27",X"FD",X"7E",X"04",
		X"DD",X"BE",X"04",X"38",X"EB",X"18",X"07",X"FD",X"7E",X"00",X"FE",X"03",X"28",X"B3",X"FD",X"7E",
		X"07",X"F6",X"1F",X"E6",X"FE",X"FD",X"77",X"07",X"C3",X"F8",X"27",X"FD",X"7E",X"03",X"FE",X"00",
		X"C8",X"DD",X"21",X"69",X"4C",X"DD",X"7E",X"03",X"FE",X"00",X"28",X"03",X"CD",X"E1",X"28",X"DD",
		X"21",X"71",X"4C",X"DD",X"7E",X"03",X"FE",X"00",X"28",X"03",X"CD",X"E1",X"28",X"DD",X"21",X"79",
		X"4C",X"DD",X"7E",X"03",X"FE",X"00",X"C8",X"CD",X"E1",X"28",X"C9",X"FD",X"7E",X"03",X"FE",X"00",
		X"C8",X"DD",X"21",X"71",X"4C",X"DD",X"7E",X"03",X"FE",X"00",X"28",X"03",X"CD",X"E1",X"28",X"DD",
		X"21",X"79",X"4C",X"DD",X"7E",X"03",X"FE",X"00",X"C8",X"CD",X"E1",X"28",X"C9",X"FD",X"7E",X"03",
		X"FE",X"00",X"C8",X"DD",X"21",X"79",X"4C",X"DD",X"7E",X"03",X"FE",X"00",X"C8",X"CD",X"E1",X"28",
		X"C9",X"DD",X"7E",X"00",X"FD",X"86",X"00",X"FE",X"05",X"28",X"05",X"FE",X"09",X"28",X"2A",X"C9",
		X"DD",X"7E",X"04",X"FD",X"96",X"04",X"DD",X"7E",X"00",X"FA",X"14",X"29",X"FE",X"02",X"C0",X"DD",
		X"7E",X"07",X"F6",X"0F",X"EE",X"04",X"DD",X"77",X"07",X"FD",X"7E",X"07",X"F6",X"0F",X"EE",X"02",
		X"FD",X"77",X"07",X"C9",X"FE",X"03",X"C0",X"18",X"E6",X"DD",X"7E",X"03",X"FD",X"96",X"03",X"DD",
		X"7E",X"00",X"FA",X"40",X"29",X"DD",X"7E",X"00",X"FE",X"05",X"C0",X"DD",X"7E",X"07",X"F6",X"0F",
		X"EE",X"01",X"DD",X"77",X"07",X"FD",X"7E",X"07",X"F6",X"0F",X"EE",X"08",X"FD",X"77",X"07",X"C9",
		X"FE",X"04",X"C0",X"18",X"E6",X"3A",X"29",X"4E",X"3C",X"32",X"29",X"4E",X"E5",X"21",X"00",X"04",
		X"19",X"3A",X"40",X"44",X"77",X"E1",X"CB",X"7E",X"20",X"48",X"2A",X"93",X"4C",X"7E",X"21",X"AE",
		X"29",X"CD",X"BA",X"15",X"7E",X"32",X"2D",X"4E",X"3E",X"40",X"32",X"86",X"4C",X"AF",X"32",X"2B",
		X"4E",X"32",X"2C",X"4E",X"3A",X"8C",X"4C",X"32",X"84",X"4C",X"3A",X"8D",X"4C",X"32",X"85",X"4C",
		X"D5",X"23",X"5E",X"23",X"56",X"2A",X"AE",X"4C",X"19",X"22",X"AE",X"4C",X"D1",X"21",X"8C",X"4D",
		X"CB",X"C6",X"AF",X"32",X"2B",X"4E",X"3A",X"29",X"4E",X"FE",X"10",X"C0",X"3E",X"FF",X"32",X"29",
		X"4E",X"C9",X"3A",X"29",X"4E",X"FE",X"10",X"C0",X"EB",X"22",X"E0",X"4E",X"EB",X"C9",X"44",X"00",
		X"10",X"48",X"00",X"20",X"4C",X"00",X"40",X"50",X"00",X"80",X"D5",X"E5",X"2A",X"0F",X"4E",X"ED",
		X"5B",X"AE",X"4C",X"19",X"22",X"AE",X"4C",X"E1",X"D1",X"C9",X"DD",X"21",X"16",X"32",X"DD",X"22",
		X"F6",X"4D",X"21",X"84",X"33",X"3E",X"1A",X"CD",X"BD",X"2E",X"CD",X"D1",X"34",X"3E",X"0E",X"32",
		X"E2",X"4E",X"3E",X"81",X"21",X"FD",X"2D",X"CD",X"EF",X"30",X"21",X"10",X"00",X"22",X"11",X"4E",
		X"3E",X"04",X"32",X"13",X"4E",X"3E",X"08",X"32",X"14",X"4E",X"3E",X"10",X"32",X"31",X"4E",X"21",
		X"F6",X"30",X"CD",X"28",X"2F",X"CD",X"31",X"2F",X"11",X"6F",X"41",X"21",X"D6",X"2F",X"3E",X"01",
		X"06",X"0B",X"CD",X"DF",X"15",X"11",X"11",X"41",X"21",X"E1",X"2F",X"3E",X"01",X"06",X"11",X"CD",
		X"DF",X"15",X"C9",X"DD",X"21",X"16",X"32",X"DD",X"22",X"F6",X"4D",X"21",X"84",X"33",X"3E",X"1A",
		X"CD",X"BD",X"2E",X"CD",X"D1",X"34",X"3E",X"0E",X"32",X"E2",X"4E",X"3E",X"87",X"21",X"FD",X"2D",
		X"CD",X"EF",X"30",X"21",X"20",X"00",X"22",X"11",X"4E",X"3E",X"05",X"32",X"13",X"4E",X"3E",X"0A",
		X"32",X"14",X"4E",X"3E",X"10",X"32",X"31",X"4E",X"21",X"F6",X"30",X"CD",X"28",X"2F",X"CD",X"31",
		X"2F",X"11",X"6F",X"41",X"21",X"D6",X"2F",X"3E",X"01",X"06",X"0B",X"CD",X"DF",X"15",X"11",X"11",
		X"41",X"21",X"F2",X"2F",X"3E",X"01",X"06",X"10",X"CD",X"DF",X"15",X"C9",X"DD",X"21",X"1F",X"32",
		X"DD",X"22",X"F6",X"4D",X"21",X"7A",X"32",X"3E",X"19",X"CD",X"BD",X"2E",X"CD",X"2A",X"35",X"3E",
		X"0E",X"32",X"E2",X"4E",X"3E",X"75",X"21",X"1D",X"2E",X"CD",X"EF",X"30",X"21",X"30",X"00",X"22",
		X"11",X"4E",X"3E",X"07",X"32",X"13",X"4E",X"3E",X"0C",X"32",X"14",X"4E",X"3E",X"0F",X"32",X"31",
		X"4E",X"21",X"26",X"31",X"CD",X"28",X"2F",X"CD",X"31",X"2F",X"11",X"6F",X"41",X"21",X"02",X"30",
		X"3E",X"01",X"06",X"0B",X"CD",X"DF",X"15",X"11",X"31",X"41",X"21",X"0D",X"30",X"3E",X"01",X"06",
		X"0F",X"CD",X"DF",X"15",X"C9",X"DD",X"21",X"1F",X"32",X"DD",X"22",X"F6",X"4D",X"21",X"7A",X"32",
		X"3E",X"19",X"CD",X"BD",X"2E",X"CD",X"2A",X"35",X"3E",X"0E",X"32",X"E2",X"4E",X"3E",X"78",X"21",
		X"1D",X"2E",X"CD",X"EF",X"30",X"21",X"40",X"00",X"22",X"11",X"4E",X"3E",X"09",X"32",X"13",X"4E",
		X"3E",X"0D",X"32",X"14",X"4E",X"3E",X"0F",X"32",X"31",X"4E",X"21",X"26",X"31",X"CD",X"28",X"2F",
		X"CD",X"31",X"2F",X"11",X"6F",X"41",X"21",X"02",X"30",X"3E",X"01",X"06",X"0B",X"CD",X"DF",X"15",
		X"11",X"31",X"41",X"21",X"1C",X"30",X"3E",X"01",X"06",X"0E",X"CD",X"DF",X"15",X"C9",X"DD",X"21",
		X"1F",X"32",X"DD",X"22",X"F6",X"4D",X"21",X"11",X"33",X"3E",X"1A",X"CD",X"BD",X"2E",X"CD",X"53",
		X"35",X"3E",X"10",X"32",X"E2",X"4E",X"3E",X"72",X"21",X"3D",X"2E",X"CD",X"EF",X"30",X"21",X"50",
		X"00",X"22",X"11",X"4E",X"3E",X"0A",X"32",X"13",X"4E",X"3E",X"0E",X"32",X"14",X"4E",X"3E",X"0F",
		X"32",X"31",X"4E",X"21",X"56",X"31",X"CD",X"28",X"2F",X"CD",X"31",X"2F",X"11",X"8F",X"41",X"21",
		X"2A",X"30",X"3E",X"01",X"06",X"09",X"CD",X"DF",X"15",X"11",X"F1",X"40",X"21",X"33",X"30",X"3E",
		X"01",X"06",X"12",X"CD",X"DF",X"15",X"C9",X"DD",X"21",X"1F",X"32",X"DD",X"22",X"F6",X"4D",X"21",
		X"11",X"33",X"3E",X"1A",X"CD",X"BD",X"2E",X"CD",X"53",X"35",X"3E",X"10",X"32",X"E2",X"4E",X"3E",
		X"6F",X"21",X"3D",X"2E",X"CD",X"EF",X"30",X"21",X"60",X"00",X"22",X"11",X"4E",X"3E",X"0B",X"32",
		X"13",X"4E",X"3E",X"0E",X"32",X"14",X"4E",X"3E",X"0F",X"32",X"31",X"4E",X"21",X"56",X"31",X"CD",
		X"28",X"2F",X"CD",X"31",X"2F",X"11",X"8F",X"41",X"21",X"2A",X"30",X"3E",X"01",X"06",X"09",X"CD",
		X"DF",X"15",X"11",X"11",X"41",X"21",X"45",X"30",X"3E",X"01",X"06",X"11",X"CD",X"DF",X"15",X"C9",
		X"DD",X"21",X"1F",X"32",X"DD",X"22",X"F6",X"4D",X"21",X"AF",X"34",X"3E",X"1A",X"CD",X"BD",X"2E",
		X"3E",X"0E",X"32",X"E2",X"4E",X"3E",X"84",X"21",X"5D",X"2E",X"CD",X"EF",X"30",X"21",X"70",X"00",
		X"22",X"11",X"4E",X"3E",X"0C",X"32",X"13",X"4E",X"3E",X"0F",X"32",X"14",X"4E",X"3E",X"0F",X"32",
		X"31",X"4E",X"21",X"86",X"31",X"CD",X"28",X"2F",X"CD",X"31",X"2F",X"11",X"4F",X"41",X"21",X"56",
		X"30",X"3E",X"01",X"06",X"0C",X"CD",X"DF",X"15",X"11",X"11",X"41",X"21",X"62",X"30",X"3E",X"01",
		X"06",X"10",X"CD",X"DF",X"15",X"C9",X"DD",X"21",X"1F",X"32",X"DD",X"22",X"F6",X"4D",X"21",X"AF",
		X"34",X"3E",X"1A",X"CD",X"BD",X"2E",X"3E",X"0E",X"32",X"E2",X"4E",X"3E",X"6C",X"21",X"5D",X"2E",
		X"CD",X"EF",X"30",X"21",X"80",X"00",X"22",X"11",X"4E",X"3E",X"0D",X"32",X"13",X"4E",X"3E",X"10",
		X"32",X"14",X"4E",X"3E",X"0F",X"32",X"31",X"4E",X"21",X"86",X"31",X"CD",X"28",X"2F",X"CD",X"31",
		X"2F",X"11",X"4F",X"41",X"21",X"56",X"30",X"3E",X"01",X"06",X"0C",X"CD",X"DF",X"15",X"11",X"31",
		X"41",X"21",X"72",X"30",X"3E",X"01",X"06",X"0F",X"CD",X"DF",X"15",X"C9",X"DD",X"21",X"1F",X"32",
		X"DD",X"22",X"F6",X"4D",X"21",X"51",X"34",X"3E",X"19",X"CD",X"BD",X"2E",X"CD",X"A0",X"35",X"3E",
		X"10",X"32",X"E2",X"4E",X"3E",X"75",X"21",X"7D",X"2E",X"CD",X"EF",X"30",X"21",X"90",X"00",X"22",
		X"11",X"4E",X"3E",X"0E",X"32",X"13",X"4E",X"3E",X"10",X"32",X"14",X"4E",X"3E",X"0E",X"32",X"31",
		X"4E",X"21",X"B6",X"31",X"CD",X"28",X"2F",X"CD",X"31",X"2F",X"11",X"6F",X"41",X"21",X"81",X"30",
		X"3E",X"01",X"06",X"0A",X"CD",X"DF",X"15",X"11",X"11",X"41",X"21",X"8B",X"30",X"3E",X"01",X"06",
		X"11",X"CD",X"DF",X"15",X"C9",X"DD",X"21",X"1F",X"32",X"DD",X"22",X"F6",X"4D",X"21",X"51",X"34",
		X"3E",X"19",X"CD",X"BD",X"2E",X"CD",X"A0",X"35",X"3E",X"10",X"32",X"E2",X"4E",X"3E",X"7B",X"21",
		X"7D",X"2E",X"CD",X"EF",X"30",X"21",X"00",X"01",X"22",X"11",X"4E",X"3E",X"0F",X"32",X"13",X"4E",
		X"3E",X"10",X"32",X"14",X"4E",X"3E",X"0E",X"32",X"31",X"4E",X"21",X"B6",X"31",X"CD",X"28",X"2F",
		X"CD",X"31",X"2F",X"11",X"6F",X"41",X"21",X"81",X"30",X"3E",X"01",X"06",X"0A",X"CD",X"DF",X"15",
		X"11",X"11",X"41",X"21",X"9C",X"30",X"3E",X"01",X"06",X"10",X"CD",X"DF",X"15",X"C9",X"DD",X"21",
		X"16",X"32",X"DD",X"22",X"F6",X"4D",X"21",X"28",X"32",X"3E",X"1A",X"CD",X"BD",X"2E",X"CD",X"C1",
		X"35",X"3E",X"10",X"32",X"E2",X"4E",X"3E",X"7E",X"21",X"9D",X"2E",X"CD",X"EF",X"30",X"21",X"10",
		X"01",X"22",X"11",X"4E",X"3E",X"10",X"32",X"13",X"4E",X"3E",X"10",X"32",X"14",X"4E",X"3E",X"0D",
		X"32",X"31",X"4E",X"21",X"E6",X"31",X"CD",X"28",X"2F",X"CD",X"31",X"2F",X"11",X"70",X"41",X"21",
		X"AC",X"30",X"3E",X"01",X"06",X"0B",X"CD",X"DF",X"15",X"C9",X"DD",X"21",X"16",X"32",X"DD",X"22",
		X"F6",X"4D",X"21",X"28",X"32",X"3E",X"1A",X"CD",X"BD",X"2E",X"CD",X"C1",X"35",X"3E",X"10",X"32",
		X"E2",X"4E",X"3E",X"66",X"21",X"9D",X"2E",X"CD",X"EF",X"30",X"21",X"20",X"01",X"22",X"11",X"4E",
		X"3E",X"10",X"32",X"13",X"4E",X"3E",X"10",X"32",X"14",X"4E",X"3E",X"0C",X"32",X"31",X"4E",X"21",
		X"E6",X"31",X"CD",X"28",X"2F",X"CD",X"31",X"2F",X"11",X"70",X"41",X"21",X"AC",X"30",X"3E",X"01",
		X"06",X"0B",X"CD",X"DF",X"15",X"C9",X"C9",X"C9",X"C9",X"C9",X"61",X"47",X"4F",X"52",X"4B",X"41",
		X"4E",X"53",X"2C",X"43",X"4F",X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"20",X"31",X"39",X"38",
		X"33",X"54",X"45",X"43",X"48",X"53",X"54",X"41",X"52",X"20",X"49",X"4E",X"43",X"A3",X"40",X"BC",
		X"40",X"8C",X"41",X"93",X"41",X"6C",X"42",X"73",X"42",X"43",X"43",X"5C",X"43",X"8B",X"40",X"94",
		X"40",X"A4",X"41",X"BB",X"41",X"44",X"42",X"5B",X"42",X"6B",X"43",X"74",X"43",X"AC",X"40",X"B3",
		X"40",X"29",X"41",X"36",X"41",X"C9",X"42",X"D6",X"42",X"4C",X"43",X"53",X"43",X"23",X"41",X"3C",
		X"41",X"8D",X"41",X"92",X"41",X"6D",X"42",X"72",X"42",X"C3",X"42",X"DC",X"42",X"CD",X"40",X"D2",
		X"40",X"46",X"41",X"59",X"41",X"A6",X"42",X"B9",X"42",X"2D",X"43",X"32",X"43",X"A3",X"40",X"BC",
		X"40",X"8A",X"41",X"95",X"41",X"6A",X"42",X"75",X"42",X"43",X"43",X"5C",X"43",X"AB",X"40",X"B4",
		X"40",X"2C",X"41",X"33",X"41",X"CC",X"42",X"D3",X"42",X"4B",X"43",X"54",X"43",X"CD",X"41",X"D2",
		X"41",X"88",X"41",X"97",X"41",X"68",X"42",X"77",X"42",X"2D",X"42",X"32",X"42",X"C5",X"40",X"DA",
		X"40",X"8B",X"41",X"94",X"41",X"6B",X"42",X"74",X"42",X"25",X"43",X"3A",X"43",X"EC",X"40",X"F3",
		X"40",X"28",X"41",X"37",X"41",X"C8",X"42",X"D7",X"42",X"0C",X"43",X"13",X"43",X"C4",X"40",X"DB",
		X"40",X"2C",X"41",X"33",X"41",X"CC",X"42",X"D3",X"42",X"24",X"43",X"3B",X"43",X"89",X"40",X"96",
		X"40",X"A8",X"41",X"B7",X"41",X"48",X"42",X"57",X"42",X"69",X"43",X"76",X"43",X"E5",X"CD",X"17",
		X"15",X"11",X"40",X"40",X"E1",X"D5",X"11",X"DF",X"4D",X"ED",X"A0",X"ED",X"A0",X"ED",X"A0",X"7E",
		X"FE",X"0F",X"38",X"F5",X"ED",X"A0",X"2B",X"D1",X"E5",X"21",X"DF",X"4D",X"23",X"46",X"DD",X"7E",
		X"00",X"12",X"13",X"10",X"FC",X"7E",X"23",X"86",X"2B",X"77",X"23",X"23",X"7E",X"FE",X"F0",X"30",
		X"18",X"12",X"13",X"23",X"46",X"DD",X"7E",X"01",X"12",X"13",X"10",X"FC",X"7E",X"23",X"86",X"2B",
		X"77",X"23",X"23",X"7E",X"12",X"13",X"C3",X"DC",X"2E",X"21",X"DF",X"4D",X"3A",X"F5",X"4D",X"3C",
		X"32",X"F5",X"4D",X"FE",X"1C",X"28",X"0B",X"7E",X"3D",X"77",X"FE",X"F1",X"D2",X"DC",X"2E",X"C3",
		X"C4",X"2E",X"E1",X"AF",X"32",X"F5",X"4D",X"C9",X"11",X"61",X"4C",X"01",X"30",X"00",X"ED",X"B0",
		X"C9",X"21",X"F8",X"4D",X"11",X"F9",X"4D",X"36",X"00",X"01",X"11",X"00",X"ED",X"B0",X"21",X"FB",
		X"4D",X"CB",X"FE",X"21",X"FE",X"4D",X"CB",X"FE",X"21",X"01",X"4E",X"CB",X"FE",X"21",X"04",X"4E",
		X"CB",X"FE",X"21",X"07",X"4E",X"CB",X"FE",X"AF",X"32",X"1B",X"4E",X"32",X"29",X"4E",X"32",X"2B",
		X"4E",X"32",X"32",X"4E",X"32",X"33",X"4E",X"21",X"00",X"00",X"22",X"AE",X"4C",X"3A",X"04",X"4D",
		X"17",X"21",X"B7",X"30",X"CD",X"BA",X"15",X"7E",X"32",X"30",X"40",X"23",X"7E",X"32",X"2F",X"40",
		X"3E",X"01",X"32",X"30",X"44",X"32",X"2F",X"44",X"3E",X"40",X"32",X"27",X"4E",X"32",X"28",X"4E",
		X"AF",X"32",X"E4",X"4E",X"21",X"DD",X"4D",X"CB",X"86",X"AF",X"32",X"9C",X"4E",X"06",X"14",X"21",
		X"CE",X"40",X"11",X"37",X"4E",X"C5",X"01",X"05",X"00",X"ED",X"B0",X"3E",X"1B",X"CD",X"BA",X"15",
		X"C1",X"10",X"F2",X"3A",X"40",X"44",X"32",X"9B",X"4E",X"11",X"CE",X"40",X"21",X"D5",X"2F",X"3E",
		X"05",X"06",X"14",X"CD",X"F5",X"15",X"11",X"CE",X"44",X"21",X"D4",X"2F",X"3E",X"05",X"06",X"14",
		X"CD",X"F5",X"15",X"C9",X"09",X"40",X"45",X"53",X"41",X"42",X"40",X"44",X"49",X"4F",X"52",X"55",
		X"51",X"47",X"47",X"49",X"4F",X"52",X"4B",X"40",X"4F",X"54",X"40",X"53",X"45",X"56",X"41",X"57",
		X"40",X"32",X"47",X"47",X"49",X"4F",X"52",X"4B",X"40",X"4F",X"54",X"40",X"45",X"56",X"41",X"57",
		X"40",X"31",X"45",X"53",X"41",X"42",X"40",X"47",X"47",X"49",X"4F",X"52",X"4B",X"4E",X"55",X"52",
		X"44",X"40",X"4F",X"54",X"40",X"53",X"45",X"56",X"41",X"57",X"40",X"32",X"4E",X"55",X"52",X"44",
		X"40",X"4F",X"54",X"40",X"45",X"56",X"41",X"57",X"40",X"31",X"45",X"53",X"41",X"42",X"40",X"4E",
		X"55",X"52",X"44",X"50",X"4C",X"4F",X"54",X"52",X"45",X"47",X"40",X"4F",X"54",X"40",X"53",X"45",
		X"56",X"41",X"57",X"40",X"32",X"50",X"4C",X"4F",X"54",X"52",X"45",X"47",X"40",X"4F",X"54",X"40",
		X"45",X"56",X"41",X"57",X"40",X"31",X"45",X"53",X"41",X"42",X"40",X"50",X"4C",X"4F",X"54",X"52",
		X"45",X"47",X"44",X"49",X"55",X"52",X"50",X"40",X"4F",X"54",X"40",X"53",X"45",X"56",X"41",X"57",
		X"40",X"32",X"44",X"49",X"55",X"52",X"50",X"40",X"4F",X"54",X"40",X"45",X"56",X"41",X"57",X"40",
		X"31",X"45",X"53",X"41",X"42",X"40",X"44",X"49",X"55",X"52",X"50",X"4E",X"41",X"4B",X"52",X"4F",
		X"47",X"40",X"4F",X"54",X"40",X"53",X"45",X"56",X"41",X"57",X"40",X"32",X"4E",X"41",X"4B",X"52",
		X"4F",X"47",X"40",X"4F",X"54",X"40",X"45",X"56",X"41",X"57",X"40",X"31",X"45",X"53",X"41",X"42",
		X"40",X"4E",X"41",X"4B",X"52",X"4F",X"47",X"40",X"01",X"40",X"02",X"40",X"03",X"40",X"04",X"40",
		X"05",X"40",X"06",X"40",X"07",X"40",X"08",X"40",X"09",X"01",X"00",X"01",X"01",X"01",X"02",X"01",
		X"03",X"01",X"04",X"01",X"05",X"01",X"06",X"01",X"07",X"01",X"08",X"01",X"09",X"02",X"00",X"02",
		X"01",X"02",X"02",X"02",X"03",X"02",X"04",X"02",X"05",X"02",X"06",X"02",X"07",X"02",X"08",X"32",
		X"34",X"4E",X"22",X"2F",X"4E",X"C9",X"03",X"02",X"00",X"3B",X"14",X"5D",X"07",X"5F",X"03",X"02",
		X"00",X"63",X"14",X"5D",X"07",X"1F",X"03",X"02",X"00",X"AB",X"14",X"5D",X"07",X"1F",X"03",X"02",
		X"00",X"D3",X"14",X"5D",X"07",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"02",X"04",
		X"00",X"8B",X"E4",X"5C",X"01",X"40",X"04",X"02",X"00",X"5B",X"3C",X"62",X"07",X"5F",X"03",X"02",
		X"00",X"D3",X"5C",X"5D",X"07",X"1F",X"02",X"02",X"00",X"3B",X"B4",X"5C",X"07",X"1F",X"05",X"02",
		X"00",X"B3",X"D4",X"60",X"07",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"02",X"04",
		X"00",X"8B",X"FC",X"5C",X"01",X"40",X"04",X"02",X"00",X"23",X"84",X"62",X"07",X"5F",X"03",X"02",
		X"00",X"73",X"24",X"5D",X"07",X"1F",X"03",X"02",X"00",X"9B",X"24",X"5D",X"07",X"1F",X"05",X"02",
		X"00",X"EB",X"84",X"60",X"07",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"02",X"04",
		X"00",X"8B",X"EC",X"5C",X"01",X"40",X"04",X"02",X"00",X"23",X"94",X"62",X"07",X"5F",X"04",X"02",
		X"00",X"23",X"7C",X"62",X"07",X"1F",X"05",X"02",X"00",X"EB",X"7C",X"60",X"07",X"1F",X"05",X"02",
		X"00",X"EB",X"94",X"60",X"07",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"02",X"04",
		X"00",X"8B",X"FC",X"5C",X"01",X"40",X"04",X"02",X"00",X"23",X"D4",X"62",X"07",X"5F",X"04",X"02",
		X"00",X"23",X"3C",X"62",X"07",X"1F",X"05",X"02",X"00",X"EB",X"3C",X"60",X"07",X"1F",X"05",X"02",
		X"00",X"EB",X"D4",X"60",X"07",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"02",X"04",
		X"00",X"8B",X"E4",X"5C",X"01",X"40",X"02",X"02",X"00",X"43",X"FC",X"5C",X"07",X"5F",X"02",X"02",
		X"00",X"5B",X"FC",X"5C",X"07",X"1F",X"02",X"02",X"00",X"B3",X"FC",X"5C",X"07",X"1F",X"02",X"02",
		X"00",X"CB",X"FC",X"5C",X"07",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"02",X"04",
		X"00",X"8B",X"DC",X"5C",X"01",X"40",X"65",X"0A",X"0B",X"0C",X"0D",X"0E",X"0F",X"10",X"14",X"65",
		X"0A",X"0B",X"0C",X"0D",X"0E",X"0F",X"10",X"16",X"F1",X"20",X"00",X"F4",X"04",X"FF",X"0B",X"06",
		X"02",X"0D",X"08",X"FE",X"0B",X"06",X"02",X"0D",X"04",X"FF",X"F4",X"01",X"00",X"0A",X"1C",X"00",
		X"0A",X"01",X"00",X"F4",X"01",X"01",X"0C",X"1C",X"FE",X"0E",X"01",X"01",X"F2",X"05",X"00",X"0A",
		X"14",X"00",X"0A",X"05",X"00",X"F4",X"04",X"FF",X"0B",X"16",X"02",X"0D",X"04",X"FF",X"F4",X"01",
		X"00",X"0A",X"1C",X"00",X"0A",X"01",X"00",X"F4",X"01",X"01",X"0C",X"0C",X"FE",X"0E",X"02",X"02",
		X"0C",X"0C",X"FE",X"0E",X"01",X"01",X"F1",X"20",X"00",X"FF",X"F1",X"20",X"00",X"F3",X"07",X"01",
		X"0C",X"10",X"FE",X"0E",X"07",X"01",X"F1",X"0A",X"00",X"0A",X"0A",X"00",X"0A",X"0A",X"00",X"F1",
		X"09",X"00",X"0B",X"0C",X"00",X"0D",X"09",X"00",X"F2",X"01",X"00",X"0A",X"02",X"01",X"0D",X"03",
		X"FE",X"0B",X"0E",X"02",X"0D",X"03",X"FE",X"0B",X"02",X"01",X"0A",X"01",X"00",X"F4",X"01",X"00",
		X"0A",X"1C",X"00",X"0A",X"01",X"00",X"F2",X"01",X"00",X"0A",X"0C",X"FF",X"0E",X"02",X"02",X"0C",
		X"0C",X"FF",X"0A",X"01",X"00",X"F2",X"01",X"00",X"0A",X"0B",X"01",X"0D",X"04",X"FE",X"0B",X"0B",
		X"01",X"0A",X"01",X"00",X"F4",X"01",X"00",X"0A",X"1C",X"00",X"0A",X"01",X"00",X"F2",X"01",X"00",
		X"0A",X"03",X"FF",X"0E",X"01",X"02",X"0C",X"10",X"FE",X"0E",X"01",X"02",X"0C",X"03",X"FF",X"0A",
		X"01",X"00",X"F1",X"09",X"00",X"0C",X"0C",X"00",X"0E",X"09",X"00",X"F1",X"0A",X"00",X"0A",X"0A",
		X"00",X"0A",X"0A",X"00",X"F3",X"09",X"FF",X"0B",X"0C",X"02",X"0D",X"09",X"FF",X"F1",X"20",X"00",
		X"FF",X"F1",X"20",X"00",X"F4",X"01",X"00",X"0A",X"02",X"01",X"0D",X"08",X"FE",X"0B",X"04",X"02",
		X"0D",X"08",X"FE",X"0B",X"02",X"01",X"0A",X"01",X"00",X"F1",X"02",X"00",X"0C",X"1A",X"00",X"0E",
		X"02",X"00",X"F5",X"03",X"00",X"0A",X"18",X"00",X"0A",X"03",X"00",X"F3",X"03",X"00",X"0A",X"0A",
		X"FF",X"0E",X"02",X"02",X"0C",X"0A",X"FF",X"0A",X"03",X"00",X"F3",X"03",X"00",X"0A",X"08",X"01",
		X"0D",X"06",X"FE",X"0B",X"08",X"01",X"0A",X"03",X"00",X"F5",X"03",X"00",X"0A",X"18",X"00",X"0A",
		X"03",X"00",X"F1",X"02",X"00",X"0B",X"1A",X"00",X"0D",X"02",X"00",X"F4",X"01",X"00",X"0A",X"05",
		X"FF",X"0E",X"02",X"02",X"0C",X"0A",X"FE",X"0E",X"02",X"02",X"0C",X"05",X"FF",X"0A",X"01",X"00",
		X"F1",X"20",X"00",X"FF",X"F1",X"20",X"00",X"F3",X"03",X"FF",X"0B",X"08",X"02",X"0D",X"06",X"FE",
		X"0B",X"08",X"02",X"0D",X"03",X"FF",X"F1",X"01",X"00",X"0A",X"1C",X"00",X"0A",X"01",X"00",X"F2",
		X"01",X"00",X"0A",X"04",X"FF",X"0E",X"02",X"02",X"0C",X"0C",X"FE",X"0E",X"02",X"02",X"0C",X"04",
		X"FF",X"0A",X"01",X"00",X"F2",X"01",X"00",X"0A",X"03",X"01",X"0D",X"04",X"FE",X"0B",X"0A",X"02",
		X"0D",X"04",X"FE",X"0B",X"03",X"01",X"0A",X"01",X"00",X"F1",X"01",X"00",X"0A",X"1C",X"00",X"0A",
		X"01",X"00",X"F2",X"01",X"01",X"0C",X"1C",X"FE",X"0E",X"01",X"01",X"F2",X"03",X"01",X"0C",X"0A",
		X"FE",X"0E",X"02",X"02",X"0C",X"0A",X"FE",X"0E",X"03",X"01",X"F2",X"04",X"FF",X"0B",X"08",X"02",
		X"0D",X"04",X"FE",X"0B",X"08",X"02",X"0D",X"04",X"FF",X"F2",X"02",X"FF",X"0B",X"1A",X"02",X"0D",
		X"02",X"FF",X"F1",X"01",X"00",X"0A",X"1C",X"00",X"0A",X"01",X"00",X"F2",X"01",X"00",X"0A",X"04",
		X"FF",X"0E",X"02",X"02",X"0C",X"0C",X"FE",X"0E",X"02",X"02",X"0C",X"04",X"FF",X"0A",X"01",X"00",
		X"F2",X"01",X"00",X"0A",X"03",X"01",X"0D",X"04",X"FE",X"0B",X"0A",X"02",X"0D",X"04",X"FE",X"0B",
		X"03",X"01",X"0A",X"01",X"00",X"F1",X"01",X"00",X"0A",X"1C",X"00",X"0A",X"01",X"00",X"F3",X"01",
		X"01",X"0C",X"0C",X"FE",X"0E",X"02",X"02",X"0C",X"0C",X"FE",X"0E",X"01",X"01",X"F1",X"20",X"00",
		X"FF",X"F1",X"20",X"00",X"F3",X"05",X"FF",X"0B",X"01",X"02",X"0D",X"06",X"FE",X"0B",X"02",X"02",
		X"0D",X"06",X"FE",X"0B",X"01",X"02",X"0D",X"05",X"FF",X"F1",X"02",X"00",X"0B",X"1A",X"00",X"0D",
		X"02",X"00",X"F3",X"01",X"01",X"0C",X"1C",X"FE",X"0E",X"01",X"01",X"FC",X"04",X"00",X"0A",X"16",
		X"00",X"0A",X"04",X"00",X"F3",X"03",X"FF",X"0B",X"18",X"02",X"0D",X"03",X"FF",X"F1",X"02",X"00",
		X"0C",X"1A",X"00",X"0E",X"02",X"00",X"F3",X"03",X"01",X"0C",X"05",X"FE",X"0E",X"02",X"02",X"0C",
		X"06",X"FE",X"0E",X"02",X"02",X"0C",X"05",X"FE",X"0E",X"03",X"01",X"F1",X"20",X"00",X"FF",X"F1",
		X"20",X"00",X"FB",X"0B",X"FF",X"0B",X"08",X"02",X"0D",X"0B",X"FF",X"F4",X"01",X"00",X"0A",X"1C",
		X"00",X"0A",X"01",X"00",X"FB",X"01",X"01",X"0C",X"1C",X"FE",X"0E",X"01",X"01",X"F1",X"20",X"00",
		X"FF",X"3E",X"0E",X"32",X"C7",X"40",X"32",X"D7",X"40",X"32",X"AF",X"41",X"32",X"87",X"42",X"32",
		X"97",X"42",X"32",X"2F",X"43",X"3E",X"0C",X"32",X"C8",X"40",X"32",X"D8",X"40",X"32",X"B0",X"41",
		X"32",X"88",X"42",X"32",X"98",X"42",X"32",X"30",X"43",X"3E",X"0D",X"32",X"CF",X"40",X"32",X"67",
		X"41",X"32",X"77",X"41",X"32",X"4F",X"42",X"32",X"27",X"43",X"32",X"37",X"43",X"3E",X"0B",X"32",
		X"D0",X"40",X"32",X"68",X"41",X"32",X"78",X"41",X"32",X"50",X"42",X"32",X"28",X"43",X"32",X"38",
		X"43",X"3E",X"0A",X"32",X"FB",X"41",X"32",X"1B",X"42",X"C9",X"3E",X"0E",X"32",X"AF",X"41",X"3E",
		X"0C",X"32",X"B0",X"41",X"3E",X"0D",X"32",X"4F",X"42",X"3E",X"0B",X"32",X"50",X"42",X"3E",X"0C",
		X"32",X"E1",X"42",X"3E",X"0B",X"32",X"01",X"41",X"3E",X"0D",X"32",X"1E",X"41",X"3E",X"0E",X"32",
		X"FE",X"42",X"C9",X"3E",X"0D",X"32",X"E8",X"40",X"32",X"F6",X"40",X"32",X"6F",X"42",X"3E",X"0B",
		X"32",X"E9",X"40",X"32",X"F7",X"40",X"32",X"70",X"42",X"3E",X"0E",X"32",X"8F",X"41",X"32",X"08",
		X"43",X"32",X"16",X"43",X"3E",X"0C",X"32",X"90",X"41",X"32",X"09",X"43",X"32",X"17",X"43",X"3E",
		X"0C",X"32",X"81",X"43",X"32",X"C1",X"40",X"3E",X"0B",X"32",X"21",X"43",X"32",X"61",X"40",X"3E",
		X"0E",X"32",X"9E",X"43",X"32",X"DE",X"40",X"3E",X"0D",X"32",X"3E",X"43",X"32",X"7E",X"40",X"C9",
		X"3E",X"0D",X"32",X"CA",X"40",X"32",X"D4",X"40",X"3E",X"0B",X"32",X"CB",X"40",X"32",X"D5",X"40",
		X"3E",X"0E",X"32",X"2A",X"43",X"32",X"34",X"43",X"3E",X"0C",X"32",X"2B",X"43",X"32",X"35",X"43",
		X"C9",X"3E",X"0D",X"32",X"EF",X"40",X"3E",X"0B",X"32",X"F0",X"40",X"32",X"05",X"42",X"3E",X"0C",
		X"32",X"E5",X"41",X"32",X"10",X"43",X"3E",X"0E",X"32",X"0F",X"43",X"C9",X"3E",X"40",X"CD",X"07",
		X"15",X"3E",X"01",X"CD",X"17",X"15",X"11",X"4D",X"44",X"21",X"47",X"37",X"3E",X"06",X"06",X"1C",
		X"CD",X"F5",X"15",X"11",X"C1",X"40",X"21",X"7B",X"37",X"3E",X"01",X"06",X"14",X"CD",X"DF",X"15",
		X"11",X"C2",X"40",X"21",X"8F",X"37",X"3E",X"01",X"06",X"14",X"CD",X"DF",X"15",X"11",X"C3",X"40",
		X"21",X"A3",X"37",X"3E",X"01",X"06",X"14",X"CD",X"DF",X"15",X"11",X"C4",X"40",X"21",X"8F",X"37",
		X"3E",X"01",X"06",X"14",X"CD",X"DF",X"15",X"11",X"C5",X"40",X"21",X"7B",X"37",X"3E",X"01",X"06",
		X"14",X"CD",X"DF",X"15",X"11",X"47",X"40",X"21",X"B7",X"37",X"3E",X"01",X"06",X"1C",X"CD",X"F5",
		X"15",X"11",X"49",X"40",X"21",X"B7",X"37",X"3E",X"01",X"06",X"1C",X"CD",X"F5",X"15",X"11",X"4B",
		X"40",X"21",X"B8",X"37",X"3E",X"01",X"06",X"1C",X"CD",X"F5",X"15",X"11",X"4D",X"40",X"21",X"B9",
		X"37",X"3E",X"01",X"06",X"1C",X"CD",X"DF",X"15",X"11",X"4E",X"40",X"21",X"D5",X"37",X"3E",X"01",
		X"06",X"1C",X"CD",X"DF",X"15",X"11",X"4F",X"40",X"21",X"F1",X"37",X"3E",X"01",X"06",X"1C",X"CD",
		X"DF",X"15",X"11",X"50",X"40",X"21",X"0D",X"38",X"3E",X"01",X"06",X"1C",X"CD",X"DF",X"15",X"11",
		X"51",X"40",X"21",X"29",X"38",X"3E",X"01",X"06",X"1C",X"CD",X"DF",X"15",X"11",X"52",X"40",X"21",
		X"45",X"38",X"3E",X"01",X"06",X"1C",X"CD",X"DF",X"15",X"11",X"54",X"40",X"21",X"B8",X"37",X"3E",
		X"01",X"06",X"1C",X"CD",X"F5",X"15",X"11",X"56",X"40",X"21",X"B7",X"37",X"3E",X"01",X"06",X"1C",
		X"CD",X"F5",X"15",X"11",X"58",X"40",X"21",X"B7",X"37",X"3E",X"01",X"06",X"1C",X"CD",X"F5",X"15",
		X"11",X"7A",X"40",X"21",X"61",X"38",X"3E",X"01",X"06",X"13",X"CD",X"DF",X"15",X"11",X"7B",X"40",
		X"21",X"74",X"38",X"3E",X"01",X"06",X"13",X"CD",X"DF",X"15",X"11",X"7C",X"40",X"21",X"87",X"38",
		X"3E",X"01",X"06",X"13",X"CD",X"DF",X"15",X"3E",X"0E",X"32",X"7C",X"46",X"11",X"7D",X"40",X"21",
		X"74",X"38",X"3E",X"01",X"06",X"13",X"CD",X"DF",X"15",X"11",X"7E",X"40",X"21",X"61",X"38",X"3E",
		X"01",X"06",X"13",X"CD",X"DF",X"15",X"AF",X"32",X"E6",X"4E",X"3E",X"9F",X"32",X"E7",X"4E",X"3E",
		X"A3",X"32",X"E8",X"4E",X"11",X"E7",X"4E",X"CD",X"48",X"37",X"11",X"E8",X"4E",X"CD",X"48",X"37",
		X"3E",X"01",X"CD",X"A5",X"15",X"3A",X"E6",X"4E",X"FE",X"B0",X"C8",X"3C",X"32",X"E6",X"4E",X"21",
		X"95",X"4C",X"CB",X"6E",X"C0",X"18",X"DD",X"03",X"1A",X"FE",X"A2",X"28",X"1C",X"FE",X"A6",X"28",
		X"21",X"C6",X"01",X"12",X"5F",X"D6",X"01",X"57",X"21",X"40",X"40",X"01",X"80",X"03",X"7A",X"ED",
		X"B1",X"78",X"B1",X"C8",X"2B",X"73",X"23",X"18",X"F5",X"3E",X"9F",X"12",X"5F",X"3E",X"A2",X"57",
		X"18",X"E6",X"3E",X"A3",X"12",X"5F",X"3E",X"A6",X"57",X"18",X"DD",X"A8",X"9F",X"9F",X"9F",X"9F",
		X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"A8",X"A3",
		X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",
		X"40",X"40",X"A3",X"A3",X"40",X"53",X"54",X"4E",X"45",X"53",X"45",X"52",X"50",X"40",X"5A",X"45",
		X"48",X"43",X"4E",X"41",X"53",X"40",X"A3",X"A7",X"9F",X"94",X"93",X"92",X"9E",X"93",X"9E",X"9E",
		X"93",X"9E",X"94",X"93",X"92",X"9E",X"9D",X"9E",X"93",X"9E",X"94",X"93",X"92",X"9E",X"94",X"93",
		X"92",X"9E",X"94",X"93",X"92",X"96",X"9E",X"93",X"9E",X"93",X"9E",X"94",X"93",X"9E",X"93",X"9E",
		X"93",X"9E",X"95",X"9E",X"93",X"9E",X"93",X"9E",X"93",X"9E",X"93",X"9E",X"93",X"9E",X"93",X"9E",
		X"93",X"9E",X"97",X"93",X"9E",X"93",X"9E",X"93",X"93",X"9E",X"93",X"9E",X"93",X"9E",X"93",X"95",
		X"93",X"9E",X"93",X"9E",X"93",X"9E",X"93",X"9E",X"93",X"9E",X"9E",X"9E",X"93",X"93",X"98",X"9E",
		X"9E",X"93",X"93",X"9E",X"93",X"9E",X"93",X"93",X"93",X"9E",X"99",X"96",X"93",X"9E",X"98",X"93",
		X"93",X"9E",X"93",X"9E",X"93",X"9E",X"93",X"96",X"93",X"93",X"9E",X"94",X"9E",X"93",X"96",X"9E",
		X"93",X"9E",X"93",X"9E",X"93",X"9E",X"9B",X"9E",X"93",X"9E",X"9A",X"9E",X"93",X"9E",X"93",X"9E",
		X"93",X"9E",X"93",X"9E",X"93",X"9C",X"93",X"96",X"9E",X"93",X"9E",X"9E",X"93",X"9E",X"93",X"9E",
		X"93",X"94",X"9D",X"9E",X"93",X"9E",X"9B",X"9E",X"93",X"9E",X"9C",X"93",X"96",X"9E",X"9C",X"93",
		X"96",X"A8",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",
		X"9F",X"9F",X"9F",X"A8",X"A3",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",
		X"40",X"40",X"40",X"40",X"40",X"40",X"A3",X"A3",X"40",X"52",X"41",X"54",X"53",X"48",X"43",X"45",
		X"54",X"40",X"33",X"38",X"39",X"31",X"40",X"1A",X"40",X"A3",X"C9",X"21",X"A0",X"4E",X"22",X"9D",
		X"4E",X"11",X"A1",X"4E",X"01",X"3F",X"00",X"36",X"00",X"ED",X"B0",X"C9",X"21",X"A0",X"4E",X"22",
		X"9D",X"4E",X"11",X"A1",X"4E",X"01",X"3F",X"00",X"36",X"00",X"ED",X"B0",X"C9",X"21",X"8F",X"39",
		X"22",X"35",X"4E",X"3E",X"EF",X"32",X"F8",X"4C",X"C9",X"C9",X"2A",X"35",X"4E",X"E5",X"21",X"8F",
		X"39",X"7D",X"E1",X"BD",X"CC",X"02",X"39",X"7E",X"FE",X"00",X"28",X"0E",X"23",X"46",X"3A",X"8C",
		X"4C",X"B8",X"28",X"14",X"2B",X"22",X"35",X"4E",X"18",X"17",X"23",X"46",X"3A",X"8D",X"4C",X"B8",
		X"28",X"06",X"2B",X"22",X"35",X"4E",X"18",X"09",X"23",X"7E",X"32",X"F8",X"4C",X"23",X"22",X"35",
		X"4E",X"C9",X"3E",X"FF",X"32",X"F8",X"4C",X"C9",X"C9",X"21",X"A0",X"4E",X"22",X"9D",X"4E",X"C9",
		X"C9",X"21",X"C0",X"4E",X"22",X"9D",X"4E",X"C9",X"C9",X"C9",X"C9",X"C9",X"3E",X"09",X"32",X"1C",
		X"4E",X"3E",X"02",X"32",X"1D",X"4E",X"3E",X"08",X"32",X"1E",X"4E",X"32",X"20",X"4E",X"32",X"1F",
		X"4E",X"32",X"23",X"4E",X"3E",X"16",X"32",X"21",X"4E",X"32",X"25",X"4E",X"3E",X"12",X"32",X"22",
		X"4E",X"32",X"24",X"4E",X"ED",X"5B",X"1E",X"4E",X"CD",X"80",X"39",X"ED",X"5B",X"20",X"4E",X"CD",
		X"80",X"39",X"ED",X"5B",X"22",X"4E",X"CD",X"80",X"39",X"ED",X"5B",X"24",X"4E",X"CD",X"80",X"39",
		X"3A",X"1D",X"4E",X"C6",X"02",X"32",X"1D",X"4E",X"06",X"08",X"21",X"1E",X"4E",X"35",X"23",X"10",
		X"FC",X"3E",X"05",X"CD",X"A5",X"15",X"3A",X"1C",X"4E",X"3D",X"32",X"1C",X"4E",X"20",X"C5",X"C9",
		X"CD",X"E9",X"14",X"21",X"8E",X"39",X"3A",X"1D",X"4E",X"47",X"CD",X"F5",X"15",X"C9",X"62",X"00",
		X"A4",X"FB",X"01",X"E3",X"F7",X"00",X"EC",X"FD",X"01",X"9B",X"FE",X"00",X"DC",X"FD",X"01",X"73",
		X"F7",X"00",X"EC",X"FD",X"01",X"2B",X"FE",X"00",X"A4",X"FB",X"01",X"6B",X"FE",X"00",X"64",X"FD",
		X"01",X"2B",X"FE",X"00",X"24",X"FB",X"01",X"73",X"F7",X"01",X"72",X"FF",X"01",X"4B",X"F7",X"00",
		X"94",X"FB",X"01",X"5B",X"F7",X"01",X"5C",X"FF",X"01",X"93",X"F7",X"01",X"94",X"FF",X"01",X"83",
		X"FE",X"01",X"82",X"FF",X"01",X"6B",X"FF",X"01",X"6B",X"FE",X"01",X"6A",X"FF",X"00",X"34",X"FB",
		X"00",X"33",X"FF",X"00",X"2C",X"FB",X"00",X"2D",X"FF",X"01",X"8B",X"F7",X"01",X"8C",X"FF",X"00",
		X"5C",X"FD",X"00",X"5D",X"FF",X"00",X"64",X"FD",X"00",X"63",X"FF",X"01",X"9B",X"FE",X"0B",X"20",
		X"4D",X"0B",X"3B",X"4D",X"0C",X"02",X"01",X"43",X"00",X"02",X"08",X"05",X"04",X"01",X"54",X"00",
		X"05",X"04",X"01",X"32",X"00",X"05",X"04",X"01",X"85",X"00",X"05",X"04",X"01",X"A7",X"00",X"05",
		X"04",X"01",X"64",X"00",X"05",X"04",X"01",X"0B",X"01",X"05",X"04",X"09",X"0B",X"05",X"4D",X"0B",
		X"3B",X"4D",X"01",X"F0",X"00",X"0C",X"02",X"06",X"02",X"08",X"05",X"03",X"02",X"00",X"05",X"03",
		X"07",X"0F",X"09",X"0B",X"05",X"4D",X"0C",X"04",X"01",X"A0",X"00",X"02",X"0F",X"06",X"06",X"03",
		X"10",X"00",X"05",X"01",X"07",X"07",X"06",X"03",X"EF",X"FF",X"05",X"01",X"07",X"07",X"04",X"FF",
		X"03",X"40",X"00",X"07",X"0A",X"09",X"0B",X"3B",X"4D",X"0B",X"71",X"4D",X"0B",X"8C",X"4D",X"0B",
		X"A7",X"4D",X"0C",X"02",X"01",X"80",X"00",X"02",X"0F",X"06",X"06",X"03",X"10",X"00",X"05",X"01",
		X"07",X"07",X"06",X"03",X"EF",X"FF",X"05",X"01",X"07",X"07",X"04",X"FF",X"03",X"FA",X"FF",X"07",
		X"0F",X"09",X"0C",X"02",X"01",X"40",X"00",X"02",X"0F",X"06",X"06",X"03",X"06",X"00",X"05",X"01",
		X"07",X"0F",X"04",X"FF",X"07",X"0A",X"05",X"01",X"08",X"A6",X"3A",X"0B",X"71",X"4D",X"0C",X"04",
		X"02",X"0F",X"01",X"40",X"00",X"06",X"06",X"03",X"10",X"00",X"05",X"01",X"07",X"0A",X"03",X"80",
		X"FF",X"07",X"04",X"09",X"0C",X"02",X"01",X"40",X"00",X"02",X"0F",X"06",X"06",X"03",X"06",X"00",
		X"05",X"01",X"07",X"0F",X"04",X"FF",X"07",X"0A",X"05",X"01",X"08",X"D8",X"3A",X"0B",X"A7",X"4D",
		X"0C",X"07",X"01",X"95",X"00",X"02",X"0F",X"06",X"05",X"02",X"04",X"FE",X"07",X"02",X"01",X"95",
		X"00",X"02",X"0F",X"06",X"05",X"02",X"04",X"FE",X"07",X"02",X"01",X"C7",X"00",X"02",X"0F",X"06",
		X"05",X"02",X"04",X"FE",X"07",X"02",X"01",X"95",X"00",X"02",X"0F",X"06",X"05",X"02",X"04",X"FE",
		X"07",X"02",X"01",X"C7",X"00",X"02",X"0F",X"06",X"05",X"02",X"04",X"FE",X"07",X"02",X"01",X"EC",
		X"00",X"02",X"0F",X"06",X"05",X"02",X"04",X"FE",X"07",X"02",X"01",X"C7",X"00",X"02",X"0F",X"06",
		X"05",X"02",X"04",X"FE",X"07",X"02",X"01",X"EC",X"00",X"02",X"0F",X"06",X"05",X"02",X"04",X"FE",
		X"07",X"02",X"01",X"2A",X"01",X"02",X"0F",X"06",X"05",X"02",X"04",X"FE",X"07",X"02",X"01",X"EC",
		X"00",X"02",X"0F",X"06",X"05",X"02",X"04",X"FE",X"07",X"02",X"01",X"2A",X"01",X"02",X"0F",X"06",
		X"05",X"02",X"04",X"FE",X"07",X"02",X"01",X"8E",X"01",X"02",X"0F",X"06",X"05",X"02",X"04",X"FE",
		X"07",X"02",X"01",X"2A",X"01",X"02",X"0F",X"06",X"05",X"02",X"04",X"FE",X"07",X"02",X"01",X"8E",
		X"01",X"02",X"0F",X"06",X"05",X"02",X"04",X"FE",X"07",X"02",X"01",X"D8",X"01",X"02",X"0F",X"06",
		X"05",X"02",X"04",X"FE",X"07",X"02",X"01",X"C0",X"01",X"02",X"0F",X"06",X"05",X"02",X"04",X"FE",
		X"07",X"02",X"01",X"8E",X"01",X"02",X"0F",X"06",X"05",X"02",X"04",X"FE",X"07",X"02",X"01",X"64",
		X"01",X"02",X"0F",X"06",X"05",X"02",X"04",X"FE",X"07",X"02",X"01",X"2A",X"01",X"02",X"0F",X"06",
		X"05",X"02",X"04",X"FE",X"07",X"02",X"01",X"64",X"01",X"02",X"0F",X"06",X"05",X"02",X"04",X"FE",
		X"07",X"02",X"01",X"8E",X"01",X"02",X"0F",X"06",X"05",X"02",X"04",X"FE",X"07",X"04",X"05",X"08",
		X"01",X"95",X"00",X"02",X"0F",X"06",X"05",X"02",X"04",X"FE",X"07",X"02",X"01",X"95",X"00",X"02",
		X"0F",X"06",X"05",X"02",X"04",X"FE",X"07",X"02",X"01",X"C7",X"00",X"02",X"0F",X"06",X"05",X"02",
		X"04",X"FE",X"07",X"02",X"01",X"95",X"00",X"02",X"0F",X"06",X"05",X"02",X"04",X"FE",X"07",X"02",
		X"01",X"C7",X"00",X"02",X"0F",X"06",X"05",X"02",X"04",X"FE",X"07",X"02",X"01",X"EC",X"00",X"02",
		X"0F",X"06",X"05",X"02",X"04",X"FE",X"07",X"02",X"01",X"C7",X"00",X"02",X"0F",X"06",X"05",X"02",
		X"04",X"FE",X"07",X"02",X"01",X"EC",X"00",X"02",X"0F",X"06",X"05",X"02",X"04",X"FE",X"07",X"02",
		X"01",X"2A",X"01",X"02",X"0F",X"06",X"05",X"02",X"04",X"FE",X"07",X"02",X"01",X"EC",X"00",X"02",
		X"0F",X"06",X"05",X"02",X"04",X"FE",X"07",X"02",X"01",X"2A",X"01",X"02",X"0F",X"06",X"05",X"02",
		X"04",X"FE",X"07",X"02",X"01",X"64",X"01",X"02",X"0F",X"06",X"05",X"02",X"04",X"FE",X"07",X"02",
		X"01",X"2A",X"01",X"02",X"0F",X"06",X"05",X"02",X"04",X"FE",X"07",X"02",X"01",X"64",X"01",X"02",
		X"0F",X"06",X"05",X"02",X"04",X"FE",X"07",X"02",X"01",X"64",X"01",X"02",X"0F",X"06",X"05",X"02",
		X"04",X"FE",X"07",X"06",X"05",X"0C",X"09",X"00",X"00",X"15",X"00",X"00",X"00",X"30",X"00",X"00",
		X"00",X"45",X"00",X"00",X"00",X"60",X"00",X"00",X"50",X"12",X"00",X"00",X"00",X"25",X"00",X"00",
		X"50",X"37",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"20",X"00",X"00",
		X"00",X"30",X"00",X"00",X"00",X"40",X"00",X"00",X"50",X"07",X"00",X"00",X"00",X"15",X"00",X"00",
		X"50",X"22",X"00",X"00",X"00",X"30",X"00",X"05",X"04",X"03",X"02",X"00",X"03",X"06",X"09",X"00",
		X"03",X"00",X"00",X"06",X"03",X"00",X"03",X"00",X"00",X"06",X"03",X"00",X"00",X"09",X"00",X"FF",
		X"4C",X"52",X"53",X"50",X"42",X"03",X"4D",X"43",X"53",X"60",X"17",X"03",X"4A",X"4D",X"53",X"20",
		X"85",X"02",X"42",X"4F",X"40",X"90",X"76",X"02",X"4A",X"53",X"40",X"50",X"31",X"02",X"4A",X"46",
		X"53",X"90",X"10",X"02",X"46",X"53",X"4D",X"00",X"05",X"02",X"43",X"53",X"4D",X"60",X"01",X"02",
		X"43",X"44",X"40",X"80",X"98",X"01",X"48",X"44",X"43",X"40",X"86",X"01",X"07",X"10",X"03",X"12",
		X"96",X"47",X"4F",X"52",X"4B",X"41",X"4E",X"53",X"2C",X"43",X"4F",X"50",X"59",X"52",X"49",X"47",
		X"48",X"54",X"20",X"31",X"39",X"38",X"33",X"54",X"45",X"43",X"48",X"53",X"54",X"41",X"52",X"20",
		X"49",X"4E",X"43",X"00",X"FF",X"00",X"FF",X"00",X"FB",X"00",X"E3",X"00",X"FF",X"00",X"FF",X"00",
		X"3E",X"00",X"3E",X"00",X"FF",X"00",X"FF",X"00",X"3E",X"00",X"3E",X"00",X"FF",X"00",X"FF",X"00",
		X"02",X"00",X"CB",X"00",X"FF",X"00",X"FF",X"00",X"DA",X"00",X"F3",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"3A",X"80",X"50",X"E6",X"80",X"FE",X"80",X"28",X"03",X"C3",X"FF",X"FF",X"C3",X"C7",X"02",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
