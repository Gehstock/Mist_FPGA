library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity tron_sp_bits_4 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of tron_sp_bits_4 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",
		X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"66",X"00",X"00",X"77",X"66",X"00",
		X"22",X"77",X"00",X"00",X"22",X"77",X"00",X"00",X"22",X"77",X"00",X"00",X"00",X"77",X"00",X"00",
		X"00",X"77",X"00",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",
		X"00",X"22",X"77",X"00",X"00",X"22",X"77",X"00",X"22",X"22",X"66",X"00",X"22",X"22",X"66",X"00",
		X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"77",X"22",X"77",X"00",X"77",X"22",X"77",X"00",
		X"66",X"77",X"66",X"00",X"66",X"77",X"66",X"00",X"22",X"27",X"22",X"00",X"22",X"77",X"22",X"00",
		X"00",X"77",X"77",X"22",X"00",X"22",X"77",X"22",X"00",X"22",X"66",X"00",X"00",X"22",X"66",X"00",
		X"77",X"22",X"22",X"00",X"77",X"22",X"22",X"00",X"77",X"22",X"77",X"00",X"77",X"22",X"77",X"00",
		X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",
		X"00",X"22",X"77",X"00",X"00",X"22",X"77",X"00",X"22",X"22",X"66",X"00",X"22",X"22",X"66",X"00",
		X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"77",X"22",X"77",X"00",X"77",X"22",X"77",X"00",
		X"66",X"77",X"66",X"00",X"66",X"77",X"66",X"00",X"22",X"27",X"22",X"00",X"22",X"77",X"22",X"00",
		X"00",X"77",X"77",X"22",X"00",X"22",X"77",X"22",X"00",X"22",X"66",X"00",X"00",X"22",X"66",X"00",
		X"77",X"22",X"22",X"00",X"77",X"22",X"22",X"00",X"77",X"22",X"77",X"00",X"77",X"22",X"77",X"00",
		X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"77",X"00",X"00",X"CC",X"77",X"00",X"00",X"CC",
		X"22",X"00",X"00",X"00",X"22",X"CC",X"00",X"00",X"77",X"77",X"CC",X"00",X"77",X"77",X"CC",X"00",
		X"CC",X"22",X"77",X"00",X"CC",X"22",X"77",X"00",X"CC",X"22",X"22",X"00",X"CC",X"22",X"72",X"00",
		X"77",X"77",X"22",X"00",X"77",X"72",X"22",X"00",X"77",X"77",X"22",X"00",X"77",X"77",X"22",X"00",
		X"22",X"77",X"77",X"C0",X"22",X"27",X"77",X"C0",X"22",X"22",X"77",X"00",X"22",X"22",X"77",X"00",
		X"77",X"22",X"77",X"00",X"77",X"22",X"77",X"00",X"CC",X"22",X"22",X"00",X"CC",X"22",X"22",X"00",
		X"CC",X"77",X"22",X"CC",X"CC",X"77",X"22",X"CC",X"77",X"CC",X"77",X"00",X"77",X"CC",X"77",X"00",
		X"77",X"00",X"CC",X"00",X"77",X"00",X"CC",X"00",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",
		X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",
		X"00",X"AA",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"CB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"CB",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"CB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"CB",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"A2",X"00",X"00",X"00",X"32",X"00",X"00",X"10",X"33",X"00",X"10",X"11",X"33",X"00",X"11",
		X"31",X"31",X"01",X"D1",X"33",X"32",X"01",X"D1",X"33",X"31",X"01",X"D1",X"33",X"31",X"11",X"D1",
		X"33",X"31",X"D1",X"D1",X"33",X"32",X"D1",X"D1",X"33",X"31",X"D1",X"D1",X"33",X"31",X"D1",X"D1",
		X"33",X"31",X"D1",X"D1",X"33",X"32",X"D1",X"D1",X"33",X"31",X"D1",X"D1",X"33",X"3A",X"D1",X"D1",
		X"33",X"31",X"21",X"D1",X"33",X"32",X"22",X"D1",X"33",X"22",X"32",X"D1",X"33",X"23",X"33",X"D1",
		X"33",X"23",X"33",X"D1",X"33",X"22",X"32",X"D1",X"33",X"32",X"22",X"D1",X"33",X"31",X"21",X"D1",
		X"33",X"1A",X"D1",X"D1",X"33",X"AD",X"D1",X"D1",X"33",X"11",X"11",X"D1",X"31",X"00",X"01",X"D1",
		X"11",X"00",X"00",X"11",X"10",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"11",X"11",X"00",X"DD",X"DD",X"DD",X"00",X"33",X"33",X"33",X"10",X"11",X"11",X"11",X"11",
		X"2A",X"22",X"22",X"11",X"11",X"11",X"11",X"10",X"33",X"33",X"33",X"00",X"33",X"33",X"33",X"00",
		X"11",X"11",X"21",X"00",X"01",X"DD",X"22",X"00",X"01",X"D2",X"D2",X"00",X"01",X"D2",X"D3",X"00",
		X"01",X"D2",X"33",X"00",X"01",X"D2",X"D3",X"00",X"01",X"D2",X"D2",X"00",X"0A",X"DD",X"22",X"00",
		X"11",X"1A",X"21",X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",X"00",X"1A",X"1A",X"11",X"00",
		X"01",X"DD",X"DD",X"00",X"01",X"DD",X"DD",X"00",X"01",X"DD",X"DD",X"00",X"11",X"11",X"11",X"00",
		X"33",X"33",X"33",X"00",X"33",X"33",X"33",X"00",X"11",X"11",X"11",X"10",X"2A",X"22",X"22",X"11",
		X"11",X"11",X"11",X"11",X"33",X"33",X"33",X"10",X"DD",X"DD",X"DD",X"00",X"11",X"11",X"11",X"00",
		X"50",X"00",X"00",X"00",X"50",X"00",X"00",X"50",X"55",X"00",X"00",X"55",X"C5",X"00",X"00",X"2C",
		X"C5",X"00",X"05",X"CC",X"6C",X"00",X"05",X"2C",X"AC",X"20",X"05",X"55",X"6C",X"C5",X"05",X"55",
		X"6C",X"C7",X"05",X"2C",X"6C",X"7C",X"25",X"CC",X"6C",X"C7",X"25",X"2C",X"AC",X"C7",X"25",X"55",
		X"6C",X"7C",X"25",X"55",X"6C",X"77",X"25",X"2C",X"6C",X"55",X"CC",X"CC",X"6C",X"55",X"7C",X"2C",
		X"AC",X"55",X"7C",X"55",X"6C",X"55",X"7C",X"55",X"6C",X"55",X"7C",X"2C",X"6C",X"55",X"7C",X"CC",
		X"6C",X"55",X"7C",X"2C",X"AC",X"55",X"7C",X"55",X"6C",X"55",X"7C",X"55",X"6C",X"55",X"CC",X"2C",
		X"6C",X"77",X"75",X"CC",X"6C",X"CC",X"55",X"2C",X"CC",X"22",X"05",X"55",X"CC",X"22",X"05",X"55",
		X"C5",X"77",X"00",X"50",X"55",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"50",X"00",X"00",X"05",
		X"25",X"2C",X"55",X"00",X"25",X"2C",X"55",X"00",X"55",X"CC",X"5C",X"50",X"5A",X"55",X"A5",X"55",
		X"CC",X"C6",X"CC",X"65",X"CC",X"CC",X"CC",X"C5",X"6A",X"66",X"A6",X"55",X"CC",X"CC",X"CC",X"50",
		X"55",X"5C",X"CC",X"00",X"00",X"5C",X"77",X"00",X"00",X"C7",X"77",X"00",X"00",X"77",X"57",X"77",
		X"00",X"77",X"55",X"C0",X"00",X"75",X"55",X"00",X"00",X"75",X"55",X"00",X"00",X"75",X"55",X"00",
		X"00",X"75",X"55",X"00",X"00",X"75",X"55",X"00",X"00",X"75",X"55",X"00",X"00",X"77",X"55",X"C0",
		X"00",X"77",X"57",X"77",X"00",X"C7",X"77",X"00",X"00",X"5C",X"77",X"00",X"55",X"5C",X"CC",X"00",
		X"CC",X"CC",X"CC",X"50",X"6A",X"66",X"A6",X"55",X"CC",X"CC",X"CC",X"C5",X"CC",X"C6",X"CC",X"65",
		X"55",X"55",X"A5",X"55",X"55",X"CC",X"5C",X"50",X"25",X"2C",X"55",X"00",X"C5",X"CC",X"55",X"C5",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"00",X"00",X"00",X"33",X"00",X"00",X"0F",X"30",X"00",X"00",X"F3",X"30",X"00",
		X"00",X"33",X"3F",X"00",X"55",X"33",X"3F",X"00",X"05",X"35",X"99",X"00",X"00",X"55",X"99",X"00",
		X"00",X"AA",X"99",X"00",X"00",X"AA",X"3F",X"00",X"00",X"9A",X"93",X"00",X"0F",X"99",X"59",X"00",
		X"F5",X"55",X"55",X"00",X"0F",X"33",X"93",X"00",X"00",X"39",X"33",X"00",X"00",X"99",X"3F",X"00",
		X"00",X"99",X"55",X"00",X"00",X"55",X"55",X"00",X"09",X"95",X"55",X"00",X"99",X"39",X"95",X"00",
		X"00",X"33",X"FF",X"00",X"00",X"F3",X"00",X"00",X"00",X"0F",X"A0",X"00",X"00",X"00",X"A0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"22",X"50",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"32",X"00",X"00",
		X"00",X"32",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"23",X"00",X"00",X"00",X"32",X"00",X"00",
		X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",
		X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E2",X"22",X"20",X"22",X"22",X"00",X"00",
		X"22",X"BB",X"00",X"00",X"22",X"EB",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"00",
		X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",
		X"00",X"32",X"00",X"00",X"00",X"23",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",
		X"32",X"30",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",
		X"02",X"00",X"00",X"00",X"02",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",
		X"00",X"2E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EB",X"00",X"00",X"00",X"77",X"00",X"00",
		X"00",X"EB",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"2E",X"00",X"00",X"00",X"22",X"00",X"00",
		X"00",X"22",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",
		X"00",X"00",X"22",X"00",X"00",X"00",X"23",X"00",X"00",X"00",X"32",X"00",X"00",X"20",X"22",X"00",
		X"00",X"20",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"20",X"00",X"00",X"00",X"A2",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"A0",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"22",X"02",X"00",X"00",X"20",X"22",X"00",X"00",X"00",X"32",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"D6",X"EE",X"00",X"00",X"26",X"BE",X"00",X"00",
		X"26",X"BE",X"00",X"00",X"27",X"BE",X"00",X"00",X"77",X"BE",X"00",X"00",X"7D",X"BE",X"00",X"00",
		X"7D",X"BE",X"00",X"00",X"DD",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"23",X"30",X"00",X"00",X"22",X"22",X"00",X"00",X"02",X"22",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"7C",X"00",
		X"00",X"00",X"7C",X"00",X"00",X"00",X"7C",X"00",X"00",X"00",X"7C",X"00",X"00",X"00",X"0C",X"00",
		X"00",X"00",X"07",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"07",X"00",
		X"00",X"00",X"07",X"00",X"00",X"00",X"7F",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"C7",X"00",X"00",X"00",X"C7",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"70",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"70",X"00",
		X"00",X"00",X"70",X"00",X"00",X"00",X"F7",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"C7",X"00",X"00",X"00",X"C7",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"07",X"00",X"00",
		X"00",X"07",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"C7",X"00",X"00",X"00",X"C7",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C7",X"00",X"00",
		X"00",X"C7",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"7C",X"00",X"00",X"00",X"7C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"C7",X"00",X"00",X"00",X"C7",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"70",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"C7",X"00",X"00",
		X"00",X"07",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"C7",X"00",X"00",X"00",X"C7",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"C7",X"00",X"00",X"00",X"C7",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"C7",X"00",X"00",X"00",X"C7",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C7",X"00",X"00",X"00",
		X"C7",X"00",X"00",X"00",X"C7",X"00",X"00",X"00",X"00",X"F7",X"F7",X"00",X"00",X"FF",X"CC",X"00",
		X"00",X"FF",X"77",X"00",X"00",X"7F",X"CC",X"00",X"00",X"00",X"C7",X"00",X"00",X"00",X"C7",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"7F",X"00",X"C7",X"00",X"FF",X"00",
		X"C7",X"F7",X"CC",X"00",X"00",X"FF",X"77",X"00",X"00",X"7F",X"CC",X"00",X"00",X"00",X"C7",X"00",
		X"00",X"00",X"C7",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"77",X"00",X"70",X"FF",X"CC",X"00",X"CC",X"FF",X"77",X"00",
		X"CC",X"FF",X"77",X"00",X"70",X"FF",X"CC",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"33",X"33",X"00",X"03",X"99",X"E9",X"00",X"03",X"99",X"E9",X"33",
		X"39",X"9E",X"EE",X"99",X"99",X"99",X"EE",X"EE",X"49",X"99",X"9E",X"99",X"C4",X"99",X"99",X"99",
		X"C4",X"99",X"EE",X"33",X"49",X"9E",X"EE",X"EE",X"33",X"99",X"99",X"99",X"03",X"33",X"99",X"33",
		X"00",X"00",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"93",X"00",X"00",X"00",
		X"E9",X"30",X"00",X"00",X"9E",X"93",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"E9",X"00",X"00",
		X"33",X"9E",X"00",X"00",X"EE",X"39",X"00",X"00",X"99",X"93",X"00",X"00",X"33",X"39",X"00",X"00",
		X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"00",X"00",X"00",X"39",X"03",X"33",X"33",X"9E",X"03",X"99",X"E9",X"EE",X"03",X"99",X"E9",X"99",
		X"39",X"9E",X"EE",X"99",X"99",X"99",X"EE",X"93",X"49",X"99",X"9E",X"30",X"C4",X"99",X"99",X"00",
		X"C4",X"99",X"EE",X"00",X"49",X"9E",X"EE",X"30",X"33",X"99",X"9E",X"93",X"03",X"33",X"99",X"99",
		X"00",X"00",X"39",X"EE",X"00",X"00",X"03",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"9E",X"30",X"00",X"00",
		X"E9",X"30",X"00",X"00",X"99",X"30",X"00",X"00",X"93",X"00",X"00",X"00",X"30",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",
		X"99",X"30",X"00",X"00",X"33",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"E0",X"00",
		X"00",X"EE",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"E0",X"00",X"00",X"99",X"E9",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"99",X"00",
		X"00",X"9E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9E",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E9",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"9E",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"4E",X"00",X"00",
		X"00",X"04",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"04",X"00",X"00",
		X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"9E",X"00",
		X"00",X"00",X"9E",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"9E",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"9E",X"00",
		X"00",X"00",X"9E",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"40",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",
		X"00",X"00",X"0E",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",
		X"00",X"E9",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",
		X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"E9",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"9E",X"00",X"00",X"99",X"EE",X"00",X"00",X"EE",X"CC",X"9E",X"00",
		X"EE",X"EE",X"CC",X"00",X"CC",X"CC",X"C1",X"00",X"EE",X"CC",X"11",X"99",X"EE",X"CC",X"11",X"99",
		X"EE",X"CC",X"11",X"99",X"EE",X"CC",X"11",X"99",X"CC",X"CC",X"C1",X"00",X"EE",X"EE",X"CC",X"00",
		X"EE",X"CC",X"9E",X"00",X"99",X"EE",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"CC",X"00",X"00",
		X"00",X"99",X"90",X"00",X"00",X"9E",X"90",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"90",X"00",
		X"00",X"CC",X"F0",X"00",X"00",X"CC",X"90",X"00",X"00",X"CC",X"90",X"00",X"00",X"CC",X"E0",X"00",
		X"00",X"CC",X"E0",X"00",X"00",X"CC",X"E0",X"00",X"00",X"CC",X"E0",X"00",X"00",X"CC",X"00",X"00",
		X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"47",X"00",X"00",X"FF",X"77",X"00",X"00",X"77",X"CC",X"47",X"00",
		X"77",X"77",X"CC",X"00",X"CC",X"CC",X"C4",X"00",X"4C",X"CC",X"44",X"44",X"4C",X"CC",X"44",X"44",
		X"4C",X"CC",X"44",X"44",X"4C",X"CC",X"44",X"44",X"CC",X"CC",X"C4",X"00",X"77",X"77",X"CC",X"00",
		X"77",X"CC",X"47",X"00",X"FF",X"77",X"00",X"00",X"00",X"47",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",
		X"00",X"FF",X"F0",X"00",X"00",X"F4",X"F0",X"00",X"00",X"44",X"00",X"00",X"00",X"CC",X"00",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"F0",X"00",
		X"00",X"CC",X"F0",X"00",X"00",X"CC",X"40",X"00",X"00",X"CC",X"40",X"00",X"00",X"CC",X"70",X"00",
		X"00",X"CC",X"70",X"00",X"00",X"CC",X"70",X"00",X"00",X"CC",X"70",X"00",X"00",X"CC",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",
		X"31",X"31",X"31",X"00",X"13",X"13",X"13",X"00",X"31",X"31",X"31",X"00",X"11",X"11",X"11",X"00",
		X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",
		X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",
		X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",
		X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"53",X"53",X"53",X"05",X"35",X"35",X"35",X"03",X"53",X"53",X"53",X"05",X"35",X"35",X"35",
		X"33",X"53",X"53",X"50",X"33",X"33",X"33",X"30",X"33",X"33",X"33",X"30",X"33",X"33",X"33",X"30",
		X"33",X"33",X"33",X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",X"00",
		X"33",X"33",X"33",X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",X"00",
		X"33",X"33",X"33",X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",X"00",
		X"13",X"13",X"13",X"00",X"31",X"31",X"31",X"00",X"13",X"13",X"13",X"00",X"31",X"31",X"31",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"05",X"B5",X"B5",X"B5",X"0B",X"5B",X"5B",X"5B",X"05",X"B5",X"B5",X"B5",X"0B",X"5B",X"5B",X"5B",
		X"05",X"B5",X"B5",X"B5",X"0B",X"5B",X"5B",X"5B",X"05",X"55",X"55",X"55",X"05",X"55",X"55",X"55",
		X"55",X"55",X"55",X"50",X"55",X"55",X"55",X"50",X"55",X"55",X"55",X"50",X"55",X"55",X"55",X"50",
		X"55",X"55",X"55",X"50",X"55",X"55",X"55",X"50",X"55",X"55",X"55",X"50",X"55",X"55",X"55",X"50",
		X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",
		X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",
		X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"35",X"35",X"35",X"00",
		X"53",X"53",X"53",X"00",X"35",X"35",X"35",X"00",X"53",X"53",X"53",X"00",X"35",X"35",X"35",X"00",
		X"DB",X"DB",X"DB",X"00",X"BD",X"BD",X"BD",X"00",X"DB",X"DB",X"DB",X"00",X"BD",X"BD",X"BD",X"00",
		X"DB",X"DB",X"DB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",
		X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",
		X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",
		X"BB",X"BB",X"BB",X"B0",X"BB",X"BB",X"BB",X"B0",X"BB",X"BB",X"BB",X"B0",X"BB",X"BB",X"BB",X"B0",
		X"BB",X"BB",X"BB",X"B0",X"BB",X"BB",X"BB",X"B0",X"BB",X"BB",X"BB",X"B0",X"BB",X"BB",X"BB",X"B0",
		X"0B",X"BB",X"BB",X"BB",X"0B",X"BB",X"BB",X"BB",X"05",X"B5",X"B5",X"B5",X"0B",X"5B",X"5B",X"5B",
		X"05",X"B5",X"B5",X"B5",X"0B",X"5B",X"5B",X"5B",X"05",X"B5",X"B5",X"B5",X"0B",X"5B",X"5B",X"5B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DF",X"DF",X"DF",X"00",X"FD",X"FD",X"FD",X"00",X"DF",X"DF",X"DF",X"00",X"FD",X"FD",X"FD",X"00",
		X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",
		X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",
		X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",
		X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",X"BD",X"BD",X"BD",X"00",
		X"DB",X"DB",X"DB",X"D0",X"BD",X"BD",X"BD",X"B0",X"DB",X"DB",X"DB",X"D0",X"BD",X"BD",X"BD",X"B0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",
		X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",
		X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",
		X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",
		X"FF",X"FF",X"FF",X"00",X"DF",X"DF",X"DF",X"00",X"FD",X"FD",X"FD",X"00",X"DF",X"DF",X"DF",X"D0",
		X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"66",X"65",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"05",X"05",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"44",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"44",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"06",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"65",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"05",X"05",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"05",X"00",X"0E",X"00",X"05",X"00",X"E0",X"0A",X"00",X"7F",X"09",X"00",X"00",X"F0",X"20",
		X"0A",X"0F",X"0F",X"0B",X"00",X"00",X"00",X"A0",X"AB",X"00",X"0B",X"00",X"F0",X"F0",X"F0",X"00",
		X"0A",X"09",X"09",X"00",X"90",X"20",X"90",X"00",X"0E",X"0B",X"00",X"B0",X"00",X"00",X"00",X"A5",
		X"0E",X"00",X"0B",X"00",X"0A",X"00",X"2E",X"A0",X"00",X"0B",X"00",X"00",X"00",X"09",X"00",X"A7",
		X"00",X"90",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"E0",X"00",X"00",X"00",X"95",X"00",X"00",X"7E",X"09",X"00",X"00",X"90",X"05",X"00",X"00",
		X"09",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",
		X"07",X"00",X"00",X"00",X"20",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2A",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"07",X"00",X"07",X"00",
		X"07",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"44",X"44",X"00",X"40",X"44",X"40",X"00",X"44",
		X"44",X"00",X"00",X"44",X"44",X"00",X"00",X"40",X"44",X"00",X"00",X"00",X"07",X"00",X"00",X"00",
		X"07",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"77",X"00",X"55",X"00",X"55",X"00",
		X"CC",X"00",X"5C",X"00",X"CC",X"00",X"05",X"00",X"C5",X"00",X"00",X"00",X"50",X"00",X"00",X"00",
		X"50",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"50",X"00",X"00",X"00",
		X"50",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"50",X"55",X"00",X"00",X"00",X"CC",X"00",X"00",
		X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"50",X"50",X"00",X"00",X"50",X"50",X"50",X"00",
		X"50",X"00",X"C5",X"00",X"55",X"50",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"57",X"00",X"00",X"00",X"05",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"75",X"55",X"55",X"00",X"75",X"CC",X"5C",X"00",
		X"75",X"CC",X"5C",X"00",X"75",X"CC",X"5C",X"00",X"75",X"55",X"55",X"00",X"75",X"00",X"00",X"00",
		X"75",X"00",X"00",X"00",X"75",X"00",X"05",X"00",X"75",X"00",X"5C",X"00",X"00",X"00",X"5C",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"50",X"00",X"00",X"00",X"75",
		X"00",X"00",X"00",X"75",X"00",X"00",X"55",X"50",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"5C",X"00",X"75",X"00",X"5C",X"00",X"75",X"00",X"05",X"00",X"75",X"00",X"00",X"00",
		X"75",X"00",X"00",X"00",X"75",X"55",X"55",X"00",X"75",X"CC",X"5C",X"00",X"75",X"CC",X"5C",X"00",
		X"75",X"CC",X"5C",X"00",X"75",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
