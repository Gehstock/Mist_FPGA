library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity draw_bg_bits_2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of draw_bg_bits_2 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"00",X"3C",X"00",X"00",
		X"00",X"00",X"03",X"00",X"0C",X"C0",X"30",X"30",X"FF",X"FC",X"C0",X"0C",X"C0",X"0C",X"00",X"00",
		X"00",X"00",X"FF",X"F0",X"C0",X"0C",X"FF",X"F0",X"C0",X"0C",X"C0",X"0C",X"FF",X"F0",X"00",X"00",
		X"00",X"00",X"FF",X"FC",X"C0",X"0C",X"C0",X"00",X"C0",X"00",X"C0",X"0C",X"FF",X"FC",X"00",X"00",
		X"00",X"00",X"FF",X"F0",X"C0",X"0C",X"C0",X"0C",X"C0",X"0C",X"C0",X"0C",X"FF",X"F0",X"00",X"00",
		X"00",X"00",X"FF",X"F0",X"C0",X"00",X"FF",X"C0",X"C0",X"00",X"C0",X"00",X"FF",X"FC",X"00",X"00",
		X"00",X"00",X"FF",X"FC",X"C0",X"00",X"FF",X"C0",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FC",X"C0",X"00",X"C3",X"FC",X"C0",X"0C",X"C0",X"0C",X"3F",X"F0",X"00",X"00",
		X"00",X"00",X"C0",X"0C",X"C0",X"0C",X"C0",X"0C",X"FF",X"FC",X"C0",X"0C",X"C0",X"0C",X"00",X"00",
		X"00",X"00",X"FF",X"FC",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"FF",X"FC",X"00",X"00",
		X"00",X"00",X"00",X"FC",X"00",X"30",X"00",X"30",X"C0",X"30",X"C0",X"30",X"FF",X"F0",X"00",X"00",
		X"00",X"00",X"C0",X"0C",X"C0",X"30",X"FF",X"C0",X"C0",X"30",X"C0",X"0C",X"C0",X"0C",X"00",X"00",
		X"00",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"0C",X"C0",X"0C",X"FF",X"FC",X"00",X"00",
		X"00",X"00",X"C0",X"0C",X"F0",X"3C",X"CC",X"CC",X"C3",X"0C",X"C0",X"0C",X"C0",X"0C",X"00",X"00",
		X"00",X"00",X"F0",X"0C",X"CC",X"0C",X"C3",X"0C",X"C0",X"CC",X"C0",X"3C",X"C0",X"0C",X"00",X"00",
		X"00",X"00",X"3F",X"F0",X"C0",X"0C",X"C0",X"0C",X"C0",X"0C",X"C0",X"0C",X"3F",X"F0",X"00",X"00",
		X"00",X"00",X"FF",X"F0",X"C0",X"0C",X"C0",X"0C",X"FF",X"F0",X"C0",X"00",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"F0",X"C0",X"0C",X"C0",X"0C",X"FF",X"F0",X"C0",X"0C",X"C0",X"0C",X"00",X"00",
		X"00",X"00",X"FF",X"FC",X"C0",X"00",X"FF",X"FC",X"00",X"0C",X"C0",X"0C",X"FF",X"FC",X"00",X"00",
		X"00",X"00",X"FF",X"FC",X"C3",X"0C",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"0C",X"C0",X"0C",X"C0",X"0C",X"C0",X"0C",X"C0",X"0C",X"3F",X"F0",X"00",X"00",
		X"00",X"00",X"C0",X"0C",X"30",X"30",X"30",X"30",X"0C",X"C0",X"0C",X"C0",X"03",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"0C",X"C3",X"0C",X"C3",X"0C",X"CC",X"CC",X"CC",X"CC",X"30",X"30",X"00",X"00",
		X"00",X"00",X"F0",X"3C",X"3C",X"F0",X"0F",X"C0",X"3C",X"F0",X"F0",X"3C",X"C0",X"0C",X"00",X"00",
		X"00",X"00",X"C0",X"0C",X"30",X"30",X"0C",X"C0",X"03",X"00",X"03",X"00",X"03",X"00",X"00",X"00",
		X"00",X"C0",X"3F",X"FC",X"30",X"C0",X"3F",X"FC",X"00",X"CC",X"00",X"CC",X"3F",X"FC",X"00",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"03",X"33",X"0C",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"CC",X"CC",X"33",X"33",X"CC",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"C0",X"CC",X"C0",X"33",X"30",X"CC",X"CC",
		X"33",X"33",X"CC",X"CC",X"33",X"33",X"CC",X"CC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"33",X"33",X"CC",X"CC",X"33",X"33",X"CC",X"CC",
		X"33",X"33",X"0C",X"CC",X"03",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"CC",X"CC",X"33",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"30",X"CC",X"C0",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"F0",X"FF",X"C0",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"03",X"FF",X"0F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"FF",X"C0",X"FF",X"F0",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",
		X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",
		X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",
		X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"0F",X"FF",X"03",X"FF",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"F1",X"FF",X"C5",X"00",X"15",
		X"00",X"00",X"03",X"FF",X"0F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"FF",X"C0",X"FF",X"F0",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",
		X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",
		X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",
		X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",X"0F",X"FF",X"03",X"FF",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"F0",X"FF",X"C0",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",
		X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",
		X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"F1",X"FF",X"C5",X"00",X"14",
		X"55",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"50",X"00",X"50",X"00",X"50",X"00",
		X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"00",
		X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"00",X"40",X"00",
		X"00",X"00",X"00",X"30",X"00",X"F0",X"00",X"30",X"00",X"30",X"00",X"30",X"00",X"FC",X"00",X"00",
		X"00",X"00",X"FF",X"FC",X"00",X"0C",X"3F",X"FC",X"C0",X"00",X"C0",X"0C",X"FF",X"FC",X"00",X"00",
		X"00",X"00",X"FF",X"FC",X"C0",X"0C",X"03",X"F0",X"00",X"0C",X"C0",X"0C",X"FF",X"FC",X"00",X"00",
		X"00",X"00",X"00",X"30",X"C0",X"30",X"C0",X"30",X"FF",X"FC",X"00",X"30",X"00",X"30",X"00",X"00",
		X"00",X"00",X"FF",X"FC",X"C0",X"00",X"FF",X"FC",X"00",X"0C",X"C0",X"0C",X"3F",X"F0",X"00",X"00",
		X"00",X"00",X"3F",X"FC",X"C0",X"00",X"FF",X"F0",X"C0",X"0C",X"C0",X"0C",X"3F",X"F0",X"00",X"00",
		X"00",X"00",X"FF",X"FC",X"C0",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"00",
		X"00",X"00",X"3F",X"F0",X"C0",X"0C",X"3F",X"F0",X"C0",X"0C",X"C0",X"0C",X"3F",X"F0",X"00",X"00",
		X"00",X"00",X"3F",X"F0",X"C0",X"0C",X"3F",X"FC",X"00",X"0C",X"C0",X"0C",X"3F",X"F0",X"00",X"00",
		X"00",X"00",X"3F",X"F0",X"C0",X"0C",X"C0",X"0C",X"C0",X"0C",X"C0",X"0C",X"3F",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"AA",X"00",X"80",X"00",X"80",X"00",X"00",
		X"00",X"00",X"08",X"AA",X"08",X"80",X"08",X"AA",X"A8",X"80",X"08",X"80",X"08",X"AA",X"00",X"00",
		X"00",X"00",X"A0",X"80",X"00",X"80",X"80",X"80",X"00",X"80",X"00",X"80",X"A8",X"AA",X"00",X"00",
		X"00",X"00",X"00",X"AA",X"00",X"80",X"00",X"80",X"00",X"80",X"08",X"80",X"A8",X"AA",X"00",X"00",
		X"00",X"00",X"A0",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"A0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"AA",X"00",X"80",X"00",X"80",X"00",X"00",
		X"00",X"00",X"08",X"AA",X"08",X"80",X"08",X"AA",X"A8",X"80",X"08",X"80",X"08",X"AA",X"00",X"00",
		X"00",X"00",X"A0",X"80",X"00",X"80",X"80",X"80",X"00",X"80",X"00",X"80",X"A8",X"AA",X"00",X"00",
		X"00",X"00",X"00",X"AA",X"00",X"80",X"00",X"80",X"00",X"80",X"08",X"80",X"A8",X"AA",X"00",X"00",
		X"00",X"00",X"A0",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"A0",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"33",X"30",X"CC",X"CC",X"33",X"30",X"CC",X"CC",X"33",X"30",X"CC",X"C1",X"33",X"05",X"00",X"15",
		X"55",X"55",X"55",X"54",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"55",X"00",X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"50",X"00",X"54",X"00",X"54",X"00",
		X"54",X"00",X"54",X"00",X"54",X"00",X"54",X"00",X"54",X"00",X"54",X"00",X"54",X"00",X"54",X"00",
		X"54",X"00",X"54",X"00",X"54",X"00",X"54",X"00",X"54",X"00",X"54",X"00",X"54",X"00",X"50",X"00",
		X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"54",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"55",X"00",X"15",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"50",X"00",X"54",X"00",X"55",X"00",
		X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",
		X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",
		X"55",X"00",X"54",X"00",X"50",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"55",X"00",X"15",X"00",X"05",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"54",X"00",X"55",X"00",
		X"55",X"40",X"55",X"40",X"55",X"40",X"55",X"40",X"55",X"40",X"55",X"40",X"55",X"40",X"55",X"40",
		X"55",X"40",X"55",X"40",X"55",X"00",X"54",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"04",X"40",X"10",X"10",X"55",X"54",X"40",X"04",X"40",X"04",X"00",X"00",
		X"00",X"00",X"55",X"50",X"40",X"04",X"55",X"50",X"40",X"04",X"40",X"04",X"55",X"50",X"00",X"00",
		X"00",X"00",X"55",X"54",X"40",X"04",X"40",X"00",X"40",X"00",X"40",X"04",X"55",X"54",X"00",X"00",
		X"00",X"00",X"55",X"50",X"40",X"04",X"40",X"04",X"40",X"04",X"40",X"04",X"55",X"50",X"00",X"00",
		X"00",X"00",X"55",X"50",X"40",X"00",X"55",X"40",X"40",X"00",X"40",X"00",X"55",X"54",X"00",X"00",
		X"00",X"00",X"55",X"50",X"40",X"00",X"55",X"40",X"40",X"00",X"40",X"00",X"40",X"00",X"00",X"00",
		X"00",X"00",X"55",X"54",X"40",X"00",X"40",X"54",X"40",X"04",X"40",X"04",X"15",X"50",X"00",X"00",
		X"00",X"00",X"40",X"04",X"40",X"04",X"40",X"04",X"55",X"54",X"40",X"04",X"40",X"04",X"00",X"00",
		X"00",X"00",X"55",X"54",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"55",X"54",X"00",X"00",
		X"00",X"00",X"05",X"54",X"00",X"10",X"00",X"10",X"40",X"10",X"40",X"10",X"15",X"40",X"00",X"00",
		X"00",X"00",X"40",X"04",X"40",X"10",X"55",X"40",X"40",X"10",X"40",X"04",X"40",X"04",X"00",X"00",
		X"00",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"55",X"54",X"00",X"00",
		X"00",X"00",X"40",X"04",X"50",X"14",X"44",X"44",X"41",X"04",X"40",X"04",X"40",X"04",X"00",X"00",
		X"00",X"00",X"50",X"04",X"44",X"04",X"41",X"04",X"40",X"44",X"40",X"14",X"40",X"04",X"00",X"00",
		X"00",X"00",X"15",X"50",X"40",X"04",X"40",X"04",X"40",X"04",X"40",X"04",X"15",X"50",X"00",X"00",
		X"00",X"00",X"55",X"50",X"40",X"04",X"40",X"04",X"55",X"50",X"40",X"00",X"40",X"00",X"00",X"00",
		X"00",X"00",X"55",X"50",X"40",X"04",X"40",X"04",X"55",X"50",X"40",X"10",X"40",X"04",X"00",X"00",
		X"00",X"00",X"55",X"54",X"40",X"00",X"55",X"54",X"00",X"04",X"40",X"04",X"55",X"54",X"00",X"00",
		X"00",X"00",X"55",X"54",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"40",X"04",X"40",X"04",X"40",X"04",X"40",X"04",X"40",X"04",X"15",X"50",X"00",X"00",
		X"00",X"00",X"40",X"04",X"10",X"10",X"10",X"10",X"04",X"40",X"04",X"40",X"01",X"00",X"00",X"00",
		X"00",X"00",X"40",X"04",X"41",X"04",X"41",X"04",X"41",X"04",X"44",X"44",X"10",X"10",X"00",X"00",
		X"00",X"00",X"40",X"04",X"10",X"10",X"04",X"40",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"50",X"14",X"14",X"50",X"05",X"40",X"14",X"50",X"50",X"14",X"40",X"04",X"00",X"00",
		X"00",X"00",X"15",X"50",X"40",X"04",X"40",X"04",X"40",X"04",X"40",X"04",X"15",X"50",X"00",X"00",
		X"00",X"00",X"00",X"10",X"00",X"50",X"00",X"10",X"00",X"10",X"00",X"10",X"00",X"54",X"00",X"00",
		X"00",X"00",X"55",X"54",X"00",X"04",X"15",X"54",X"40",X"00",X"40",X"04",X"55",X"54",X"00",X"00",
		X"00",X"00",X"55",X"54",X"40",X"04",X"01",X"50",X"00",X"04",X"40",X"04",X"55",X"54",X"00",X"00",
		X"00",X"00",X"00",X"10",X"40",X"10",X"40",X"10",X"55",X"54",X"00",X"10",X"00",X"10",X"00",X"00",
		X"00",X"00",X"55",X"54",X"40",X"00",X"55",X"54",X"00",X"04",X"40",X"04",X"15",X"50",X"00",X"00",
		X"00",X"00",X"15",X"54",X"40",X"00",X"55",X"50",X"40",X"04",X"40",X"04",X"15",X"50",X"00",X"00",
		X"00",X"00",X"55",X"54",X"40",X"04",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"00",
		X"00",X"00",X"15",X"50",X"40",X"04",X"15",X"50",X"40",X"04",X"40",X"04",X"15",X"50",X"00",X"00",
		X"00",X"00",X"15",X"50",X"40",X"04",X"15",X"54",X"00",X"04",X"40",X"04",X"15",X"50",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"14",X"00",X"14",X"00",X"00",
		X"01",X"00",X"15",X"54",X"11",X"00",X"15",X"54",X"01",X"04",X"01",X"04",X"15",X"54",X"01",X"00",
		X"AA",X"80",X"AA",X"A0",X"A0",X"A8",X"A0",X"28",X"A0",X"28",X"A0",X"28",X"A0",X"28",X"A0",X"28",
		X"A0",X"28",X"A0",X"28",X"A0",X"28",X"A0",X"28",X"A0",X"28",X"A0",X"A8",X"AA",X"A0",X"AA",X"80",
		X"AA",X"A8",X"AA",X"A8",X"A0",X"28",X"A0",X"28",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"AA",X"A0",
		X"AA",X"A0",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"28",X"A0",X"28",X"AA",X"A8",X"AA",X"A8",
		X"0A",X"80",X"2A",X"A0",X"28",X"A0",X"A0",X"28",X"A0",X"28",X"A0",X"28",X"A0",X"28",X"AA",X"A8",
		X"AA",X"A8",X"A0",X"28",X"A0",X"28",X"A0",X"28",X"A0",X"28",X"A0",X"28",X"A0",X"28",X"A0",X"28",
		X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",
		X"AA",X"80",X"AA",X"A0",X"A0",X"A8",X"A0",X"28",X"A0",X"28",X"A0",X"28",X"A0",X"28",X"AA",X"A0",
		X"A0",X"0A",X"A0",X"0A",X"A0",X"0A",X"A0",X"0A",X"A2",X"8A",X"A2",X"8A",X"A2",X"8A",X"A2",X"8A",
		X"A2",X"8A",X"A2",X"8A",X"AA",X"AA",X"AA",X"AA",X"A8",X"2A",X"A8",X"2A",X"A0",X"0A",X"A0",X"0A",
		X"AA",X"A8",X"AA",X"A8",X"A0",X"28",X"A0",X"28",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"AA",X"A8",
		X"AA",X"A8",X"00",X"28",X"00",X"28",X"00",X"28",X"A0",X"28",X"A0",X"28",X"AA",X"A8",X"AA",X"A8",
		X"AA",X"AA",X"AA",X"AA",X"82",X"82",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",
		X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",
		X"A0",X"28",X"A0",X"28",X"A0",X"28",X"A8",X"28",X"A8",X"28",X"A8",X"28",X"AA",X"28",X"A2",X"28",
		X"A2",X"28",X"A2",X"A8",X"A0",X"A8",X"A0",X"A8",X"A0",X"A8",X"A0",X"28",X"A0",X"28",X"A0",X"28",
		X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"28",X"A0",X"28",X"AA",X"A8",X"AA",X"A8",
		X"0A",X"80",X"2A",X"A0",X"A8",X"A8",X"A0",X"28",X"A0",X"00",X"A8",X"00",X"2A",X"00",X"0A",X"80",
		X"02",X"A0",X"00",X"A8",X"00",X"28",X"A0",X"28",X"A0",X"28",X"A8",X"A8",X"2A",X"A0",X"0A",X"80",
		X"AA",X"AA",X"AA",X"AA",X"82",X"82",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",
		X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",
		X"A0",X"28",X"A0",X"28",X"A0",X"28",X"A8",X"28",X"A8",X"28",X"A8",X"28",X"AA",X"28",X"A2",X"28",
		X"A2",X"28",X"A2",X"A8",X"A0",X"A8",X"A0",X"A8",X"A0",X"A8",X"A0",X"28",X"A0",X"28",X"A0",X"28",
		X"0A",X"80",X"0A",X"80",X"28",X"A0",X"A0",X"28",X"A0",X"28",X"A0",X"28",X"A0",X"28",X"AA",X"A8",
		X"AA",X"A8",X"A0",X"28",X"A0",X"28",X"A0",X"28",X"A0",X"28",X"A0",X"28",X"A0",X"28",X"A0",X"28",
		X"AA",X"00",X"AA",X"80",X"A0",X"A0",X"A0",X"28",X"A0",X"28",X"A0",X"28",X"A0",X"28",X"A0",X"28",
		X"A0",X"28",X"A0",X"28",X"A0",X"28",X"A0",X"28",X"A0",X"28",X"A0",X"A8",X"AA",X"A0",X"AA",X"80",
		X"00",X"15",X"00",X"15",X"00",X"05",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"54",X"00",X"55",X"00",
		X"55",X"40",X"55",X"50",X"55",X"50",X"55",X"50",X"55",X"50",X"55",X"50",X"55",X"50",X"55",X"50",
		X"55",X"50",X"55",X"50",X"55",X"50",X"55",X"50",X"55",X"50",X"55",X"50",X"55",X"50",X"55",X"50",
		X"55",X"50",X"55",X"50",X"55",X"50",X"55",X"40",X"55",X"00",X"54",X"00",X"00",X"00",X"00",X"00",
		X"00",X"A0",X"02",X"A0",X"0A",X"A0",X"0A",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",
		X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",
		X"0A",X"80",X"2A",X"A0",X"A8",X"A8",X"A0",X"28",X"00",X"28",X"00",X"28",X"00",X"28",X"00",X"A0",
		X"02",X"A0",X"0A",X"80",X"2A",X"00",X"A8",X"00",X"A0",X"00",X"A0",X"28",X"AA",X"A8",X"AA",X"A8",
		X"0A",X"80",X"2A",X"A0",X"A8",X"A8",X"A0",X"28",X"00",X"28",X"00",X"28",X"00",X"A8",X"0A",X"A0",
		X"0A",X"A0",X"00",X"A8",X"00",X"28",X"00",X"28",X"A0",X"28",X"A8",X"A8",X"2A",X"A0",X"0A",X"80",
		X"00",X"A0",X"00",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",
		X"AA",X"A8",X"AA",X"A8",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",
		X"AA",X"A8",X"AA",X"A8",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A2",X"80",X"AA",X"A0",
		X"A8",X"A8",X"A0",X"28",X"00",X"28",X"00",X"28",X"A0",X"28",X"A8",X"A8",X"2A",X"A0",X"0A",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"FC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"FC",X"FC",X"00",X"00",X"FF",X"FC",
		X"FC",X"FC",X"0C",X"C0",X"FC",X"FC",X"C0",X"0C",X"C0",X"0C",X"FC",X"FC",X"00",X"00",X"FF",X"FC",
		X"FC",X"FC",X"C0",X"CC",X"FC",X"CC",X"0C",X"CC",X"0C",X"CC",X"FC",X"FC",X"00",X"00",X"FF",X"FC",
		X"FC",X"FC",X"0C",X"C0",X"0C",X"FC",X"0C",X"0C",X"0C",X"0C",X"0C",X"FC",X"00",X"00",X"FF",X"FC",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"15",X"55",X"00",X"00",X"00",X"00",
		X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"54",X"54",X"44",X"44",X"44",X"44",X"44",X"44",X"54",X"54",X"00",X"00",X"55",X"54",X"00",X"00",
		X"FF",X"C0",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",
		X"F0",X"3C",X"F0",X"3C",X"F0",X"3C",X"F0",X"3C",X"F0",X"3C",X"F0",X"3C",X"FC",X"FC",X"3C",X"F0",
		X"0F",X"C0",X"0F",X"C0",X"0F",X"C0",X"0F",X"C0",X"0F",X"C0",X"0F",X"C0",X"0F",X"C0",X"0F",X"C0",
		X"15",X"54",X"17",X"D7",X"17",X"17",X"17",X"17",X"15",X"5F",X"17",X"17",X"17",X"17",X"17",X"17",
		X"14",X"14",X"17",X"17",X"17",X"17",X"17",X"17",X"17",X"17",X"17",X"17",X"17",X"17",X"17",X"17",
		X"15",X"54",X"17",X"D7",X"17",X"3F",X"17",X"03",X"15",X"57",X"0F",X"D7",X"17",X"17",X"17",X"17",
		X"15",X"54",X"1D",X"74",X"1D",X"74",X"01",X"70",X"01",X"70",X"01",X"70",X"01",X"70",X"01",X"70",
		X"17",X"17",X"17",X"17",X"15",X"57",X"3F",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"70",X"01",X"70",X"01",X"70",X"03",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"17",X"17",X"17",X"17",X"15",X"57",X"3F",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"FF",X"0F",X"AE",X"3F",X"FF",X"3A",X"AF",X"3F",X"FF",X"3F",X"FF",X"3F",X"FF",
		X"FC",X"00",X"F0",X"CC",X"C3",X"33",X"0C",X"CC",X"33",X"33",X"0C",X"CC",X"33",X"33",X"0C",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"54",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FC",X"FC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"FC",X"FC",X"00",X"00",X"FF",X"FC",
		X"00",X"00",X"FC",X"FC",X"0C",X"C0",X"FC",X"FC",X"C0",X"0C",X"FC",X"FC",X"00",X"00",X"FF",X"FC",
		X"00",X"00",X"FC",X"FC",X"C0",X"CC",X"FC",X"CC",X"0C",X"CC",X"FC",X"FC",X"00",X"00",X"FF",X"FC",
		X"0A",X"80",X"2A",X"A0",X"A8",X"A8",X"A0",X"28",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",
		X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"28",X"A8",X"A8",X"2A",X"A0",X"0A",X"80",
		X"0A",X"80",X"2A",X"A0",X"A8",X"A8",X"A0",X"28",X"A0",X"28",X"A0",X"28",X"A0",X"28",X"A0",X"28",
		X"A0",X"28",X"A0",X"28",X"A0",X"28",X"A0",X"28",X"A0",X"28",X"A8",X"A8",X"2A",X"A0",X"0A",X"80",
		X"2A",X"A8",X"2A",X"A8",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",
		X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"2A",X"A8",X"2A",X"A8",
		X"AA",X"80",X"AA",X"A0",X"A0",X"A8",X"A0",X"28",X"A0",X"28",X"A0",X"28",X"A0",X"A8",X"AA",X"A0",
		X"AA",X"A0",X"A0",X"A8",X"A0",X"28",X"A0",X"28",X"A0",X"28",X"A0",X"A8",X"AA",X"A0",X"AA",X"80",
		X"AA",X"A8",X"AA",X"A8",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"AA",X"A0",
		X"AA",X"A0",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"AA",X"A8",X"AA",X"A8",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"F0",X"30",X"0C",X"C3",X"C3",X"CC",X"03",X"CC",X"03",X"C3",X"C3",X"30",X"0C",X"0F",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"FF",X"03",X"FF",X"03",X"C0",X"03",X"C0",X"03",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"03",X"C0",X"03",X"C0",X"03",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"C0",X"FF",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",
		X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",
		X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"FF",X"03",X"FF",X"03",X"C0",X"03",X"C0",X"03",X"C0",
		X"03",X"C0",X"03",X"C0",X"03",X"C0",X"FF",X"FF",X"FF",X"FF",X"03",X"C0",X"03",X"C0",X"03",X"C0",
		X"03",X"C0",X"03",X"C0",X"03",X"C0",X"FF",X"C0",X"FF",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",
		X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"FF",X"03",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"C0",X"03",X"C0",X"03",X"C0",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"C0",X"03",X"C0",X"03",X"C0",X"FF",X"C0",X"FF",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FC",X"FC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"FC",X"FC",X"00",X"00",X"FF",X"FC",
		X"00",X"00",X"FC",X"FC",X"0C",X"C0",X"FC",X"FC",X"C0",X"0C",X"FC",X"FC",X"00",X"00",X"FF",X"FC",
		X"00",X"00",X"FC",X"FC",X"C0",X"CC",X"FC",X"CC",X"0C",X"CC",X"FC",X"FC",X"00",X"00",X"FF",X"FC",
		X"00",X"00",X"FC",X"FC",X"0C",X"C0",X"0C",X"FC",X"0C",X"0C",X"0C",X"FC",X"00",X"00",X"FF",X"FC",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
