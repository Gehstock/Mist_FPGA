library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity obj2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of obj2 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"31",X"31",X"10",X"00",X"00",X"00",X"02",X"00",X"88",X"EE",X"FF",X"E6",X"E6",X"50",X"00",
		X"00",X"00",X"00",X"66",X"FF",X"CC",X"E0",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"13",X"11",X"00",X"00",X"01",X"12",X"12",X"99",X"DD",X"C9",X"6A",X"6A",X"79",X"E0",X"80",
		X"B8",X"9E",X"2C",X"C0",X"F0",X"60",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"33",X"F7",X"70",X"00",X"00",X"00",X"00",X"00",X"AA",X"FF",X"D4",X"40",
		X"00",X"00",X"00",X"77",X"EE",X"E8",X"F0",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"C0",
		X"01",X"33",X"01",X"00",X"00",X"01",X"01",X"12",X"00",X"EE",X"EE",X"FC",X"3D",X"E2",X"C0",X"00",
		X"CF",X"CF",X"3C",X"F0",X"88",X"00",X"00",X"00",X"08",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"32",X"00",X"00",X"00",X"00",X"00",X"11",X"FE",X"CC",
		X"00",X"00",X"00",X"00",X"44",X"F8",X"F0",X"01",X"00",X"00",X"00",X"00",X"30",X"C0",X"80",X"08",
		X"60",X"81",X"11",X"11",X"00",X"00",X"01",X"00",X"00",X"44",X"FF",X"5E",X"12",X"24",X"08",X"00",
		X"CD",X"CF",X"36",X"C4",X"88",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"77",X"00",X"00",X"00",X"11",X"33",X"FE",X"CC",X"CC",
		X"00",X"00",X"88",X"88",X"F0",X"F0",X"03",X"47",X"00",X"00",X"40",X"80",X"00",X"00",X"00",X"C0",
		X"FC",X"C0",X"00",X"01",X"11",X"00",X"00",X"00",X"00",X"22",X"77",X"FF",X"2B",X"01",X"03",X"12",
		X"DE",X"B8",X"E2",X"E2",X"E2",X"C0",X"80",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"70",X"00",X"00",X"60",X"E0",X"70",X"A9",X"C5",X"D1",
		X"00",X"10",X"10",X"24",X"3C",X"38",X"B8",X"98",X"80",X"00",X"00",X"00",X"00",X"44",X"66",X"EE",
		X"E1",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"2C",X"7F",X"77",X"26",X"23",X"00",X"00",X"00",
		X"31",X"22",X"73",X"33",X"31",X"10",X"10",X"00",X"CC",X"44",X"88",X"CC",X"CC",X"CC",X"CC",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"61",X"61",X"42",X"DB",
		X"20",X"20",X"40",X"48",X"68",X"38",X"30",X"B9",X"00",X"00",X"00",X"44",X"44",X"CC",X"CC",X"88",
		X"00",X"11",X"32",X"30",X"43",X"04",X"00",X"00",X"C8",X"F3",X"F7",X"7F",X"13",X"11",X"00",X"00",
		X"B9",X"11",X"77",X"33",X"39",X"31",X"31",X"10",X"00",X"88",X"00",X"88",X"88",X"88",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"54",X"61",X"43",X"53",
		X"80",X"80",X"80",X"80",X"D1",X"F1",X"71",X"B9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"57",X"CC",X"F9",X"F9",X"F3",X"C1",X"08",X"08",
		X"B9",X"11",X"31",X"B8",X"98",X"9C",X"88",X"00",X"00",X"88",X"88",X"88",X"88",X"88",X"80",X"08",
		X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"00",X"20",X"20",X"10",X"10",X"12",X"86",X"97",X"D3",
		X"00",X"00",X"11",X"91",X"F3",X"F3",X"31",X"B9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"53",X"C8",X"61",X"D3",X"D3",X"C2",X"42",X"04",
		X"11",X"10",X"CC",X"CC",X"4E",X"44",X"00",X"00",X"88",X"CC",X"EE",X"E6",X"71",X"10",X"00",X"00",
		X"10",X"00",X"00",X"00",X"00",X"20",X"60",X"70",X"00",X"80",X"80",X"42",X"C3",X"C1",X"C0",X"A2",
		X"00",X"00",X"66",X"77",X"EE",X"5D",X"3B",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"EE",
		X"30",X"20",X"11",X"32",X"30",X"30",X"30",X"01",X"F3",X"40",X"DB",X"B7",X"95",X"08",X"08",X"00",
		X"71",X"10",X"88",X"CE",X"4C",X"00",X"00",X"00",X"F7",X"70",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"20",X"10",X"00",X"00",X"00",X"30",X"00",X"00",X"11",X"11",X"F0",X"F0",X"0C",X"2E",
		X"00",X"00",X"00",X"88",X"CC",X"F7",X"33",X"33",X"00",X"00",X"00",X"00",X"00",X"88",X"CC",X"EE",
		X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B7",X"D1",X"74",X"74",X"74",X"30",X"10",X"00",
		X"00",X"44",X"EE",X"FF",X"4D",X"08",X"0C",X"84",X"F3",X"30",X"00",X"08",X"88",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"30",X"10",X"01",X"00",X"00",X"00",X"00",X"22",X"F1",X"F0",X"08",
		X"00",X"00",X"00",X"00",X"00",X"88",X"F7",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C4",
		X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"3B",X"3F",X"C6",X"32",X"11",X"00",X"00",X"00",
		X"00",X"22",X"FF",X"A7",X"84",X"42",X"01",X"00",X"60",X"18",X"88",X"88",X"00",X"00",X"08",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"30",X"00",X"00",X"00",X"EE",X"77",X"71",X"F0",X"80",
		X"00",X"00",X"00",X"00",X"55",X"FF",X"B2",X"20",X"00",X"00",X"00",X"00",X"CC",X"FE",X"E0",X"00",
		X"01",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"3F",X"3F",X"C3",X"F0",X"11",X"00",X"00",X"00",
		X"00",X"77",X"77",X"F3",X"CB",X"74",X"30",X"00",X"08",X"CC",X"08",X"00",X"00",X"08",X"08",X"84",
		X"00",X"00",X"00",X"F7",X"73",X"30",X"00",X"02",X"00",X"00",X"00",X"88",X"EE",X"F7",X"50",X"00",
		X"00",X"00",X"00",X"00",X"FB",X"EE",X"E0",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"13",X"11",X"03",X"34",X"F0",X"00",X"00",X"99",X"DD",X"8D",X"7B",X"E2",X"88",X"00",X"00",
		X"B8",X"9E",X"2C",X"E2",X"F9",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"73",X"78",X"00",X"02",X"00",X"00",X"00",X"00",X"CC",X"F7",X"D0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"66",X"E0",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"13",X"11",X"78",X"34",X"00",X"00",X"00",X"99",X"DD",X"C1",X"F3",X"CC",X"00",X"00",X"00",
		X"B8",X"9E",X"2C",X"60",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"81",X"00",X"0A",X"42",X"E1",
		X"00",X"50",X"01",X"16",X"81",X"DA",X"22",X"F7",X"00",X"C0",X"3C",X"C3",X"0A",X"49",X"52",X"EE",
		X"0F",X"01",X"00",X"00",X"00",X"40",X"00",X"00",X"0F",X"0F",X"01",X"00",X"14",X"02",X"40",X"00",
		X"77",X"D7",X"25",X"4E",X"90",X"C2",X"12",X"04",X"CE",X"AB",X"4E",X"81",X"06",X"68",X"4D",X"07",
		X"00",X"00",X"40",X"00",X"00",X"40",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"A0",X"08",X"00",X"00",X"08",X"28",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"77",X"00",X"00",X"01",X"F0",X"80",X"00",X"30",X"F9",
		X"00",X"00",X"F0",X"00",X"12",X"60",X"C0",X"F8",X"00",X"00",X"E0",X"00",X"C0",X"00",X"00",X"80",
		X"00",X"77",X"33",X"00",X"00",X"01",X"00",X"00",X"1E",X"9F",X"8B",X"66",X"80",X"3C",X"01",X"00",
		X"E0",X"AD",X"0C",X"24",X"03",X"00",X"0F",X"00",X"00",X"80",X"00",X"00",X"48",X"00",X"2C",X"00",
		X"00",X"00",X"00",X"12",X"10",X"00",X"00",X"33",X"00",X"12",X"60",X"C0",X"00",X"30",X"F9",X"BC",
		X"70",X"C0",X"30",X"04",X"08",X"F0",X"E8",X"E1",X"80",X"00",X"80",X"00",X"00",X"80",X"00",X"80",
		X"44",X"33",X"77",X"00",X"00",X"00",X"00",X"00",X"1F",X"8F",X"BB",X"22",X"40",X"0F",X"00",X"00",
		X"8C",X"0C",X"01",X"01",X"81",X"0F",X"00",X"00",X"00",X"00",X"2C",X"10",X"0E",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"30",X"24",X"02",X"00",X"10",X"70",X"48",X"80",X"01",X"30",X"73",X"34",
		X"80",X"60",X"C0",X"80",X"20",X"C0",X"E1",X"C2",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",
		X"11",X"77",X"00",X"33",X"00",X"00",X"00",X"00",X"9F",X"0F",X"89",X"FF",X"20",X"01",X"02",X"00",
		X"8F",X"0F",X"00",X"00",X"0F",X"0A",X"00",X"00",X"24",X"0C",X"12",X"0C",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"10",X"20",X"34",X"30",X"60",X"D0",X"90",X"90",X"10",X"30",X"71",
		X"80",X"60",X"80",X"20",X"60",X"D0",X"F8",X"E4",X"00",X"00",X"00",X"00",X"00",X"82",X"02",X"05",
		X"00",X"00",X"11",X"33",X"00",X"00",X"00",X"00",X"70",X"34",X"8F",X"00",X"EE",X"88",X"00",X"00",
		X"E9",X"48",X"08",X"01",X"83",X"0C",X"08",X"00",X"0D",X"03",X"06",X"0C",X"00",X"00",X"00",X"00",
		X"00",X"10",X"10",X"30",X"20",X"20",X"20",X"24",X"C0",X"B0",X"60",X"40",X"60",X"30",X"71",X"72",
		X"00",X"00",X"00",X"80",X"A0",X"E0",X"C0",X"F8",X"00",X"00",X"00",X"00",X"00",X"50",X"D0",X"A0",
		X"06",X"00",X"11",X"33",X"11",X"00",X"00",X"00",X"70",X"07",X"8F",X"88",X"00",X"66",X"00",X"00",
		X"C8",X"80",X"10",X"30",X"24",X"06",X"00",X"00",X"60",X"40",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"10",X"10",X"20",X"20",X"20",X"02",X"40",X"24",X"00",X"00",X"40",X"90",X"D0",X"50",X"70",X"72",
		X"00",X"00",X"00",X"40",X"40",X"C0",X"F0",X"CA",X"00",X"00",X"00",X"B0",X"A0",X"A0",X"A0",X"40",
		X"20",X"60",X"24",X"04",X"00",X"00",X"00",X"00",X"72",X"16",X"07",X"02",X"DD",X"BB",X"AA",X"00",
		X"C8",X"C0",X"80",X"10",X"9A",X"89",X"00",X"00",X"40",X"40",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"00",X"00",X"80",X"90",X"90",X"58",X"70",X"31",
		X"00",X"00",X"00",X"40",X"40",X"D0",X"E1",X"E4",X"00",X"20",X"A0",X"A0",X"A0",X"A0",X"20",X"20",
		X"12",X"10",X"10",X"10",X"01",X"00",X"00",X"00",X"13",X"03",X"01",X"80",X"22",X"22",X"11",X"00",
		X"E4",X"E0",X"48",X"08",X"44",X"44",X"44",X"00",X"60",X"40",X"40",X"48",X"40",X"00",X"00",X"00",
		X"00",X"00",X"00",X"A0",X"A0",X"82",X"49",X"40",X"00",X"00",X"00",X"50",X"50",X"70",X"70",X"7A",
		X"10",X"20",X"20",X"20",X"30",X"24",X"C0",X"C8",X"00",X"80",X"80",X"80",X"48",X"40",X"40",X"48",
		X"40",X"24",X"12",X"10",X"10",X"01",X"00",X"00",X"36",X"16",X"03",X"00",X"A2",X"00",X"00",X"00",
		X"C8",X"C0",X"C0",X"80",X"44",X"44",X"88",X"00",X"40",X"40",X"48",X"40",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"40",X"24",X"1A",X"00",X"00",X"00",X"20",X"A0",X"38",X"70",X"70",
		X"20",X"82",X"58",X"41",X"C0",X"C0",X"C0",X"C8",X"00",X"00",X"00",X"80",X"80",X"C0",X"80",X"C0",
		X"0C",X"04",X"24",X"12",X"00",X"00",X"00",X"00",X"B6",X"27",X"03",X"44",X"19",X"68",X"04",X"00",
		X"E8",X"C0",X"C0",X"62",X"00",X"88",X"44",X"00",X"40",X"28",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"05",X"04",X"28",X"01",X"24",X"01",X"40",X"60",X"B0",X"F1",X"36",
		X"C0",X"24",X"92",X"90",X"81",X"80",X"C0",X"E8",X"00",X"00",X"00",X"00",X"80",X"08",X"40",X"68",
		X"0B",X"0C",X"06",X"12",X"00",X"00",X"00",X"00",X"1F",X"03",X"23",X"91",X"1C",X"12",X"01",X"00",
		X"E0",X"E0",X"3D",X"00",X"44",X"11",X"00",X"00",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"24",X"10",X"24",X"12",X"10",X"D0",X"70",X"79",
		X"00",X"80",X"68",X"30",X"12",X"01",X"80",X"C8",X"00",X"00",X"00",X"00",X"00",X"C0",X"48",X"00",
		X"04",X"06",X"0B",X"0C",X"07",X"01",X"00",X"00",X"36",X"1F",X"0B",X"11",X"00",X"0F",X"01",X"00",
		X"E0",X"F1",X"68",X"00",X"AA",X"19",X"08",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"00",
		X"10",X"01",X"00",X"01",X"00",X"00",X"10",X"00",X"00",X"E0",X"01",X"E0",X"20",X"12",X"78",X"71",
		X"00",X"00",X"E0",X"02",X"01",X"00",X"C0",X"F9",X"00",X"00",X"00",X"00",X"C0",X"08",X"00",X"00",
		X"01",X"00",X"02",X"01",X"0C",X"03",X"00",X"00",X"1E",X"13",X"0F",X"08",X"00",X"0D",X"03",X"00",
		X"F1",X"F8",X"68",X"CC",X"44",X"0E",X"07",X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"77",X"00",X"00",X"78",X"C0",X"80",X"00",X"30",X"F9",
		X"00",X"00",X"F0",X"00",X"12",X"60",X"C0",X"F8",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"80",
		X"00",X"77",X"33",X"00",X"00",X"01",X"00",X"00",X"1E",X"9F",X"8B",X"66",X"80",X"3C",X"01",X"00",
		X"E0",X"AD",X"0C",X"04",X"1E",X"00",X"0F",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"2C",X"00",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"77",X"00",X"00",X"01",X"F0",X"80",X"00",X"30",X"F9",
		X"00",X"00",X"F0",X"00",X"78",X"40",X"C0",X"F8",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"80",
		X"00",X"77",X"33",X"00",X"00",X"00",X"01",X"00",X"1E",X"9F",X"8B",X"66",X"80",X"C0",X"0F",X"00",
		X"E0",X"AD",X"0C",X"24",X"03",X"00",X"1E",X"00",X"00",X"80",X"00",X"00",X"48",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"20",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"20",
		X"00",X"00",X"00",X"20",X"10",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"00",X"00",X"00",X"10",X"0F",X"01",X"84",X"00",X"0D",X"1E",X"0E",X"0E",X"C3",X"3D",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"0B",X"00",X"00",X"00",X"40",X"00",X"00",X"1C",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"80",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"68",
		X"2D",X"1C",X"62",X"75",X"FC",X"FE",X"FF",X"FF",X"0F",X"87",X"E9",X"FF",X"EF",X"8F",X"CE",X"07",
		X"10",X"20",X"6C",X"CE",X"8C",X"8C",X"18",X"28",X"2C",X"24",X"02",X"00",X"00",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"60",X"24",
		X"00",X"00",X"00",X"30",X"E0",X"00",X"CC",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"71",X"24",X"23",X"11",X"00",X"00",X"00",
		X"00",X"33",X"CC",X"00",X"0E",X"CF",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"20",X"31",X"60",
		X"00",X"40",X"C0",X"80",X"00",X"FF",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"00",X"24",X"00",X"30",X"01",X"00",X"00",X"00",X"00",
		X"11",X"EE",X"80",X"CF",X"33",X"00",X"00",X"00",X"00",X"00",X"0E",X"3F",X"CC",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"60",X"40",X"73",X"62",
		X"00",X"00",X"00",X"00",X"00",X"88",X"22",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"60",X"04",X"10",X"00",X"00",X"88",X"00",
		X"22",X"CC",X"C3",X"3B",X"00",X"00",X"00",X"00",X"1F",X"6E",X"88",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"44",X"46",X"47",X"23",X"23",X"00",X"00",X"00",X"00",X"22",X"22",X"44",X"44",
		X"00",X"00",X"00",X"00",X"88",X"98",X"54",X"54",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",
		X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2A",X"E8",X"24",X"00",X"00",X"00",X"11",X"00",
		X"20",X"C0",X"48",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"11",X"44",X"44",
		X"00",X"00",X"20",X"20",X"60",X"20",X"EC",X"64",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"8F",X"67",X"11",X"00",X"00",X"00",X"00",X"00",X"44",X"33",X"3C",X"CD",X"00",X"00",X"00",X"00",
		X"20",X"60",X"02",X"80",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"20",X"30",X"10",X"00",X"FF",X"00",X"88",
		X"00",X"00",X"00",X"00",X"80",X"40",X"C8",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"07",X"CF",X"33",X"00",X"00",X"00",X"88",X"77",X"10",X"3F",X"CC",X"00",X"00",X"00",
		X"42",X"00",X"C0",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"70",X"00",X"33",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"80",X"60",X"42",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"CC",X"33",X"00",X"07",X"3F",X"CC",X"00",
		X"00",X"E8",X"42",X"4C",X"88",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"70",X"70",X"00",X"EE",X"00",
		X"00",X"00",X"08",X"0C",X"D2",X"E0",X"C0",X"84",X"00",X"00",X"00",X"00",X"00",X"88",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"EE",X"00",X"70",X"61",X"03",X"00",
		X"00",X"C0",X"84",X"0E",X"1E",X"59",X"C4",X"00",X"44",X"00",X"00",X"00",X"88",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"12",X"00",X"88",X"54",X"10",
		X"00",X"00",X"87",X"F0",X"70",X"C0",X"80",X"08",X"00",X"00",X"6A",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"32",X"54",X"88",X"00",X"03",X"00",X"00",
		X"00",X"80",X"08",X"C0",X"34",X"1E",X"0F",X"00",X"88",X"00",X"00",X"00",X"00",X"C4",X"6A",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"70",X"70",X"00",X"EE",X"00",
		X"00",X"00",X"08",X"0C",X"D2",X"E0",X"C0",X"84",X"00",X"00",X"00",X"00",X"00",X"88",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"EE",X"00",X"70",X"61",X"03",X"00",
		X"00",X"C0",X"84",X"0E",X"1E",X"59",X"C4",X"00",X"44",X"00",X"00",X"00",X"88",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"70",X"00",X"33",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"80",X"60",X"42",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"CC",X"33",X"00",X"07",X"3F",X"CC",X"00",
		X"00",X"E8",X"42",X"4C",X"88",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"50",X"70",X"00",X"EE",X"00",
		X"00",X"00",X"08",X"0C",X"D2",X"E0",X"C0",X"84",X"00",X"00",X"00",X"00",X"00",X"88",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"EE",X"00",X"70",X"61",X"03",X"00",
		X"00",X"C0",X"84",X"0E",X"1E",X"59",X"C4",X"00",X"44",X"00",X"00",X"00",X"88",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"52",X"B8",X"10",X"01",
		X"00",X"00",X"0E",X"78",X"F0",X"80",X"B3",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"00",
		X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"01",X"03",X"CB",X"54",X"11",X"00",
		X"00",X"C4",X"B3",X"08",X"78",X"3C",X"86",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"12",
		X"00",X"00",X"00",X"10",X"70",X"80",X"66",X"11",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"88",
		X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"12",X"11",X"00",X"00",X"00",X"00",
		X"00",X"99",X"66",X"08",X"8F",X"67",X"11",X"00",X"00",X"88",X"00",X"00",X"00",X"08",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"80",X"00",
		X"03",X"00",X"B4",X"08",X"02",X"00",X"10",X"00",X"07",X"0B",X"1A",X"04",X"03",X"07",X"09",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"20",X"40",X"00",X"10",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"DB",X"7C",X"D3",X"BC",X"0F",X"87",X"B4",X"DA",X"96",X"A5",X"4B",X"0E",X"3C",X"C3",X"1E",
		X"84",X"8C",X"8A",X"09",X"87",X"40",X"48",X"84",X"00",X"40",X"00",X"00",X"08",X"60",X"00",X"00",
		X"49",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"69",X"0F",X"24",X"60",X"20",X"20",X"80",X"00",
		X"28",X"10",X"00",X"40",X"00",X"20",X"00",X"00",X"20",X"10",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"20",X"00",X"88",X"89",X"00",X"20",X"70",X"3C",X"5E",X"16",X"DE",X"CE",
		X"00",X"00",X"10",X"70",X"F0",X"F0",X"71",X"F7",X"00",X"00",X"E0",X"C0",X"80",X"00",X"00",X"CC",
		X"77",X"89",X"88",X"00",X"20",X"00",X"00",X"00",X"FF",X"EC",X"FC",X"16",X"1E",X"5E",X"16",X"02",
		X"FF",X"7F",X"17",X"87",X"87",X"07",X"01",X"00",X"F8",X"CC",X"00",X"00",X"08",X"0C",X"0E",X"00",
		X"00",X"00",X"00",X"00",X"01",X"41",X"00",X"11",X"00",X"80",X"E0",X"2C",X"BC",X"3C",X"FC",X"EC",
		X"00",X"30",X"F0",X"F0",X"E0",X"F3",X"F7",X"F7",X"C0",X"80",X"00",X"00",X"00",X"00",X"E8",X"CC",
		X"89",X"BB",X"45",X"44",X"44",X"10",X"00",X"00",X"FF",X"EE",X"FE",X"DE",X"07",X"27",X"03",X"00",
		X"FF",X"07",X"C3",X"C3",X"C3",X"C0",X"08",X"08",X"88",X"00",X"0C",X"0E",X"0F",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"30",X"03",X"03",X"40",X"00",X"00",X"10",X"90",X"F0",X"78",X"AC",X"2C",
		X"60",X"E0",X"C0",X"C0",X"E2",X"F3",X"F7",X"F7",X"00",X"00",X"00",X"00",X"A8",X"C0",X"CC",X"88",
		X"11",X"01",X"99",X"77",X"22",X"22",X"00",X"00",X"FD",X"FF",X"FE",X"6F",X"01",X"13",X"41",X"00",
		X"EF",X"03",X"C3",X"E1",X"68",X"2C",X"2C",X"20",X"88",X"0F",X"0F",X"0E",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"70",X"34",X"16",X"17",X"10",X"30",X"70",X"70",X"70",X"F0",X"F0",X"D0",
		X"80",X"00",X"00",X"33",X"FF",X"F7",X"FF",X"DF",X"00",X"00",X"40",X"80",X"88",X"88",X"00",X"01",
		X"01",X"91",X"01",X"00",X"99",X"66",X"22",X"11",X"D9",X"EE",X"FE",X"FF",X"27",X"00",X"00",X"20",
		X"0F",X"07",X"E1",X"E0",X"78",X"7C",X"1E",X"00",X"0F",X"0E",X"0C",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"30",X"34",X"07",X"60",X"E0",X"E0",X"F0",X"F1",X"F0",X"D0",X"E0",
		X"00",X"10",X"20",X"64",X"EE",X"EE",X"EF",X"CF",X"00",X"00",X"00",X"00",X"00",X"01",X"0F",X"0F",
		X"03",X"02",X"40",X"00",X"00",X"22",X"11",X"00",X"BD",X"7D",X"FF",X"7F",X"57",X"CC",X"44",X"22",
		X"89",X"F8",X"3C",X"9E",X"9F",X"07",X"40",X"00",X"0E",X"0C",X"80",X"C0",X"C0",X"08",X"00",X"00",
		X"10",X"10",X"10",X"10",X"10",X"10",X"00",X"70",X"80",X"80",X"C0",X"C0",X"F1",X"F1",X"D1",X"E0",
		X"40",X"40",X"EA",X"EE",X"EE",X"EF",X"CF",X"8F",X"00",X"00",X"00",X"01",X"07",X"0E",X"0E",X"0C",
		X"07",X"13",X"03",X"00",X"20",X"00",X"00",X"00",X"F1",X"7D",X"77",X"77",X"27",X"22",X"EE",X"11",
		X"30",X"F0",X"8F",X"DF",X"03",X"00",X"20",X"88",X"80",X"C0",X"C0",X"68",X"00",X"00",X"00",X"00",
		X"00",X"02",X"03",X"03",X"03",X"01",X"01",X"00",X"00",X"00",X"11",X"19",X"3F",X"1F",X"1F",X"C1",
		X"80",X"80",X"C4",X"CC",X"FE",X"FC",X"FC",X"D8",X"00",X"20",X"60",X"E0",X"E0",X"C0",X"C0",X"80",
		X"30",X"07",X"13",X"01",X"00",X"00",X"00",X"00",X"E0",X"3C",X"3F",X"3B",X"01",X"80",X"00",X"33",
		X"B8",X"8F",X"EF",X"EE",X"8C",X"88",X"88",X"66",X"E0",X"78",X"AC",X"0C",X"00",X"80",X"00",X"00",
		X"00",X"00",X"08",X"0C",X"07",X"07",X"03",X"03",X"20",X"20",X"31",X"33",X"77",X"7F",X"3F",X"1D",
		X"00",X"10",X"30",X"B8",X"F8",X"F8",X"F8",X"B8",X"80",X"80",X"80",X"80",X"80",X"80",X"C0",X"F0",
		X"00",X"30",X"03",X"07",X"00",X"00",X"00",X"00",X"E0",X"F0",X"3F",X"BF",X"1D",X"00",X"40",X"00",
		X"8B",X"EF",X"FF",X"FF",X"4E",X"44",X"33",X"CC",X"68",X"AC",X"0C",X"00",X"40",X"00",X"88",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"0F",X"07",X"00",X"80",X"62",X"FB",X"77",X"FF",X"3F",X"0F",
		X"60",X"70",X"70",X"F8",X"F0",X"F8",X"B8",X"8B",X"00",X"00",X"00",X"00",X"00",X"F0",X"E0",X"AC",
		X"03",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"48",X"F0",X"78",X"3C",X"8E",X"0E",X"10",X"00",
		X"CF",X"F7",X"FF",X"EF",X"BF",X"11",X"11",X"22",X"2C",X"04",X"20",X"00",X"00",X"CC",X"00",X"00",
		X"00",X"00",X"20",X"10",X"11",X"11",X"00",X"08",X"10",X"00",X"00",X"CC",X"FF",X"FE",X"FF",X"BF",
		X"80",X"C0",X"E0",X"E0",X"E0",X"F0",X"C3",X"83",X"00",X"00",X"00",X"00",X"E0",X"E0",X"E0",X"AC",
		X"0F",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"0F",X"0E",X"78",X"70",X"1E",X"5E",X"1E",X"00",
		X"9B",X"77",X"F7",X"FF",X"4E",X"00",X"00",X"40",X"08",X"98",X"08",X"00",X"99",X"66",X"44",X"88",
		X"00",X"00",X"00",X"40",X"30",X"11",X"11",X"00",X"70",X"30",X"30",X"30",X"FE",X"FE",X"FF",X"FF",
		X"00",X"80",X"D0",X"F0",X"96",X"07",X"27",X"DF",X"00",X"00",X"80",X"C0",X"C0",X"C0",X"E0",X"88",
		X"01",X"0F",X"0F",X"25",X"00",X"00",X"00",X"00",X"8E",X"1C",X"3C",X"4B",X"07",X"27",X"03",X"00",
		X"FF",X"F3",X"F7",X"E3",X"80",X"48",X"20",X"00",X"88",X"19",X"EE",X"44",X"22",X"44",X"00",X"00",
		X"10",X"00",X"00",X"00",X"00",X"33",X"F1",X"33",X"80",X"E0",X"F0",X"70",X"70",X"FC",X"EE",X"FF",
		X"00",X"10",X"70",X"F0",X"3C",X"5E",X"97",X"37",X"00",X"00",X"00",X"00",X"80",X"A0",X"00",X"11",
		X"00",X"00",X"03",X"0F",X"0F",X"00",X"00",X"00",X"EE",X"1C",X"3C",X"0F",X"0D",X"01",X"01",X"00",
		X"FF",X"F3",X"F7",X"48",X"68",X"AC",X"08",X"00",X"19",X"EE",X"2A",X"22",X"00",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"20",X"00",X"88",X"89",X"00",X"20",X"34",X"3C",X"5E",X"16",X"DE",X"CE",
		X"00",X"00",X"00",X"10",X"F0",X"F0",X"70",X"F1",X"00",X"00",X"00",X"C0",X"E0",X"C0",X"80",X"CC",
		X"77",X"89",X"88",X"00",X"20",X"00",X"00",X"00",X"FF",X"EC",X"FC",X"16",X"1E",X"5E",X"16",X"02",
		X"FF",X"1F",X"07",X"87",X"87",X"01",X"00",X"00",X"F8",X"CC",X"08",X"0C",X"0E",X"0C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"20",X"00",X"88",X"89",X"00",X"20",X"34",X"3C",X"5E",X"16",X"DE",X"CE",
		X"00",X"00",X"00",X"00",X"90",X"B0",X"70",X"F0",X"00",X"00",X"00",X"00",X"C0",X"E0",X"C0",X"CC",
		X"77",X"89",X"88",X"00",X"20",X"00",X"00",X"00",X"FF",X"EC",X"FC",X"16",X"1E",X"5E",X"16",X"02",
		X"FF",X"0F",X"07",X"83",X"81",X"00",X"00",X"00",X"F8",X"CC",X"0C",X"0E",X"0C",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"20",X"00",X"88",X"89",X"00",X"20",X"34",X"3C",X"5E",X"16",X"DE",X"CE",
		X"00",X"00",X"00",X"00",X"80",X"B0",X"70",X"F0",X"00",X"00",X"00",X"00",X"00",X"E0",X"F0",X"C0",
		X"77",X"89",X"88",X"00",X"20",X"00",X"00",X"00",X"FF",X"EC",X"FC",X"16",X"1E",X"5E",X"16",X"02",
		X"3F",X"0F",X"07",X"83",X"80",X"00",X"00",X"00",X"F8",X"0C",X"0F",X"0E",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"20",X"00",X"88",X"89",X"00",X"20",X"34",X"3C",X"5E",X"16",X"DE",X"CE",
		X"00",X"00",X"00",X"00",X"80",X"B0",X"70",X"F0",X"00",X"00",X"00",X"00",X"00",X"80",X"E0",X"F0",
		X"77",X"89",X"88",X"00",X"20",X"00",X"00",X"00",X"FF",X"EC",X"FC",X"16",X"1E",X"5E",X"16",X"02",
		X"0F",X"0F",X"07",X"83",X"80",X"00",X"00",X"00",X"3C",X"0F",X"0E",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"11",X"77",X"11",X"01",X"00",X"00",X"00",X"33",X"FF",X"FF",X"FF",X"03",
		X"00",X"00",X"66",X"FF",X"CD",X"CF",X"1E",X"78",X"00",X"00",X"00",X"04",X"0C",X"08",X"00",X"80",
		X"30",X"01",X"11",X"77",X"33",X"00",X"00",X"00",X"83",X"03",X"CC",X"EE",X"FF",X"BF",X"33",X"00",
		X"1E",X"0F",X"1E",X"03",X"89",X"EE",X"FF",X"FF",X"84",X"80",X"00",X"08",X"0C",X"04",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"11",X"33",X"FF",X"00",X"00",X"00",X"33",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"88",X"EE",X"CD",X"8F",X"16",X"3C",X"00",X"00",X"00",X"08",X"00",X"00",X"84",X"80",
		X"01",X"30",X"01",X"00",X"00",X"33",X"00",X"00",X"01",X"A2",X"77",X"77",X"FF",X"DF",X"77",X"00",
		X"1E",X"0F",X"00",X"FF",X"FF",X"FF",X"88",X"00",X"80",X"0E",X"00",X"CC",X"88",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"FF",X"00",X"00",X"00",X"33",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"FF",X"FF",X"FF",X"CC",X"33",X"00",X"00",X"00",X"CC",X"88",X"66",X"CC",X"CC",
		X"00",X"01",X"10",X"00",X"00",X"00",X"00",X"00",X"88",X"51",X"91",X"7F",X"33",X"77",X"44",X"88",
		X"FF",X"FF",X"FF",X"FF",X"6E",X"88",X"00",X"00",X"CC",X"88",X"88",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"11",X"11",X"33",X"33",X"33",X"00",X"00",X"FF",X"FF",X"FF",X"EE",X"EF",X"EE",
		X"00",X"04",X"04",X"24",X"2D",X"3C",X"4B",X"0F",X"00",X"00",X"00",X"80",X"00",X"80",X"1F",X"22",
		X"77",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"AB",X"00",X"48",X"95",X"11",X"33",X"33",X"22",
		X"04",X"33",X"FF",X"FF",X"FF",X"BF",X"00",X"00",X"EE",X"CC",X"CC",X"CC",X"88",X"00",X"00",X"00",
		X"00",X"11",X"11",X"33",X"77",X"77",X"77",X"57",X"CC",X"8A",X"8E",X"8A",X"9A",X"8B",X"8B",X"8B",
		X"00",X"00",X"00",X"02",X"E0",X"68",X"69",X"4B",X"00",X"00",X"00",X"00",X"00",X"04",X"0E",X"08",
		X"33",X"33",X"33",X"22",X"44",X"00",X"00",X"00",X"8B",X"89",X"88",X"48",X"53",X"11",X"11",X"33",
		X"1D",X"7F",X"FF",X"FF",X"FF",X"EE",X"88",X"00",X"EE",X"CC",X"CC",X"CC",X"88",X"00",X"00",X"00",
		X"00",X"00",X"00",X"11",X"33",X"33",X"77",X"77",X"44",X"46",X"CE",X"9A",X"9A",X"8B",X"CD",X"CD",
		X"00",X"00",X"04",X"E1",X"C3",X"97",X"1D",X"7F",X"00",X"00",X"00",X"08",X"00",X"88",X"CC",X"CC",
		X"77",X"57",X"33",X"33",X"33",X"22",X"00",X"00",X"CD",X"CC",X"CC",X"20",X"25",X"20",X"00",X"00",
		X"77",X"FF",X"77",X"FF",X"77",X"66",X"66",X"44",X"CC",X"CC",X"88",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"33",X"00",X"22",X"66",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"00",X"88",X"88",X"88",X"CC",X"CC",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"23",X"11",X"11",X"11",X"11",X"22",X"00",X"EE",X"EE",X"CC",X"DC",X"9A",X"10",X"00",X"00",
		X"FF",X"FF",X"77",X"77",X"3B",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"00",
		X"00",X"00",X"22",X"23",X"22",X"33",X"33",X"33",X"00",X"00",X"02",X"30",X"3C",X"16",X"07",X"89",
		X"00",X"04",X"26",X"B7",X"B7",X"3F",X"3F",X"3F",X"00",X"00",X"00",X"00",X"88",X"88",X"CC",X"CC",
		X"33",X"33",X"11",X"11",X"00",X"00",X"00",X"00",X"CC",X"EE",X"FF",X"7F",X"EE",X"66",X"22",X"22",
		X"3B",X"77",X"33",X"40",X"4A",X"40",X"00",X"00",X"EE",X"EE",X"EE",X"CC",X"44",X"44",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"8F",X"89",X"00",X"00",X"00",X"04",X"70",X"70",X"4B",X"0F",
		X"00",X"26",X"17",X"37",X"B7",X"B7",X"3F",X"3F",X"00",X"00",X"00",X"88",X"CC",X"CC",X"EE",X"EE",
		X"EE",X"77",X"33",X"33",X"11",X"00",X"00",X"00",X"03",X"CD",X"EE",X"FF",X"BF",X"77",X"11",X"00",
		X"3F",X"19",X"11",X"21",X"AC",X"88",X"88",X"CC",X"EE",X"CC",X"CC",X"44",X"22",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"00",X"10",X"8F",X"44",X"00",X"02",X"02",X"42",X"4B",X"C3",X"2D",X"0F",
		X"00",X"00",X"FF",X"FF",X"FF",X"77",X"7F",X"77",X"00",X"00",X"00",X"88",X"88",X"CC",X"CC",X"CC",
		X"77",X"33",X"33",X"33",X"11",X"00",X"00",X"00",X"02",X"CC",X"FF",X"FF",X"FF",X"DF",X"00",X"00",
		X"5D",X"00",X"21",X"9A",X"88",X"CC",X"CC",X"44",X"EE",X"77",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"33",X"11",X"66",X"33",X"33",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"33",X"CC",
		X"00",X"00",X"00",X"CC",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"88",X"CC",X"FF",
		X"33",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"67",X"11",X"00",X"00",
		X"11",X"A8",X"98",X"EF",X"CC",X"EE",X"22",X"11",X"00",X"08",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"00",X"00",X"12",X"10",X"00",X"00",X"11",X"77",X"3B",X"1F",X"86",X"C3",
		X"00",X"00",X"CC",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"88",X"CC",X"FF",X"00",
		X"10",X"07",X"00",X"33",X"11",X"00",X"00",X"00",X"87",X"0F",X"00",X"FF",X"FF",X"FF",X"11",X"00",
		X"08",X"54",X"EE",X"EE",X"FF",X"BF",X"EE",X"00",X"08",X"C0",X"08",X"00",X"00",X"CC",X"00",X"00",
		X"00",X"00",X"00",X"00",X"77",X"11",X"00",X"01",X"00",X"00",X"33",X"FF",X"FF",X"FF",X"FF",X"33",
		X"00",X"00",X"88",X"EE",X"FF",X"EE",X"8B",X"1E",X"00",X"00",X"00",X"00",X"00",X"0C",X"08",X"80",
		X"30",X"01",X"00",X"11",X"77",X"00",X"00",X"00",X"81",X"22",X"FF",X"FF",X"FF",X"BF",X"33",X"00",
		X"3C",X"1E",X"03",X"CC",X"FF",X"FF",X"CC",X"00",X"84",X"80",X"08",X"0C",X"EE",X"88",X"00",X"00",
		X"00",X"00",X"00",X"44",X"33",X"11",X"00",X"01",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"33",
		X"00",X"00",X"00",X"00",X"00",X"CC",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",
		X"30",X"01",X"00",X"11",X"33",X"44",X"00",X"00",X"80",X"33",X"FF",X"FF",X"DF",X"33",X"00",X"00",
		X"00",X"FF",X"FF",X"FF",X"EE",X"88",X"00",X"00",X"00",X"EE",X"CC",X"88",X"00",X"00",X"00",X"00",
		X"00",X"40",X"20",X"00",X"00",X"00",X"08",X"16",X"00",X"80",X"24",X"52",X"43",X"01",X"01",X"87",
		X"80",X"40",X"04",X"06",X"0E",X"0F",X"0F",X"4F",X"00",X"40",X"02",X"02",X"0E",X"0A",X"17",X"3F",
		X"03",X"21",X"10",X"43",X"01",X"00",X"10",X"00",X"4B",X"0F",X"0E",X"0F",X"0E",X"07",X"97",X"43",
		X"8F",X"1B",X"1F",X"4E",X"1F",X"37",X"19",X"3F",X"77",X"77",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"08",X"0C",X"C2",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"41",X"16",X"1A",X"0D",X"07",X"8B",
		X"00",X"06",X"0F",X"86",X"C2",X"0F",X"0F",X"06",X"00",X"00",X"08",X"00",X"40",X"0C",X"06",X"02",
		X"66",X"FF",X"DF",X"FF",X"FF",X"FF",X"FE",X"FF",X"EE",X"77",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",
		X"83",X"86",X"87",X"DB",X"DF",X"CF",X"EF",X"65",X"00",X"14",X"04",X"0A",X"0C",X"0C",X"86",X"82",
		X"00",X"00",X"00",X"33",X"00",X"01",X"43",X"13",X"00",X"00",X"66",X"11",X"F9",X"78",X"DE",X"EF",
		X"00",X"00",X"11",X"33",X"FF",X"FF",X"F1",X"F0",X"00",X"00",X"EE",X"00",X"00",X"88",X"CC",X"E6",
		X"13",X"40",X"00",X"00",X"33",X"00",X"00",X"00",X"67",X"CF",X"07",X"8F",X"11",X"66",X"00",X"00",
		X"78",X"78",X"1A",X"2D",X"33",X"11",X"00",X"00",X"E2",X"C0",X"80",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"00",X"00",X"00",X"22",X"55",X"10",X"01",X"00",X"00",X"00",X"FF",X"32",X"F1",X"78",X"DE",
		X"00",X"33",X"FF",X"F7",X"F1",X"3D",X"F7",X"F7",X"00",X"CC",X"88",X"88",X"80",X"E0",X"E0",X"84",
		X"53",X"13",X"00",X"20",X"00",X"00",X"00",X"00",X"67",X"EF",X"47",X"03",X"46",X"CC",X"11",X"00",
		X"78",X"69",X"0F",X"8D",X"DC",X"88",X"00",X"00",X"C8",X"C0",X"6A",X"7B",X"E2",X"00",X"00",X"00",
		X"00",X"00",X"00",X"11",X"00",X"22",X"55",X"10",X"00",X"10",X"32",X"B8",X"65",X"F0",X"F1",X"D2",
		X"EE",X"E6",X"E2",X"7A",X"F2",X"F4",X"ED",X"FC",X"00",X"00",X"00",X"C0",X"E0",X"2C",X"04",X"48",
		X"30",X"53",X"21",X"01",X"10",X"00",X"00",X"00",X"EF",X"EF",X"AB",X"01",X"23",X"22",X"66",X"00",
		X"F0",X"1E",X"0D",X"5E",X"22",X"44",X"00",X"00",X"CC",X"E6",X"7B",X"E2",X"CC",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"10",X"11",X"30",X"74",X"61",X"43",X"FC",X"F0",X"3C",
		X"88",X"C4",X"C4",X"F4",X"E5",X"F6",X"F8",X"E1",X"00",X"00",X"00",X"80",X"80",X"80",X"E6",X"F1",
		X"67",X"01",X"01",X"21",X"00",X"00",X"00",X"00",X"6F",X"BB",X"FF",X"6F",X"01",X"91",X"11",X"00",
		X"4B",X"0E",X"2F",X"2E",X"2A",X"22",X"00",X"00",X"79",X"2C",X"4C",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"44",X"44",X"44",X"99",X"77",X"77",X"FE",X"FE",X"F0",
		X"00",X"00",X"FF",X"FC",X"F0",X"F0",X"C3",X"C3",X"00",X"00",X"00",X"00",X"00",X"99",X"AA",X"EE",
		X"10",X"33",X"45",X"00",X"10",X"00",X"00",X"00",X"C3",X"F7",X"7F",X"5D",X"2E",X"02",X"20",X"00",
		X"58",X"1E",X"1F",X"1D",X"55",X"44",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"10",X"10",X"10",X"00",X"11",X"33",X"88",X"CC",X"F0",X"3D",X"1E",X"34",X"3C",X"8F",
		X"00",X"60",X"68",X"F0",X"FF",X"FC",X"DE",X"D2",X"00",X"00",X"22",X"EE",X"EE",X"EE",X"CC",X"C4",
		X"44",X"01",X"33",X"22",X"00",X"00",X"00",X"00",X"0F",X"3F",X"77",X"22",X"33",X"83",X"10",X"00",
		X"F2",X"79",X"E8",X"AC",X"6A",X"11",X"22",X"00",X"88",X"88",X"88",X"88",X"00",X"00",X"00",X"00",
		X"00",X"22",X"22",X"33",X"74",X"74",X"21",X"10",X"00",X"10",X"21",X"CA",X"E5",X"F2",X"3D",X"17",
		X"00",X"80",X"C0",X"79",X"F2",X"F4",X"E9",X"DA",X"00",X"00",X"44",X"CC",X"E6",X"E2",X"C0",X"80",
		X"33",X"22",X"00",X"00",X"11",X"11",X"00",X"00",X"E1",X"97",X"3F",X"AA",X"11",X"01",X"20",X"00",
		X"7B",X"BC",X"FC",X"DF",X"8E",X"0C",X"40",X"00",X"88",X"44",X"44",X"88",X"88",X"00",X"00",X"00",
		X"00",X"00",X"44",X"77",X"77",X"77",X"33",X"32",X"00",X"60",X"61",X"F0",X"FF",X"F3",X"B7",X"B4",
		X"11",X"33",X"F0",X"CB",X"87",X"C2",X"C3",X"1F",X"00",X"88",X"80",X"80",X"80",X"00",X"88",X"CC",
		X"11",X"11",X"11",X"11",X"00",X"00",X"00",X"00",X"F4",X"E9",X"71",X"53",X"65",X"88",X"44",X"00",
		X"0F",X"CF",X"EE",X"44",X"CC",X"1C",X"80",X"00",X"22",X"08",X"CC",X"44",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"55",X"77",X"00",X"00",X"FF",X"F3",X"F0",X"F0",X"3C",X"3C",
		X"22",X"22",X"99",X"EE",X"EE",X"F7",X"F7",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"22",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A1",X"87",X"8F",X"8B",X"AA",X"22",X"22",X"00",
		X"3C",X"FE",X"EF",X"AB",X"47",X"04",X"40",X"00",X"80",X"CC",X"2A",X"00",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"10",X"10",X"76",X"F8",X"11",X"32",X"32",X"F2",X"7A",X"F6",X"F1",X"78",
		X"88",X"C0",X"E2",X"68",X"2C",X"F3",X"F0",X"C3",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"80",
		X"E9",X"43",X"23",X"00",X"00",X"00",X"00",X"00",X"2D",X"07",X"4F",X"47",X"45",X"44",X"00",X"00",
		X"6F",X"DD",X"FF",X"6F",X"08",X"98",X"88",X"00",X"6E",X"08",X"08",X"48",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"30",X"70",X"43",X"02",X"21",X"77",X"76",X"74",X"E5",X"F4",X"F2",X"7B",X"F3",
		X"00",X"80",X"C4",X"D1",X"6A",X"F0",X"F8",X"B4",X"00",X"00",X"00",X"88",X"00",X"44",X"AA",X"80",
		X"33",X"76",X"ED",X"74",X"33",X"00",X"00",X"00",X"F0",X"87",X"0B",X"A7",X"44",X"22",X"00",X"00",
		X"7F",X"7F",X"5D",X"08",X"4C",X"44",X"66",X"00",X"C0",X"AC",X"48",X"08",X"80",X"00",X"00",X"00",
		X"00",X"33",X"11",X"11",X"10",X"70",X"70",X"12",X"00",X"CC",X"FF",X"FE",X"F8",X"CB",X"FE",X"FE",
		X"00",X"00",X"00",X"FF",X"C4",X"F8",X"E1",X"B7",X"00",X"00",X"00",X"00",X"44",X"AA",X"80",X"08",
		X"31",X"30",X"65",X"ED",X"74",X"00",X"00",X"00",X"E1",X"69",X"0F",X"1B",X"B3",X"11",X"00",X"00",
		X"6E",X"7F",X"2E",X"0C",X"26",X"33",X"88",X"00",X"AC",X"8C",X"00",X"40",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"33",X"00",X"01",X"43",X"13",X"00",X"00",X"66",X"11",X"F9",X"78",X"DE",X"67",
		X"00",X"00",X"33",X"73",X"B4",X"F8",X"F5",X"F7",X"00",X"00",X"EE",X"CC",X"CC",X"88",X"C8",X"E0",
		X"13",X"40",X"00",X"00",X"33",X"00",X"00",X"00",X"EF",X"CF",X"07",X"9F",X"11",X"66",X"00",X"00",
		X"7B",X"78",X"1A",X"2D",X"07",X"30",X"00",X"00",X"A4",X"C8",X"80",X"C4",X"C4",X"E6",X"00",X"00",
		X"00",X"00",X"00",X"33",X"00",X"01",X"43",X"13",X"00",X"00",X"66",X"11",X"F9",X"79",X"DE",X"EF",
		X"00",X"33",X"71",X"F1",X"B5",X"79",X"F6",X"FC",X"00",X"00",X"EE",X"88",X"88",X"80",X"C0",X"E0",
		X"13",X"40",X"00",X"00",X"33",X"00",X"00",X"00",X"67",X"DE",X"07",X"9E",X"11",X"66",X"00",X"00",
		X"FC",X"7A",X"3D",X"38",X"B4",X"70",X"33",X"00",X"2C",X"48",X"80",X"88",X"88",X"EE",X"00",X"00",
		X"00",X"21",X"00",X"00",X"00",X"20",X"00",X"00",X"87",X"03",X"0B",X"85",X"83",X"81",X"91",X"05",
		X"B7",X"B7",X"97",X"4B",X"2D",X"A5",X"F8",X"3C",X"FF",X"FF",X"7F",X"BF",X"3F",X"5B",X"69",X"96",
		X"00",X"12",X"03",X"00",X"00",X"10",X"00",X"00",X"43",X"A1",X"4B",X"2C",X"80",X"00",X"00",X"00",
		X"87",X"0F",X"0C",X"08",X"00",X"00",X"00",X"10",X"C3",X"2D",X"0F",X"07",X"02",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"3F",X"0F",X"1E",X"A5",X"F7",X"FF",X"EE",X"CC",X"21",X"42",X"94",X"28",
		X"16",X"70",X"30",X"61",X"03",X"83",X"03",X"D0",X"00",X"10",X"20",X"08",X"84",X"08",X"00",X"40",
		X"49",X"B4",X"1A",X"C2",X"0E",X"06",X"02",X"10",X"60",X"90",X"2C",X"43",X"10",X"70",X"03",X"00",
		X"41",X"A1",X"48",X"E0",X"C3",X"0F",X"0E",X"00",X"68",X"24",X"90",X"00",X"00",X"40",X"20",X"10",
		X"00",X"00",X"00",X"10",X"00",X"01",X"03",X"73",X"00",X"00",X"00",X"80",X"50",X"58",X"8F",X"CF",
		X"00",X"00",X"00",X"80",X"10",X"20",X"0E",X"0F",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"08",
		X"30",X"70",X"03",X"01",X"00",X"10",X"00",X"00",X"E6",X"C0",X"80",X"58",X"50",X"80",X"00",X"00",
		X"01",X"00",X"00",X"20",X"10",X"80",X"00",X"00",X"0C",X"08",X"00",X"00",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"30",X"00",X"01",X"03",X"00",X"00",X"00",X"00",X"10",X"C3",X"C0",X"EE",
		X"00",X"00",X"00",X"B0",X"07",X"0C",X"33",X"75",X"00",X"00",X"00",X"84",X"08",X"4C",X"88",X"CC",
		X"13",X"70",X"30",X"21",X"00",X"00",X"00",X"00",X"FA",X"E0",X"E0",X"78",X"2C",X"20",X"40",X"00",
		X"F3",X"07",X"00",X"00",X"40",X"20",X"00",X"00",X"EE",X"0F",X"00",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"12",X"03",X"01",X"05",X"00",X"11",X"19",X"33",X"10",
		X"08",X"00",X"71",X"C4",X"CC",X"FF",X"F3",X"F9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",
		X"13",X"16",X"70",X"30",X"21",X"00",X"00",X"00",X"FC",X"E1",X"E0",X"E0",X"2C",X"1C",X"20",X"40",
		X"F7",X"FF",X"07",X"00",X"00",X"00",X"00",X"00",X"CC",X"C8",X"80",X"0E",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"50",X"00",X"00",X"10",X"41",X"42",X"40",X"04",X"80",
		X"00",X"86",X"1B",X"22",X"77",X"FD",X"FB",X"E3",X"00",X"00",X"00",X"00",X"44",X"8E",X"0A",X"20",
		X"01",X"03",X"12",X"30",X"00",X"00",X"00",X"00",X"FF",X"F4",X"F0",X"F0",X"C3",X"86",X"00",X"00",
		X"02",X"00",X"30",X"80",X"80",X"40",X"80",X"00",X"40",X"00",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"20",X"20",X"A1",X"41",X"43",X"03",
		X"00",X"00",X"00",X"03",X"07",X"0C",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"C0",
		X"30",X"40",X"01",X"00",X"00",X"00",X"00",X"00",X"87",X"7E",X"7E",X"7C",X"F0",X"A1",X"20",X"00",
		X"00",X"10",X"A0",X"A0",X"2C",X"18",X"20",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"01",X"43",X"41",X"41",X"01",X"04",X"80",X"00",
		X"00",X"00",X"DD",X"EF",X"EE",X"EA",X"CE",X"84",X"00",X"00",X"04",X"0C",X"48",X"48",X"00",X"40",
		X"00",X"10",X"20",X"20",X"00",X"00",X"00",X"00",X"80",X"B3",X"7E",X"7E",X"3C",X"30",X"50",X"00",
		X"80",X"88",X"E0",X"F0",X"86",X"0C",X"00",X"00",X"80",X"00",X"00",X"00",X"80",X"80",X"00",X"00",
		X"00",X"04",X"02",X"01",X"00",X"00",X"00",X"00",X"44",X"C4",X"F7",X"F6",X"7E",X"37",X"37",X"02",
		X"11",X"99",X"FF",X"F7",X"F7",X"EE",X"66",X"80",X"00",X"81",X"81",X"81",X"02",X"02",X"04",X"08",
		X"00",X"00",X"10",X"10",X"00",X"00",X"00",X"00",X"10",X"F0",X"34",X"16",X"12",X"10",X"00",X"00",
		X"CD",X"FE",X"E7",X"C7",X"C6",X"40",X"00",X"00",X"00",X"80",X"40",X"40",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"10",X"10",X"10",X"00",X"10",X"00",X"00",X"5D",X"3F",X"37",X"32",X"13",X"01",
		X"04",X"AC",X"9E",X"9A",X"8A",X"89",X"81",X"80",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"10",X"70",X"52",X"83",X"81",X"00",X"00",
		X"90",X"F6",X"F3",X"E3",X"E3",X"78",X"40",X"00",X"00",X"C0",X"28",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"20",X"10",X"00",X"00",X"00",X"00",X"07",X"01",X"00",X"00",X"80",
		X"00",X"40",X"40",X"40",X"48",X"3C",X"06",X"16",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"C0",
		X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"80",X"20",X"20",X"41",X"40",X"20",X"00",
		X"07",X"73",X"F3",X"F1",X"78",X"2C",X"20",X"00",X"A0",X"18",X"0C",X"08",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"22",X"17",X"01",X"40",X"00",X"16",X"89",X"44",X"EE",X"FB",X"FD",X"7C",
		X"00",X"00",X"80",X"28",X"24",X"24",X"02",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"A0",
		X"20",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"07",X"01",X"C0",X"10",X"10",X"20",X"10",X"00",
		X"F7",X"F3",X"F1",X"F0",X"3C",X"16",X"00",X"00",X"08",X"0C",X"8C",X"C8",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"FC",X"76",X"77",X"FF",X"FC",
		X"08",X"08",X"04",X"04",X"02",X"02",X"8A",X"89",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"80",
		X"77",X"73",X"30",X"03",X"00",X"00",X"00",X"00",X"F9",X"FE",X"AF",X"0F",X"00",X"00",X"00",X"00",
		X"91",X"F3",X"78",X"70",X"70",X"C3",X"83",X"40",X"8C",X"8E",X"C6",X"E4",X"C0",X"48",X"00",X"00",
		X"00",X"00",X"03",X"00",X"22",X"11",X"33",X"77",X"00",X"00",X"D0",X"0E",X"03",X"CC",X"EA",X"FC",
		X"00",X"00",X"00",X"80",X"1C",X"34",X"77",X"F5",X"00",X"00",X"00",X"C0",X"00",X"08",X"0C",X"8C",
		X"0F",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"20",X"40",X"00",X"00",X"00",
		X"78",X"70",X"21",X"C3",X"40",X"20",X"00",X"00",X"E0",X"C0",X"28",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"00",X"01",X"03",X"73",X"00",X"00",X"00",X"80",X"40",X"69",X"CC",X"EE",
		X"00",X"00",X"00",X"40",X"83",X"0F",X"00",X"33",X"00",X"00",X"00",X"00",X"0E",X"0C",X"44",X"88",
		X"30",X"70",X"03",X"01",X"00",X"10",X"00",X"00",X"F6",X"E0",X"C0",X"68",X"40",X"80",X"00",X"00",
		X"F1",X"3F",X"03",X"00",X"82",X"40",X"00",X"00",X"CC",X"88",X"4C",X"04",X"02",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"00",X"01",X"03",X"73",X"00",X"00",X"00",X"80",X"41",X"48",X"CC",X"DD",
		X"00",X"01",X"06",X"08",X"10",X"33",X"FF",X"FF",X"00",X"0C",X"08",X"00",X"C0",X"EE",X"88",X"88",
		X"30",X"70",X"03",X"01",X"00",X"10",X"00",X"00",X"F4",X"D1",X"C1",X"48",X"40",X"80",X"00",X"00",
		X"F1",X"F0",X"FF",X"3F",X"12",X"01",X"00",X"00",X"CC",X"88",X"88",X"EE",X"C0",X"00",X"08",X"04",
		X"00",X"40",X"24",X"16",X"07",X"03",X"43",X"10",X"80",X"40",X"30",X"10",X"90",X"0A",X"14",X"03",
		X"00",X"00",X"C0",X"40",X"84",X"40",X"4A",X"2C",X"00",X"00",X"08",X"01",X"0C",X"0D",X"AE",X"E9",
		X"00",X"80",X"60",X"01",X"00",X"00",X"00",X"20",X"81",X"86",X"04",X"02",X"00",X"A1",X"20",X"50",
		X"07",X"24",X"20",X"02",X"53",X"37",X"A7",X"97",X"80",X"33",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"A0",X"04",X"84",X"02",X"04",X"82",X"10",X"40",X"20",X"82",X"52",X"50",X"2B",X"48",
		X"00",X"00",X"A0",X"61",X"87",X"0A",X"24",X"49",X"20",X"40",X"08",X"00",X"0C",X"2C",X"3C",X"1E",
		X"FF",X"DD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"70",X"03",X"9E",X"CD",X"AF",X"EF",X"FC",
		X"01",X"0E",X"83",X"04",X"92",X"0D",X"83",X"D2",X"16",X"43",X"81",X"09",X"40",X"08",X"20",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"13",X"00",X"00",X"20",X"A0",X"60",X"4C",X"DD",X"EE",
		X"00",X"00",X"00",X"0F",X"03",X"01",X"88",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"08",X"00",
		X"30",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"B3",X"69",X"48",X"59",X"60",X"A0",X"20",X"00",
		X"ED",X"0F",X"01",X"00",X"89",X"09",X"00",X"00",X"80",X"00",X"08",X"08",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"01",X"00",X"00",X"01",X"42",X"40",X"D1",X"CC",X"EE",
		X"00",X"0E",X"03",X"01",X"01",X"99",X"13",X"36",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"13",X"30",X"33",X"00",X"00",X"00",X"00",X"00",X"FF",X"B1",X"2C",X"2C",X"24",X"30",X"20",X"00",
		X"FC",X"0F",X"03",X"88",X"CC",X"00",X"84",X"00",X"88",X"88",X"08",X"0C",X"04",X"04",X"08",X"00",
		X"00",X"00",X"00",X"10",X"00",X"30",X"00",X"01",X"00",X"07",X"0F",X"08",X"00",X"22",X"AA",X"8D",
		X"00",X"00",X"00",X"44",X"66",X"77",X"21",X"FE",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"88",
		X"01",X"11",X"11",X"11",X"00",X"00",X"00",X"00",X"FF",X"D1",X"96",X"BD",X"12",X"10",X"10",X"00",
		X"BF",X"0F",X"00",X"44",X"66",X"00",X"42",X"00",X"88",X"88",X"4C",X"04",X"04",X"04",X"08",X"00",
		X"00",X"00",X"00",X"00",X"00",X"20",X"10",X"70",X"00",X"07",X"0C",X"08",X"08",X"3B",X"2A",X"0C",
		X"00",X"00",X"08",X"00",X"76",X"57",X"76",X"8F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",
		X"01",X"01",X"01",X"11",X"00",X"00",X"00",X"00",X"FF",X"DD",X"DA",X"96",X"87",X"00",X"00",X"00",
		X"0C",X"08",X"33",X"2A",X"C0",X"A0",X"80",X"00",X"0E",X"02",X"02",X"04",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"03",X"07",X"0C",X"08",X"11",X"A2",
		X"00",X"00",X"08",X"0C",X"24",X"47",X"46",X"8C",X"00",X"00",X"00",X"00",X"00",X"0C",X"02",X"02",
		X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"89",X"7F",X"6E",X"6D",X"4B",X"02",X"00",X"00",
		X"9D",X"BB",X"AA",X"D4",X"E4",X"20",X"00",X"00",X"02",X"00",X"04",X"00",X"80",X"00",X"00",X"00",
		X"00",X"00",X"01",X"02",X"00",X"00",X"02",X"20",X"00",X"00",X"0C",X"17",X"03",X"03",X"89",X"CD",
		X"00",X"00",X"00",X"C8",X"F3",X"C6",X"8C",X"99",X"00",X"00",X"00",X"00",X"0E",X"03",X"01",X"01",
		X"10",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"F0",X"0E",X"16",X"32",X"32",X"00",X"00",
		X"99",X"CC",X"FE",X"FE",X"8C",X"08",X"00",X"00",X"02",X"04",X"C0",X"00",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"03",X"04",X"04",X"00",X"00",X"00",X"00",X"DC",X"3E",X"17",X"03",
		X"00",X"00",X"00",X"80",X"5D",X"E7",X"CC",X"88",X"00",X"00",X"00",X"00",X"88",X"0E",X"07",X"03",
		X"15",X"20",X"00",X"10",X"00",X"00",X"00",X"00",X"CD",X"10",X"F0",X"07",X"03",X"01",X"00",X"00",
		X"BB",X"CC",X"77",X"E7",X"C6",X"84",X"00",X"00",X"03",X"24",X"80",X"40",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"06",X"04",X"04",X"00",X"00",X"00",X"10",X"7E",X"13",X"01",X"44",
		X"00",X"00",X"01",X"CF",X"86",X"86",X"8C",X"9D",X"00",X"00",X"0C",X"02",X"00",X"00",X"8A",X"A8",
		X"02",X"01",X"10",X"00",X"00",X"00",X"00",X"00",X"44",X"11",X"F3",X"73",X"81",X"00",X"00",X"00",
		X"CC",X"F8",X"8B",X"CB",X"EA",X"6A",X"00",X"00",X"40",X"E0",X"08",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"03",X"04",X"04",X"00",X"00",X"01",X"03",X"42",X"2E",X"26",X"13",
		X"00",X"00",X"0C",X"0E",X"03",X"01",X"88",X"54",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",
		X"04",X"00",X"02",X"00",X"10",X"00",X"00",X"00",X"9B",X"DD",X"55",X"B2",X"72",X"40",X"00",X"00",
		X"19",X"EF",X"67",X"6B",X"2D",X"04",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"01",X"00",X"E6",X"AE",X"E6",X"1F",
		X"00",X"0E",X"03",X"01",X"01",X"CD",X"45",X"03",X"00",X"00",X"00",X"00",X"00",X"40",X"80",X"E0",
		X"07",X"04",X"04",X"02",X"00",X"00",X"00",X"00",X"03",X"01",X"CC",X"45",X"30",X"50",X"10",X"00",
		X"FF",X"BB",X"B5",X"96",X"1E",X"00",X"00",X"00",X"08",X"08",X"08",X"88",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"11",X"00",X"00",X"00",X"22",X"66",X"EE",X"48",X"F7",
		X"00",X"0E",X"0F",X"01",X"00",X"44",X"55",X"1B",X"00",X"00",X"00",X"80",X"00",X"C0",X"00",X"08",
		X"11",X"11",X"23",X"02",X"02",X"02",X"01",X"00",X"DF",X"0F",X"00",X"22",X"66",X"00",X"24",X"00",
		X"FF",X"B8",X"96",X"DB",X"84",X"80",X"80",X"00",X"08",X"88",X"88",X"88",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"07",X"0C",X"08",X"08",X"99",X"8C",X"C6",
		X"00",X"00",X"08",X"24",X"20",X"B8",X"33",X"77",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"08",
		X"11",X"11",X"01",X"03",X"02",X"02",X"01",X"00",X"F3",X"0F",X"0C",X"11",X"33",X"00",X"12",X"00",
		X"FF",X"D8",X"43",X"43",X"42",X"C0",X"40",X"00",X"8C",X"C0",X"CC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"13",X"00",X"00",X"20",X"A1",X"42",X"4C",X"DD",X"EE",
		X"00",X"00",X"0F",X"09",X"00",X"00",X"9B",X"33",X"00",X"00",X"00",X"08",X"08",X"00",X"00",X"00",
		X"30",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"B0",X"69",X"48",X"59",X"51",X"A0",X"20",X"00",
		X"E5",X"3E",X"17",X"03",X"89",X"00",X"09",X"00",X"80",X"00",X"00",X"00",X"08",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"13",X"00",X"01",X"21",X"82",X"40",X"5D",X"DD",X"EE",
		X"00",X"0C",X"0E",X"06",X"13",X"13",X"33",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"B0",X"69",X"48",X"59",X"51",X"91",X"20",X"01",
		X"E5",X"7C",X"3F",X"17",X"13",X"02",X"02",X"0C",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"30",X"80",X"10",X"30",X"40",X"01",X"70",X"86",X"0B",X"87",X"0A",X"04",X"0B",X"14",
		X"C2",X"C2",X"61",X"61",X"16",X"40",X"29",X"18",X"FF",X"77",X"11",X"86",X"4B",X"B4",X"40",X"68",
		X"03",X"40",X"80",X"10",X"42",X"30",X"20",X"40",X"20",X"01",X"82",X"43",X"E0",X"90",X"00",X"00",
		X"09",X"01",X"1A",X"50",X"A0",X"40",X"10",X"10",X"49",X"A1",X"E0",X"40",X"83",X"96",X"07",X"00",
		X"FF",X"FF",X"EE",X"03",X"A5",X"4B",X"D2",X"E0",X"01",X"40",X"82",X"16",X"A4",X"C2",X"80",X"40",
		X"B4",X"A0",X"49",X"16",X"28",X"04",X"08",X"03",X"00",X"80",X"C0",X"80",X"00",X"00",X"00",X"A0",
		X"92",X"04",X"18",X"06",X"4A",X"E1",X"0F",X"2C",X"02",X"29",X"40",X"84",X"42",X"38",X"10",X"00",
		X"10",X"4D",X"1C",X"60",X"B0",X"14",X"21",X"F0",X"40",X"80",X"40",X"80",X"C0",X"C0",X"C2",X"10");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
