module rom();


localparam ROM = {
	8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h7E,8'h81,8'hA5,8'h81,8'h81,8'hBD,8'h99,8'h81,8'h81,8'h7E,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h7E,8'hFF,8'hDB,8'hFF,8'hFF,8'hC3,8'hE7,8'hFF,8'hFF,8'h7E,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h00,8'h00,8'h6C,8'hFE,8'hFE,8'hFE,8'hFE,8'h7C,8'h38,8'h10,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h00,8'h00,8'h10,8'h38,8'h7C,8'hFE,8'h7C,8'h38,8'h10,8'h00,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h00,8'h18,8'h3C,8'h3C,8'hE7,8'hE7,8'hE7,8'h18,8'h18,8'h3C,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h00,8'h18,8'h3C,8'h7E,8'hFF,8'hFF,8'h7E,8'h18,8'h18,8'h3C,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h18,8'h3C,8'h3C,8'h18,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
	8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hE7,8'hC3,8'hC3,8'hE7,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,
	8'h00,8'h00,8'h00,8'h00,8'h00,8'h3C,8'h66,8'h42,8'h42,8'h66,8'h3C,8'h00,8'h00,8'h00,8'h00,8'h00,
	8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hC3,8'h99,8'hBD,8'hBD,8'h99,8'hC3,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,
	8'h00,8'h00,8'h1E,8'h0E,8'h1A,8'h32,8'h78,"11001100","11001100","11001100","11001100",8'h78,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h3C,8'h66,8'h66,8'h66,8'h66,8'h3C,8'h18,8'h7E,8'h18,8'h18,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,"00111111","00110011","00111111","00110000","00110000","00110000","00110000","01110000","11110000","11100000",8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,"01111111","01100011","01111111","01100011","01100011","01100011","01100011","01100111",8'hE7,"11100110","11000000",8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h00,8'h18,8'h18,8'hDB,8'h3C,8'hE7,8'h3C,8'hDB,8'h18,8'h18,8'h00,8'h00,8'h00,8'h00,
	8'h00,"10000000","11000000","11100000","11110000","11111000",8'hFE,"11111000","11110000","11100000","11000000","10000000",8'h00,8'h00,8'h00,8'h00,
	8'h00,"00000010","00000110",8'h0E,8'h1E,"00111110",8'hFE,"00111110",8'h1E,8'h0E,"00000110","00000010",8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h18,8'h3C,8'h7E,8'h18,8'h18,8'h18,8'h7E,8'h3C,8'h18,8'h00,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h66,8'h66,8'h66,8'h66,8'h66,8'h66,8'h66,8'h00,8'h66,8'h66,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,"01111111",8'hDB,8'hDB,8'hDB,"01111011","00011011","00011011","00011011","00011011","00011011",8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h7C,8'hC6,"01100000",8'h38,8'h6C,8'hC6,8'hC6,8'h6C,8'h38,"00001100",8'hC6,8'h7C,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hFE,8'hFE,8'hFE,8'hFE,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h18,8'h3C,8'h7E,8'h18,8'h18,8'h18,8'h7E,8'h3C,8'h18,8'h7E,"00110000",8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h18,8'h3C,8'h7E,8'h18,8'h18,8'h18,8'h18,8'h18,8'h18,8'h18,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h18,8'h18,8'h18,8'h18,8'h18,8'h18,8'h18,8'h7E,8'h3C,8'h18,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h00,8'h00,8'h00,8'h18,"00001100",8'hFE,"00001100",8'h18,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h00,8'h00,8'h00,"00110000","01100000",8'hFE,"01100000","00110000",8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,"11000000","11000000","11000000",8'hFE,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h00,8'h00,8'h00,"00100100",8'h66,8'hFF,8'h66,"00100100",8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h00,8'h00,8'h10,8'h38,8'h38,8'h7C,8'h7C,8'hFE,8'hFE,8'h00,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h00,8'h00,8'hFE,8'hFE,8'h7C,8'h7C,8'h38,8'h38,8'h10,8'h00,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h18,8'h3C,8'h3C,8'h3C,8'h18,8'h18,8'h18,8'h00,8'h18,8'h18,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h66,8'h66,8'h66,"00100100",8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h00,8'h6C,8'h6C,8'hFE,8'h6C,8'h6C,8'h6C,8'hFE,8'h6C,8'h6C,8'h00,8'h00,8'h00,8'h00,
	8'h18,8'h18,8'h7C,8'hC6,"11000010","11000000",8'h7C,"00000110","00000110","10000110",8'hC6,8'h7C,8'h18,8'h18,8'h00,8'h00,
	8'h00,8'h00,8'h00,8'h00,"11000010",8'hC6,"00001100",8'h18,"00110000","01100000",8'hC6,"10000110",8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h38,8'h6C,8'h6C,8'h38,"01110110","11011100","11001100","11001100","11001100","01110110",8'h00,8'h00,8'h00,8'h00,
	8'h00,"00110000","00110000","00110000","01100000",8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,"00001100",8'h18,"00110000","00110000","00110000","00110000","00110000","00110000",8'h18,"00001100",8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,"00110000",8'h18,"00001100","00001100","00001100","00001100","00001100","00001100",8'h18,"00110000",8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h00,8'h00,8'h00,8'h66,8'h3C,8'hFF,8'h3C,8'h66,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h00,8'h00,8'h00,8'h18,8'h18,8'h7E,8'h18,8'h18,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h18,8'h18,8'h18,"00110000",8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h7E,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h18,8'h18,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h00,8'h00,"00000010","00000110","00001100",8'h18,"00110000","01100000","11000000","10000000",8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h7C,8'hC6,8'hC6,"11001110","11011110","11110110","11100110",8'hC6,8'hC6,8'h7C,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h18,8'h38,8'h78,8'h18,8'h18,8'h18,8'h18,8'h18,8'h18,8'h7E,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h7C,8'hC6,"00000110","00001100",8'h18,"00110000","01100000","11000000",8'hC6,8'hFE,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h7C,8'hC6,"00000110","00000110",8'h3C,"00000110","00000110","00000110",8'hC6,8'h7C,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,"00001100","00011100",8'h3C,8'h6C,"11001100",8'hFE,"00001100","00001100","00001100",8'h1E,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'hFE,"11000000","11000000","11000000","11111100","00000110","00000110","00000110",8'hC6,8'h7C,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h38,"01100000","11000000","11000000","11111100",8'hC6,8'hC6,8'hC6,8'hC6,8'h7C,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'hFE,8'hC6,"00000110","00000110","00001100",8'h18,"00110000","00110000","00110000","00110000",8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h7C,8'hC6,8'hC6,8'hC6,8'h7C,8'hC6,8'hC6,8'hC6,8'hC6,8'h7C,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h7C,8'hC6,8'hC6,8'hC6,8'h7E,"00000110","00000110","00000110","00001100",8'h78,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h00,8'h00,8'h18,8'h18,8'h00,8'h00,8'h00,8'h18,8'h18,8'h00,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h00,8'h00,8'h18,8'h18,8'h00,8'h00,8'h00,8'h18,8'h18,"00110000",8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h00,"00000110","00001100",8'h18,"00110000","01100000","00110000",8'h18,"00001100","00000110",8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h00,8'h00,8'h00,8'h7E,8'h00,8'h00,8'h7E,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h00,"01100000","00110000",8'h18,"00001100","00000110","00001100",8'h18,"00110000","01100000",8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h7C,8'hC6,8'hC6,"00001100",8'h18,8'h18,8'h18,8'h00,8'h18,8'h18,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h7C,8'hC6,8'hC6,8'hC6,"11011110","11011110","11011110","11011100","11000000",8'h7C,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h10,8'h38,8'h6C,8'hC6,8'hC6,8'hFE,8'hC6,8'hC6,8'hC6,8'hC6,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,"11111100",8'h66,8'h66,8'h66,8'h7C,8'h66,8'h66,8'h66,8'h66,"11111100",8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h3C,8'h66,"11000010","11000000","11000000","11000000","11000000","11000010",8'h66,8'h3C,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,"11111000",8'h6C,8'h66,8'h66,8'h66,8'h66,8'h66,8'h66,8'h6C,"11111000",8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'hFE,8'h66,"01100010","01101000",8'h78,"01101000","01100000","01100010",8'h66,8'hFE,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'hFE,8'h66,"01100010","01101000",8'h78,"01101000","01100000","01100000","01100000","11110000",8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h3C,8'h66,"11000010","11000000","11000000","11011110",8'hC6,8'hC6,8'h66,"00111010",8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'hC6,8'hC6,8'hC6,8'hC6,8'hFE,8'hC6,8'hC6,8'hC6,8'hC6,8'hC6,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h3C,8'h18,8'h18,8'h18,8'h18,8'h18,8'h18,8'h18,8'h18,8'h3C,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h1E,"00001100","00001100","00001100","00001100","00001100","11001100","11001100","11001100",8'h78,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,"11100110",8'h66,8'h66,8'h6C,8'h78,8'h78,8'h6C,8'h66,8'h66,"11100110",8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,"11110000","01100000","01100000","01100000","01100000","01100000","01100000","01100010",8'h66,8'hFE,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'hC3,8'hE7,8'hFF,8'hFF,8'hDB,8'hC3,8'hC3,8'hC3,8'hC3,8'hC3,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'hC6,"11100110","11110110",8'hFE,"11011110","11001110",8'hC6,8'hC6,8'hC6,8'hC6,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h7C,8'hC6,8'hC6,8'hC6,8'hC6,8'hC6,8'hC6,8'hC6,8'hC6,8'h7C,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,"11111100",8'h66,8'h66,8'h66,8'h7C,"01100000","01100000","01100000","01100000","11110000",8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h7C,8'hC6,8'hC6,8'hC6,8'hC6,8'hC6,8'hC6,"11010110","11011110",8'h7C,"00001100",8'h0E,8'h00,8'h00,
	8'h00,8'h00,"11111100",8'h66,8'h66,8'h66,8'h7C,8'h6C,8'h66,8'h66,8'h66,"11100110",8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h7C,8'hC6,8'hC6,"01100000",8'h38,"00001100","00000110",8'hC6,8'hC6,8'h7C,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'hFF,8'hDB,8'h99,8'h18,8'h18,8'h18,8'h18,8'h18,8'h18,8'h3C,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'hC6,8'hC6,8'hC6,8'hC6,8'hC6,8'hC6,8'hC6,8'hC6,8'hC6,8'h7C,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'hC3,8'hC3,8'hC3,8'hC3,8'hC3,8'hC3,8'hC3,8'h66,8'h3C,8'h18,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'hC3,8'hC3,8'hC3,8'hC3,8'hC3,8'hDB,8'hDB,8'hFF,8'h66,8'h66,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'hC3,8'hC3,8'h66,8'h3C,8'h18,8'h18,8'h3C,8'h66,8'hC3,8'hC3,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'hC3,8'hC3,8'hC3,8'h66,8'h3C,8'h18,8'h18,8'h18,8'h18,8'h3C,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'hFF,8'hC3,"10000110","00001100",8'h18,"00110000","01100000","11000001",8'hC3,8'hFF,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h3C,"00110000","00110000","00110000","00110000","00110000","00110000","00110000","00110000",8'h3C,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h00,"10000000","11000000","11100000","01110000",8'h38,"00011100",8'h0E,"00000110","00000010",8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h3C,"00001100","00001100","00001100","00001100","00001100","00001100","00001100","00001100",8'h3C,8'h00,8'h00,8'h00,8'h00,
	8'h10,8'h38,8'h6C,8'hC6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hFF,8'h00,8'h00,
	"00110000","00110000",8'h18,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h00,8'h00,8'h00,8'h78,"00001100",8'h7C,"11001100","11001100","11001100","01110110",8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,"11100000","01100000","01100000",8'h78,8'h6C,8'h66,8'h66,8'h66,8'h66,8'h7C,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h00,8'h00,8'h00,8'h7C,8'hC6,"11000000","11000000","11000000",8'hC6,8'h7C,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,"00011100","00001100","00001100",8'h3C,8'h6C,"11001100","11001100","11001100","11001100","01110110",8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h00,8'h00,8'h00,8'h7C,8'hC6,8'hFE,"11000000","11000000",8'hC6,8'h7C,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h38,8'h6C,"01100100","01100000","11110000","01100000","01100000","01100000","01100000","11110000",8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h00,8'h00,8'h00,"01110110","11001100","11001100","11001100","11001100","11001100",8'h7C,"00001100","11001100",8'h78,8'h00,
	8'h00,8'h00,"11100000","01100000","01100000",8'h6C,"01110110",8'h66,8'h66,8'h66,8'h66,"11100110",8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h18,8'h18,8'h00,8'h38,8'h18,8'h18,8'h18,8'h18,8'h18,8'h3C,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,"00000110","00000110",8'h00,8'h0E,"00000110","00000110","00000110","00000110","00000110","00000110",8'h66,8'h66,8'h3C,8'h00,
	8'h00,8'h00,"11100000","01100000","01100000",8'h66,8'h6C,8'h78,8'h78,8'h6C,8'h66,"11100110",8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h38,8'h18,8'h18,8'h18,8'h18,8'h18,8'h18,8'h18,8'h18,8'h3C,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h00,8'h00,8'h00,"11100110",8'hFF,8'hDB,8'hDB,8'hDB,8'hDB,8'hDB,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h00,8'h00,8'h00,"11011100",8'h66,8'h66,8'h66,8'h66,8'h66,8'h66,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h00,8'h00,8'h00,8'h7C,8'hC6,8'hC6,8'hC6,8'hC6,8'hC6,8'h7C,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h00,8'h00,8'h00,"11011100",8'h66,8'h66,8'h66,8'h66,8'h66,8'h7C,"01100000","01100000","11110000",8'h00,
	8'h00,8'h00,8'h00,8'h00,8'h00,"01110110","11001100","11001100","11001100","11001100","11001100",8'h7C,"00001100","00001100",8'h1E,8'h00,
	8'h00,8'h00,8'h00,8'h00,8'h00,"11011100","01110110",8'h66,"01100000","01100000","01100000","11110000",8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h00,8'h00,8'h00,8'h7C,8'hC6,"01100000",8'h38,"00001100",8'hC6,8'h7C,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h10,"00110000","00110000","11111100","00110000","00110000","00110000","00110000","00110110","00011100",8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h00,8'h00,8'h00,"11001100","11001100","11001100","11001100","11001100","11001100","01110110",8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h00,8'h00,8'h00,8'hC3,8'hC3,8'hC3,8'hC3,8'h66,8'h3C,8'h18,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h00,8'h00,8'h00,8'hC3,8'hC3,8'hC3,8'hDB,8'hDB,8'hFF,8'h66,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h00,8'h00,8'h00,8'hC3,8'h66,8'h3C,8'h18,8'h3C,8'h66,8'hC3,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h00,8'h00,8'h00,8'hC6,8'hC6,8'hC6,8'hC6,8'hC6,8'hC6,8'h7E,"00000110","00001100","11111000",8'h00,
	8'h00,8'h00,8'h00,8'h00,8'h00,8'hFE,"11001100",8'h18,"00110000","01100000",8'hC6,8'hFE,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h0E,8'h18,8'h18,8'h18,"01110000",8'h18,8'h18,8'h18,8'h18,8'h0E,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h18,8'h18,8'h18,8'h18,8'h00,8'h18,8'h18,8'h18,8'h18,8'h18,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,"01110000",8'h18,8'h18,8'h18,8'h0E,8'h18,8'h18,8'h18,8'h18,"01110000",8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,"01110110","11011100",8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
	8'h00,8'h00,8'h00,8'h00,8'h10,8'h38,8'h6C,8'hC6,8'hC6,8'hC6,8'hFE,8'h00,8'h00,8'h00,8'h00,8'h00
	};
	
	endmodule