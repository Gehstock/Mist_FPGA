`define BUILD_DATE "180708"
`define BUILD_TIME "073707"
