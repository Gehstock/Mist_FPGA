library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ckong_tile_bit1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ckong_tile_bit1 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"38",X"7C",X"C2",X"82",X"86",X"7C",X"38",X"00",X"02",X"02",X"FE",X"FE",X"42",X"02",X"00",X"00",
		X"62",X"F2",X"BA",X"9A",X"9E",X"CE",X"46",X"00",X"8C",X"DE",X"F2",X"B2",X"92",X"86",X"04",X"00",
		X"08",X"FE",X"FE",X"C8",X"68",X"38",X"18",X"00",X"1C",X"BE",X"A2",X"A2",X"A2",X"E6",X"E4",X"00",
		X"0C",X"9E",X"92",X"92",X"D2",X"7E",X"3C",X"00",X"C0",X"E0",X"B0",X"9E",X"8E",X"C0",X"C0",X"00",
		X"0C",X"6E",X"9A",X"9A",X"B2",X"F2",X"6C",X"00",X"78",X"FC",X"96",X"92",X"92",X"F2",X"60",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"18",X"24",X"62",X"51",X"85",X"46",X"24",X"18",X"18",X"24",X"46",X"89",X"91",X"62",X"24",X"18",
		X"18",X"24",X"42",X"D5",X"AB",X"42",X"24",X"18",X"00",X"00",X"80",X"80",X"80",X"80",X"FF",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"7E",X"C8",X"88",X"C8",X"7E",X"3E",X"00",
		X"6C",X"FE",X"92",X"92",X"92",X"FE",X"FE",X"00",X"44",X"C6",X"82",X"82",X"C6",X"7C",X"38",X"00",
		X"38",X"7C",X"C6",X"82",X"82",X"FE",X"FE",X"00",X"82",X"92",X"92",X"92",X"FE",X"FE",X"00",X"00",
		X"80",X"90",X"90",X"90",X"90",X"FE",X"FE",X"00",X"9E",X"9E",X"92",X"82",X"C6",X"7C",X"38",X"00",
		X"FE",X"FE",X"10",X"10",X"10",X"FE",X"FE",X"00",X"82",X"82",X"FE",X"FE",X"82",X"82",X"00",X"00",
		X"FC",X"FE",X"02",X"02",X"02",X"06",X"04",X"00",X"82",X"C6",X"6E",X"3C",X"18",X"FE",X"FE",X"00",
		X"02",X"02",X"02",X"02",X"FE",X"FE",X"00",X"00",X"FE",X"FE",X"70",X"38",X"70",X"FE",X"FE",X"00",
		X"FE",X"FE",X"1C",X"38",X"70",X"FE",X"FE",X"00",X"7C",X"FE",X"82",X"82",X"82",X"FE",X"7C",X"00",
		X"70",X"F8",X"88",X"88",X"88",X"FE",X"FE",X"00",X"7A",X"FC",X"8E",X"8A",X"82",X"FE",X"7C",X"00",
		X"72",X"F6",X"9E",X"8C",X"88",X"FE",X"FE",X"00",X"0C",X"5E",X"D2",X"92",X"92",X"F6",X"64",X"00",
		X"80",X"80",X"FE",X"FE",X"80",X"80",X"00",X"00",X"FC",X"FE",X"02",X"02",X"02",X"FE",X"FC",X"00",
		X"F0",X"F8",X"1C",X"0E",X"1C",X"F8",X"F0",X"00",X"F8",X"FE",X"1C",X"38",X"1C",X"FE",X"F8",X"00",
		X"C6",X"EE",X"7C",X"38",X"7C",X"EE",X"C6",X"00",X"C0",X"F0",X"1E",X"1E",X"F0",X"C0",X"00",X"00",
		X"C2",X"E2",X"F2",X"BA",X"9E",X"8E",X"86",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"00",X"00",
		X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"00",X"00",X"40",X"40",X"40",X"40",X"40",X"40",X"00",
		X"00",X"00",X"00",X"00",X"28",X"00",X"00",X"00",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",
		X"00",X"00",X"82",X"C6",X"6C",X"38",X"00",X"00",X"00",X"00",X"38",X"6C",X"C6",X"82",X"00",X"00",
		X"00",X"00",X"82",X"FE",X"FE",X"82",X"00",X"00",X"82",X"FE",X"FE",X"82",X"82",X"FE",X"FE",X"82",
		X"00",X"28",X"28",X"28",X"28",X"28",X"28",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"00",
		X"F6",X"F6",X"00",X"00",X"F6",X"F6",X"00",X"00",X"FA",X"FA",X"00",X"00",X"FA",X"FA",X"00",X"00",
		X"00",X"00",X"00",X"F6",X"F6",X"00",X"00",X"00",X"00",X"00",X"00",X"FA",X"FA",X"00",X"00",X"00",
		X"00",X"00",X"00",X"E0",X"C0",X"00",X"00",X"00",X"00",X"E0",X"C0",X"00",X"E0",X"C0",X"00",X"00",
		X"00",X"60",X"E0",X"00",X"60",X"E0",X"00",X"00",X"00",X"00",X"C0",X"00",X"C0",X"00",X"00",X"00",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"FF",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"FF",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"FF",
		X"00",X"00",X"00",X"00",X"06",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"06",X"00",X"00",
		X"38",X"28",X"3E",X"00",X"00",X"00",X"00",X"00",X"3E",X"00",X"3C",X"02",X"02",X"3C",X"00",X"0E",
		X"22",X"2A",X"3E",X"00",X"00",X"0E",X"3A",X"2A",X"22",X"3E",X"00",X"3E",X"08",X"10",X"3E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"22",X"A5",X"BD",X"81",X"42",X"3C",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"3C",X"42",X"81",X"A5",X"7C",X"40",X"00",X"38",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"04",X"02",X"84",X"48",X"12",X"12",X"12",X"12",
		X"FE",X"44",X"44",X"44",X"44",X"44",X"44",X"FF",X"17",X"14",X"14",X"52",X"42",X"42",X"44",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"A2",X"00",X"F0",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",
		X"00",X"01",X"0F",X"3F",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"0F",
		X"54",X"A6",X"02",X"02",X"62",X"73",X"77",X"FF",X"FF",X"8F",X"76",X"7C",X"4E",X"A6",X"D7",X"A3",
		X"FF",X"FF",X"FE",X"FD",X"7F",X"87",X"03",X"80",X"1F",X"3F",X"78",X"F0",X"F1",X"F6",X"F8",X"6F",
		X"BF",X"5F",X"AF",X"4F",X"2A",X"90",X"40",X"A8",X"C1",X"61",X"51",X"25",X"35",X"A1",X"B2",X"AE",
		X"CE",X"9A",X"31",X"3B",X"BF",X"3F",X"1D",X"08",X"1F",X"33",X"61",X"C0",X"C0",X"C7",X"C7",X"65",
		X"40",X"A8",X"50",X"AA",X"4F",X"AF",X"5F",X"BF",X"AE",X"AE",X"B2",X"A1",X"25",X"55",X"41",X"61",
		X"05",X"07",X"03",X"02",X"80",X"00",X"81",X"C1",X"61",X"C5",X"C7",X"C7",X"C0",X"61",X"33",X"1F",
		X"FF",X"77",X"73",X"62",X"02",X"02",X"A6",X"54",X"51",X"E3",X"92",X"66",X"CC",X"76",X"0F",X"FF",
		X"81",X"00",X"81",X"41",X"E0",X"FE",X"FF",X"FF",X"6F",X"F8",X"F6",X"F1",X"F0",X"78",X"3F",X"1F",
		X"A2",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"F0",X"00",
		X"FF",X"FF",X"FF",X"7F",X"1F",X"07",X"01",X"00",X"0F",X"07",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"72",X"02",X"52",X"AA",X"AA",X"FA",X"FA",X"FA",X"FA",X"FA",X"02",X"72",X"8A",X"8A",X"FA",X"FA",
		X"FA",X"FA",X"F2",X"02",X"FA",X"12",X"22",X"7A",X"BA",X"AA",X"EA",X"6A",X"02",X"F2",X"0A",X"0A",
		X"38",X"7C",X"C2",X"82",X"86",X"7C",X"38",X"00",X"02",X"02",X"FE",X"FE",X"42",X"02",X"00",X"00",
		X"62",X"F2",X"BA",X"9A",X"9E",X"4E",X"46",X"00",X"8C",X"DE",X"F2",X"B2",X"92",X"86",X"04",X"00",
		X"08",X"FE",X"FE",X"C8",X"68",X"38",X"18",X"00",X"1C",X"BE",X"B2",X"B2",X"B2",X"E6",X"E4",X"00",
		X"0C",X"9E",X"92",X"92",X"D2",X"7E",X"3C",X"00",X"C0",X"E0",X"B0",X"9E",X"8E",X"C0",X"C0",X"00",
		X"0C",X"6E",X"9A",X"9A",X"B2",X"F2",X"6C",X"00",X"78",X"FC",X"96",X"92",X"92",X"F2",X"60",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"00",X"00",X"FF",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"FF",X"00",X"00",X"00",
		X"FF",X"BE",X"BC",X"F8",X"E0",X"C0",X"C0",X"E0",X"03",X"01",X"01",X"03",X"07",X"0F",X"1F",X"3F",
		X"FF",X"FF",X"FF",X"FF",X"FE",X"F8",X"E0",X"C0",X"F3",X"E2",X"C4",X"07",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"0F",X"A8",X"E8",X"F9",X"FB",X"FF",X"FF",X"FF",X"FF",
		X"7E",X"FC",X"FE",X"FF",X"FF",X"FE",X"FF",X"FE",X"AA",X"AA",X"AA",X"AA",X"EA",X"FA",X"FE",X"FF",
		X"00",X"80",X"80",X"A0",X"A0",X"A0",X"A8",X"A8",X"01",X"01",X"03",X"07",X"0F",X"1F",X"1F",X"7F",
		X"80",X"80",X"80",X"A0",X"A0",X"A8",X"A8",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"20",X"A0",X"A0",X"A0",X"A0",X"00",X"00",X"7F",X"80",X"83",X"82",X"02",X"B2",
		X"A0",X"A0",X"A0",X"20",X"C0",X"00",X"00",X"00",X"02",X"82",X"83",X"80",X"7F",X"00",X"00",X"00",
		X"FF",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"FF",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"04",X"02",X"84",X"54",X"12",X"12",X"12",X"12",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"14",X"14",X"14",X"12",X"02",X"02",X"04",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"02",X"00",X"00",X"00",X"00",X"DE",X"2E",X"76",X"6A",
		X"02",X"02",X"02",X"01",X"00",X"00",X"00",X"00",X"6A",X"6A",X"76",X"2E",X"DE",X"00",X"00",X"00",
		X"07",X"0F",X"18",X"30",X"20",X"47",X"1E",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"02",
		X"FE",X"1E",X"47",X"20",X"30",X"18",X"0F",X"07",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"0F",X"1F",X"3F",X"3F",X"3F",X"3F",X"1F",X"0F",X"00",X"C0",X"E0",X"F0",X"F0",X"F8",X"FC",X"FE",
		X"1F",X"3F",X"3F",X"3F",X"3F",X"1F",X"0F",X"00",X"FC",X"F8",X"F0",X"F0",X"E0",X"C0",X"00",X"00",
		X"0F",X"1F",X"3F",X"3F",X"3F",X"3F",X"1D",X"08",X"00",X"C0",X"E0",X"F0",X"F0",X"F8",X"F4",X"E0",
		X"02",X"17",X"3F",X"3F",X"3F",X"3F",X"1F",X"0F",X"4A",X"1C",X"B8",X"F0",X"F0",X"E0",X"C0",X"00",
		X"03",X"07",X"0F",X"3C",X"3D",X"3E",X"3F",X"3D",X"38",X"BC",X"9C",X"CC",X"80",X"40",X"00",X"80",
		X"3D",X"3F",X"3E",X"3D",X"3C",X"0F",X"07",X"03",X"80",X"00",X"46",X"86",X"CE",X"8C",X"8C",X"00",
		X"00",X"00",X"07",X"0F",X"1F",X"5F",X"E6",X"ED",X"00",X"00",X"F0",X"F8",X"FC",X"FE",X"33",X"DF",
		X"7D",X"08",X"02",X"30",X"38",X"3C",X"3C",X"1C",X"DE",X"88",X"20",X"03",X"07",X"0F",X"0E",X"0C",
		X"BE",X"A6",X"82",X"82",X"82",X"82",X"A6",X"BE",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"86",X"FF",X"FF",X"3F",X"3F",X"FF",X"FF",X"8E",
		X"80",X"F7",X"F7",X"F4",X"F4",X"F7",X"F4",X"F4",X"01",X"DF",X"5F",X"5F",X"5F",X"DF",X"5F",X"5F",
		X"F7",X"F4",X"F5",X"F4",X"F7",X"FF",X"F7",X"80",X"DF",X"5F",X"5F",X"5F",X"DF",X"FF",X"DF",X"01",
		X"20",X"50",X"88",X"88",X"88",X"88",X"88",X"56",X"00",X"00",X"1F",X"7F",X"FF",X"7F",X"3F",X"2F",
		X"26",X"0C",X"0C",X"0C",X"0C",X"00",X"00",X"00",X"5E",X"0F",X"47",X"07",X"07",X"0F",X"07",X"03",
		X"07",X"08",X"08",X"08",X"07",X"00",X"07",X"08",X"C0",X"20",X"20",X"20",X"C0",X"00",X"C0",X"20",
		X"08",X"08",X"07",X"00",X"00",X"0F",X"04",X"00",X"20",X"20",X"C0",X"00",X"20",X"E0",X"20",X"00",
		X"FF",X"44",X"44",X"44",X"44",X"44",X"44",X"FF",X"7F",X"44",X"44",X"44",X"44",X"44",X"44",X"7F",
		X"BF",X"84",X"84",X"84",X"84",X"84",X"84",X"BF",X"DF",X"C4",X"44",X"44",X"44",X"44",X"44",X"DF",
		X"6F",X"E4",X"A4",X"24",X"24",X"24",X"A4",X"EF",X"37",X"74",X"D4",X"94",X"14",X"94",X"D4",X"77",
		X"1B",X"38",X"68",X"C8",X"88",X"C8",X"68",X"3B",X"0D",X"1C",X"34",X"64",X"44",X"64",X"34",X"1D",
		X"07",X"08",X"08",X"07",X"00",X"07",X"08",X"08",X"C0",X"20",X"20",X"C0",X"00",X"C0",X"20",X"20",
		X"07",X"00",X"06",X"09",X"08",X"08",X"04",X"00",X"C0",X"00",X"20",X"20",X"A0",X"60",X"20",X"00",
		X"07",X"08",X"08",X"07",X"00",X"07",X"08",X"08",X"C0",X"20",X"20",X"C0",X"00",X"C0",X"20",X"20",
		X"07",X"00",X"08",X"0D",X"0B",X"09",X"08",X"00",X"C0",X"00",X"C0",X"20",X"20",X"20",X"20",X"00",
		X"86",X"8E",X"9A",X"B2",X"A2",X"B2",X"9A",X"8E",X"C3",X"47",X"4D",X"59",X"51",X"59",X"4D",X"C7",
		X"E1",X"63",X"66",X"6C",X"68",X"6C",X"66",X"E3",X"F0",X"51",X"53",X"56",X"54",X"56",X"53",X"F1",
		X"F8",X"48",X"49",X"4B",X"4A",X"4B",X"49",X"F8",X"FC",X"44",X"44",X"45",X"45",X"45",X"44",X"FC",
		X"FE",X"46",X"46",X"46",X"46",X"46",X"46",X"FE",X"FF",X"45",X"45",X"45",X"45",X"45",X"45",X"FF",
		X"07",X"08",X"08",X"07",X"00",X"07",X"08",X"08",X"C0",X"20",X"20",X"C0",X"00",X"C0",X"20",X"20",
		X"07",X"00",X"09",X"0A",X"0A",X"0A",X"0E",X"00",X"C0",X"00",X"C0",X"20",X"20",X"20",X"40",X"00",
		X"07",X"08",X"08",X"07",X"00",X"07",X"08",X"08",X"C0",X"20",X"20",X"C0",X"00",X"C0",X"20",X"20",
		X"07",X"00",X"06",X"09",X"09",X"09",X"06",X"00",X"C0",X"00",X"C0",X"20",X"20",X"20",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"C0",X"C0",X"40",X"40",X"40",X"40",X"40",X"C0",
		X"60",X"E0",X"A0",X"20",X"20",X"20",X"A0",X"E0",X"30",X"70",X"D0",X"90",X"10",X"90",X"D0",X"70",
		X"18",X"38",X"68",X"C8",X"88",X"C8",X"68",X"38",X"0C",X"1C",X"34",X"64",X"44",X"64",X"34",X"1C",
		X"00",X"00",X"00",X"02",X"01",X"02",X"0A",X"08",X"60",X"70",X"70",X"70",X"70",X"F0",X"70",X"70",
		X"05",X"00",X"05",X"05",X"02",X"00",X"01",X"00",X"70",X"F0",X"70",X"70",X"F0",X"70",X"70",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"F0",X"00",X"F0",X"40",X"40",X"E0",X"E0",
		X"00",X"04",X"04",X"FC",X"F8",X"00",X"A8",X"A8",X"E0",X"F8",X"7D",X"01",X"70",X"88",X"FE",X"FE",
		X"86",X"8E",X"9A",X"B2",X"A2",X"B2",X"9A",X"8E",X"43",X"47",X"4D",X"59",X"51",X"59",X"4D",X"47",
		X"21",X"23",X"26",X"2C",X"28",X"2C",X"26",X"23",X"10",X"11",X"13",X"16",X"14",X"16",X"13",X"11",
		X"08",X"08",X"09",X"0B",X"0A",X"0B",X"09",X"08",X"04",X"04",X"04",X"05",X"05",X"05",X"04",X"04",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"42",X"24",X"00",X"00",X"24",X"42",X"00",X"26",X"6F",X"71",X"78",X"78",X"71",X"35",X"00",
		X"08",X"00",X"01",X"24",X"00",X"00",X"05",X"08",X"00",X"18",X"38",X"9F",X"37",X"25",X"09",X"5E",
		X"40",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"17",X"0E",X"10",X"21",X"0F",X"13",X"04",X"00",
		X"02",X"08",X"40",X"20",X"04",X"40",X"01",X"04",X"00",X"00",X"00",X"07",X"13",X"03",X"38",X"7F",
		X"08",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"02",X"43",X"07",X"06",X"10",X"00",
		X"80",X"10",X"08",X"04",X"06",X"03",X"10",X"2F",X"20",X"04",X"02",X"0B",X"37",X"FF",X"FF",X"FF",
		X"03",X"01",X"01",X"0A",X"05",X"00",X"00",X"20",X"FF",X"FF",X"FF",X"F9",X"13",X"21",X"42",X"00",
		X"01",X"40",X"00",X"00",X"02",X"01",X"00",X"00",X"00",X"00",X"03",X"03",X"7F",X"FF",X"7F",X"7F",
		X"01",X"03",X"06",X"00",X"10",X"01",X"00",X"10",X"FF",X"FF",X"7F",X"7F",X"8D",X"00",X"22",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"20",X"00",X"20",X"A3",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",
		X"20",X"20",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"02",X"02",X"02",X"02",X"02",X"02",X"03",
		X"07",X"04",X"04",X"04",X"04",X"04",X"04",X"07",X"0F",X"08",X"08",X"08",X"08",X"08",X"08",X"0F",
		X"1F",X"11",X"11",X"11",X"11",X"11",X"11",X"1F",X"3F",X"22",X"22",X"22",X"22",X"22",X"22",X"3F",
		X"7F",X"44",X"44",X"44",X"44",X"44",X"44",X"7F",X"FF",X"88",X"88",X"88",X"88",X"88",X"88",X"FF",
		X"18",X"24",X"62",X"51",X"85",X"46",X"24",X"18",X"18",X"24",X"46",X"89",X"91",X"62",X"24",X"18",
		X"18",X"2C",X"52",X"A9",X"D5",X"4A",X"34",X"18",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"FF",
		X"FF",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"40",X"C0",X"40",X"40",X"C0",X"40",X"40",X"FF",
		X"FF",X"40",X"40",X"C0",X"40",X"40",X"C0",X"40",X"20",X"E0",X"20",X"20",X"E0",X"20",X"20",X"FF",
		X"FF",X"20",X"20",X"E0",X"20",X"20",X"E0",X"20",X"10",X"F0",X"10",X"10",X"F0",X"10",X"10",X"FF",
		X"FF",X"10",X"10",X"F0",X"10",X"10",X"F0",X"10",X"08",X"F8",X"08",X"08",X"F8",X"08",X"08",X"FF",
		X"FF",X"08",X"08",X"F8",X"08",X"08",X"F8",X"08",X"04",X"FC",X"04",X"04",X"FC",X"04",X"04",X"FF",
		X"FF",X"04",X"04",X"FC",X"04",X"04",X"FC",X"04",X"02",X"FE",X"02",X"02",X"FE",X"02",X"02",X"FF",
		X"FF",X"02",X"02",X"FE",X"02",X"02",X"FE",X"02",X"81",X"FF",X"81",X"81",X"FF",X"81",X"81",X"FF",
		X"FF",X"81",X"81",X"FF",X"81",X"81",X"FF",X"81",X"40",X"7F",X"40",X"40",X"7F",X"40",X"40",X"FF",
		X"FF",X"40",X"40",X"7F",X"40",X"40",X"7F",X"40",X"20",X"3F",X"20",X"20",X"3F",X"20",X"20",X"FF",
		X"FF",X"20",X"20",X"3F",X"20",X"20",X"3F",X"20",X"10",X"1F",X"10",X"10",X"1F",X"10",X"10",X"FF",
		X"FF",X"10",X"10",X"1F",X"10",X"10",X"1F",X"10",X"08",X"0F",X"08",X"08",X"0F",X"08",X"08",X"FF",
		X"FF",X"08",X"08",X"0F",X"08",X"08",X"0F",X"08",X"04",X"07",X"04",X"04",X"07",X"04",X"04",X"FF",
		X"FF",X"04",X"04",X"07",X"04",X"04",X"07",X"04",X"02",X"03",X"02",X"02",X"03",X"02",X"02",X"FF",
		X"FF",X"02",X"02",X"03",X"02",X"02",X"03",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"FF",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"02",X"84",X"48",X"12",X"12",X"12",X"12",
		X"17",X"14",X"14",X"52",X"42",X"42",X"44",X"FF",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",
		X"FE",X"44",X"44",X"44",X"44",X"44",X"44",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"03",X"07",X"0E",X"1C",X"38",X"70",X"E0",X"C0",X"83",X"87",X"8E",X"9C",X"B8",X"F0",X"E0",X"C0",
		X"C0",X"E0",X"70",X"38",X"1C",X"0E",X"07",X"03",X"C0",X"E0",X"F0",X"B8",X"9C",X"8E",X"87",X"83",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"08",X"08",X"09",X"0B",X"0A",X"0B",X"09",X"08",X"60",X"E0",X"A0",X"20",X"20",X"20",X"A0",X"E0",
		X"08",X"08",X"09",X"0B",X"0A",X"0B",X"09",X"08",X"60",X"E0",X"A0",X"20",X"20",X"20",X"A0",X"E0",
		X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"80",X"80",X"A0",X"83",X"81",X"E1",X"D3",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"6F",X"0E",X"0E",X"1F",X"36",X"25",X"00",
		X"00",X"40",X"6C",X"6F",X"7F",X"FF",X"DF",X"DF",X"00",X"00",X"00",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"DF",X"9F",X"1F",X"0F",X"0F",X"07",X"06",X"04",X"C0",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",
		X"01",X"01",X"3B",X"7F",X"FF",X"BF",X"BF",X"BF",X"00",X"00",X"80",X"80",X"80",X"C0",X"C0",X"C0",
		X"BF",X"BF",X"DF",X"67",X"31",X"10",X"10",X"00",X"C0",X"C0",X"C0",X"C0",X"C0",X"40",X"00",X"00",
		X"10",X"10",X"3F",X"77",X"DF",X"BF",X"BF",X"BF",X"00",X"40",X"C0",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"BF",X"BF",X"FF",X"5F",X"77",X"3F",X"10",X"10",X"E0",X"E0",X"E0",X"E0",X"E0",X"C0",X"40",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"BE",X"A6",X"82",X"82",X"82",X"82",X"A6",X"BE",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"86",X"FF",X"FF",X"3F",X"3F",X"FF",X"FF",X"8E",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"44",X"44",X"44",X"44",X"44",X"44",X"FF",X"7F",X"44",X"44",X"44",X"44",X"44",X"44",X"7F",
		X"BF",X"84",X"84",X"84",X"84",X"84",X"84",X"BF",X"DF",X"C4",X"44",X"44",X"44",X"44",X"44",X"DF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"04",X"1C",X"65",X"E1",X"F9",X"E9",X"00",X"00",X"00",X"FF",X"FF",X"E7",X"E5",X"E8",
		X"C1",X"55",X"4C",X"44",X"04",X"00",X"00",X"00",X"BF",X"FF",X"FF",X"39",X"00",X"00",X"00",X"00",
		X"00",X"00",X"05",X"1D",X"65",X"E1",X"F9",X"D9",X"00",X"06",X"8F",X"9F",X"FD",X"FC",X"F8",X"B8",
		X"C1",X"55",X"4C",X"44",X"04",X"00",X"00",X"00",X"F8",X"FC",X"FC",X"BC",X"5C",X"3C",X"00",X"00",
		X"00",X"00",X"00",X"02",X"0E",X"32",X"70",X"7C",X"1E",X"1C",X"1C",X"1C",X"FC",X"FC",X"F8",X"FB",
		X"74",X"60",X"2A",X"26",X"22",X"02",X"00",X"00",X"FF",X"FF",X"1D",X"18",X"00",X"00",X"00",X"00",
		X"00",X"03",X"07",X"07",X"1F",X"7B",X"7B",X"7B",X"00",X"00",X"00",X"F0",X"FE",X"FF",X"FF",X"FF",
		X"7B",X"7B",X"7B",X"3F",X"3F",X"1C",X"00",X"00",X"F7",X"FB",X"F8",X"F8",X"F8",X"60",X"00",X"00",
		X"00",X"07",X"1F",X"3F",X"3F",X"3F",X"3F",X"3F",X"00",X"80",X"C0",X"F0",X"FE",X"FF",X"FF",X"BF",
		X"3F",X"7F",X"7F",X"3F",X"1F",X"03",X"00",X"00",X"FF",X"F3",X"F0",X"E0",X"80",X"00",X"00",X"00",
		X"00",X"03",X"07",X"07",X"0F",X"1F",X"1F",X"1F",X"80",X"80",X"F0",X"F8",X"FC",X"FE",X"FE",X"DE",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"0F",X"07",X"03",X"44",X"C0",X"C0",X"C0",X"80",X"80",X"00",X"00",
		X"00",X"00",X"01",X"03",X"1B",X"7B",X"7B",X"7B",X"00",X"C0",X"C0",X"FD",X"FF",X"FF",X"FF",X"FB",
		X"7B",X"7B",X"7B",X"1B",X"03",X"01",X"00",X"00",X"FB",X"FF",X"FF",X"FF",X"FD",X"C0",X"C0",X"00",
		X"00",X"00",X"00",X"FF",X"44",X"44",X"44",X"44",X"00",X"00",X"00",X"FF",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"FF",X"00",X"00",X"00",X"44",X"44",X"44",X"44",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"04",X"1C",X"65",X"E3",X"1F",X"1F",X"00",X"00",X"00",X"1F",X"FF",X"FF",X"FD",X"F8",
		X"1F",X"55",X"4C",X"44",X"04",X"00",X"00",X"00",X"BF",X"FF",X"FF",X"39",X"00",X"00",X"00",X"00",
		X"00",X"00",X"04",X"1C",X"65",X"E1",X"F9",X"E9",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FD",X"F8",
		X"C1",X"55",X"4C",X"44",X"04",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"F9",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"04",X"1C",X"65",X"E7",X"1F",X"1F",X"00",X"06",X"0F",X"1F",X"FD",X"FC",X"F8",X"F8",
		X"1F",X"55",X"4C",X"44",X"04",X"00",X"00",X"00",X"B8",X"FC",X"7C",X"1C",X"1C",X"3C",X"00",X"00",
		X"00",X"00",X"04",X"1C",X"64",X"E1",X"F9",X"E9",X"00",X"06",X"0F",X"1F",X"FD",X"FC",X"F8",X"F8",
		X"C1",X"55",X"4C",X"44",X"04",X"00",X"00",X"00",X"F8",X"FC",X"FC",X"DC",X"1C",X"1C",X"00",X"00",
		X"00",X"00",X"00",X"02",X"0E",X"32",X"71",X"1F",X"1E",X"1C",X"1C",X"1C",X"FC",X"FC",X"F8",X"FB",
		X"1F",X"1F",X"2A",X"26",X"22",X"02",X"00",X"00",X"FF",X"DF",X"FD",X"38",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"02",X"0E",X"32",X"70",X"7C",X"1E",X"1C",X"1C",X"1C",X"FC",X"FC",X"F8",X"FB",
		X"74",X"60",X"2A",X"26",X"22",X"02",X"00",X"00",X"FF",X"FF",X"FD",X"78",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"02",X"0E",X"32",X"70",X"7C",X"04",X"0C",X"18",X"9C",X"CE",X"FF",X"FF",X"FE",
		X"74",X"60",X"2A",X"26",X"22",X"02",X"00",X"00",X"DC",X"FC",X"FC",X"7C",X"4C",X"CC",X"4C",X"1C",
		X"01",X"03",X"07",X"1F",X"65",X"E1",X"F9",X"E9",X"80",X"80",X"00",X"F8",X"FC",X"FE",X"FE",X"BF",
		X"C1",X"55",X"4D",X"45",X"05",X"01",X"00",X"00",X"FF",X"FF",X"FE",X"9F",X"0F",X"06",X"0C",X"00",
		X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"80",X"80",X"A0",X"83",X"81",X"E1",X"D3",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"6F",X"0E",X"0E",X"1F",X"36",X"25",X"00",
		X"00",X"40",X"6C",X"6F",X"7F",X"FF",X"DF",X"DF",X"00",X"00",X"00",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"DF",X"9F",X"1F",X"0F",X"0F",X"07",X"06",X"04",X"C0",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",
		X"01",X"01",X"3B",X"7F",X"FF",X"BF",X"BF",X"BF",X"00",X"00",X"80",X"80",X"80",X"C0",X"C0",X"C0",
		X"BF",X"BF",X"DF",X"67",X"31",X"10",X"10",X"00",X"C0",X"C0",X"C0",X"C0",X"C0",X"40",X"00",X"00",
		X"10",X"10",X"3F",X"77",X"DF",X"BF",X"BF",X"BF",X"00",X"40",X"C0",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"BF",X"BF",X"FF",X"5F",X"77",X"3F",X"10",X"10",X"E0",X"E0",X"E0",X"E0",X"E0",X"C0",X"40",X"00",
		X"00",X"01",X"07",X"0F",X"1F",X"1F",X"1F",X"1F",X"60",X"E0",X"E0",X"E0",X"F0",X"E0",X"C0",X"C0",
		X"1F",X"1F",X"1F",X"0F",X"06",X"06",X"03",X"01",X"E0",X"E0",X"C0",X"00",X"00",X"00",X"80",X"80",
		X"00",X"00",X"03",X"07",X"0F",X"0D",X"1E",X"1F",X"00",X"00",X"C0",X"E0",X"F0",X"F0",X"F8",X"78",
		X"1F",X"19",X"09",X"0F",X"07",X"03",X"00",X"00",X"B8",X"F8",X"F0",X"F0",X"E0",X"C0",X"00",X"00",
		X"07",X"00",X"0F",X"1F",X"1F",X"1F",X"1F",X"1F",X"E0",X"00",X"F0",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"0F",X"00",X"07",X"F8",X"F8",X"F8",X"F8",X"F8",X"F0",X"00",X"E0",
		X"07",X"00",X"0F",X"1F",X"1F",X"1F",X"1F",X"1F",X"E0",X"00",X"F0",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"0F",X"00",X"07",X"F8",X"F8",X"F8",X"F8",X"F8",X"F0",X"00",X"E0",
		X"00",X"00",X"00",X"1F",X"3F",X"BF",X"BF",X"BF",X"00",X"00",X"00",X"F8",X"FC",X"FD",X"FD",X"FD",
		X"BF",X"BF",X"BF",X"3F",X"1F",X"00",X"00",X"00",X"FD",X"FD",X"FD",X"FC",X"F8",X"00",X"00",X"00",
		X"00",X"00",X"03",X"07",X"0F",X"0C",X"1B",X"1A",X"00",X"00",X"C0",X"E0",X"70",X"B0",X"58",X"B8",
		X"19",X"18",X"0C",X"0F",X"07",X"03",X"00",X"00",X"B8",X"38",X"70",X"F0",X"E0",X"C0",X"00",X"00",
		X"07",X"00",X"0F",X"1F",X"1F",X"1F",X"1F",X"1F",X"E0",X"00",X"F0",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"0F",X"00",X"07",X"F8",X"F8",X"F8",X"F8",X"F8",X"F0",X"00",X"E0",
		X"07",X"00",X"0F",X"1F",X"1F",X"1F",X"1F",X"1F",X"E0",X"00",X"F0",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"0F",X"00",X"07",X"F8",X"F8",X"F8",X"F8",X"F8",X"F0",X"00",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"80",X"00",X"80",X"8F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"42",X"48",X"44",X"42",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"78",X"02",X"42",X"0A",X"14",X"02",
		X"00",X"1E",X"3F",X"3F",X"3F",X"7D",X"7F",X"3E",X"CC",X"E6",X"EF",X"C3",X"E7",X"E7",X"E7",X"C3",
		X"1E",X"3F",X"7D",X"3F",X"1F",X"0C",X"00",X"0F",X"F7",X"F7",X"E7",X"C3",X"E7",X"F6",X"E6",X"FC",
		X"00",X"1E",X"3F",X"3F",X"3F",X"6F",X"7F",X"3E",X"CC",X"E6",X"EF",X"C3",X"E7",X"E7",X"E7",X"C3",
		X"1E",X"3F",X"7F",X"3F",X"1B",X"0C",X"00",X"0F",X"F7",X"F7",X"E7",X"C3",X"E7",X"F6",X"E6",X"FC",
		X"00",X"1E",X"3B",X"3F",X"3F",X"7F",X"7F",X"3E",X"CC",X"E6",X"EF",X"C3",X"E7",X"E7",X"E7",X"C3",
		X"1E",X"3F",X"77",X"3F",X"1F",X"0C",X"00",X"0F",X"F7",X"F7",X"E7",X"C3",X"E7",X"F6",X"E6",X"FC",
		X"0F",X"01",X"09",X"1F",X"3F",X"3F",X"1A",X"0E",X"E0",X"D8",X"B8",X"BC",X"BC",X"BC",X"BC",X"BC",
		X"1A",X"3F",X"3F",X"1F",X"09",X"01",X"01",X"0F",X"BC",X"BC",X"BC",X"BC",X"B8",X"D8",X"E0",X"E0",
		X"0F",X"01",X"09",X"1F",X"3F",X"3F",X"1A",X"0E",X"D0",X"F8",X"D8",X"8C",X"DC",X"FC",X"DC",X"8C",
		X"1A",X"3F",X"3F",X"1F",X"09",X"01",X"01",X"0F",X"DC",X"FC",X"DC",X"8C",X"D8",X"F8",X"D8",X"F0",
		X"38",X"FC",X"FF",X"EF",X"FF",X"FF",X"FF",X"7F",X"00",X"00",X"40",X"80",X"80",X"C0",X"00",X"80",
		X"7F",X"FF",X"FF",X"FF",X"EF",X"FF",X"FC",X"38",X"C0",X"80",X"C0",X"80",X"80",X"40",X"00",X"00",
		X"00",X"00",X"09",X"00",X"00",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"04",X"04",X"04",
		X"08",X"04",X"04",X"03",X"00",X"00",X"00",X"00",X"04",X"08",X"0C",X"0C",X"14",X"1C",X"1C",X"0C",
		X"00",X"00",X"00",X"00",X"01",X"02",X"04",X"08",X"01",X"03",X"07",X"E3",X"07",X"05",X"03",X"03",
		X"00",X"00",X"48",X"B4",X"00",X"00",X"00",X"00",X"03",X"07",X"05",X"03",X"06",X"00",X"00",X"00",
		X"00",X"00",X"38",X"3C",X"7C",X"7F",X"FF",X"FC",X"00",X"00",X"00",X"00",X"40",X"80",X"00",X"00",
		X"FC",X"FC",X"78",X"20",X"00",X"00",X"06",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"EE",X"60",X"00",X"0E",X"1A",X"1D",X"18",X"00",X"10",X"30",X"30",
		X"10",X"08",X"08",X"04",X"02",X"02",X"01",X"00",X"60",X"40",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"3C",X"60",X"C0",
		X"01",X"03",X"06",X"04",X"04",X"01",X"06",X"0E",X"80",X"00",X"00",X"00",X"00",X"01",X"03",X"E0",
		X"00",X"00",X"00",X"00",X"C0",X"78",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"17",X"E7",X"87",X"06",X"06",X"00",X"40",X"E0",X"70",X"B0",X"F8",X"18",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"78",X"FE",X"33",
		X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"40",X"07",X"81",X"83",X"03",X"03",X"01",X"00",X"00",
		X"0F",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"03",X"03",X"05",X"07",X"07",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0E",X"5E",X"FF",X"FF",X"CF",X"C6",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"E0",X"E0",
		X"01",X"01",X"03",X"03",X"87",X"C7",X"7F",X"3F",X"E0",X"E0",X"C0",X"C1",X"83",X"87",X"07",X"03",
		X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"04",X"00",X"01",X"07",X"3C",X"C0",X"00",X"00",X"00",
		X"04",X"08",X"09",X"09",X"08",X"10",X"10",X"10",X"00",X"00",X"FC",X"07",X"01",X"00",X"00",X"00",
		X"03",X"07",X"07",X"03",X"08",X"1C",X"1E",X"3F",X"00",X"00",X"C0",X"60",X"30",X"1C",X"3E",X"7E",
		X"3F",X"3B",X"1F",X"03",X"03",X"03",X"01",X"00",X"F6",X"EE",X"DC",X"DC",X"DC",X"D8",X"D0",X"60",
		X"00",X"00",X"01",X"01",X"02",X"02",X"02",X"04",X"40",X"80",X"00",X"00",X"00",X"42",X"33",X"07",
		X"04",X"04",X"08",X"08",X"08",X"08",X"08",X"08",X"07",X"07",X"07",X"07",X"00",X"00",X"00",X"00",
		X"00",X"80",X"C0",X"40",X"61",X"3A",X"0E",X"07",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"0A",X"32",X"41",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",
		X"60",X"F0",X"A0",X"80",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"60",X"20",X"20",
		X"00",X"08",X"08",X"04",X"0E",X"08",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"0C",X"06",X"06",X"06",X"04",X"08",X"10",X"00",X"00",X"0C",X"0E",X"0F",X"0F",X"0F",X"07",
		X"20",X"00",X"80",X"60",X"18",X"0C",X"00",X"00",X"07",X"03",X"03",X"01",X"00",X"00",X"00",X"00",
		X"00",X"18",X"20",X"40",X"80",X"00",X"00",X"21",X"00",X"00",X"10",X"70",X"70",X"F0",X"F0",X"F0",
		X"11",X"09",X"04",X"04",X"06",X"06",X"06",X"06",X"F0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"01",X"03",X"06",X"0C",X"15",X"00",X"00",X"80",X"40",X"E0",X"30",X"18",X"54",
		X"15",X"0C",X"06",X"03",X"01",X"00",X"00",X"00",X"54",X"18",X"30",X"E0",X"40",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"20",X"50",X"70",X"50",X"D8",X"88",X"88",X"04",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"88",X"88",X"D8",X"50",X"70",X"50",X"20",
		X"00",X"44",X"02",X"01",X"05",X"43",X"0F",X"16",X"00",X"00",X"00",X"78",X"FE",X"86",X"03",X"73",
		X"03",X"0E",X"5B",X"21",X"00",X"00",X"00",X"00",X"7B",X"3B",X"33",X"86",X"FE",X"3C",X"00",X"00",
		X"00",X"00",X"28",X"87",X"33",X"1E",X"0C",X"44",X"00",X"80",X"78",X"FC",X"86",X"03",X"71",X"F9",
		X"32",X"1E",X"0D",X"03",X"01",X"00",X"00",X"00",X"F9",X"79",X"7B",X"32",X"86",X"FC",X"38",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"30",X"30",X"30",X"30",X"00",X"00",X"00",X"00",X"C0",X"C0",X"C0",X"C0",
		X"30",X"30",X"3F",X"3F",X"00",X"00",X"00",X"00",X"C0",X"C0",X"FC",X"FC",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"3F",X"3F",X"30",X"30",X"00",X"00",X"00",X"00",X"FC",X"FC",X"C0",X"C0",
		X"30",X"30",X"3F",X"3F",X"00",X"00",X"00",X"00",X"C0",X"C0",X"FC",X"FC",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0C",X"0C",X"0C",
		X"00",X"00",X"3F",X"3F",X"00",X"00",X"00",X"00",X"0C",X"0C",X"FC",X"FC",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"3C",X"3C",X"30",X"30",X"00",X"00",X"00",X"00",X"3C",X"3C",X"0C",X"0C",
		X"30",X"30",X"3F",X"3F",X"00",X"00",X"00",X"00",X"0C",X"0C",X"FC",X"FC",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"3F",X"3F",X"30",X"30",X"00",X"00",X"00",X"00",X"FC",X"FC",X"0C",X"0C",
		X"30",X"30",X"3F",X"3F",X"00",X"00",X"00",X"00",X"0C",X"0C",X"FC",X"FC",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"3F",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"FC",X"30",X"C0",
		X"03",X"0C",X"3F",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"FC",X"00",X"00",X"00",X"00",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"FF",X"FF",X"03",X"03",X"03",X"03",X"03",X"03",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"03",X"1F",X"FC",
		X"00",X"00",X"01",X"0F",X"7E",X"F0",X"80",X"00",X"0F",X"3F",X"FB",X"C3",X"03",X"03",X"03",X"03",
		X"00",X"00",X"00",X"00",X"00",X"03",X"1F",X"FC",X"00",X"00",X"01",X"0F",X"7E",X"F0",X"80",X"00",
		X"07",X"3F",X"F8",X"C0",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C3",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"FF",X"F0",X"00",X"00",X"00",X"00",X"3F",X"FF",X"C0",X"00",
		X"00",X"00",X"03",X"FF",X"FC",X"00",X"00",X"00",X"00",X"0F",X"FF",X"F0",X"00",X"00",X"00",X"00",
		X"3F",X"FF",X"C3",X"03",X"03",X"03",X"03",X"03",X"FC",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"FC",X"FF",X"C3",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"F0",X"FF",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"FF",X"3F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FC",X"FF",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"FF",X"0F",X"00",
		X"03",X"03",X"03",X"03",X"03",X"C3",X"FF",X"3F",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"E0",
		X"FC",X"1F",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"F0",X"7E",X"0F",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"F8",X"3F",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",
		X"FC",X"1F",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"F0",X"7E",X"0F",X"01",X"00",X"00",
		X"03",X"03",X"03",X"03",X"C3",X"FD",X"3F",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"03",X"03",X"03",X"03",X"03",X"03",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"03",X"03",X"03",X"03",X"03",X"03",X"FF",X"FF",
		X"C0",X"C0",X"FF",X"FF",X"C0",X"C0",X"C0",X"C0",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"03",X"03",X"03",X"03",X"FF",X"FF",X"03",X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
