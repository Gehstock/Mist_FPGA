library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity fg_sp_graphx_3 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of fg_sp_graphx_3 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"7C",X"C2",X"82",X"86",X"7C",X"38",
		X"00",X"00",X"80",X"84",X"FE",X"FE",X"80",X"80",X"00",X"C4",X"E6",X"F2",X"B2",X"BA",X"9E",X"8C",
		X"00",X"40",X"C2",X"92",X"9A",X"9E",X"F6",X"62",X"00",X"30",X"38",X"2C",X"26",X"FE",X"FE",X"20",
		X"00",X"4E",X"CE",X"8A",X"8A",X"8A",X"FA",X"70",X"00",X"78",X"FC",X"96",X"92",X"92",X"F2",X"60",
		X"00",X"06",X"06",X"E2",X"F2",X"1A",X"0E",X"06",X"00",X"6C",X"9E",X"9A",X"B2",X"B2",X"EC",X"60",
		X"00",X"0C",X"9E",X"92",X"92",X"D2",X"7E",X"3C",X"00",X"00",X"00",X"00",X"00",X"16",X"0E",X"00",
		X"00",X"10",X"10",X"10",X"10",X"10",X"00",X"00",X"00",X"F8",X"FC",X"26",X"22",X"26",X"FC",X"F8",
		X"00",X"FE",X"FE",X"92",X"92",X"92",X"FE",X"6C",X"00",X"38",X"7C",X"C6",X"82",X"82",X"C6",X"44",
		X"00",X"FE",X"FE",X"82",X"82",X"C6",X"7C",X"38",X"00",X"00",X"FE",X"FE",X"92",X"92",X"92",X"82",
		X"00",X"FE",X"FE",X"12",X"12",X"12",X"12",X"02",X"00",X"38",X"7C",X"C6",X"82",X"92",X"F2",X"F2",
		X"00",X"FE",X"FE",X"10",X"10",X"10",X"FE",X"FE",X"00",X"00",X"82",X"82",X"FE",X"FE",X"82",X"82",
		X"00",X"40",X"C0",X"80",X"80",X"80",X"FE",X"7E",X"00",X"FE",X"FE",X"30",X"78",X"EC",X"C6",X"82",
		X"00",X"00",X"FE",X"FE",X"80",X"80",X"80",X"80",X"00",X"FE",X"FE",X"1C",X"38",X"1C",X"FE",X"FE",
		X"00",X"FE",X"FE",X"1C",X"38",X"70",X"FE",X"FE",X"00",X"7C",X"FE",X"82",X"82",X"82",X"FE",X"7C",
		X"00",X"FE",X"FE",X"22",X"22",X"22",X"3E",X"1C",X"00",X"7C",X"FE",X"82",X"A2",X"E2",X"7E",X"BC",
		X"00",X"FE",X"FE",X"22",X"62",X"F2",X"DE",X"9C",X"00",X"4C",X"DE",X"92",X"92",X"96",X"F4",X"60",
		X"00",X"00",X"02",X"02",X"FE",X"FE",X"02",X"02",X"00",X"7E",X"FE",X"80",X"80",X"80",X"FE",X"7E",
		X"00",X"1E",X"3E",X"70",X"E0",X"70",X"3E",X"1E",X"00",X"3E",X"FE",X"70",X"38",X"70",X"FE",X"3E",
		X"00",X"C6",X"EE",X"7C",X"38",X"7C",X"EE",X"C6",X"00",X"00",X"06",X"1E",X"F0",X"F0",X"1E",X"06",
		X"00",X"C2",X"E2",X"F2",X"BA",X"9E",X"8E",X"86",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7E",X"81",X"BD",X"BD",X"A5",X"A5",X"81",X"7E",
		X"00",X"FF",X"FF",X"C3",X"C3",X"E7",X"7E",X"7E",X"FF",X"DB",X"DB",X"DB",X"7E",X"FF",X"C3",X"C3",
		X"F7",X"76",X"7E",X"FF",X"C3",X"C3",X"FF",X"7E",X"00",X"76",X"81",X"81",X"81",X"81",X"81",X"76",
		X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"00",X"70",X"89",X"89",X"89",X"89",X"89",X"06",
		X"00",X"00",X"81",X"89",X"89",X"89",X"89",X"76",X"00",X"06",X"08",X"08",X"08",X"08",X"F7",X"00",
		X"00",X"06",X"89",X"89",X"89",X"89",X"89",X"70",X"00",X"76",X"89",X"89",X"89",X"89",X"89",X"70",
		X"00",X"06",X"01",X"01",X"01",X"01",X"01",X"76",X"00",X"76",X"89",X"89",X"89",X"89",X"89",X"76",
		X"00",X"06",X"89",X"89",X"89",X"89",X"89",X"76",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"1F",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"1F",X"00",X"00",X"00",
		X"00",X"00",X"00",X"F8",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"F8",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"00",X"00",X"00",X"66",X"66",X"00",X"00",X"00",X"00",X"00",X"50",X"30",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"70",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"42",X"20",X"E8",X"E0",X"D8",X"78",X"FC",X"D8",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"C0",X"D2",X"65",X"E6",X"43",X"7F",X"1D",X"3B",X"7E",X"24",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"84",X"40",X"D0",X"C0",X"B0",X"F0",X"F8",X"B0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"08",X"80",X"A4",X"CA",X"CD",X"87",X"FF",X"3A",X"77",X"FD",X"48",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"08",X"80",X"A0",X"80",X"60",X"E0",X"F0",X"60",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"49",X"94",X"9B",X"0F",X"FF",X"75",X"EF",X"FB",X"90",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"01",X"03",X"01",X"01",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"10",X"00",X"40",X"00",X"C0",X"C0",X"E0",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"92",X"29",X"37",X"1F",X"FE",X"EB",X"DF",X"F6",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"03",X"07",X"02",X"03",X"00",X"01",X"03",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"80",X"00",X"80",X"80",X"C0",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"40",X"01",X"24",X"52",X"6E",X"3E",X"FD",X"D7",X"BF",X"ED",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0D",X"06",X"0E",X"04",X"07",X"01",X"03",X"07",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"02",X"48",X"A4",X"DD",X"7C",X"FB",X"AF",X"7F",X"DB",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"1A",X"0C",X"1C",X"08",X"0F",X"03",X"07",X"0F",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"90",X"48",X"BA",X"F8",X"F6",X"5E",X"FF",X"B6",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"30",X"34",X"19",X"39",X"10",X"1F",X"07",X"0E",X"1F",X"09",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"21",X"90",X"74",X"F0",X"EC",X"BC",X"FE",X"6C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"60",X"69",X"32",X"73",X"21",X"3F",X"0E",X"1D",X"3F",X"12",
		X"08",X"1C",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7C",X"44",X"30",X"00",
		X"00",X"1C",X"06",X"0E",X"00",X"00",X"0F",X"1C",X"1C",X"0C",X"0F",X"40",X"18",X"70",X"44",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"20",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"10",X"60",X"40",X"38",X"00",X"3C",X"70",
		X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"21",X"00",X"04",X"00",X"00",X"00",X"18",X"77",X"01",
		X"70",X"3C",X"00",X"38",X"40",X"60",X"10",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"47",X"08",X"00",X"00",X"00",X"04",X"00",X"20",X"00",X"00",X"04",X"00",X"00",X"00",X"00",
		X"C0",X"80",X"00",X"80",X"80",X"00",X"80",X"C0",X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"00",
		X"01",X"03",X"02",X"07",X"02",X"05",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"C0",X"80",X"00",X"80",X"80",X"00",X"80",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"05",X"02",X"07",X"02",X"03",X"01",
		X"00",X"00",X"00",X"00",X"70",X"80",X"70",X"A0",X"C0",X"40",X"3E",X"0C",X"18",X"10",X"34",X"F6",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"02",X"02",X"02",X"02",
		X"F6",X"34",X"10",X"18",X"0C",X"3E",X"80",X"C0",X"D0",X"80",X"A0",X"70",X"00",X"00",X"00",X"00",
		X"02",X"02",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"40",X"80",X"80",X"40",X"00",X"E0",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"03",X"07",
		X"03",X"02",X"0D",X"05",X"01",X"0C",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"03",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"E0",X"00",X"40",X"80",X"80",X"40",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"0C",X"01",X"05",X"0D",X"02",X"03",
		X"00",X"C0",X"00",X"80",X"50",X"40",X"00",X"00",X"80",X"00",X"00",X"00",X"80",X"C2",X"FF",X"FB",
		X"00",X"07",X"04",X"09",X"0F",X"14",X"0F",X"38",X"3F",X"1C",X"0E",X"07",X"03",X"03",X"07",X"07",
		X"FB",X"FF",X"C2",X"80",X"00",X"00",X"00",X"80",X"80",X"80",X"00",X"80",X"00",X"00",X"C0",X"00",
		X"07",X"07",X"03",X"03",X"07",X"0E",X"1C",X"3F",X"35",X"08",X"02",X"15",X"0A",X"04",X"07",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"1F",X"02",X"2A",X"10",X"1A",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"1A",X"10",X"2A",X"02",X"1F",X"00",X"00",X"00",X"00",
		X"00",X"80",X"00",X"00",X"80",X"00",X"00",X"00",X"9C",X"38",X"70",X"E0",X"C0",X"84",X"FE",X"F6",
		X"00",X"0F",X"04",X"12",X"34",X"08",X"3E",X"2A",X"0F",X"00",X"00",X"00",X"01",X"01",X"03",X"03",
		X"F6",X"FE",X"84",X"C0",X"E0",X"70",X"38",X"9C",X"00",X"00",X"00",X"80",X"00",X"00",X"80",X"00",
		X"03",X"03",X"01",X"01",X"00",X"00",X"00",X"0F",X"2A",X"3E",X"08",X"34",X"12",X"04",X"0F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"50",X"60",X"50",X"38",X"00",X"00",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"00",X"00",X"38",X"50",X"60",X"50",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"04",X"00",X"78",X"82",X"34",X"D1",X"E0",X"70",X"00",X"00",X"1E",X"30",X"F6",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F6",X"30",X"1E",X"00",X"00",X"70",X"80",X"51",X"84",X"A0",X"70",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"1C",X"14",X"6A",X"20",X"5A",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"40",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"5A",X"20",X"6A",X"14",X"1C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"30",X"10",X"1C",X"00",X"00",X"1E",X"38",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",
		X"38",X"1E",X"00",X"00",X"1C",X"30",X"28",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"00",X"00",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"00",X"00",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"10",X"20",X"1C",X"00",X"00",X"1E",X"38",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"38",X"1E",X"00",X"00",X"1C",X"20",X"10",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"02",X"06",X"00",X"F8",X"03",X"03",X"03",X"78",X"78",X"00",X"F8",X"00",X"1E",X"10",X"1C",
		X"0E",X"1E",X"02",X"00",X"7F",X"7F",X"3F",X"33",X"3F",X"3F",X"7F",X"7F",X"00",X"60",X"70",X"40",
		X"2C",X"60",X"74",X"68",X"38",X"30",X"00",X"FC",X"FC",X"00",X"2C",X"36",X"0E",X"1E",X"24",X"00",
		X"00",X"58",X"3C",X"18",X"10",X"30",X"00",X"7F",X"7F",X"00",X"60",X"60",X"E0",X"E8",X"F0",X"68",
		X"00",X"0C",X"06",X"00",X"00",X"0E",X"1C",X"00",X"00",X"00",X"00",X"00",X"22",X"1A",X"14",X"00",
		X"00",X"28",X"34",X"1C",X"14",X"00",X"18",X"20",X"20",X"18",X"00",X"00",X"C0",X"E8",X"F0",X"68",
		X"70",X"7E",X"62",X"00",X"00",X"70",X"40",X"FC",X"FC",X"70",X"00",X"00",X"00",X"06",X"16",X"0E",
		X"60",X"26",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"62",X"06",
		X"08",X"10",X"00",X"00",X"00",X"78",X"C8",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"21",X"42",X"00",X"00",X"00",X"01",X"12",X"05",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"84",X"C4",X"FC",X"F0",X"D0",X"90",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"1F",X"7F",X"7B",X"77",X"77",X"7B",X"7F",X"1F",X"00",X"00",X"00",X"00",
		X"60",X"20",X"60",X"E0",X"20",X"E0",X"80",X"80",X"80",X"80",X"E0",X"20",X"E0",X"00",X"00",X"00",
		X"00",X"80",X"80",X"31",X"3F",X"37",X"27",X"07",X"3F",X"3F",X"3F",X"3F",X"31",X"11",X"00",X"11",
		X"00",X"F0",X"F0",X"68",X"28",X"3F",X"1F",X"BF",X"9F",X"DF",X"BF",X"62",X"62",X"F0",X"F0",X"00",
		X"00",X"7F",X"FD",X"F8",X"C0",X"D8",X"B0",X"B6",X"BD",X"EE",X"FF",X"F3",X"FE",X"FF",X"7F",X"00",
		X"80",X"80",X"00",X"08",X"08",X"0F",X"1F",X"1F",X"1F",X"1F",X"0F",X"02",X"02",X"00",X"00",X"80",
		X"00",X"7F",X"FF",X"FB",X"2B",X"DB",X"33",X"37",X"BF",X"6F",X"7F",X"33",X"F7",X"F7",X"7F",X"00",
		X"80",X"C0",X"00",X"08",X"08",X"0F",X"1F",X"1F",X"1F",X"1F",X"0F",X"02",X"02",X"00",X"C0",X"80",
		X"01",X"78",X"F8",X"F8",X"38",X"F8",X"38",X"3E",X"BE",X"78",X"78",X"38",X"F8",X"F8",X"78",X"01",
		X"80",X"C0",X"00",X"08",X"08",X"0F",X"FF",X"1F",X"1F",X"FF",X"0F",X"02",X"02",X"00",X"C0",X"80",
		X"01",X"F0",X"F0",X"F8",X"F8",X"F8",X"FF",X"FE",X"FE",X"FF",X"F8",X"F8",X"F8",X"F0",X"F0",X"01",
		X"00",X"20",X"60",X"50",X"50",X"10",X"78",X"C8",X"C8",X"78",X"88",X"0C",X"0C",X"0C",X"08",X"00",
		X"00",X"08",X"0C",X"1C",X"1C",X"3C",X"78",X"10",X"16",X"7B",X"3D",X"48",X"48",X"60",X"20",X"00",
		X"14",X"14",X"00",X"30",X"60",X"F8",X"1C",X"1E",X"1E",X"1C",X"F8",X"60",X"30",X"00",X"08",X"08",
		X"00",X"00",X"04",X"0C",X"00",X"3F",X"20",X"20",X"20",X"20",X"3F",X"00",X"00",X"20",X"20",X"00",
		X"00",X"00",X"00",X"08",X"80",X"40",X"90",X"40",X"00",X"00",X"80",X"00",X"00",X"00",X"10",X"00",
		X"00",X"00",X"00",X"20",X"00",X"30",X"02",X"08",X"02",X"13",X"08",X"14",X"02",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"10",X"20",X"10",X"08",X"10",X"28",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"2E",X"32",X"20",X"00",
		X"00",X"00",X"00",X"00",X"90",X"80",X"C0",X"00",X"10",X"00",X"20",X"30",X"70",X"28",X"40",X"00",
		X"00",X"00",X"00",X"00",X"07",X"1F",X"1F",X"0E",X"0E",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"F8",X"DC",X"EC",X"7E",X"77",X"F8",X"D4",X"B8",X"F8",X"E0",X"C0",X"00",X"00",
		X"00",X"00",X"04",X"0E",X"1B",X"18",X"35",X"3F",X"1F",X"1F",X"3F",X"7F",X"0F",X"1C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"08",X"40",X"E0",X"51",X"A1",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E1",X"B3",X"84",X"08",X"08",X"00",X"48",X"2C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"03",X"05",X"0D",X"27",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"09",X"03",X"91",X"40",X"84",X"12",X"2C",X"28",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"80",X"C8",X"70",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"2C",X"68",X"9D",X"C0",X"92",X"0C",X"D8",X"C0",X"E0",X"F0",X"FE",
		X"00",X"80",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"3A",X"51",X"8A",X"12",X"00",X"00",X"30",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"0C",X"1E",X"51",X"1C",X"40",X"3A",X"33",X"07",X"0F",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"2B",X"0C",X"14",X"08",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"70",X"F8",X"D0",X"F8",X"50",X"20",X"00",X"00",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"0B",X"2B",X"60",X"FA",X"71",X"7A",X"4C",X"4E",X"82",X"6C",X"70",X"9C",
		X"00",X"00",X"60",X"10",X"08",X"04",X"80",X"C0",X"80",X"DA",X"90",X"08",X"18",X"80",X"00",X"00",
		X"BC",X"DE",X"BE",X"ED",X"DA",X"B4",X"FA",X"FF",X"7F",X"B7",X"EF",X"AF",X"F2",X"61",X"01",X"00",
		X"00",X"00",X"28",X"00",X"2A",X"54",X"82",X"9E",X"27",X"9E",X"F5",X"BB",X"7F",X"5F",X"3F",X"3F",
		X"00",X"00",X"01",X"00",X"00",X"00",X"02",X"04",X"01",X"2A",X"47",X"6D",X"22",X"00",X"02",X"18",
		X"0F",X"17",X"25",X"5B",X"F7",X"FF",X"EE",X"FB",X"FF",X"FF",X"27",X"EA",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"04",X"05",X"03",X"0D",X"0F",X"1B",X"09",X"07",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"40",X"10",X"08",X"04",X"00",X"00",X"00",X"0A",X"90",X"00",X"18",X"00",
		X"01",X"00",X"14",X"08",X"00",X"00",X"08",X"20",X"28",X"48",X"20",X"00",X"00",X"01",X"00",X"00",
		X"00",X"00",X"00",X"20",X"42",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"80",X"70",X"70",X"00",X"00",X"00",X"04",X"00",
		X"00",X"00",X"10",X"10",X"01",X"02",X"80",X"08",X"86",X"25",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"44",X"80",X"20",X"24",X"08",X"80",X"44",X"60",X"00",X"58",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"10",X"82",X"46",X"00",X"14",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"4E",X"FE",X"DE",X"85",X"87",X"C7",X"A7",X"8B",X"FF",
		X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"07",X"47",X"CE",X"CD",X"C6",X"7C",X"7E",X"AC",X"50",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"1A",X"3E",X"7E",X"2F",X"7F",X"FF",X"20",X"EF",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",
		X"FE",X"7F",X"E2",X"7F",X"7F",X"7F",X"FF",X"FE",X"54",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"A0",X"60",X"A0",X"50",X"A0",X"F0",X"58",X"A8",X"70",X"A8",X"D4",X"F8",
		X"00",X"00",X"C4",X"AE",X"77",X"AF",X"D6",X"FF",X"FF",X"FF",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"FA",X"B4",X"3C",X"F8",X"D4",X"F8",X"94",X"58",X"B0",X"60",X"C0",X"00",X"00",X"00",X"00",
		X"FF",X"47",X"6F",X"FF",X"FD",X"FE",X"7D",X"7F",X"AE",X"76",X"BD",X"FA",X"94",X"08",X"00",X"00",
		X"00",X"00",X"00",X"0A",X"15",X"7F",X"FD",X"FB",X"FF",X"7F",X"FF",X"7F",X"FF",X"BF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"03",X"02",X"07",X"0F",X"19",X"0F",X"0F",X"0F",X"1F",X"1C",X"0E",
		X"FF",X"FF",X"FF",X"7F",X"7F",X"FF",X"FF",X"FE",X"FF",X"57",X"2B",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0B",X"07",X"03",X"07",X"02",X"04",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"70",X"88",X"B4",X"D8",X"F8",X"74",X"EA",X"7E",X"7E",X"B3",X"4D",X"CA",X"B4",X"9A",X"D6",X"FC",
		X"00",X"71",X"CE",X"FD",X"2A",X"F7",X"EC",X"D7",X"B7",X"57",X"2D",X"26",X"41",X"6B",X"83",X"DB",
		X"FE",X"FE",X"FC",X"FE",X"7B",X"9D",X"CA",X"C4",X"92",X"3C",X"C0",X"C0",X"A0",X"40",X"80",X"00",
		X"F7",X"EB",X"FD",X"FB",X"FF",X"EF",X"FF",X"FD",X"FE",X"7F",X"B7",X"CB",X"FC",X"BA",X"11",X"00",
		X"00",X"00",X"00",X"01",X"A1",X"65",X"77",X"8B",X"6D",X"3E",X"1A",X"15",X"CB",X"EB",X"B4",X"79",
		X"00",X"00",X"00",X"00",X"08",X"00",X"02",X"00",X"01",X"02",X"04",X"02",X"01",X"4B",X"67",X"0F",
		X"DF",X"FF",X"FF",X"5F",X"3F",X"D7",X"ED",X"FF",X"7F",X"EE",X"55",X"0E",X"1D",X"08",X"00",X"00",
		X"1F",X"1E",X"0C",X"09",X"12",X"04",X"01",X"10",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"C0",X"60",X"80",X"00",X"00",X"80",X"B8",X"70",X"64",X"18",X"B0",
		X"00",X"80",X"00",X"00",X"24",X"56",X"83",X"04",X"37",X"50",X"BA",X"D5",X"B6",X"68",X"6B",X"9C",
		X"24",X"2A",X"00",X"86",X"0A",X"11",X"82",X"04",X"12",X"18",X"40",X"80",X"20",X"40",X"80",X"00",
		X"D4",X"0A",X"54",X"09",X"28",X"00",X"0A",X"21",X"18",X"56",X"A5",X"02",X"10",X"22",X"01",X"00",
		X"00",X"00",X"00",X"00",X"20",X"00",X"20",X"82",X"28",X"10",X"0A",X"14",X"08",X"02",X"24",X"59",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"01",X"00",X"04",X"02",X"00",X"48",X"64",X"0C",
		X"55",X"2A",X"18",X"06",X"1A",X"94",X"0D",X"0B",X"02",X"40",X"10",X"00",X"09",X"00",X"00",X"00",
		X"10",X"1A",X"0C",X"09",X"10",X"04",X"00",X"10",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"F0",X"70",X"28",X"28",X"3F",X"1B",X"19",X"19",X"1B",X"3F",X"22",X"22",X"70",X"F0",X"00",
		X"00",X"7F",X"C0",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"C0",X"7F",X"00",
		X"00",X"FC",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"FC",X"00",
		X"00",X"0F",X"1C",X"10",X"10",X"F0",X"90",X"90",X"90",X"90",X"F0",X"10",X"10",X"1C",X"0F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"A0",X"48",X"12",X"BA",X"5B",X"E6",X"F4",X"F8",X"B0",X"90",X"D8",X"48",X"02",X"08",X"00",
		X"00",X"02",X"07",X"0C",X"0F",X"06",X"E7",X"3F",X"F6",X"03",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"F0",X"08",X"08",X"08",X"08",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"80",X"BF",X"BE",X"BE",X"BE",X"BE",X"BF",X"80",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"60",X"30",X"18",X"00",X"00",X"00",X"00",
		X"C0",X"60",X"30",X"18",X"0C",X"06",X"03",X"23",X"63",X"63",X"00",X"00",X"63",X"63",X"22",X"00",
		X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"10",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"FC",X"FF",X"F1",X"F8",X"FE",X"F1",X"F9",X"FC",X"FC",X"04",X"04",X"00",X"04",X"00",X"00",
		X"00",X"04",X"50",X"04",X"30",X"69",X"C0",X"80",X"00",X"40",X"24",X"00",X"80",X"60",X"00",X"00",
		X"00",X"00",X"00",X"06",X"04",X"05",X"04",X"FF",X"7F",X"06",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"77",X"77",X"77",X"77",X"7F",X"7F",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"60",X"F0",X"D0",X"74",X"7C",X"74",X"D4",X"F8",X"70",X"00",X"00",X"00",X"00",
		X"00",X"00",X"9C",X"BE",X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"BE",X"9C",X"80",X"00",X"00",
		X"00",X"E0",X"F0",X"E0",X"E0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"7C",X"FD",X"FD",X"FD",X"FD",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"08",X"08",X"F8",X"08",X"08",X"00",X"F8",X"10",X"20",X"10",X"F8",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"81",X"01",X"01",X"01",X"01",X"01",X"01",X"FF",
		X"FF",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"FF",
		X"00",X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"FF",X"80",X"80",X"80",X"80",X"80",X"80",
		X"7F",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"7F",
		X"00",X"7F",X"40",X"40",X"40",X"40",X"40",X"40",X"FF",X"81",X"81",X"81",X"81",X"81",X"81",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
