library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity cclimber_tile_bit1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of cclimber_tile_bit1 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"1C",X"26",X"63",X"63",X"63",X"32",X"1C",X"00",X"0C",X"1C",X"0C",X"0C",X"0C",X"0C",X"3F",X"00",
		X"3E",X"63",X"07",X"1E",X"3C",X"70",X"7F",X"00",X"3F",X"06",X"0C",X"1E",X"03",X"63",X"3E",X"00",
		X"0E",X"1E",X"36",X"66",X"7F",X"06",X"06",X"00",X"3E",X"30",X"3E",X"03",X"03",X"33",X"1E",X"00",
		X"1E",X"30",X"60",X"7E",X"63",X"63",X"3E",X"00",X"3F",X"23",X"06",X"0C",X"18",X"18",X"18",X"00",
		X"3C",X"62",X"72",X"3C",X"4F",X"43",X"3E",X"00",X"3E",X"63",X"63",X"3F",X"03",X"06",X"3C",X"00",
		X"1C",X"36",X"63",X"63",X"7F",X"63",X"63",X"00",X"7E",X"63",X"63",X"7E",X"63",X"63",X"7E",X"00",
		X"1E",X"33",X"60",X"60",X"60",X"33",X"1E",X"00",X"7C",X"66",X"63",X"63",X"63",X"66",X"7C",X"00",
		X"3F",X"30",X"30",X"3E",X"30",X"30",X"3F",X"00",X"7F",X"60",X"60",X"7E",X"60",X"60",X"60",X"00",
		X"1F",X"30",X"60",X"67",X"63",X"33",X"1F",X"00",X"63",X"63",X"63",X"7F",X"63",X"63",X"63",X"00",
		X"3F",X"0C",X"0C",X"0C",X"0C",X"0C",X"3F",X"00",X"03",X"03",X"03",X"03",X"03",X"63",X"3E",X"00",
		X"63",X"66",X"6C",X"78",X"7C",X"6E",X"67",X"00",X"30",X"30",X"30",X"30",X"30",X"30",X"3F",X"00",
		X"63",X"77",X"7F",X"7F",X"6B",X"63",X"63",X"00",X"63",X"73",X"7B",X"7F",X"6F",X"67",X"63",X"00",
		X"3E",X"63",X"63",X"63",X"63",X"63",X"3E",X"00",X"7E",X"63",X"63",X"63",X"7E",X"60",X"60",X"00",
		X"3E",X"63",X"63",X"63",X"6F",X"66",X"3D",X"00",X"7E",X"63",X"63",X"67",X"7C",X"6E",X"67",X"00",
		X"3C",X"66",X"60",X"3E",X"03",X"63",X"3E",X"00",X"3F",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"00",
		X"63",X"63",X"63",X"63",X"63",X"63",X"3E",X"00",X"63",X"63",X"63",X"77",X"3E",X"1C",X"08",X"00",
		X"63",X"63",X"6B",X"7F",X"7F",X"36",X"22",X"00",X"63",X"77",X"3E",X"1C",X"3E",X"77",X"63",X"00",
		X"33",X"33",X"12",X"1E",X"0C",X"0C",X"0C",X"00",X"7F",X"07",X"0E",X"1C",X"38",X"70",X"7F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"06",X"06",X"00",X"00",X"18",X"30",X"30",X"30",X"30",X"30",X"18",X"00",
		X"18",X"0C",X"0C",X"0C",X"0C",X"0C",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",
		X"00",X"00",X"00",X"18",X"1C",X"04",X"08",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"0F",X"0F",X"0E",X"09",X"03",X"06",X"02",X"00",X"F0",X"F0",X"70",X"90",X"C0",X"60",X"20",X"00",
		X"00",X"01",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"80",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"07",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"1F",X"F8",X"F8",X"F8",X"F0",X"F0",X"F0",X"F0",X"E0",
		X"1F",X"1C",X"10",X"27",X"29",X"01",X"00",X"00",X"E0",X"E0",X"60",X"20",X"A0",X"A0",X"A0",X"00",
		X"00",X"01",X"0F",X"0F",X"1F",X"1F",X"1F",X"1F",X"00",X"80",X"E0",X"E0",X"F0",X"F0",X"E0",X"E0",
		X"3F",X"3F",X"3F",X"3F",X"7F",X"7F",X"7F",X"7F",X"E0",X"E0",X"C0",X"C0",X"C0",X"C0",X"00",X"C0",
		X"10",X"10",X"10",X"10",X"10",X"18",X"1F",X"1F",X"08",X"08",X"08",X"08",X"08",X"18",X"F8",X"F8",
		X"0F",X"0F",X"07",X"07",X"03",X"03",X"01",X"00",X"F0",X"F0",X"E0",X"E0",X"C0",X"C0",X"80",X"00",
		X"00",X"00",X"0F",X"1F",X"1F",X"1F",X"1F",X"1F",X"00",X"00",X"F0",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"1F",X"1F",X"1F",X"1F",X"18",X"10",X"10",X"10",X"F8",X"F8",X"F8",X"F8",X"18",X"08",X"08",X"08",
		X"04",X"0C",X"0C",X"1E",X"1F",X"0F",X"0F",X"0F",X"02",X"06",X"04",X"04",X"84",X"FC",X"F8",X"F8",
		X"0F",X"0F",X"0F",X"0F",X"07",X"02",X"00",X"00",X"F0",X"E0",X"C0",X"80",X"80",X"00",X"00",X"00",
		X"00",X"03",X"07",X"0F",X"0F",X"0F",X"0F",X"1F",X"00",X"C0",X"F8",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"1F",X"1F",X"37",X"20",X"20",X"20",X"60",X"40",X"F8",X"F8",X"F8",X"F0",X"30",X"10",X"20",X"20",
		X"0E",X"09",X"07",X"0F",X"0F",X"0F",X"0E",X"09",X"38",X"C8",X"F0",X"F8",X"F8",X"F8",X"38",X"C8",
		X"07",X"07",X"07",X"03",X"01",X"00",X"00",X"00",X"70",X"F0",X"F0",X"E0",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"00",X"00",X"00",X"00",X"00",X"C0",X"F0",X"F8",
		X"0F",X"0F",X"0E",X"09",X"07",X"0F",X"0F",X"0F",X"F8",X"F8",X"38",X"C8",X"F0",X"F8",X"F8",X"F8",
		X"00",X"07",X"0F",X"0F",X"1F",X"00",X"1F",X"1D",X"3E",X"DE",X"EC",X"F4",X"F8",X"F8",X"70",X"B0",
		X"3F",X"1F",X"1F",X"1F",X"07",X"00",X"00",X"00",X"C0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",
		X"07",X"07",X"0F",X"00",X"1F",X"1F",X"3F",X"3F",X"F8",X"FC",X"FC",X"7C",X"B8",X"D8",X"E0",X"F0",
		X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"08",X"06",X"03",X"00",X"00",X"00",
		X"00",X"00",X"01",X"0E",X"F0",X"00",X"00",X"00",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"10",X"10",X"10",X"08",X"08",X"08",X"04",X"08",X"08",X"84",X"82",X"40",X"40",X"30",X"0C",
		X"00",X"10",X"21",X"C1",X"02",X"02",X"0C",X"30",X"88",X"88",X"00",X"00",X"00",X"10",X"10",X"20",
		X"04",X"01",X"01",X"00",X"00",X"00",X"11",X"11",X"0C",X"30",X"40",X"40",X"83",X"84",X"08",X"00",
		X"30",X"0C",X"02",X"02",X"41",X"21",X"10",X"10",X"20",X"10",X"10",X"10",X"08",X"08",X"08",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"02",X"00",X"00",X"00",X"0F",X"70",X"80",X"00",X"00",
		X"00",X"00",X"00",X"C0",X"06",X"01",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"80",X"F0",X"1E",X"01",X"00",X"00",
		X"E0",X"00",X"01",X"0F",X"78",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"08",X"10",X"08",X"08",X"04",X"04",X"00",X"88",X"88",X"00",X"07",X"80",X"40",X"30",X"08",
		X"11",X"11",X"00",X"E0",X"01",X"02",X"0C",X"10",X"08",X"10",X"08",X"10",X"10",X"20",X"20",X"00",
		X"00",X"04",X"04",X"08",X"08",X"10",X"08",X"10",X"08",X"30",X"40",X"80",X"07",X"00",X"88",X"88",
		X"10",X"0C",X"02",X"01",X"E0",X"00",X"11",X"11",X"00",X"20",X"20",X"10",X"10",X"08",X"10",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"1E",X"F0",X"80",X"00",X"07",
		X"00",X"00",X"80",X"71",X"0F",X"01",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"80",X"00",X"18",X"07",X"00",X"00",
		X"C0",X"00",X"01",X"00",X"18",X"E0",X"00",X"00",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"10",X"10",X"10",X"00",X"00",X"00",X"04",X"08",X"88",X"84",X"C3",X"00",X"00",X"20",X"1C",
		X"10",X"11",X"21",X"C3",X"00",X"00",X"04",X"31",X"88",X"08",X"08",X"08",X"10",X"10",X"10",X"20",
		X"04",X"08",X"08",X"08",X"10",X"10",X"10",X"11",X"1C",X"20",X"00",X"00",X"C3",X"84",X"88",X"08",
		X"38",X"04",X"00",X"00",X"C3",X"21",X"11",X"10",X"20",X"10",X"10",X"10",X"08",X"08",X"08",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"00",X"00",X"07",X"18",X"00",X"80",X"00",X"03",
		X"00",X"00",X"E0",X"18",X"00",X"01",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",
		X"06",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"80",X"70",X"00",X"01",X"00",X"00",
		X"F0",X"00",X"01",X"0E",X"00",X"80",X"00",X"00",X"60",X"00",X"80",X"00",X"00",X"00",X"00",X"00",
		X"11",X"11",X"11",X"10",X"10",X"08",X"08",X"08",X"08",X"08",X"04",X"84",X"81",X"60",X"00",X"00",
		X"10",X"10",X"20",X"21",X"81",X"06",X"00",X"00",X"88",X"88",X"88",X"08",X"08",X"10",X"10",X"10",
		X"08",X"08",X"08",X"10",X"10",X"11",X"11",X"11",X"00",X"00",X"60",X"81",X"84",X"04",X"08",X"08",
		X"00",X"00",X"06",X"81",X"21",X"20",X"10",X"10",X"10",X"10",X"10",X"08",X"08",X"88",X"88",X"88",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"06",X"00",X"00",X"01",X"00",X"70",X"80",X"00",X"0F",
		X"00",X"00",X"80",X"00",X"0E",X"01",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"60",
		X"07",X"07",X"07",X"3F",X"23",X"77",X"2F",X"0F",X"E8",X"FC",X"E8",X"F8",X"C0",X"E0",X"F0",X"F0",
		X"09",X"01",X"07",X"03",X"03",X"03",X"03",X"01",X"90",X"80",X"E0",X"C0",X"C0",X"C0",X"C0",X"80",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"30",X"60",X"60",X"C0",X"C0",X"80",X"C0",X"C0",
		X"13",X"3B",X"13",X"1F",X"07",X"07",X"07",X"07",X"C0",X"C0",X"C4",X"FE",X"E4",X"E0",X"E0",X"E0",
		X"1F",X"1F",X"1F",X"3F",X"2F",X"77",X"2F",X"0F",X"A0",X"F0",X"A0",X"E0",X"80",X"E0",X"F0",X"90",
		X"1F",X"09",X"09",X"03",X"01",X"00",X"00",X"00",X"80",X"E0",X"E0",X"F0",X"F0",X"F8",X"70",X"20",
		X"30",X"18",X"18",X"0C",X"0C",X"06",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"4F",X"EF",X"4F",X"7F",X"1F",X"1F",X"1F",X"1F",X"00",X"00",X"20",X"F0",X"A0",X"80",X"80",X"80",
		X"17",X"3F",X"17",X"1F",X"03",X"07",X"0F",X"0F",X"E0",X"E0",X"E0",X"FC",X"C4",X"EE",X"F4",X"F0",
		X"09",X"01",X"07",X"03",X"03",X"03",X"03",X"01",X"90",X"80",X"E0",X"C0",X"C0",X"C0",X"C0",X"80",
		X"0C",X"06",X"06",X"03",X"03",X"01",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",
		X"03",X"03",X"43",X"7F",X"47",X"07",X"07",X"07",X"C8",X"DC",X"C8",X"F8",X"E0",X"E0",X"E0",X"E0",
		X"01",X"01",X"09",X"1F",X"09",X"07",X"0F",X"09",X"FA",X"FF",X"FA",X"FE",X"F0",X"E0",X"E0",X"F0",
		X"01",X"07",X"07",X"0F",X"0F",X"1F",X"0E",X"04",X"F8",X"90",X"90",X"C0",X"80",X"00",X"00",X"00",
		X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"60",X"F0",X"F0",
		X"04",X"0E",X"04",X"07",X"01",X"01",X"01",X"01",X"F0",X"F0",X"F2",X"FF",X"FA",X"F8",X"F8",X"F8",
		X"8C",X"08",X"DD",X"CB",X"0A",X"76",X"28",X"05",X"CD",X"E7",X"31",X"28",X"0F",X"01",X"04",X"00",
		X"21",X"11",X"39",X"11",X"15",X"39",X"ED",X"B0",X"DD",X"CB",X"09",X"C6",X"DD",X"CB",X"0E",X"5E",
		X"20",X"C7",X"CD",X"F9",X"18",X"28",X"C5",X"18",X"62",X"DD",X"CB",X"0E",X"E6",X"CD",X"49",X"1F",
		X"DA",X"F6",X"11",X"EF",X"3A",X"CA",X"DD",X"11",X"CD",X"0D",X"19",X"0E",X"01",X"CD",X"C0",X"2D",
		X"0E",X"13",X"DD",X"CB",X"0F",X"56",X"20",X"1E",X"21",X"FB",X"0C",X"CD",X"30",X"00",X"38",X"14",
		X"DD",X"CB",X"09",X"D6",X"CD",X"0D",X"19",X"0E",X"00",X"CD",X"D8",X"18",X"0E",X"82",X"CD",X"C0",
		X"2D",X"C3",X"8C",X"08",X"0E",X"07",X"CD",X"73",X"24",X"2E",X"2D",X"41",X"2B",X"DD",X"CB",X"0F",
		X"56",X"28",X"08",X"21",X"FB",X"0C",X"CD",X"30",X"00",X"28",X"D5",X"0E",X"11",X"CD",X"73",X"19",
		X"18",X"15",X"DD",X"CB",X"0E",X"66",X"20",X"0F",X"CD",X"F9",X"18",X"16",X"E1",X"CD",X"83",X"1C",
		X"DD",X"CB",X"09",X"D6",X"C3",X"1D",X"12",X"0E",X"01",X"CD",X"C0",X"2D",X"16",X"E2",X"CD",X"83",
		X"1C",X"DD",X"CB",X"09",X"F6",X"DD",X"CB",X"09",X"D6",X"C3",X"1C",X"10",X"2A",X"37",X"39",X"DD",
		X"CB",X"76",X"66",X"C2",X"2C",X"12",X"E5",X"CD",X"E5",X"04",X"E1",X"22",X"37",X"39",X"DD",X"CB",
		X"0A",X"6E",X"20",X"E1",X"DD",X"36",X"0C",X"07",X"DD",X"CB",X"0A",X"76",X"28",X"05",X"0E",X"6B",
		X"CD",X"56",X"2B",X"0E",X"6D",X"CD",X"56",X"2B",X"0E",X"02",X"CD",X"59",X"1A",X"CD",X"B8",X"34",
		X"CD",X"E3",X"18",X"28",X"C0",X"EF",X"2C",X"28",X"14",X"CD",X"F1",X"34",X"CD",X"9E",X"33",X"CD",
		X"E3",X"18",X"28",X"B1",X"EF",X"2C",X"38",X"F1",X"CD",X"E3",X"18",X"38",X"E8",X"CD",X"8F",X"31",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7C",X"7C",X"00",X"00",X"00",X"00",X"00",X"00",X"7C",X"7C",X"7C",X"00",X"00",X"00",X"00",X"00",
		X"7C",X"7C",X"7C",X"7C",X"00",X"00",X"00",X"00",X"7C",X"7C",X"7C",X"7C",X"7C",X"00",X"00",X"00",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"00",X"00",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"00",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"CB",X"0A",X"5E",X"20",X"05",X"16",X"49",X"CD",
		X"83",X"1C",X"DD",X"7E",X"07",X"CD",X"21",X"00",X"18",X"1F",X"26",X"48",X"4B",X"B3",X"9D",X"CB",
		X"77",X"28",X"3C",X"DD",X"CB",X"08",X"F6",X"DD",X"CB",X"09",X"EE",X"CD",X"49",X"1F",X"28",X"48",
		X"21",X"8F",X"14",X"CD",X"61",X"14",X"28",X"C2",X"21",X"9A",X"14",X"CD",X"61",X"14",X"28",X"BA",
		X"CD",X"49",X"1F",X"28",X"33",X"EF",X"24",X"28",X"25",X"CD",X"22",X"1E",X"28",X"25",X"EF",X"28",
		X"28",X"02",X"37",X"DF",X"CD",X"46",X"13",X"EF",X"29",X"DF",X"CD",X"5E",X"14",X"28",X"9B",X"AF",
		X"C3",X"31",X"22",X"1E",X"08",X"18",X"02",X"1E",X"FF",X"CD",X"15",X"20",X"18",X"EC",X"CD",X"BA",
		X"1F",X"18",X"E7",X"CD",X"0D",X"20",X"18",X"E2",X"DD",X"CB",X"08",X"FE",X"0E",X"02",X"CD",X"73",
		X"24",X"30",X"2F",X"33",X"0B",X"0E",X"11",X"CD",X"73",X"19",X"CD",X"04",X"20",X"18",X"CB",X"DD",
		X"CB",X"08",X"56",X"20",X"1C",X"DD",X"CB",X"08",X"C6",X"DD",X"CB",X"0A",X"5E",X"20",X"12",X"DD",
		X"7E",X"03",X"E6",X"0F",X"20",X"06",X"DD",X"CB",X"09",X"6E",X"28",X"05",X"16",X"29",X"CD",X"83",
		X"1C",X"CD",X"F3",X"1F",X"18",X"A4",X"CD",X"15",X"25",X"18",X"CF",X"CD",X"46",X"13",X"CD",X"3F",
		X"20",X"EF",X"2C",X"38",X"06",X"CD",X"46",X"13",X"CD",X"5C",X"20",X"EF",X"5D",X"DF",X"18",X"8A",
		X"CD",X"49",X"1F",X"DF",X"DD",X"CB",X"08",X"FE",X"0E",X"0A",X"CD",X"73",X"24",X"0A",X"09",X"08",
		X"01",X"0E",X"08",X"11",X"68",X"84",X"92",X"A1",X"E0",X"20",X"10",X"2C",X"43",X"91",X"0A",X"21",
		X"92",X"85",X"48",X"21",X"12",X"0C",X"02",X"01",X"11",X"0A",X"92",X"04",X"22",X"5E",X"40",X"80",
		X"19",X"26",X"40",X"92",X"A5",X"88",X"80",X"94",X"00",X"E8",X"34",X"02",X"09",X"91",X"22",X"42",
		X"AA",X"41",X"50",X"2D",X"02",X"04",X"04",X"03",X"24",X"54",X"8A",X"04",X"18",X"60",X"80",X"80",
		X"0C",X"13",X"20",X"45",X"4A",X"91",X"80",X"89",X"C0",X"30",X"8C",X"04",X"22",X"12",X"49",X"11",
		X"92",X"44",X"2A",X"11",X"20",X"16",X"09",X"00",X"29",X"02",X"22",X"44",X"88",X"10",X"90",X"60",
		X"00",X"00",X"00",X"01",X"03",X"04",X"02",X"00",X"00",X"00",X"00",X"80",X"C0",X"20",X"40",X"04",
		X"01",X"00",X"04",X"40",X"80",X"1B",X"24",X"00",X"80",X"00",X"20",X"42",X"00",X"A2",X"5C",X"00",
		X"00",X"00",X"00",X"01",X"03",X"04",X"02",X"00",X"00",X"00",X"00",X"80",X"C0",X"20",X"40",X"00",
		X"01",X"00",X"00",X"04",X"01",X"4B",X"10",X"00",X"80",X"00",X"00",X"40",X"00",X"66",X"92",X"00",
		X"00",X"07",X"08",X"11",X"0F",X"04",X"22",X"70",X"00",X"E0",X"10",X"88",X"F0",X"20",X"44",X"0E",
		X"F9",X"FC",X"F0",X"E0",X"F1",X"F1",X"DF",X"80",X"9F",X"3F",X"0F",X"07",X"8F",X"8F",X"FB",X"01",
		X"03",X"04",X"09",X"14",X"63",X"A4",X"9C",X"42",X"B0",X"50",X"0C",X"B2",X"45",X"3A",X"C5",X"11",
		X"4A",X"24",X"43",X"2D",X"42",X"28",X"15",X"02",X"8A",X"66",X"19",X"85",X"EA",X"14",X"60",X"80",
		X"0C",X"13",X"2A",X"15",X"24",X"A2",X"A2",X"99",X"D0",X"28",X"54",X"24",X"AB",X"29",X"52",X"49",
		X"4C",X"95",X"4A",X"29",X"40",X"2A",X"15",X"00",X"15",X"91",X"6A",X"44",X"48",X"30",X"90",X"60",
		X"01",X"06",X"28",X"57",X"A1",X"98",X"66",X"51",X"40",X"A8",X"14",X"42",X"B4",X"C2",X"24",X"52",
		X"88",X"A3",X"5C",X"A2",X"4D",X"30",X"0A",X"0D",X"42",X"39",X"25",X"C6",X"28",X"90",X"20",X"C0",
		X"06",X"09",X"0C",X"12",X"22",X"56",X"89",X"A8",X"00",X"A8",X"54",X"02",X"94",X"52",X"A9",X"32",
		X"92",X"4A",X"94",X"D5",X"24",X"2A",X"14",X"0B",X"99",X"4A",X"4A",X"24",X"A8",X"54",X"C8",X"30",
		X"00",X"00",X"60",X"F0",X"70",X"38",X"18",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",
		X"79",X"70",X"20",X"02",X"00",X"01",X"03",X"00",X"72",X"3E",X"1C",X"8C",X"C4",X"90",X"88",X"84",
		X"84",X"14",X"48",X"08",X"28",X"88",X"10",X"50",X"8C",X"24",X"08",X"50",X"90",X"08",X"58",X"04",
		X"89",X"22",X"04",X"54",X"4A",X"82",X"26",X"04",X"15",X"22",X"82",X"0A",X"05",X"A1",X"45",X"01",
		X"2C",X"84",X"08",X"28",X"88",X"06",X"2A",X"01",X"90",X"50",X"28",X"08",X"28",X"C8",X"14",X"84",
		X"50",X"10",X"B0",X"10",X"20",X"60",X"A0",X"10",X"4A",X"06",X"94",X"04",X"58",X"28",X"10",X"90",
		X"84",X"20",X"02",X"90",X"4A",X"04",X"91",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DD",X"CB",X"09",X"46",X"CD",X"BF",X"26",X"CD",X"09",X"27",X"DD",X"CB",X"09",X"66",X"CD",X"BF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"40",X"40",X"40",X"40",X"80",X"80",X"80",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"20",X"20",X"20",X"20",
		X"04",X"04",X"04",X"04",X"08",X"08",X"08",X"08",X"20",X"20",X"40",X"40",X"40",X"80",X"80",X"80",
		X"04",X"08",X"08",X"08",X"10",X"10",X"10",X"20",X"00",X"00",X"00",X"00",X"00",X"C0",X"38",X"07",
		X"00",X"00",X"80",X"70",X"0E",X"01",X"00",X"00",X"E0",X"1C",X"03",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"38",X"07",X"00",X"00",X"80",X"70",X"0E",X"01",X"00",X"00",
		X"E0",X"1C",X"03",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"80",X"40",X"20",X"10",X"08",X"04",X"02",X"01",X"80",X"40",X"20",X"10",X"08",X"04",X"02",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"C0",X"30",X"0C",X"03",
		X"C0",X"30",X"0C",X"03",X"00",X"00",X"00",X"00",X"FF",X"FE",X"FC",X"F8",X"F0",X"F8",X"FC",X"FF",
		X"80",X"C0",X"E0",X"F0",X"F8",X"FC",X"FE",X"FF",X"01",X"01",X"01",X"02",X"02",X"02",X"04",X"04",
		X"E0",X"1C",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"70",X"0E",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"38",X"07",X"4F",X"41",X"79",X"A7",X"28",X"EF",X"3E",X"20",
		X"77",X"23",X"10",X"FC",X"C9",X"3A",X"06",X"00",X"5F",X"C6",X"10",X"CD",X"D0",X"26",X"3A",X"07",
		X"00",X"93",X"4F",X"11",X"18",X"39",X"E5",X"21",X"13",X"39",X"CD",X"EA",X"27",X"E1",X"A7",X"C8",
		X"4F",X"06",X"00",X"EB",X"ED",X"B0",X"EB",X"C9",X"11",X"17",X"39",X"E5",X"0E",X"04",X"21",X"15",
		X"39",X"CD",X"EA",X"27",X"E1",X"18",X"02",X"3E",X"22",X"4F",X"E6",X"1F",X"C3",X"07",X"01",X"2A",
		X"47",X"39",X"3E",X"84",X"5E",X"BB",X"C8",X"23",X"56",X"ED",X"53",X"11",X"39",X"23",X"22",X"47",
		X"39",X"21",X"7F",X"39",X"3E",X"09",X"11",X"01",X"28",X"CD",X"FF",X"26",X"3A",X"11",X"39",X"57",
		X"3E",X"E1",X"CD",X"1A",X"27",X"36",X"20",X"23",X"E5",X"11",X"0E",X"00",X"21",X"0A",X"28",X"3A",
		X"11",X"39",X"D6",X"3F",X"28",X"15",X"47",X"19",X"7E",X"FE",X"04",X"28",X"07",X"A7",X"20",X"09",
		X"05",X"23",X"18",X"F4",X"21",X"43",X"29",X"18",X"02",X"10",X"EC",X"7B",X"EB",X"E1",X"CD",X"FF",
		X"26",X"E5",X"21",X"07",X"00",X"7E",X"2B",X"96",X"4F",X"2B",X"2B",X"11",X"40",X"39",X"3A",X"12",
		X"39",X"A7",X"ED",X"52",X"EB",X"06",X"04",X"BE",X"28",X"14",X"38",X"11",X"23",X"10",X"F8",X"2B",
		X"96",X"19",X"2B",X"91",X"28",X"03",X"30",X"FB",X"81",X"1E",X"23",X"18",X"05",X"2B",X"96",X"19",
		X"1E",X"2A",X"86",X"E1",X"CD",X"D7",X"26",X"01",X"0A",X"00",X"B7",X"ED",X"42",X"73",X"23",X"C3",
		X"AE",X"26",X"3A",X"07",X"39",X"A1",X"28",X"0C",X"79",X"FE",X"08",X"0E",X"72",X"28",X"02",X"0E",
		X"44",X"CD",X"56",X"2B",X"3C",X"C9",X"2A",X"17",X"39",X"BF",X"DD",X"CB",X"08",X"56",X"C8",X"AF",
		X"BD",X"20",X"05",X"BC",X"C8",X"3C",X"BC",X"C8",X"21",X"7F",X"39",X"0E",X"05",X"CD",X"DA",X"26",
		X"CD",X"09",X"27",X"CD",X"E6",X"26",X"C3",X"AE",X"26",X"1A",X"B9",X"30",X"01",X"4F",X"91",X"12",
		X"5E",X"23",X"56",X"79",X"E5",X"69",X"26",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"38",X"38",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"1E",X"3F",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"07",X"0F",X"1C",X"38",X"30",X"00",X"00",X"FC",X"FE",X"FF",X"71",X"61",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"81",X"C3",X"C3",X"00",X"00",X"00",X"00",X"E0",X"F0",X"F8",X"39",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"01",X"00",X"00",X"00",X"08",X"38",X"3C",X"DC",X"CE",
		X"00",X"1C",X"18",X"38",X"38",X"38",X"39",X"38",X"3C",X"FC",X"E0",X"E0",X"E4",X"FC",X"F8",X"E0",
		X"31",X"30",X"30",X"30",X"30",X"30",X"31",X"33",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"C0",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"70",X"70",X"70",X"30",X"39",X"1D",X"0D",
		X"E0",X"E1",X"E1",X"C3",X"FE",X"FC",X"F0",X"C0",X"C7",X"9E",X"8F",X"0F",X"0C",X"1C",X"18",X"18",
		X"18",X"18",X"F8",X"F0",X"70",X"30",X"30",X"61",X"3F",X"30",X"30",X"60",X"60",X"E0",X"C0",X"C0",
		X"0C",X"1F",X"1F",X"3B",X"30",X"70",X"70",X"E0",X"00",X"00",X"80",X"C0",X"C0",X"E0",X"E0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"03",
		X"07",X"1F",X"7F",X"F8",X"D8",X"9C",X"9C",X"0E",X"81",X"E1",X"F0",X"78",X"38",X"38",X"38",X"38",
		X"CF",X"C7",X"C7",X"E3",X"E1",X"E1",X"60",X"70",X"38",X"38",X"A8",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"60",X"60",X"60",X"60",X"60",X"70",X"70",X"76",X"3F",X"3E",X"3E",X"37",X"33",X"31",X"30",X"30",
		X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"03",X"03",X"03",X"03",X"06",X"04",X"00",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",
		X"38",X"30",X"30",X"70",X"70",X"71",X"01",X"00",X"61",X"E1",X"C3",X"C3",X"C3",X"87",X"86",X"01",
		X"C0",X"81",X"81",X"03",X"03",X"07",X"0E",X"0E",X"E1",X"C1",X"C7",X"FF",X"F8",X"60",X"70",X"70",
		X"C3",X"C7",X"8C",X"1C",X"38",X"30",X"70",X"70",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"E0",X"70",X"38",X"38",X"3C",X"3C",X"3C",X"00",X"00",X"00",X"00",X"00",X"10",X"38",X"70",
		X"03",X"03",X"03",X"03",X"03",X"01",X"00",X"00",X"0E",X"0E",X"0E",X"87",X"87",X"E7",X"F3",X"7B",
		X"38",X"70",X"E0",X"E0",X"E0",X"F8",X"3C",X"8F",X"70",X"70",X"30",X"38",X"38",X"38",X"38",X"20",
		X"70",X"70",X"30",X"20",X"00",X"00",X"00",X"00",X"3E",X"3E",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"70",X"30",X"38",X"08",X"00",X"00",X"00",X"00",X"70",X"70",X"38",X"38",X"1C",X"0F",X"07",X"01",
		X"00",X"00",X"00",X"00",X"01",X"8F",X"FE",X"F8",X"38",X"38",X"71",X"E3",X"C7",X"0E",X"0C",X"1C",
		X"60",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"87",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"38",X"70",X"F8",X"7C",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"2C",X"7E",X"4F",X"3C",X"C8",X"E5",X"CD",X"56",X"2B",X"E1",X"23",X"18",X"F4",X"CD",X"4E",X"1A",
		X"2A",X"6F",X"39",X"EB",X"CD",X"AE",X"2D",X"C4",X"60",X"2D",X"3E",X"C0",X"CD",X"E5",X"33",X"11",
		X"AF",X"3B",X"18",X"63",X"CD",X"7C",X"2D",X"2A",X"73",X"39",X"73",X"23",X"72",X"C9",X"2A",X"9C",
		X"37",X"3E",X"67",X"CD",X"E0",X"33",X"2A",X"C0",X"37",X"3E",X"69",X"CD",X"E0",X"33",X"2A",X"61",
		X"39",X"3E",X"6D",X"CD",X"E0",X"33",X"CD",X"7C",X"2D",X"ED",X"53",X"61",X"39",X"C9",X"ED",X"5B",
		X"6F",X"39",X"2A",X"61",X"39",X"CD",X"60",X"2D",X"3E",X"CD",X"CD",X"E5",X"33",X"22",X"61",X"39",
		X"3E",X"C7",X"CD",X"E5",X"33",X"EB",X"3E",X"C9",X"CD",X"E5",X"33",X"18",X"1A",X"18",X"48",X"FD",
		X"6E",X"02",X"FD",X"66",X"03",X"2B",X"22",X"5F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
