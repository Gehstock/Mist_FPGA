library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity mpa_43j is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of mpa_43j is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"01",X"02",X"02",X"03",X"03",X"04",X"04",X"05",X"60",X"01",X"58",X"01",X"50",X"01",X"48",X"01",
		X"40",X"01",X"38",X"01",X"39",X"10",X"39",X"20",X"39",X"30",X"39",X"48",X"39",X"60",X"39",X"70",
		X"39",X"80",X"39",X"98",X"39",X"B0",X"39",X"D0",X"B4",X"38",X"FF",X"58",X"8E",X"28",X"B4",X"38",
		X"00",X"19",X"24",X"2C",X"33",X"39",X"3E",X"43",X"48",X"4C",X"50",X"54",X"58",X"5B",X"5F",X"62",
		X"65",X"68",X"6B",X"6E",X"71",X"74",X"77",X"79",X"7C",X"7E",X"50",X"5E",X"6B",X"87",X"87",X"A2",
		X"A2",X"A3",X"02",X"00",X"A4",X"A5",X"02",X"00",X"A6",X"A7",X"02",X"A8",X"A9",X"01",X"AA",X"02",
		X"AB",X"AC",X"AD",X"02",X"00",X"AE",X"AF",X"02",X"B0",X"B1",X"01",X"B2",X"B3",X"B4",X"02",X"00",
		X"B5",X"B6",X"B7",X"02",X"00",X"00",X"00",X"B8",X"B9",X"02",X"00",X"00",X"00",X"BA",X"02",X"00",
		X"BB",X"BC",X"BD",X"02",X"BE",X"BF",X"01",X"C0",X"C1",X"02",X"00",X"C2",X"C3",X"C4",X"02",X"00",
		X"00",X"00",X"C5",X"C6",X"02",X"00",X"00",X"00",X"C7",X"C8",X"02",X"00",X"C9",X"CA",X"CB",X"02",
		X"CC",X"01",X"DA",X"DB",X"DC",X"02",X"00",X"00",X"F0",X"03",X"00",X"00",X"F0",X"02",X"00",X"00",
		X"F0",X"02",X"DD",X"DE",X"DF",X"01",X"0F",X"04",X"05",X"0F",X"24",X"27",X"0F",X"43",X"48",X"11",
		X"48",X"4E",X"12",X"4E",X"53",X"10",X"63",X"68",X"13",X"68",X"6C",X"0F",X"6C",X"6D",X"14",X"6D",
		X"6E",X"12",X"6E",X"74",X"10",X"89",X"8E",X"FF",X"0C",X"03",X"03",X"03",X"02",X"01",X"FF",X"3B",
		X"FF",X"70",X"FC",X"24",X"B9",X"FF",X"10",X"FC",X"24",X"3B",X"01",X"A0",X"FC",X"53",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"0A",X"0D",X"0F",X"11",X"13",X"15",X"16",X"18",X"19",X"1A",X"1B",X"1D",X"1E",X"1F",X"20",
		X"21",X"22",X"23",X"24",X"25",X"26",X"27",X"28",X"28",X"28",X"28",X"28",X"FF",X"1F",X"01",X"1C",
		X"04",X"0C",X"00",X"24",X"02",X"1D",X"05",X"20",X"08",X"0C",X"04",X"34",X"05",X"21",X"06",X"07",
		X"07",X"0C",X"0C",X"14",X"05",X"1E",X"08",X"1E",X"0F",X"0C",X"12",X"34",X"02",X"1B",X"03",X"1A",
		X"06",X"10",X"21",X"42",X"02",X"1D",X"04",X"1D",X"08",X"0F",X"27",X"42",X"05",X"20",X"06",X"20",
		X"0B",X"0C",X"2F",X"42",X"09",X"16",X"02",X"22",X"06",X"1C",X"3A",X"4E",X"0E",X"19",X"03",X"26",
		X"07",X"1C",X"40",X"4E",X"12",X"1D",X"05",X"2A",X"0A",X"1C",X"47",X"4E",X"05",X"20",X"05",X"26",
		X"08",X"0C",X"51",X"45",X"05",X"19",X"05",X"1F",X"11",X"0C",X"58",X"7F",X"08",X"1E",X"04",X"1E",
		X"09",X"0C",X"69",X"00",X"00",X"1B",X"16",X"1C",X"17",X"1A",X"72",X"20",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"04",X"03",X"01",X"01",X"03",X"04",X"06",X"07",X"08",X"07",X"05",X"02",X"04",X"06",X"08",
		X"09",X"0B",X"01",X"03",X"04",X"06",X"07",X"09",X"0A",X"0C",X"0D",X"0C",X"0A",X"08",X"07",X"05",
		X"03",X"01",X"02",X"04",X"05",X"04",X"02",X"01",X"03",X"05",X"06",X"08",X"07",X"05",X"03",X"02",
		X"04",X"06",X"08",X"0A",X"0B",X"0D",X"0B",X"09",X"07",X"05",X"01",X"02",X"03",X"02",X"02",X"01",
		X"04",X"06",X"07",X"08",X"06",X"04",X"01",X"02",X"04",X"06",X"08",X"0A",X"0C",X"0B",X"0A",X"05",
		X"02",X"03",X"07",X"09",X"0A",X"0C",X"0B",X"09",X"03",X"03",X"07",X"09",X"09",X"0B",X"0A",X"0A",
		X"0A",X"09",X"08",X"08",X"07",X"06",X"06",X"04",X"04",X"02",X"04",X"05",X"07",X"08",X"07",X"05",
		X"03",X"00",X"02",X"02",X"02",X"02",X"02",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"02",X"02",
		X"02",X"02",X"02",X"F8",X"F8",X"F8",X"F8",X"F8",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3E",X"FF",X"D3",X"C0",X"32",X"C5",X"E1",X"21",X"00",X"E1",X"36",X"00",X"54",X"5D",X"13",X"01",
		X"CF",X"00",X"ED",X"B0",X"3E",X"01",X"57",X"01",X"00",X"08",X"21",X"00",X"E0",X"7A",X"77",X"5E",
		X"BB",X"C2",X"BB",X"34",X"23",X"0B",X"79",X"B0",X"20",X"F3",X"7A",X"07",X"30",X"E8",X"16",X"55",
		X"7A",X"01",X"00",X"08",X"21",X"00",X"E0",X"77",X"23",X"3C",X"5F",X"0B",X"79",X"B0",X"28",X"09",
		X"7B",X"FE",X"AB",X"20",X"F2",X"3E",X"55",X"18",X"EE",X"7A",X"01",X"00",X"08",X"21",X"00",X"E0",
		X"BE",X"20",X"19",X"23",X"3C",X"5F",X"0B",X"79",X"B0",X"28",X"09",X"7B",X"FE",X"AB",X"20",X"F0",
		X"3E",X"55",X"18",X"EC",X"14",X"7A",X"FE",X"AB",X"20",X"C6",X"18",X"09",X"5E",X"57",X"AF",X"C3",
		X"BB",X"34",X"7A",X"18",X"DE",X"31",X"00",X"E8",X"3E",X"01",X"57",X"01",X"00",X"08",X"21",X"00",
		X"80",X"7A",X"77",X"5E",X"BB",X"28",X"08",X"CD",X"3B",X"35",X"CB",X"4F",X"CA",X"F5",X"33",X"23",
		X"0B",X"79",X"B0",X"20",X"EC",X"7A",X"07",X"30",X"E1",X"16",X"55",X"7A",X"01",X"00",X"08",X"21",
		X"00",X"80",X"77",X"23",X"3C",X"5F",X"0B",X"79",X"B0",X"28",X"09",X"7B",X"FE",X"AB",X"20",X"F2",
		X"3E",X"55",X"18",X"EE",X"7A",X"01",X"00",X"08",X"21",X"00",X"80",X"BE",X"20",X"19",X"23",X"3C",
		X"5F",X"0B",X"79",X"B0",X"28",X"09",X"7B",X"FE",X"AB",X"20",X"F0",X"3E",X"55",X"18",X"EC",X"14",
		X"7A",X"FE",X"AB",X"20",X"C6",X"18",X"0D",X"5E",X"57",X"CD",X"37",X"35",X"CB",X"4F",X"CA",X"F5",
		X"33",X"7A",X"18",X"DA",X"DD",X"21",X"EB",X"33",X"C3",X"B1",X"35",X"21",X"66",X"3A",X"DD",X"21",
		X"F5",X"33",X"C3",X"65",X"34",X"21",X"00",X"E1",X"36",X"00",X"54",X"5D",X"13",X"01",X"CF",X"00",
		X"ED",X"B0",X"21",X"00",X"00",X"AF",X"32",X"00",X"E7",X"06",X"00",X"0E",X"10",X"AF",X"AE",X"23",
		X"10",X"FC",X"0D",X"20",X"F9",X"E5",X"CD",X"35",X"34",X"E1",X"3A",X"00",X"E7",X"3C",X"FE",X"04",
		X"20",X"E4",X"AF",X"D3",X"1C",X"FB",X"3A",X"00",X"D0",X"CB",X"4F",X"20",X"F9",X"3E",X"03",X"32",
		X"01",X"E7",X"C3",X"CD",X"35",X"F5",X"FE",X"FF",X"28",X"02",X"0E",X"08",X"21",X"86",X"3A",X"09",
		X"EB",X"3A",X"00",X"E7",X"0F",X"0F",X"4F",X"21",X"C4",X"80",X"09",X"E5",X"EB",X"0E",X"08",X"ED",
		X"B0",X"13",X"13",X"D5",X"FD",X"E1",X"DD",X"E1",X"F1",X"CD",X"9A",X"34",X"3A",X"00",X"E7",X"C6",
		X"30",X"DD",X"77",X"03",X"C9",X"7E",X"23",X"FE",X"00",X"28",X"0B",X"5E",X"23",X"56",X"23",X"4F",
		X"06",X"00",X"ED",X"B0",X"18",X"EF",X"DD",X"E9",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"C6",X"30",
		X"FE",X"3A",X"38",X"02",X"C6",X"07",X"FD",X"77",X"00",X"DD",X"E9",X"E6",X"0F",X"C6",X"30",X"FE",
		X"3A",X"38",X"02",X"C6",X"07",X"FD",X"77",X"01",X"DD",X"E9",X"F5",X"0F",X"0F",X"0F",X"0F",X"E6",
		X"0F",X"C6",X"30",X"FE",X"3A",X"38",X"02",X"C6",X"07",X"FD",X"77",X"00",X"F1",X"E6",X"0F",X"C6",
		X"30",X"FE",X"3A",X"38",X"02",X"C6",X"07",X"FD",X"77",X"01",X"C9",X"08",X"D9",X"DD",X"21",X"C4",
		X"34",X"C3",X"B1",X"35",X"21",X"72",X"3A",X"DD",X"21",X"CE",X"34",X"C3",X"65",X"34",X"D9",X"FD",
		X"21",X"8F",X"80",X"DD",X"21",X"DB",X"34",X"7C",X"C3",X"78",X"34",X"DD",X"21",X"E3",X"34",X"7C",
		X"C3",X"8B",X"34",X"FD",X"23",X"FD",X"23",X"DD",X"21",X"EF",X"34",X"7D",X"C3",X"78",X"34",X"DD",
		X"21",X"F7",X"34",X"7D",X"C3",X"8B",X"34",X"FD",X"21",X"95",X"80",X"DD",X"21",X"03",X"35",X"7A",
		X"C3",X"78",X"34",X"DD",X"21",X"0B",X"35",X"7A",X"C3",X"8B",X"34",X"FD",X"21",X"99",X"80",X"DD",
		X"21",X"17",X"35",X"7B",X"C3",X"78",X"34",X"7B",X"DD",X"21",X"1F",X"35",X"C3",X"8B",X"34",X"3A",
		X"00",X"D0",X"CB",X"47",X"CA",X"2F",X"35",X"CB",X"4F",X"20",X"F4",X"08",X"C3",X"F5",X"33",X"08",
		X"B7",X"CA",X"72",X"33",X"C3",X"24",X"33",X"E5",X"D9",X"18",X"09",X"E5",X"D9",X"DD",X"21",X"44",
		X"35",X"C3",X"B1",X"35",X"21",X"00",X"80",X"11",X"00",X"E0",X"01",X"A0",X"04",X"ED",X"B0",X"21",
		X"00",X"80",X"36",X"00",X"54",X"5D",X"13",X"01",X"9F",X"04",X"ED",X"B0",X"21",X"72",X"3A",X"DD",
		X"21",X"66",X"35",X"C3",X"65",X"34",X"D9",X"FD",X"21",X"8F",X"80",X"7C",X"CD",X"9A",X"34",X"FD",
		X"23",X"FD",X"23",X"7D",X"CD",X"9A",X"34",X"FD",X"21",X"95",X"80",X"7A",X"CD",X"9A",X"34",X"FD",
		X"21",X"99",X"80",X"7B",X"CD",X"9A",X"34",X"E1",X"3A",X"00",X"D0",X"CB",X"47",X"28",X"06",X"CB",
		X"4F",X"28",X"10",X"18",X"F3",X"D9",X"21",X"00",X"E0",X"11",X"00",X"80",X"01",X"A0",X"04",X"ED",
		X"B0",X"D9",X"C9",X"21",X"A0",X"84",X"36",X"00",X"54",X"5D",X"13",X"01",X"5F",X"03",X"ED",X"B0",
		X"C9",X"21",X"00",X"84",X"01",X"FF",X"03",X"36",X"00",X"54",X"5D",X"13",X"ED",X"B0",X"21",X"00",
		X"80",X"01",X"FF",X"03",X"36",X"00",X"54",X"5D",X"13",X"ED",X"B0",X"DD",X"E9",X"CD",X"AD",X"38",
		X"21",X"BF",X"3E",X"CD",X"08",X"39",X"3A",X"01",X"E7",X"06",X"02",X"CD",X"1C",X"39",X"3A",X"00",
		X"D0",X"CB",X"47",X"20",X"14",X"3A",X"01",X"E7",X"07",X"4F",X"06",X"00",X"DD",X"21",X"96",X"3A",
		X"DD",X"09",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"E9",X"DD",X"21",X"02",X"E7",X"CD",X"DD",X"38",
		X"47",X"E6",X"55",X"FE",X"55",X"28",X"09",X"78",X"E6",X"AA",X"FE",X"AA",X"28",X"13",X"18",X"CE",
		X"DD",X"36",X"00",X"55",X"DD",X"36",X"01",X"08",X"DD",X"36",X"02",X"01",X"CD",X"32",X"36",X"18",
		X"BD",X"DD",X"36",X"00",X"AA",X"DD",X"36",X"01",X"03",X"DD",X"36",X"02",X"FF",X"CD",X"32",X"36",
		X"18",X"AC",X"DD",X"56",X"00",X"1E",X"02",X"CD",X"C8",X"38",X"28",X"0E",X"CD",X"4E",X"36",X"DD",
		X"56",X"00",X"1E",X"01",X"CD",X"C8",X"38",X"20",X"F3",X"C9",X"CD",X"4E",X"36",X"C9",X"3A",X"01",
		X"E7",X"DD",X"BE",X"01",X"C8",X"06",X"00",X"CD",X"1C",X"39",X"DD",X"86",X"02",X"32",X"01",X"E7",
		X"06",X"02",X"CD",X"1C",X"39",X"C9",X"CD",X"AD",X"38",X"21",X"10",X"3B",X"CD",X"08",X"39",X"3A",
		X"03",X"D0",X"21",X"CB",X"80",X"CD",X"B2",X"36",X"3A",X"04",X"D0",X"21",X"0B",X"81",X"CD",X"B2",
		X"36",X"DD",X"21",X"AC",X"3A",X"FD",X"21",X"A8",X"3A",X"3A",X"03",X"D0",X"EE",X"FF",X"06",X"02",
		X"CD",X"C6",X"36",X"DD",X"21",X"F8",X"3A",X"FD",X"21",X"F4",X"3A",X"3A",X"04",X"D0",X"EE",X"FF",
		X"06",X"01",X"CD",X"C5",X"36",X"CD",X"EC",X"36",X"3A",X"00",X"D0",X"CB",X"4F",X"20",X"C0",X"C3",
		X"CD",X"35",X"EE",X"FF",X"06",X"08",X"0F",X"38",X"04",X"36",X"30",X"18",X"02",X"36",X"31",X"23",
		X"23",X"10",X"F3",X"C9",X"0F",X"0F",X"4F",X"C5",X"DD",X"A6",X"00",X"DD",X"86",X"01",X"DD",X"23",
		X"DD",X"23",X"4F",X"06",X"00",X"FD",X"6E",X"00",X"FD",X"66",X"01",X"09",X"4E",X"FD",X"6E",X"02",
		X"FD",X"66",X"03",X"09",X"CD",X"11",X"39",X"C1",X"79",X"10",X"D9",X"C9",X"3A",X"04",X"D0",X"CB",
		X"57",X"CA",X"06",X"37",X"21",X"77",X"3B",X"CD",X"08",X"39",X"DD",X"21",X"99",X"3B",X"FD",X"21",
		X"9B",X"3B",X"06",X"01",X"18",X"10",X"21",X"7F",X"3C",X"CD",X"08",X"39",X"DD",X"21",X"92",X"3C",
		X"FD",X"21",X"96",X"3C",X"06",X"02",X"3A",X"03",X"D0",X"EE",X"FF",X"0F",X"0F",X"CD",X"C4",X"36",
		X"C9",X"AF",X"32",X"0F",X"E7",X"67",X"6F",X"22",X"0D",X"E7",X"CD",X"AD",X"38",X"21",X"22",X"3D",
		X"CD",X"08",X"39",X"3A",X"00",X"D0",X"21",X"CB",X"80",X"CD",X"B2",X"36",X"3A",X"01",X"D0",X"21",
		X"0B",X"81",X"CD",X"B2",X"36",X"3A",X"02",X"D0",X"21",X"4B",X"81",X"CD",X"B2",X"36",X"CD",X"8C",
		X"37",X"3A",X"0D",X"E7",X"21",X"8C",X"81",X"CD",X"7A",X"37",X"23",X"3A",X"0E",X"E7",X"CD",X"7A",
		X"37",X"3A",X"00",X"D0",X"CB",X"4F",X"20",X"CB",X"3A",X"01",X"D0",X"CB",X"4F",X"20",X"C4",X"CD",
		X"AD",X"38",X"3E",X"01",X"CD",X"3C",X"39",X"C3",X"CD",X"35",X"F5",X"0F",X"0F",X"0F",X"0F",X"E6",
		X"0F",X"C6",X"30",X"77",X"23",X"F1",X"E6",X"0F",X"C6",X"30",X"77",X"C9",X"21",X"0F",X"E7",X"3A",
		X"4E",X"E0",X"E6",X"C0",X"BE",X"C8",X"32",X"0F",X"E7",X"3A",X"0E",X"E7",X"C6",X"01",X"27",X"32",
		X"0E",X"E7",X"D0",X"3A",X"0D",X"E7",X"C6",X"01",X"27",X"32",X"0D",X"E7",X"C9",X"2A",X"53",X"3D",
		X"22",X"06",X"E7",X"21",X"68",X"3D",X"FD",X"21",X"57",X"3D",X"CD",X"C0",X"37",X"C3",X"CD",X"35",
		X"FD",X"22",X"0B",X"E7",X"E5",X"CD",X"AD",X"38",X"E1",X"CD",X"08",X"39",X"DD",X"21",X"08",X"E7",
		X"3E",X"01",X"32",X"05",X"E7",X"06",X"02",X"CD",X"23",X"39",X"3E",X"01",X"0E",X"40",X"CD",X"3E",
		X"39",X"CD",X"72",X"38",X"CD",X"7D",X"38",X"3E",X"FF",X"32",X"11",X"E7",X"3A",X"00",X"D0",X"CB",
		X"4F",X"28",X"4A",X"CD",X"F2",X"38",X"E6",X"AA",X"FE",X"2A",X"28",X"13",X"CD",X"DD",X"38",X"47",
		X"E6",X"55",X"FE",X"55",X"28",X"11",X"78",X"E6",X"AA",X"FE",X"AA",X"28",X"1D",X"18",X"DD",X"CD",
		X"72",X"38",X"CD",X"7D",X"38",X"18",X"D5",X"DD",X"36",X"00",X"55",X"3A",X"06",X"E7",X"DD",X"77",
		X"01",X"DD",X"36",X"02",X"01",X"CD",X"4F",X"38",X"18",X"C2",X"DD",X"36",X"00",X"AA",X"3A",X"07",
		X"E7",X"DD",X"77",X"01",X"DD",X"36",X"02",X"FF",X"CD",X"4F",X"38",X"18",X"AF",X"CD",X"72",X"38",
		X"3E",X"01",X"0E",X"20",X"CD",X"3E",X"39",X"3A",X"00",X"D0",X"CB",X"4F",X"20",X"9E",X"C9",X"CD",
		X"72",X"38",X"DD",X"56",X"00",X"1E",X"02",X"CD",X"C8",X"38",X"28",X"0F",X"CD",X"95",X"38",X"DD",
		X"56",X"00",X"1E",X"01",X"CD",X"C8",X"38",X"20",X"F3",X"18",X"03",X"CD",X"95",X"38",X"CD",X"7D",
		X"38",X"C9",X"3E",X"00",X"32",X"00",X"D0",X"CB",X"FF",X"32",X"00",X"D0",X"C9",X"3A",X"05",X"E7",
		X"4F",X"06",X"00",X"FD",X"2A",X"0B",X"E7",X"FD",X"09",X"FD",X"7E",X"00",X"32",X"00",X"D0",X"CB",
		X"FF",X"32",X"00",X"D0",X"C9",X"3A",X"05",X"E7",X"DD",X"BE",X"01",X"C8",X"06",X"00",X"CD",X"23",
		X"39",X"DD",X"86",X"02",X"32",X"05",X"E7",X"06",X"02",X"CD",X"23",X"39",X"C9",X"21",X"00",X"80",
		X"01",X"FF",X"03",X"36",X"00",X"54",X"5D",X"13",X"ED",X"B0",X"21",X"00",X"84",X"01",X"FF",X"03",
		X"36",X"00",X"54",X"5D",X"13",X"ED",X"B0",X"C9",X"0E",X"00",X"06",X"0C",X"CD",X"E2",X"38",X"A2",
		X"C8",X"10",X"F9",X"0D",X"20",X"F4",X"1D",X"20",X"EF",X"3E",X"FF",X"A2",X"C9",X"CD",X"E2",X"38",
		X"18",X"1F",X"21",X"10",X"E7",X"3A",X"01",X"D0",X"1F",X"CB",X"16",X"1F",X"CB",X"16",X"7E",X"EE",
		X"FF",X"C9",X"21",X"11",X"E7",X"3A",X"00",X"D0",X"1F",X"CB",X"16",X"1F",X"CB",X"16",X"7E",X"EE",
		X"FF",X"F5",X"AF",X"3D",X"20",X"FD",X"F1",X"C9",X"7E",X"FE",X"00",X"C8",X"CD",X"11",X"39",X"18",
		X"F7",X"4E",X"06",X"00",X"23",X"5E",X"23",X"56",X"23",X"ED",X"B0",X"C9",X"4F",X"D6",X"03",X"07",
		X"3C",X"18",X"01",X"4F",X"C5",X"0E",X"64",X"06",X"00",X"60",X"07",X"07",X"07",X"6F",X"29",X"29",
		X"09",X"EB",X"21",X"00",X"84",X"19",X"C1",X"70",X"23",X"70",X"79",X"C9",X"0E",X"00",X"06",X"00",
		X"10",X"FE",X"0D",X"20",X"F9",X"3D",X"20",X"F4",X"C9",X"C5",X"0E",X"00",X"06",X"00",X"10",X"FE",
		X"F5",X"3A",X"00",X"D0",X"CB",X"4F",X"28",X"09",X"F1",X"0D",X"20",X"F0",X"3D",X"20",X"EB",X"C1",
		X"C9",X"F1",X"C1",X"06",X"01",X"C9",X"CD",X"AD",X"38",X"11",X"00",X"E1",X"21",X"6D",X"3E",X"01",
		X"10",X"00",X"ED",X"B0",X"11",X"60",X"E1",X"21",X"7D",X"3E",X"01",X"10",X"00",X"ED",X"B0",X"3A",
		X"00",X"D0",X"CB",X"4F",X"20",X"F9",X"21",X"00",X"E1",X"36",X"00",X"54",X"5D",X"13",X"01",X"BF",
		X"00",X"ED",X"B0",X"C3",X"CD",X"35",X"3E",X"01",X"32",X"12",X"E7",X"AF",X"32",X"11",X"E7",X"18",
		X"2A",X"3A",X"00",X"D0",X"CB",X"4F",X"CA",X"CD",X"35",X"CD",X"F2",X"38",X"E6",X"AA",X"FE",X"2A",
		X"20",X"EF",X"3A",X"12",X"E7",X"3C",X"32",X"12",X"E7",X"FE",X"01",X"28",X"0E",X"FE",X"02",X"CA",
		X"E8",X"39",X"FE",X"03",X"CA",X"13",X"3A",X"D6",X"03",X"18",X"EB",X"CD",X"AD",X"38",X"21",X"1C",
		X"81",X"06",X"1A",X"3E",X"5A",X"77",X"2B",X"3D",X"10",X"FB",X"21",X"0C",X"82",X"06",X"0A",X"3E",
		X"39",X"77",X"2B",X"3D",X"10",X"FB",X"18",X"B9",X"CD",X"BA",X"38",X"21",X"20",X"80",X"36",X"F3",
		X"54",X"5D",X"13",X"01",X"BF",X"03",X"ED",X"B0",X"21",X"8D",X"3E",X"06",X"0A",X"C5",X"5E",X"23",
		X"56",X"23",X"46",X"23",X"4E",X"23",X"7E",X"23",X"EB",X"CD",X"23",X"3A",X"EB",X"C1",X"10",X"ED",
		X"C3",X"A1",X"39",X"21",X"20",X"84",X"36",X"0C",X"54",X"5D",X"13",X"01",X"BF",X"03",X"ED",X"B0",
		X"C3",X"A1",X"39",X"C5",X"E5",X"77",X"23",X"10",X"FC",X"E1",X"0E",X"20",X"09",X"C1",X"0D",X"20",
		X"F2",X"C9",X"CD",X"AD",X"38",X"21",X"20",X"80",X"0E",X"1E",X"06",X"0F",X"C5",X"06",X"00",X"36",
		X"94",X"54",X"5D",X"23",X"36",X"93",X"23",X"EB",X"ED",X"B0",X"EB",X"0E",X"1E",X"36",X"96",X"54",
		X"5D",X"23",X"36",X"95",X"23",X"EB",X"ED",X"B0",X"EB",X"C1",X"10",X"E0",X"3A",X"00",X"D0",X"CB",
		X"4F",X"20",X"F9",X"C3",X"CD",X"35",X"08",X"84",X"80",X"52",X"41",X"4D",X"00",X"00",X"00",X"4F",
		X"4B",X"00",X"10",X"84",X"80",X"52",X"41",X"4D",X"00",X"00",X"00",X"4E",X"47",X"00",X"00",X"5D",
		X"00",X"00",X"00",X"00",X"5D",X"00",X"52",X"4F",X"4D",X"00",X"00",X"00",X"4F",X"4B",X"52",X"4F",
		X"4D",X"00",X"00",X"00",X"4E",X"47",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"36",X"21",X"37",
		X"AD",X"37",X"66",X"39",X"96",X"39",X"32",X"3A",X"B0",X"3A",X"B8",X"3A",X"03",X"00",X"03",X"04",
		X"00",X"04",X"08",X"0C",X"10",X"1B",X"26",X"31",X"01",X"73",X"81",X"35",X"01",X"73",X"81",X"33",
		X"01",X"73",X"81",X"32",X"01",X"73",X"81",X"31",X"08",X"ED",X"81",X"31",X"30",X"00",X"33",X"30",
		X"00",X"35",X"30",X"08",X"ED",X"81",X"32",X"30",X"00",X"34",X"30",X"00",X"36",X"30",X"08",X"ED",
		X"81",X"00",X"00",X"00",X"00",X"00",X"00",X"31",X"30",X"08",X"ED",X"81",X"00",X"00",X"00",X"00",
		X"00",X"00",X"4E",X"4F",X"FA",X"3A",X"FC",X"3A",X"01",X"00",X"00",X"0A",X"07",X"B1",X"82",X"54",
		X"41",X"42",X"4C",X"45",X"00",X"00",X"07",X"B1",X"82",X"55",X"50",X"52",X"49",X"47",X"48",X"54",
		X"16",X"84",X"80",X"44",X"49",X"50",X"00",X"53",X"57",X"00",X"31",X"00",X"32",X"00",X"33",X"00",
		X"34",X"00",X"35",X"00",X"36",X"00",X"37",X"00",X"38",X"03",X"C6",X"80",X"53",X"57",X"31",X"03",
		X"06",X"81",X"53",X"57",X"32",X"0B",X"64",X"81",X"50",X"41",X"54",X"52",X"4F",X"4C",X"00",X"43",
		X"41",X"52",X"53",X"0D",X"A4",X"81",X"45",X"58",X"54",X"45",X"4E",X"44",X"00",X"50",X"4F",X"49",
		X"4E",X"54",X"53",X"08",X"F6",X"81",X"54",X"48",X"4F",X"55",X"53",X"41",X"4E",X"44",X"09",X"24",
		X"82",X"43",X"4F",X"49",X"4E",X"00",X"4D",X"4F",X"44",X"45",X"09",X"A4",X"82",X"42",X"4F",X"44",
		X"59",X"00",X"54",X"59",X"50",X"45",X"00",X"01",X"2E",X"82",X"00",X"1A",X"64",X"82",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"9F",X"3B",X"AF",X"3B",X"00",
		X"10",X"20",X"30",X"40",X"50",X"60",X"60",X"70",X"80",X"90",X"A0",X"B0",X"60",X"60",X"C0",X"0D",
		X"31",X"82",X"31",X"43",X"4F",X"49",X"4E",X"00",X"00",X"31",X"50",X"4C",X"41",X"59",X"00",X"0D",
		X"31",X"82",X"32",X"43",X"4F",X"49",X"4E",X"53",X"00",X"31",X"50",X"4C",X"41",X"59",X"00",X"0D",
		X"31",X"82",X"33",X"43",X"4F",X"49",X"4E",X"53",X"00",X"31",X"50",X"4C",X"41",X"59",X"00",X"0D",
		X"31",X"82",X"34",X"43",X"4F",X"49",X"4E",X"53",X"00",X"31",X"50",X"4C",X"41",X"59",X"00",X"0D",
		X"31",X"82",X"35",X"43",X"4F",X"49",X"4E",X"53",X"00",X"31",X"50",X"4C",X"41",X"59",X"00",X"0D",
		X"31",X"82",X"36",X"43",X"4F",X"49",X"4E",X"53",X"00",X"31",X"50",X"4C",X"41",X"59",X"00",X"0D",
		X"31",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",
		X"31",X"82",X"31",X"43",X"4F",X"49",X"4E",X"00",X"00",X"32",X"50",X"4C",X"41",X"59",X"53",X"0D",
		X"31",X"82",X"31",X"43",X"4F",X"49",X"4E",X"00",X"00",X"33",X"50",X"4C",X"41",X"59",X"53",X"0D",
		X"31",X"82",X"31",X"43",X"4F",X"49",X"4E",X"00",X"00",X"34",X"50",X"4C",X"41",X"59",X"53",X"0D",
		X"31",X"82",X"31",X"43",X"4F",X"49",X"4E",X"00",X"00",X"35",X"50",X"4C",X"41",X"59",X"53",X"0D",
		X"31",X"82",X"31",X"43",X"4F",X"49",X"4E",X"00",X"00",X"36",X"50",X"4C",X"41",X"59",X"53",X"0D",
		X"31",X"82",X"00",X"46",X"52",X"45",X"45",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"2E",X"82",X"41",X"0B",X"64",X"82",X"43",X"4F",X"49",X"4E",X"00",X"4D",X"4F",X"44",X"45",X"00",
		X"42",X"00",X"03",X"00",X"03",X"04",X"9A",X"3C",X"A2",X"3C",X"00",X"10",X"20",X"30",X"40",X"50",
		X"60",X"70",X"0D",X"31",X"82",X"31",X"43",X"4F",X"49",X"4E",X"00",X"00",X"31",X"50",X"4C",X"41",
		X"59",X"00",X"0D",X"31",X"82",X"32",X"43",X"4F",X"49",X"4E",X"53",X"00",X"31",X"50",X"4C",X"41",
		X"59",X"00",X"0D",X"31",X"82",X"33",X"43",X"4F",X"49",X"4E",X"53",X"00",X"31",X"50",X"4C",X"41",
		X"59",X"00",X"0D",X"31",X"82",X"00",X"46",X"52",X"45",X"45",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0D",X"71",X"82",X"31",X"43",X"4F",X"49",X"4E",X"00",X"00",X"32",X"50",X"4C",X"41",
		X"59",X"53",X"0D",X"71",X"82",X"31",X"43",X"4F",X"49",X"4E",X"00",X"00",X"33",X"50",X"4C",X"41",
		X"59",X"53",X"0D",X"71",X"82",X"31",X"43",X"4F",X"49",X"4E",X"00",X"00",X"35",X"50",X"4C",X"41",
		X"59",X"53",X"0D",X"71",X"82",X"31",X"43",X"4F",X"49",X"4E",X"00",X"00",X"36",X"50",X"4C",X"41",
		X"59",X"53",X"0F",X"8B",X"80",X"31",X"00",X"32",X"00",X"33",X"00",X"34",X"00",X"35",X"00",X"36",
		X"00",X"37",X"00",X"38",X"04",X"C4",X"80",X"4B",X"45",X"59",X"30",X"04",X"04",X"81",X"4B",X"45",
		X"59",X"31",X"04",X"44",X"81",X"4B",X"45",X"59",X"32",X"06",X"84",X"81",X"54",X"49",X"4D",X"49",
		X"4E",X"47",X"00",X"0E",X"01",X"00",X"00",X"00",X"01",X"10",X"11",X"12",X"13",X"14",X"16",X"17",
		X"18",X"1B",X"1C",X"1D",X"1E",X"1F",X"00",X"00",X"0B",X"27",X"80",X"53",X"00",X"4F",X"00",X"55",
		X"00",X"4E",X"00",X"44",X"00",X"53",X"0E",X"44",X"81",X"30",X"37",X"00",X"53",X"50",X"41",X"43",
		X"45",X"00",X"50",X"4C",X"41",X"4E",X"54",X"0D",X"64",X"81",X"30",X"38",X"00",X"55",X"46",X"4F",
		X"00",X"46",X"4C",X"59",X"49",X"4E",X"47",X"0C",X"84",X"80",X"30",X"31",X"00",X"45",X"58",X"50",
		X"4C",X"4F",X"53",X"49",X"4F",X"4E",X"0E",X"E4",X"80",X"30",X"34",X"00",X"43",X"41",X"52",X"00",
		X"4D",X"49",X"53",X"53",X"49",X"4C",X"45",X"10",X"C4",X"80",X"30",X"33",X"00",X"55",X"46",X"4F",
		X"00",X"45",X"58",X"50",X"4C",X"4F",X"53",X"49",X"4F",X"4E",X"10",X"A4",X"80",X"30",X"32",X"00",
		X"50",X"4F",X"49",X"4E",X"54",X"00",X"50",X"41",X"53",X"53",X"41",X"47",X"45",X"07",X"04",X"81",
		X"30",X"35",X"00",X"43",X"4F",X"49",X"4E",X"0B",X"24",X"81",X"30",X"36",X"00",X"43",X"41",X"52",
		X"00",X"4A",X"55",X"4D",X"50",X"14",X"84",X"81",X"30",X"39",X"00",X"42",X"41",X"43",X"4B",X"00",
		X"47",X"52",X"4F",X"55",X"4E",X"44",X"00",X"4D",X"55",X"53",X"49",X"43",X"0F",X"A4",X"81",X"31",
		X"30",X"00",X"45",X"4E",X"44",X"49",X"4E",X"47",X"00",X"4D",X"55",X"53",X"49",X"43",X"10",X"C4",
		X"81",X"31",X"31",X"00",X"4F",X"50",X"45",X"4E",X"49",X"4E",X"47",X"00",X"4D",X"55",X"53",X"49",
		X"43",X"0F",X"E4",X"81",X"31",X"32",X"00",X"53",X"54",X"45",X"50",X"00",X"50",X"41",X"53",X"53",
		X"41",X"47",X"45",X"11",X"04",X"82",X"31",X"33",X"00",X"43",X"4F",X"4E",X"47",X"52",X"41",X"54",
		X"55",X"4C",X"41",X"54",X"49",X"4F",X"4E",X"10",X"24",X"82",X"31",X"34",X"00",X"43",X"41",X"52",
		X"00",X"45",X"58",X"50",X"4C",X"4F",X"53",X"49",X"4F",X"4E",X"00",X"00",X"00",X"A8",X"01",X"38",
		X"60",X"A8",X"41",X"38",X"98",X"90",X"81",X"38",X"60",X"90",X"C1",X"38",X"98",X"68",X"01",X"38",
		X"60",X"68",X"41",X"38",X"98",X"50",X"81",X"38",X"60",X"50",X"C1",X"38",X"98",X"20",X"84",X"20",
		X"07",X"00",X"00",X"87",X"20",X"07",X"08",X"00",X"85",X"20",X"08",X"02",X"00",X"86",X"05",X"08",
		X"05",X"05",X"86",X"04",X"08",X"0C",X"09",X"86",X"05",X"08",X"06",X"0E",X"86",X"04",X"08",X"04",
		X"12",X"86",X"05",X"08",X"03",X"17",X"86",X"04",X"08",X"00",X"1B",X"86",X"05",X"08",X"08",X"0E",
		X"84",X"80",X"30",X"31",X"00",X"00",X"44",X"49",X"50",X"00",X"53",X"57",X"49",X"54",X"43",X"48",
		X"0C",X"C4",X"80",X"30",X"32",X"00",X"00",X"49",X"3F",X"4F",X"00",X"50",X"4F",X"52",X"54",X"0A",
		X"04",X"81",X"30",X"33",X"00",X"00",X"53",X"4F",X"55",X"4E",X"44",X"53",X"0D",X"44",X"81",X"30",
		X"34",X"00",X"00",X"43",X"48",X"41",X"52",X"41",X"43",X"54",X"45",X"52",X"09",X"84",X"81",X"30",
		X"35",X"00",X"00",X"43",X"4F",X"4C",X"4F",X"52",X"0F",X"C4",X"81",X"30",X"36",X"00",X"00",X"42",
		X"45",X"41",X"4D",X"00",X"41",X"44",X"4A",X"55",X"53",X"54",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
