library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity travusa_chr_bit1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of travusa_chr_bit1 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"3F",X"60",X"40",X"40",X"40",X"40",X"40",X"00",X"FC",X"06",X"02",X"02",X"02",X"02",X"02",
		X"40",X"40",X"40",X"40",X"40",X"60",X"3F",X"00",X"02",X"02",X"02",X"02",X"02",X"06",X"FC",X"00",
		X"77",X"67",X"6D",X"7D",X"7B",X"3F",X"1E",X"00",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",
		X"38",X"7D",X"7D",X"6D",X"6F",X"6F",X"67",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"00",X"00",
		X"7F",X"3F",X"00",X"1C",X"3E",X"77",X"63",X"63",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"7F",X"00",X"00",X"00",X"00",X"18",X"3B",X"F8",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"7F",X"7F",X"60",X"60",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"10",X"82",X"22",X"A1",X"04",X"46",X"00",X"C9",X"00",X"64",X"01",X"00",X"48",X"90",X"82",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"FE",X"FF",X"7F",X"9F",X"5F",X"3F",X"0F",X"3F",X"0F",X"57",X"42",X"00",X"24",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"7F",X"1F",X"A7",X"09",X"0F",X"17",X"03",X"09",X"42",X"00",X"00",X"84",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C3",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C3",
		X"50",X"0A",X"00",X"88",X"A4",X"14",X"BE",X"DF",X"FC",X"FE",X"FF",X"7F",X"7F",X"3F",X"4F",X"17",
		X"07",X"0F",X"21",X"04",X"91",X"21",X"00",X"08",X"4B",X"F4",X"BA",X"F6",X"3F",X"52",X"3E",X"7F",
		X"BF",X"EA",X"54",X"83",X"28",X"C1",X"06",X"A0",X"FF",X"A6",X"50",X"24",X"54",X"08",X"A2",X"44",
		X"FF",X"FF",X"7F",X"FF",X"FF",X"7F",X"7F",X"FF",X"0F",X"2F",X"03",X"0A",X"03",X"40",X"01",X"00",
		X"84",X"00",X"09",X"40",X"00",X"24",X"46",X"00",X"00",X"02",X"80",X"48",X"00",X"00",X"44",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"7F",X"7F",X"3F",X"3F",X"03",
		X"80",X"C0",X"C0",X"C0",X"E0",X"E0",X"F0",X"F0",X"DF",X"1F",X"6F",X"4F",X"87",X"77",X"4F",X"67",
		X"FE",X"FE",X"7F",X"3F",X"BF",X"3F",X"5F",X"1F",X"FA",X"E0",X"A8",X"01",X"82",X"00",X"20",X"04",
		X"9D",X"73",X"84",X"94",X"64",X"89",X"20",X"12",X"DD",X"A5",X"B0",X"C6",X"09",X"5A",X"22",X"85",
		X"FB",X"2D",X"DA",X"2B",X"D6",X"D5",X"77",X"22",X"F5",X"A5",X"3A",X"9C",X"A5",X"5E",X"E0",X"04",
		X"BB",X"E5",X"29",X"7C",X"D6",X"8F",X"6A",X"79",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",
		X"81",X"C4",X"E0",X"F8",X"FE",X"FF",X"FF",X"FF",X"00",X"80",X"02",X"50",X"44",X"84",X"E0",X"F8",
		X"AE",X"49",X"BD",X"26",X"6A",X"B9",X"0E",X"6F",X"7F",X"3F",X"9F",X"DF",X"7F",X"CF",X"47",X"77",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"07",X"CB",X"93",X"3F",X"E7",X"2D",X"79",X"C4",X"16",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"FF",X"3F",X"7F",X"9F",X"DF",X"0F",X"5F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"07",X"07",X"07",X"07",X"07",X"00",X"00",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"00",X"00",X"00",X"00",X"07",X"07",X"07",X"07",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"E0",X"E0",X"E0",X"E0",X"00",X"00",X"00",X"0D",X"7B",X"81",X"64",X"0E",X"30",X"4F",
		X"FF",X"00",X"18",X"3C",X"3C",X"18",X"00",X"FF",X"FF",X"80",X"80",X"80",X"80",X"80",X"80",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FC",X"F8",X"E0",X"80",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"F8",X"E0",X"80",X"00",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"DF",X"77",X"1A",X"07",X"00",X"00",
		X"07",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FC",X"F8",X"E0",X"80",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"F8",X"E0",X"80",X"00",X"00",X"00",X"00",
		X"37",X"67",X"9B",X"D3",X"3F",X"7B",X"51",X"11",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"F8",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E7",X"2A",X"9F",X"D5",X"F0",X"E2",X"FC",X"C2",
		X"F9",X"FB",X"FE",X"FC",X"FF",X"FF",X"FF",X"FF",X"08",X"03",X"03",X"83",X"C1",X"E0",X"F0",X"F8",
		X"FF",X"01",X"61",X"F1",X"F1",X"61",X"01",X"FF",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"88",X"8A",X"DF",X"F9",X"CB",X"DE",X"E4",X"F7",X"FB",X"F8",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"DB",X"85",X"48",X"20",X"90",X"E6",X"E2",X"E0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FD",X"FF",X"FE",X"FE",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FC",X"F8",X"E0",X"80",X"FF",X"E3",X"83",X"03",X"03",X"03",X"03",X"03",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"F8",
		X"FF",X"FC",X"F8",X"E0",X"80",X"00",X"00",X"00",X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"FF",X"FF",X"FF",X"FC",X"F8",X"E0",X"80",X"00",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"7F",X"7F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"01",X"07",X"1F",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"FC",X"FE",X"7F",X"7F",X"3F",X"4F",X"17",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"E0",X"E0",X"80",X"40",X"80",X"00",
		X"07",X"0D",X"07",X"03",X"03",X"01",X"01",X"00",X"C0",X"C0",X"E0",X"E0",X"60",X"70",X"F0",X"70",
		X"07",X"07",X"07",X"07",X"0F",X"0F",X"05",X"07",X"C0",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",
		X"03",X"00",X"00",X"00",X"01",X"03",X"03",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"07",X"07",X"07",X"03",X"03",X"01",X"00",X"80",X"C0",X"E0",X"E0",X"C0",X"C0",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"C3",X"00",X"00",X"00",X"00",X"00",X"00",X"FB",X"C2",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"4C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"E0",X"F0",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",X"F0",X"FC",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"F0",X"F8",X"FC",X"FF",X"7F",X"5F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"F0",X"00",X"00",X"C0",X"F8",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"80",X"F8",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"F0",X"C0",X"06",X"9E",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"03",
		X"FF",X"FF",X"FF",X"FF",X"0F",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"01",X"00",X"00",X"00",X"FE",
		X"FF",X"FF",X"FF",X"FF",X"7F",X"1F",X"0F",X"03",X"7F",X"1F",X"07",X"01",X"80",X"E0",X"F8",X"FE",
		X"00",X"00",X"E0",X"FC",X"FF",X"FF",X"1F",X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",
		X"FF",X"7F",X"3F",X"0F",X"07",X"81",X"C0",X"F0",X"7F",X"3F",X"1F",X"8F",X"C7",X"E3",X"F1",X"78",
		X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"0F",X"07",X"1F",X"0F",X"03",X"81",X"E0",X"F0",X"FC",X"7E",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"03",X"00",X"FF",X"7F",X"1F",X"07",X"01",X"80",X"E0",X"F8",
		X"7F",X"00",X"00",X"00",X"80",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"E0",X"FF",X"FF",X"FF",X"1F",
		X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"C0",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",
		X"00",X"00",X"0F",X"FF",X"FF",X"FF",X"F0",X"00",X"F0",X"00",X"00",X"00",X"0F",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"F0",X"00",X"00",X"00",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",X"00",X"00",
		X"FF",X"FF",X"F8",X"C0",X"00",X"00",X"07",X"3F",X"FF",X"FF",X"FF",X"FF",X"FE",X"F0",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"C0",X"00",X"00",X"07",X"3F",X"FF",X"FF",X"FF",
		X"FF",X"FE",X"F0",X"00",X"00",X"01",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"C0",X"00",X"00",
		X"00",X"3F",X"FF",X"FF",X"FF",X"C0",X"00",X"00",X"00",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"FF",X"FF",X"FF",X"F0",X"00",X"00",X"00",
		X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"C0",X"00",X"00",X"07",X"3F",
		X"01",X"0F",X"FF",X"FF",X"FE",X"F0",X"00",X"00",X"01",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"00",X"00",X"07",X"3F",X"FF",X"FF",X"FF",X"FF",X"F0",X"80",X"00",X"00",X"0F",X"7F",X"FF",
		X"00",X"00",X"03",X"1F",X"FF",X"FF",X"FC",X"E0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"E0",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"7F",X"01",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"3F",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FC",X"7E",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C0",X"E0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F9",X"FF",X"FF",X"7F",X"1F",X"0F",X"07",X"03",X"81",
		X"C7",X"E1",X"F0",X"F8",X"FC",X"7E",X"3F",X"1F",X"0F",X"07",X"03",X"81",X"C0",X"E0",X"F0",X"F8",
		X"FC",X"7E",X"3F",X"1F",X"0F",X"07",X"03",X"01",X"FC",X"FC",X"FC",X"FC",X"FC",X"FE",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"9F",
		X"CF",X"E7",X"F3",X"F9",X"FC",X"7E",X"3F",X"1F",X"C0",X"E0",X"F0",X"F8",X"FC",X"7E",X"3F",X"1F",
		X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"FF",X"FF",X"FD",X"FC",X"FC",X"FC",X"FC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"9F",
		X"FF",X"FF",X"FF",X"FB",X"FC",X"7E",X"3F",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"1F",X"FF",X"FF",X"7F",X"8F",X"C1",X"E0",X"F0",X"F8",
		X"FF",X"7F",X"3F",X"1F",X"0F",X"07",X"03",X"81",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C1",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"01",X"00",X"00",X"00",X"FC",X"FF",X"FF",X"07",X"83",X"83",X"C1",X"C1",X"E0",X"E0",X"F0",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"F1",X"11",X"11",X"11",X"1F",X"11",X"11",X"11",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"1F",X"1F",X"1F",X"1F",X"11",X"11",X"11",X"FF",X"1F",X"1F",X"1F",X"1F",X"11",X"11",X"11",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"10",X"10",X"10",X"1F",X"11",X"11",X"11",
		X"F0",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"FF",X"01",X"93",X"FF",X"01",X"9D",X"63",X"01",
		X"FD",X"03",X"FD",X"01",X"6D",X"93",X"FF",X"01",X"C3",X"E1",X"F0",X"F8",X"FC",X"DE",X"CF",X"C7",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"FF",X"F5",X"BF",X"FF",X"ED",X"FF",
		X"B9",X"F7",X"9D",X"32",X"EB",X"AE",X"76",X"DB",X"5C",X"89",X"A9",X"C6",X"2D",X"37",X"5F",X"FF",
		X"3F",X"96",X"69",X"D1",X"F4",X"D9",X"77",X"FF",X"F7",X"A1",X"D2",X"45",X"A8",X"14",X"7A",X"FF",
		X"FF",X"FE",X"D4",X"FA",X"A0",X"51",X"A2",X"08",X"FF",X"DF",X"16",X"AF",X"4D",X"1A",X"05",X"50",
		X"FF",X"7E",X"AE",X"54",X"29",X"88",X"22",X"49",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"42",X"25",X"56",X"AD",X"F7",X"DF",X"EF",X"20",X"52",X"24",X"53",X"BD",X"77",X"DF",X"FD",
		X"21",X"44",X"2A",X"B5",X"5B",X"BD",X"EB",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",
		X"10",X"BF",X"A0",X"A8",X"8F",X"BF",X"C0",X"FF",X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"40",X"60",
		X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"04",X"09",X"F1",X"01",X"07",X"FF",X"FD",X"03",X"FF",
		X"5A",X"48",X"7E",X"7E",X"40",X"7E",X"7E",X"64",X"7E",X"7E",X"7E",X"7E",X"00",X"00",X"24",X"66",
		X"66",X"66",X"66",X"18",X"66",X"66",X"66",X"66",X"6E",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"6E",
		X"FF",X"FF",X"D7",X"BD",X"D7",X"4B",X"81",X"00",X"38",X"D1",X"95",X"4B",X"DE",X"F7",X"FF",X"FF",
		X"AE",X"97",X"59",X"BB",X"27",X"D7",X"58",X"D0",X"EA",X"B0",X"41",X"2D",X"C8",X"0E",X"0C",X"05",
		X"34",X"C2",X"0A",X"40",X"48",X"84",X"A0",X"28",X"04",X"20",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"28",X"01",X"21",X"64",X"64",X"F6",X"F6",X"98",X"D4",X"DC",X"E9",X"EB",X"A2",X"23",X"23",
		X"A2",X"DA",X"C8",X"89",X"01",X"01",X"1B",X"FE",X"05",X"06",X"CA",X"FD",X"B6",X"2A",X"6B",X"9D",
		X"90",X"9C",X"8A",X"CA",X"C2",X"C0",X"C0",X"E9",X"00",X"08",X"8A",X"19",X"41",X"C5",X"EB",X"D3",
		X"3D",X"BC",X"F6",X"F2",X"4F",X"6A",X"D7",X"B5",X"D2",X"99",X"1C",X"14",X"40",X"C0",X"F0",X"BF",
		X"EB",X"6D",X"03",X"0A",X"1B",X"18",X"0D",X"1C",X"09",X"B2",X"56",X"5D",X"67",X"69",X"8A",X"22",
		X"2A",X"50",X"08",X"D8",X"91",X"54",X"50",X"26",X"22",X"54",X"BF",X"AC",X"E9",X"CA",X"93",X"6D",
		X"E0",X"DF",X"BF",X"7F",X"78",X"78",X"73",X"72",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"45",X"90",
		X"00",X"FF",X"FF",X"FF",X"00",X"00",X"94",X"22",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"A9",X"CA",
		X"07",X"FB",X"FD",X"FE",X"1E",X"0E",X"8E",X"CE",X"75",X"72",X"70",X"74",X"72",X"73",X"76",X"71",
		X"0E",X"CE",X"8E",X"8E",X"4E",X"0E",X"CE",X"4E",X"74",X"72",X"73",X"78",X"3F",X"9F",X"CF",X"E0",
		X"74",X"AA",X"D1",X"02",X"FF",X"FF",X"FF",X"00",X"33",X"D6",X"29",X"00",X"FF",X"FF",X"FF",X"00",
		X"2C",X"6A",X"D8",X"41",X"FF",X"FF",X"FF",X"00",X"CE",X"4E",X"8E",X"3E",X"FE",X"FD",X"FB",X"17",
		X"00",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"00",X"00",X"C3",X"C3",X"C3",X"C3",
		X"C0",X"9F",X"3E",X"7C",X"78",X"79",X"7B",X"7F",X"03",X"F9",X"7C",X"3E",X"1E",X"9E",X"DE",X"FE",
		X"EE",X"1A",X"81",X"38",X"9C",X"01",X"E3",X"10",X"AB",X"E4",X"B9",X"6E",X"4D",X"3B",X"8B",X"8E",
		X"89",X"02",X"05",X"41",X"46",X"82",X"00",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"33",X"49",X"98",X"55",X"8A",X"A9",X"15",X"68",X"98",X"1A",X"CD",X"23",X"10",X"98",X"B9",X"FD",
		X"4A",X"92",X"39",X"20",X"04",X"95",X"BF",X"FF",X"92",X"48",X"B1",X"56",X"08",X"01",X"43",X"EF",
		X"FF",X"FF",X"CF",X"A7",X"0A",X"15",X"42",X"E8",X"FF",X"FF",X"FF",X"FF",X"33",X"4D",X"84",X"53",
		X"FF",X"FD",X"FD",X"FD",X"94",X"2D",X"91",X"66",X"FF",X"FF",X"FF",X"DF",X"DF",X"DF",X"DF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"5A",X"B7",X"FE",X"F7",X"6F",X"BE",X"DF",X"ED",X"00",X"EF",X"EF",X"10",X"10",X"EF",X"EF",X"00",
		X"00",X"FC",X"FA",X"0E",X"16",X"C6",X"A6",X"66",X"66",X"24",X"00",X"00",X"7E",X"66",X"72",X"7A",
		X"7E",X"7E",X"40",X"7E",X"7E",X"72",X"5E",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"DA",X"92",X"DA",X"52",X"52",X"DA",X"00",X"00",X"CA",X"AA",X"CA",X"AA",X"AA",X"CE",X"00",
		X"00",X"A4",X"AA",X"AA",X"CA",X"AE",X"AA",X"00",X"00",X"A9",X"AA",X"AA",X"BA",X"AB",X"AA",X"00",
		X"00",X"3B",X"92",X"93",X"91",X"91",X"93",X"00",X"00",X"51",X"51",X"51",X"55",X"51",X"71",X"00",
		X"00",X"4B",X"6A",X"6A",X"5A",X"5A",X"4B",X"00",X"C0",X"FF",X"EF",X"E8",X"EE",X"EE",X"EE",X"FE",
		X"C1",X"FC",X"BE",X"BE",X"BE",X"8E",X"FE",X"FF",X"C0",X"FF",X"EF",X"E1",X"FC",X"FE",X"8F",X"FF",
		X"C1",X"FC",X"BE",X"BE",X"BE",X"BE",X"CF",X"FF",X"8F",X"EF",X"EF",X"EF",X"EF",X"EF",X"E0",X"FF",
		X"E3",X"FB",X"BB",X"39",X"39",X"39",X"BB",X"FF",X"81",X"FC",X"8E",X"BE",X"BE",X"BE",X"BE",X"FF",
		X"F1",X"11",X"11",X"11",X"1F",X"11",X"11",X"11",X"00",X"00",X"1C",X"FC",X"FC",X"E1",X"0A",X"51",
		X"FF",X"F0",X"80",X"00",X"0F",X"7F",X"FF",X"F0",X"F8",X"C0",X"00",X"07",X"3F",X"FF",X"FF",X"F8",
		X"11",X"B6",X"64",X"92",X"C0",X"4F",X"3F",X"FF",X"9A",X"28",X"81",X"0F",X"FF",X"FE",X"F0",X"00",
		X"07",X"3F",X"FF",X"F8",X"C0",X"00",X"07",X"3F",X"C3",X"C0",X"00",X"00",X"0F",X"FF",X"FF",X"FF",
		X"00",X"00",X"0F",X"FF",X"FF",X"FF",X"F0",X"00",X"89",X"6A",X"30",X"9B",X"C2",X"00",X"03",X"C3",
		X"88",X"9C",X"30",X"00",X"0F",X"FF",X"FF",X"F0",X"A4",X"20",X"0F",X"FF",X"FF",X"F0",X"00",X"00",
		X"0F",X"FF",X"FF",X"F0",X"00",X"00",X"0F",X"FF",X"FF",X"F0",X"00",X"00",X"0F",X"FF",X"FF",X"FF",
		X"00",X"00",X"0F",X"FF",X"FF",X"FF",X"F0",X"00",X"FF",X"0F",X"10",X"8A",X"D9",X"46",X"60",X"1A",
		X"CF",X"C3",X"C3",X"03",X"00",X"80",X"69",X"2D",X"C0",X"FF",X"FF",X"FF",X"3F",X"80",X"A1",X"1C",
		X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"11",X"FF",X"03",X"01",X"00",X"80",X"84",X"86",X"07",
		X"FF",X"3F",X"38",X"00",X"05",X"57",X"98",X"A2",X"F0",X"01",X"26",X"4C",X"66",X"28",X"A2",X"26",
		X"07",X"3F",X"FF",X"FF",X"F8",X"C0",X"00",X"07",X"FF",X"FE",X"F0",X"00",X"01",X"0F",X"FF",X"FE",
		X"C0",X"00",X"07",X"3F",X"FF",X"F8",X"C2",X"02",X"0F",X"FF",X"FE",X"F0",X"05",X"6A",X"4B",X"AC",
		X"F8",X"C1",X"07",X"29",X"D0",X"15",X"6C",X"49",X"01",X"0F",X"FF",X"FF",X"FE",X"F0",X"00",X"01",
		X"FF",X"FF",X"F8",X"80",X"00",X"07",X"7F",X"FF",X"F0",X"00",X"00",X"03",X"C3",X"C3",X"C0",X"82",
		X"00",X"0F",X"FF",X"FF",X"F0",X"00",X"4C",X"84",X"FF",X"FF",X"F0",X"02",X"A5",X"B4",X"32",X"46",
		X"F0",X"02",X"08",X"24",X"20",X"90",X"C2",X"0C",X"0F",X"FF",X"FF",X"FF",X"F0",X"00",X"00",X"0F",
		X"FF",X"FF",X"F0",X"00",X"00",X"0F",X"FF",X"FF",X"F0",X"00",X"00",X"0F",X"FF",X"FF",X"F0",X"00",
		X"00",X"03",X"C3",X"C3",X"C0",X"02",X"42",X"C9",X"3F",X"FF",X"FF",X"C0",X"16",X"89",X"DA",X"22",
		X"FF",X"FF",X"00",X"45",X"42",X"90",X"CA",X"23",X"0C",X"00",X"00",X"61",X"11",X"58",X"B6",X"03",
		X"00",X"3F",X"FF",X"FF",X"FF",X"C0",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",
		X"FF",X"FF",X"FF",X"03",X"01",X"00",X"08",X"0C",X"9F",X"47",X"89",X"60",X"66",X"9A",X"C8",X"57",
		X"C0",X"FC",X"FF",X"3F",X"83",X"20",X"99",X"48",X"00",X"00",X"E0",X"FF",X"FF",X"1F",X"40",X"84",
		X"7F",X"00",X"00",X"80",X"C3",X"C3",X"43",X"00",X"B3",X"51",X"50",X"68",X"F5",X"F7",X"F6",X"2C",
		X"C1",X"E0",X"60",X"20",X"03",X"87",X"61",X"50",X"FE",X"7F",X"1F",X"07",X"81",X"E0",X"F8",X"7E",
		X"00",X"C0",X"FC",X"FF",X"FF",X"3F",X"03",X"00",X"0E",X"47",X"83",X"A1",X"14",X"50",X"C1",X"9A",
		X"1F",X"0F",X"83",X"E1",X"F0",X"7C",X"1E",X"4F",X"81",X"C0",X"F0",X"F8",X"7E",X"3F",X"0F",X"87",
		X"4E",X"46",X"60",X"C8",X"2C",X"9A",X"51",X"44",X"3C",X"1E",X"0F",X"07",X"63",X"71",X"38",X"DC",
		X"3F",X"8F",X"A7",X"11",X"D0",X"46",X"66",X"54",X"3C",X"1E",X"8F",X"C7",X"E3",X"71",X"38",X"9C",
		X"43",X"A1",X"08",X"46",X"B2",X"45",X"B2",X"91",X"E1",X"F0",X"7C",X"9E",X"4F",X"43",X"F9",X"94",
		X"F8",X"7E",X"3F",X"0F",X"87",X"C1",X"F0",X"78",X"62",X"CE",X"B7",X"35",X"CA",X"2D",X"C6",X"59",
		X"C3",X"00",X"42",X"06",X"F5",X"B2",X"CF",X"70",X"FF",X"FF",X"0F",X"40",X"64",X"07",X"2A",X"94",
		X"00",X"E0",X"FC",X"FF",X"1F",X"83",X"84",X"A6",X"7F",X"1F",X"07",X"81",X"C8",X"C0",X"42",X"03",
		X"80",X"E0",X"F0",X"FC",X"7E",X"1F",X"0F",X"83",X"F6",X"7D",X"DB",X"DD",X"2E",X"B7",X"49",X"BB",
		X"FF",X"FF",X"FF",X"01",X"00",X"00",X"C2",X"C3",X"F0",X"FF",X"FF",X"FF",X"0F",X"00",X"00",X"F0",
		X"FF",X"FF",X"FE",X"FC",X"F8",X"F8",X"F9",X"FB",X"FF",X"FF",X"7F",X"3F",X"1F",X"1F",X"9F",X"DF",
		X"FF",X"FF",X"00",X"00",X"00",X"C3",X"C3",X"00",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BE",X"B6",X"79",X"FB",X"57",X"4E",X"AA",X"FD",
		X"BF",X"D4",X"DE",X"FF",X"BE",X"67",X"73",X"FF",X"D9",X"AD",X"BB",X"FF",X"FD",X"75",X"EF",X"EF",
		X"BD",X"FB",X"BB",X"9F",X"77",X"7C",X"FE",X"B2",X"FB",X"BB",X"D7",X"EF",X"F6",X"F5",X"FE",X"FA",
		X"6F",X"7F",X"F7",X"DE",X"AC",X"EE",X"DE",X"DF",X"73",X"7F",X"E9",X"7D",X"3E",X"3E",X"6C",X"F5",
		X"82",X"F2",X"AB",X"FE",X"83",X"57",X"E7",X"DF",X"BD",X"FB",X"F9",X"FD",X"EF",X"2F",X"7F",X"4D",
		X"ED",X"DF",X"FE",X"F7",X"E3",X"F3",X"B5",X"F9",X"FF",X"62",X"EB",X"BF",X"A3",X"3F",X"F5",X"F8",
		X"B9",X"33",X"2E",X"5C",X"86",X"D3",X"9B",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"87",X"C7",X"27",X"2D",X"29",X"29",X"4A",X"6C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"0A",X"E5",X"E4",X"0A",X"04",X"00",X"80",X"40",X"02",X"07",X"07",X"02",X"40",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"0F",X"1F",X"3F",X"3F",X"7F",X"7F",X"00",X"00",X"10",X"1C",X"38",X"1C",X"10",X"00",
		X"7F",X"7F",X"3F",X"3F",X"1F",X"0F",X"03",X"00",X"00",X"00",X"00",X"00",X"20",X"18",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"DF",X"DD",X"FF",X"FB",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"EF",X"DF",X"FE",X"FF",X"FF",
		X"FF",X"FC",X"FD",X"FB",X"FF",X"FF",X"FF",X"BF",X"FF",X"FF",X"EF",X"DE",X"FF",X"FF",X"DF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"7A",X"7B",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"90",
		X"00",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"00",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"00",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"00",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"FF",X"F7",X"E1",X"C1",X"C1",X"E1",X"F7",X"FF",X"FF",X"F7",X"E1",X"C1",X"C1",X"E1",X"F7",X"FF",
		X"00",X"00",X"00",X"60",X"7A",X"7B",X"60",X"00",X"00",X"00",X"00",X"00",X"90",X"90",X"00",X"00",
		X"00",X"00",X"3A",X"7A",X"70",X"70",X"7A",X"7B",X"00",X"00",X"10",X"90",X"80",X"80",X"90",X"90",
		X"FF",X"FF",X"FF",X"FE",X"FC",X"F8",X"F0",X"E0",X"FF",X"FF",X"7F",X"3F",X"1F",X"0F",X"07",X"03",
		X"C0",X"F8",X"F8",X"F9",X"FB",X"FB",X"FB",X"FB",X"01",X"07",X"07",X"F7",X"F7",X"07",X"F7",X"F7",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"F8",X"FB",X"FB",X"F8",X"F8",X"F8",X"F8",X"07",X"07",X"77",X"77",X"07",X"07",X"07",X"07",
		X"F8",X"F8",X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"07",X"07",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"00",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"00",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"00",
		X"00",X"00",X"02",X"18",X"70",X"18",X"02",X"00",X"00",X"00",X"10",X"90",X"00",X"90",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"78",X"78",X"79",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",
		X"00",X"00",X"38",X"78",X"70",X"70",X"79",X"38",X"00",X"00",X"10",X"90",X"80",X"80",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"00",X"00",X"78",X"79",X"00",X"00",X"78",X"79",X"00",X"00",X"90",X"90",X"00",X"00",X"90",X"90",
		X"00",X"00",X"38",X"78",X"70",X"70",X"78",X"39",X"00",X"00",X"10",X"10",X"00",X"00",X"90",X"90",
		X"00",X"00",X"60",X"60",X"78",X"79",X"60",X"60",X"00",X"00",X"00",X"00",X"90",X"90",X"00",X"00",
		X"00",X"00",X"38",X"78",X"70",X"70",X"78",X"39",X"00",X"00",X"90",X"90",X"80",X"80",X"90",X"90",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"00",X"00",X"38",X"78",X"71",X"70",X"78",X"39",X"00",X"00",X"90",X"90",X"80",X"00",X"90",X"90",
		X"00",X"00",X"78",X"78",X"00",X"08",X"78",X"79",X"00",X"00",X"90",X"90",X"90",X"80",X"90",X"90",
		X"00",X"00",X"38",X"79",X"70",X"70",X"78",X"39",X"00",X"00",X"90",X"90",X"00",X"00",X"90",X"90",
		X"FA",X"FA",X"FA",X"FA",X"FA",X"FB",X"FB",X"FB",X"22",X"14",X"48",X"80",X"40",X"32",X"00",X"00",
		X"FB",X"FB",X"FB",X"FA",X"FA",X"FA",X"FA",X"FA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"DD",X"C9",X"81",X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"03",X"81",X"C9",X"DD",X"FF",X"FF",X"FF",X"FF",X"F9",X"F8",X"BC",X"F0",X"FC",X"F9",X"F2",X"F8",
		X"00",X"7F",X"7F",X"7F",X"7E",X"79",X"77",X"77",X"00",X"FF",X"FF",X"80",X"7F",X"FF",X"FF",X"FE",
		X"6F",X"5F",X"5F",X"5F",X"3E",X"3F",X"3F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",
		X"00",X"FF",X"FF",X"03",X"FC",X"7F",X"7F",X"FF",X"00",X"FE",X"FE",X"FE",X"FE",X"1E",X"E6",X"F8",
		X"7F",X"7F",X"3F",X"3F",X"7F",X"7F",X"BF",X"FF",X"FE",X"FE",X"FE",X"FE",X"BE",X"DE",X"9E",X"96",
		X"3F",X"3F",X"3F",X"3E",X"5E",X"5F",X"5D",X"69",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"6F",X"77",X"79",X"7E",X"7F",X"7F",X"7F",X"00",X"FF",X"FF",X"FF",X"3F",X"C0",X"FF",X"FF",X"00",
		X"FF",X"BF",X"7F",X"7F",X"27",X"27",X"79",X"79",X"96",X"9E",X"DE",X"BE",X"FE",X"FE",X"FE",X"FC",
		X"FF",X"FF",X"FF",X"F8",X"07",X"FF",X"FF",X"00",X"F2",X"CE",X"3E",X"FE",X"FE",X"FE",X"FE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"07",X"07",X"00",X"00",X"07",X"07",X"07",X"F0",X"F8",X"FC",X"1C",X"1C",X"FC",X"F8",X"F0",
		X"00",X"00",X"01",X"01",X"01",X"1F",X"1F",X"1F",X"00",X"F8",X"FC",X"FC",X"8C",X"FC",X"FC",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"38",
		X"07",X"07",X"06",X"06",X"07",X"03",X"01",X"00",X"9C",X"CC",X"EC",X"7C",X"3C",X"F8",X"F0",X"00",
		X"0C",X"1C",X"1C",X"19",X"19",X"1F",X"1F",X"0F",X"78",X"FC",X"FC",X"CC",X"CC",X"9C",X"9C",X"18",
		X"FF",X"FF",X"F0",X"80",X"23",X"3F",X"9F",X"8F",X"FF",X"FF",X"7F",X"1F",X"0F",X"CF",X"E7",X"F7",
		X"C7",X"00",X"00",X"00",X"01",X"03",X"E7",X"FF",X"F7",X"57",X"13",X"03",X"83",X"83",X"C3",X"E3",
		X"EF",X"EF",X"E7",X"A2",X"00",X"00",X"00",X"30",X"F3",X"E3",X"E3",X"43",X"03",X"03",X"07",X"07",
		X"1C",X"80",X"C0",X"00",X"80",X"FF",X"FF",X"FF",X"07",X"0F",X"0F",X"1F",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"BB",X"FF",X"FF",X"F6",X"DF",X"FA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"FD",X"F9",X"FD",X"BD",X"E9",X"FD",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"7F",X"7E",X"3C",X"3C",X"18",X"10",X"00",
		X"FE",X"DE",X"7E",X"6E",X"3E",X"3C",X"10",X"00",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",
		X"1F",X"1F",X"FE",X"FF",X"7D",X"83",X"FF",X"FE",X"BC",X"DF",X"EF",X"73",X"3C",X"1F",X"07",X"00",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"34",X"84",X"84",X"FC",X"00",X"00",X"00",X"00",X"0F",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"F8",X"F0",X"F0",X"E0",X"C0",X"C0",X"80",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"87",X"C7",X"E7",X"F3",X"F3",X"79",X"FD",X"BC",X"EF",X"F7",X"3B",X"1D",X"0E",X"07",X"03",X"01",
		X"7F",X"5E",X"7C",X"7E",X"2E",X"3F",X"3F",X"17",X"00",X"80",X"80",X"C0",X"C0",X"E0",X"F0",X"78",
		X"17",X"1F",X"1F",X"0B",X"0F",X"0D",X"06",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F4",X"F4",X"F4",X"F4",X"F4",X"F4",X"74",X"34",X"FF",X"FF",X"FF",X"FF",X"FF",X"03",X"00",X"F8",
		X"FF",X"FF",X"FF",X"3F",X"00",X"80",X"FE",X"03",X"FF",X"FF",X"07",X"00",X"E0",X"3F",X"00",X"00",
		X"FF",X"03",X"00",X"F8",X"FF",X"F8",X"F8",X"FC",X"00",X"80",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"6C",X"2D",X"A1",X"A1",X"3F",X"1F",X"0F",X"0F",X"FF",X"7F",X"C3",X"FF",X"F0",X"FC",X"7E",X"9F",
		X"1F",X"F0",X"3F",X"00",X"0F",X"3F",X"3C",X"7B",X"FC",X"0F",X"00",X"E0",X"E0",X"60",X"E0",X"E0",
		X"03",X"00",X"00",X"07",X"0F",X"1E",X"1D",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"FC",X"84",X"84",X"34",X"34",X"74",X"F4",X"00",X"00",X"FF",X"7F",X"01",X"00",X"FC",X"FF",
		X"C0",X"00",X"1F",X"00",X"C0",X"FF",X"FF",X"FF",X"9F",X"1F",X"1E",X"FE",X"FF",X"FF",X"FF",X"FF",
		X"01",X"00",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"C0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",
		X"6F",X"6F",X"EF",X"EF",X"EF",X"EF",X"EF",X"6C",X"F6",X"03",X"03",X"01",X"01",X"00",X"C0",X"FE",
		X"8F",X"80",X"C0",X"C0",X"C0",X"F0",X"FF",X"FF",X"1B",X"0B",X"0D",X"0D",X"FD",X"FE",X"FE",X"06",
		X"00",X"00",X"00",X"7F",X"7F",X"7F",X"71",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F4",X"F4",X"F4",X"E4",X"E4",X"C4",X"8C",X"18",X"01",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",
		X"80",X"00",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",X"FA",X"78",X"78",X"39",X"3B",X"BF",X"9F",
		X"71",X"38",X"2C",X"26",X"23",X"21",X"C1",X"7F",X"60",X"C0",X"C0",X"E0",X"E0",X"F0",X"1F",X"00",
		X"EE",X"EC",X"EC",X"ED",X"ED",X"ED",X"EC",X"EC",X"23",X"03",X"01",X"01",X"C1",X"E0",X"E0",X"74",
		X"0E",X"FC",X"00",X"FC",X"FF",X"FF",X"07",X"FC",X"FE",X"C7",X"FF",X"FF",X"7F",X"C1",X"FA",X"1B",
		X"F9",X"FF",X"FF",X"CF",X"F0",X"1F",X"00",X"00",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"FA",X"28",X"80",X"02",X"03",X"D1",X"20",
		X"7C",X"C8",X"E4",X"F0",X"C4",X"80",X"15",X"CA",X"50",X"A8",X"10",X"28",X"5C",X"28",X"14",X"0A",
		X"5F",X"36",X"1F",X"0F",X"0D",X"86",X"07",X"A3",X"66",X"F7",X"DF",X"BE",X"CC",X"FC",X"67",X"FE",
		X"C1",X"49",X"80",X"8A",X"29",X"21",X"61",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"14",X"14",X"34",X"2C",X"69",X"70",X"C4",X"88",X"21",X"19",X"59",X"13",X"02",X"81",X"A1",X"03",
		X"08",X"38",X"F0",X"E0",X"C7",X"8E",X"FD",X"F7",X"02",X"8E",X"0F",X"99",X"3A",X"FF",X"FE",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"F8",X"FF",X"FF",X"FF",X"E0",X"80",X"07",X"1F",X"7F",
		X"F0",X"C1",X"03",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"02",X"0E",X"03",X"00",X"0F",X"0F",X"0B",X"0B",
		X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"0B",X"0B",X"0F",X"0F",X"00",X"00",X"00",X"00",
		X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"01",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"0F",X"07",X"C3",X"E3",
		X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"F1",X"F1",X"F8",X"F8",X"FC",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"01",X"80",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"01",X"80",X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"01",X"80",X"F8",X"FF",X"FF",X"FF",
		X"F3",X"F3",X"F3",X"F3",X"03",X"03",X"FF",X"FF",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FC",X"F9",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F1",X"F1",X"E1",X"E1",X"E1",X"E1",X"E1",X"F1",
		X"F1",X"F9",X"FC",X"FE",X"00",X"98",X"00",X"08",X"FF",X"FF",X"FF",X"00",X"00",X"96",X"08",X"40",
		X"00",X"00",X"6A",X"00",X"00",X"B1",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"0F",
		X"0F",X"0F",X"1F",X"1F",X"1F",X"1F",X"1F",X"0F",X"83",X"2B",X"07",X"17",X"97",X"E7",X"FF",X"FD",
		X"3C",X"3C",X"3C",X"3C",X"3C",X"3F",X"3F",X"3F",X"10",X"00",X"20",X"02",X"00",X"44",X"B6",X"00",
		X"E0",X"18",X"C0",X"82",X"00",X"02",X"11",X"04",X"C8",X"C0",X"D0",X"C2",X"D0",X"D0",X"C4",X"D0",
		X"0F",X"0F",X"07",X"03",X"00",X"00",X"00",X"00",X"FE",X"FC",X"F8",X"F0",X"E0",X"C0",X"80",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"A4",X"C1",X"87",X"0D",X"57",X"9F",X"2F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"1E",X"3E",X"20",X"3E",X"00",X"1C",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"22",X"3E",X"1C",X"00",X"3E",X"00",X"20",X"3E",X"03",X"0F",X"06",X"00",X"00",X"00",X"00",X"00",
		X"50",X"50",X"58",X"18",X"00",X"07",X"8F",X"8F",X"7E",X"6E",X"46",X"46",X"46",X"06",X"82",X"C2",
		X"C7",X"00",X"00",X"00",X"01",X"03",X"E7",X"FF",X"E2",X"42",X"02",X"02",X"82",X"82",X"C2",X"E2",
		X"20",X"00",X"3E",X"02",X"3E",X"3E",X"00",X"3E",X"01",X"03",X"13",X"3B",X"31",X"38",X"18",X"0C",
		X"24",X"3C",X"0E",X"00",X"22",X"3E",X"1C",X"00",X"0F",X"07",X"01",X"00",X"00",X"00",X"00",X"00",
		X"EF",X"EF",X"E7",X"A2",X"00",X"00",X"00",X"30",X"F2",X"E2",X"E2",X"42",X"02",X"02",X"06",X"06",
		X"1C",X"80",X"C0",X"00",X"00",X"74",X"34",X"24",X"06",X"0E",X"0E",X"1E",X"3E",X"3E",X"3E",X"3E",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"FF",X"E3",X"C3",X"83",X"8F",X"9E",X"8C",X"80",X"FF",X"C3",X"81",X"00",X"18",X"3C",X"78",X"60",
		X"C0",X"E1",X"FF",X"C0",X"80",X"80",X"9F",X"9F",X"E1",X"E3",X"FF",X"00",X"00",X"00",X"3F",X"3F",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"8F",X"80",X"C0",X"F0",X"FF",X"E3",X"C3",X"83",X"3F",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"8F",X"9F",X"9F",X"8F",X"80",X"C0",X"E0",X"FF",X"3C",X"3C",X"3C",X"F8",X"00",X"01",X"03",X"FF",
		X"00",X"38",X"3E",X"3F",X"31",X"3F",X"36",X"32",X"00",X"9F",X"FF",X"FF",X"1F",X"FF",X"DF",X"5B",
		X"3F",X"3F",X"36",X"37",X"30",X"3F",X"3F",X"38",X"DD",X"FC",X"1E",X"DF",X"5F",X"FF",X"FF",X"1F",
		X"00",X"FF",X"FE",X"DF",X"DF",X"CF",X"CF",X"E7",X"00",X"FC",X"FC",X"FC",X"7C",X"7C",X"7C",X"3C",
		X"E7",X"E2",X"30",X"10",X"88",X"C0",X"E0",X"80",X"3C",X"3C",X"1C",X"1C",X"0C",X"0C",X"0C",X"0C",
		X"3F",X"3F",X"30",X"3F",X"38",X"3F",X"3F",X"30",X"DF",X"FF",X"1C",X"FB",X"1F",X"DF",X"FF",X"9F",
		X"3F",X"38",X"3F",X"3F",X"30",X"3F",X"3F",X"00",X"FF",X"3F",X"9F",X"DF",X"5F",X"FF",X"FF",X"00",
		X"00",X"30",X"F8",X"F0",X"F1",X"E3",X"E6",X"CE",X"0C",X"8C",X"1C",X"1C",X"3C",X"3C",X"7C",X"7C",
		X"DE",X"BE",X"FE",X"7E",X"FF",X"FB",X"FF",X"00",X"7C",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"00",X"C0",X"20",X"00",X"F0",X"F0",X"F0",X"F0",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"FF",X"FF",X"FF",X"0F",X"03",X"C1",X"F0",X"F8",X"1F",X"0F",X"87",X"C3",X"E0",X"F0",X"FF",X"7F",
		X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"07",X"80",X"E0",X"FF",X"FF",X"FF",X"FF",
		X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"FE",
		X"00",X"1E",X"3F",X"20",X"3F",X"11",X"1E",X"22",X"F8",X"E1",X"DF",X"FD",X"FD",X"FE",X"FE",X"FF",
		X"22",X"7E",X"7C",X"60",X"3E",X"00",X"20",X"3E",X"FC",X"7E",X"3F",X"0F",X"03",X"09",X"48",X"41",
		X"FF",X"FF",X"EF",X"E1",X"B8",X"BE",X"4F",X"F2",X"C2",X"82",X"82",X"02",X"42",X"C2",X"82",X"82",
		X"EC",X"FC",X"F9",X"8E",X"C0",X"79",X"30",X"80",X"02",X"06",X"06",X"0E",X"0E",X"1C",X"36",X"A4",
		X"20",X"00",X"3E",X"02",X"3E",X"3E",X"00",X"1E",X"40",X"C2",X"C2",X"C2",X"C2",X"C6",X"44",X"01",
		X"24",X"3E",X"0E",X"04",X"22",X"3E",X"1C",X"0C",X"02",X"0F",X"0E",X"1E",X"1F",X"37",X"3E",X"3B",
		X"B8",X"9A",X"89",X"2A",X"39",X"0A",X"60",X"98",X"00",X"00",X"40",X"D2",X"D0",X"C0",X"EA",X"C4",
		X"04",X"62",X"F2",X"BA",X"78",X"CC",X"A4",X"F2",X"4C",X"70",X"60",X"2A",X"30",X"3A",X"3C",X"14",
		X"1C",X"7C",X"7C",X"7C",X"5C",X"0C",X"04",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"74",X"74",X"7C",X"7C",X"7C",X"7C",X"7C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"12",X"10",X"08",X"08",X"02",X"00",X"11",X"11",X"60",X"C0",X"60",X"40",X"20",X"A0",X"20",X"60",
		X"00",X"00",X"02",X"10",X"10",X"10",X"08",X"11",X"C0",X"60",X"C0",X"60",X"60",X"A0",X"60",X"40",
		X"7C",X"7C",X"7C",X"7C",X"6C",X"4C",X"0C",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"6C",X"7C",X"7C",X"5C",X"1C",X"0C",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"08",X"08",X"00",X"10",X"00",X"00",X"10",X"20",X"20",X"90",X"50",X"30",X"A0",X"60",X"40",
		X"09",X"08",X"08",X"20",X"20",X"20",X"10",X"11",X"60",X"20",X"50",X"30",X"90",X"30",X"60",X"20",
		X"1D",X"05",X"00",X"1D",X"05",X"00",X"19",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"13",X"01",X"00",X"11",X"11",X"1D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"04",X"10",X"34",X"34",X"34",X"3A",X"00",X"00",X"00",X"60",X"F0",X"D0",X"D0",X"00",
		X"2A",X"02",X"03",X"03",X"0B",X"1A",X"18",X"39",X"40",X"40",X"00",X"40",X"60",X"68",X"48",X"18",
		X"15",X"15",X"15",X"01",X"00",X"1F",X"00",X"1B",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",
		X"01",X"00",X"11",X"11",X"1D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3A",X"36",X"36",X"AE",X"8E",X"CC",X"D9",X"FB",X"F8",X"E8",X"E8",X"18",X"08",X"C0",X"80",X"E0",
		X"6B",X"3A",X"3A",X"02",X"00",X"00",X"00",X"00",X"90",X"D0",X"F0",X"60",X"00",X"00",X"00",X"00",
		X"7F",X"40",X"40",X"40",X"40",X"47",X"40",X"40",X"FF",X"00",X"00",X"20",X"20",X"A0",X"20",X"20",
		X"40",X"41",X"40",X"40",X"40",X"44",X"43",X"40",X"00",X"E0",X"20",X"20",X"00",X"40",X"60",X"00",
		X"FF",X"00",X"68",X"68",X"68",X"68",X"68",X"40",X"FE",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"00",X"00",X"60",X"68",X"60",X"40",X"00",X"00",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"43",X"40",X"44",X"47",X"40",X"40",X"40",X"44",X"C0",X"20",X"20",X"A0",X"20",X"00",X"00",X"E0",
		X"44",X"44",X"47",X"40",X"40",X"40",X"40",X"7F",X"20",X"20",X"A0",X"20",X"00",X"00",X"00",X"FF",
		X"20",X"10",X"40",X"68",X"28",X"00",X"00",X"00",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"68",X"68",X"68",X"68",X"68",X"68",X"00",X"FF",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"FE",
		X"00",X"C0",X"0B",X"84",X"11",X"C0",X"30",X"49",X"02",X"85",X"2A",X"05",X"0A",X"84",X"18",X"67",
		X"00",X"2E",X"C0",X"2A",X"21",X"4C",X"B3",X"08",X"90",X"6F",X"90",X"02",X"A4",X"01",X"08",X"80",
		X"00",X"02",X"20",X"00",X"50",X"00",X"08",X"10",X"10",X"02",X"54",X"01",X"4A",X"02",X"A0",X"30",
		X"00",X"00",X"4A",X"20",X"35",X"40",X"66",X"E0",X"10",X"80",X"0A",X"08",X"03",X"54",X"20",X"10",
		X"E0",X"74",X"79",X"B0",X"02",X"4C",X"10",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"BE",X"3F",X"7F",X"1F",X"BF",X"1F",X"4F",X"0D",X"A4",X"42",X"A0",X"D2",X"A1",X"D2",X"E8",X"D0",
		X"1F",X"86",X"0D",X"03",X"53",X"84",X"10",X"02",X"F8",X"90",X"D8",X"F0",X"E2",X"C8",X"12",X"80",
		X"00",X"20",X"10",X"90",X"00",X"60",X"1A",X"75",X"7A",X"7D",X"FA",X"BD",X"FE",X"7D",X"7E",X"7F",
		X"83",X"0F",X"1D",X"7F",X"7F",X"EF",X"FF",X"F7",X"C8",X"86",X"3E",X"FC",X"F0",X"C4",X"BE",X"FF",
		X"FE",X"F9",X"F8",X"FE",X"FC",X"F8",X"A0",X"E3",X"1F",X"87",X"03",X"41",X"21",X"10",X"08",X"00",
		X"E3",X"E3",X"E1",X"C0",X"D8",X"FE",X"FB",X"FF",X"00",X"C0",X"89",X"09",X"1F",X"3F",X"FF",X"BF",
		X"FF",X"FF",X"EF",X"7E",X"7F",X"3E",X"1F",X"87",X"FF",X"DA",X"E0",X"F8",X"FC",X"3C",X"8E",X"C0",
		X"0B",X"00",X"80",X"02",X"90",X"40",X"80",X"49",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"F8",X"F8",X"FE",X"9C",X"8C",X"84",X"80",X"D0",X"11",X"84",
		X"FC",X"FC",X"FC",X"FE",X"FE",X"F8",X"C0",X"C2",X"8F",X"6D",X"28",X"08",X"10",X"10",X"E0",X"60",
		X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"F8",X"FA",X"F8",X"D0",X"82",X"04",X"20",X"00",X"00",X"48",
		X"F8",X"F0",X"F8",X"F0",X"E0",X"E0",X"E1",X"E8",X"00",X"40",X"00",X"00",X"41",X"03",X"07",X"07",
		X"FF",X"FF",X"FD",X"FD",X"F7",X"FE",X"EE",X"FC",X"EF",X"BC",X"E0",X"80",X"00",X"00",X"00",X"05",
		X"FC",X"C8",X"F8",X"F8",X"F0",X"D1",X"F1",X"F3",X"0D",X"1B",X"39",X"3B",X"66",X"40",X"10",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"F8",X"C0",X"02",X"17",
		X"FC",X"FC",X"F8",X"F8",X"F8",X"F0",X"F0",X"F0",X"1F",X"0F",X"06",X"00",X"00",X"00",X"00",X"00",
		X"77",X"D5",X"F3",X"F7",X"F7",X"D1",X"D1",X"F0",X"00",X"21",X"08",X"88",X"84",X"83",X"48",X"E0",
		X"E8",X"E8",X"F8",X"F4",X"FC",X"FA",X"FB",X"FE",X"F0",X"E8",X"DB",X"5B",X"3A",X"09",X"01",X"80",
		X"F0",X"F0",X"F0",X"FA",X"FB",X"FB",X"F9",X"FC",X"01",X"03",X"13",X"7B",X"E9",X"E0",X"C8",X"9C",
		X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"3F",X"13",X"C0",X"F8",X"FF",X"FF",X"FF",
		X"FC",X"F8",X"F0",X"F0",X"70",X"00",X"40",X"50",X"FF",X"7F",X"1F",X"03",X"00",X"00",X"00",X"00",
		X"18",X"1C",X"5F",X"9F",X"5F",X"1F",X"5F",X"5F",X"00",X"00",X"00",X"E0",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FE",X"FE",X"FE",X"FD",X"3D",X"1A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"7F",X"7F",X"7F",X"7F",X"3F",X"9F",X"C0",
		X"00",X"00",X"00",X"10",X"FE",X"DC",X"EE",X"FE",X"00",X"00",X"00",X"10",X"C2",X"84",X"C2",X"EE",
		X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"03",X"03",X"01",X"00",X"00",X"C0",X"C0",X"E0",X"E0");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
