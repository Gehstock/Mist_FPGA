library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity gfx2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of gfx2 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"08",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"02",X"20",X"20",X"20",
		X"10",X"10",X"10",X"30",X"30",X"21",X"61",X"43",X"00",X"00",X"00",X"80",X"80",X"80",X"C0",X"48",
		X"A0",X"A8",X"E0",X"E8",X"86",X"80",X"00",X"00",X"A0",X"B2",X"F0",X"E2",X"2C",X"20",X"00",X"00",
		X"C3",X"D2",X"F0",X"74",X"76",X"70",X"30",X"03",X"68",X"78",X"F0",X"C4",X"CC",X"C0",X"80",X"08",
		X"00",X"00",X"00",X"00",X"08",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"02",X"20",X"20",X"20",
		X"10",X"10",X"10",X"30",X"30",X"21",X"61",X"43",X"00",X"00",X"00",X"80",X"80",X"80",X"C0",X"48",
		X"A0",X"A8",X"E0",X"E8",X"80",X"80",X"00",X"00",X"A0",X"B2",X"F0",X"E2",X"20",X"20",X"00",X"00",
		X"C3",X"D2",X"F0",X"74",X"76",X"70",X"30",X"03",X"68",X"78",X"F0",X"C4",X"CC",X"C0",X"80",X"08",
		X"00",X"00",X"80",X"40",X"60",X"E1",X"C6",X"20",X"00",X"00",X"20",X"10",X"11",X"11",X"00",X"00",
		X"00",X"00",X"00",X"CC",X"F1",X"B4",X"C3",X"CB",X"00",X"08",X"40",X"20",X"11",X"F6",X"78",X"3C",
		X"00",X"88",X"80",X"84",X"08",X"00",X"00",X"00",X"04",X"20",X"10",X"00",X"20",X"10",X"00",X"00",
		X"43",X"65",X"74",X"F8",X"60",X"E2",X"D2",X"04",X"F1",X"F1",X"F0",X"FC",X"74",X"01",X"00",X"00",
		X"00",X"00",X"80",X"40",X"60",X"E0",X"C4",X"20",X"00",X"00",X"20",X"10",X"11",X"11",X"00",X"00",
		X"00",X"00",X"00",X"CC",X"F1",X"B4",X"C3",X"CB",X"00",X"08",X"40",X"20",X"11",X"F6",X"78",X"3C",
		X"00",X"88",X"80",X"84",X"08",X"00",X"00",X"00",X"04",X"20",X"10",X"00",X"20",X"10",X"00",X"00",
		X"43",X"65",X"74",X"F8",X"60",X"E2",X"D0",X"00",X"F1",X"F1",X"F0",X"FC",X"74",X"01",X"00",X"00",
		X"08",X"08",X"C0",X"00",X"00",X"C8",X"E9",X"E1",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"F0",
		X"00",X"00",X"78",X"00",X"00",X"30",X"E1",X"87",X"F0",X"30",X"F5",X"60",X"E0",X"F1",X"3C",X"78",
		X"E9",X"C8",X"00",X"00",X"C0",X"08",X"08",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E1",X"30",X"00",X"00",X"78",X"00",X"00",X"00",X"3C",X"F1",X"E0",X"60",X"F5",X"30",X"F0",X"00",
		X"00",X"00",X"C0",X"00",X"00",X"C8",X"E9",X"E1",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"F0",
		X"00",X"00",X"78",X"00",X"00",X"30",X"E1",X"87",X"F0",X"30",X"F5",X"60",X"E0",X"F1",X"3C",X"78",
		X"E9",X"C8",X"00",X"00",X"C0",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E1",X"30",X"00",X"00",X"78",X"00",X"00",X"00",X"3C",X"F1",X"E0",X"60",X"F5",X"30",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"06",X"03",X"03",X"00",X"00",X"00",X"00",X"01",X"03",X"06",X"06",
		X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"01",X"03",X"06",X"06",
		X"0F",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"06",X"03",X"01",X"00",X"00",X"00",X"00",X"00",
		X"03",X"03",X"0F",X"00",X"00",X"00",X"00",X"00",X"07",X"06",X"06",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"06",X"07",X"07",X"07",
		X"00",X"00",X"00",X"00",X"03",X"07",X"0F",X"0F",X"00",X"00",X"00",X"00",X"07",X"06",X"06",X"07",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"06",X"00",X"00",X"00",X"00",X"00",
		X"0B",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"07",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"03",X"03",X"52",X"52",X"03",X"07",X"00",X"00",X"88",X"88",X"C8",X"C8",X"88",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"17",X"96",X"96",X"96",X"96",X"77",X"33",X"11",X"CC",X"EC",X"EC",X"EC",X"EC",X"CC",X"88",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"26",X"17",X"17",X"35",X"52",X"43",X"03",X"00",X"00",X"00",X"00",X"80",X"C8",X"88",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"07",X"43",X"43",X"43",X"21",X"00",X"00",X"EC",X"F6",X"F6",X"F6",X"F7",X"EE",X"EE",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"01",X"01",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"4C",X"3E",X"7B",X"B5",X"87",X"03",X"00",X"00",X"00",X"00",X"80",X"00",X"CC",X"EC",
		X"00",X"80",X"80",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"03",X"43",X"21",X"21",X"10",X"00",X"00",X"F6",X"F7",X"7B",X"7B",X"7F",X"FF",X"33",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"13",X"03",X"01",X"01",X"10",X"00",
		X"00",X"00",X"00",X"EC",X"7E",X"7B",X"3D",X"87",X"00",X"00",X"00",X"00",X"00",X"00",X"EC",X"FE",
		X"80",X"C8",X"CC",X"CC",X"88",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"03",X"21",X"10",X"00",X"00",X"00",X"00",X"F7",X"7B",X"3D",X"1E",X"B7",X"73",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C8",X"00",X"00",X"08",X"37",X"03",X"03",X"01",X"10",
		X"00",X"00",X"00",X"00",X"E8",X"E6",X"7B",X"1F",X"00",X"00",X"00",X"00",X"00",X"A8",X"FE",X"FF",
		X"CC",X"CC",X"EE",X"EE",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"83",X"03",X"10",X"00",X"00",X"00",X"00",X"00",X"F3",X"3C",X"0F",X"87",X"71",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"C8",X"CC",X"00",X"00",X"00",X"00",X"00",X"1F",X"07",X"03",
		X"00",X"00",X"00",X"00",X"00",X"E8",X"F7",X"5B",X"00",X"00",X"00",X"00",X"00",X"FC",X"FF",X"FF",
		X"E6",X"7F",X"6E",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"87",X"41",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"0F",X"87",X"70",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"CC",X"EE",X"F7",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"D1",X"FF",X"C3",X"00",X"00",X"00",X"00",X"70",X"FF",X"FF",X"F8",
		X"6E",X"4C",X"80",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"C1",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"70",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"03",X"03",X"07",X"00",X"00",X"00",X"00",X"03",X"06",X"06",X"06",
		X"00",X"00",X"00",X"00",X"0E",X"03",X"03",X"03",X"00",X"00",X"00",X"00",X"06",X"06",X"06",X"07",
		X"0E",X"0C",X"08",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"03",X"00",X"00",X"00",X"00",X"00",
		X"03",X"03",X"0E",X"00",X"00",X"00",X"00",X"00",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"01",X"01",X"01",X"03",X"13",X"17",X"00",X"80",X"80",X"80",X"80",X"48",X"C8",X"AC",
		X"00",X"C0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"30",X"00",X"00",X"00",X"00",
		X"1F",X"0F",X"0F",X"0F",X"B4",X"24",X"24",X"00",X"9E",X"0F",X"0F",X"3C",X"B4",X"24",X"24",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"24",X"42",X"12",X"03",X"13",X"53",X"00",X"00",X"00",X"00",X"00",X"48",X"AC",X"9E",
		X"F0",X"68",X"C0",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"01",X"03",X"10",X"00",X"00",X"00",
		X"07",X"0F",X"0F",X"0F",X"87",X"21",X"01",X"00",X"8F",X"0F",X"1E",X"1E",X"E1",X"81",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"68",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"80",X"48",X"24",X"24",X"03",X"17",X"53",X"00",X"00",X"00",X"00",X"80",X"1C",X"9E",X"8F",
		X"68",X"C0",X"C0",X"48",X"48",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"01",X"00",X"00",
		X"07",X"07",X"07",X"0F",X"2D",X"50",X"00",X"00",X"8F",X"0F",X"0F",X"2D",X"48",X"68",X"24",X"00",
		X"00",X"00",X"00",X"20",X"60",X"E0",X"68",X"C0",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"C0",X"78",X"16",X"17",X"17",X"00",X"00",X"00",X"00",X"00",X"F0",X"8F",X"CF",
		X"C0",X"68",X"24",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"03",X"03",X"03",X"43",X"16",X"A4",X"00",X"8F",X"0F",X"1E",X"3C",X"3C",X"52",X"00",X"00",
		X"00",X"00",X"00",X"40",X"C0",X"C0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"24",X"12",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"B0",X"0F",X"B7",X"00",X"00",X"00",X"00",X"00",X"F0",X"1E",X"0F",
		X"C0",X"68",X"24",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"07",X"03",X"43",X"03",X"03",X"03",X"02",X"8F",X"0F",X"1E",X"1E",X"1E",X"69",X"80",X"00",
		X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"E0",X"00",X"00",X"00",X"00",X"00",X"34",X"21",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"0F",X"B7",X"00",X"00",X"10",X"30",X"52",X"87",X"0F",X"1E",
		X"0E",X"80",X"80",X"C0",X"48",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"37",X"43",X"03",X"21",X"01",X"01",X"00",X"00",X"8F",X"0F",X"0F",X"0F",X"0F",X"2C",X"48",X"08",
		X"00",X"00",X"00",X"00",X"80",X"E0",X"0E",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",
		X"00",X"00",X"00",X"00",X"00",X"10",X"61",X"B7",X"00",X"20",X"70",X"70",X"96",X"1E",X"0F",X"8F",
		X"80",X"E0",X"0E",X"80",X"00",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"07",X"01",X"00",X"00",X"00",X"00",X"00",X"8F",X"0F",X"0F",X"0F",X"16",X"16",X"02",X"00",
		X"00",X"00",X"00",X"00",X"0E",X"03",X"03",X"07",X"00",X"00",X"00",X"00",X"07",X"06",X"06",X"07",
		X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"07",X"06",X"06",X"06",
		X"0C",X"0E",X"07",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"07",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"07",X"06",X"06",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",
		X"00",X"00",X"03",X"17",X"3F",X"3F",X"1F",X"78",X"00",X"00",X"80",X"C0",X"E8",X"BC",X"1E",X"1E",
		X"80",X"C0",X"48",X"48",X"04",X"04",X"00",X"00",X"03",X"16",X"34",X"24",X"04",X"04",X"00",X"00",
		X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
		X"00",X"00",X"16",X"36",X"3F",X"3F",X"1F",X"78",X"00",X"00",X"00",X"C0",X"F0",X"1E",X"1E",X"0F",
		X"2C",X"3C",X"12",X"01",X"00",X"00",X"00",X"00",X"21",X"03",X"03",X"12",X"12",X"02",X"00",X"00",
		X"68",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"2C",X"00",X"00",X"00",X"00",X"01",X"01",X"21",X"21",
		X"00",X"00",X"70",X"3C",X"7F",X"7F",X"6F",X"3C",X"00",X"00",X"00",X"C0",X"68",X"3C",X"0F",X"43",
		X"87",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"21",X"01",X"01",X"01",X"01",X"01",X"10",X"00",
		X"68",X"68",X"48",X"C0",X"C0",X"80",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"C0",X"4A",X"01",X"00",X"00",X"00",X"10",X"13",X"03",X"13",X"03",X"03",
		X"00",X"00",X"F0",X"D6",X"CF",X"CF",X"68",X"48",X"00",X"00",X"C0",X"F0",X"1E",X"0F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"21",X"21",X"30",X"01",X"00",X"00",X"00",
		X"48",X"48",X"48",X"48",X"48",X"48",X"04",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"C0",X"0F",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"03",X"03",
		X"00",X"00",X"30",X"E1",X"C3",X"EF",X"FE",X"DE",X"00",X"00",X"E0",X"78",X"0F",X"3C",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"3C",X"1E",X"16",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"80",X"08",X"08",X"84",
		X"00",X"00",X"0C",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"13",X"03",
		X"00",X"00",X"00",X"30",X"C3",X"87",X"CF",X"FE",X"00",X"00",X"F0",X"87",X"1E",X"68",X"08",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1E",X"1E",X"1E",X"1E",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"2C",X"86",
		X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"30",
		X"00",X"00",X"00",X"10",X"70",X"C3",X"87",X"CF",X"00",X"00",X"70",X"C3",X"0E",X"0C",X"08",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"13",X"03",X"01",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"DE",X"1E",X"0F",X"07",X"01",X"00",X"00",X"00",X"00",X"80",X"C0",X"68",X"3C",X"07",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
		X"00",X"01",X"03",X"07",X"0D",X"0D",X"0F",X"0F",X"00",X"00",X"80",X"C0",X"60",X"60",X"3C",X"3C",
		X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"03",X"03",X"12",X"02",X"02",X"00",X"00",X"00",
		X"0F",X"CB",X"B8",X"10",X"10",X"10",X"00",X"00",X"78",X"F2",X"B2",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"21",
		X"00",X"04",X"34",X"16",X"0A",X"0A",X"0F",X"0F",X"00",X"00",X"00",X"C0",X"C0",X"F0",X"3C",X"78",
		X"80",X"C0",X"40",X"00",X"00",X"00",X"00",X"00",X"21",X"21",X"03",X"01",X"01",X"01",X"00",X"00",
		X"0F",X"0F",X"D8",X"C4",X"00",X"00",X"00",X"00",X"7A",X"D1",X"C0",X"80",X"80",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"00",X"00",X"01",X"10",X"10",X"10",X"01",X"00",
		X"00",X"00",X"00",X"3C",X"1C",X"0A",X"0B",X"0F",X"00",X"00",X"00",X"80",X"E0",X"78",X"3C",X"79",
		X"E0",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"6D",X"2E",X"48",X"04",X"04",X"00",X"79",X"68",X"C0",X"40",X"20",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"20",X"00",X"00",X"00",X"01",X"10",X"01",X"10",X"10",
		X"00",X"00",X"00",X"E0",X"38",X"05",X"0B",X"0F",X"00",X"00",X"00",X"00",X"E0",X"78",X"7A",X"79",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"3E",X"97",X"24",X"02",X"01",X"00",X"68",X"68",X"E0",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"E0",X"00",X"00",X"00",X"00",X"00",X"12",X"01",X"01",X"01",X"01",
		X"00",X"00",X"00",X"E0",X"F0",X"09",X"07",X"0B",X"00",X"00",X"00",X"C0",X"F0",X"7A",X"79",X"68",
		X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"87",X"17",X"43",X"01",X"00",X"00",X"68",X"78",X"C0",X"88",X"80",X"80",X"48",X"00",
		X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"07",X"03",X"03",
		X"00",X"00",X"10",X"70",X"E1",X"03",X"0F",X"03",X"00",X"00",X"F0",X"F0",X"7A",X"3D",X"48",X"68",
		X"80",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"07",X"01",X"00",X"00",X"00",X"78",X"E0",X"88",X"4C",X"48",X"24",X"00",X"00",
		X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"30",
		X"00",X"00",X"00",X"00",X"30",X"F0",X"C3",X"03",X"00",X"00",X"00",X"F0",X"E0",X"E6",X"C0",X"68",
		X"C0",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"03",X"0F",X"0F",X"03",X"00",X"00",X"00",X"3C",X"2C",X"48",X"6E",X"2C",X"0F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"08",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"02",X"30",X"01",X"00",X"01",
		X"00",X"00",X"02",X"02",X"38",X"D3",X"91",X"6E",X"00",X"00",X"00",X"05",X"61",X"C6",X"61",X"23",
		X"00",X"00",X"08",X"80",X"04",X"00",X"00",X"00",X"00",X"00",X"01",X"30",X"00",X"00",X"00",X"00",
		X"26",X"59",X"D2",X"20",X"04",X"00",X"00",X"00",X"46",X"CB",X"69",X"68",X"04",X"00",X"00",X"00",
		X"00",X"20",X"68",X"48",X"80",X"8C",X"08",X"00",X"04",X"61",X"30",X"10",X"10",X"00",X"00",X"71",
		X"00",X"00",X"1A",X"F2",X"D4",X"B9",X"EE",X"CC",X"00",X"00",X"40",X"F8",X"CC",X"77",X"33",X"31",
		X"88",X"08",X"4C",X"88",X"C0",X"60",X"20",X"00",X"00",X"01",X"11",X"00",X"10",X"30",X"42",X"00",
		X"EA",X"EF",X"9D",X"B0",X"7D",X"60",X"00",X"00",X"74",X"33",X"AE",X"7C",X"26",X"42",X"12",X"00",
		X"33",X"46",X"8C",X"CC",X"0C",X"88",X"8C",X"EF",X"88",X"66",X"37",X"13",X"11",X"01",X"32",X"67",
		X"00",X"00",X"19",X"0F",X"37",X"D8",X"80",X"D0",X"44",X"88",X"08",X"8D",X"1F",X"42",X"10",X"39",
		X"88",X"C4",X"EE",X"00",X"88",X"CC",X"66",X"13",X"DE",X"10",X"11",X"23",X"67",X"66",X"CC",X"88",
		X"84",X"09",X"5F",X"A1",X"4F",X"44",X"00",X"00",X"B0",X"03",X"41",X"B7",X"9F",X"8D",X"88",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"06",X"02",X"02",X"00",X"00",X"00",X"00",X"07",X"08",X"00",X"01",
		X"00",X"00",X"00",X"00",X"01",X"0A",X"0A",X"02",X"00",X"00",X"00",X"00",X"08",X"0D",X"05",X"05",
		X"02",X"0A",X"0C",X"00",X"00",X"00",X"00",X"00",X"02",X"04",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"02",X"03",X"09",X"00",X"00",X"00",X"00",X"00",X"05",X"05",X"08",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"06",X"02",X"02",X"00",X"00",X"00",X"00",X"01",X"03",X"05",X"09",
		X"00",X"00",X"00",X"00",X"01",X"02",X"02",X"02",X"00",X"00",X"00",X"00",X"08",X"0D",X"05",X"05",
		X"02",X"0A",X"0C",X"00",X"00",X"00",X"00",X"00",X"0F",X"01",X"01",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"05",X"05",X"08",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"06",X"02",X"02",X"00",X"00",X"00",X"00",X"07",X"08",X"08",X"07",
		X"00",X"00",X"00",X"00",X"01",X"0A",X"0A",X"02",X"00",X"00",X"00",X"00",X"08",X"0D",X"05",X"05",
		X"02",X"0A",X"0C",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"07",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"0B",X"01",X"00",X"00",X"00",X"00",X"00",X"05",X"05",X"08",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"06",X"02",X"02",X"00",X"00",X"00",X"00",X"0F",X"08",X"0F",X"00",
		X"00",X"00",X"00",X"00",X"09",X"02",X"02",X"0A",X"00",X"00",X"00",X"00",X"08",X"0D",X"05",X"05",
		X"02",X"0A",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"07",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"0B",X"01",X"00",X"00",X"00",X"00",X"00",X"05",X"05",X"08",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"06",X"0B",X"09",X"09",X"00",X"00",X"00",X"00",X"09",X"0A",X"0A",X"0A",
		X"00",X"00",X"00",X"00",X"08",X"0D",X"05",X"05",X"00",X"00",X"00",X"00",X"0C",X"06",X"02",X"02",
		X"09",X"0D",X"06",X"00",X"00",X"00",X"00",X"00",X"0A",X"0B",X"09",X"00",X"00",X"00",X"00",X"00",
		X"05",X"05",X"08",X"00",X"00",X"00",X"00",X"00",X"02",X"0A",X"0C",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"06",X"0B",X"09",X"09",X"00",X"00",X"00",X"00",X"0B",X"0A",X"0B",X"08",
		X"00",X"00",X"00",X"00",X"0C",X"01",X"09",X"05",X"00",X"00",X"00",X"00",X"0C",X"06",X"02",X"02",
		X"09",X"0D",X"06",X"00",X"00",X"00",X"00",X"00",X"08",X"0A",X"09",X"00",X"00",X"00",X"00",X"00",
		X"05",X"05",X"08",X"00",X"00",X"00",X"00",X"00",X"02",X"0A",X"0C",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"16",X"29",X"66",X"CC",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"60",X"10",X"00",X"00",X"00",X"00",X"01",X"06",X"08",X"19",
		X"83",X"07",X"0F",X"1E",X"3C",X"1E",X"0F",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"10",
		X"01",X"01",X"02",X"02",X"00",X"03",X"04",X"B7",X"13",X"52",X"94",X"84",X"08",X"00",X"88",X"8A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"1A",X"14",X"00",X"00",
		X"00",X"00",X"08",X"06",X"67",X"FF",X"33",X"11",X"00",X"00",X"00",X"10",X"20",X"48",X"04",X"84",
		X"00",X"00",X"00",X"20",X"48",X"04",X"02",X"02",X"0E",X"87",X"87",X"C3",X"69",X"C3",X"87",X"0F",
		X"30",X"01",X"0A",X"08",X"08",X"08",X"08",X"02",X"08",X"00",X"06",X"01",X"66",X"32",X"33",X"13",
		X"03",X"00",X"03",X"0F",X"0D",X"01",X"01",X"01",X"00",X"00",X"01",X"02",X"02",X"01",X"00",X"00",
		X"2A",X"6E",X"64",X"C8",X"8C",X"66",X"3B",X"06",X"03",X"03",X"03",X"03",X"03",X"03",X"00",X"00",
		X"77",X"03",X"10",X"14",X"28",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"10",X"30",X"40",X"80",X"00",X"00",X"00",X"08",X"80",X"08",X"06",X"01",X"00",X"00",X"00",
		X"04",X"04",X"08",X"00",X"08",X"08",X"04",X"04",X"0E",X"08",X"0E",X"0F",X"0D",X"0C",X"0C",X"04",
		X"06",X"06",X"06",X"0E",X"0E",X"06",X"00",X"00",X"33",X"00",X"00",X"03",X"00",X"22",X"22",X"13",
		X"08",X"00",X"00",X"80",X"40",X"00",X"00",X"00",X"88",X"EC",X"3A",X"15",X"03",X"00",X"00",X"00",
		X"00",X"00",X"CC",X"F3",X"03",X"0C",X"00",X"00",X"77",X"45",X"12",X"1C",X"00",X"00",X"00",X"00",
		X"00",X"11",X"00",X"00",X"90",X"E9",X"5A",X"F1",X"00",X"66",X"11",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"EE",X"11",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"98",X"A9",X"D2",
		X"F2",X"F0",X"E1",X"A1",X"43",X"87",X"0F",X"07",X"00",X"00",X"00",X"00",X"88",X"44",X"21",X"30",
		X"10",X"21",X"53",X"21",X"10",X"21",X"D2",X"B4",X"2C",X"DC",X"98",X"BA",X"F1",X"5E",X"A4",X"8E",
		X"22",X"44",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"CC",X"7C",X"C3",X"FC",X"B4",
		X"00",X"00",X"00",X"00",X"80",X"E8",X"BC",X"87",X"00",X"00",X"00",X"00",X"11",X"66",X"4C",X"0E",
		X"11",X"22",X"44",X"08",X"00",X"00",X"00",X"00",X"68",X"48",X"C0",X"08",X"19",X"93",X"93",X"0F",
		X"E0",X"51",X"32",X"BA",X"DF",X"BC",X"3C",X"F8",X"C2",X"E1",X"E9",X"D2",X"A5",X"A5",X"A4",X"68",
		X"03",X"07",X"0F",X"04",X"0F",X"C3",X"C3",X"A5",X"10",X"10",X"21",X"21",X"10",X"00",X"00",X"00",
		X"7B",X"7A",X"F4",X"79",X"B4",X"43",X"30",X"00",X"03",X"80",X"C0",X"4A",X"B4",X"69",X"B4",X"9E",
		X"E1",X"F0",X"3E",X"D3",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"11",X"11",X"33",X"22",X"44",X"88",X"E9",X"ED",X"B8",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"0B",X"09",X"03",X"01",X"0C",X"5B",X"E0",X"F0",
		X"E7",X"7B",X"68",X"C1",X"38",X"16",X"DF",X"FD",X"C0",X"80",X"80",X"C0",X"79",X"86",X"C2",X"68",
		X"00",X"00",X"00",X"00",X"88",X"CC",X"22",X"11",X"4B",X"78",X"90",X"00",X"88",X"88",X"88",X"00",
		X"F3",X"4B",X"F0",X"36",X"11",X"00",X"00",X"00",X"C8",X"C6",X"6B",X"97",X"0D",X"88",X"00",X"00",
		X"C8",X"00",X"00",X"11",X"11",X"22",X"22",X"01",X"C0",X"22",X"00",X"04",X"20",X"00",X"10",X"00",
		X"40",X"02",X"00",X"20",X"8C",X"46",X"46",X"23",X"00",X"00",X"00",X"24",X"22",X"00",X"00",X"0C",
		X"01",X"A1",X"44",X"20",X"80",X"04",X"80",X"54",X"00",X"00",X"00",X"45",X"08",X"00",X"10",X"00",
		X"00",X"40",X"08",X"00",X"04",X"33",X"00",X"00",X"02",X"07",X"37",X"04",X"04",X"80",X"54",X"02",
		X"11",X"22",X"40",X"22",X"66",X"00",X"00",X"18",X"44",X"44",X"80",X"11",X"00",X"CC",X"00",X"00",
		X"02",X"00",X"10",X"01",X"00",X"22",X"08",X"11",X"01",X"00",X"88",X"10",X"02",X"44",X"00",X"00",
		X"10",X"22",X"00",X"86",X"44",X"40",X"00",X"10",X"22",X"14",X"0C",X"00",X"A8",X"00",X"C1",X"C0",
		X"33",X"A3",X"47",X"04",X"00",X"58",X"68",X"40",X"22",X"00",X"00",X"00",X"00",X"13",X"80",X"00",
		X"10",X"22",X"10",X"54",X"10",X"80",X"00",X"30",X"00",X"22",X"00",X"80",X"88",X"00",X"01",X"00",
		X"20",X"00",X"08",X"04",X"00",X"88",X"41",X"03",X"40",X"51",X"40",X"10",X"06",X"04",X"28",X"FC",
		X"0C",X"00",X"11",X"11",X"02",X"04",X"88",X"00",X"44",X"22",X"00",X"00",X"11",X"20",X"00",X"00",
		X"91",X"00",X"21",X"82",X"08",X"11",X"22",X"22",X"88",X"00",X"10",X"00",X"80",X"00",X"00",X"00",
		X"03",X"04",X"80",X"00",X"00",X"98",X"33",X"00",X"22",X"11",X"44",X"02",X"00",X"06",X"02",X"01",
		X"91",X"04",X"04",X"18",X"00",X"44",X"18",X"26",X"44",X"CC",X"00",X"00",X"44",X"20",X"04",X"04",
		X"00",X"18",X"00",X"22",X"88",X"00",X"04",X"22",X"A0",X"08",X"00",X"00",X"88",X"00",X"01",X"03",
		X"04",X"10",X"00",X"C4",X"00",X"46",X"00",X"00",X"00",X"40",X"60",X"11",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
