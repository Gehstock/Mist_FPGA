library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity kbe3_IC6 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of kbe3_IC6 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"A9",X"99",X"98",X"87",X"76",X"66",X"66",X"78",X"9A",X"BC",X"CB",X"A9",X"87",X"66",X"68",X"99",
		X"AA",X"A9",X"87",X"77",X"77",X"89",X"AA",X"99",X"98",X"88",X"99",X"88",X"77",X"66",X"67",X"78",
		X"89",X"AB",X"CB",X"AA",X"98",X"77",X"78",X"89",X"9A",X"99",X"88",X"88",X"88",X"89",X"99",X"98",
		X"88",X"88",X"88",X"99",X"99",X"87",X"76",X"66",X"77",X"89",X"AA",X"BB",X"B9",X"98",X"77",X"77",
		X"89",X"9A",X"99",X"98",X"77",X"78",X"89",X"99",X"99",X"88",X"88",X"88",X"99",X"99",X"87",X"66",
		X"77",X"78",X"99",X"9A",X"AA",X"A9",X"98",X"88",X"78",X"88",X"99",X"99",X"98",X"88",X"88",X"89",
		X"99",X"99",X"88",X"88",X"88",X"99",X"99",X"88",X"87",X"77",X"78",X"88",X"88",X"99",X"9A",X"AA",
		X"99",X"88",X"77",X"78",X"99",X"99",X"99",X"88",X"88",X"88",X"99",X"99",X"98",X"88",X"88",X"88",
		X"89",X"99",X"99",X"98",X"87",X"77",X"77",X"78",X"89",X"99",X"AA",X"AA",X"98",X"87",X"77",X"78",
		X"88",X"88",X"88",X"98",X"88",X"88",X"99",X"98",X"88",X"87",X"89",X"AA",X"A9",X"76",X"66",X"8C",
		X"EC",X"96",X"44",X"68",X"DF",X"D8",X"63",X"46",X"8D",X"FC",X"76",X"43",X"7A",X"9D",X"D9",X"67",
		X"44",X"8A",X"8D",X"D9",X"66",X"35",X"A9",X"BE",X"B6",X"65",X"48",X"B8",X"DC",X"96",X"64",X"69",
		X"9A",X"EC",X"86",X"54",X"8B",X"8D",X"D8",X"56",X"46",X"A9",X"BE",X"A6",X"64",X"5A",X"A7",X"EB",
		X"77",X"64",X"7B",X"7D",X"E8",X"57",X"37",X"C8",X"AF",X"95",X"74",X"4A",X"A9",X"FA",X"46",X"64",
		X"BB",X"5F",X"D5",X"58",X"37",X"C6",X"EF",X"63",X"84",X"7D",X"6A",X"F9",X"37",X"56",X"B7",X"BF",
		X"83",X"66",X"8D",X"59",X"F9",X"45",X"78",X"C5",X"BF",X"75",X"65",X"9C",X"3A",X"F7",X"47",X"6A",
		X"C2",X"CF",X"63",X"84",X"AC",X"3D",X"F4",X"27",X"7B",X"A4",X"FE",X"42",X"68",X"BA",X"9F",X"93",
		X"26",X"BD",X"4B",X"F8",X"33",X"5B",X"C6",X"FC",X"44",X"56",X"E7",X"5F",X"C4",X"35",X"7C",X"5C",
		X"F7",X"46",X"4A",X"B2",X"FE",X"54",X"77",X"B5",X"7F",X"95",X"56",X"9B",X"2F",X"D5",X"47",X"9D",
		X"55",X"F8",X"25",X"8A",X"B5",X"FA",X"43",X"69",X"E6",X"9F",X"73",X"47",X"DA",X"4F",X"A5",X"52",
		X"5F",X"8E",X"E3",X"47",X"5B",X"78",X"F8",X"35",X"48",X"D5",X"FF",X"54",X"44",X"B9",X"CF",X"42",
		X"87",X"97",X"7F",X"B3",X"45",X"6D",X"7F",X"C5",X"75",X"4A",X"6F",X"F4",X"17",X"88",X"47",X"FA",
		X"35",X"48",X"B6",X"FC",X"55",X"78",X"93",X"FE",X"64",X"67",X"B5",X"CF",X"48",X"55",X"B9",X"6F",
		X"64",X"57",X"9A",X"5F",X"91",X"64",X"6D",X"3F",X"F0",X"34",X"7C",X"58",X"F6",X"53",X"2A",X"A4",
		X"F8",X"37",X"49",X"A1",X"FF",X"46",X"47",X"C5",X"AF",X"67",X"47",X"C6",X"5F",X"96",X"54",X"BB",
		X"0F",X"F2",X"81",X"3F",X"82",X"F9",X"64",X"1C",X"D1",X"AF",X"7E",X"00",X"FE",X"1F",X"A7",X"D0",
		X"4F",X"4A",X"F2",X"D0",X"0F",X"90",X"F8",X"CC",X"08",X"E3",X"FF",X"2F",X"00",X"F9",X"2F",X"8E",
		X"D0",X"8B",X"5B",X"F2",X"F0",X"2E",X"83",X"F8",X"F6",X"0A",X"A6",X"FF",X"3F",X"02",X"EB",X"4F",
		X"9E",X"A0",X"89",X"5F",X"F1",X"F0",X"0C",X"B5",X"FB",X"8E",X"08",X"95",X"BF",X"6E",X"60",X"9A",
		X"5F",X"F3",X"F0",X"28",X"4E",X"F6",X"9B",X"0A",X"87",X"8F",X"8F",X"10",X"95",X"BF",X"F2",X"F1",
		X"0B",X"8C",X"8D",X"AF",X"05",X"78",X"CF",X"99",X"60",X"DA",X"C5",X"C8",X"F0",X"08",X"4D",X"DF",
		X"8C",X"07",X"8F",X"48",X"DC",X"D0",X"90",X"D5",X"FE",X"64",X"0A",X"DA",X"2F",X"5F",X"40",X"83",
		X"6C",X"FF",X"C0",X"0F",X"79",X"DB",X"4F",X"07",X"60",X"BF",X"F3",X"F0",X"97",X"DA",X"D5",X"CB",
		X"0F",X"0D",X"6F",X"9E",X"40",X"77",X"F3",X"F7",X"F3",X"37",X"4B",X"5F",X"5F",X"00",X"9B",X"87",
		X"F3",X"F0",X"59",X"08",X"EF",X"7F",X"05",X"79",X"8C",X"F6",X"F0",X"84",X"28",X"EF",X"3F",X"03",
		X"77",X"BB",X"F5",X"F1",X"55",X"1B",X"CF",X"BF",X"03",X"6B",X"A8",X"F5",X"F3",X"46",X"36",X"EF",
		X"1F",X"02",X"3A",X"78",X"FB",X"E6",X"24",X"46",X"BF",X"7F",X"81",X"0D",X"09",X"FD",X"FA",X"03",
		X"60",X"BF",X"FB",X"F0",X"29",X"07",X"CF",X"AF",X"35",X"33",X"49",X"FB",X"F8",X"40",X"32",X"9F",
		X"FB",X"E4",X"16",X"06",X"CF",X"FF",X"61",X"30",X"99",X"ED",X"FA",X"64",X"26",X"3E",X"EE",X"B6",
		X"36",X"66",X"D7",X"F8",X"B5",X"47",X"5B",X"CB",X"6A",X"76",X"88",X"69",X"A9",X"C8",X"57",X"88",
		X"89",X"88",X"9B",X"79",X"A5",X"9A",X"88",X"A5",X"9A",X"87",X"87",X"9C",X"79",X"89",X"69",X"88",
		X"88",X"A8",X"C6",X"77",X"6B",X"98",X"9A",X"5A",X"65",X"A9",X"B8",X"A5",X"B6",X"68",X"9B",X"7C",
		X"89",X"77",X"49",X"E7",X"C7",X"88",X"95",X"7A",X"9D",X"99",X"76",X"55",X"BA",X"D9",X"B5",X"87",
		X"27",X"AE",X"EB",X"54",X"86",X"67",X"DD",X"C7",X"77",X"43",X"7C",X"FD",X"A5",X"67",X"55",X"7D",
		X"DC",X"D6",X"05",X"84",X"AE",X"DC",X"95",X"27",X"36",X"BF",X"FA",X"71",X"65",X"66",X"FD",X"FB",
		X"51",X"27",X"5B",X"FF",X"B8",X"32",X"44",X"7D",X"FF",X"B3",X"23",X"65",X"9F",X"FF",X"84",X"03",
		X"57",X"DF",X"F7",X"53",X"34",X"77",X"FF",X"D8",X"32",X"27",X"7B",X"FE",X"C7",X"30",X"69",X"5E",
		X"FE",X"75",X"03",X"77",X"9F",X"FD",X"61",X"15",X"78",X"CF",X"CB",X"70",X"09",X"94",X"FF",X"E6",
		X"20",X"38",X"B8",X"FF",X"D1",X"13",X"58",X"8D",X"FD",X"86",X"01",X"AA",X"6D",X"FC",X"83",X"03",
		X"AA",X"5F",X"FA",X"42",X"16",X"A7",X"AF",X"F9",X"51",X"19",X"A7",X"AF",X"E7",X"41",X"2A",X"A4",
		X"FF",X"B6",X"30",X"3D",X"A6",X"FF",X"85",X"30",X"5C",X"97",X"FF",X"62",X"02",X"9C",X"7B",X"FB",
		X"46",X"00",X"DD",X"6C",X"F8",X"44",X"03",X"CE",X"7E",X"F6",X"14",X"28",X"E9",X"4F",X"F2",X"64",
		X"0C",X"F6",X"5F",X"D1",X"94",X"0B",X"F7",X"5F",X"C0",X"64",X"6C",X"D3",X"6F",X"93",X"A1",X"3F",
		X"B1",X"BF",X"44",X"B0",X"5E",X"D0",X"BF",X"13",X"B3",X"7F",X"70",X"FF",X"07",X"80",X"BF",X"70",
		X"FF",X"2B",X"60",X"CD",X"52",X"FC",X"09",X"73",X"DB",X"32",X"F7",X"2B",X"37",X"F9",X"07",X"F7",
		X"4B",X"19",X"F7",X"18",X"F4",X"99",X"1B",X"A9",X"0A",X"F5",X"78",X"4B",X"C4",X"0F",X"F1",X"99",
		X"2D",X"B3",X"0F",X"F4",X"A5",X"6B",X"96",X"0F",X"E2",X"97",X"3D",X"C0",X"3F",X"82",X"F4",X"1F",
		X"90",X"AF",X"06",X"F0",X"3F",X"90",X"FF",X"0A",X"E0",X"AE",X"00",X"FF",X"0E",X"A0",X"DD",X"04",
		X"FF",X"2F",X"40",X"FA",X"0E",X"F1",X"6F",X"05",X"F1",X"0F",X"F0",X"CC",X"09",X"F0",X"3F",X"F4",
		X"C6",X"0D",X"F0",X"AF",X"45",X"E3",X"0F",X"40",X"FF",X"0C",X"C0",X"6F",X"00",X"FF",X"2C",X"70",
		X"9F",X"06",X"FF",X"3E",X"50",X"F9",X"0F",X"F0",X"8E",X"02",X"F4",X"0F",X"F0",X"B8",X"08",X"F0",
		X"1F",X"F2",X"B6",X"0E",X"C0",X"FF",X"F4",X"C1",X"1F",X"A0",X"FF",X"16",X"B0",X"4F",X"50",X"FF",
		X"09",X"B0",X"AF",X"08",X"FF",X"1B",X"50",X"CC",X"0F",X"F4",X"3B",X"30",X"FA",X"0F",X"F0",X"4E",
		X"06",X"F1",X"2F",X"F0",X"A9",X"0A",X"E0",X"9F",X"50",X"97",X"0C",X"E0",X"FF",X"20",X"D4",X"3E",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
