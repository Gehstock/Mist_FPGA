library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity burger_time_sound_prog is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of burger_time_sound_prog is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"4C",X"7A",X"F0",X"4C",X"09",X"F0",X"4C",X"55",X"F2",X"78",X"D8",X"A2",X"FF",X"9A",X"A2",X"EF",
		X"A9",X"00",X"95",X"00",X"CA",X"D0",X"FB",X"20",X"2A",X"F0",X"A9",X"08",X"85",X"1E",X"A9",X"FF",
		X"8D",X"00",X"C0",X"58",X"20",X"4A",X"F0",X"4C",X"27",X"F0",X"A9",X"00",X"85",X"05",X"AA",X"A5",
		X"05",X"8D",X"00",X"40",X"8D",X"00",X"80",X"BD",X"64",X"F0",X"8D",X"00",X"20",X"8D",X"00",X"60",
		X"E8",X"E6",X"05",X"A5",X"05",X"C9",X"10",X"90",X"E6",X"60",X"A9",X"00",X"85",X"05",X"AA",X"A5",
		X"05",X"8D",X"00",X"80",X"BD",X"64",X"F0",X"8D",X"00",X"60",X"E8",X"E6",X"05",X"A5",X"05",X"C9",
		X"0B",X"90",X"EC",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"68",X"A8",X"68",X"AA",X"68",X"40",X"48",X"8A",X"48",X"98",X"48",X"A5",
		X"01",X"F0",X"F1",X"A5",X"04",X"C9",X"05",X"D0",X"04",X"A9",X"00",X"85",X"04",X"E6",X"04",X"0A",
		X"AA",X"BD",X"9E",X"F0",X"85",X"1C",X"BD",X"9F",X"F0",X"85",X"1D",X"6C",X"1C",X"00",X"AA",X"F0",
		X"FE",X"F0",X"3F",X"F1",X"80",X"F1",X"74",X"F0",X"74",X"F0",X"A5",X"12",X"D0",X"38",X"A4",X"0C",
		X"E6",X"0C",X"B1",X"06",X"F0",X"3F",X"C9",X"FF",X"D0",X"07",X"A9",X"FF",X"85",X"15",X"4C",X"E9",
		X"F0",X"20",X"1E",X"F2",X"A9",X"00",X"8D",X"00",X"40",X"A5",X"1A",X"8D",X"00",X"20",X"A9",X"01",
		X"8D",X"00",X"40",X"A5",X"1B",X"8D",X"00",X"20",X"A5",X"1E",X"85",X"17",X"A9",X"08",X"8D",X"00",
		X"40",X"A5",X"17",X"8D",X"00",X"20",X"4C",X"74",X"F0",X"A9",X"0C",X"85",X"1E",X"A9",X"0B",X"85",
		X"20",X"A9",X"00",X"85",X"43",X"A9",X"00",X"85",X"1A",X"85",X"1B",X"4C",X"C4",X"F0",X"A5",X"15",
		X"D0",X"34",X"A5",X"13",X"D0",X"2D",X"A4",X"0D",X"E6",X"0D",X"B1",X"08",X"F0",X"28",X"20",X"1E",
		X"F2",X"A9",X"02",X"8D",X"00",X"40",X"A5",X"1A",X"8D",X"00",X"20",X"A9",X"03",X"8D",X"00",X"40",
		X"A5",X"1B",X"8D",X"00",X"20",X"A5",X"1F",X"85",X"18",X"A9",X"09",X"8D",X"00",X"40",X"A5",X"18",
		X"8D",X"00",X"20",X"4C",X"74",X"F0",X"A9",X"00",X"85",X"1A",X"85",X"1B",X"4C",X"11",X"F1",X"A5",
		X"15",X"D0",X"34",X"A5",X"14",X"D0",X"2D",X"A4",X"0E",X"E6",X"0E",X"B1",X"0A",X"F0",X"28",X"20",
		X"1E",X"F2",X"A9",X"04",X"8D",X"00",X"40",X"A5",X"1A",X"8D",X"00",X"20",X"A9",X"05",X"8D",X"00",
		X"40",X"A5",X"1B",X"8D",X"00",X"20",X"A5",X"20",X"85",X"19",X"A9",X"0A",X"8D",X"00",X"40",X"A5",
		X"19",X"8D",X"00",X"20",X"4C",X"74",X"F0",X"A9",X"00",X"85",X"1A",X"85",X"1B",X"4C",X"52",X"F1",
		X"4C",X"8C",X"F1",X"4C",X"DE",X"F1",X"4C",X"FE",X"F1",X"4C",X"74",X"F0",X"A5",X"15",X"D0",X"20",
		X"A5",X"0F",X"D0",X"0F",X"A4",X"0C",X"B1",X"06",X"85",X"0F",X"E6",X"0C",X"A9",X"FF",X"85",X"12",
		X"4C",X"83",X"F1",X"C6",X"0F",X"A5",X"0F",X"D0",X"F7",X"A9",X"00",X"85",X"12",X"4C",X"A0",X"F1",
		X"A9",X"00",X"AA",X"95",X"0C",X"E8",X"E0",X"0B",X"D0",X"F9",X"A2",X"00",X"A5",X"03",X"D0",X"0D",
		X"BD",X"80",X"F3",X"95",X"06",X"E8",X"E0",X"06",X"D0",X"F6",X"4C",X"89",X"F1",X"BD",X"86",X"F3",
		X"95",X"06",X"E8",X"E0",X"06",X"D0",X"F6",X"A9",X"0C",X"85",X"1F",X"4C",X"89",X"F1",X"A5",X"10",
		X"D0",X"0F",X"A4",X"0D",X"B1",X"08",X"85",X"10",X"E6",X"0D",X"A9",X"FF",X"85",X"13",X"4C",X"86",
		X"F1",X"C6",X"10",X"A5",X"10",X"D0",X"F7",X"A9",X"00",X"85",X"13",X"4C",X"EE",X"F1",X"A5",X"11",
		X"D0",X"0F",X"A4",X"0E",X"B1",X"0A",X"85",X"11",X"E6",X"0E",X"A9",X"FF",X"85",X"14",X"4C",X"89",
		X"F1",X"C6",X"11",X"A5",X"11",X"D0",X"F7",X"A9",X"00",X"85",X"14",X"4C",X"0E",X"F2",X"48",X"29",
		X"0F",X"AA",X"BD",X"3D",X"F2",X"85",X"1A",X"BD",X"49",X"F2",X"85",X"1B",X"68",X"4A",X"4A",X"4A",
		X"4A",X"F0",X"09",X"AA",X"18",X"46",X"1B",X"66",X"1A",X"CA",X"D0",X"F8",X"60",X"F2",X"1B",X"51",
		X"91",X"DD",X"32",X"91",X"F9",X"6A",X"E3",X"63",X"EB",X"0E",X"0E",X"0D",X"0C",X"0B",X"0B",X"0A",
		X"09",X"09",X"08",X"08",X"07",X"48",X"8A",X"48",X"98",X"48",X"AD",X"00",X"A0",X"85",X"3D",X"29",
		X"F0",X"F0",X"34",X"C9",X"10",X"D0",X"2D",X"A5",X"3D",X"29",X"0F",X"F0",X"27",X"C9",X"0F",X"B0",
		X"23",X"AA",X"A5",X"3E",X"DD",X"C6",X"F2",X"F0",X"02",X"B0",X"19",X"BD",X"C6",X"F2",X"85",X"3E",
		X"8A",X"0A",X"AA",X"BD",X"E1",X"F2",X"85",X"3F",X"BD",X"E2",X"F2",X"85",X"40",X"A2",X"FF",X"9A",
		X"58",X"6C",X"3F",X"00",X"4C",X"74",X"F0",X"A5",X"01",X"85",X"02",X"A9",X"00",X"85",X"01",X"A9",
		X"0F",X"85",X"1E",X"A9",X"0E",X"85",X"1F",X"A9",X"0E",X"85",X"20",X"A5",X"3D",X"0A",X"C9",X"0C",
		X"90",X"03",X"4C",X"FF",X"F2",X"AA",X"BD",X"D5",X"F2",X"85",X"41",X"BD",X"D6",X"F2",X"85",X"42",
		X"20",X"06",X"F3",X"6C",X"41",X"00",X"00",X"03",X"03",X"02",X"07",X"04",X"09",X"09",X"06",X"0A",
		X"08",X"0C",X"0B",X"05",X"01",X"09",X"F0",X"8C",X"F3",X"AA",X"F3",X"30",X"F3",X"30",X"F3",X"58",
		X"F3",X"74",X"F0",X"3A",X"F6",X"DB",X"F3",X"12",X"F4",X"33",X"F6",X"49",X"F4",X"AE",X"F4",X"41",
		X"F6",X"D8",X"F6",X"48",X"F6",X"4F",X"F6",X"60",X"F5",X"56",X"F6",X"EF",X"F4",X"5D",X"F6",X"A5",
		X"02",X"85",X"01",X"4C",X"74",X"F0",X"A9",X"07",X"8D",X"00",X"40",X"A9",X"F8",X"8D",X"00",X"20",
		X"60",X"A9",X"08",X"8D",X"00",X"40",X"A5",X"1E",X"8D",X"00",X"20",X"A9",X"09",X"8D",X"00",X"40",
		X"A5",X"1F",X"8D",X"00",X"20",X"A9",X"0A",X"8D",X"00",X"40",X"A5",X"20",X"8D",X"00",X"20",X"60",
		X"A9",X"00",X"85",X"03",X"A5",X"43",X"D0",X"C7",X"A2",X"00",X"BD",X"80",X"F3",X"95",X"06",X"E8",
		X"E0",X"06",X"D0",X"F6",X"A9",X"0C",X"85",X"1E",X"A9",X"00",X"85",X"1F",X"A9",X"0B",X"85",X"20",
		X"85",X"01",X"20",X"11",X"F3",X"4C",X"74",X"F0",X"A9",X"FF",X"85",X"03",X"A5",X"43",X"D0",X"9F",
		X"A2",X"00",X"BD",X"86",X"F3",X"95",X"06",X"E8",X"E0",X"06",X"D0",X"F6",X"A9",X"0C",X"85",X"1E",
		X"A9",X"0C",X"85",X"1F",X"A9",X"0B",X"85",X"20",X"85",X"01",X"20",X"11",X"F3",X"4C",X"74",X"F0",
		X"F9",X"F8",X"8A",X"F9",X"9C",X"F9",X"F9",X"F8",X"0A",X"FA",X"9C",X"F9",X"20",X"C8",X"F3",X"A2",
		X"00",X"BD",X"A4",X"F3",X"95",X"06",X"E8",X"E0",X"06",X"D0",X"F6",X"A9",X"0F",X"85",X"01",X"85",
		X"43",X"4C",X"74",X"F0",X"A3",X"F7",X"D4",X"F7",X"04",X"F8",X"20",X"C8",X"F3",X"A2",X"00",X"BD",
		X"C2",X"F3",X"95",X"06",X"E8",X"E0",X"06",X"D0",X"F6",X"A9",X"0F",X"85",X"01",X"85",X"43",X"4C",
		X"74",X"F0",X"42",X"F8",X"A1",X"F8",X"C3",X"F8",X"20",X"2A",X"F0",X"20",X"06",X"F3",X"A2",X"00",
		X"8A",X"85",X"04",X"95",X"0C",X"E8",X"E0",X"0B",X"D0",X"F9",X"60",X"20",X"68",X"F7",X"A0",X"20",
		X"A9",X"24",X"20",X"53",X"F7",X"A9",X"D2",X"85",X"2F",X"A9",X"F5",X"85",X"30",X"A9",X"00",X"85",
		X"25",X"A9",X"00",X"85",X"29",X"A9",X"08",X"85",X"2A",X"20",X"A4",X"F5",X"A5",X"22",X"C9",X"FF",
		X"F0",X"06",X"20",X"B8",X"F5",X"4C",X"F9",X"F3",X"20",X"68",X"F7",X"A9",X"00",X"85",X"3E",X"4C",
		X"23",X"F0",X"20",X"68",X"F7",X"A0",X"0C",X"A9",X"10",X"20",X"53",X"F7",X"A9",X"07",X"85",X"2F",
		X"A9",X"F6",X"85",X"30",X"A9",X"00",X"85",X"25",X"A9",X"02",X"85",X"29",X"A9",X"09",X"85",X"2A",
		X"20",X"A4",X"F5",X"A5",X"22",X"C9",X"FF",X"F0",X"06",X"20",X"B8",X"F5",X"4C",X"30",X"F4",X"20",
		X"68",X"F7",X"A9",X"00",X"85",X"3E",X"4C",X"23",X"F0",X"20",X"68",X"F7",X"A0",X"24",X"A9",X"2A",
		X"20",X"53",X"F7",X"A9",X"10",X"85",X"27",X"A9",X"0F",X"85",X"22",X"A9",X"57",X"85",X"2B",X"A9",
		X"74",X"85",X"2D",X"A5",X"2B",X"38",X"E9",X"0F",X"85",X"2B",X"A5",X"2D",X"38",X"E9",X"06",X"85",
		X"2D",X"20",X"75",X"F7",X"A9",X"09",X"85",X"21",X"20",X"83",X"F7",X"E6",X"21",X"20",X"83",X"F7",
		X"A0",X"02",X"20",X"8E",X"F7",X"E6",X"2B",X"E6",X"2D",X"E6",X"2D",X"E6",X"2D",X"20",X"75",X"F7",
		X"A0",X"01",X"20",X"8E",X"F7",X"A5",X"27",X"29",X"01",X"F0",X"02",X"C6",X"22",X"C6",X"27",X"F0",
		X"03",X"4C",X"63",X"F4",X"20",X"68",X"F7",X"A9",X"00",X"85",X"3E",X"4C",X"23",X"F0",X"20",X"68",
		X"F7",X"A0",X"10",X"A9",X"14",X"20",X"53",X"F7",X"A9",X"03",X"85",X"27",X"85",X"23",X"A9",X"02",
		X"85",X"29",X"A9",X"09",X"85",X"2A",X"A9",X"07",X"85",X"22",X"20",X"B8",X"F5",X"E6",X"22",X"A5",
		X"22",X"C9",X"0F",X"D0",X"F5",X"A9",X"00",X"85",X"22",X"20",X"B8",X"F5",X"A0",X"0F",X"20",X"8E",
		X"F7",X"C6",X"27",X"D0",X"E1",X"20",X"68",X"F7",X"A9",X"00",X"85",X"3E",X"4C",X"23",X"F0",X"20",
		X"68",X"F7",X"A0",X"2A",X"A9",X"36",X"20",X"53",X"F7",X"A9",X"01",X"85",X"27",X"A9",X"00",X"85",
		X"22",X"20",X"27",X"F5",X"38",X"A5",X"2B",X"E9",X"20",X"85",X"2D",X"20",X"75",X"F7",X"A4",X"21",
		X"20",X"8E",X"F7",X"A5",X"2B",X"C9",X"00",X"D0",X"E8",X"C6",X"27",X"D0",X"E0",X"20",X"68",X"F7",
		X"A9",X"00",X"85",X"3E",X"4C",X"23",X"F0",X"A6",X"22",X"BD",X"38",X"F5",X"85",X"2B",X"E8",X"BD",
		X"38",X"F5",X"85",X"21",X"E8",X"86",X"22",X"60",X"29",X"08",X"2C",X"08",X"2E",X"08",X"34",X"08",
		X"37",X"08",X"3A",X"08",X"3F",X"08",X"47",X"08",X"52",X"08",X"58",X"08",X"60",X"08",X"68",X"08",
		X"74",X"08",X"80",X"08",X"90",X"08",X"A0",X"08",X"B4",X"08",X"D0",X"08",X"F0",X"08",X"00",X"01",
		X"20",X"68",X"F7",X"A0",X"00",X"A9",X"0C",X"20",X"53",X"F7",X"A9",X"E0",X"85",X"2B",X"A9",X"90",
		X"85",X"2D",X"A5",X"2B",X"38",X"E9",X"04",X"85",X"2B",X"A5",X"2D",X"38",X"E9",X"04",X"85",X"2D",
		X"20",X"75",X"F7",X"A0",X"01",X"20",X"8E",X"F7",X"E6",X"2B",X"E6",X"2D",X"20",X"75",X"F7",X"A0",
		X"01",X"20",X"8E",X"F7",X"A5",X"2B",X"C9",X"64",X"D0",X"D8",X"20",X"68",X"F7",X"A9",X"00",X"85",
		X"3E",X"4C",X"23",X"F0",X"A6",X"25",X"A4",X"26",X"B1",X"2F",X"95",X"21",X"E6",X"26",X"E8",X"E0",
		X"03",X"D0",X"F3",X"A2",X"00",X"86",X"25",X"60",X"A5",X"29",X"8D",X"00",X"80",X"A5",X"21",X"8D",
		X"00",X"60",X"A5",X"2A",X"8D",X"00",X"80",X"A5",X"22",X"8D",X"00",X"60",X"A4",X"23",X"20",X"8E",
		X"F7",X"60",X"E0",X"0F",X"04",X"E2",X"0F",X"04",X"E0",X"0E",X"03",X"E2",X"0E",X"03",X"E0",X"0D",
		X"03",X"E2",X"0D",X"02",X"E0",X"0C",X"02",X"E2",X"0C",X"02",X"20",X"09",X"01",X"22",X"08",X"01",
		X"00",X"09",X"01",X"00",X"09",X"01",X"20",X"09",X"01",X"FF",X"0F",X"0A",X"FD",X"0D",X"02",X"FF",
		X"0A",X"02",X"FD",X"08",X"02",X"FF",X"FF",X"E0",X"0E",X"0E",X"E2",X"0E",X"0E",X"E0",X"0D",X"0D",
		X"E2",X"0D",X"0D",X"E0",X"0C",X"0D",X"E2",X"0C",X"0D",X"E0",X"0B",X"0D",X"E2",X"0B",X"0D",X"E0",
		X"0A",X"07",X"E2",X"0A",X"07",X"E0",X"09",X"07",X"E2",X"07",X"03",X"DE",X"08",X"03",X"DD",X"08",
		X"03",X"FF",X"FF",X"A9",X"05",X"85",X"44",X"4C",X"64",X"F6",X"A9",X"04",X"85",X"44",X"4C",X"64",
		X"F6",X"A9",X"01",X"85",X"44",X"4C",X"64",X"F6",X"A9",X"00",X"85",X"44",X"4C",X"64",X"F6",X"A9",
		X"02",X"85",X"44",X"4C",X"64",X"F6",X"A9",X"06",X"85",X"44",X"4C",X"64",X"F6",X"A9",X"03",X"85",
		X"44",X"4C",X"64",X"F6",X"20",X"68",X"F7",X"A5",X"44",X"0A",X"AA",X"BD",X"A8",X"FA",X"85",X"45",
		X"BD",X"A9",X"FA",X"85",X"46",X"BD",X"9A",X"FA",X"85",X"47",X"BD",X"9B",X"FA",X"85",X"48",X"A0",
		X"00",X"B1",X"45",X"8D",X"00",X"80",X"C8",X"B1",X"45",X"8D",X"00",X"60",X"C8",X"B1",X"45",X"C9",
		X"80",X"D0",X"EE",X"C8",X"84",X"26",X"A0",X"00",X"A9",X"00",X"8D",X"00",X"80",X"B1",X"47",X"8D",
		X"00",X"60",X"C8",X"A9",X"02",X"8D",X"00",X"80",X"B1",X"47",X"8D",X"00",X"60",X"20",X"C1",X"F6",
		X"C8",X"B1",X"47",X"C9",X"81",X"D0",X"E1",X"20",X"68",X"F7",X"A9",X"00",X"85",X"3E",X"4C",X"23",
		X"F0",X"98",X"48",X"A4",X"26",X"B1",X"45",X"85",X"21",X"A9",X"FC",X"85",X"22",X"C6",X"22",X"D0",
		X"FC",X"C6",X"21",X"D0",X"F8",X"68",X"A8",X"60",X"20",X"68",X"F7",X"A0",X"00",X"A9",X"0C",X"20",
		X"53",X"F7",X"A9",X"E3",X"85",X"2B",X"A9",X"A0",X"85",X"2D",X"A5",X"2B",X"38",X"E9",X"04",X"85",
		X"2B",X"A5",X"2D",X"38",X"E9",X"03",X"85",X"2D",X"20",X"75",X"F7",X"A0",X"01",X"20",X"8E",X"F7",
		X"18",X"E6",X"2B",X"E6",X"2D",X"20",X"75",X"F7",X"A0",X"01",X"20",X"8E",X"F7",X"A5",X"2B",X"C9",
		X"30",X"B0",X"D7",X"20",X"68",X"F7",X"A9",X"00",X"85",X"3E",X"4C",X"23",X"F0",X"07",X"F9",X"09",
		X"1D",X"0A",X"1D",X"0B",X"00",X"0C",X"40",X"0D",X"09",X"07",X"FD",X"03",X"02",X"06",X"0F",X"07",
		X"EF",X"07",X"F9",X"09",X"10",X"0A",X"10",X"0B",X"00",X"0D",X"09",X"0C",X"40",X"07",X"FE",X"01",
		X"03",X"07",X"F9",X"03",X"01",X"05",X"01",X"07",X"F9",X"09",X"10",X"0A",X"10",X"0B",X"00",X"0C",
		X"37",X"0D",X"09",X"85",X"31",X"B9",X"1D",X"F7",X"8D",X"00",X"80",X"C8",X"B9",X"1D",X"F7",X"8D",
		X"00",X"60",X"C8",X"C4",X"31",X"D0",X"EE",X"60",X"A9",X"00",X"A2",X"10",X"95",X"21",X"CA",X"10",
		X"FB",X"20",X"4A",X"F0",X"60",X"A2",X"05",X"B5",X"29",X"8E",X"00",X"80",X"8D",X"00",X"60",X"CA",
		X"10",X"F5",X"60",X"A5",X"21",X"8D",X"00",X"80",X"A5",X"22",X"8D",X"00",X"60",X"60",X"A9",X"F0",
		X"85",X"32",X"20",X"99",X"F7",X"88",X"D0",X"F6",X"60",X"A2",X"00",X"CA",X"D0",X"FD",X"C6",X"32",
		X"10",X"F9",X"60",X"44",X"20",X"47",X"0E",X"00",X"0A",X"47",X"28",X"45",X"10",X"44",X"10",X"45",
		X"20",X"49",X"0E",X"00",X"0A",X"49",X"28",X"47",X"10",X"45",X"10",X"47",X"20",X"4B",X"0E",X"00",
		X"0A",X"4B",X"28",X"49",X"10",X"4B",X"10",X"50",X"18",X"47",X"08",X"49",X"18",X"47",X"08",X"00",
		X"40",X"00",X"FF",X"FF",X"40",X"20",X"44",X"0E",X"00",X"0A",X"44",X"28",X"42",X"10",X"40",X"10",
		X"42",X"20",X"45",X"0E",X"00",X"0A",X"45",X"28",X"44",X"10",X"42",X"10",X"44",X"20",X"47",X"0E",
		X"00",X"0A",X"47",X"28",X"45",X"10",X"47",X"10",X"47",X"18",X"44",X"08",X"45",X"18",X"44",X"08",
		X"00",X"40",X"00",X"FF",X"30",X"10",X"00",X"10",X"34",X"10",X"00",X"10",X"37",X"10",X"00",X"10",
		X"40",X"10",X"00",X"10",X"32",X"10",X"00",X"10",X"35",X"10",X"00",X"10",X"39",X"10",X"00",X"10",
		X"42",X"10",X"00",X"10",X"3B",X"10",X"00",X"10",X"32",X"10",X"00",X"10",X"35",X"10",X"00",X"10",
		X"37",X"10",X"00",X"10",X"40",X"10",X"00",X"10",X"39",X"10",X"00",X"10",X"37",X"10",X"00",X"30",
		X"00",X"FF",X"44",X"2A",X"00",X"02",X"37",X"09",X"00",X"02",X"39",X"09",X"00",X"0D",X"40",X"09",
		X"00",X"02",X"45",X"2A",X"00",X"02",X"44",X"2A",X"00",X"02",X"42",X"1F",X"00",X"02",X"41",X"09",
		X"00",X"02",X"42",X"09",X"00",X"02",X"00",X"16",X"49",X"2A",X"00",X"02",X"47",X"09",X"00",X"02",
		X"45",X"1F",X"00",X"02",X"44",X"09",X"00",X"02",X"00",X"16",X"47",X"14",X"00",X"02",X"47",X"1D",
		X"00",X"04",X"47",X"09",X"00",X"02",X"49",X"2A",X"00",X"02",X"4B",X"2A",X"00",X"02",X"50",X"1F",
		X"00",X"02",X"47",X"09",X"00",X"02",X"4B",X"1D",X"00",X"04",X"50",X"09",X"00",X"5A",X"00",X"FF",
		X"FF",X"00",X"58",X"42",X"2A",X"00",X"02",X"40",X"2A",X"00",X"B2",X"44",X"14",X"00",X"02",X"44",
		X"1D",X"00",X"04",X"44",X"09",X"00",X"02",X"45",X"2A",X"00",X"02",X"47",X"2A",X"00",X"4F",X"00",
		X"FF",X"00",X"FF",X"30",X"24",X"00",X"08",X"30",X"24",X"00",X"08",X"32",X"24",X"00",X"08",X"34",
		X"24",X"00",X"08",X"35",X"24",X"00",X"08",X"35",X"24",X"00",X"08",X"35",X"24",X"00",X"08",X"35",
		X"24",X"00",X"08",X"34",X"24",X"00",X"08",X"34",X"24",X"00",X"08",X"32",X"24",X"00",X"08",X"32",
		X"24",X"00",X"08",X"30",X"24",X"00",X"8C",X"00",X"FF",X"4A",X"0D",X"00",X"05",X"4A",X"0D",X"00",
		X"05",X"4B",X"0D",X"00",X"05",X"4B",X"0D",X"00",X"05",X"50",X"0D",X"00",X"05",X"50",X"0D",X"00",
		X"05",X"51",X"0D",X"00",X"05",X"51",X"0D",X"00",X"05",X"52",X"0E",X"00",X"16",X"49",X"0E",X"00",
		X"16",X"52",X"0E",X"00",X"16",X"49",X"0E",X"00",X"16",X"50",X"0D",X"00",X"05",X"55",X"0D",X"00",
		X"05",X"54",X"0D",X"00",X"05",X"52",X"0D",X"00",X"05",X"50",X"0D",X"00",X"05",X"4B",X"0D",X"00",
		X"05",X"50",X"0D",X"00",X"05",X"4B",X"0D",X"00",X"05",X"50",X"0E",X"00",X"16",X"55",X"0E",X"00",
		X"16",X"50",X"0E",X"00",X"16",X"55",X"0E",X"00",X"16",X"50",X"0E",X"00",X"16",X"59",X"0E",X"00",
		X"16",X"50",X"0E",X"00",X"16",X"59",X"0E",X"00",X"16",X"4A",X"10",X"00",X"14",X"57",X"0D",X"00",
		X"17",X"49",X"10",X"00",X"14",X"55",X"0D",X"00",X"17",X"4A",X"10",X"00",X"14",X"57",X"0D",X"00",
		X"17",X"49",X"10",X"00",X"14",X"55",X"0D",X"00",X"17",X"FF",X"00",X"20",X"00",X"90",X"00",X"90",
		X"00",X"90",X"00",X"90",X"00",X"90",X"00",X"90",X"00",X"98",X"00",X"F0",X"3A",X"0D",X"00",X"05",
		X"3A",X"0D",X"00",X"05",X"39",X"0D",X"00",X"05",X"39",X"0D",X"00",X"05",X"38",X"0D",X"00",X"05",
		X"38",X"0D",X"00",X"05",X"37",X"0D",X"00",X"05",X"37",X"0D",X"00",X"05",X"36",X"24",X"00",X"12",
		X"36",X"0D",X"00",X"05",X"36",X"1C",X"00",X"2C",X"35",X"12",X"00",X"12",X"37",X"12",X"00",X"12",
		X"39",X"0D",X"00",X"05",X"38",X"0D",X"00",X"05",X"39",X"0D",X"00",X"05",X"38",X"0D",X"00",X"05",
		X"39",X"24",X"00",X"12",X"39",X"0D",X"00",X"05",X"39",X"1C",X"00",X"2C",X"35",X"24",X"00",X"12",
		X"35",X"0D",X"00",X"05",X"35",X"1C",X"00",X"2C",X"37",X"12",X"00",X"36",X"35",X"12",X"00",X"36",
		X"37",X"12",X"00",X"36",X"35",X"12",X"00",X"36",X"00",X"F0",X"67",X"0D",X"00",X"05",X"64",X"0D",
		X"00",X"05",X"67",X"0D",X"00",X"05",X"64",X"0D",X"00",X"05",X"00",X"48",X"67",X"0D",X"00",X"05",
		X"64",X"0D",X"00",X"05",X"67",X"0D",X"00",X"05",X"64",X"0D",X"00",X"05",X"00",X"48",X"67",X"0D",
		X"00",X"05",X"64",X"0D",X"00",X"05",X"67",X"0D",X"00",X"05",X"64",X"0D",X"00",X"05",X"00",X"48",
		X"67",X"0D",X"00",X"05",X"64",X"0D",X"00",X"05",X"67",X"0D",X"00",X"05",X"64",X"0D",X"00",X"05",
		X"00",X"48",X"67",X"0D",X"00",X"05",X"64",X"0D",X"00",X"05",X"67",X"0D",X"00",X"05",X"64",X"0D",
		X"00",X"05",X"00",X"48",X"67",X"0D",X"00",X"05",X"64",X"0D",X"00",X"05",X"67",X"0D",X"00",X"05",
		X"64",X"0D",X"00",X"05",X"00",X"48",X"67",X"0D",X"00",X"05",X"64",X"0D",X"00",X"05",X"67",X"0D",
		X"00",X"05",X"64",X"0D",X"00",X"05",X"00",X"48",X"67",X"0D",X"00",X"05",X"64",X"0D",X"00",X"05",
		X"67",X"0D",X"00",X"05",X"64",X"0D",X"00",X"05",X"00",X"48",X"12",X"FB",X"3B",X"FB",X"49",X"FB",
		X"58",X"FB",X"DF",X"FB",X"EC",X"FB",X"15",X"FC",X"B6",X"FA",X"C2",X"FA",X"D6",X"FA",X"E2",X"FA",
		X"EE",X"FA",X"FA",X"FA",X"06",X"FB",X"07",X"F8",X"08",X"0F",X"09",X"0F",X"01",X"00",X"03",X"01",
		X"80",X"11",X"07",X"F8",X"08",X"10",X"09",X"10",X"0A",X"10",X"01",X"01",X"03",X"01",X"0B",X"04",
		X"0C",X"02",X"0D",X"0F",X"80",X"03",X"07",X"F8",X"08",X"0F",X"09",X"0F",X"01",X"00",X"03",X"00",
		X"80",X"0A",X"07",X"F8",X"08",X"0F",X"09",X"0F",X"01",X"00",X"03",X"00",X"80",X"0A",X"07",X"F8",
		X"08",X"0D",X"09",X"0B",X"01",X"01",X"03",X"03",X"80",X"08",X"07",X"F8",X"08",X"0F",X"09",X"0F",
		X"01",X"00",X"03",X"00",X"80",X"08",X"07",X"F8",X"08",X"0F",X"09",X"0F",X"01",X"00",X"03",X"00",
		X"80",X"0A",X"7E",X"FA",X"00",X"00",X"64",X"92",X"00",X"00",X"54",X"52",X"00",X"00",X"3F",X"FA",
		X"00",X"00",X"54",X"52",X"00",X"00",X"64",X"92",X"00",X"00",X"7E",X"FA",X"00",X"00",X"64",X"92",
		X"00",X"00",X"43",X"0C",X"00",X"00",X"3F",X"FA",X"3F",X"FA",X"81",X"43",X"2F",X"43",X"2F",X"43",
		X"2F",X"43",X"2F",X"43",X"2F",X"43",X"2F",X"43",X"81",X"C9",X"C9",X"00",X"00",X"C9",X"C9",X"00",
		X"00",X"A9",X"A9",X"00",X"00",X"64",X"64",X"81",X"A9",X"54",X"96",X"4B",X"86",X"43",X"A9",X"54",
		X"96",X"4B",X"86",X"43",X"7F",X"3F",X"A9",X"54",X"96",X"4B",X"86",X"43",X"7E",X"3F",X"A9",X"54",
		X"96",X"4B",X"86",X"43",X"A9",X"54",X"96",X"4B",X"86",X"43",X"7F",X"3F",X"A9",X"54",X"96",X"4B",
		X"86",X"43",X"7E",X"3F",X"A9",X"54",X"96",X"4B",X"86",X"43",X"A9",X"54",X"96",X"4B",X"86",X"43",
		X"7F",X"3F",X"A9",X"54",X"96",X"4B",X"86",X"43",X"7E",X"3F",X"A9",X"54",X"96",X"4B",X"86",X"43",
		X"A9",X"54",X"96",X"4B",X"86",X"43",X"7F",X"3F",X"A9",X"54",X"96",X"4B",X"86",X"43",X"7E",X"3F",
		X"A9",X"54",X"96",X"4B",X"86",X"43",X"A9",X"54",X"96",X"4B",X"86",X"43",X"7F",X"3F",X"A9",X"54",
		X"96",X"4B",X"86",X"43",X"7E",X"3F",X"A9",X"54",X"96",X"4B",X"86",X"43",X"A9",X"54",X"96",X"4B",
		X"86",X"43",X"7F",X"3F",X"A9",X"54",X"96",X"4B",X"86",X"43",X"7E",X"3F",X"00",X"00",X"81",X"FD",
		X"FD",X"FD",X"FD",X"FD",X"FD",X"A9",X"A9",X"A9",X"A9",X"A9",X"A9",X"81",X"54",X"2A",X"54",X"2A",
		X"00",X"00",X"54",X"2A",X"54",X"2A",X"00",X"00",X"64",X"32",X"64",X"32",X"00",X"00",X"64",X"32",
		X"64",X"32",X"00",X"00",X"7E",X"3F",X"7E",X"3F",X"00",X"00",X"7E",X"3F",X"7E",X"3F",X"00",X"00",
		X"7E",X"3F",X"7E",X"3F",X"81",X"A9",X"54",X"00",X"00",X"3F",X"2A",X"00",X"00",X"3F",X"2A",X"00",
		X"00",X"3F",X"2A",X"00",X"00",X"3F",X"2A",X"00",X"00",X"3F",X"2A",X"00",X"00",X"3F",X"2A",X"00",
		X"00",X"3F",X"2A",X"81",X"4C",X"EC",X"FC",X"78",X"D8",X"A2",X"FF",X"9A",X"AD",X"00",X"A0",X"A9",
		X"00",X"8D",X"00",X"C0",X"A0",X"00",X"A2",X"00",X"B9",X"55",X"F2",X"95",X"00",X"C8",X"E8",X"D0",
		X"F7",X"B9",X"55",X"F2",X"9D",X"00",X"01",X"C8",X"E8",X"D0",X"F6",X"B5",X"00",X"D9",X"55",X"F2",
		X"D0",X"D2",X"C8",X"E8",X"D0",X"F5",X"BD",X"00",X"01",X"D9",X"55",X"F2",X"D0",X"7E",X"C8",X"E8",
		X"D0",X"F4",X"C8",X"C0",X"20",X"D0",X"CF",X"A2",X"00",X"A0",X"00",X"98",X"85",X"49",X"A9",X"02",
		X"85",X"4A",X"BD",X"55",X"F2",X"91",X"49",X"E8",X"C8",X"D0",X"F7",X"E6",X"4A",X"A5",X"4A",X"C9",
		X"04",X"90",X"EF",X"A9",X"00",X"85",X"49",X"A9",X"02",X"85",X"4A",X"B1",X"49",X"DD",X"55",X"F2",
		X"D0",X"4A",X"E8",X"C8",X"D0",X"F5",X"E6",X"4A",X"A5",X"4A",X"C9",X"04",X"90",X"ED",X"E8",X"E0",
		X"20",X"D0",X"C6",X"A2",X"00",X"BD",X"D4",X"FC",X"8D",X"00",X"40",X"E8",X"BD",X"D4",X"FC",X"8D",
		X"00",X"20",X"E8",X"E0",X"18",X"D0",X"EE",X"A2",X"80",X"A0",X"00",X"88",X"D0",X"FD",X"CA",X"D0",
		X"FA",X"4C",X"03",X"F0",X"00",X"66",X"01",X"01",X"02",X"1C",X"03",X"01",X"04",X"EF",X"05",X"00",
		X"07",X"F8",X"08",X"10",X"09",X"10",X"0A",X"10",X"0C",X"30",X"0D",X"09",X"A0",X"00",X"B9",X"0D",
		X"FD",X"8D",X"00",X"40",X"C8",X"B9",X"0D",X"FD",X"8D",X"00",X"20",X"C8",X"C0",X"18",X"D0",X"EE",
		X"A2",X"A0",X"A0",X"00",X"88",X"D0",X"FD",X"CA",X"D0",X"FA",X"4C",X"EC",X"FC",X"00",X"CC",X"01",
		X"02",X"02",X"A4",X"03",X"02",X"04",X"7E",X"05",X"02",X"07",X"38",X"08",X"10",X"09",X"10",X"0A",
		X"10",X"0C",X"30",X"0D",X"09",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"F0",X"37",X"FC",X"06",X"F0");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
