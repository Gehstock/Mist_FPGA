library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity GFX1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of GFX1 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"CC",X"EE",X"11",X"11",X"33",X"EE",X"CC",X"00",X"11",X"33",X"66",X"44",X"44",X"33",X"11",X"00",
		X"11",X"11",X"FF",X"FF",X"11",X"11",X"00",X"00",X"00",X"00",X"77",X"77",X"22",X"00",X"00",X"00",
		X"11",X"99",X"DD",X"DD",X"FF",X"77",X"33",X"00",X"33",X"77",X"55",X"44",X"44",X"66",X"22",X"00",
		X"66",X"FF",X"99",X"99",X"99",X"33",X"22",X"00",X"44",X"66",X"77",X"55",X"44",X"44",X"00",X"00",
		X"44",X"FF",X"FF",X"44",X"44",X"CC",X"CC",X"00",X"00",X"77",X"77",X"66",X"33",X"11",X"00",X"00",
		X"EE",X"FF",X"11",X"11",X"11",X"33",X"22",X"00",X"00",X"55",X"55",X"55",X"55",X"77",X"77",X"00",
		X"66",X"FF",X"99",X"99",X"99",X"FF",X"EE",X"00",X"00",X"44",X"44",X"44",X"66",X"33",X"11",X"00",
		X"00",X"00",X"88",X"FF",X"77",X"00",X"00",X"00",X"66",X"77",X"55",X"44",X"44",X"66",X"66",X"00",
		X"66",X"77",X"DD",X"DD",X"99",X"99",X"66",X"00",X"00",X"33",X"44",X"44",X"55",X"77",X"33",X"00",
		X"CC",X"EE",X"BB",X"99",X"99",X"99",X"00",X"00",X"33",X"77",X"44",X"44",X"44",X"77",X"33",X"00",
		X"F0",X"F0",X"F0",X"FF",X"FF",X"F0",X"F0",X"F0",X"F1",X"F1",X"F1",X"FF",X"FF",X"F1",X"F1",X"F1",
		X"F0",X"F0",X"F0",X"FF",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F1",X"F1",X"F1",X"F1",X"F1",
		X"F0",X"F0",X"F0",X"FF",X"FF",X"F0",X"F0",X"F0",X"F1",X"F1",X"F1",X"F1",X"F1",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"FF",X"FF",X"F1",X"F1",X"F1",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F1",X"F1",X"F1",X"FF",X"FF",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",
		X"F0",X"F0",X"F0",X"FF",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"FF",X"FF",X"F0",X"F0",X"F0",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"26",X"79",X"5B",X"5B",X"79",X"26",X"00",X"00",X"00",X"11",X"77",X"77",X"11",X"00",X"00",
		X"00",X"66",X"66",X"00",X"00",X"66",X"66",X"00",X"00",X"66",X"66",X"00",X"00",X"66",X"66",X"00",
		X"FC",X"F2",X"F1",X"F5",X"F5",X"F9",X"F2",X"FC",X"F3",X"F4",X"F8",X"FA",X"FA",X"F9",X"F4",X"F3",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"EF",X"00",X"EF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"EF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"EF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"EF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"88",X"CC",X"22",X"22",X"66",X"CC",X"88",X"00",X"33",X"77",X"CC",X"88",X"88",X"77",X"33",X"00",
		X"22",X"22",X"EE",X"EE",X"22",X"22",X"00",X"00",X"00",X"00",X"FF",X"FF",X"44",X"00",X"00",X"00",
		X"22",X"22",X"AA",X"AA",X"EE",X"EE",X"66",X"00",X"66",X"FF",X"BB",X"99",X"99",X"CC",X"44",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"66",X"44",X"00",X"88",X"DD",X"FF",X"BB",X"99",X"88",X"00",X"00",
		X"88",X"EE",X"EE",X"88",X"88",X"88",X"88",X"00",X"00",X"FF",X"FF",X"CC",X"66",X"33",X"11",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"66",X"44",X"00",X"11",X"BB",X"AA",X"AA",X"AA",X"EE",X"EE",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"EE",X"CC",X"00",X"00",X"99",X"99",X"99",X"DD",X"77",X"33",X"00",
		X"00",X"00",X"00",X"EE",X"EE",X"00",X"00",X"00",X"CC",X"EE",X"BB",X"99",X"88",X"CC",X"CC",X"00",
		X"CC",X"EE",X"AA",X"AA",X"22",X"22",X"CC",X"00",X"00",X"66",X"99",X"99",X"BB",X"FF",X"66",X"00",
		X"88",X"CC",X"66",X"22",X"22",X"22",X"00",X"00",X"77",X"FF",X"99",X"99",X"99",X"FF",X"66",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"EE",X"88",X"88",X"88",X"EE",X"EE",X"00",X"33",X"77",X"CC",X"88",X"CC",X"77",X"33",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"EE",X"EE",X"00",X"66",X"FF",X"99",X"99",X"99",X"FF",X"FF",X"00",
		X"44",X"66",X"22",X"22",X"66",X"CC",X"88",X"00",X"44",X"CC",X"88",X"88",X"CC",X"77",X"33",X"00",
		X"88",X"CC",X"66",X"22",X"22",X"EE",X"EE",X"00",X"33",X"77",X"CC",X"88",X"88",X"FF",X"FF",X"00",
		X"22",X"22",X"22",X"22",X"EE",X"EE",X"00",X"00",X"88",X"99",X"99",X"99",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"00",X"88",X"99",X"99",X"99",X"99",X"FF",X"FF",X"00",
		X"EE",X"EE",X"22",X"22",X"66",X"CC",X"88",X"00",X"99",X"99",X"99",X"88",X"CC",X"77",X"33",X"00",
		X"EE",X"EE",X"00",X"00",X"00",X"EE",X"EE",X"00",X"FF",X"FF",X"11",X"11",X"11",X"FF",X"FF",X"00",
		X"22",X"22",X"EE",X"EE",X"22",X"22",X"00",X"00",X"88",X"88",X"FF",X"FF",X"88",X"88",X"00",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"66",X"44",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"22",X"66",X"EE",X"CC",X"88",X"EE",X"EE",X"00",X"88",X"CC",X"66",X"33",X"11",X"FF",X"FF",X"00",
		X"22",X"22",X"22",X"22",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"EE",X"EE",X"00",X"88",X"00",X"EE",X"EE",X"00",X"FF",X"FF",X"77",X"33",X"77",X"FF",X"FF",X"00",
		X"EE",X"EE",X"CC",X"88",X"00",X"EE",X"EE",X"00",X"FF",X"FF",X"11",X"33",X"77",X"FF",X"FF",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"EE",X"CC",X"00",X"77",X"FF",X"88",X"88",X"88",X"FF",X"77",X"00",
		X"00",X"88",X"88",X"88",X"88",X"EE",X"EE",X"00",X"77",X"FF",X"88",X"88",X"88",X"FF",X"FF",X"00",
		X"AA",X"CC",X"EE",X"AA",X"22",X"EE",X"CC",X"00",X"77",X"FF",X"88",X"88",X"88",X"FF",X"77",X"00",
		X"22",X"66",X"EE",X"CC",X"88",X"EE",X"EE",X"00",X"77",X"FF",X"99",X"88",X"88",X"FF",X"FF",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"66",X"44",X"00",X"00",X"55",X"DD",X"99",X"99",X"FF",X"66",X"00",
		X"00",X"00",X"EE",X"EE",X"00",X"00",X"00",X"00",X"88",X"88",X"FF",X"FF",X"88",X"88",X"00",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"EE",X"CC",X"00",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"00",
		X"00",X"88",X"CC",X"EE",X"CC",X"88",X"00",X"00",X"FF",X"FF",X"11",X"00",X"11",X"FF",X"FF",X"00",
		X"EE",X"EE",X"CC",X"88",X"CC",X"EE",X"EE",X"00",X"FF",X"FF",X"11",X"33",X"11",X"FF",X"FF",X"00",
		X"66",X"EE",X"CC",X"88",X"CC",X"EE",X"66",X"00",X"CC",X"EE",X"77",X"33",X"77",X"EE",X"CC",X"00",
		X"00",X"00",X"EE",X"EE",X"00",X"00",X"00",X"00",X"EE",X"FF",X"11",X"11",X"FF",X"EE",X"00",X"00",
		X"22",X"22",X"22",X"AA",X"EE",X"EE",X"66",X"00",X"CC",X"EE",X"FF",X"BB",X"99",X"88",X"88",X"00",
		X"00",X"ED",X"98",X"1A",X"C0",X"50",X"09",X"48",X"50",X"11",X"49",X"50",X"01",X"27",X"00",X"1E",
		X"00",X"ED",X"98",X"1A",X"C0",X"50",X"09",X"D8",X"67",X"11",X"D9",X"67",X"01",X"27",X"00",X"1E",
		X"00",X"ED",X"98",X"1A",X"C0",X"50",X"09",X"40",X"50",X"11",X"41",X"50",X"01",X"37",X"00",X"1E",
		X"00",X"ED",X"98",X"09",X"24",X"64",X"11",X"25",X"64",X"01",X"67",X"00",X"1E",X"FF",X"ED",X"98",
		X"3C",X"DE",X"EF",X"6F",X"6F",X"EF",X"DE",X"3C",X"C3",X"B7",X"7F",X"6F",X"6F",X"7F",X"B7",X"C3",
		X"3C",X"DE",X"2F",X"2F",X"2F",X"2F",X"DE",X"3C",X"C3",X"B7",X"4F",X"4F",X"4F",X"4F",X"B7",X"C3",
		X"3C",X"1E",X"0F",X"0F",X"0F",X"0F",X"1E",X"3C",X"C3",X"87",X"0F",X"0F",X"0F",X"0F",X"87",X"C3",
		X"F0",X"F8",X"FC",X"7F",X"7F",X"FC",X"F8",X"F0",X"F1",X"F3",X"E7",X"CF",X"CF",X"E7",X"F3",X"F1",
		X"F0",X"F0",X"F0",X"FF",X"FF",X"F0",X"F0",X"F0",X"F1",X"F1",X"F1",X"FF",X"FF",X"F1",X"F1",X"F1",
		X"F0",X"F0",X"F0",X"2D",X"2D",X"F0",X"F0",X"F0",X"F0",X"96",X"69",X"78",X"78",X"78",X"B4",X"F0",
		X"00",X"04",X"01",X"0A",X"00",X"04",X"01",X"00",X"00",X"02",X"08",X"00",X"02",X"09",X"04",X"01",
		X"F0",X"F0",X"F0",X"78",X"78",X"F0",X"F0",X"78",X"C3",X"E1",X"E1",X"C3",X"C3",X"E1",X"E1",X"E1",
		X"B4",X"D2",X"B4",X"78",X"78",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E1",X"E1",X"D2",X"B4",X"D2",
		X"F0",X"F0",X"F0",X"78",X"78",X"A5",X"D2",X"F0",X"F0",X"B4",X"5A",X"E1",X"E1",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"78",X"78",X"F0",X"F0",X"F0",X"F0",X"F0",X"E1",X"D2",X"D2",X"E1",X"F0",X"F0",
		X"F0",X"F0",X"78",X"B4",X"B4",X"78",X"F0",X"F0",X"F0",X"E1",X"D2",X"B4",X"B4",X"D2",X"E1",X"F0",
		X"F0",X"78",X"B4",X"D2",X"D2",X"B4",X"78",X"F0",X"E1",X"D2",X"B4",X"78",X"78",X"B4",X"D2",X"E1",
		X"B4",X"B4",X"C3",X"F0",X"F0",X"C3",X"B4",X"B4",X"D2",X"D2",X"3C",X"F0",X"F0",X"3C",X"D2",X"D2",
		X"78",X"78",X"B4",X"C3",X"C3",X"B4",X"78",X"78",X"E1",X"E1",X"D2",X"3C",X"3C",X"D2",X"E1",X"E1",
		X"78",X"78",X"78",X"87",X"87",X"78",X"78",X"78",X"E1",X"E1",X"E1",X"1E",X"1E",X"E1",X"E1",X"E1",
		X"F0",X"F0",X"78",X"3C",X"3C",X"78",X"F0",X"F0",X"1E",X"87",X"C3",X"E1",X"E1",X"C3",X"87",X"1E",
		X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",
		X"87",X"1E",X"3C",X"78",X"78",X"3C",X"1E",X"87",X"F0",X"F0",X"E1",X"C3",X"C3",X"E1",X"F0",X"F0",
		X"3C",X"D2",X"E1",X"E1",X"E1",X"E1",X"D2",X"3C",X"C3",X"B4",X"78",X"78",X"78",X"78",X"B4",X"C3",
		X"F0",X"F0",X"1E",X"E1",X"E1",X"1E",X"F0",X"F0",X"F0",X"F0",X"87",X"78",X"78",X"87",X"F0",X"F0",
		X"F0",X"F0",X"C3",X"2D",X"2D",X"C3",X"F0",X"F0",X"F0",X"F0",X"3C",X"4B",X"4B",X"3C",X"F0",X"F0",
		X"F0",X"78",X"B4",X"3C",X"3C",X"B4",X"78",X"F0",X"F0",X"E1",X"D2",X"C3",X"C3",X"D2",X"E1",X"F0",
		X"F0",X"B4",X"D2",X"5A",X"5A",X"D2",X"B4",X"F0",X"F0",X"D2",X"B4",X"A5",X"A5",X"B4",X"D2",X"F0",
		X"96",X"E1",X"E1",X"69",X"69",X"E1",X"E1",X"96",X"96",X"78",X"78",X"69",X"69",X"78",X"78",X"96",
		X"78",X"78",X"D2",X"E1",X"E1",X"D2",X"78",X"78",X"E1",X"E1",X"B4",X"78",X"78",X"B4",X"E1",X"E1",
		X"96",X"69",X"69",X"F0",X"F0",X"78",X"78",X"F0",X"F0",X"E1",X"E1",X"F0",X"F0",X"69",X"69",X"96",
		X"F0",X"F0",X"78",X"78",X"78",X"69",X"E1",X"96",X"96",X"78",X"69",X"E1",X"E1",X"E1",X"F0",X"F0",
		X"F0",X"F0",X"1E",X"E1",X"E1",X"1E",X"F0",X"F0",X"F0",X"F0",X"87",X"78",X"78",X"87",X"F0",X"F0",
		X"F0",X"1E",X"E1",X"E1",X"E1",X"E1",X"1E",X"F0",X"F0",X"87",X"78",X"78",X"78",X"78",X"87",X"F0",
		X"1E",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"1E",X"87",X"78",X"78",X"78",X"78",X"78",X"78",X"87",
		X"F0",X"F0",X"78",X"3C",X"3C",X"78",X"F0",X"F0",X"F0",X"F0",X"E1",X"C3",X"C3",X"E1",X"F0",X"F0",
		X"F0",X"78",X"3C",X"1E",X"1E",X"3C",X"78",X"F0",X"F0",X"E1",X"C3",X"87",X"87",X"C3",X"E1",X"F0",
		X"78",X"3C",X"1E",X"0F",X"0F",X"1E",X"3C",X"78",X"E1",X"C3",X"87",X"0F",X"0F",X"87",X"C3",X"E1",
		X"96",X"C3",X"E1",X"F0",X"F0",X"E1",X"C3",X"96",X"96",X"3C",X"78",X"F0",X"F0",X"78",X"3C",X"96",
		X"1E",X"87",X"C3",X"E1",X"E1",X"C3",X"87",X"1E",X"87",X"1E",X"3C",X"78",X"78",X"3C",X"1E",X"87",
		X"3C",X"0F",X"87",X"C3",X"C3",X"87",X"0F",X"3C",X"87",X"0F",X"1E",X"3C",X"3C",X"1E",X"0F",X"87",
		X"C3",X"E1",X"B4",X"F0",X"F0",X"B4",X"E1",X"C3",X"3C",X"78",X"D2",X"F0",X"F0",X"D2",X"78",X"3C",
		X"F0",X"96",X"D2",X"78",X"78",X"D2",X"96",X"F0",X"F0",X"96",X"B4",X"E1",X"E1",X"B4",X"96",X"F0",
		X"F0",X"F0",X"3C",X"3C",X"3C",X"3C",X"F0",X"F0",X"F0",X"F0",X"C3",X"C3",X"C3",X"C3",X"F0",X"F0",
		X"F0",X"F0",X"D2",X"0F",X"0F",X"D2",X"F0",X"F0",X"F0",X"F0",X"B4",X"0F",X"0F",X"B4",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"78",X"78",X"87",X"87",X"96",X"96",X"1E",X"1E",X"E1",X"E1",X"F0",X"F0",X"F0",
		X"96",X"87",X"87",X"78",X"78",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E1",X"E1",X"1E",X"1E",X"96",
		X"E0",X"D0",X"B0",X"70",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"D0",X"B0",X"70",
		X"F1",X"F3",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"F0",X"F0",X"F0",X"F1",X"F3",X"F7",X"FF",
		X"F0",X"F0",X"F0",X"F0",X"F8",X"FC",X"FE",X"FF",X"F8",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F0",X"F0",X"F0",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"F0",X"F0",X"F0",
		X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"F3",X"F1",X"FF",X"F7",X"F3",X"F1",X"F0",X"F0",X"F0",X"F0",
		X"FF",X"FE",X"FC",X"F8",X"F0",X"F0",X"F0",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"F8",
		X"FC",X"FC",X"FC",X"FC",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",
		X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"30",X"30",X"30",X"30",X"FC",X"FC",X"FC",X"FC",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",
		X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"30",X"30",X"30",X"30",
		X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"FC",X"FC",X"FC",X"FC",X"30",X"30",X"30",X"30",
		X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",
		X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"30",X"30",X"30",X"30",X"FC",X"FC",X"FC",X"FC",X"30",X"30",X"30",X"30",X"FC",X"FC",X"FC",X"FC",
		X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"30",X"30",X"30",X"30",X"FC",X"FC",X"FC",X"FC",
		X"FC",X"FC",X"FC",X"FC",X"30",X"30",X"30",X"30",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"FC",X"FC",X"FC",X"FC",
		X"FC",X"FC",X"FC",X"FC",X"30",X"30",X"30",X"30",X"FC",X"FC",X"FC",X"FC",X"30",X"30",X"30",X"30",
		X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"06",X"06",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"06",X"06",X"00",X"00",X"00",X"00",X"06",X"06",X"00",X"00",X"00",X"00",
		X"00",X"00",X"06",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"00",X"00",
		X"06",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"06",
		X"00",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"00",
		X"00",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"00",X"00",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"0C",X"00",X"00",X"03",X"03",X"00",X"00",X"00",X"00",X"00",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"C0",X"E0",X"F4",X"F8",X"F8",X"F4",X"E0",X"C0",X"30",X"70",X"F2",X"F1",X"F1",X"F2",X"70",X"30",
		X"47",X"4F",X"52",X"4B",X"41",X"4E",X"53",X"2C",X"43",X"4F",X"50",X"59",X"52",X"49",X"47",X"48",
		X"54",X"20",X"31",X"39",X"38",X"33",X"54",X"45",X"43",X"48",X"53",X"54",X"41",X"52",X"20",X"49",
		X"4E",X"43",X"1A",X"04",X"65",X"E5",X"AC",X"38",X"E5",X"E1",X"38",X"09",X"97",X"64",X"E3",X"E6",
		X"09",X"96",X"64",X"E3",X"4E",X"28",X"02",X"30",X"32",X"3E",X"00",X"1A",X"03",X"50",X"E5",X"66",
		X"15",X"11",X"50",X"41",X"09",X"DD",X"30",X"3E",X"01",X"06",X"25",X"E5",X"F7",X"15",X"3E",X"03",
		X"E5",X"71",X"15",X"09",X"96",X"64",X"E3",X"EE",X"3A",X"8E",X"64",X"3D",X"1A",X"8E",X"64",X"3E",
		X"40",X"09",X"16",X"40",X"11",X"17",X"40",X"01",X"20",X"00",X"5F",X"ED",X"98",X"E5",X"13",X"00",
		X"3A",X"FF",X"64",X"1A",X"03",X"65",X"3A",X"00",X"65",X"1A",X"04",X"65",X"E5",X"21",X"39",X"C3",
		X"B2",X"23",X"09",X"96",X"64",X"E3",X"4E",X"08",X"E2",X"E3",X"6E",X"28",X"AC",X"3A",X"96",X"64",
		X"E3",X"7F",X"08",X"43",X"E5",X"66",X"15",X"11",X"50",X"41",X"09",X"02",X"31",X"3E",X"01",X"06",
		X"25",X"E5",X"F7",X"15",X"3E",X"03",X"E5",X"71",X"15",X"09",X"96",X"64",X"E3",X"AE",X"3A",X"8F",
		X"64",X"3D",X"1A",X"8F",X"64",X"3E",X"40",X"09",X"02",X"40",X"11",X"03",X"40",X"01",X"20",X"00",
		X"5F",X"ED",X"98",X"E5",X"0C",X"00",X"3A",X"01",X"65",X"1A",X"03",X"65",X"3A",X"02",X"65",X"1A",
		X"04",X"65",X"E5",X"11",X"39",X"30",X"1B",X"3E",X"01",X"1A",X"03",X"50",X"30",X"9E",X"E5",X"66",
		X"15",X"09",X"96",X"64",X"E3",X"4E",X"C2",X"E8",X"22",X"11",X"10",X"41",X"09",X"27",X"31",X"3E",
		X"01",X"06",X"11",X"E5",X"F7",X"15",X"09",X"08",X"65",X"E3",X"C6",X"3E",X"01",X"E5",X"71",X"15",
		X"09",X"96",X"64",X"E3",X"6E",X"28",X"8F",X"C3",X"E8",X"22",X"E5",X"EF",X"26",X"09",X"97",X"64",
		X"E3",X"66",X"28",X"13",X"E3",X"A6",X"09",X"C2",X"65",X"E3",X"C6",X"1A",X"C0",X"50",X"3A",X"C2",
		X"65",X"FE",X"00",X"08",X"DE",X"30",X"05",X"3E",X"02",X"E5",X"71",X"15",X"E5",X"C5",X"33",X"ED",
		X"73",X"AE",X"64",X"7B",X"9A",X"28",X"21",X"09",X"00",X"00",X"0A",X"AE",X"64",X"E5",X"73",X"27",
		X"1A",X"C0",X"50",X"E5",X"37",X"16",X"09",X"96",X"64",X"E3",X"66",X"28",X"F7",X"E3",X"A6",X"E5",
		X"14",X"16",X"09",X"96",X"64",X"E3",X"56",X"08",X"27",X"E5",X"33",X"39",X"E5",X"14",X"16",X"09",
		X"96",X"64",X"E3",X"76",X"08",X"21",X"30",X"4F",X"E3",X"96",X"E5",X"32",X"39",X"30",X"EA",X"E3",
		X"B6",X"09",X"97",X"64",X"E3",X"E6",X"09",X"96",X"64",X"E3",X"6E",X"08",X"29",X"3A",X"01",X"65",
		X"3C",X"FE",X"24",X"08",X"02",X"3E",X"23",X"1A",X"01",X"65",X"1A",X"03",X"65",X"3A",X"02",X"65",
		X"3C",X"FE",X"31",X"08",X"02",X"3E",X"30",X"1A",X"02",X"65",X"1A",X"04",X"65",X"E5",X"34",X"39",
		X"E5",X"31",X"39",X"C3",X"B2",X"23",X"3A",X"FF",X"64",X"3C",X"FE",X"24",X"08",X"02",X"3E",X"23",
		X"1A",X"FF",X"64",X"1A",X"03",X"65",X"3A",X"00",X"65",X"3C",X"FE",X"31",X"08",X"02",X"3E",X"30",
		X"1A",X"00",X"65",X"1A",X"04",X"65",X"E5",X"34",X"39",X"E5",X"30",X"39",X"C3",X"B2",X"23",X"3A",
		X"98",X"64",X"FE",X"00",X"08",X"2E",X"09",X"96",X"64",X"E3",X"6E",X"08",X"2F",X"3A",X"8F",X"64",
		X"FE",X"00",X"08",X"66",X"E5",X"66",X"15",X"11",X"90",X"41",X"09",X"08",X"31",X"3E",X"01",X"06",
		X"21",X"E5",X"F7",X"15",X"3E",X"02",X"E5",X"71",X"15",X"E5",X"F8",X"11",X"09",X"95",X"64",X"E3",
		X"DE",X"C3",X"7D",X"07",X"D6",X"01",X"1A",X"98",X"64",X"C3",X"6E",X"23",X"3A",X"8E",X"64",X"FE",
		X"00",X"08",X"0D",X"09",X"96",X"64",X"E3",X"4E",X"08",X"E2",X"E5",X"66",X"15",X"11",X"D8",X"40",
		X"09",X"29",X"31",X"3E",X"01",X"06",X"14",X"E5",X"F7",X"15",X"3E",X"03",X"E5",X"71",X"15",X"C3",
		X"35",X"23",X"E5",X"10",X"39",X"C3",X"12",X"23",X"E5",X"20",X"39",X"C3",X"12",X"23",X"2A",X"91",
		X"64",X"EB",X"F5",X"09",X"00",X"00",X"F5",X"31",X"F5",X"7E",X"01",X"F5",X"86",X"02",X"47",X"CE",
		X"27",X"F5",X"5F",X"02",X"E3",X"38",X"E3",X"38",X"E3",X"38",X"E3",X"38",X"F5",X"7E",X"00",X"09",
		X"FC",X"24",X"E3",X"0F",X"E5",X"BA",X"15",X"76",X"0B",X"56",X"EB",X"E9",X"20",X"25",X"20",X"25",
		X"21",X"25",X"11",X"25",X"31",X"25",X"09",X"25",X"E1",X"F5",X"7E",X"04",X"90",X"F5",X"5F",X"04",
		X"E1",X"F5",X"7E",X"04",X"80",X"F5",X"5F",X"04",X"E1",X"F5",X"7E",X"03",X"80",X"F5",X"5F",X"03",
		X"E1",X"F5",X"7E",X"03",X"90",X"F5",X"5F",X"03",X"E1",X"2A",X"76",X"64",X"EB",X"F5",X"09",X"00",
		X"00",X"F5",X"31",X"EB",X"01",X"00",X"64",X"1F",X"3F",X"ED",X"42",X"CD",X"F5",X"7E",X"00",X"09",
		X"64",X"25",X"E3",X"0F",X"E5",X"BA",X"15",X"76",X"0B",X"56",X"EB",X"E9",X"34",X"26",X"70",X"25",
		X"B3",X"25",X"2B",X"26",X"1D",X"26",X"60",X"26",X"F5",X"7E",X"03",X"1A",X"74",X"64",X"F5",X"7E",
		X"04",X"1A",X"75",X"64",X"E5",X"9A",X"26",X"F5",X"7E",X"06",X"12",X"3A",X"22",X"64",X"FE",X"00",
		X"08",X"17",X"3A",X"23",X"64",X"FE",X"00",X"08",X"17",X"C1",X"09",X"24",X"64",X"21",X"CD",X"D1",
		X"13",X"01",X"05",X"00",X"1E",X"FF",X"ED",X"98",X"E1",X"F5",X"7E",X"06",X"13",X"12",X"30",X"E9",
		X"F5",X"7E",X"06",X"09",X"08",X"00",X"31",X"EB",X"12",X"30",X"F6",X"E5",X"F2",X"26",X"F5",X"7E",
		X"03",X"90",X"1A",X"74",X"64",X"F5",X"7E",X"04",X"1A",X"75",X"64",X"E5",X"9A",X"26",X"3A",X"22",
		X"64",X"FE",X"00",X"28",X"1A",X"3A",X"22",X"64",X"E3",X"0F",X"F5",X"46",X"05",X"80",X"3D",X"C1",
		X"FD",X"09",X"24",X"64",X"FD",X"21",X"FD",X"5B",X"00",X"FD",X"5A",X"01",X"FD",X"5F",X"02",X"3C",
		X"13",X"FD",X"5B",X"03",X"FD",X"5A",X"04",X"FD",X"5F",X"05",X"3A",X"74",X"64",X"F5",X"5F",X"03",
		X"3A",X"75",X"64",X"F5",X"5F",X"04",X"E1",X"3A",X"23",X"64",X"FE",X"00",X"E2",X"51",X"26",X"3A",
		X"23",X"64",X"E3",X"0F",X"C6",X"27",X"F5",X"46",X"05",X"80",X"C1",X"FD",X"09",X"24",X"64",X"FD",
		X"21",X"FD",X"5B",X"00",X"FD",X"5A",X"01",X"FD",X"5F",X"02",X"3C",X"09",X"08",X"00",X"31",X"EB",
		X"FD",X"5B",X"03",X"FD",X"5A",X"04",X"FD",X"5F",X"05",X"C3",X"F2",X"25",X"F5",X"7E",X"03",X"1A",
		X"74",X"64",X"F5",X"7E",X"04",X"1A",X"75",X"64",X"C3",X"AB",X"25",X"E5",X"F2",X"26",X"F5",X"7E",
		X"03",X"80",X"C3",X"8A",X"25",X"E5",X"F2",X"26",X"F5",X"7E",X"04",X"90",X"1A",X"75",X"64",X"F5",
		X"7E",X"03",X"1A",X"74",X"64",X"C3",X"AB",X"25",X"E5",X"F2",X"26",X"F5",X"7E",X"04",X"80",X"30",
		X"EB",X"F5",X"7E",X"05",X"C1",X"FD",X"09",X"24",X"64",X"FD",X"21",X"FD",X"5B",X"00",X"FD",X"5A",
		X"01",X"FD",X"5F",X"02",X"3A",X"74",X"64",X"F5",X"5F",X"03",X"3A",X"75",X"64",X"F5",X"5F",X"04",
		X"F5",X"7E",X"00",X"09",X"85",X"26",X"E3",X"0F",X"E5",X"BA",X"15",X"D5",X"76",X"0B",X"56",X"EB",
		X"D1",X"F5",X"7E",X"06",X"E9",X"91",X"26",X"91",X"26",X"92",X"26",X"B5",X"26",X"88",X"26",X"8F",
		X"26",X"E1",X"13",X"FD",X"5B",X"03",X"FD",X"5A",X"04",X"FD",X"5F",X"05",X"E1",X"33",X"30",X"DB",
		X"09",X"08",X"00",X"31",X"EB",X"30",X"EC",X"EB",X"11",X"08",X"00",X"1F",X"3F",X"ED",X"52",X"EB",
		X"30",X"C9",X"3A",X"74",X"64",X"CE",X"07",X"1A",X"22",X"64",X"3A",X"75",X"64",X"CE",X"07",X"1A",
		X"23",X"64",X"3A",X"74",X"64",X"E3",X"3F",X"E3",X"3F",X"E3",X"3F",X"57",X"3A",X"75",X"64",X"E3",
		X"3F",X"E3",X"3F",X"E3",X"3F",X"77",X"E5",X"E9",X"14",X"E1",X"F5",X"7E",X"01",X"F5",X"86",X"02",
		X"47",X"CE",X"27",X"F5",X"5F",X"02",X"E3",X"38",X"E3",X"38",X"E3",X"38",X"E3",X"38",X"E1",X"3A",
		X"03",X"65",X"09",X"FD",X"26",X"E3",X"0F",X"E3",X"0F",X"E5",X"BA",X"15",X"E9",X"E5",X"E2",X"29",
		X"E1",X"E5",X"0B",X"2A",X"E1",X"E5",X"7C",X"2A",X"E1",X"E5",X"D5",X"2A",X"E1",X"E5",X"2E",X"2B",
		X"E1",X"E5",X"87",X"2B",X"E1",X"E5",X"C8",X"2B",X"E1",X"E5",X"1E",X"2C",X"E1",X"E5",X"A4",X"2C",
		X"E1",X"E5",X"CD",X"2C",X"E1",X"E5",X"3E",X"2D",X"E1",X"E5",X"A2",X"2D",X"E1",X"E5",X"D6",X"2D",
		X"E1",X"E5",X"D7",X"2D",X"E1",X"E5",X"F0",X"2D",X"E1",X"E5",X"F1",X"2D",X"E1",X"D5",X"1F",X"3F",
		X"09",X"26",X"01",X"16",X"00",X"ED",X"52",X"7D",X"1F",X"3F",X"09",X"10",X"01",X"D1",X"72",X"16",
		X"00",X"ED",X"52",X"55",X"77",X"E1",X"7D",X"EE",X"03",X"6F",X"E1",X"09",X"96",X"64",X"E3",X"46",
		X"E0",X"E3",X"6E",X"28",X"43",X"09",X"A8",X"64",X"7B",X"86",X"0F",X"5F",X"0B",X"7A",X"A6",X"0F",
		X"5F",X"0B",X"3E",X"00",X"A6",X"0F",X"5F",X"38",X"02",X"30",X"1A",X"09",X"96",X"64",X"E3",X"6E",
		X"28",X"13",X"09",X"DE",X"43",X"11",X"DF",X"43",X"01",X"05",X"00",X"1E",X"40",X"ED",X"98",X"AF",
		X"1A",X"DE",X"43",X"30",X"30",X"09",X"CC",X"43",X"11",X"CD",X"43",X"01",X"05",X"00",X"1E",X"40",
		X"ED",X"98",X"AF",X"1A",X"CC",X"43",X"30",X"05",X"09",X"AB",X"64",X"30",X"BB",X"09",X"96",X"64",
		X"E3",X"6E",X"28",X"74",X"09",X"AA",X"64",X"11",X"FB",X"43",X"3A",X"99",X"64",X"DD",X"E5",X"33",
		X"10",X"0B",X"0B",X"0B",X"EB",X"2A",X"8B",X"64",X"D9",X"FE",X"04",X"D0",X"E3",X"0F",X"E3",X"0F",
		X"3C",X"3C",X"E5",X"BA",X"15",X"E5",X"98",X"11",X"D0",X"3A",X"98",X"64",X"3C",X"1A",X"98",X"64",
		X"09",X"08",X"65",X"E3",X"C6",X"09",X"96",X"64",X"E3",X"6E",X"28",X"12",X"3A",X"99",X"64",X"3C",
		X"1A",X"99",X"64",X"3A",X"8E",X"64",X"3C",X"1A",X"8E",X"64",X"E5",X"13",X"00",X"E1",X"3A",X"9A",
		X"9C",X"63",X"41",X"9C",X"BE",X"BE",X"41",X"00",X"41",X"14",X"36",X"41",X"63",X"63",X"14",X"00",
		X"41",X"41",X"FF",X"00",X"41",X"41",X"FF",X"00",X"00",X"22",X"77",X"00",X"00",X"00",X"77",X"00",
		X"41",X"FF",X"DD",X"63",X"C9",X"77",X"DD",X"00",X"63",X"14",X"55",X"22",X"77",X"36",X"14",X"00",
		X"36",X"C9",X"C9",X"22",X"FF",X"63",X"C9",X"00",X"14",X"14",X"77",X"00",X"36",X"14",X"55",X"00",
		X"00",X"00",X"88",X"CC",X"66",X"22",X"33",X"FF",X"00",X"00",X"11",X"33",X"66",X"00",X"00",X"77",
		X"33",X"EE",X"88",X"00",X"00",X"00",X"00",X"FF",X"CC",X"77",X"11",X"00",X"00",X"00",X"00",X"FF",
		X"EE",X"00",X"00",X"66",X"CC",X"88",X"00",X"00",X"FF",X"CC",X"44",X"66",X"33",X"11",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"88",X"EE",X"33",X"FF",X"00",X"00",X"00",X"00",X"11",X"77",X"CC",
		X"00",X"00",X"00",X"88",X"88",X"CC",X"44",X"44",X"00",X"00",X"33",X"77",X"55",X"44",X"44",X"66",
		X"00",X"33",X"11",X"88",X"CC",X"EE",X"77",X"33",X"00",X"00",X"EE",X"33",X"00",X"00",X"00",X"88",
		X"66",X"22",X"22",X"AA",X"EE",X"CC",X"00",X"00",X"22",X"22",X"33",X"11",X"11",X"00",X"00",X"00",
		X"11",X"00",X"00",X"00",X"CC",X"77",X"00",X"00",X"CC",X"EE",X"77",X"33",X"11",X"77",X"CC",X"00",
		X"00",X"00",X"00",X"88",X"88",X"CC",X"44",X"66",X"00",X"00",X"00",X"11",X"11",X"33",X"22",X"66",
		X"77",X"DD",X"99",X"99",X"11",X"11",X"11",X"11",X"00",X"99",X"99",X"99",X"88",X"88",X"88",X"88",
		X"66",X"44",X"CC",X"88",X"88",X"00",X"00",X"00",X"66",X"22",X"33",X"11",X"11",X"00",X"00",X"00",
		X"11",X"11",X"11",X"11",X"99",X"99",X"99",X"44",X"88",X"88",X"88",X"88",X"99",X"99",X"BB",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"88",X"CC",X"CC",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"11",
		X"00",X"00",X"33",X"66",X"EE",X"00",X"00",X"FF",X"00",X"00",X"CC",X"66",X"77",X"11",X"00",X"FF",
		X"88",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"33",X"33",X"11",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"88",X"EE",X"66",X"33",X"00",X"00",X"FF",X"00",X"00",X"77",X"66",X"CC",X"00",X"00",
		X"00",X"00",X"00",X"00",X"88",X"88",X"44",X"44",X"00",X"00",X"00",X"00",X"00",X"11",X"22",X"22",
		X"00",X"00",X"33",X"00",X"88",X"44",X"22",X"11",X"00",X"00",X"CC",X"33",X"00",X"00",X"00",X"00",
		X"44",X"44",X"88",X"00",X"00",X"00",X"00",X"00",X"22",X"22",X"11",X"11",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"CC",X"33",X"00",X"00",X"88",X"44",X"22",X"11",X"00",X"CC",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"88",X"CC",X"44",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"22",
		X"00",X"00",X"33",X"FF",X"DD",X"99",X"11",X"11",X"00",X"00",X"00",X"33",X"99",X"99",X"88",X"88",
		X"44",X"CC",X"88",X"00",X"00",X"00",X"00",X"00",X"22",X"33",X"11",X"00",X"00",X"00",X"00",X"00",
		X"11",X"11",X"99",X"99",X"DD",X"00",X"00",X"00",X"88",X"88",X"99",X"BB",X"FF",X"CC",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",
		X"00",X"00",X"00",X"33",X"66",X"CC",X"00",X"FF",X"00",X"00",X"00",X"CC",X"66",X"33",X"11",X"FF",
		X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"88",X"CC",X"66",X"33",X"00",X"00",X"00",X"FF",X"00",X"33",X"66",X"CC",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"99",X"CC",X"AA",X"99",X"00",X"00",X"00",X"00",X"CC",X"66",X"33",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"CC",X"66",X"33",X"00",X"00",X"00",X"00",X"99",X"55",X"33",X"88",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",
		X"00",X"00",X"00",X"33",X"77",X"DD",X"99",X"11",X"00",X"00",X"00",X"22",X"AA",X"BB",X"99",X"88",
		X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"99",X"DD",X"55",X"44",X"00",X"00",X"00",X"88",X"99",X"BB",X"AA",X"CC",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"33",X"EE",X"00",X"77",X"00",X"00",X"00",X"00",X"CC",X"66",X"33",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"CC",X"66",X"33",X"00",X"00",X"00",X"00",X"EE",X"00",X"77",X"CC",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"11",X"44",X"AA",X"99",X"00",X"00",X"00",X"00",X"CC",X"22",X"11",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"88",X"44",X"33",X"00",X"00",X"00",X"00",X"99",X"55",X"22",X"88",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"33",X"55",X"55",X"99",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"99",X"AA",X"AA",X"CC",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"33",X"00",X"00",X"00",X"00",X"00",X"CC",X"22",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"44",X"33",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"11",X"44",X"66",X"55",X"00",X"00",X"00",X"00",X"00",X"88",X"44",X"22",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"22",X"11",X"00",X"00",X"00",X"00",X"00",X"AA",X"66",X"22",X"88",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"77",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"EE",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"88",X"CC",X"EE",X"EE",X"FF",X"FF",X"00",X"00",X"11",X"33",X"77",X"77",X"FF",X"FF",
		X"33",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"EE",X"EE",X"CC",X"88",X"00",X"00",X"FF",X"FF",X"77",X"77",X"33",X"11",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"33",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CC",
		X"00",X"00",X"88",X"88",X"88",X"CC",X"CC",X"CC",X"00",X"00",X"11",X"11",X"11",X"33",X"33",X"33",
		X"FB",X"F8",X"FB",X"FF",X"FC",X"FB",X"FC",X"FF",X"FB",X"F1",X"FF",X"FF",X"F3",X"FD",X"F3",X"FF",
		X"CC",X"CC",X"88",X"88",X"88",X"00",X"00",X"00",X"33",X"33",X"11",X"11",X"11",X"00",X"00",X"00",
		X"FC",X"FB",X"FC",X"FF",X"FC",X"FB",X"FC",X"00",X"F3",X"FD",X"F3",X"FF",X"F3",X"FD",X"F3",X"00",
		X"00",X"00",X"88",X"88",X"88",X"CC",X"CC",X"CC",X"00",X"00",X"11",X"11",X"11",X"33",X"33",X"33",
		X"F9",X"FA",X"FB",X"FB",X"FF",X"FC",X"FB",X"FC",X"FB",X"FD",X"F5",X"FB",X"FF",X"F3",X"FD",X"F3",
		X"CC",X"CC",X"CC",X"88",X"88",X"88",X"00",X"00",X"33",X"33",X"33",X"11",X"11",X"11",X"00",X"00",
		X"FF",X"FC",X"FB",X"FC",X"FF",X"FC",X"FB",X"FC",X"FF",X"F3",X"FD",X"F3",X"FF",X"F3",X"FD",X"F3",
		X"00",X"00",X"88",X"88",X"88",X"CC",X"CC",X"CC",X"00",X"00",X"11",X"11",X"11",X"33",X"33",X"33",
		X"FF",X"FE",X"FE",X"F8",X"FE",X"FC",X"FB",X"FC",X"FF",X"F7",X"FB",X"F1",X"FF",X"F3",X"FD",X"F3",
		X"CC",X"CC",X"CC",X"88",X"88",X"88",X"00",X"00",X"33",X"33",X"33",X"11",X"11",X"11",X"00",X"00",
		X"FF",X"FC",X"FB",X"FC",X"FF",X"FC",X"FB",X"FC",X"FF",X"F3",X"FD",X"F3",X"FF",X"F3",X"FD",X"F3",
		X"00",X"00",X"88",X"88",X"88",X"CC",X"CC",X"CC",X"00",X"00",X"11",X"11",X"11",X"33",X"33",X"33",
		X"FC",X"FB",X"FB",X"FC",X"FF",X"FC",X"FB",X"FC",X"FB",X"F5",X"F5",X"FB",X"FF",X"F3",X"FD",X"F3",
		X"CC",X"CC",X"CC",X"88",X"88",X"88",X"00",X"00",X"33",X"33",X"33",X"11",X"11",X"11",X"00",X"00",
		X"FF",X"FC",X"FB",X"FC",X"FF",X"FC",X"FB",X"FC",X"FF",X"F3",X"FD",X"F3",X"FF",X"F3",X"FD",X"F3",
		X"00",X"00",X"00",X"00",X"88",X"CC",X"EE",X"FF",X"00",X"00",X"00",X"00",X"32",X"76",X"EF",X"CF",
		X"00",X"00",X"02",X"70",X"67",X"91",X"08",X"0C",X"00",X"00",X"22",X"33",X"19",X"0C",X"37",X"37",
		X"FF",X"EE",X"CC",X"88",X"00",X"00",X"00",X"00",X"8F",X"EF",X"76",X"32",X"00",X"00",X"00",X"00",
		X"0C",X"08",X"91",X"E7",X"70",X"02",X"00",X"00",X"37",X"37",X"0C",X"19",X"33",X"22",X"00",X"00",
		X"00",X"00",X"00",X"00",X"88",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"00",X"00",
		X"11",X"33",X"77",X"FF",X"BB",X"33",X"07",X"0C",X"88",X"CC",X"EE",X"FF",X"DD",X"CC",X"0E",X"03",
		X"80",X"84",X"80",X"00",X"00",X"00",X"00",X"00",X"10",X"12",X"10",X"00",X"00",X"00",X"00",X"00",
		X"4C",X"88",X"89",X"C3",X"C3",X"EF",X"77",X"33",X"23",X"11",X"19",X"3C",X"3C",X"7F",X"EE",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"EE",X"00",X"00",X"11",X"33",X"76",X"BA",X"AB",X"CF",
		X"00",X"00",X"8A",X"70",X"E7",X"91",X"08",X"0C",X"00",X"00",X"00",X"00",X"08",X"2E",X"37",X"37",
		X"EE",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"CF",X"AB",X"BA",X"76",X"33",X"11",X"00",X"00",
		X"0C",X"08",X"91",X"E7",X"70",X"8A",X"00",X"00",X"37",X"37",X"2E",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"11",X"33",X"33",X"77",X"07",X"0C",X"00",X"88",X"88",X"CC",X"CC",X"EE",X"0E",X"03",
		X"80",X"84",X"80",X"44",X"CC",X"88",X"00",X"00",X"10",X"12",X"10",X"22",X"33",X"11",X"00",X"00",
		X"4C",X"88",X"89",X"C3",X"C3",X"EF",X"99",X"77",X"23",X"11",X"19",X"3C",X"3C",X"7F",X"99",X"EE",
		X"47",X"4F",X"52",X"4B",X"41",X"4E",X"53",X"2C",X"43",X"4F",X"50",X"59",X"52",X"49",X"47",X"48",
		X"54",X"20",X"31",X"39",X"38",X"33",X"54",X"45",X"43",X"48",X"53",X"54",X"41",X"52",X"20",X"49",
		X"4E",X"43",X"F0",X"F0",X"F0",X"F0",X"78",X"78",X"93",X"93",X"B1",X"B1",X"B1",X"B1",X"93",X"B1",
		X"E4",X"78",X"E4",X"F0",X"D2",X"F0",X"78",X"F0",X"F0",X"B1",X"F0",X"E4",X"F0",X"D2",X"B1",X"D2",
		X"F0",X"78",X"F0",X"D2",X"F0",X"A5",X"78",X"F0",X"F0",X"B1",X"5A",X"F0",X"E4",X"F0",X"B1",X"F0",
		X"F0",X"78",X"F0",X"F0",X"F0",X"F0",X"78",X"F0",X"F0",X"D2",X"B1",X"F0",X"F0",X"B1",X"D2",X"F0",
		X"F0",X"E4",X"78",X"F0",X"F0",X"78",X"E4",X"F0",X"F0",X"E4",X"D2",X"B1",X"B1",X"D2",X"E4",X"F0",
		X"F0",X"D2",X"E4",X"78",X"78",X"E4",X"D2",X"F0",X"B1",X"78",X"E4",X"D2",X"D2",X"E4",X"78",X"B1",
		X"E4",X"F0",X"93",X"E4",X"E4",X"93",X"F0",X"E4",X"D2",X"F0",X"6C",X"D2",X"D2",X"6C",X"F0",X"D2",
		X"78",X"93",X"E4",X"78",X"78",X"E4",X"93",X"78",X"B1",X"6C",X"D2",X"B1",X"B1",X"D2",X"6C",X"B1",
		X"78",X"87",X"78",X"78",X"78",X"78",X"87",X"78",X"B1",X"4E",X"B1",X"B1",X"B1",X"B1",X"4E",X"B1",
		X"F0",X"6C",X"78",X"F0",X"F0",X"78",X"6C",X"F0",X"4E",X"B1",X"93",X"87",X"87",X"93",X"B1",X"4E",
		X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"B1",X"B1",X"B1",X"B1",X"B1",X"B1",X"B1",X"B1",
		X"87",X"78",X"6C",X"4E",X"4E",X"6C",X"78",X"87",X"F0",X"93",X"B1",X"F0",X"F0",X"B1",X"93",X"F0",
		X"6C",X"B1",X"B1",X"D2",X"D2",X"B1",X"B1",X"6C",X"93",X"78",X"78",X"E4",X"E4",X"78",X"78",X"93",
		X"F0",X"B1",X"4E",X"F0",X"F0",X"4E",X"B1",X"F0",X"F0",X"78",X"87",X"F0",X"F0",X"87",X"78",X"F0",
		X"F0",X"2D",X"93",X"F0",X"F0",X"93",X"2D",X"F0",X"F0",X"1B",X"6C",X"F0",X"F0",X"6C",X"1B",X"F0",
		X"F0",X"6C",X"E4",X"78",X"78",X"E4",X"6C",X"F0",X"F0",X"93",X"D2",X"B1",X"B1",X"D2",X"93",X"F0",
		X"F0",X"5A",X"D2",X"E4",X"E4",X"D2",X"5A",X"F0",X"F0",X"A5",X"E4",X"D2",X"D2",X"E4",X"A5",X"F0",
		X"C6",X"39",X"B1",X"B1",X"B1",X"B1",X"39",X"C6",X"C6",X"39",X"78",X"78",X"78",X"78",X"39",X"C6",
		X"78",X"B1",X"D2",X"78",X"78",X"D2",X"B1",X"78",X"B1",X"78",X"E4",X"B1",X"B1",X"E4",X"78",X"B1",
		X"C6",X"F0",X"39",X"78",X"39",X"78",X"F0",X"F0",X"F0",X"F0",X"B1",X"39",X"B1",X"39",X"F0",X"C6",
		X"F0",X"78",X"78",X"B1",X"F0",X"39",X"78",X"C6",X"C6",X"B1",X"39",X"F0",X"78",X"B1",X"B1",X"F0",
		X"F0",X"B1",X"4E",X"F0",X"F0",X"4E",X"B1",X"F0",X"F0",X"78",X"87",X"F0",X"F0",X"87",X"78",X"F0",
		X"F0",X"B1",X"B1",X"4E",X"4E",X"B1",X"B1",X"F0",X"F0",X"78",X"78",X"87",X"87",X"78",X"78",X"F0",
		X"4E",X"B1",X"B1",X"B1",X"B1",X"B1",X"B1",X"4E",X"87",X"78",X"78",X"78",X"78",X"78",X"78",X"87",
		X"F0",X"6C",X"78",X"F0",X"F0",X"78",X"6C",X"F0",X"F0",X"93",X"B1",X"F0",X"F0",X"B1",X"93",X"F0",
		X"F0",X"4E",X"6C",X"78",X"78",X"6C",X"4E",X"F0",X"F0",X"87",X"93",X"B1",X"B1",X"93",X"87",X"F0",
		X"78",X"0F",X"4E",X"6C",X"6C",X"4E",X"0F",X"78",X"B1",X"0F",X"87",X"93",X"93",X"87",X"0F",X"B1",
		X"C6",X"F0",X"B1",X"93",X"93",X"B1",X"F0",X"C6",X"C6",X"F0",X"78",X"6C",X"6C",X"78",X"F0",X"C6",
		X"4E",X"B1",X"93",X"87",X"87",X"93",X"B1",X"4E",X"87",X"78",X"6C",X"4E",X"4E",X"6C",X"78",X"87",
		X"6C",X"93",X"87",X"0F",X"0F",X"87",X"93",X"6C",X"87",X"6C",X"4E",X"0F",X"0F",X"4E",X"6C",X"87",
		X"93",X"F0",X"E4",X"B1",X"B1",X"E4",X"F0",X"93",X"6C",X"F0",X"D2",X"78",X"78",X"D2",X"F0",X"6C",
		X"F0",X"78",X"D2",X"C6",X"C6",X"D2",X"78",X"F0",X"F0",X"B1",X"E4",X"C6",X"C6",X"E4",X"B1",X"F0",
		X"F0",X"6C",X"6C",X"F0",X"F0",X"6C",X"6C",X"F0",X"F0",X"93",X"93",X"F0",X"F0",X"93",X"93",X"F0",
		X"F0",X"0F",X"D2",X"F0",X"F0",X"D2",X"0F",X"F0",X"F0",X"0F",X"E4",X"F0",X"F0",X"E4",X"0F",X"F0",
		X"F0",X"78",X"F0",X"87",X"F0",X"87",X"78",X"C6",X"C6",X"B1",X"4E",X"F0",X"4E",X"F0",X"B1",X"F0",
		X"C6",X"78",X"87",X"F0",X"87",X"F0",X"78",X"F0",X"F0",X"B1",X"F0",X"4E",X"F0",X"4E",X"B1",X"C6",
		X"B0",X"F0",X"E0",X"F0",X"D0",X"F0",X"70",X"F0",X"F0",X"B0",X"F0",X"E0",X"F0",X"D0",X"F0",X"70",
		X"F1",X"FF",X"F7",X"FF",X"F3",X"FF",X"FF",X"FF",X"F0",X"F1",X"F0",X"F7",X"F0",X"F3",X"F0",X"FF",
		X"F0",X"F8",X"F0",X"FE",X"F0",X"FC",X"F0",X"FF",X"F8",X"FF",X"FE",X"FF",X"FC",X"FF",X"FF",X"FF",
		X"F0",X"00",X"F0",X"F0",X"F0",X"F0",X"00",X"F0",X"F0",X"00",X"F0",X"F0",X"F0",X"F0",X"00",X"F0",
		X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"B0",X"B0",X"B0",X"B0",X"B0",X"B0",X"B0",X"B0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"F3",X"FF",X"F7",X"FF",X"F1",X"FF",X"F0",X"F3",X"F0",X"F7",X"F0",X"F1",X"F0",
		X"FF",X"F0",X"FC",X"F0",X"FE",X"F0",X"F8",X"F0",X"FF",X"FF",X"FF",X"FC",X"FF",X"FE",X"FF",X"F8",
		X"FC",X"60",X"FC",X"60",X"FC",X"60",X"FC",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",
		X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"60",X"FC",X"60",X"FC",X"60",X"FC",X"60",X"FC",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",
		X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"60",X"FC",X"60",X"FC",X"60",X"FC",X"60",
		X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"FC",X"60",X"FC",X"60",X"FC",X"60",X"FC",X"60",
		X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",
		X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"60",X"FC",X"60",X"FC",X"60",X"FC",X"60",X"FC",X"60",X"FC",X"60",X"FC",X"60",X"FC",X"60",X"FC",
		X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"60",X"FC",X"60",X"FC",X"60",X"FC",X"60",X"FC",
		X"FC",X"60",X"FC",X"60",X"FC",X"60",X"FC",X"60",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"FC",X"60",X"FC",X"60",X"FC",X"60",X"FC",
		X"FC",X"60",X"FC",X"60",X"FC",X"60",X"FC",X"60",X"FC",X"60",X"FC",X"60",X"FC",X"60",X"FC",X"60",
		X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",
		X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"06",X"06",X"00",X"00",X"00",X"06",X"00",X"00",X"00",
		X"00",X"06",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"06",X"00",
		X"00",X"00",X"06",X"00",X"00",X"00",X"06",X"00",X"00",X"06",X"00",X"00",X"00",X"06",X"00",X"00",
		X"06",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"06",
		X"00",X"00",X"0C",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"03",X"00",X"00",
		X"00",X"00",X"03",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"0C",X"00",X"00",
		X"00",X"00",X"00",X"03",X"00",X"03",X"00",X"00",X"00",X"00",X"0C",X"00",X"0C",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0C",X"00",X"0C",X"00",X"00",X"00",X"00",X"03",X"00",X"03",X"00",X"00",X"00",
		X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"90",X"F8",X"F4",X"B0",X"B0",X"F4",X"F8",X"90",X"60",X"F1",X"F2",X"70",X"70",X"F2",X"F1",X"60",
		X"17",X"11",X"52",X"53",X"1F",X"1E",X"1B",X"2C",X"13",X"52",X"50",X"17",X"1F",X"19",X"59",X"18",
		X"54",X"68",X"61",X"54",X"20",X"63",X"69",X"15",X"13",X"11",X"53",X"20",X"18",X"52",X"54",X"19",
		X"1E",X"35",X"4A",X"AC",X"13",X"B5",X"04",X"68",X"B5",X"C7",X"68",X"B3",X"B1",X"34",X"09",X"B6",
		X"09",X"1E",X"34",X"02",X"C6",X"28",X"B3",X"60",X"62",X"03",X"00",X"B5",X"6E",X"50",X"4A",X"36",
		X"45",X"09",X"50",X"60",X"41",X"DD",X"11",X"6E",X"01",X"F7",X"25",X"6E",X"06",X"45",X"B5",X"03",
		X"B5",X"C6",X"45",X"B3",X"71",X"34",X"09",X"BE",X"6A",X"4A",X"34",X"34",X"8E",X"8E",X"6D",X"6E",
		X"10",X"41",X"46",X"10",X"09",X"47",X"10",X"01",X"20",X"C8",X"5F",X"43",X"00",X"B5",X"BD",X"00",
		X"6A",X"03",X"34",X"6A",X"FF",X"35",X"4A",X"00",X"35",X"B5",X"04",X"69",X"4A",X"21",X"35",X"93",
		X"E2",X"34",X"09",X"1E",X"23",X"B3",X"C6",X"08",X"B2",X"AC",X"3E",X"C6",X"B3",X"6A",X"28",X"34",
		X"B3",X"B5",X"08",X"45",X"7F",X"36",X"13",X"41",X"50",X"61",X"09",X"01",X"11",X"6E",X"02",X"06",
		X"25",X"6E",X"F7",X"B5",X"B5",X"03",X"45",X"71",X"45",X"B3",X"C6",X"6A",X"09",X"AE",X"34",X"8F",
		X"34",X"34",X"4A",X"10",X"6D",X"6E",X"8F",X"09",X"02",X"10",X"41",X"20",X"10",X"01",X"03",X"00",
		X"5F",X"0C",X"C8",X"6A",X"BD",X"00",X"B5",X"01",X"35",X"6A",X"03",X"35",X"4A",X"02",X"35",X"4A",
		X"04",X"69",X"B5",X"4B",X"35",X"60",X"41",X"6E",X"01",X"60",X"03",X"B5",X"4A",X"CE",X"50",X"36",
		X"45",X"B3",X"C6",X"92",X"09",X"1E",X"34",X"B8",X"22",X"09",X"40",X"61",X"41",X"27",X"11",X"6E",
		X"01",X"F7",X"41",X"09",X"06",X"45",X"B5",X"08",X"35",X"01",X"96",X"71",X"B3",X"B5",X"6E",X"45",
		X"09",X"3E",X"34",X"8F",X"C6",X"28",X"B3",X"93",X"B8",X"26",X"B5",X"C7",X"22",X"09",X"BF",X"34",
		X"B3",X"B3",X"28",X"09",X"36",X"A6",X"43",X"92",X"35",X"90",X"96",X"6A",X"B3",X"50",X"4A",X"92",
		X"35",X"DE",X"00",X"05",X"FE",X"60",X"08",X"6E",X"02",X"B5",X"71",X"63",X"B5",X"95",X"45",X"BD",
		X"73",X"CA",X"34",X"21",X"AE",X"28",X"7B",X"09",X"00",X"34",X"0A",X"73",X"00",X"B5",X"AE",X"27",
		X"4A",X"67",X"50",X"09",X"90",X"46",X"B5",X"C6",X"34",X"F7",X"36",X"A6",X"B3",X"B3",X"28",X"B5",
		X"44",X"34",X"09",X"56",X"46",X"B3",X"C6",X"08",X"27",X"B5",X"63",X"46",X"B5",X"44",X"69",X"09",
		X"C6",X"08",X"B3",X"60",X"34",X"21",X"76",X"1F",X"B3",X"69",X"B5",X"BA",X"C6",X"60",X"62",X"B3",
		X"E6",X"B3",X"C7",X"09",X"09",X"B6",X"34",X"C6",X"34",X"29",X"3E",X"01",X"B3",X"6A",X"08",X"35",
		X"6C",X"02",X"24",X"23",X"FE",X"6E",X"08",X"4A",X"01",X"35",X"4A",X"02",X"35",X"6A",X"03",X"35",
		X"6C",X"02",X"61",X"60",X"FE",X"6E",X"08",X"4A",X"02",X"35",X"4A",X"64",X"35",X"B5",X"04",X"69",
		X"B5",X"E2",X"69",X"6A",X"61",X"23",X"93",X"FF",X"34",X"08",X"FE",X"6E",X"6C",X"02",X"24",X"23",
		X"4A",X"03",X"34",X"6A",X"FF",X"35",X"4A",X"00",X"35",X"08",X"FE",X"6E",X"6C",X"02",X"61",X"60",
		X"4A",X"04",X"35",X"B5",X"00",X"35",X"4A",X"64",X"69",X"93",X"60",X"23",X"B5",X"E2",X"69",X"6A",
		X"C8",X"08",X"FE",X"09",X"34",X"2E",X"00",X"C6",X"34",X"2F",X"3E",X"8F",X"B3",X"6A",X"08",X"34",
		X"FE",X"B5",X"08",X"45",X"00",X"36",X"36",X"41",X"C0",X"61",X"09",X"01",X"11",X"6E",X"08",X"06",
		X"21",X"6E",X"F7",X"B5",X"B5",X"02",X"45",X"71",X"45",X"09",X"F8",X"34",X"B5",X"C5",X"41",X"B3",
		X"DE",X"D6",X"7D",X"4A",X"93",X"01",X"07",X"C8",X"34",X"6A",X"3E",X"34",X"93",X"8E",X"23",X"FE",
		X"00",X"C6",X"0D",X"B3",X"08",X"34",X"09",X"1E",X"08",X"45",X"B5",X"D8",X"B2",X"41",X"36",X"10",
		X"09",X"01",X"61",X"44",X"29",X"06",X"6E",X"B5",X"F7",X"B5",X"6E",X"45",X"45",X"71",X"03",X"93",
		X"65",X"69",X"B5",X"42",X"23",X"93",X"40",X"23",X"B5",X"42",X"69",X"2A",X"20",X"23",X"93",X"C1",
		X"34",X"00",X"F5",X"F5",X"BB",X"00",X"09",X"61",X"F5",X"86",X"01",X"17",X"7E",X"02",X"F5",X"9E",
		X"27",X"B3",X"5F",X"B3",X"F5",X"68",X"02",X"68",X"B3",X"F5",X"B3",X"00",X"68",X"7E",X"68",X"09",
		X"FC",X"B5",X"B3",X"45",X"24",X"EA",X"0F",X"76",X"0B",X"20",X"BB",X"20",X"56",X"25",X"B9",X"25",
		X"21",X"61",X"41",X"09",X"25",X"25",X"25",X"25",X"B1",X"C0",X"7E",X"5F",X"F5",X"F5",X"04",X"04",
		X"B1",X"80",X"7E",X"5F",X"F5",X"F5",X"04",X"04",X"B1",X"80",X"7E",X"5F",X"F5",X"F5",X"03",X"03",
		X"B1",X"C0",X"7E",X"5F",X"F5",X"F5",X"03",X"03",X"B1",X"BB",X"76",X"09",X"2A",X"F5",X"34",X"00",
		X"00",X"01",X"61",X"34",X"F5",X"00",X"BB",X"4F",X"6F",X"F5",X"12",X"00",X"BD",X"7E",X"9D",X"09",
		X"34",X"B5",X"B3",X"45",X"25",X"EA",X"0F",X"76",X"0B",X"64",X"BB",X"70",X"56",X"26",X"B9",X"25",
		X"E3",X"4D",X"2B",X"30",X"25",X"26",X"26",X"26",X"F5",X"74",X"03",X"F5",X"7E",X"34",X"4A",X"7E",
		X"04",X"B5",X"75",X"26",X"4A",X"CA",X"34",X"F5",X"7E",X"22",X"42",X"FE",X"06",X"34",X"6A",X"00",
		X"08",X"34",X"6A",X"00",X"47",X"FE",X"23",X"08",X"47",X"34",X"09",X"9D",X"91",X"21",X"24",X"D1",
		X"43",X"4E",X"05",X"BD",X"01",X"FF",X"00",X"C8",X"B1",X"43",X"7E",X"60",X"F5",X"42",X"06",X"B9",
		X"F5",X"08",X"06",X"61",X"7E",X"00",X"09",X"BB",X"42",X"F2",X"F6",X"F5",X"60",X"26",X"B5",X"7E",
		X"03",X"34",X"4A",X"7E",X"C0",X"F5",X"74",X"04",X"4A",X"CA",X"34",X"6A",X"75",X"26",X"B5",X"22",
		X"34",X"4A",X"00",X"22",X"FE",X"6A",X"28",X"34",X"B3",X"05",X"F5",X"6D",X"0F",X"80",X"16",X"91",
		X"FD",X"FD",X"24",X"FD",X"09",X"21",X"34",X"5B",X"00",X"FD",X"5A",X"02",X"FD",X"5F",X"01",X"6C",
		X"43",X"FD",X"5B",X"04",X"FD",X"5A",X"03",X"FD",X"5F",X"34",X"6A",X"5F",X"05",X"F5",X"74",X"03",
		X"6A",X"5F",X"34",X"B1",X"75",X"04",X"F5",X"6A",X"23",X"B2",X"FE",X"26",X"34",X"51",X"00",X"6A",
		X"23",X"96",X"B3",X"F5",X"34",X"27",X"0F",X"16",X"05",X"09",X"91",X"34",X"80",X"24",X"FD",X"FD",
		X"21",X"FD",X"5B",X"01",X"FD",X"5A",X"00",X"FD",X"5F",X"08",X"6C",X"61",X"02",X"00",X"09",X"BB",
		X"FD",X"5A",X"03",X"FD",X"5B",X"04",X"FD",X"5F",X"05",X"F5",X"F2",X"03",X"93",X"7E",X"25",X"4A",
		X"74",X"04",X"F5",X"75",X"34",X"4A",X"7E",X"34",X"93",X"F2",X"25",X"F5",X"AB",X"26",X"B5",X"7E",
		X"03",X"25",X"93",X"F2",X"80",X"B5",X"8A",X"26",X"F5",X"4A",X"04",X"34",X"7E",X"75",X"C0",X"F5",
		X"7E",X"34",X"4A",X"AB",X"03",X"93",X"74",X"25",X"B5",X"7E",X"26",X"80",X"F2",X"04",X"F5",X"60",
		X"BB",X"91",X"7E",X"09",X"F5",X"FD",X"05",X"24",X"34",X"5B",X"21",X"FD",X"FD",X"00",X"FD",X"5A",
		X"01",X"6A",X"5F",X"34",X"FD",X"74",X"02",X"F5",X"5F",X"34",X"6A",X"5F",X"03",X"F5",X"75",X"04",
		X"F5",X"85",X"00",X"B3",X"7E",X"26",X"09",X"0F",X"B5",X"76",X"45",X"56",X"EA",X"0B",X"D5",X"BB",
		X"D1",X"B9",X"7E",X"26",X"F5",X"C1",X"06",X"C1",X"26",X"26",X"26",X"26",X"C2",X"88",X"E5",X"8F",
		X"26",X"5B",X"43",X"FD",X"B1",X"03",X"FD",X"5A",X"04",X"B1",X"5F",X"60",X"FD",X"63",X"05",X"DB",
		X"09",X"BB",X"00",X"BC",X"08",X"60",X"61",X"BB",X"41",X"6F",X"00",X"52",X"08",X"BD",X"4F",X"BB",
		X"60",X"34",X"6A",X"07",X"99",X"9E",X"74",X"4A",X"22",X"34",X"6A",X"07",X"34",X"9E",X"75",X"4A",
		X"23",X"34",X"6A",X"6F",X"34",X"B3",X"74",X"B3",X"6F",X"6A",X"6F",X"34",X"B3",X"75",X"57",X"B3",
		X"6F",X"6F",X"6F",X"B5",X"B3",X"77",X"B3",X"B9",X"44",X"01",X"F5",X"86",X"B1",X"F5",X"7E",X"02",
		X"17",X"5F",X"27",X"B3",X"9E",X"02",X"F5",X"68",X"B3",X"B3",X"B3",X"B1",X"68",X"68",X"68",X"6A",
		X"03",X"26",X"09",X"0F",X"35",X"B3",X"FD",X"B3",X"0F",X"B9",X"EA",X"B2",X"B5",X"B5",X"45",X"29",
		X"B1",X"B1",X"0B",X"7C",X"B5",X"B5",X"2A",X"2A",X"B1",X"B1",X"D5",X"2E",X"B5",X"B5",X"2A",X"2B",
		X"B1",X"B1",X"87",X"98",X"B5",X"B5",X"2B",X"2B",X"B1",X"B1",X"4E",X"A4",X"B5",X"B5",X"2C",X"2C",
		X"B1",X"B1",X"9D",X"6E",X"B5",X"B5",X"2C",X"2D",X"B1",X"B1",X"A2",X"D6",X"B5",X"B5",X"2D",X"2D",
		X"B1",X"B1",X"D7",X"F0",X"B5",X"B5",X"2D",X"2D",X"B1",X"B1",X"F1",X"4F",X"B5",X"D5",X"2D",X"6F",
		X"09",X"00",X"01",X"52",X"26",X"BD",X"46",X"7D",X"4F",X"01",X"09",X"72",X"6F",X"D1",X"40",X"46",
		X"00",X"77",X"52",X"7D",X"BD",X"B1",X"55",X"BE",X"03",X"C6",X"B1",X"B3",X"3F",X"34",X"09",X"16",
		X"B0",X"13",X"3E",X"A8",X"B3",X"09",X"28",X"34",X"7B",X"0B",X"0F",X"A6",X"86",X"7A",X"5F",X"0F",
		X"5F",X"A6",X"6E",X"5F",X"0B",X"0F",X"00",X"68",X"02",X"C6",X"4A",X"B3",X"60",X"34",X"09",X"3E",
		X"28",X"13",X"09",X"DF",X"43",X"41",X"DE",X"13",X"01",X"10",X"00",X"C8",X"05",X"BD",X"4E",X"AF",
		X"4A",X"60",X"13",X"9C",X"DE",X"09",X"60",X"13",X"41",X"05",X"13",X"4E",X"9D",X"00",X"01",X"10",
		X"BD",X"9C",X"AF",X"60",X"C8",X"13",X"4A",X"05",X"09",X"EB",X"34",X"C6",X"AB",X"09",X"60",X"34",
		X"B3",X"09",X"28",X"34",X"3E",X"AA",X"74",X"41",X"FB",X"34",X"6A",X"B5",X"13",X"DD",X"C9",X"63",
		X"40",X"BB",X"0B",X"8B",X"0B",X"2A",X"0B",X"34",X"D9",X"B3",X"04",X"B3",X"FE",X"0F",X"D0",X"0F",
		X"6C",X"45",X"B5",X"C8",X"6C",X"B5",X"EA",X"41",X"D0",X"6C",X"C8",X"C8",X"6A",X"4A",X"34",X"34",
		X"09",X"96",X"35",X"C6",X"08",X"09",X"B3",X"34",X"B3",X"6A",X"28",X"34",X"3E",X"C9",X"42",X"6C",
		X"4A",X"8E",X"34",X"6C",X"C9",X"34",X"6A",X"4A",X"8E",X"00",X"B5",X"6A",X"34",X"B1",X"43",X"CA");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
