library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_7M is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_7M is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"3C",X"62",X"62",X"73",X"00",X"00",X"00",X"60",X"72",X"7E",X"7E",X"7E",
		X"7F",X"73",X"73",X"3F",X"1E",X"00",X"00",X"00",X"78",X"CE",X"EE",X"F2",X"72",X"30",X"00",X"00",
		X"00",X"00",X"00",X"00",X"78",X"C4",X"C4",X"E6",X"00",X"00",X"08",X"34",X"76",X"77",X"7E",X"78",
		X"FE",X"E6",X"E6",X"7E",X"3C",X"00",X"00",X"00",X"78",X"E8",X"F4",X"F2",X"73",X"3E",X"0C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"12",X"23",X"3F",X"00",X"00",X"00",X"00",X"10",X"30",X"32",X"22",
		X"63",X"63",X"73",X"7F",X"7F",X"3F",X"1E",X"00",X"72",X"76",X"36",X"F6",X"F6",X"38",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"23",X"3F",X"00",X"00",X"00",X"00",X"14",X"34",X"36",X"26",
		X"63",X"63",X"73",X"7F",X"7F",X"3F",X"1E",X"00",X"76",X"72",X"74",X"F6",X"F6",X"3E",X"06",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"23",X"3F",X"00",X"00",X"00",X"00",X"12",X"36",X"36",X"26",
		X"63",X"63",X"73",X"7F",X"7F",X"3F",X"1E",X"00",X"76",X"70",X"30",X"F6",X"F6",X"3E",X"0E",X"0C",
		X"00",X"1E",X"3F",X"7F",X"7F",X"73",X"63",X"63",X"00",X"00",X"38",X"F6",X"F6",X"36",X"76",X"72",
		X"23",X"3F",X"12",X"00",X"00",X"00",X"00",X"00",X"22",X"32",X"30",X"10",X"00",X"00",X"00",X"00",
		X"00",X"1E",X"3F",X"7F",X"7F",X"73",X"63",X"63",X"00",X"06",X"3E",X"F6",X"F6",X"74",X"72",X"76",
		X"23",X"3F",X"02",X"00",X"00",X"00",X"00",X"00",X"26",X"36",X"34",X"14",X"00",X"00",X"00",X"00",
		X"00",X"1E",X"3F",X"7F",X"7F",X"73",X"63",X"63",X"0C",X"0E",X"3E",X"F6",X"F6",X"30",X"70",X"76",
		X"23",X"3F",X"02",X"00",X"00",X"00",X"00",X"00",X"26",X"36",X"36",X"12",X"00",X"00",X"00",X"00",
		X"00",X"07",X"0F",X"1C",X"3B",X"37",X"34",X"34",X"00",X"F0",X"F8",X"1C",X"6E",X"F6",X"96",X"96",
		X"34",X"37",X"3F",X"1C",X"0F",X"07",X"00",X"00",X"96",X"F6",X"FE",X"1C",X"F8",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"0F",X"1C",X"34",X"00",X"00",X"00",X"00",X"F0",X"F8",X"9C",X"96",
		X"34",X"37",X"37",X"18",X"0F",X"07",X"00",X"00",X"96",X"F6",X"F6",X"0C",X"F8",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"07",X"3F",X"3F",X"00",X"00",X"00",X"00",X"60",X"F0",X"F0",X"F0",
		X"3F",X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"07",X"04",X"04",X"00",X"00",X"00",X"00",X"F0",X"F8",X"98",X"90",
		X"04",X"27",X"30",X"18",X"0F",X"07",X"00",X"00",X"90",X"F0",X"00",X"00",X"F0",X"F0",X"00",X"00",
		X"00",X"07",X"0F",X"1C",X"3C",X"34",X"34",X"34",X"00",X"F0",X"F8",X"1C",X"1E",X"96",X"96",X"96",
		X"34",X"37",X"3F",X"1C",X"0F",X"07",X"00",X"00",X"96",X"F6",X"FE",X"1C",X"F8",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"0F",X"1C",X"34",X"00",X"00",X"00",X"00",X"F0",X"F8",X"9C",X"96",
		X"34",X"37",X"37",X"18",X"0F",X"07",X"00",X"00",X"96",X"F6",X"F6",X"0C",X"F8",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"04",X"3F",X"3F",X"00",X"00",X"00",X"00",X"10",X"90",X"F0",X"F0",
		X"3F",X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"07",X"04",X"04",X"00",X"00",X"00",X"00",X"F0",X"F8",X"98",X"90",
		X"04",X"27",X"30",X"18",X"0F",X"07",X"00",X"00",X"90",X"F0",X"00",X"00",X"F0",X"F0",X"00",X"00",
		X"00",X"07",X"0F",X"1C",X"3A",X"36",X"34",X"34",X"00",X"F0",X"F8",X"1C",X"6E",X"F6",X"96",X"96",
		X"34",X"37",X"3B",X"1C",X"0F",X"07",X"00",X"00",X"96",X"B6",X"2E",X"1C",X"F8",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"0F",X"1C",X"34",X"00",X"00",X"00",X"00",X"F0",X"F8",X"9C",X"96",
		X"34",X"37",X"33",X"18",X"0F",X"07",X"00",X"00",X"96",X"B6",X"26",X"0C",X"F8",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"06",X"3F",X"3F",X"00",X"00",X"00",X"00",X"60",X"F0",X"F0",X"F0",
		X"3F",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"F0",X"B0",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"07",X"04",X"04",X"00",X"00",X"00",X"00",X"F0",X"F8",X"98",X"90",
		X"04",X"27",X"30",X"18",X"0F",X"07",X"00",X"00",X"90",X"B0",X"00",X"00",X"F0",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"E0",X"71",X"79",X"F8",X"E0",X"00",X"00",X"00",X"80",X"C0",X"F8",X"FC",X"7C",
		X"F8",X"E0",X"F8",X"79",X"71",X"E0",X"00",X"00",X"F8",X"7C",X"FC",X"F8",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"E2",X"77",X"79",X"F8",X"C8",X"00",X"00",X"00",X"00",X"00",X"F8",X"FC",X"7C",
		X"F0",X"C8",X"F8",X"79",X"77",X"E2",X"00",X"00",X"F8",X"7C",X"FC",X"F8",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"1C",X"0E",X"0F",X"1F",X"3E",X"00",X"00",X"20",X"60",X"EC",X"7C",X"3C",X"18",
		X"3F",X"3E",X"1F",X"0F",X"0E",X"1C",X"00",X"00",X"38",X"18",X"3C",X"7C",X"EC",X"60",X"20",X"00",
		X"00",X"00",X"00",X"38",X"60",X"F8",X"FE",X"F0",X"00",X"00",X"C0",X"CC",X"5C",X"FC",X"78",X"F0",
		X"F2",X"7C",X"79",X"E1",X"00",X"00",X"00",X"00",X"F8",X"FC",X"FC",X"C8",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"38",X"60",X"F8",X"FE",X"F0",X"00",X"00",X"00",X"18",X"78",X"F8",X"7C",X"FC",
		X"F2",X"7C",X"79",X"E0",X"00",X"00",X"00",X"00",X"FC",X"EC",X"E0",X"60",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"38",X"60",X"F8",X"FE",X"F0",X"00",X"00",X"40",X"CC",X"5C",X"FC",X"78",X"F0",
		X"F2",X"7C",X"78",X"E0",X"00",X"00",X"00",X"00",X"F8",X"7C",X"18",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"38",X"60",X"F8",X"FE",X"F0",X"00",X"00",X"00",X"D8",X"78",X"F8",X"7C",X"EC",
		X"F2",X"7C",X"78",X"F0",X"00",X"00",X"00",X"00",X"E4",X"E0",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"F1",X"79",X"7C",X"F2",X"00",X"00",X"80",X"C0",X"C8",X"FC",X"FC",X"F8",
		X"F0",X"FE",X"F8",X"60",X"38",X"00",X"00",X"00",X"F0",X"78",X"FC",X"5C",X"CC",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"F0",X"79",X"7C",X"F2",X"00",X"00",X"00",X"00",X"60",X"E0",X"EC",X"FC",
		X"F0",X"FE",X"F8",X"60",X"38",X"00",X"00",X"00",X"FC",X"7C",X"F8",X"78",X"18",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"F0",X"78",X"7C",X"F2",X"00",X"00",X"00",X"C0",X"00",X"18",X"7C",X"F8",
		X"F0",X"FE",X"F8",X"60",X"38",X"00",X"00",X"00",X"F0",X"78",X"FC",X"5C",X"CC",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"F0",X"78",X"7C",X"F2",X"00",X"00",X"00",X"00",X"60",X"60",X"E0",X"E4",
		X"F0",X"FE",X"F8",X"60",X"38",X"00",X"00",X"00",X"EC",X"7C",X"FC",X"78",X"D8",X"00",X"00",X"00",
		X"00",X"00",X"00",X"71",X"3B",X"3C",X"7C",X"E4",X"00",X"00",X"00",X"00",X"80",X"FC",X"7E",X"3E",
		X"F8",X"E4",X"7C",X"3C",X"3B",X"71",X"00",X"00",X"7C",X"3E",X"7E",X"FC",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"38",X"1D",X"1E",X"3E",X"7C",X"00",X"00",X"00",X"80",X"C0",X"7C",X"3E",X"1E",
		X"7C",X"7C",X"3E",X"1E",X"1D",X"38",X"00",X"00",X"3C",X"1E",X"3E",X"7C",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"38",X"48",X"FB",X"FE",X"F8",X"F8",X"40",X"E0",X"C0",X"48",X"7C",X"7E",X"7E",X"7E",
		X"7E",X"3C",X"39",X"71",X"00",X"00",X"00",X"00",X"7C",X"FC",X"9C",X"C0",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"01",X"03",X"E3",X"7A",X"79",X"E0",X"00",X"00",X"0C",X"9E",X"BE",X"FC",X"F8",X"FC",
		X"F8",X"F0",X"FC",X"FC",X"7D",X"3C",X"38",X"70",X"FC",X"FC",X"FC",X"F8",X"C8",X"E0",X"60",X"00",
		X"00",X"00",X"00",X"00",X"01",X"71",X"3C",X"3E",X"00",X"00",X"00",X"C0",X"C0",X"9C",X"FC",X"7C",
		X"79",X"F8",X"FE",X"FB",X"48",X"38",X"00",X"00",X"7E",X"7E",X"7E",X"7C",X"48",X"C0",X"E0",X"40",
		X"70",X"38",X"3C",X"73",X"FC",X"FC",X"F0",X"F8",X"00",X"60",X"E0",X"C0",X"F8",X"FC",X"FC",X"FC",
		X"E0",X"79",X"7A",X"E3",X"03",X"01",X"00",X"00",X"FC",X"F8",X"FC",X"BE",X"9E",X"0C",X"00",X"00",
		X"43",X"47",X"41",X"64",X"66",X"67",X"67",X"77",X"0F",X"FC",X"F0",X"40",X"00",X"80",X"80",X"80",
		X"77",X"63",X"63",X"42",X"06",X"07",X"04",X"04",X"80",X"80",X"00",X"00",X"00",X"00",X"C0",X"20",
		X"04",X"27",X"27",X"37",X"37",X"3F",X"3F",X"3F",X"00",X"E0",X"FE",X"F0",X"80",X"80",X"80",X"80",
		X"3F",X"3B",X"33",X"00",X"06",X"07",X"04",X"04",X"80",X"80",X"00",X"00",X"00",X"00",X"C0",X"20",
		X"00",X"17",X"19",X"1C",X"1F",X"1F",X"1F",X"1F",X"00",X"80",X"C0",X"70",X"58",X"00",X"80",X"80",
		X"1F",X"1F",X"1F",X"12",X"06",X"07",X"04",X"04",X"80",X"80",X"00",X"00",X"00",X"00",X"C0",X"20",
		X"10",X"20",X"20",X"40",X"60",X"18",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2F",
		X"04",X"0F",X"7F",X"40",X"20",X"20",X"10",X"00",X"FC",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"06",X"08",X"10",X"10",X"18",X"08",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2E",
		X"04",X"0F",X"1F",X"10",X"10",X"08",X"06",X"00",X"F8",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"07",X"18",X"10",X"10",X"18",X"08",X"0C",X"0C",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"2C",
		X"04",X"0F",X"1F",X"10",X"10",X"18",X"07",X"00",X"F0",X"C0",X"80",X"00",X"00",X"00",X"80",X"00",
		X"40",X"47",X"60",X"67",X"77",X"77",X"63",X"43",X"00",X"FE",X"F8",X"60",X"80",X"80",X"80",X"80",
		X"67",X"7B",X"7A",X"67",X"07",X"04",X"04",X"00",X"80",X"00",X"00",X"00",X"80",X"C0",X"20",X"00",
		X"00",X"04",X"04",X"07",X"67",X"7A",X"7B",X"67",X"00",X"20",X"C0",X"80",X"00",X"00",X"00",X"80",
		X"43",X"63",X"77",X"77",X"67",X"60",X"47",X"40",X"80",X"80",X"80",X"80",X"60",X"F8",X"FE",X"00",
		X"00",X"00",X"00",X"E0",X"71",X"79",X"F8",X"E0",X"00",X"00",X"40",X"E0",X"80",X"98",X"FC",X"7C",
		X"F0",X"E0",X"F8",X"79",X"71",X"E0",X"00",X"00",X"F8",X"7C",X"FC",X"98",X"80",X"E0",X"40",X"00",
		X"00",X"00",X"01",X"71",X"39",X"3D",X"7F",X"F8",X"00",X"00",X"80",X"80",X"8C",X"FC",X"FC",X"F8",
		X"F8",X"E0",X"F0",X"60",X"78",X"F0",X"00",X"00",X"78",X"F8",X"7C",X"DC",X"CC",X"C0",X"C0",X"00",
		X"00",X"00",X"00",X"E2",X"77",X"79",X"F8",X"C8",X"00",X"00",X"00",X"00",X"00",X"F8",X"FC",X"7C",
		X"F0",X"C8",X"F8",X"79",X"77",X"E2",X"00",X"00",X"F8",X"7C",X"FC",X"F8",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0E",X"1E",X"3E",X"7C",X"7D",X"7B",X"00",X"00",X"00",X"00",X"40",X"C0",X"C0",X"80",
		X"7B",X"7D",X"7D",X"3E",X"1E",X"0F",X"03",X"00",X"80",X"C0",X"C0",X"E0",X"F0",X"90",X"E0",X"00",
		X"00",X"00",X"0E",X"1E",X"3E",X"7C",X"7D",X"7B",X"00",X"00",X"00",X"00",X"43",X"C1",X"C1",X"80",
		X"7B",X"7D",X"7D",X"3E",X"1E",X"0F",X"03",X"00",X"80",X"C1",X"C1",X"E3",X"F7",X"91",X"E0",X"00",
		X"00",X"00",X"0E",X"1F",X"3F",X"7F",X"7F",X"7F",X"00",X"00",X"00",X"80",X"C0",X"C0",X"E0",X"E0",
		X"7F",X"7F",X"7F",X"3F",X"1F",X"0F",X"03",X"00",X"E0",X"E0",X"E0",X"F0",X"F0",X"F0",X"E0",X"00",
		X"00",X"00",X"1C",X"3C",X"58",X"09",X"9B",X"F7",X"00",X"00",X"00",X"00",X"84",X"82",X"88",X"04",
		X"F7",X"FB",X"FB",X"7D",X"3D",X"1F",X"07",X"00",X"0A",X"94",X"84",X"C2",X"EC",X"24",X"CA",X"00",
		X"C0",X"C0",X"30",X"30",X"37",X"2E",X"0E",X"1D",X"00",X"02",X"04",X"0A",X"04",X"82",X"C6",X"CE",
		X"0D",X"0B",X"02",X"05",X"02",X"00",X"00",X"00",X"8E",X"7E",X"FE",X"3C",X"1C",X"1C",X"38",X"00",
		X"C0",X"80",X"70",X"68",X"1E",X"1D",X"1B",X"1B",X"00",X"00",X"02",X"04",X"02",X"84",X"A6",X"8E",
		X"07",X"07",X"06",X"05",X"02",X"00",X"00",X"00",X"0E",X"7E",X"FE",X"3C",X"1C",X"1C",X"38",X"00",
		X"40",X"C0",X"60",X"58",X"1C",X"3B",X"1B",X"17",X"00",X"00",X"00",X"02",X"04",X"82",X"66",X"4E",
		X"06",X"0D",X"04",X"04",X"02",X"00",X"00",X"00",X"BE",X"7E",X"FE",X"1C",X"1C",X"1C",X"18",X"00",
		X"C0",X"C0",X"50",X"5C",X"3A",X"37",X"16",X"0E",X"00",X"00",X"00",X"00",X"02",X"00",X"E6",X"CE",
		X"0D",X"0D",X"02",X"01",X"02",X"00",X"00",X"00",X"8E",X"7E",X"FE",X"3C",X"1C",X"1C",X"38",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"3B",X"00",X"00",X"40",X"70",X"78",X"78",X"7C",X"7C",
		X"3A",X"38",X"18",X"1E",X"0E",X"02",X"00",X"00",X"7C",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"07",X"0F",X"1F",X"3F",X"3F",X"3E",X"00",X"00",X"E0",X"F0",X"D8",X"DC",X"8C",X"0C",
		X"3F",X"3F",X"3E",X"1F",X"0F",X"07",X"00",X"00",X"8C",X"8C",X"1C",X"D8",X"F0",X"E0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"E2",X"77",X"79",X"F8",X"C8",X"00",X"00",X"00",X"00",X"00",X"F8",X"FC",X"7C",
		X"F0",X"C8",X"F8",X"79",X"77",X"E2",X"00",X"00",X"F8",X"7C",X"FC",X"F8",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"1D",X"0F",X"1F",X"3F",X"3F",X"00",X"00",X"C0",X"C0",X"80",X"F8",X"FC",X"7C",
		X"3F",X"3F",X"3F",X"1F",X"0F",X"1D",X"00",X"00",X"78",X"7C",X"FC",X"F8",X"80",X"C0",X"C0",X"00",
		X"00",X"00",X"00",X"01",X"00",X"41",X"63",X"43",X"00",X"00",X"00",X"C0",X"FC",X"FE",X"F4",X"E0",
		X"03",X"63",X"43",X"41",X"00",X"01",X"00",X"00",X"E0",X"E0",X"F4",X"FE",X"FC",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"0F",X"00",X"00",X"00",X"40",X"E0",X"E0",X"F0",X"E0",
		X"03",X"0F",X"0F",X"07",X"01",X"00",X"00",X"00",X"F0",X"E0",X"E0",X"F0",X"E0",X"40",X"00",X"00",
		X"00",X"00",X"00",X"70",X"3B",X"3E",X"7C",X"EC",X"00",X"00",X"00",X"80",X"D8",X"FC",X"7E",X"3E",
		X"F8",X"EC",X"7C",X"3E",X"3B",X"70",X"00",X"00",X"7E",X"3E",X"7E",X"FC",X"D8",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"1F",X"3F",X"3F",X"7F",X"7F",X"00",X"00",X"00",X"00",X"C0",X"E0",X"F0",X"F0",
		X"7F",X"7F",X"3F",X"3F",X"1F",X"0F",X"03",X"00",X"F8",X"F8",X"F8",X"F8",X"F8",X"F0",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"0F",X"1F",X"17",X"00",X"00",X"00",X"00",X"00",X"1C",X"22",X"41",
		X"17",X"17",X"1F",X"0F",X"07",X"09",X"11",X"01",X"51",X"59",X"22",X"3C",X"BC",X"B8",X"80",X"80",
		X"00",X"00",X"00",X"00",X"04",X"27",X"17",X"17",X"00",X"00",X"00",X"00",X"00",X"1C",X"22",X"41",
		X"1F",X"1F",X"1F",X"1F",X"27",X"01",X"01",X"00",X"51",X"59",X"22",X"3C",X"BC",X"B8",X"80",X"00",
		X"00",X"00",X"00",X"00",X"04",X"0F",X"1F",X"1F",X"00",X"00",X"00",X"00",X"00",X"1C",X"22",X"41",
		X"7F",X"1F",X"1F",X"0F",X"07",X"00",X"00",X"00",X"51",X"59",X"22",X"3C",X"BC",X"38",X"00",X"00",
		X"00",X"00",X"00",X"40",X"24",X"1F",X"1F",X"1F",X"00",X"00",X"00",X"00",X"00",X"1C",X"22",X"41",
		X"1F",X"17",X"17",X"27",X"07",X"01",X"00",X"00",X"51",X"59",X"62",X"3C",X"BC",X"B8",X"00",X"00",
		X"00",X"00",X"02",X"02",X"03",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"E0",X"00",X"00",X"00",
		X"00",X"08",X"0C",X"06",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",
		X"00",X"00",X"03",X"02",X"02",X"02",X"03",X"00",X"00",X"00",X"E0",X"20",X"20",X"20",X"E0",X"00",
		X"00",X"08",X"0C",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"02",X"02",X"02",X"00",X"00",X"00",X"00",X"E0",X"20",X"20",X"20",
		X"03",X"08",X"0C",X"06",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"20",
		X"02",X"0A",X"0F",X"06",X"00",X"00",X"00",X"00",X"20",X"20",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"0A",X"0E",X"06",X"03",X"00",X"00",X"00",X"E0",X"20",X"20",X"20",X"E0",X"00",X"00",X"00",
		X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"0F",X"06",X"02",X"02",X"01",X"00",X"00",X"00",X"E0",X"20",X"20",X"20",X"C0",X"00",
		X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"0C",X"06",X"03",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"20",X"00",X"00",
		X"00",X"00",X"02",X"02",X"03",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"E0",X"00",X"00",X"00",
		X"00",X"08",X"0C",X"06",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",
		X"00",X"00",X"00",X"1F",X"3F",X"3F",X"7F",X"7F",X"00",X"00",X"00",X"00",X"C0",X"E0",X"F0",X"F0",
		X"7C",X"7E",X"3F",X"3F",X"1F",X"0F",X"03",X"00",X"F8",X"F8",X"F8",X"F8",X"F8",X"F0",X"C0",X"00",
		X"00",X"00",X"00",X"1F",X"3F",X"3F",X"7F",X"7E",X"00",X"00",X"00",X"00",X"C0",X"E0",X"F0",X"F0",
		X"78",X"7C",X"3E",X"3F",X"1F",X"0F",X"03",X"00",X"78",X"F8",X"F8",X"F8",X"F8",X"F0",X"C0",X"00",
		X"00",X"00",X"00",X"1F",X"3F",X"3F",X"7F",X"78",X"00",X"00",X"00",X"00",X"C0",X"E0",X"F0",X"70",
		X"78",X"78",X"3C",X"3F",X"1F",X"0F",X"03",X"00",X"78",X"78",X"78",X"F8",X"F8",X"F0",X"C0",X"00",
		X"00",X"00",X"00",X"1F",X"3F",X"3F",X"7C",X"70",X"00",X"00",X"00",X"00",X"C0",X"E0",X"70",X"30",
		X"70",X"70",X"38",X"3C",X"1F",X"0F",X"03",X"00",X"38",X"38",X"78",X"78",X"F8",X"F0",X"C0",X"00",
		X"00",X"00",X"00",X"0A",X"1E",X"1E",X"3A",X"3A",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"C0",
		X"3A",X"3A",X"1E",X"1E",X"0A",X"02",X"00",X"00",X"C0",X"C0",X"C0",X"E0",X"F0",X"F0",X"E0",X"C0",
		X"00",X"00",X"00",X"0E",X"1E",X"1A",X"3A",X"3A",X"00",X"20",X"30",X"30",X"20",X"C0",X"C0",X"C0",
		X"3A",X"3E",X"1E",X"1A",X"0A",X"02",X"00",X"00",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"00",X"00",X"04",X"0E",X"1A",X"1A",X"3A",X"3A",X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",X"F0",
		X"3E",X"3E",X"1A",X"1A",X"0A",X"02",X"00",X"00",X"F0",X"E0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"00",X"00",X"04",X"0A",X"1A",X"1A",X"3A",X"3E",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"C0",
		X"3E",X"3A",X"1A",X"1A",X"0A",X"06",X"00",X"00",X"C0",X"C0",X"C0",X"E0",X"F0",X"F0",X"E0",X"C0",
		X"00",X"00",X"00",X"08",X"18",X"1A",X"3E",X"3E",X"00",X"20",X"30",X"30",X"20",X"C0",X"C0",X"C0",
		X"3A",X"3A",X"1A",X"1A",X"0E",X"06",X"00",X"00",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"00",X"00",X"00",X"00",X"1A",X"1E",X"3E",X"3A",X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",X"F0",
		X"3A",X"3A",X"1A",X"1E",X"0E",X"02",X"00",X"00",X"F0",X"E0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"04",X"07",X"0F",X"0F",X"7E",X"78",X"00",X"00",X"20",X"00",X"C0",X"EC",X"70",X"10",
		X"78",X"7C",X"3E",X"07",X"07",X"07",X"03",X"00",X"18",X"38",X"7C",X"F0",X"C0",X"C0",X"C0",X"00",
		X"00",X"02",X"01",X"01",X"21",X"33",X"7F",X"1F",X"00",X"00",X"00",X"00",X"C0",X"E0",X"90",X"08",
		X"1E",X"3F",X"37",X"23",X"01",X"01",X"03",X"00",X"08",X"08",X"98",X"F8",X"F0",X"F0",X"C0",X"00",
		X"00",X"00",X"00",X"10",X"38",X"3C",X"1F",X"0F",X"00",X"80",X"40",X"40",X"C0",X"F8",X"E4",X"82",
		X"0F",X"0F",X"1F",X"38",X"10",X"00",X"00",X"00",X"82",X"C4",X"E0",X"F8",X"78",X"70",X"C0",X"00",
		X"00",X"00",X"00",X"1C",X"3E",X"3F",X"0F",X"07",X"00",X"00",X"10",X"10",X"20",X"24",X"F8",X"E0",
		X"07",X"07",X"0F",X"3E",X"1C",X"0C",X"02",X"00",X"E0",X"F0",X"F8",X"38",X"18",X"10",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"1F",X"3F",X"79",X"70",X"00",X"40",X"80",X"08",X"88",X"C0",X"F0",X"F0",
		X"60",X"70",X"39",X"1F",X"0F",X"0F",X"03",X"00",X"F8",X"F8",X"F8",X"88",X"00",X"00",X"80",X"00",
		X"00",X"02",X"01",X"03",X"27",X"3F",X"78",X"78",X"00",X"00",X"00",X"00",X"C0",X"E0",X"70",X"30",
		X"78",X"7C",X"2E",X"07",X"07",X"07",X"03",X"00",X"3C",X"22",X"64",X"C0",X"C0",X"C0",X"C0",X"00",
		X"00",X"01",X"01",X"03",X"33",X"3E",X"7F",X"7F",X"00",X"00",X"00",X"60",X"10",X"08",X"08",X"00",
		X"7F",X"67",X"23",X"21",X"13",X"0F",X"03",X"00",X"8E",X"F8",X"E0",X"C0",X"C0",X"E0",X"C0",X"00",
		X"00",X"02",X"02",X"03",X"07",X"07",X"7F",X"7F",X"00",X"00",X"30",X"08",X"04",X"84",X"C0",X"E0",
		X"63",X"41",X"20",X"30",X"19",X"0F",X"03",X"00",X"FC",X"F2",X"E0",X"C0",X"C0",X"C0",X"C0",X"00",
		X"00",X"02",X"02",X"03",X"07",X"0F",X"0F",X"7F",X"00",X"00",X"00",X"00",X"C0",X"E0",X"F0",X"F0",
		X"60",X"60",X"20",X"10",X"08",X"07",X"03",X"00",X"F8",X"78",X"64",X"C0",X"80",X"80",X"C0",X"00",
		X"03",X"07",X"07",X"07",X"03",X"07",X"07",X"07",X"E0",X"E0",X"E0",X"C0",X"E0",X"E0",X"E0",X"C0",
		X"00",X"03",X"07",X"04",X"00",X"00",X"00",X"00",X"20",X"E0",X"E0",X"40",X"00",X"00",X"00",X"00",
		X"03",X"07",X"07",X"07",X"03",X"07",X"07",X"07",X"E0",X"E0",X"E0",X"C0",X"E0",X"E0",X"E0",X"C0",
		X"03",X"07",X"07",X"05",X"00",X"00",X"00",X"00",X"A0",X"E0",X"E0",X"C0",X"00",X"00",X"00",X"00",
		X"03",X"07",X"07",X"07",X"03",X"07",X"07",X"07",X"E0",X"E0",X"E0",X"C0",X"E0",X"E0",X"E0",X"C0",
		X"03",X"07",X"07",X"05",X"00",X"00",X"00",X"00",X"E0",X"E0",X"E0",X"40",X"00",X"00",X"00",X"00",
		X"03",X"07",X"07",X"07",X"03",X"07",X"07",X"07",X"E0",X"E0",X"E0",X"C0",X"E0",X"E0",X"E0",X"C0",
		X"02",X"07",X"07",X"07",X"00",X"00",X"00",X"00",X"E0",X"E0",X"E0",X"40",X"00",X"00",X"00",X"00",
		X"03",X"07",X"07",X"07",X"03",X"07",X"07",X"07",X"E0",X"E0",X"E0",X"C0",X"E0",X"E0",X"E0",X"C0",
		X"02",X"07",X"07",X"07",X"00",X"00",X"00",X"00",X"E0",X"E0",X"E0",X"40",X"00",X"00",X"00",X"00",
		X"03",X"07",X"07",X"07",X"03",X"07",X"07",X"07",X"E0",X"E0",X"E0",X"C0",X"E0",X"E0",X"E0",X"C0",
		X"03",X"07",X"07",X"07",X"00",X"03",X"07",X"04",X"E0",X"E0",X"E0",X"C0",X"20",X"E0",X"E0",X"40",
		X"03",X"07",X"07",X"07",X"03",X"07",X"07",X"07",X"E0",X"E0",X"E0",X"C0",X"E0",X"E0",X"E0",X"C0",
		X"03",X"07",X"07",X"07",X"00",X"00",X"00",X"00",X"E0",X"E0",X"E0",X"C0",X"00",X"00",X"00",X"00",
		X"03",X"07",X"07",X"07",X"03",X"07",X"07",X"07",X"E0",X"E0",X"E0",X"C0",X"E0",X"E0",X"E0",X"C0",
		X"03",X"07",X"07",X"07",X"00",X"03",X"07",X"04",X"E0",X"E0",X"E0",X"C0",X"20",X"E0",X"E0",X"40",
		X"03",X"07",X"07",X"07",X"03",X"07",X"07",X"07",X"E0",X"E0",X"E0",X"C0",X"E0",X"E0",X"E0",X"C0",
		X"03",X"07",X"07",X"05",X"00",X"03",X"07",X"04",X"A0",X"E0",X"E0",X"C0",X"20",X"E0",X"E0",X"40",
		X"03",X"07",X"07",X"07",X"03",X"07",X"07",X"07",X"E0",X"E0",X"E0",X"C0",X"E0",X"E0",X"E0",X"C0",
		X"03",X"07",X"07",X"07",X"03",X"07",X"07",X"05",X"E0",X"E0",X"E0",X"C0",X"E0",X"E0",X"E0",X"40",
		X"03",X"07",X"07",X"07",X"03",X"07",X"07",X"07",X"E0",X"E0",X"E0",X"C0",X"E0",X"E0",X"E0",X"C0",
		X"03",X"07",X"07",X"07",X"03",X"07",X"07",X"05",X"E0",X"E0",X"E0",X"C0",X"A0",X"E0",X"E0",X"C0",
		X"03",X"07",X"07",X"07",X"03",X"07",X"07",X"07",X"E0",X"E0",X"E0",X"C0",X"E0",X"E0",X"E0",X"C0",
		X"03",X"07",X"07",X"07",X"03",X"07",X"07",X"07",X"E0",X"E0",X"E0",X"C0",X"E0",X"E0",X"E0",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"07",X"07",X"05",X"00",X"01",X"00",X"01",X"A0",X"E0",X"E0",X"C0",X"A0",X"40",X"A0",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"07",X"07",X"05",X"00",X"01",X"00",X"01",X"E0",X"E0",X"E0",X"40",X"A0",X"40",X"A0",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"03",X"03",X"07",X"00",X"01",X"00",X"01",X"E0",X"C0",X"C0",X"80",X"A0",X"40",X"A0",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"07",X"07",X"07",X"00",X"01",X"00",X"01",X"E0",X"E0",X"E0",X"40",X"A0",X"40",X"A0",X"40",
		X"00",X"00",X"00",X"00",X"08",X"04",X"02",X"01",X"00",X"00",X"00",X"10",X"11",X"11",X"01",X"01",
		X"00",X"00",X"00",X"1C",X"00",X"00",X"00",X"0F",X"08",X"08",X"25",X"11",X"C9",X"20",X"03",X"3B",
		X"00",X"00",X"00",X"08",X"88",X"88",X"80",X"80",X"00",X"00",X"00",X"00",X"10",X"20",X"40",X"80",
		X"10",X"10",X"A4",X"88",X"93",X"04",X"C0",X"DC",X"00",X"00",X"00",X"38",X"00",X"00",X"00",X"F0",
		X"0F",X"00",X"00",X"00",X"1C",X"00",X"00",X"00",X"3B",X"03",X"20",X"C9",X"11",X"25",X"08",X"08",
		X"01",X"02",X"04",X"08",X"00",X"00",X"00",X"00",X"01",X"01",X"11",X"11",X"10",X"00",X"00",X"00",
		X"DC",X"C0",X"04",X"93",X"88",X"A4",X"10",X"10",X"F0",X"00",X"00",X"00",X"38",X"00",X"00",X"00",
		X"80",X"80",X"88",X"88",X"08",X"00",X"00",X"00",X"80",X"40",X"20",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"20",X"10",X"08",X"04",X"00",X"00",X"00",X"01",X"21",X"21",X"20",X"01",X"01",X"11",
		X"00",X"00",X"1C",X"01",X"00",X"00",X"00",X"73",X"90",X"48",X"20",X"80",X"40",X"00",X"00",X"80",
		X"00",X"80",X"80",X"84",X"04",X"04",X"80",X"88",X"00",X"00",X"04",X"08",X"10",X"20",X"00",X"00",
		X"89",X"12",X"04",X"01",X"02",X"00",X"00",X"00",X"00",X"00",X"1C",X"80",X"00",X"00",X"00",X"EE",
		X"77",X"00",X"00",X"00",X"01",X"38",X"00",X"00",X"00",X"00",X"00",X"40",X"80",X"20",X"48",X"91",
		X"00",X"00",X"04",X"08",X"10",X"20",X"00",X"00",X"11",X"01",X"20",X"20",X"21",X"01",X"01",X"00",
		X"01",X"00",X"00",X"02",X"01",X"04",X"12",X"09",X"CE",X"00",X"00",X"00",X"80",X"38",X"00",X"00",
		X"88",X"80",X"80",X"04",X"84",X"84",X"80",X"00",X"00",X"00",X"20",X"10",X"08",X"04",X"00",X"00",
		X"00",X"40",X"20",X"10",X"00",X"00",X"02",X"01",X"81",X"81",X"01",X"00",X"21",X"21",X"00",X"00",
		X"60",X"00",X"0C",X"00",X"00",X"00",X"00",X"EC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"81",X"81",X"00",X"84",X"84",X"00",X"00",X"00",X"02",X"04",X"08",X"00",X"00",X"40",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"30",X"00",X"00",X"00",X"00",X"37",
		X"EC",X"00",X"00",X"00",X"00",X"0C",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"02",X"00",X"00",X"10",X"20",X"40",X"00",X"00",X"00",X"21",X"21",X"00",X"81",X"81",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"37",X"00",X"00",X"00",X"00",X"30",X"00",X"06",
		X"00",X"00",X"84",X"84",X"00",X"80",X"81",X"81",X"80",X"40",X"00",X"00",X"08",X"04",X"02",X"00",
		X"00",X"40",X"20",X"10",X"00",X"00",X"00",X"00",X"81",X"81",X"01",X"00",X"00",X"00",X"00",X"00",
		X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"81",X"81",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"04",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"07",
		X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"20",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"81",X"81",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"06",
		X"00",X"00",X"00",X"00",X"00",X"80",X"81",X"81",X"00",X"00",X"00",X"00",X"08",X"04",X"02",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"1F",X"3F",X"3E",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"E7",X"CE",X"9E",X"1F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"3F",X"1F",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"1F",X"9E",X"CE",X"E7",X"40",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"3F",X"1F",X"0E",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"47",X"EE",X"9E",X"1F",X"0B",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"1F",X"3F",X"18",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0B",X"1F",X"9E",X"EE",X"47",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"78",X"38",X"08",X"04",X"0E",X"0A",X"00",X"00",X"01",X"03",X"06",X"04",X"47",X"57",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"8F",X"1F",X"6F",X"CF",X"8D",X"87",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"04",X"08",X"38",X"78",X"F0",X"F0",X"A0",X"47",X"04",X"06",X"03",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"8D",X"CF",X"6F",X"1F",X"8F",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"07",X"07",X"0E",X"00",X"00",X"00",X"00",X"C0",X"00",X"80",X"00",
		X"0C",X"0C",X"0C",X"08",X"08",X"04",X"0E",X"0A",X"00",X"00",X"00",X"06",X"07",X"07",X"43",X"51",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"1F",X"3F",X"EF",X"CF",X"8D",X"87",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"04",X"08",X"08",X"0C",X"0C",X"0C",X"0E",X"43",X"07",X"07",X"06",X"00",X"00",X"00",X"00",
		X"07",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"8D",X"CF",X"EF",X"3F",X"1F",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"F8",X"F9",X"F1",X"F1",X"F3",X"F3",X"E3",X"E7",
		X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"E7",X"EF",X"EF",X"EF",X"EF",X"EF",X"E7",X"F7",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"FC",X"C0",X"C0",X"C0",X"C0",X"00",X"40",X"00",X"00",
		X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"F7",X"F7",X"F3",X"F8",X"FE",X"FF",X"FF",X"FF",
		X"5F",X"5F",X"4F",X"27",X"33",X"18",X"07",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"00",
		X"FC",X"FC",X"FC",X"FC",X"38",X"88",X"E0",X"F8",X"00",X"00",X"00",X"1C",X"1F",X"1F",X"7F",X"7F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"00",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"07",X"01",X"1C",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"06",X"00",X"00",X"00",X"3C",X"3F",X"7F",X"7F",X"70",X"30",X"10",X"10",X"00",X"80",X"F0",X"F0",
		X"0F",X"0F",X"0F",X"07",X"07",X"07",X"03",X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"03",X"03",X"03",X"01",X"01",X"01",X"01",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"7F",X"7F",X"3F",X"87",X"F0",X"FE",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"10",X"C0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"00",X"F8",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"03",X"C3",X"FF",X"FF",X"00",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"00",
		X"5F",X"5F",X"5E",X"5E",X"5A",X"5B",X"59",X"5C",X"F8",X"F9",X"FB",X"FB",X"7B",X"38",X"3F",X"9F",
		X"5C",X"5E",X"58",X"5E",X"5F",X"40",X"58",X"5C",X"8F",X"45",X"01",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"F8",X"F8",X"F0",X"F0",X"60",X"00",X"E0",X"07",X"0F",X"0F",X"1F",X"1F",X"1F",X"3F",X"3E",
		X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"04",X"20",X"80",X"40",X"00",X"00",X"00",X"00",X"00",
		X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"80",X"80",X"00",X"E0",X"E0",X"E4",X"E5",X"F7",
		X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"F7",X"FF",X"FF",X"FE",X"FE",X"FC",X"FC",X"F8",
		X"0E",X"1E",X"3E",X"9E",X"CF",X"6F",X"3F",X"B8",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",
		X"E0",X"80",X"1E",X"3F",X"7F",X"7F",X"7F",X"FF",X"00",X"00",X"00",X"80",X"C0",X"E0",X"E0",X"E0",
		X"C1",X"C0",X"00",X"C0",X"81",X"81",X"83",X"00",X"00",X"3F",X"00",X"00",X"00",X"F0",X"F0",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"FF",X"FF",X"0F",X"0F",X"0F",X"0F",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"1F",X"1F",X"3F",X"3F",X"1F",X"1F",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"41",X"49",X"49",X"49",X"7F",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"7F",X"38",X"1C",X"38",X"7F",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"39",X"7B",X"4F",X"46",X"44",X"7F",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"41",X"49",X"49",X"49",X"7F",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"3F",X"64",X"44",X"64",X"3F",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"4F",X"4F",X"49",X"49",X"63",X"3E",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"78",X"7C",X"0E",X"07",X"0E",X"7C",X"78",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3E",X"7F",X"41",X"41",X"41",X"7F",X"3E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"03",X"07",X"0F",X"1F",X"3F",X"7E",X"FC",X"FF",X"FF",X"FF",X"FF",X"80",X"00",X"00",X"00",
		X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"00",X"00",X"80",X"C0",X"E0",X"F0",X"F8",X"FC",X"7E",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"7E",X"3F",X"1F",X"0F",X"07",X"03",X"01",X"00",X"00",X"00",X"80",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"1F",
		X"00",X"00",X"00",X"01",X"FF",X"FF",X"FF",X"FF",X"3F",X"7E",X"FC",X"F8",X"F0",X"E0",X"C0",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"F7",X"F7",X"F6",X"F0",X"F0",X"F0",X"F8",X"F9",
		X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"FC",X"FE",X"FE",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"F8",X"C0",X"00",X"00",X"04",X"1C",X"7C",X"FE",X"03",X"08",X"3E",X"F8",X"E1",X"43",X"07",X"0E",
		X"78",X"10",X"00",X"00",X"00",X"04",X"1F",X"3E",X"00",X"38",X"7F",X"00",X"00",X"00",X"00",X"07",
		X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"F8",X"F8",X"FB",X"FB",X"F9",X"FC",X"FF",X"FF",
		X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"FF",X"FF",X"FF",X"FE",X"FE",X"F8",X"F8",X"F8",
		X"7C",X"F8",X"F0",X"E0",X"C0",X"00",X"00",X"C1",X"0F",X"0F",X"1E",X"3C",X"7C",X"F8",X"F0",X"F0",
		X"F1",X"FC",X"E0",X"00",X"00",X"3F",X"7E",X"FC",X"E0",X"41",X"01",X"01",X"03",X"03",X"07",X"07",
		X"00",X"00",X"00",X"60",X"C0",X"85",X"09",X"09",X"54",X"54",X"54",X"14",X"94",X"94",X"B2",X"B2",
		X"13",X"33",X"07",X"01",X"00",X"00",X"00",X"90",X"32",X"32",X"32",X"32",X"32",X"02",X"00",X"00",
		X"7F",X"7F",X"7F",X"3F",X"3F",X"3F",X"3F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"C0",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"FF",X"3F",X"3F",X"C1",X"01",X"70",X"78",X"3C",X"3E",X"1F",X"0F",
		X"1C",X"1C",X"3C",X"3C",X"78",X"78",X"38",X"88",X"40",X"70",X"70",X"70",X"70",X"70",X"F0",X"F0",
		X"E0",X"F0",X"F0",X"F0",X"E0",X"E0",X"E1",X"E1",X"30",X"00",X"00",X"80",X"E0",X"F0",X"F0",X"F0",
		X"3F",X"3F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"07",X"03",X"03",X"41",X"60",X"60",X"00",X"FF",
		X"7F",X"7F",X"FF",X"3F",X"0F",X"0F",X"0F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"FC",X"F8",
		X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"F8",X"FB",X"F3",X"F7",X"F0",X"F0",X"F0",X"F7",
		X"F0",X"C0",X"80",X"18",X"7F",X"FF",X"3F",X"07",X"7F",X"1F",X"07",X"02",X"00",X"C1",X"E0",X"F6",
		X"00",X"C0",X"FE",X"FC",X"00",X"00",X"3C",X"FC",X"77",X"07",X"60",X"3F",X"80",X"0F",X"08",X"01",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"CC",X"CE",X"CE",X"CE",X"CE",X"86",X"80",X"00",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"80",X"8C",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"03",X"00",X"00",X"00",X"38",X"38",X"30",X"38",X"F3",X"77",X"F0",X"1E",X"10",X"00",X"00",X"20",
		X"19",X"01",X"11",X"1C",X"07",X"00",X"00",X"C0",X"60",X"40",X"80",X"03",X"07",X"C6",X"10",X"00",
		X"E0",X"80",X"00",X"3A",X"9C",X"CC",X"76",X"1A",X"4D",X"4D",X"69",X"69",X"2B",X"AA",X"AA",X"AB",
		X"84",X"E2",X"3C",X"FF",X"00",X"85",X"33",X"08",X"AA",X"AA",X"47",X"08",X"07",X"D0",X"64",X"B4",
		X"98",X"10",X"21",X"43",X"06",X"8C",X"19",X"33",X"00",X"00",X"C0",X"84",X"1F",X"7E",X"E0",X"07",
		X"64",X"87",X"40",X"07",X"C7",X"07",X"1F",X"1F",X"7F",X"FC",X"00",X"00",X"F1",X"FC",X"FE",X"FF",
		X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"0F",X"0F",X"01",X"00",X"88",X"0E",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"0F",X"0F",X"0F",X"8F",X"8F",X"CF",X"CF",
		X"F0",X"F0",X"E0",X"E0",X"E0",X"00",X"00",X"80",X"1F",X"1F",X"1F",X"1F",X"3F",X"3F",X"1F",X"C0",
		X"E1",X"E3",X"C7",X"87",X"81",X"80",X"C0",X"C0",X"FF",X"FE",X"F8",X"F3",X"F9",X"3C",X"03",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",X"E7",X"F3",X"F9",X"FC",X"FE",X"F0",X"F0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C0",X"CF",X"CF",X"CF",X"CF",X"CF",X"CF",X"CF",
		X"C0",X"C1",X"81",X"81",X"83",X"03",X"03",X"03",X"00",X"E0",X"F8",X"F8",X"F8",X"F0",X"F0",X"E0",
		X"01",X"84",X"07",X"07",X"07",X"01",X"00",X"06",X"E0",X"60",X"00",X"C0",X"81",X"80",X"21",X"E1",
		X"00",X"07",X"18",X"33",X"27",X"4F",X"5F",X"5F",X"00",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"00",X"FF",X"FF",X"C7",X"C3",X"01",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"08",X"0C",X"0E",X"0F",X"0F",
		X"00",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"7F",X"3F",X"1F",X"0F",X"07",X"01",X"80",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"0F",X"0F",X"CF",X"E7",X"F3",X"F8",X"C2",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C0",X"00",X"00",X"0E",X"0F",X"0F",X"0F",X"0F",
		X"C0",X"F0",X"F8",X"F8",X"F8",X"F8",X"F8",X"78",X"7F",X"3F",X"0E",X"04",X"00",X"03",X"03",X"03",
		X"18",X"08",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"07",X"07",X"07",X"07",X"0F",X"0E",X"08",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"03",X"01",X"02",X"00",X"00",X"00",X"78",X"FC",X"FE",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"F6",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"1A",
		X"0F",X"1F",X"1F",X"1F",X"3F",X"1D",X"03",X"01",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F9",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"73",X"07",X"06",X"00",X"00",X"00",X"00",X"00",
		X"EF",X"FB",X"FD",X"FC",X"FC",X"FC",X"F0",X"E0",X"F0",X"50",X"B0",X"E0",X"00",X"00",X"00",X"00",
		X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"40",X"F8",X"F0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"06",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"FC",X"70",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"10",X"00",X"00",X"00",X"00",
		X"04",X"00",X"11",X"00",X"08",X"00",X"00",X"40",X"01",X"10",X"00",X"00",X"24",X"00",X"00",X"82",
		X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",
		X"00",X"10",X"01",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"12",X"00",X"00",
		X"00",X"08",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"40",X"00",X"00",X"04",X"20",X"00",X"00",
		X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"20",X"00",X"01",X"00",X"00",
		X"00",X"81",X"00",X"10",X"00",X"00",X"80",X"00",X"10",X"00",X"00",X"00",X"90",X"00",X"00",X"10",
		X"01",X"10",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
