library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity obj4 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of obj4 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"13",X"13",X"21",X"20",X"20",X"41",X"41",X"80",X"08",X"1E",X"2F",X"2E",X"2E",X"4C",X"4F",
		X"80",X"00",X"10",X"26",X"2F",X"2C",X"40",X"48",X"80",X"00",X"10",X"20",X"20",X"20",X"40",X"40",
		X"40",X"40",X"40",X"80",X"80",X"81",X"83",X"83",X"46",X"42",X"44",X"8E",X"8E",X"8F",X"8E",X"88",
		X"44",X"40",X"40",X"8C",X"8F",X"86",X"80",X"80",X"40",X"40",X"40",X"80",X"80",X"80",X"80",X"80",
		X"E0",X"10",X"10",X"20",X"23",X"2F",X"47",X"41",X"E0",X"10",X"90",X"A0",X"6A",X"6F",X"6C",X"6F",
		X"E0",X"10",X"80",X"87",X"4E",X"48",X"20",X"2E",X"00",X"00",X"80",X"80",X"40",X"40",X"20",X"20",
		X"40",X"40",X"40",X"80",X"80",X"81",X"81",X"83",X"6F",X"61",X"60",X"93",X"9F",X"9E",X"9C",X"90",
		X"20",X"20",X"23",X"1F",X"18",X"10",X"10",X"10",X"20",X"20",X"20",X"1C",X"10",X"10",X"10",X"10",
		X"80",X"80",X"80",X"80",X"80",X"40",X"40",X"43",X"80",X"80",X"80",X"80",X"80",X"41",X"4E",X"4D",
		X"80",X"80",X"80",X"80",X"84",X"48",X"40",X"4E",X"80",X"80",X"80",X"80",X"80",X"40",X"40",X"40",
		X"47",X"48",X"20",X"20",X"20",X"10",X"11",X"00",X"4F",X"4B",X"20",X"23",X"23",X"16",X"08",X"80",
		X"42",X"40",X"23",X"2C",X"28",X"10",X"00",X"80",X"40",X"48",X"20",X"20",X"20",X"10",X"00",X"80",
		X"80",X"80",X"80",X"80",X"80",X"41",X"43",X"47",X"90",X"90",X"90",X"91",X"93",X"6E",X"6D",X"6F",
		X"10",X"10",X"18",X"18",X"10",X"20",X"2C",X"28",X"10",X"10",X"10",X"10",X"10",X"20",X"20",X"2C",
		X"4F",X"4D",X"21",X"20",X"20",X"10",X"10",X"E0",X"6F",X"6D",X"68",X"60",X"A5",X"91",X"13",X"E3",
		X"21",X"23",X"4E",X"4E",X"8E",X"8C",X"18",X"E0",X"28",X"20",X"40",X"40",X"80",X"80",X"00",X"00",
		X"00",X"10",X"10",X"20",X"20",X"20",X"43",X"47",X"80",X"00",X"16",X"2E",X"27",X"2A",X"4C",X"4C",
		X"80",X"00",X"10",X"20",X"20",X"24",X"44",X"46",X"80",X"00",X"10",X"20",X"20",X"24",X"46",X"4E",
		X"4F",X"4E",X"40",X"80",X"80",X"80",X"80",X"80",X"4F",X"48",X"40",X"81",X"80",X"80",X"80",X"80",
		X"4D",X"4A",X"4F",X"8F",X"8B",X"81",X"81",X"80",X"4C",X"44",X"48",X"8C",X"8C",X"8C",X"8C",X"88",
		X"E0",X"10",X"10",X"20",X"20",X"20",X"40",X"40",X"E0",X"10",X"94",X"A4",X"66",X"66",X"65",X"6C",
		X"E0",X"10",X"80",X"80",X"50",X"54",X"2C",X"25",X"00",X"00",X"80",X"84",X"44",X"4C",X"2C",X"38",
		X"40",X"41",X"43",X"83",X"87",X"84",X"80",X"80",X"6D",X"6C",X"68",X"98",X"90",X"90",X"90",X"90",
		X"25",X"2D",X"2F",X"3F",X"37",X"33",X"33",X"31",X"30",X"38",X"30",X"38",X"38",X"38",X"30",X"30",
		X"80",X"80",X"80",X"80",X"80",X"40",X"40",X"40",X"80",X"80",X"80",X"80",X"84",X"44",X"44",X"44",
		X"80",X"80",X"80",X"80",X"81",X"41",X"49",X"45",X"80",X"80",X"80",X"80",X"80",X"40",X"40",X"40",
		X"40",X"40",X"20",X"20",X"20",X"10",X"10",X"00",X"44",X"4D",X"2E",X"2E",X"2C",X"1C",X"08",X"88",
		X"45",X"4D",X"2F",X"27",X"27",X"11",X"00",X"80",X"40",X"48",X"28",X"28",X"28",X"18",X"08",X"88",
		X"80",X"80",X"80",X"80",X"81",X"41",X"41",X"40",X"90",X"90",X"90",X"90",X"90",X"69",X"68",X"6C",
		X"30",X"30",X"31",X"31",X"33",X"23",X"2D",X"25",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"38",
		X"40",X"40",X"20",X"20",X"20",X"10",X"10",X"E0",X"64",X"6D",X"67",X"6E",X"AE",X"9E",X"16",X"E4",
		X"2D",X"2F",X"53",X"53",X"80",X"80",X"10",X"E0",X"38",X"2C",X"4E",X"4E",X"87",X"81",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"86",X"07",X"00",X"00",X"00",X"00",X"00",X"02",X"03",X"05",
		X"00",X"00",X"06",X"07",X"0E",X"05",X"03",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0E",
		X"03",X"02",X"11",X"13",X"13",X"13",X"13",X"11",X"08",X"05",X"0E",X"0C",X"0C",X"08",X"08",X"00",
		X"0F",X"0F",X"06",X"00",X"00",X"00",X"00",X"00",X"0F",X"07",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"10",X"10",X"20",X"20",X"20",X"40",X"43",X"80",X"00",X"01",X"01",X"00",X"00",X"03",X"01",
		X"00",X"00",X"00",X"08",X"0C",X"07",X"0B",X"0F",X"00",X"00",X"00",X"00",X"00",X"08",X"0C",X"0E",
		X"41",X"40",X"40",X"80",X"80",X"80",X"80",X"80",X"08",X"0C",X"07",X"07",X"07",X"03",X"01",X"00",
		X"0F",X"0B",X"01",X"00",X"0A",X"08",X"0C",X"0C",X"0F",X"0B",X"08",X"00",X"00",X"00",X"00",X"00",
		X"10",X"10",X"10",X"10",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"01",X"00",X"07",
		X"00",X"00",X"00",X"00",X"00",X"08",X"07",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",
		X"00",X"81",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"0C",X"03",X"01",X"00",X"00",X"00",
		X"0F",X"0D",X"00",X"0C",X"0C",X"06",X"01",X"00",X"0E",X"01",X"00",X"00",X"00",X"00",X"08",X"00",
		X"80",X"80",X"80",X"80",X"80",X"40",X"40",X"40",X"00",X"00",X"00",X"0E",X"07",X"01",X"00",X"07",
		X"00",X"00",X"00",X"00",X"05",X"0F",X"03",X"0F",X"00",X"00",X"00",X"00",X"0C",X"0F",X"0E",X"08",
		X"40",X"40",X"20",X"23",X"20",X"10",X"10",X"00",X"00",X"00",X"0C",X"0F",X"01",X"00",X"00",X"80",
		X"0F",X"08",X"00",X"0C",X"0F",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"0C",
		X"00",X"00",X"00",X"0F",X"07",X"03",X"01",X"01",X"00",X"00",X"00",X"08",X"0E",X"0F",X"0C",X"1F",
		X"00",X"00",X"00",X"00",X"0F",X"8E",X"80",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"07",X"0F",X"00",X"00",X"16",X"12",X"14",X"2F",X"2E",X"28",X"20",X"20",
		X"04",X"00",X"00",X"0E",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"0F",X"01",X"01",X"00",X"00",X"00",X"00",X"0C",X"0F",X"0C",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"1F",X"17",X"10",X"10",X"10",X"86",X"82",X"0C",X"0F",X"0C",X"00",X"00",X"00",
		X"04",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"20",X"20",X"20",X"20",X"20",X"18",X"16",X"1F",
		X"00",X"01",X"03",X"01",X"07",X"01",X"05",X"00",X"00",X"0C",X"0F",X"0F",X"0A",X"01",X"08",X"09",
		X"0F",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"1E",X"0E",X"03",X"03",X"04",X"02",X"00",X"00",
		X"0B",X"83",X"8B",X"01",X"04",X"01",X"00",X"00",X"0D",X"0D",X"02",X"06",X"09",X"00",X"03",X"07",
		X"10",X"10",X"10",X"10",X"10",X"10",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"00",X"00",X"00",X"00",X"00",X"08",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"81",X"80",X"00",X"43",X"30",X"40",X"30",X"31",X"1F",X"18",X"06",X"2C",X"E1",
		X"00",X"80",X"FF",X"F0",X"F3",X"F6",X"F0",X"A8",X"10",X"70",X"FE",X"E0",X"EC",X"C0",X"A0",X"B0",
		X"00",X"40",X"00",X"80",X"80",X"01",X"00",X"00",X"00",X"01",X"04",X"10",X"18",X"3F",X"31",X"60",
		X"00",X"F8",X"F0",X"F6",X"F3",X"F0",X"8F",X"00",X"00",X"00",X"C0",X"E0",X"EC",X"F0",X"7E",X"10",
		X"00",X"00",X"10",X"03",X"01",X"80",X"81",X"00",X"00",X"03",X"F6",X"FC",X"30",X"1C",X"11",X"20",
		X"37",X"FC",X"F3",X"F4",X"F8",X"F0",X"E8",X"80",X"08",X"80",X"C8",X"E0",X"E0",X"30",X"80",X"10",
		X"70",X"00",X"00",X"40",X"00",X"40",X"20",X"00",X"C1",X"00",X"04",X"00",X"04",X"1F",X"10",X"10",
		X"08",X"F0",X"71",X"F1",X"F9",X"FF",X"C0",X"80",X"30",X"F0",X"FE",X"F1",X"FE",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"06",X"02",X"01",X"01",X"17",X"3C",X"78",X"F1",X"5C",X"1B",X"08",
		X"E8",X"F6",X"FC",X"F8",X"F0",X"D0",X"40",X"90",X"00",X"00",X"80",X"E0",X"40",X"00",X"00",X"F0",
		X"82",X"A0",X"30",X"00",X"10",X"00",X"10",X"00",X"61",X"80",X"06",X"00",X"02",X"01",X"02",X"80",
		X"79",X"73",X"70",X"70",X"FF",X"0A",X"00",X"00",X"F6",X"FC",X"F3",X"EC",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"02",X"07",X"03",X"06",X"1D",X"39",X"79",X"F0",X"94",X"19",
		X"68",X"F6",X"F8",X"E0",X"E0",X"C0",X"18",X"34",X"00",X"00",X"80",X"00",X"20",X"72",X"F2",X"E5",
		X"00",X"81",X"80",X"30",X"00",X"00",X"00",X"00",X"28",X"48",X"80",X"07",X"00",X"80",X"00",X"60",
		X"79",X"30",X"34",X"69",X"0B",X"0C",X"08",X"00",X"CD",X"83",X"06",X"0C",X"00",X"00",X"00",X"00",
		X"00",X"01",X"01",X"03",X"12",X"12",X"12",X"16",X"7C",X"FB",X"F6",X"F4",X"F6",X"F0",X"F1",X"0A",
		X"80",X"80",X"90",X"80",X"B0",X"10",X"70",X"BB",X"00",X"80",X"80",X"C0",X"E0",X"F5",X"FD",X"FA",
		X"07",X"00",X"00",X"80",X"50",X"00",X"00",X"00",X"08",X"18",X"10",X"23",X"67",X"60",X"00",X"30",
		X"78",X"10",X"3D",X"1B",X"06",X"06",X"00",X"00",X"E6",X"C4",X"8C",X"08",X"00",X"00",X"00",X"00",
		X"11",X"11",X"12",X"32",X"32",X"32",X"74",X"F6",X"F0",X"F0",X"E4",X"E8",X"EC",X"E4",X"E0",X"A2",
		X"A0",X"30",X"10",X"50",X"30",X"70",X"73",X"FA",X"00",X"80",X"C0",X"EB",X"FA",X"FA",X"EA",X"E4",
		X"E2",X"07",X"06",X"04",X"00",X"40",X"20",X"00",X"0A",X"08",X"18",X"1D",X"10",X"10",X"90",X"00",
		X"78",X"90",X"04",X"0D",X"03",X"01",X"00",X"60",X"C4",X"C4",X"CC",X"C0",X"40",X"00",X"00",X"00",
		X"E0",X"72",X"72",X"32",X"32",X"32",X"32",X"72",X"00",X"80",X"C8",X"C8",X"E8",X"EC",X"E4",X"E1",
		X"80",X"D0",X"30",X"F0",X"70",X"F1",X"71",X"F4",X"70",X"E2",X"EA",X"CA",X"CA",X"CA",X"C2",X"E2",
		X"73",X"E1",X"81",X"01",X"01",X"00",X"00",X"10",X"81",X"04",X"06",X"0B",X"01",X"01",X"20",X"80",
		X"14",X"C1",X"83",X"86",X"82",X"82",X"40",X"10",X"E6",X"64",X"14",X"0C",X"04",X"00",X"00",X"80",
		X"00",X"10",X"30",X"7A",X"FA",X"FA",X"7D",X"74",X"50",X"90",X"00",X"90",X"80",X"C0",X"E0",X"EA",
		X"F1",X"F2",X"72",X"F2",X"73",X"F6",X"70",X"D8",X"80",X"88",X"88",X"C8",X"CC",X"C4",X"E4",X"FC",
		X"34",X"36",X"33",X"31",X"21",X"01",X"00",X"00",X"E2",X"80",X"04",X"07",X"09",X"01",X"00",X"60",
		X"0A",X"43",X"42",X"46",X"42",X"22",X"92",X"00",X"74",X"04",X"0C",X"04",X"00",X"20",X"40",X"00",
		X"00",X"00",X"00",X"20",X"70",X"F4",X"F6",X"FB",X"10",X"70",X"10",X"30",X"10",X"90",X"C0",X"C0",
		X"E2",X"FA",X"FD",X"F5",X"FC",X"F4",X"F0",X"88",X"00",X"00",X"00",X"08",X"88",X"8C",X"88",X"8C",
		X"7C",X"34",X"16",X"03",X"00",X"00",X"00",X"00",X"EA",X"82",X"C4",X"83",X"08",X"0E",X"04",X"00",
		X"49",X"43",X"23",X"29",X"1D",X"65",X"00",X"C0",X"04",X"0A",X"00",X"10",X"A0",X"00",X"00",X"00",
		X"00",X"00",X"10",X"00",X"40",X"E4",X"F4",X"7A",X"61",X"F6",X"F1",X"70",X"70",X"30",X"81",X"C2",
		X"0C",X"06",X"8B",X"C9",X"E9",X"F0",X"92",X"89",X"00",X"00",X"00",X"00",X"08",X"08",X"04",X"0E",
		X"3B",X"1C",X"06",X"03",X"00",X"00",X"00",X"00",X"E9",X"C0",X"C0",X"68",X"0D",X"03",X"01",X"00",
		X"41",X"21",X"10",X"0E",X"03",X"10",X"00",X"60",X"00",X"18",X"18",X"C4",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"70",X"20",X"00",X"00",X"F0",X"76",X"F1",X"F6",X"F3",X"F1",X"B1",X"20",X"91",
		X"00",X"88",X"CE",X"E3",X"F3",X"A1",X"82",X"0B",X"00",X"00",X"00",X"00",X"00",X"0C",X"0C",X"00",
		X"F4",X"F6",X"FB",X"7C",X"07",X"01",X"00",X"00",X"E2",X"E9",X"E8",X"E0",X"F0",X"0F",X"01",X"00",
		X"61",X"10",X"00",X"0F",X"01",X"08",X"08",X"10",X"18",X"DC",X"C4",X"00",X"88",X"00",X"80",X"00",
		X"01",X"11",X"30",X"71",X"70",X"C0",X"10",X"80",X"C0",X"FE",X"F1",X"FE",X"F2",X"F3",X"70",X"11",
		X"00",X"00",X"FE",X"F2",X"C1",X"80",X"83",X"48",X"00",X"00",X"80",X"00",X"0C",X"18",X"10",X"0C",
		X"C0",X"F0",X"F2",X"F1",X"FC",X"13",X"00",X"00",X"00",X"F1",X"EC",X"F8",X"F0",X"FD",X"33",X"10",
		X"30",X"08",X"01",X"03",X"00",X"8E",X"87",X"80",X"E4",X"06",X"08",X"2E",X"00",X"20",X"40",X"00",
		X"00",X"00",X"01",X"80",X"80",X"00",X"43",X"30",X"00",X"70",X"3F",X"1C",X"18",X"06",X"2C",X"E1",
		X"00",X"10",X"FF",X"F0",X"F3",X"F6",X"F0",X"A8",X"70",X"F0",X"F0",X"E0",X"EC",X"C0",X"A0",X"B0",
		X"00",X"40",X"00",X"80",X"80",X"01",X"00",X"00",X"00",X"01",X"04",X"10",X"18",X"3F",X"71",X"00",
		X"00",X"F8",X"F0",X"F4",X"FF",X"F0",X"1F",X"00",X"00",X"00",X"C0",X"E0",X"E0",X"F0",X"FE",X"70",
		X"00",X"00",X"00",X"81",X"80",X"00",X"43",X"30",X"00",X"00",X"01",X"3F",X"18",X"06",X"2C",X"E1",
		X"00",X"10",X"FF",X"F0",X"FF",X"F4",X"F0",X"A8",X"00",X"E0",X"FE",X"F0",X"E0",X"E0",X"A0",X"B0",
		X"00",X"40",X"00",X"80",X"80",X"00",X"01",X"00",X"00",X"01",X"04",X"10",X"38",X"0C",X"0F",X"00",
		X"00",X"F8",X"F0",X"F6",X"F3",X"F0",X"1F",X"00",X"00",X"00",X"E0",X"E0",X"FC",X"F0",X"E0",X"00",
		X"00",X"00",X"00",X"80",X"80",X"00",X"40",X"30",X"00",X"00",X"00",X"10",X"30",X"00",X"20",X"E0",
		X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"A0",X"00",X"00",X"00",X"F0",X"F0",X"E0",X"A0",X"B0",
		X"00",X"40",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"10",X"00",X"00",X"00",
		X"00",X"F0",X"F0",X"F0",X"F1",X"0F",X"01",X"00",X"00",X"00",X"E0",X"FD",X"F7",X"0F",X"0E",X"0E",
		X"00",X"00",X"00",X"80",X"80",X"00",X"40",X"33",X"00",X"00",X"00",X"00",X"30",X"30",X"2C",X"EF",
		X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"A8",X"00",X"00",X"00",X"00",X"F0",X"F0",X"E0",X"BE",
		X"03",X"43",X"0F",X"8A",X"87",X"07",X"07",X"0B",X"0F",X"0F",X"36",X"30",X"09",X"06",X"02",X"0E",
		X"00",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"04",X"0E",X"E6",X"F2",X"F0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"20",X"40",X"40",X"20",X"B0",X"00",X"00",X"00",X"30",X"11",X"03",X"10",X"F1",
		X"00",X"00",X"13",X"3F",X"FE",X"F0",X"DC",X"53",X"00",X"00",X"C8",X"E0",X"E0",X"E0",X"40",X"40",
		X"63",X"A0",X"20",X"40",X"40",X"20",X"00",X"00",X"0F",X"00",X"00",X"01",X"00",X"00",X"00",X"00",
		X"AC",X"A3",X"5C",X"70",X"7E",X"33",X"10",X"00",X"80",X"80",X"40",X"E0",X"E0",X"E0",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"00",X"01",X"01",X"63",X"F3",X"06",X"07",X"11",
		X"04",X"3C",X"7C",X"78",X"F0",X"EF",X"D0",X"65",X"00",X"80",X"C0",X"C0",X"C0",X"C0",X"40",X"88",
		X"A0",X"60",X"10",X"51",X"20",X"20",X"00",X"00",X"21",X"07",X"0C",X"00",X"00",X"00",X"00",X"00",
		X"A9",X"86",X"70",X"33",X"00",X"00",X"00",X"00",X"80",X"70",X"FE",X"EC",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0C",X"0C",X"0E",X"1C",X"7F",X"FE",
		X"00",X"00",X"70",X"F0",X"F0",X"E8",X"F2",X"CA",X"00",X"00",X"80",X"80",X"80",X"E0",X"80",X"40",
		X"00",X"20",X"10",X"10",X"30",X"20",X"00",X"00",X"C9",X"01",X"03",X"02",X"84",X"C4",X"80",X"80",
		X"1A",X"44",X"33",X"30",X"00",X"00",X"00",X"00",X"5E",X"B8",X"E0",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"03",X"01",X"11",X"00",X"00",X"00",X"10",X"12",X"52",X"95",X"75",
		X"00",X"60",X"F0",X"F0",X"F8",X"E9",X"B5",X"E5",X"00",X"00",X"00",X"04",X"CC",X"0C",X"98",X"68",
		X"00",X"00",X"00",X"10",X"10",X"00",X"10",X"00",X"C9",X"81",X"81",X"81",X"81",X"C1",X"20",X"40",
		X"1B",X"52",X"20",X"00",X"00",X"00",X"00",X"00",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"20",X"10",X"71",X"F4",X"F5",
		X"00",X"72",X"63",X"F3",X"E7",X"D3",X"AF",X"E7",X"00",X"00",X"00",X"E0",X"80",X"40",X"00",X"80",
		X"07",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"E5",X"C2",X"0C",X"00",X"20",X"70",X"30",X"20",
		X"19",X"08",X"0C",X"04",X"02",X"82",X"00",X"80",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"11",X"02",X"73",X"B3",X"B1",X"F0",X"3F",X"C0",X"5A",
		X"00",X"28",X"78",X"FC",X"EC",X"F6",X"EE",X"88",X"00",X"00",X"80",X"00",X"C0",X"00",X"80",X"00",
		X"10",X"00",X"07",X"03",X"00",X"00",X"00",X"00",X"59",X"26",X"A0",X"2C",X"10",X"00",X"00",X"00",
		X"38",X"0E",X"03",X"00",X"00",X"80",X"E0",X"A0",X"80",X"00",X"00",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"11",X"10",X"10",X"10",X"00",X"10",X"00",X"60",X"FC",X"FF",X"F7",X"F0",X"73",X"9C",
		X"00",X"40",X"80",X"70",X"88",X"6C",X"80",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"83",X"8C",X"A3",X"A0",X"17",X"1C",X"10",X"00",
		X"0F",X"00",X"00",X"08",X"00",X"C0",X"30",X"80",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"20",X"20",X"30",X"00",X"00",X"30",X"33",X"B5",X"B0",X"90",X"CE",X"11",
		X"80",X"C0",X"BC",X"CF",X"AF",X"CF",X"B2",X"80",X"00",X"00",X"00",X"00",X"08",X"00",X"80",X"00",
		X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"D7",X"50",X"4E",X"20",X"00",X"05",X"03",X"00",
		X"0F",X"00",X"82",X"4F",X"1F",X"1E",X"18",X"00",X"08",X"00",X"00",X"08",X"C0",X"60",X"00",X"00",
		X"00",X"00",X"00",X"30",X"30",X"50",X"51",X"20",X"00",X"20",X"60",X"D3",X"E0",X"D8",X"F4",X"F2",
		X"00",X"00",X"8F",X"0F",X"C7",X"3F",X"44",X"00",X"00",X"00",X"0C",X"0C",X"08",X"00",X"00",X"00",
		X"20",X"10",X"11",X"00",X"00",X"00",X"00",X"00",X"3F",X"D0",X"54",X"A8",X"60",X"03",X"00",X"00",
		X"0F",X"00",X"04",X"0F",X"87",X"0F",X"0F",X"00",X"00",X"00",X"30",X"40",X"E8",X"88",X"0C",X"00",
		X"00",X"00",X"00",X"00",X"30",X"70",X"70",X"30",X"00",X"00",X"93",X"A5",X"80",X"D0",X"DE",X"F1",
		X"00",X"00",X"0C",X"0F",X"8F",X"2F",X"42",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",
		X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B7",X"20",X"6E",X"20",X"10",X"05",X"03",X"00",
		X"0F",X"00",X"02",X"0F",X"1F",X"0E",X"08",X"00",X"08",X"30",X"40",X"E8",X"40",X"00",X"00",X"00",
		X"00",X"00",X"01",X"10",X"10",X"30",X"70",X"70",X"F0",X"70",X"7C",X"5F",X"17",X"60",X"D3",X"FC",
		X"00",X"80",X"80",X"C0",X"48",X"4C",X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"20",
		X"70",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"F3",X"BC",X"13",X"00",X"07",X"0C",X"00",X"00",
		X"0F",X"00",X"80",X"F8",X"00",X"00",X"00",X"00",X"2C",X"70",X"C0",X"A0",X"80",X"00",X"00",X"00",
		X"00",X"10",X"30",X"10",X"00",X"10",X"60",X"20",X"00",X"C0",X"E3",X"E5",X"B0",X"20",X"4E",X"B1",
		X"00",X"00",X"0C",X"0F",X"0F",X"8F",X"82",X"00",X"00",X"00",X"00",X"00",X"08",X"10",X"20",X"40",
		X"60",X"F0",X"F0",X"70",X"00",X"00",X"00",X"00",X"E7",X"F0",X"FE",X"B0",X"10",X"05",X"03",X"00",
		X"8F",X"00",X"02",X"CF",X"EF",X"0E",X"08",X"00",X"78",X"40",X"60",X"48",X"40",X"00",X"00",X"00",
		X"00",X"00",X"00",X"20",X"40",X"40",X"20",X"B0",X"00",X"00",X"01",X"37",X"1F",X"07",X"12",X"F0",
		X"00",X"00",X"0E",X"0D",X"B8",X"F8",X"D3",X"54",X"00",X"00",X"00",X"00",X"C0",X"E0",X"48",X"40",
		X"60",X"A0",X"20",X"40",X"40",X"20",X"00",X"00",X"0F",X"00",X"02",X"0F",X"07",X"03",X"00",X"00",
		X"AF",X"A0",X"53",X"78",X"38",X"0D",X"0E",X"00",X"80",X"80",X"48",X"E0",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"20",X"40",X"40",X"20",X"B0",X"00",X"00",X"00",X"30",X"10",X"01",X"10",X"F0",
		X"00",X"00",X"01",X"07",X"8F",X"F8",X"F6",X"59",X"00",X"00",X"0C",X"08",X"00",X"E0",X"E0",X"C8",
		X"61",X"A0",X"20",X"40",X"40",X"20",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"BE",X"B1",X"76",X"78",X"07",X"01",X"00",X"00",X"C0",X"C8",X"E0",X"E0",X"00",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"10",X"10",X"10",X"00",
		X"00",X"00",X"00",X"38",X"00",X"F0",X"E0",X"00",X"08",X"04",X"04",X"E3",X"60",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",
		X"02",X"00",X"00",X"00",X"04",X"06",X"00",X"79",X"02",X"04",X"00",X"00",X"01",X"03",X"0F",X"EF",
		X"00",X"00",X"04",X"06",X"00",X"08",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"8D",X"74",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"E3",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"40",X"20",X"11",X"00",X"02",X"07",X"0F",X"0F",X"07",X"13",X"F3",
		X"00",X"60",X"F0",X"F0",X"F8",X"78",X"69",X"57",X"00",X"00",X"C0",X"C0",X"80",X"00",X"00",X"4C",
		X"00",X"21",X"40",X"00",X"02",X"00",X"00",X"00",X"00",X"03",X"03",X"07",X"0F",X"0F",X"07",X"02",
		X"0F",X"67",X"79",X"F8",X"F8",X"F0",X"60",X"00",X"0F",X"0C",X"00",X"80",X"C0",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"05",X"00",X"10",X"00",X"08",X"0E",X"1E",X"1F",X"1F",X"03",X"03",
		X"00",X"00",X"C0",X"F0",X"F0",X"F3",X"77",X"67",X"00",X"00",X"00",X"80",X"80",X"40",X"0E",X"0C",
		X"71",X"00",X"11",X"10",X"20",X"01",X"00",X"00",X"00",X"01",X"01",X"83",X"07",X"07",X"03",X"00",
		X"1F",X"18",X"3C",X"7C",X"3C",X"0C",X"08",X"08",X"08",X"E0",X"E0",X"C0",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"03",X"03",X"03",X"14",X"00",X"00",X"00",X"18",X"1E",X"1F",X"9F",X"0F",
		X"00",X"00",X"F0",X"F0",X"F2",X"F3",X"67",X"47",X"00",X"00",X"80",X"80",X"0A",X"8C",X"0C",X"48",
		X"10",X"11",X"70",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"41",X"09",X"81",X"83",X"05",X"00",
		X"1E",X"1C",X"3C",X"1E",X"0E",X"0E",X"0E",X"02",X"E8",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"07",X"07",X"07",X"00",X"00",X"00",X"00",X"10",X"1C",X"6C",X"8E",
		X"00",X"00",X"20",X"E3",X"FF",X"E7",X"EF",X"5D",X"00",X"00",X"04",X"88",X"08",X"08",X"C0",X"80",
		X"11",X"18",X"11",X"20",X"10",X"00",X"00",X"00",X"06",X"01",X"01",X"00",X"85",X"80",X"00",X"02",
		X"10",X"38",X"0E",X"0E",X"0F",X"0F",X"0F",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"07",X"00",X"00",X"00",X"00",X"01",X"10",X"1E",X"6F",
		X"00",X"01",X"22",X"E6",X"CE",X"CE",X"8E",X"4C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"02",X"04",X"00",X"00",X"00",X"00",X"00",X"CE",X"8A",X"80",X"88",X"42",X"80",X"00",X"00",
		X"0E",X"47",X"0F",X"07",X"07",X"07",X"04",X"00",X"00",X"00",X"08",X"0C",X"0C",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"01",X"11",X"3B",X"4F",
		X"04",X"04",X"4E",X"CE",X"EE",X"EE",X"EC",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"03",X"03",X"00",X"02",X"00",X"00",X"00",X"4E",X"CA",X"C0",X"40",X"65",X"10",X"20",X"00",
		X"0F",X"0F",X"07",X"03",X"03",X"00",X"02",X"00",X"08",X"0C",X"0C",X"0E",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"01",X"13",X"01",X"11",X"0E",
		X"08",X"08",X"2C",X"6C",X"6E",X"FC",X"FC",X"6B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",
		X"03",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"2F",X"4F",X"4C",X"68",X"31",X"08",X"00",X"00",
		X"07",X"07",X"01",X"00",X"04",X"80",X"40",X"00",X"0E",X"0F",X"0E",X"0C",X"00",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"33",X"33",X"17",X"17",X"13",X"03",
		X"00",X"00",X"00",X"88",X"88",X"C8",X"CB",X"CF",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0F",
		X"00",X"03",X"03",X"07",X"00",X"00",X"00",X"00",X"2F",X"6F",X"6C",X"3C",X"1C",X"00",X"04",X"00",
		X"07",X"01",X"00",X"00",X"CA",X"40",X"20",X"00",X"0E",X"0E",X"0C",X"00",X"04",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"08",X"06",X"0F",X"C7",X"FF",X"73",X"70",
		X"00",X"00",X"00",X"08",X"00",X"09",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"0F",X"0E",X"0E",
		X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"07",X"4F",X"4F",X"3F",X"1E",X"0E",X"01",X"00",
		X"0B",X"08",X"00",X"11",X"E4",X"20",X"00",X"00",X"0E",X"04",X"02",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"11",X"01",X"31",X"30",X"10",X"00",X"00",X"20",X"3C",X"9F",X"EE",X"FF",X"EB",
		X"00",X"00",X"00",X"00",X"80",X"03",X"03",X"07",X"00",X"00",X"00",X"00",X"0E",X"0E",X"0E",X"0E",
		X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"E1",X"27",X"17",X"0F",X"0F",X"0F",X"00",
		X"06",X"08",X"08",X"00",X"EA",X"10",X"00",X"04",X"08",X"01",X"08",X"C0",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"04",X"03",X"01",X"31",X"70",X"00",X"00",X"F0",X"70",X"3E",X"0E",X"BF",X"EF",
		X"00",X"00",X"01",X"83",X"87",X"0F",X"0F",X"8A",X"00",X"00",X"08",X"0C",X"0C",X"0C",X"0E",X"00",
		X"30",X"30",X"10",X"00",X"00",X"00",X"00",X"00",X"F9",X"C3",X"83",X"13",X"07",X"07",X"03",X"00",
		X"20",X"0C",X"08",X"0D",X"E8",X"0C",X"02",X"00",X"20",X"48",X"00",X"80",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"00",X"03",X"2F",X"03",X"00",X"00",X"70",X"F0",X"F0",X"3C",X"0F",X"8F",
		X"00",X"01",X"07",X"8F",X"8F",X"0F",X"06",X"0C",X"00",X"00",X"00",X"00",X"08",X"0A",X"00",X"20",
		X"00",X"10",X"30",X"10",X"00",X"00",X"00",X"00",X"6F",X"E3",X"F3",X"F3",X"F1",X"61",X"01",X"00",
		X"C0",X"8C",X"08",X"0C",X"0E",X"0E",X"08",X"00",X"48",X"00",X"88",X"40",X"00",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"40",X"20",X"11",X"00",X"02",X"07",X"0F",X"0F",X"07",X"13",X"F3",
		X"00",X"00",X"F0",X"F0",X"F8",X"78",X"78",X"51",X"00",X"00",X"00",X"80",X"80",X"80",X"00",X"4C",
		X"00",X"21",X"40",X"00",X"02",X"00",X"00",X"00",X"00",X"03",X"03",X"07",X"0F",X"0F",X"07",X"02",
		X"0F",X"71",X"78",X"F8",X"F8",X"F0",X"00",X"00",X"0F",X"0C",X"80",X"80",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"40",X"20",X"11",X"00",X"02",X"07",X"0F",X"0F",X"07",X"13",X"F3",
		X"00",X"00",X"00",X"01",X"3A",X"7C",X"78",X"50",X"00",X"00",X"00",X"0C",X"C0",X"E0",X"C0",X"4C",
		X"00",X"21",X"40",X"00",X"02",X"00",X"00",X"00",X"00",X"03",X"03",X"07",X"0F",X"0F",X"07",X"02",
		X"0F",X"70",X"78",X"3C",X"0A",X"01",X"00",X"00",X"0F",X"CC",X"E0",X"C0",X"00",X"0C",X"00",X"00",
		X"00",X"90",X"60",X"90",X"02",X"00",X"00",X"01",X"00",X"02",X"07",X"0F",X"0F",X"07",X"03",X"03",
		X"00",X"00",X"00",X"01",X"0A",X"0C",X"08",X"00",X"00",X"60",X"90",X"6C",X"00",X"00",X"00",X"00",
		X"00",X"01",X"00",X"00",X"02",X"90",X"60",X"90",X"00",X"03",X"03",X"07",X"0F",X"0F",X"07",X"02",
		X"03",X"00",X"08",X"0C",X"0A",X"01",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"6C",X"90",X"60",
		X"00",X"60",X"90",X"60",X"02",X"00",X"00",X"01",X"00",X"02",X"07",X"0F",X"0F",X"07",X"03",X"03",
		X"00",X"00",X"00",X"01",X"0A",X"0C",X"08",X"00",X"00",X"90",X"60",X"9C",X"00",X"00",X"00",X"00",
		X"00",X"01",X"00",X"00",X"02",X"60",X"90",X"60",X"00",X"03",X"03",X"07",X"0F",X"0F",X"07",X"02",
		X"00",X"00",X"08",X"0C",X"0A",X"01",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"9C",X"60",X"90",
		X"00",X"00",X"00",X"00",X"02",X"40",X"30",X"10",X"00",X"00",X"07",X"0C",X"00",X"00",X"10",X"FF",
		X"00",X"0F",X"39",X"30",X"33",X"63",X"7E",X"58",X"00",X"00",X"8E",X"8C",X"0C",X"08",X"00",X"40",
		X"13",X"30",X"40",X"00",X"00",X"00",X"00",X"00",X"FC",X"1F",X"03",X"01",X"08",X"04",X"04",X"00",
		X"50",X"38",X"2E",X"3F",X"07",X"01",X"00",X"00",X"40",X"00",X"00",X"08",X"8C",X"0C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"04",X"00",X"70",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"10",
		X"00",X"0C",X"27",X"31",X"63",X"37",X"3E",X"3C",X"00",X"00",X"0C",X"08",X"00",X"00",X"40",X"40",
		X"10",X"13",X"10",X"20",X"01",X"00",X"00",X"00",X"3F",X"FD",X"E8",X"00",X"00",X"06",X"08",X"00",
		X"5E",X"DF",X"1F",X"00",X"00",X"00",X"04",X"00",X"00",X"8E",X"CF",X"C2",X"00",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"10",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",
		X"00",X"00",X"40",X"60",X"E0",X"40",X"13",X"4C",X"00",X"00",X"00",X"00",X"86",X"48",X"00",X"80",
		X"16",X"10",X"31",X"00",X"00",X"10",X"00",X"00",X"07",X"1E",X"FE",X"F0",X"81",X"00",X"02",X"00",
		X"30",X"80",X"80",X"00",X"08",X"04",X"00",X"00",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"04",X"00",X"04",X"00",X"05",X"00",X"00",X"00",X"01",X"61",X"E1",
		X"04",X"0C",X"0C",X"5C",X"4C",X"6C",X"7B",X"0F",X"00",X"00",X"00",X"00",X"80",X"00",X"0E",X"8C",
		X"10",X"10",X"10",X"00",X"10",X"00",X"00",X"00",X"85",X"8F",X"87",X"FA",X"D0",X"00",X"00",X"00",
		X"6F",X"8C",X"C0",X"80",X"00",X"0C",X"0A",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"02",X"00",X"06",X"06",X"06",X"06",X"06",X"06",X"66",
		X"00",X"00",X"00",X"30",X"40",X"50",X"51",X"63",X"00",X"00",X"00",X"00",X"00",X"04",X"8F",X"0F",
		X"06",X"04",X"04",X"04",X"00",X"00",X"00",X"00",X"F6",X"C6",X"C7",X"C7",X"74",X"00",X"00",X"00",
		X"0E",X"48",X"00",X"00",X"80",X"01",X"04",X"00",X"01",X"02",X"02",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"02",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"16",X"06",X"17",X"33",X"43",
		X"00",X"00",X"C0",X"01",X"E3",X"86",X"4E",X"08",X"00",X"00",X"04",X"0C",X"0C",X"04",X"00",X"00",
		X"00",X"02",X"06",X"00",X"00",X"00",X"00",X"00",X"73",X"F3",X"E3",X"77",X"72",X"12",X"00",X"00",
		X"88",X"00",X"08",X"00",X"80",X"01",X"00",X"00",X"00",X"00",X"04",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"11",X"01",X"31",X"01",X"31",X"01",
		X"00",X"00",X"84",X"06",X"E2",X"63",X"C1",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",
		X"00",X"01",X"03",X"00",X"00",X"00",X"00",X"00",X"71",X"71",X"73",X"73",X"31",X"09",X"00",X"00",
		X"C0",X"80",X"88",X"88",X"C0",X"82",X"00",X"00",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"01",X"00",X"04",X"04",X"00",X"00",X"30",X"00",X"6C",X"1E",X"3F",X"07",
		X"02",X"07",X"05",X"04",X"84",X"0C",X"4C",X"0C",X"00",X"00",X"00",X"08",X"04",X"04",X"02",X"02",
		X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"33",X"71",X"70",X"38",X"18",X"08",X"04",X"00",
		X"8C",X"08",X"8C",X"EE",X"C4",X"44",X"00",X"00",X"00",X"00",X"00",X"02",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"07",X"07",X"00",X"00",X"00",X"C0",X"50",X"70",X"08",X"6C",
		X"03",X"05",X"06",X"84",X"04",X"04",X"84",X"24",X"00",X"08",X"0C",X"04",X"02",X"02",X"00",X"00",
		X"01",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"1F",X"73",X"71",X"30",X"14",X"0A",X"02",X"00",
		X"04",X"16",X"1E",X"FE",X"E2",X"00",X"00",X"00",X"00",X"02",X"02",X"02",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"10",X"07",X"03",X"02",X"03",X"03",X"93",X"23",X"73",X"ED",X"0F",
		X"00",X"0A",X"00",X"80",X"00",X"88",X"28",X"78",X"00",X"00",X"00",X"00",X"04",X"02",X"00",X"02",
		X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"0F",X"33",X"30",X"10",X"00",X"03",X"05",X"00",
		X"1A",X"1F",X"1E",X"F5",X"E0",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"16",X"21",X"00",X"10",X"00",X"00",X"60",X"20",X"50",X"50",X"DC",X"C3",
		X"00",X"00",X"00",X"02",X"00",X"00",X"60",X"F0",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"80",
		X"30",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"01",X"02",X"00",X"00",
		X"1E",X"17",X"17",X"30",X"08",X"00",X"04",X"00",X"A6",X"C0",X"08",X"80",X"80",X"00",X"00",X"00",
		X"00",X"00",X"03",X"01",X"00",X"00",X"20",X"20",X"00",X"23",X"CE",X"C8",X"6C",X"AE",X"A7",X"A3",
		X"00",X"00",X"02",X"00",X"00",X"00",X"C0",X"F0",X"00",X"00",X"00",X"00",X"04",X"02",X"00",X"A0",
		X"00",X"17",X"3F",X"34",X"00",X"01",X"00",X"00",X"87",X"8F",X"0F",X"00",X"00",X"00",X"02",X"00",
		X"BF",X"0B",X"11",X"00",X"00",X"06",X"01",X"00",X"C0",X"8C",X"80",X"40",X"48",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"00",X"42",X"30",X"10",X"00",X"00",X"04",X"00",X"00",X"00",X"10",X"FC",
		X"00",X"00",X"06",X"01",X"30",X"31",X"77",X"5E",X"00",X"00",X"00",X"88",X"CE",X"8C",X"08",X"40",
		X"13",X"30",X"40",X"02",X"00",X"01",X"00",X"00",X"FF",X"1D",X"00",X"00",X"08",X"04",X"04",X"00",
		X"5C",X"3E",X"3F",X"03",X"00",X"00",X"02",X"00",X"40",X"00",X"88",X"8C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"40",X"42",X"30",X"10",X"00",X"00",X"00",X"07",X"00",X"00",X"10",X"FC",
		X"00",X"00",X"00",X"08",X"0E",X"03",X"30",X"50",X"00",X"00",X"00",X"00",X"00",X"08",X"8C",X"40",
		X"13",X"30",X"40",X"42",X"00",X"00",X"00",X"00",X"FF",X"1C",X"00",X"00",X"06",X"04",X"00",X"00",
		X"5F",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"4E",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"04",X"08",X"C0",
		X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"1C",X"0C",X"0D",X"00",X"01",X"00",X"00",X"00",
		X"80",X"74",X"00",X"01",X"00",X"08",X"06",X"00",X"18",X"C9",X"01",X"07",X"07",X"0F",X"0F",X"0F",
		X"08",X"0C",X"0E",X"01",X"00",X"00",X"00",X"0F",X"00",X"00",X"01",X"01",X"75",X"82",X"88",X"8C",
		X"00",X"06",X"0F",X"0E",X"EC",X"10",X"10",X"18",X"00",X"00",X"08",X"00",X"00",X"04",X"06",X"02",
		X"0F",X"0F",X"0D",X"0F",X"0F",X"0F",X"0F",X"0F",X"8F",X"8E",X"8E",X"7F",X"0F",X"0E",X"0E",X"0F",
		X"1C",X"1D",X"1E",X"E6",X"06",X"00",X"0C",X"0C",X"00",X"02",X"08",X"04",X"00",X"00",X"01",X"04",
		X"00",X"00",X"00",X"03",X"00",X"21",X"13",X"12",X"00",X"00",X"06",X"01",X"0E",X"0F",X"13",X"F1",
		X"00",X"00",X"31",X"33",X"30",X"60",X"78",X"5C",X"00",X"00",X"8E",X"80",X"00",X"00",X"00",X"40",
		X"12",X"13",X"21",X"00",X"03",X"00",X"00",X"00",X"F9",X"13",X"0F",X"0E",X"01",X"06",X"00",X"00",
		X"FC",X"B8",X"24",X"30",X"03",X"01",X"00",X"00",X"C0",X"00",X"00",X"00",X"80",X"0E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"05",X"01",X"31",X"00",X"00",X"00",X"0E",X"00",X"0E",X"0F",X"33",
		X"00",X"00",X"50",X"B0",X"70",X"70",X"58",X"78",X"00",X"0C",X"00",X"80",X"08",X"0E",X"4E",X"CC",
		X"32",X"12",X"11",X"10",X"00",X"00",X"00",X"00",X"F9",X"C1",X"8B",X"8F",X"06",X"0C",X"01",X"00",
		X"B8",X"B8",X"08",X"02",X"08",X"08",X"00",X"00",X"04",X"E0",X"60",X"01",X"02",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"00",X"02",X"05",X"11",X"00",X"00",X"00",X"08",X"04",X"0C",X"0E",X"3F",
		X"02",X"00",X"00",X"41",X"31",X"63",X"B3",X"F3",X"00",X"00",X"00",X"0C",X"8E",X"8E",X"8C",X"8C",
		X"33",X"12",X"03",X"01",X"00",X"00",X"00",X"00",X"F1",X"C1",X"85",X"8F",X"87",X"02",X"06",X"00",
		X"88",X"88",X"0A",X"08",X"02",X"04",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"01",X"00",X"00",X"10",X"10",X"10",X"08",X"2F",X"3F",
		X"00",X"C0",X"C0",X"D3",X"F3",X"B1",X"F0",X"F8",X"00",X"00",X"00",X"08",X"88",X"88",X"C0",X"C0",
		X"07",X"01",X"31",X"01",X"00",X"00",X"00",X"00",X"39",X"74",X"E0",X"C9",X"4F",X"41",X"01",X"00",
		X"CC",X"CD",X"0C",X"0E",X"0A",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"04",X"04",X"44",X"E8",X"F4",X"70",X"30",X"01",X"2F",
		X"00",X"00",X"00",X"30",X"E0",X"60",X"F8",X"CC",X"00",X"00",X"00",X"00",X"00",X"01",X"E2",X"F6",
		X"01",X"03",X"05",X"10",X"00",X"00",X"00",X"00",X"3F",X"38",X"78",X"EA",X"3D",X"13",X"10",X"00",
		X"CE",X"8C",X"0D",X"0D",X"0D",X"04",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"03",X"08",X"60",X"61",X"20",X"30",X"38",X"00",X"37",
		X"00",X"06",X"CE",X"8F",X"F0",X"B0",X"F0",X"0C",X"00",X"00",X"02",X"82",X"C0",X"80",X"40",X"80",
		X"04",X"01",X"03",X"02",X"00",X"00",X"00",X"00",X"1F",X"1C",X"38",X"FD",X"F4",X"13",X"00",X"00",
		X"8C",X"8E",X"06",X"06",X"8E",X"81",X"02",X"00",X"00",X"08",X"08",X"08",X"00",X"00",X"00",X"00",
		X"00",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"13",X"37",X"33",X"31",X"10",X"38",
		X"00",X"08",X"8C",X"4E",X"CC",X"48",X"80",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",
		X"03",X"02",X"00",X"00",X"01",X"01",X"00",X"00",X"33",X"1E",X"1C",X"1D",X"36",X"43",X"00",X"00",
		X"CC",X"87",X"83",X"83",X"C6",X"2C",X"00",X"00",X"08",X"04",X"04",X"08",X"08",X"00",X"00",X"00",
		X"00",X"00",X"04",X"14",X"30",X"10",X"20",X"10",X"00",X"06",X"37",X"1F",X"F0",X"D0",X"F0",X"03",
		X"01",X"60",X"68",X"40",X"C0",X"C1",X"00",X"CE",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"0C",
		X"00",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"13",X"17",X"06",X"06",X"17",X"18",X"04",X"00",
		X"8F",X"83",X"C1",X"FB",X"F2",X"8C",X"00",X"00",X"02",X"08",X"0C",X"04",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"08",X"74",X"F6",X"00",X"00",X"00",X"C0",X"70",X"60",X"F1",X"33",
		X"02",X"22",X"71",X"F2",X"E0",X"C0",X"08",X"4F",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"37",X"13",X"0B",X"0B",X"0B",X"02",X"02",X"00",
		X"CF",X"C1",X"E1",X"75",X"CB",X"8C",X"80",X"00",X"08",X"0C",X"0A",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"11",X"01",X"70",X"70",X"00",X"00",X"30",X"FC",X"FC",X"F8",X"B0",X"F1",
		X"00",X"00",X"00",X"00",X"00",X"01",X"CF",X"CF",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"08",
		X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"93",X"3B",X"03",X"07",X"05",X"04",X"00",X"00",
		X"C9",X"E2",X"70",X"39",X"2F",X"28",X"08",X"00",X"0E",X"08",X"C8",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"17",X"17",X"13",X"13",X"04",X"00",X"00",X"28",X"C8",X"6C",X"DC",X"FC",
		X"00",X"00",X"00",X"01",X"02",X"03",X"07",X"CF",X"00",X"00",X"00",X"08",X"00",X"04",X"0A",X"88",
		X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"05",X"01",X"04",X"02",X"00",X"00",
		X"F8",X"38",X"1A",X"1F",X"1E",X"04",X"06",X"00",X"CC",X"84",X"0C",X"08",X"00",X"00",X"00",X"00",
		X"00",X"03",X"00",X"10",X"01",X"07",X"27",X"33",X"00",X"00",X"A0",X"D0",X"E0",X"E0",X"A1",X"E1",
		X"00",X"00",X"00",X"07",X"00",X"07",X"0F",X"CC",X"00",X"00",X"00",X"00",X"04",X"0A",X"08",X"C8",
		X"02",X"70",X"60",X"08",X"04",X"00",X"00",X"00",X"D1",X"D1",X"01",X"04",X"01",X"01",X"00",X"00",
		X"F9",X"38",X"1D",X"1F",X"06",X"03",X"08",X"00",X"C4",X"84",X"88",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"00",X"21",X"13",X"12",X"00",X"00",X"06",X"01",X"0E",X"0F",X"13",X"F9",
		X"00",X"00",X"00",X"00",X"30",X"30",X"78",X"58",X"00",X"00",X"06",X"80",X"C0",X"80",X"04",X"4E",
		X"12",X"13",X"21",X"00",X"03",X"00",X"00",X"00",X"F1",X"13",X"0F",X"0E",X"01",X"06",X"00",X"00",
		X"F8",X"B8",X"34",X"00",X"00",X"00",X"00",X"00",X"CE",X"04",X"80",X"80",X"00",X"06",X"00",X"00",
		X"00",X"00",X"00",X"03",X"00",X"21",X"13",X"12",X"00",X"00",X"06",X"01",X"0E",X"0E",X"12",X"F1",
		X"00",X"00",X"00",X"00",X"00",X"00",X"31",X"53",X"00",X"00",X"06",X"00",X"00",X"08",X"8C",X"4E",
		X"12",X"13",X"21",X"00",X"03",X"00",X"00",X"00",X"F9",X"12",X"0E",X"0E",X"01",X"06",X"00",X"00",
		X"F3",X"31",X"00",X"04",X"00",X"00",X"00",X"00",X"CE",X"8C",X"08",X"00",X"00",X"06",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"04",X"02",X"04",X"06",X"16",X"32",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"CE",X"0F",X"07",X"01",X"01",X"00",X"00",X"00",X"00",
		X"00",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"30",X"18",X"0C",X"0C",X"00",X"00",X"00",X"00",
		X"CE",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"05",X"0A",X"07",X"00",X"00",X"00",X"10",X"0D",X"0A",X"09",X"17",X"2C",X"48",X"80",X"00",
		X"08",X"08",X"0C",X"8B",X"43",X"20",X"10",X"00",X"00",X"02",X"04",X"00",X"00",X"00",X"00",X"80",
		X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"20",X"11",X"07",X"03",X"00",
		X"00",X"10",X"20",X"4E",X"8F",X"0F",X"0E",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"00",X"60",X"60",X"F4",X"00",X"00",X"00",X"08",X"05",X"05",X"07",X"C3",
		X"00",X"00",X"00",X"08",X"01",X"02",X"0E",X"7F",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"88",
		X"00",X"E4",X"60",X"60",X"00",X"01",X"00",X"00",X"C1",X"03",X"07",X"05",X"05",X"08",X"00",X"00",
		X"2F",X"0F",X"0E",X"02",X"01",X"08",X"00",X"00",X"7C",X"88",X"00",X"00",X"0C",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"01",X"0F",X"0F",X"01",
		X"00",X"00",X"00",X"0B",X"07",X"0F",X"3F",X"4C",X"00",X"00",X"00",X"0C",X"08",X"0C",X"F8",X"00",
		X"70",X"C4",X"20",X"72",X"30",X"00",X"00",X"00",X"E0",X"41",X"01",X"03",X"02",X"02",X"04",X"00",
		X"03",X"0F",X"0F",X"0C",X"04",X"02",X"00",X"00",X"8E",X"0F",X"0E",X"0C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"01",X"03",X"03",X"07",X"07",X"07",X"0F",X"0F",X"0E",
		X"08",X"00",X"07",X"0C",X"1C",X"7C",X"C0",X"40",X"00",X"00",X"00",X"00",X"60",X"C0",X"00",X"02",
		X"60",X"70",X"24",X"50",X"32",X"10",X"00",X"00",X"60",X"61",X"01",X"81",X"83",X"C1",X"02",X"04",
		X"07",X"0F",X"0F",X"0F",X"0F",X"01",X"00",X"00",X"0C",X"0C",X"08",X"0E",X"0E",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"05",X"00",X"00",X"01",X"05",X"07",X"07",X"07",X"0F",
		X"00",X"0E",X"0F",X"2E",X"7E",X"4D",X"43",X"03",X"00",X"00",X"40",X"80",X"04",X"8E",X"0E",X"0E",
		X"00",X"00",X"70",X"32",X"20",X"10",X"00",X"00",X"40",X"E0",X"40",X"00",X"C0",X"C8",X"40",X"00",
		X"0F",X"0F",X"0F",X"08",X"08",X"04",X"08",X"00",X"0C",X"00",X"08",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"02",X"0B",X"05",X"07",X"03",
		X"00",X"10",X"30",X"23",X"37",X"2F",X"EF",X"4F",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"0C",
		X"03",X"04",X"20",X"30",X"30",X"10",X"00",X"00",X"0F",X"30",X"30",X"80",X"A0",X"78",X"B2",X"00",
		X"0E",X"0F",X"06",X"06",X"02",X"01",X"02",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"01",X"07",X"07",X"17",X"03",X"07",X"0F",X"07",
		X"40",X"40",X"49",X"4B",X"4B",X"4B",X"87",X"07",X"00",X"00",X"04",X"0C",X"0C",X"0C",X"00",X"04",
		X"00",X"01",X"02",X"02",X"10",X"10",X"00",X"00",X"0F",X"1C",X"30",X"10",X"90",X"D0",X"B5",X"20",
		X"07",X"07",X"02",X"03",X"00",X"80",X"80",X"00",X"08",X"00",X"00",X"00",X"08",X"08",X"00",X"00",
		X"00",X"04",X"06",X"07",X"03",X"03",X"01",X"00",X"04",X"0C",X"0E",X"1E",X"0E",X"0F",X"0F",X"0F",
		X"81",X"81",X"83",X"43",X"43",X"C7",X"4F",X"07",X"00",X"09",X"0B",X"0F",X"0E",X"0E",X"0C",X"08",
		X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"06",X"0C",X"00",X"00",X"00",X"71",X"70",X"10",
		X"03",X"01",X"C0",X"C0",X"40",X"74",X"70",X"40",X"00",X"08",X"04",X"04",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"01",X"01",X"01",X"00",X"01",X"20",X"20",X"2C",X"2E",X"2E",X"2E",X"1F",X"07",
		X"04",X"0E",X"0F",X"8F",X"0E",X"0F",X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"02",X"06",X"04",X"08",X"18",X"10",X"00",
		X"07",X"81",X"C0",X"80",X"90",X"B1",X"D4",X"40",X"00",X"0C",X"02",X"00",X"80",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"01",X"00",X"00",X"80",X"C0",X"67",X"17",X"17",X"17",X"0F",
		X"00",X"04",X"04",X"04",X"0C",X"8F",X"0E",X"0F",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"0C",
		X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"0B",X"03",X"03",X"04",X"04",X"02",X"00",
		X"0F",X"68",X"60",X"10",X"50",X"E0",X"D2",X"00",X"0A",X"01",X"40",X"C0",X"C8",X"80",X"00",X"00",
		X"00",X"00",X"20",X"10",X"02",X"17",X"07",X"07",X"00",X"07",X"0F",X"47",X"E7",X"2B",X"2C",X"0C",
		X"00",X"00",X"08",X"0A",X"0E",X"0E",X"0E",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0A",
		X"03",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"01",X"01",X"02",X"01",X"00",
		X"20",X"70",X"20",X"00",X"30",X"31",X"20",X"00",X"00",X"00",X"E0",X"C4",X"40",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"60",X"30",X"00",X"00",X"01",X"01",X"01",X"0F",X"87",X"E7",X"33",X"20",
		X"08",X"08",X"0C",X"0C",X"0E",X"0E",X"0E",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"08",
		X"07",X"07",X"03",X"03",X"0F",X"07",X"00",X"00",X"08",X"0E",X"0F",X"0F",X"0F",X"0C",X"00",X"00",
		X"66",X"60",X"08",X"18",X"18",X"3C",X"08",X"04",X"60",X"E0",X"40",X"A2",X"C0",X"84",X"00",X"00",
		X"00",X"00",X"03",X"01",X"03",X"01",X"F0",X"07",X"00",X"00",X"0D",X"0E",X"0F",X"0F",X"C3",X"2C",
		X"00",X"00",X"00",X"08",X"0D",X"0F",X"08",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"60",
		X"1F",X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"03",X"02",X"04",X"00",X"00",X"00",
		X"78",X"28",X"0C",X"0C",X"04",X"02",X"00",X"00",X"E2",X"30",X"42",X"E0",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"00",X"60",X"60",X"F4",X"00",X"00",X"00",X"08",X"04",X"07",X"03",X"C1",
		X"00",X"00",X"00",X"04",X"0B",X"0F",X"0F",X"7F",X"00",X"00",X"00",X"00",X"0E",X"0C",X"0C",X"88",
		X"00",X"E4",X"60",X"60",X"00",X"01",X"00",X"00",X"C0",X"01",X"83",X"07",X"04",X"08",X"00",X"00",
		X"20",X"0F",X"0F",X"0F",X"0B",X"04",X"00",X"00",X"70",X"88",X"0C",X"0C",X"0E",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"00",X"60",X"60",X"F4",X"00",X"00",X"00",X"08",X"05",X"07",X"03",X"C3",
		X"00",X"01",X"07",X"0F",X"0F",X"0F",X"0F",X"70",X"00",X"0C",X"08",X"00",X"0C",X"0E",X"08",X"80",
		X"00",X"E4",X"60",X"60",X"00",X"01",X"00",X"00",X"C0",X"03",X"83",X"07",X"05",X"08",X"00",X"00",
		X"20",X"00",X"0F",X"0F",X"0F",X"0F",X"07",X"01",X"70",X"80",X"08",X"0E",X"0C",X"00",X"08",X"0C",
		X"00",X"00",X"04",X"06",X"06",X"63",X"61",X"F0",X"00",X"01",X"00",X"00",X"00",X"04",X"02",X"C0",
		X"00",X"01",X"00",X"09",X"02",X"09",X"00",X"71",X"00",X"00",X"01",X"08",X"01",X"02",X"01",X"80",
		X"00",X"E0",X"60",X"60",X"00",X"00",X"00",X"00",X"C0",X"00",X"01",X"08",X"00",X"00",X"00",X"00",
		X"28",X"09",X"05",X"09",X"08",X"08",X"00",X"00",X"77",X"8F",X"07",X"07",X"0B",X"0F",X"0F",X"07",
		X"00",X"00",X"00",X"00",X"02",X"69",X"6A",X"F5",X"00",X"00",X"00",X"00",X"00",X"02",X"04",X"C3",
		X"00",X"00",X"00",X"00",X"00",X"04",X"08",X"72",X"00",X"00",X"00",X"00",X"0C",X"0C",X"03",X"87",
		X"00",X"EE",X"6E",X"6E",X"0F",X"0F",X"0F",X"0F",X"CE",X"08",X"0C",X"08",X"0A",X"08",X"08",X"08",
		X"2C",X"00",X"04",X"0A",X"04",X"02",X"0C",X"0C",X"77",X"83",X"01",X"01",X"00",X"00",X"00",X"00",
		X"00",X"60",X"30",X"10",X"00",X"21",X"23",X"12",X"00",X"00",X"C2",X"FA",X"77",X"1B",X"13",X"01",
		X"00",X"00",X"10",X"EF",X"CF",X"9F",X"0F",X"7F",X"00",X"00",X"00",X"00",X"C8",X"08",X"08",X"80",
		X"00",X"12",X"23",X"21",X"00",X"10",X"30",X"60",X"04",X"01",X"13",X"1B",X"77",X"FA",X"C2",X"00",
		X"D0",X"0F",X"0F",X"9F",X"CF",X"EF",X"10",X"00",X"E0",X"80",X"08",X"08",X"C8",X"00",X"00",X"00",
		X"00",X"00",X"00",X"F0",X"71",X"00",X"01",X"23",X"00",X"00",X"01",X"F7",X"F7",X"FF",X"13",X"01",
		X"00",X"6E",X"4F",X"9F",X"AF",X"0E",X"7E",X"7C",X"00",X"00",X"00",X"80",X"00",X"00",X"E0",X"80",
		X"12",X"00",X"00",X"11",X"10",X"00",X"00",X"00",X"00",X"04",X"81",X"19",X"1F",X"33",X"72",X"E0",
		X"80",X"0F",X"8F",X"EF",X"FF",X"EF",X"0F",X"00",X"80",X"00",X"A8",X"4C",X"8C",X"4C",X"08",X"00",
		X"00",X"00",X"00",X"01",X"30",X"F3",X"60",X"01",X"00",X"07",X"1F",X"3F",X"FF",X"EF",X"E7",X"07",
		X"00",X"80",X"28",X"4C",X"4C",X"3C",X"FC",X"C0",X"00",X"00",X"00",X"00",X"00",X"C0",X"80",X"80",
		X"43",X"32",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"84",X"8F",X"81",X"11",X"30",
		X"87",X"0F",X"CF",X"FF",X"FF",X"E7",X"87",X"80",X"00",X"E8",X"0C",X"EC",X"8C",X"0C",X"08",X"00",
		X"00",X"00",X"00",X"00",X"00",X"72",X"F1",X"C7",X"00",X"27",X"2F",X"6F",X"EF",X"EF",X"4F",X"0F",
		X"00",X"80",X"88",X"A8",X"78",X"F8",X"C8",X"87",X"00",X"00",X"00",X"80",X"00",X"80",X"00",X"EC",
		X"01",X"23",X"13",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"80",X"40",X"47",X"26",X"00",X"00",
		X"0F",X"3F",X"7F",X"3F",X"6C",X"6A",X"E8",X"C0",X"0E",X"EE",X"8E",X"0C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"33",X"70",X"00",X"90",X"A3",X"D7",X"CF",X"CF",X"CF",X"6F",
		X"00",X"00",X"18",X"6C",X"FC",X"E9",X"AB",X"87",X"00",X"00",X"00",X"00",X"00",X"2C",X"CE",X"0E",
		X"F3",X"C0",X"01",X"31",X"00",X"00",X"00",X"00",X"07",X"08",X"09",X"88",X"28",X"13",X"10",X"00",
		X"07",X"77",X"17",X"33",X"32",X"3A",X"30",X"30",X"FE",X"CC",X"8C",X"80",X"08",X"80",X"00",X"00",
		X"00",X"00",X"01",X"13",X"03",X"03",X"13",X"13",X"00",X"20",X"4C",X"2E",X"8F",X"CF",X"CF",X"EF",
		X"00",X"20",X"60",X"E0",X"E0",X"63",X"27",X"87",X"00",X"00",X"00",X"40",X"4E",X"8F",X"1F",X"EF",
		X"31",X"73",X"60",X"E0",X"80",X"00",X"00",X"00",X"8E",X"88",X"09",X"0C",X"C4",X"00",X"00",X"00",
		X"17",X"33",X"11",X"11",X"86",X"4C",X"40",X"00",X"CE",X"CC",X"CC",X"C0",X"C8",X"C0",X"C0",X"40",
		X"00",X"00",X"00",X"00",X"20",X"13",X"17",X"17",X"00",X"00",X"80",X"90",X"4C",X"0E",X"8F",X"CF",
		X"00",X"80",X"80",X"C0",X"D1",X"43",X"C7",X"97",X"00",X"00",X"80",X"80",X"28",X"4E",X"CF",X"CF",
		X"17",X"13",X"30",X"31",X"30",X"60",X"40",X"00",X"EF",X"8E",X"88",X"04",X"16",X"63",X"00",X"00",
		X"37",X"03",X"08",X"01",X"43",X"36",X"00",X"00",X"CF",X"CE",X"E8",X"64",X"60",X"30",X"10",X"00",
		X"00",X"00",X"00",X"10",X"13",X"47",X"67",X"17",X"00",X"20",X"20",X"30",X"38",X"8E",X"2F",X"8F",
		X"00",X"20",X"11",X"A3",X"87",X"97",X"97",X"B7",X"00",X"00",X"4C",X"8E",X"8E",X"CE",X"CE",X"CE",
		X"13",X"11",X"11",X"10",X"10",X"10",X"10",X"10",X"EF",X"CE",X"CC",X"C4",X"8B",X"91",X"80",X"00",
		X"13",X"00",X"04",X"21",X"91",X"08",X"00",X"00",X"EC",X"7E",X"38",X"18",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"23",X"17",X"47",X"00",X"00",X"41",X"73",X"73",X"19",X"8D",X"1E",
		X"00",X"50",X"5C",X"5E",X"1F",X"9F",X"BF",X"BF",X"00",X"00",X"00",X"80",X"80",X"C0",X"CC",X"F0",
		X"37",X"13",X"03",X"00",X"01",X"00",X"00",X"00",X"8E",X"EE",X"EE",X"EC",X"C4",X"E5",X"60",X"40",
		X"0E",X"01",X"09",X"11",X"41",X"4C",X"80",X"00",X"3C",X"10",X"08",X"C8",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"73",X"00",X"10",X"11",X"51",X"E1",X"71",X"31",X"3E",
		X"00",X"4E",X"4F",X"6F",X"7F",X"7F",X"2F",X"0F",X"00",X"00",X"00",X"00",X"00",X"E4",X"F8",X"3E",
		X"07",X"77",X"17",X"03",X"00",X"00",X"00",X"00",X"0F",X"CF",X"EF",X"CF",X"63",X"65",X"71",X"30",
		X"00",X"04",X"10",X"20",X"2E",X"46",X"00",X"00",X"08",X"4C",X"8C",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"20",X"10",X"00",X"00",X"00",X"40",X"21",X"23",X"83",X"E3",X"73",X"30",
		X"80",X"8E",X"CF",X"FF",X"7F",X"5F",X"4E",X"0E",X"00",X"00",X"00",X"48",X"F0",X"FC",X"00",X"08",
		X"50",X"21",X"13",X"73",X"03",X"03",X"01",X"00",X"0E",X"1F",X"FF",X"EF",X"7F",X"3E",X"1E",X"00",
		X"00",X"04",X"00",X"12",X"9F",X"98",X"C8",X"C0",X"6C",X"84",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"00",X"00",X"70",X"00",X"00",X"20",X"17",X"9F",X"5F",X"0F",X"E7",X"E7",X"73",
		X"00",X"00",X"F8",X"FE",X"FE",X"4F",X"0C",X"08",X"00",X"00",X"F0",X"E0",X"08",X"00",X"68",X"8C",
		X"00",X"50",X"21",X"03",X"13",X"03",X"01",X"00",X"00",X"1F",X"7F",X"FF",X"3F",X"0F",X"0F",X"00",
		X"00",X"02",X"08",X"C9",X"CF",X"FC",X"74",X"10",X"04",X"00",X"80",X"88",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"70",X"31",X"23",X"12",X"00",X"00",X"02",X"0B",X"E7",X"FB",X"33",X"01",
		X"00",X"00",X"0F",X"0F",X"3F",X"FF",X"EE",X"7C",X"00",X"00",X"00",X"08",X"C8",X"00",X"00",X"80",
		X"00",X"12",X"23",X"31",X"70",X"00",X"00",X"00",X"04",X"01",X"33",X"FB",X"E7",X"0B",X"02",X"00",
		X"D0",X"0C",X"EE",X"FF",X"3F",X"0F",X"0F",X"00",X"E0",X"80",X"00",X"00",X"C8",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"71",X"33",X"12",X"00",X"01",X"03",X"0B",X"07",X"FB",X"F3",X"31",
		X"00",X"0C",X"0E",X"0E",X"0F",X"9F",X"FE",X"FC",X"00",X"00",X"00",X"00",X"00",X"C0",X"80",X"80",
		X"00",X"12",X"33",X"71",X"00",X"00",X"00",X"00",X"04",X"31",X"F3",X"FB",X"07",X"0B",X"03",X"01",
		X"D0",X"FC",X"FE",X"9F",X"0F",X"0E",X"0E",X"0C",X"E0",X"80",X"80",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"01",X"00",X"00",X"01",X"03",X"74",X"08",
		X"01",X"01",X"38",X"08",X"08",X"0A",X"07",X"07",X"07",X"E8",X"0E",X"81",X"00",X"00",X"0B",X"09",
		X"60",X"10",X"00",X"00",X"04",X"02",X"00",X"00",X"10",X"00",X"61",X"00",X"70",X"00",X"00",X"00",
		X"06",X"0C",X"00",X"00",X"C0",X"00",X"30",X"00",X"80",X"00",X"01",X"01",X"00",X"E1",X"07",X"80",
		X"0D",X"0A",X"01",X"0C",X"00",X"00",X"00",X"01",X"0E",X"0A",X"05",X"08",X"00",X"01",X"33",X"82",
		X"04",X"01",X"02",X"30",X"00",X"00",X"06",X"0C",X"00",X"00",X"C0",X"00",X"80",X"00",X"00",X"00",
		X"30",X"0B",X"06",X"09",X"05",X"0E",X"0F",X"0E",X"19",X"80",X"28",X"30",X"00",X"08",X"00",X"00",
		X"1E",X"02",X"02",X"81",X"00",X"31",X"03",X"07",X"00",X"00",X"00",X"00",X"C0",X"0C",X"8C",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
