library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity tron_sp_bits_1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of tron_sp_bits_1 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",
		X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"22",X"00",X"00",X"77",X"22",
		X"00",X"66",X"77",X"00",X"00",X"66",X"77",X"00",X"00",X"66",X"77",X"00",X"00",X"00",X"77",X"00",
		X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"66",X"00",
		X"00",X"02",X"66",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"00",X"00",
		X"00",X"00",X"00",X"62",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",
		X"00",X"22",X"77",X"00",X"00",X"22",X"77",X"00",X"00",X"66",X"66",X"00",X"00",X"66",X"27",X"00",
		X"72",X"66",X"22",X"77",X"72",X"66",X"22",X"67",X"00",X"22",X"77",X"22",X"00",X"22",X"77",X"26",
		X"20",X"66",X"77",X"66",X"20",X"66",X"77",X"66",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",
		X"00",X"66",X"22",X"66",X"00",X"66",X"22",X"26",X"00",X"22",X"77",X"22",X"00",X"22",X"77",X"22",
		X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"00",X"00",
		X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"20",X"00",X"22",X"00",X"00",X"00",X"22",
		X"00",X"22",X"77",X"00",X"00",X"22",X"77",X"00",X"00",X"66",X"66",X"00",X"00",X"66",X"27",X"00",
		X"72",X"66",X"22",X"77",X"72",X"66",X"22",X"67",X"00",X"22",X"77",X"22",X"00",X"22",X"77",X"26",
		X"20",X"66",X"77",X"66",X"20",X"66",X"77",X"66",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",
		X"00",X"66",X"22",X"66",X"00",X"66",X"22",X"26",X"00",X"22",X"77",X"22",X"00",X"22",X"77",X"22",
		X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",
		X"00",X"77",X"00",X"00",X"00",X"77",X"CC",X"00",X"00",X"22",X"77",X"77",X"00",X"22",X"77",X"77",
		X"CC",X"77",X"22",X"22",X"CC",X"77",X"22",X"72",X"CC",X"77",X"22",X"22",X"CC",X"77",X"22",X"77",
		X"67",X"77",X"22",X"77",X"67",X"77",X"22",X"77",X"CC",X"22",X"27",X"77",X"CC",X"22",X"77",X"77",
		X"00",X"22",X"27",X"22",X"00",X"22",X"27",X"22",X"00",X"22",X"77",X"77",X"00",X"22",X"77",X"77",
		X"00",X"77",X"22",X"CC",X"00",X"77",X"22",X"00",X"CC",X"77",X"22",X"77",X"CC",X"77",X"22",X"77",
		X"CC",X"77",X"77",X"22",X"CC",X"77",X"77",X"22",X"00",X"22",X"CC",X"77",X"00",X"22",X"CC",X"77",
		X"00",X"77",X"CC",X"CC",X"00",X"77",X"CC",X"CC",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"AA",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",
		X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"AA",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"BC",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BC",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"00",X"00",X"00",X"BC",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BC",X"00",X"00",X"00",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"01",X"00",X"22",X"01",X"11",X"00",X"C1",X"11",
		X"1D",X"10",X"1A",X"13",X"1D",X"10",X"00",X"33",X"1D",X"10",X"00",X"33",X"1D",X"11",X"A1",X"33",
		X"1D",X"1D",X"DD",X"33",X"1D",X"1D",X"AD",X"33",X"1D",X"1D",X"DD",X"33",X"1D",X"1D",X"DD",X"33",
		X"1D",X"1D",X"DD",X"33",X"1D",X"1D",X"DD",X"33",X"1D",X"1D",X"DD",X"33",X"1D",X"1D",X"D2",X"33",
		X"1D",X"1D",X"22",X"33",X"1D",X"1D",X"2D",X"33",X"1D",X"1D",X"3D",X"23",X"1D",X"1D",X"33",X"23",
		X"1D",X"1D",X"33",X"23",X"1D",X"1D",X"3D",X"23",X"1D",X"1D",X"2D",X"33",X"1D",X"1D",X"22",X"33",
		X"1D",X"1D",X"D2",X"33",X"1D",X"1D",X"DD",X"33",X"1D",X"11",X"11",X"33",X"1D",X"10",X"00",X"13",
		X"11",X"00",X"00",X"11",X"01",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"11",X"11",X"00",X"DD",X"DD",X"DD",X"01",X"33",X"33",X"33",X"11",X"11",X"11",X"11",
		X"11",X"22",X"A2",X"2A",X"01",X"11",X"11",X"11",X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",
		X"00",X"11",X"12",X"11",X"00",X"DD",X"22",X"DD",X"00",X"DD",X"2D",X"2D",X"00",X"DD",X"3D",X"2D",
		X"00",X"DD",X"33",X"2D",X"00",X"DD",X"3D",X"2D",X"00",X"DD",X"2D",X"2D",X"02",X"DD",X"22",X"DD",
		X"22",X"12",X"12",X"AD",X"A3",X"33",X"33",X"1A",X"A3",X"33",X"33",X"32",X"22",X"12",X"12",X"1D",
		X"02",X"DD",X"DD",X"AD",X"00",X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",X"11",X"11",X"11",
		X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",X"01",X"11",X"11",X"11",X"11",X"22",X"A2",X"2A",
		X"11",X"11",X"11",X"11",X"01",X"33",X"33",X"33",X"00",X"DD",X"DD",X"DD",X"00",X"11",X"11",X"11",
		X"00",X"00",X"00",X"05",X"05",X"00",X"00",X"05",X"55",X"00",X"00",X"55",X"C2",X"00",X"00",X"5C",
		X"CC",X"50",X"00",X"5C",X"C2",X"50",X"00",X"C6",X"55",X"50",X"02",X"CA",X"55",X"50",X"5C",X"C6",
		X"C2",X"50",X"7C",X"C6",X"CC",X"52",X"C7",X"C6",X"C2",X"52",X"7C",X"C6",X"55",X"52",X"7C",X"CA",
		X"55",X"52",X"C7",X"C6",X"C2",X"52",X"77",X"C6",X"CC",X"CC",X"55",X"C6",X"C2",X"C7",X"55",X"C6",
		X"55",X"C7",X"55",X"CA",X"55",X"C7",X"55",X"C6",X"C2",X"C7",X"55",X"C6",X"CC",X"C7",X"55",X"C6",
		X"C2",X"C7",X"55",X"C6",X"55",X"C7",X"55",X"CA",X"55",X"C7",X"55",X"C6",X"C2",X"CC",X"55",X"C6",
		X"CC",X"57",X"77",X"C6",X"C2",X"55",X"CC",X"C6",X"55",X"50",X"22",X"CA",X"55",X"50",X"22",X"CC",
		X"05",X"00",X"77",X"5C",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",
		X"00",X"52",X"25",X"2C",X"00",X"52",X"25",X"2C",X"05",X"CC",X"55",X"CC",X"55",X"55",X"5A",X"55",
		X"56",X"CC",X"CC",X"C6",X"5C",X"CC",X"CC",X"CC",X"55",X"66",X"6A",X"66",X"00",X"CC",X"CC",X"CC",
		X"00",X"55",X"CC",X"C5",X"00",X"00",X"77",X"C7",X"00",X"00",X"77",X"CC",X"00",X"05",X"75",X"77",
		X"00",X"05",X"55",X"77",X"00",X"55",X"55",X"57",X"00",X"CC",X"55",X"57",X"00",X"57",X"55",X"57",
		X"00",X"57",X"55",X"57",X"00",X"CC",X"55",X"57",X"00",X"55",X"55",X"57",X"00",X"05",X"55",X"77",
		X"00",X"05",X"75",X"77",X"00",X"00",X"77",X"CC",X"00",X"00",X"77",X"C7",X"00",X"55",X"CC",X"C5",
		X"00",X"CC",X"CC",X"CC",X"55",X"66",X"6A",X"66",X"5C",X"CC",X"CC",X"CC",X"56",X"CC",X"CC",X"C6",
		X"55",X"55",X"5A",X"55",X"05",X"CC",X"55",X"CC",X"00",X"52",X"25",X"2C",X"00",X"5C",X"C5",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"3F",X"00",X"00",X"00",X"33",X"00",
		X"00",X"0F",X"93",X"00",X"00",X"55",X"59",X"00",X"00",X"55",X"55",X"99",X"00",X"55",X"55",X"99",
		X"00",X"0F",X"AA",X"90",X"00",X"FF",X"AA",X"00",X"00",X"F3",X"AA",X"F0",X"00",X"33",X"A5",X"3F",
		X"00",X"55",X"F5",X"55",X"00",X"39",X"99",X"3F",X"00",X"F3",X"9A",X"F0",X"00",X"FF",X"9A",X"00",
		X"00",X"0F",X"9A",X"50",X"00",X"99",X"55",X"55",X"00",X"99",X"55",X"55",X"00",X"99",X"55",X"00",
		X"00",X"0F",X"93",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"3F",X"00",X"00",X"03",X"F0",X"00",
		X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"05",X"20",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"23",X"00",
		X"00",X"00",X"23",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"32",X"00",
		X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"EE",X"22",X"00",X"00",X"BE",X"22",X"00",X"00",X"BB",X"22",
		X"22",X"22",X"22",X"00",X"00",X"00",X"2E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",
		X"00",X"00",X"32",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"00",X"02",X"00",X"22",X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",
		X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"02",X"00",X"00",
		X"00",X"00",X"20",X"00",X"00",X"00",X"E2",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"7E",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"E2",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"20",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",
		X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"23",X"00",X"00",X"02",X"22",X"00",X"00",X"72",X"02",
		X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"A6",X"33",X"00",X"00",X"A6",X"3B",
		X"00",X"00",X"A6",X"AA",X"00",X"00",X"A7",X"3A",X"00",X"00",X"AA",X"3A",X"00",X"00",X"0A",X"AA",
		X"00",X"00",X"00",X"3B",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",
		X"00",X"00",X"72",X"02",X"00",X"00",X"02",X"22",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"02",X"00",X"00",X"22",X"22",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"00",X"00",X"D0",X"20",X"00",X"00",X"D0",X"00",X"00",X"00",X"D0",X"00",X"00",
		X"00",X"DD",X"70",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"DD",X"70",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"02",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"22",X"22",X"00",X"00",X"00",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"C7",
		X"00",X"00",X"00",X"C7",X"00",X"00",X"00",X"C7",X"00",X"00",X"00",X"C7",X"00",X"00",X"00",X"C0",
		X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"70",
		X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"F7",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"CC",
		X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"7C",X"00",X"00",X"00",X"7C",
		X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",
		X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"CC",
		X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"7C",X"00",X"00",X"00",X"7C",
		X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"20",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"07",X"00",
		X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"CC",
		X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"7C",X"00",X"00",X"00",X"7C",
		X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"C0",X"00",
		X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"07",X"00",
		X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"CC",
		X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"7C",X"00",X"00",X"00",X"7C",
		X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",
		X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"7F",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F7",X"00",X"00",X"00",X"CC",
		X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"7C",X"00",X"00",X"00",X"7C",
		X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"20",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"77",X"00",X"00",
		X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F7",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"7F",X"00",X"00",X"0F",X"CC",
		X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"7C",X"00",X"00",X"00",X"7C",
		X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"2C",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"77",X"00",X"00",
		X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F7",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"7F",X"00",X"00",X"0F",X"CC",
		X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"7C",X"00",X"00",X"00",X"7C",
		X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"00",X"00",
		X"00",X"70",X"00",X"00",X"00",X"77",X"00",X"FF",X"00",X"07",X"FF",X"FF",X"00",X"00",X"FF",X"CC",
		X"00",X"00",X"FF",X"77",X"00",X"00",X"FF",X"CC",X"00",X"00",X"0F",X"7C",X"00",X"00",X"00",X"7C",
		X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"2C",X"00",X"00",X"FF",X"2C",X"77",X"00",X"FF",
		X"00",X"77",X"FF",X"CC",X"00",X"07",X"FF",X"77",X"00",X"00",X"FF",X"CC",X"00",X"00",X"FF",X"7C",
		X"00",X"00",X"00",X"7C",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",
		X"00",X"00",X"00",X"F7",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F7",
		X"00",X"00",X"00",X"CF",X"00",X"00",X"00",X"7C",X"00",X"00",X"FF",X"C7",X"02",X"77",X"FF",X"C7",
		X"02",X"77",X"FF",X"C7",X"00",X"00",X"FF",X"C7",X"00",X"00",X"00",X"7C",X"00",X"00",X"00",X"CF",
		X"00",X"00",X"00",X"F7",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"33",X"00",X"EE",X"33",X"99",X"00",X"EE",X"EE",X"99",
		X"33",X"E9",X"EE",X"99",X"3E",X"99",X"EE",X"EE",X"9E",X"99",X"9E",X"99",X"99",X"9E",X"9E",X"E9",
		X"99",X"9E",X"EE",X"33",X"9E",X"E9",X"EE",X"EE",X"33",X"EE",X"E3",X"99",X"00",X"EE",X"30",X"99",
		X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"33",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"EE",X"00",X"00",X"99",X"99",X"30",X"00",X"9E",X"93",X"30",X"00",
		X"EE",X"3E",X"30",X"00",X"33",X"E9",X"30",X"00",X"EE",X"33",X"30",X"00",X"33",X"00",X"30",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"33",X"00",X"EE",X"33",X"99",X"00",X"EE",X"EE",X"99",
		X"33",X"E9",X"EE",X"EE",X"3E",X"99",X"EE",X"99",X"9E",X"99",X"9E",X"99",X"99",X"9E",X"9E",X"E9",
		X"99",X"9E",X"EE",X"33",X"3E",X"E9",X"EE",X"99",X"03",X"EE",X"E3",X"EE",X"00",X"EE",X"30",X"99",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"39",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"33",X"00",X"00",X"33",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",
		X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",
		X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"93",X"00",X"00",X"00",
		X"EE",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"EE",X"33",X"00",X"00",X"33",X"EE",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"03",X"00",X"00",
		X"00",X"03",X"00",X"00",X"00",X"39",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0E",X"00",X"00",X"00",X"9E",X"00",
		X"00",X"00",X"EE",X"99",X"00",X"00",X"EE",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"99",X"99",
		X"00",X"44",X"EE",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"99",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"E0",X"00",X"00",X"04",X"00",X"00",X"00",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E9",
		X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"E4",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E9",
		X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"E9",
		X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E9",
		X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"E9",
		X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"9E",
		X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"EE",
		X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"44",X"00",
		X"00",X"99",X"94",X"00",X"00",X"9E",X"94",X"00",X"00",X"9E",X"44",X"00",X"00",X"9E",X"00",X"00",
		X"00",X"9E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E4",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"CC",X"CC",X"EE",
		X"0E",X"EE",X"EE",X"CC",X"EE",X"CC",X"CC",X"CC",X"EE",X"CC",X"CC",X"CF",X"EE",X"CC",X"CC",X"CF",
		X"EE",X"CC",X"CC",X"CF",X"EE",X"CC",X"CC",X"CF",X"1E",X"CC",X"CC",X"CC",X"0E",X"EE",X"EE",X"CC",
		X"00",X"CC",X"CC",X"EE",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"09",X"99",X"00",X"00",X"09",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"09",X"CC",X"00",
		X"00",X"0F",X"CC",X"00",X"00",X"09",X"CC",X"00",X"00",X"09",X"CC",X"00",X"00",X"0E",X"CC",X"00",
		X"00",X"0E",X"CC",X"00",X"00",X"0E",X"CC",X"00",X"00",X"0E",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"CC",X"CC",X"77",
		X"07",X"77",X"77",X"CC",X"77",X"CC",X"CC",X"CC",X"77",X"CC",X"CC",X"CF",X"77",X"CC",X"CC",X"CF",
		X"77",X"CC",X"CC",X"CF",X"77",X"CC",X"CC",X"CF",X"77",X"CC",X"CC",X"CC",X"07",X"77",X"77",X"CC",
		X"00",X"CC",X"CC",X"77",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"0F",X"FF",X"00",X"00",X"0F",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"0F",X"CC",X"00",
		X"00",X"0F",X"CC",X"00",X"00",X"04",X"CC",X"00",X"00",X"04",X"CC",X"00",X"00",X"07",X"CC",X"00",
		X"00",X"07",X"CC",X"00",X"00",X"07",X"CC",X"00",X"00",X"07",X"CC",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",
		X"00",X"31",X"31",X"31",X"00",X"13",X"13",X"13",X"00",X"31",X"31",X"31",X"00",X"11",X"11",X"11",
		X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",
		X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",
		X"00",X"11",X"11",X"11",X"01",X"11",X"11",X"11",X"01",X"11",X"11",X"11",X"11",X"11",X"11",X"10",
		X"FF",X"FF",X"FF",X"F0",X"FF",X"FF",X"FF",X"00",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"53",X"53",X"53",X"00",X"35",X"35",X"35",X"00",X"53",X"53",X"53",X"00",X"35",X"35",X"35",
		X"00",X"53",X"53",X"53",X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",
		X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",
		X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",
		X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"33",
		X"00",X"13",X"13",X"13",X"00",X"31",X"31",X"31",X"03",X"13",X"13",X"13",X"01",X"31",X"31",X"31",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"B5",X"B5",X"B5",X"00",X"5B",X"5B",X"5B",X"00",X"B5",X"B5",X"B5",X"00",X"5B",X"5B",X"5B",
		X"00",X"B5",X"B5",X"B5",X"00",X"5B",X"5B",X"5B",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",
		X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",
		X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",
		X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",
		X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",
		X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"35",X"35",X"35",
		X"00",X"53",X"53",X"53",X"00",X"35",X"35",X"35",X"00",X"53",X"53",X"53",X"00",X"35",X"35",X"35",
		X"00",X"DB",X"DB",X"DB",X"00",X"BD",X"BD",X"BD",X"00",X"DB",X"DB",X"DB",X"00",X"BD",X"BD",X"BD",
		X"00",X"DB",X"DB",X"DB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",
		X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",
		X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",
		X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",
		X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",
		X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"B5",X"B5",X"B5",X"00",X"5B",X"5B",X"5B",
		X"00",X"B5",X"B5",X"B5",X"00",X"5B",X"5B",X"5B",X"00",X"B5",X"B5",X"B5",X"00",X"5B",X"5B",X"5B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DF",X"DF",X"DF",X"D0",X"FD",X"FD",X"FD",X"F0",X"0F",X"DF",X"DF",X"DF",X"0D",X"FD",X"FD",X"FD",
		X"00",X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",
		X"00",X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",
		X"00",X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",
		X"00",X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",X"DD",X"DD",X"DD",X"00",X"BD",X"BD",X"BD",
		X"00",X"DB",X"DB",X"DB",X"00",X"BD",X"BD",X"BD",X"00",X"DB",X"DB",X"DB",X"00",X"BD",X"BD",X"BD",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"10",
		X"FF",X"FF",X"FF",X"F0",X"0F",X"FF",X"FF",X"FF",X"0F",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",
		X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",
		X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",
		X"00",X"FF",X"FF",X"FF",X"00",X"DF",X"DF",X"DF",X"00",X"FD",X"FD",X"FD",X"00",X"DF",X"DF",X"DF",
		X"60",X"66",X"66",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"60",X"55",X"55",X"65",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"60",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"50",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"54",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"04",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"04",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"40",X"40",
		X"60",X"66",X"66",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"65",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"54",X"55",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"65",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"50",X"50",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"54",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"44",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"FA",X"00",
		X"00",X"00",X"0B",X"00",X"00",X"00",X"50",X"00",X"00",X"0A",X"AF",X"7F",X"00",X"A0",X"A0",X"00",
		X"0A",X"00",X"07",X"0F",X"A5",X"00",X"70",X"00",X"50",X"00",X"00",X"0F",X"00",X"00",X"50",X"F0",
		X"90",X"0E",X"0E",X"0E",X"0E",X"90",X"A0",X"E0",X"20",X"09",X"0A",X"0B",X"0E",X"E0",X"E0",X"A0",
		X"00",X"0E",X"4B",X"09",X"00",X"E0",X"A0",X"2A",X"00",X"0A",X"0B",X"00",X"00",X"00",X"EA",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"02",X"00",X"00",
		X"2E",X"A0",X"00",X"00",X"90",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"50",X"00",X"00",X"00",X"7B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"20",X"00",X"00",
		X"02",X"0B",X"00",X"00",X"00",X"25",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"79",X"00",X"00",
		X"00",X"79",X"07",X"00",X"00",X"79",X"00",X"00",X"00",X"97",X"00",X"00",X"00",X"97",X"00",X"00",
		X"00",X"97",X"00",X"07",X"00",X"97",X"00",X"00",X"00",X"47",X"40",X"00",X"70",X"44",X"00",X"00",
		X"03",X"44",X"00",X"00",X"70",X"47",X"00",X"00",X"00",X"47",X"00",X"00",X"00",X"97",X"00",X"07",
		X"00",X"97",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"79",X"00",X"00",X"00",X"79",X"07",X"00",
		X"00",X"07",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"77",X"00",X"55",X"00",X"55",
		X"00",X"C5",X"00",X"CC",X"00",X"50",X"00",X"CC",X"00",X"00",X"00",X"5C",X"00",X"00",X"00",X"05",
		X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",
		X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",X"00",X"00",X"55",X"05",X"00",X"00",X"CC",X"00",
		X"00",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"05",X"00",X"05",X"05",X"05",
		X"00",X"5C",X"00",X"05",X"55",X"55",X"05",X"55",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"75",X"00",X"00",X"00",X"50",X"00",
		X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",X"00",X"55",X"55",X"55",X"00",X"CC",X"CC",X"C5",
		X"00",X"CC",X"CC",X"C5",X"00",X"CC",X"CC",X"C5",X"00",X"CC",X"55",X"55",X"00",X"CC",X"00",X"05",
		X"00",X"C5",X"00",X"55",X"00",X"50",X"00",X"C5",X"00",X"00",X"00",X"C5",X"00",X"00",X"00",X"55",
		X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",
		X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"C5",X"00",X"50",X"00",X"C5",X"00",X"C5",X"00",X"55",
		X"00",X"CC",X"00",X"05",X"00",X"CC",X"55",X"55",X"00",X"CC",X"CC",X"C5",X"00",X"CC",X"CC",X"C5",
		X"00",X"CC",X"CC",X"C5",X"00",X"55",X"55",X"55",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
