`define BUILD_DATE "190416"
`define BUILD_TIME "173104"
