library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity mpb_13n is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of mpb_13n is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"A0",X"A0",X"00",X"A0",X"A0",X"B8",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"7F",X"FF",X"F8",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"00",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F2",X"1E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"18",X"7E",X"7E",X"FF",X"FF",X"FF",X"7E",X"7E",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"18",X"7E",X"7E",X"FF",X"FF",X"FF",X"7E",X"7E",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"30",X"78",X"78",X"FC",X"FC",X"78",X"78",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"30",X"78",X"78",X"FC",X"FC",X"78",X"78",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"04",X"00",X"03",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"03",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0C",X"3E",X"78",X"F3",X"E7",X"EC",X"C8",X"00",X"01",X"01",X"03",X"03",X"01",
		X"00",X"00",X"00",X"20",X"70",X"F8",X"E0",X"40",X"40",X"00",X"80",X"C0",X"E0",X"F0",X"F0",X"E0",
		X"03",X"06",X"00",X"00",X"00",X"01",X"03",X"07",X"07",X"07",X"07",X"03",X"01",X"00",X"00",X"00",
		X"C3",X"87",X"0F",X"0F",X"0F",X"CF",X"E7",X"E3",X"F0",X"F0",X"E0",X"E0",X"C0",X"00",X"00",X"00",
		X"81",X"C0",X"C0",X"E0",X"E0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"1F",X"3F",X"3F",X"3F",X"3F",
		X"00",X"00",X"00",X"08",X"00",X"12",X"B0",X"E8",X"38",X"1C",X"04",X"00",X"00",X"80",X"8E",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"1E",X"1F",X"0F",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"E0",X"E0",
		X"1F",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"3F",X"3F",X"3F",X"1F",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"83",X"80",X"00",X"00",X"00",X"02",X"07",X"07",X"0F",X"0F",X"07",X"07",X"03",X"00",X"00",
		X"20",X"80",X"E0",X"70",X"78",X"30",X"10",X"00",X"80",X"C0",X"C0",X"80",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"06",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"60",X"19",X"07",X"03",
		X"02",X"01",X"21",X"11",X"10",X"08",X"0D",X"CF",X"E7",X"7F",X"7F",X"FF",X"FC",X"F0",X"C0",X"80",
		X"00",X"00",X"10",X"10",X"89",X"89",X"0B",X"1F",X"1F",X"BE",X"1C",X"08",X"00",X"00",X"00",X"00",
		X"40",X"44",X"82",X"82",X"8E",X"DF",X"FF",X"FF",X"81",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"08",X"10",X"10",X"30",X"60",X"E1",X"F3",X"FF",X"7F",X"3F",X"0F",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"80",X"00",X"80",X"80",X"C6",X"F8",X"E0",X"80",X"80",
		X"03",X"01",X"01",X"03",X"07",X"1D",X"61",X"01",X"00",X"03",X"03",X"04",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"F3",X"7F",X"38",X"30",X"10",X"20",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"E0",X"E0",X"F9",X"FF",X"7F",X"12",X"10",X"08",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"7E",X"7E",X"FF",X"BD",X"39",X"10",X"10",X"20",X"20",
		X"03",X"03",X"03",X"03",X"07",X"07",X"0E",X"1C",X"1C",X"3E",X"F6",X"F3",X"60",X"20",X"20",X"10",
		X"C0",X"80",X"00",X"80",X"C0",X"60",X"20",X"18",X"00",X"00",X"00",X"00",X"80",X"80",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"1F",X"1F",X"3F",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"7C",X"FD",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"F0",X"F8",X"FC",X"FC",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"3F",X"3F",X"3F",X"1F",X"0F",X"07",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"B1",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"F0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FC",X"FC",X"F8",X"F0",X"F8",X"F8",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"33",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"E6",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"3C",X"7D",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",X"EC",X"FE",X"FE",X"FC",X"FC",X"F8",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"3F",X"7F",X"FF",X"FF",X"7D",X"38",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7C",X"78",X"30",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"F3",X"E0",X"60",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FE",X"FE",X"FC",X"D8",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"03",X"0F",X"1F",X"1F",X"1F",X"0F",X"0F",X"06",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"8E",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"30",X"00",X"00",X"00",
		X"00",X"00",X"00",X"30",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C6",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"F0",X"F8",X"F8",X"F8",X"F0",X"F0",X"30",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"1F",X"1F",X"1F",X"0F",X"03",X"01",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"9C",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F3",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"70",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",X"60",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"E0",X"F0",X"F0",X"F0",X"F0",X"E0",X"E0",X"40",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"3F",X"7F",X"7F",X"3F",X"0C",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"F0",X"FC",X"FE",X"FE",X"F4",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"2C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"20",X"70",X"F0",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"32",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"60",X"F0",X"70",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"60",X"F0",X"F8",X"F8",X"F8",X"F0",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"03",X"03",X"03",X"01",X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"D0",X"F8",X"FC",X"F8",X"FC",X"FC",X"FC",X"FC",X"F8",X"D0",X"00",X"00",X"00",X"00",
		X"00",X"03",X"07",X"07",X"0F",X"0F",X"07",X"0F",X"0F",X"0F",X"07",X"03",X"03",X"01",X"00",X"00",
		X"F0",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"FE",X"FC",X"B8",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"38",X"78",X"78",X"7C",X"FE",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0E",X"1F",X"1F",X"1F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"60",X"E0",X"E0",X"E0",X"E0",X"F0",X"F0",X"F0",X"F8",X"FC",X"FC",
		X"00",X"03",X"03",X"07",X"07",X"0F",X"0F",X"3F",X"3F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"C0",X"E0",X"E0",X"F0",X"E0",X"E0",X"F0",X"F0",X"F0",X"E0",X"F0",X"F0",X"F8",X"FC",X"FE",
		X"07",X"07",X"0F",X"1F",X"1F",X"3F",X"3F",X"3F",X"3F",X"7F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",
		X"00",X"00",X"80",X"80",X"80",X"80",X"E0",X"F0",X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"07",X"07",X"07",X"03",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"E0",X"E0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"0F",X"0F",X"1F",X"1F",X"1F",X"1F",X"1F",X"0F",X"0F",X"03",X"00",X"00",
		X"00",X"00",X"00",X"80",X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"E0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"03",X"0F",X"0F",X"1F",X"1F",X"1F",X"1F",X"1F",X"0F",X"0F",X"03",X"00",X"00",
		X"00",X"00",X"00",X"80",X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"E0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"03",X"0F",X"0F",X"1F",X"1F",X"1F",X"1F",X"1F",X"0F",X"0F",X"03",X"00",X"00",
		X"00",X"00",X"00",X"80",X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"E0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"0F",X"0F",X"1F",X"1F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"1F",X"1F",X"0F",X"0F",X"03",
		X"C0",X"F0",X"F0",X"F8",X"F8",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"F8",X"F8",X"F0",X"F0",X"C0",
		X"03",X"0F",X"0F",X"1F",X"1F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"1F",X"1F",X"0F",X"0F",X"03",
		X"C0",X"F0",X"F0",X"F8",X"F8",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"F8",X"F8",X"F0",X"F0",X"C0",
		X"03",X"07",X"FF",X"FF",X"0F",X"0F",X"00",X"03",X"37",X"7B",X"CE",X"84",X"84",X"CE",X"7B",X"31",
		X"E0",X"F0",X"F0",X"F8",X"F8",X"F8",X"00",X"C0",X"E6",X"DE",X"73",X"21",X"21",X"73",X"DE",X"8C",
		X"00",X"00",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"78",X"7E",X"3F",X"1E",X"0C",X"00",X"3C",X"3C",X"00",X"07",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"1F",X"1F",X"3F",X"00",X"00",X"01",X"00",X"03",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"80",X"00",X"F8",X"F8",X"00",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"84",X"84",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"07",X"0F",X"0F",X"07",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"E0",X"E0",X"F0",X"F0",X"F0",X"E0",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"07",X"0F",X"1F",X"3F",X"3F",X"1F",X"1F",X"1F",X"0F",X"03",X"01",X"00",X"00",
		X"00",X"00",X"C0",X"C0",X"E0",X"F0",X"E0",X"F0",X"F0",X"F0",X"E0",X"E0",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"07",X"0F",X"0F",X"1F",X"1F",X"1F",X"0F",X"1F",X"06",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"E0",X"F0",X"F8",X"F8",X"F8",X"F0",X"F8",X"F0",X"40",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0D",X"0F",X"3F",X"3F",X"3F",X"7F",X"3F",X"1F",X"1F",X"0F",X"03",X"00",X"00",
		X"00",X"00",X"60",X"F0",X"F8",X"FC",X"FC",X"FC",X"F8",X"F8",X"FC",X"F8",X"F8",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"3C",X"7F",X"FC",X"38",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"78",X"FC",X"7E",X"38",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"10",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"20",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"08",X"00",X"00",X"00",X"02",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"10",X"10",X"00",X"00",X"00",X"40",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"0F",X"3F",X"FF",X"FF",X"3F",X"07",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"F0",X"FC",X"FF",X"FF",X"FC",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"0F",X"3F",X"FF",X"FF",X"3F",X"07",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"F0",X"FC",X"FF",X"FF",X"FC",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"0F",X"3F",X"FF",X"FF",X"3F",X"07",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"F0",X"FC",X"FF",X"FF",X"FC",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"03",X"01",X"03",X"02",X"04",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"60",X"C0",X"C0",X"E0",X"80",X"80",X"40",X"40",X"20",X"00",X"00",
		X"00",X"08",X"04",X"00",X"00",X"06",X"03",X"07",X"2F",X"0F",X"1B",X"23",X"49",X"21",X"02",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"80",X"C0",X"E0",X"80",X"80",X"00",X"80",X"40",X"00",X"00",
		X"02",X"81",X"44",X"32",X"09",X"0D",X"07",X"03",X"07",X"4D",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"20",X"88",X"B0",X"E1",X"F4",X"F8",X"F0",X"A6",X"10",X"8C",X"02",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"14",X"0F",X"5C",X"30",X"E6",X"2F",X"DF",X"0F",X"07",X"03",X"01",X"00",X"00",X"00",X"00",
		X"00",X"A0",X"C0",X"E4",X"38",X"8D",X"E6",X"F7",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"0F",X"2F",X"39",X"F0",X"C0",X"82",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"F4",X"FE",X"9F",X"0F",X"03",X"41",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",
		X"03",X"07",X"07",X"06",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"1F",X"3F",X"3C",X"78",X"3C",X"0E",X"07",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"F8",X"FC",X"FC",X"3E",X"78",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"60",X"70",X"38",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"07",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"27",X"3F",X"3F",X"FF",X"F9",X"F0",X"E0",X"C5",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"60",X"FB",X"FF",X"7F",X"1F",X"0B",X"82",X"A0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"C0",X"E0",X"E0",
		X"0F",X"0E",X"1E",X"1E",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"87",X"1F",X"3F",X"3F",X"7F",X"7F",X"1F",X"0F",X"07",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F8",X"F8",X"FC",X"FE",X"FC",X"F8",X"F0",X"E0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"F0",X"7C",X"FC",X"3C",X"1E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"05",X"07",X"07",X"0F",X"0F",X"1F",X"1F",X"7D",
		X"08",X"04",X"0D",X"8F",X"5F",X"FF",X"FF",X"FF",X"FF",X"EF",X"F7",X"F2",X"E0",X"E0",X"C0",X"00",
		X"20",X"40",X"E0",X"F8",X"FC",X"FE",X"FF",X"FF",X"DF",X"BF",X"3F",X"1D",X"0B",X"07",X"03",X"01",
		X"00",X"00",X"00",X"00",X"00",X"40",X"80",X"90",X"E0",X"E0",X"E0",X"F4",X"F8",X"F8",X"F8",X"BC",
		X"3E",X"3E",X"3E",X"1C",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"08",X"05",X"0F",X"1F",X"07",X"02",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"90",X"A0",X"F0",X"E0",X"C0",X"C0",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"78",X"3C",X"3C",X"1A",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"01",X"01",X"03",X"0B",X"07",X"07",X"0F",X"0F",X"1F",
		X"01",X"27",X"1F",X"3F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"F8",
		X"20",X"E4",X"F8",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"D0",X"E0",X"E0",X"F0",X"F0",X"F8",X"F8",X"F8",
		X"1F",X"1F",X"1F",X"0F",X"07",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"E0",X"F0",X"F4",X"FC",X"FE",X"FF",X"FF",X"7F",X"3F",X"3F",X"0F",X"03",X"01",X"01",X"00",
		X"03",X"0F",X"1F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FE",X"FC",X"F8",X"F8",X"F0",X"C0",X"80",X"00",
		X"F8",X"F0",X"E0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"01",X"21",X"14",X"14",X"42",X"22",X"14",X"98",X"38",X"04",X"80",X"00",X"00",
		X"00",X"00",X"00",X"50",X"00",X"A4",X"28",X"40",X"42",X"44",X"2C",X"01",X"02",X"0C",X"00",X"00",
		X"00",X"00",X"10",X"10",X"09",X"0D",X"86",X"10",X"48",X"08",X"08",X"04",X"00",X"00",X"00",X"00",
		X"80",X"00",X"80",X"80",X"04",X"A8",X"48",X"11",X"10",X"12",X"24",X"00",X"00",X"00",X"00",X"00",
		X"01",X"25",X"10",X"09",X"09",X"45",X"47",X"2E",X"32",X"80",X"10",X"00",X"00",X"08",X"00",X"00",
		X"00",X"10",X"94",X"A0",X"E2",X"F4",X"34",X"1D",X"0E",X"04",X"08",X"00",X"00",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"04",X"82",X"52",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"40",X"41",X"82",X"CA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"07",X"01",X"00",X"12",X"28",X"06",X"04",X"00",X"00",X"00",X"00",
		X"51",X"29",X"BB",X"5F",X"3F",X"BE",X"FC",X"98",X"08",X"04",X"00",X"00",X"00",X"00",X"00",X"00",
		X"D4",X"DC",X"FE",X"FC",X"99",X"1A",X"0E",X"0C",X"12",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"00",X"00",X"00",X"80",X"00",X"00",X"20",X"D0",X"80",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"01",X"01",X"01",X"08",X"08",X"04",X"24",X"14",X"95",X"55",X"4F",X"2F",X"BF",X"7F",X"7F",
		X"00",X"00",X"00",X"00",X"80",X"88",X"C2",X"42",X"C4",X"CC",X"CC",X"D8",X"F8",X"F9",X"FE",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"26",X"03",X"23",X"10",X"08",X"08",X"F7",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"FF",X"7F",X"3C",X"B8",X"38",X"0C",X"88",X"08",X"04",X"00",X"00",X"10",X"00",X"20",X"00",
		X"FE",X"FC",X"FF",X"7F",X"26",X"20",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",
		X"00",X"40",X"80",X"00",X"20",X"40",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"18",X"3F",X"7F",X"EF",X"8D",X"18",X"11",X"01",X"02",X"00",X"00",X"00",X"00",
		X"00",X"20",X"10",X"20",X"00",X"F0",X"F0",X"E0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"18",X"00",X"00",X"00",X"18",X"38",X"30",X"91",X"81",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"03",X"03",X"01",X"00",X"18",X"7C",X"FF",X"8F",X"3F",X"3C",X"61",X"01",X"03",X"02",
		X"80",X"40",X"40",X"60",X"60",X"20",X"00",X"00",X"80",X"F0",X"F0",X"F0",X"E0",X"C0",X"00",X"00",
		X"01",X"08",X"04",X"0C",X"03",X"01",X"00",X"18",X"7C",X"FF",X"8F",X"3F",X"3C",X"61",X"01",X"03",
		X"00",X"80",X"C0",X"40",X"60",X"60",X"20",X"00",X"00",X"80",X"E0",X"F0",X"F0",X"E0",X"C0",X"00",
		X"01",X"08",X"04",X"06",X"02",X"07",X"01",X"00",X"18",X"7C",X"7F",X"CF",X"9F",X"1C",X"31",X"21",
		X"00",X"80",X"C0",X"C0",X"60",X"60",X"60",X"20",X"00",X"00",X"80",X"E0",X"F0",X"F0",X"E0",X"C0",
		X"00",X"00",X"03",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"40",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"04",X"01",X"08",X"02",X"00",X"04",X"02",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"00",X"20",X"00",X"A0",X"00",X"40",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"3E",X"FF",X"1E",X"0C",X"00",X"00",X"00",
		X"00",X"00",X"00",X"78",X"7E",X"3F",X"1E",X"0C",X"00",X"3C",X"3C",X"00",X"07",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"3F",X"06",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"78",X"7E",X"3F",X"1E",X"0C",X"00",X"3C",X"3C",X"00",X"07",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"25",X"05",X"09",X"05",X"25",X"18",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C6",X"29",X"29",X"29",X"29",X"29",X"C6",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"25",X"25",X"19",X"25",X"25",X"18",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C6",X"29",X"29",X"29",X"29",X"29",X"C6",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
