library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity crater_bg_bits_2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of crater_bg_bits_2 is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"04",X"0A",X"AA",X"80",X"00",X"00",X"00",X"00",X"02",X"08",X"AA",X"A0",X"00",
		X"00",X"00",X"01",X"12",X"8A",X"AA",X"8A",X"AA",X"00",X"00",X"00",X"00",X"20",X"AA",X"20",X"AA",
		X"00",X"00",X"01",X"48",X"08",X"2A",X"A8",X"8A",X"00",X"00",X"01",X"00",X"42",X"2A",X"A0",X"AA",
		X"00",X"00",X"05",X"00",X"18",X"2A",X"8A",X"AA",X"00",X"00",X"40",X"00",X"1A",X"08",X"8A",X"A8",
		X"00",X"00",X"10",X"00",X"18",X"28",X"A2",X"A8",X"00",X"00",X"00",X"00",X"04",X"82",X"AA",X"AA",
		X"00",X"01",X"00",X"00",X"04",X"82",X"AA",X"85",X"00",X"20",X"00",X"00",X"40",X"A2",X"AA",X"00",
		X"01",X"20",X"00",X"00",X"00",X"A0",X"2A",X"92",X"00",X"00",X"00",X"00",X"40",X"A2",X"00",X"9A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"A8",
		X"A8",X"28",X"00",X"02",X"A0",X"A2",X"AA",X"AA",X"2A",X"A0",X"08",X"00",X"0A",X"0A",X"AA",X"8A",
		X"82",X"AA",X"18",X"2A",X"2A",X"AA",X"AA",X"8A",X"AA",X"A8",X"6A",X"22",X"2A",X"AA",X"AA",X"22",
		X"A8",X"02",X"9A",X"2A",X"8A",X"AA",X"A8",X"82",X"AA",X"26",X"02",X"82",X"A2",X"AA",X"AA",X"2A",
		X"82",X"AA",X"22",X"8A",X"AA",X"AA",X"AA",X"8A",X"02",X"08",X"28",X"AA",X"2A",X"AA",X"8A",X"A0",
		X"06",X"22",X"8A",X"8A",X"AA",X"AA",X"A8",X"AA",X"82",X"82",X"02",X"AA",X"AA",X"AA",X"22",X"AA",
		X"8A",X"AA",X"A2",X"A8",X"22",X"AA",X"2A",X"AA",X"0A",X"A8",X"2A",X"0A",X"AA",X"2A",X"AA",X"A8",
		X"A0",X"A0",X"AA",X"AA",X"AA",X"A8",X"AA",X"A2",X"AA",X"A8",X"80",X"8A",X"AA",X"A8",X"A8",X"82",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"AA",
		X"A9",X"40",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"00",X"00",X"02",X"AA",X"2A",X"AA",X"2A",
		X"AA",X"AA",X"AA",X"00",X"0A",X"AA",X"A8",X"2A",X"8A",X"AA",X"A0",X"AA",X"22",X"8A",X"A8",X"AA",
		X"80",X"8A",X"8A",X"AA",X"22",X"AA",X"29",X"8A",X"AA",X"A2",X"82",X"AA",X"22",X"AA",X"A0",X"AA",
		X"AA",X"A2",X"8A",X"0A",X"A2",X"A2",X"80",X"82",X"AA",X"A2",X"AA",X"0A",X"AA",X"A2",X"00",X"A2",
		X"AA",X"28",X"2A",X"A8",X"AA",X"AA",X"11",X"20",X"AA",X"8A",X"A2",X"AA",X"20",X"AA",X"02",X"20",
		X"A0",X"0A",X"AA",X"02",X"2A",X"A8",X"02",X"28",X"2A",X"2A",X"28",X"28",X"2A",X"A8",X"04",X"28",
		X"AA",X"AA",X"A2",X"A2",X"08",X"88",X"04",X"2A",X"2A",X"02",X"82",X"A0",X"AA",X"A8",X"10",X"2A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"A8",X"08",X"00",X"00",X"09",X"00",X"00",X"00",X"AA",X"94",X"00",X"14",X"2A",X"55",X"55",X"50",
		X"AA",X"00",X"0A",X"20",X"0A",X"A8",X"15",X"92",X"AA",X"92",X"6A",X"80",X"8A",X"2A",X"AA",X"25",
		X"AA",X"0A",X"AA",X"00",X"AA",X"A2",X"28",X"AA",X"A8",X"02",X"AA",X"02",X"A2",X"AA",X"2A",X"AA",
		X"AA",X"5A",X"08",X"00",X"2A",X"AA",X"A2",X"AA",X"AA",X"02",X"88",X"42",X"2A",X"AA",X"AA",X"AA",
		X"A8",X"48",X"80",X"0A",X"AA",X"AA",X"AA",X"AA",X"A8",X"0A",X"82",X"AA",X"AA",X"AA",X"AA",X"A8",
		X"20",X"28",X"A2",X"2A",X"AA",X"AA",X"AA",X"A8",X"28",X"28",X"A2",X"2A",X"AA",X"22",X"AA",X"AA",
		X"08",X"82",X"A0",X"8A",X"AA",X"2A",X"AA",X"AA",X"0A",X"0A",X"88",X"A2",X"AA",X"88",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"10",X"00",X"00",X"00",X"00",
		X"04",X"25",X"40",X"29",X"90",X"10",X"00",X"00",X"24",X"A2",X"A8",X"A0",X"AA",X"A5",X"40",X"00",
		X"95",X"05",X"02",X"88",X"88",X"00",X"08",X"00",X"5A",X"22",X"2A",X"A2",X"AA",X"42",X"00",X"2A",
		X"22",X"22",X"82",X"A1",X"14",X"02",X"A2",X"00",X"AA",X"22",X"AA",X"AA",X"81",X"0A",X"A2",X"20",
		X"2A",X"A2",X"22",X"A0",X"A0",X"02",X"88",X"28",X"AA",X"AA",X"A8",X"AA",X"8A",X"2A",X"22",X"28",
		X"A8",X"AA",X"AA",X"2A",X"A8",X"8A",X"8A",X"AA",X"A2",X"88",X"AA",X"A8",X"A2",X"6A",X"82",X"A2",
		X"AA",X"AA",X"AA",X"2A",X"A2",X"AA",X"82",X"AA",X"28",X"AA",X"AA",X"AA",X"A8",X"AA",X"A2",X"8A",
		X"22",X"AA",X"8A",X"2A",X"AA",X"88",X"A0",X"AA",X"0A",X"2A",X"A8",X"AA",X"AA",X"22",X"20",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"01",X"00",X"00",X"00",X"01",
		X"02",X"95",X"44",X"00",X"10",X"01",X"A6",X"A0",X"AA",X"AA",X"A4",X"5A",X"2A",X"00",X"AA",X"91",
		X"A8",X"2A",X"AA",X"AA",X"29",X"AA",X"88",X"AA",X"AA",X"82",X"AA",X"A0",X"15",X"0A",X"AA",X"A8",
		X"AA",X"A2",X"A8",X"AA",X"18",X"AA",X"80",X"A8",X"AA",X"A8",X"8A",X"AA",X"A0",X"A0",X"A8",X"88",
		X"A8",X"AA",X"AA",X"A0",X"82",X"A0",X"A0",X"0A",X"A2",X"8A",X"AA",X"AA",X"A2",X"AA",X"88",X"82",
		X"AA",X"82",X"A8",X"AA",X"8A",X"82",X"A0",X"AA",X"AA",X"8A",X"08",X"AA",X"18",X"A0",X"20",X"0A",
		X"AA",X"8A",X"AA",X"8A",X"28",X"82",X"28",X"8A",X"A0",X"AA",X"0A",X"AA",X"28",X"A0",X"A8",X"A2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A8",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"50",X"00",X"00",X"00",X"00",X"00",X"00",
		X"28",X"48",X"00",X"00",X"00",X"00",X"00",X"00",X"28",X"46",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A8",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"A8",X"52",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A8",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"A5",X"16",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A4",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"25",X"02",X"80",X"00",X"00",X"00",X"00",X"00",
		X"24",X"06",X"80",X"00",X"00",X"00",X"00",X"00",X"A5",X"02",X"80",X"00",X"00",X"00",X"00",X"00",
		X"08",X"00",X"00",X"00",X"08",X"00",X"01",X"55",X"00",X"00",X"10",X"05",X"A5",X"55",X"55",X"55",
		X"00",X"00",X"05",X"55",X"55",X"55",X"55",X"54",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"50",
		X"00",X"91",X"55",X"55",X"55",X"55",X"55",X"40",X"02",X"95",X"55",X"55",X"55",X"55",X"55",X"40",
		X"15",X"55",X"55",X"55",X"55",X"55",X"55",X"40",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"10",X"55",X"55",X"55",X"55",X"55",X"55",X"54",X"40",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"50",X"55",X"55",X"51",X"55",X"55",X"55",X"41",X"00",
		X"55",X"55",X"40",X"95",X"55",X"40",X"00",X"00",X"55",X"55",X"41",X"85",X"40",X"00",X"10",X"11",
		X"55",X"55",X"10",X"0A",X"00",X"00",X"01",X"00",X"55",X"54",X"00",X"12",X"80",X"00",X"41",X"10",
		X"00",X"90",X"00",X"00",X"00",X"8A",X"00",X"8A",X"00",X"10",X"00",X"00",X"22",X"2A",X"86",X"9A",
		X"00",X"40",X"00",X"00",X"28",X"2A",X"8A",X"20",X"01",X"00",X"00",X"00",X"A0",X"88",X"29",X"08",
		X"00",X"00",X"00",X"06",X"28",X"82",X"88",X"22",X"00",X"00",X"00",X"02",X"22",X"08",X"2A",X"08",
		X"00",X"00",X"00",X"12",X"84",X"88",X"88",X"08",X"00",X"00",X"00",X"18",X"82",X"08",X"22",X"0A",
		X"00",X"00",X"10",X"18",X"00",X"12",X"20",X"82",X"01",X"08",X"40",X"20",X"41",X"00",X"0A",X"28",
		X"04",X"24",X"00",X"00",X"00",X"00",X"0A",X"A0",X"40",X"24",X"00",X"00",X"00",X"00",X"00",X"A0",
		X"10",X"A0",X"00",X"00",X"00",X"00",X"08",X"A8",X"08",X"20",X"00",X"00",X"00",X"14",X"28",X"28",
		X"08",X"10",X"00",X"00",X"00",X"00",X"A8",X"A8",X"00",X"40",X"00",X"00",X"04",X"4A",X"22",X"A8",
		X"08",X"2A",X"80",X"8A",X"00",X"2A",X"A0",X"0A",X"02",X"A2",X"02",X"A2",X"AA",X"AA",X"28",X"AA",
		X"8A",X"AA",X"02",X"2A",X"AA",X"AA",X"AA",X"0A",X"AA",X"8A",X"82",X"AA",X"82",X"80",X"AA",X"88",
		X"A8",X"8A",X"00",X"AA",X"AA",X"AA",X"AA",X"A8",X"AA",X"A2",X"02",X"A8",X"AA",X"AA",X"80",X"82",
		X"8A",X"A2",X"A0",X"A0",X"AA",X"88",X"AA",X"AA",X"A2",X"A8",X"A0",X"08",X"AA",X"AA",X"A8",X"8A",
		X"AA",X"28",X"A8",X"8A",X"AA",X"88",X"88",X"AA",X"8A",X"AA",X"2A",X"A2",X"08",X"28",X"A2",X"8A",
		X"A2",X"A8",X"8A",X"AA",X"22",X"A2",X"82",X"88",X"A8",X"A8",X"82",X"0A",X"A0",X"28",X"A2",X"AA",
		X"8A",X"2A",X"A0",X"2A",X"20",X"AA",X"82",X"2A",X"22",X"A8",X"0A",X"2A",X"A0",X"2A",X"0A",X"82",
		X"8A",X"00",X"2A",X"80",X"08",X"8A",X"80",X"A0",X"8A",X"28",X"A8",X"00",X"00",X"28",X"AA",X"AA",
		X"A0",X"AA",X"8A",X"0A",X"A2",X"A8",X"10",X"A2",X"A2",X"0A",X"88",X"AA",X"AA",X"88",X"10",X"A8",
		X"A2",X"02",X"82",X"AA",X"2A",X"80",X"40",X"AA",X"2A",X"AA",X"82",X"2A",X"AA",X"80",X"00",X"2A",
		X"A8",X"2A",X"A0",X"A8",X"AA",X"04",X"00",X"A8",X"AA",X"A8",X"2A",X"82",X"A2",X"00",X"02",X"A8",
		X"A8",X"A8",X"2A",X"AA",X"A8",X"80",X"02",X"A2",X"28",X"2A",X"2A",X"AA",X"A8",X"00",X"0A",X"88",
		X"0A",X"8A",X"AA",X"2A",X"22",X"00",X"0A",X"0A",X"8A",X"0A",X"AA",X"2A",X"22",X"00",X"08",X"2A",
		X"2A",X"0A",X"AA",X"AA",X"22",X"00",X"28",X"A2",X"AA",X"2A",X"AA",X"AA",X"A8",X"00",X"22",X"2A",
		X"AA",X"AA",X"AA",X"AA",X"88",X"02",X"A0",X"62",X"A8",X"AA",X"82",X"A8",X"00",X"00",X"A0",X"0A",
		X"0A",X"A2",X"AA",X"A8",X"10",X"00",X"01",X"0A",X"A0",X"20",X"A8",X"A8",X"04",X"00",X"00",X"88",
		X"02",X"AA",X"A8",X"22",X"28",X"AA",X"AA",X"AA",X"A0",X"AA",X"AA",X"80",X"AA",X"AA",X"AA",X"AA",
		X"A0",X"A8",X"2A",X"AA",X"8A",X"A8",X"AA",X"AA",X"00",X"A2",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"82",X"8A",X"88",X"AA",X"2A",X"0A",X"A8",X"AA",X"22",X"AA",X"8A",X"AA",X"2A",X"AA",X"AA",X"AA",
		X"20",X"AA",X"A8",X"8A",X"A2",X"02",X"AA",X"AA",X"A0",X"8A",X"AA",X"8A",X"AA",X"AA",X"AA",X"A8",
		X"20",X"2A",X"2A",X"AA",X"28",X"22",X"AA",X"AA",X"28",X"0A",X"AA",X"AA",X"AA",X"A2",X"AA",X"AA",
		X"8A",X"82",X"A8",X"AA",X"AA",X"AA",X"A2",X"AA",X"2A",X"82",X"AA",X"AA",X"AA",X"AA",X"AA",X"8A",
		X"2A",X"A8",X"2A",X"AA",X"2A",X"A8",X"AA",X"AA",X"AA",X"8A",X"0A",X"8A",X"A2",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"A2",X"AA",X"2A",X"A8",X"AA",X"AA",X"AA",X"22",X"AA",X"A8",X"AA",X"AA",X"22",X"AA",
		X"AA",X"2A",X"2A",X"AA",X"A8",X"00",X"2A",X"A8",X"AA",X"AA",X"AA",X"AA",X"2A",X"02",X"8A",X"88",
		X"A2",X"88",X"A8",X"A2",X"00",X"8A",X"0A",X"8A",X"AA",X"AA",X"AA",X"A2",X"AA",X"A0",X"2A",X"2A",
		X"AA",X"AA",X"A8",X"AA",X"AA",X"A0",X"AA",X"2A",X"AA",X"AA",X"AA",X"AA",X"A2",X"82",X"02",X"2A",
		X"AA",X"AA",X"A8",X"AA",X"AA",X"08",X"2A",X"28",X"A2",X"AA",X"A2",X"A8",X"20",X"58",X"2A",X"2A",
		X"AA",X"A8",X"AA",X"AA",X"09",X"2A",X"A8",X"A2",X"A8",X"AA",X"AA",X"2A",X"A5",X"A0",X"A2",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"6A",X"00",X"20",X"A0",X"AA",X"AA",X"AA",X"2A",X"80",X"82",X"2A",X"8A",
		X"AA",X"A2",X"AA",X"8A",X"28",X"A0",X"AA",X"8A",X"AA",X"AA",X"8A",X"88",X"08",X"8A",X"A2",X"A2",
		X"AA",X"AA",X"8A",X"82",X"20",X"82",X"2A",X"28",X"A2",X"AA",X"08",X"A8",X"02",X"2A",X"28",X"AA",
		X"A0",X"A8",X"AA",X"AA",X"20",X"A2",X"A8",X"A2",X"8A",X"A2",X"A8",X"AA",X"04",X"22",X"A8",X"AA",
		X"8A",X"A2",X"AA",X"A8",X"A8",X"22",X"A0",X"82",X"A8",X"8A",X"A8",X"AA",X"82",X"28",X"88",X"AA",
		X"8A",X"8A",X"8A",X"0A",X"1A",X"08",X"AA",X"AA",X"AA",X"8A",X"A8",X"AA",X"A8",X"2A",X"AA",X"AA",
		X"8A",X"22",X"AA",X"8A",X"16",X"AA",X"A2",X"AA",X"8A",X"2A",X"AA",X"AA",X"2A",X"8A",X"A2",X"AA",
		X"8A",X"28",X"A8",X"A2",X"0A",X"4A",X"22",X"AA",X"88",X"28",X"AA",X"A0",X"2A",X"88",X"A2",X"AA",
		X"A8",X"2A",X"8A",X"A2",X"AA",X"A8",X"AA",X"AA",X"A8",X"2A",X"8A",X"88",X"2A",X"A8",X"AA",X"8A",
		X"A8",X"0A",X"82",X"80",X"A8",X"20",X"A8",X"8A",X"A8",X"0A",X"28",X"88",X"2A",X"A2",X"A8",X"8A",
		X"A2",X"0A",X"20",X"AA",X"20",X"92",X"80",X"8A",X"A2",X"2A",X"28",X"AA",X"2A",X"62",X"AA",X"AA",
		X"A1",X"11",X"80",X"00",X"00",X"00",X"00",X"00",X"A4",X"04",X"20",X"00",X"00",X"00",X"00",X"00",
		X"A4",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"12",X"00",X"00",X"00",X"00",X"00",
		X"20",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"02",X"00",X"00",X"00",X"00",X"20",
		X"A0",X"08",X"02",X"00",X"00",X"00",X"00",X"20",X"A0",X"00",X"02",X"80",X"00",X"00",X"00",X"28",
		X"A0",X"00",X"42",X"80",X"00",X"00",X"00",X"A0",X"80",X"00",X"40",X"80",X"00",X"00",X"2A",X"A0",
		X"84",X"00",X"50",X"A0",X"00",X"02",X"AA",X"A8",X"94",X"00",X"40",X"20",X"00",X"2A",X"8A",X"80",
		X"10",X"00",X"40",X"28",X"00",X"00",X"0A",X"05",X"A0",X"00",X"40",X"28",X"00",X"00",X"01",X"50",
		X"90",X"00",X"40",X"28",X"00",X"00",X"55",X"02",X"40",X"00",X"44",X"2A",X"00",X"05",X"54",X"02",
		X"55",X"54",X"00",X"02",X"00",X"00",X"00",X"00",X"55",X"50",X"08",X"1A",X"88",X"00",X"00",X"00",
		X"55",X"44",X"00",X"48",X"6A",X"00",X"00",X"0A",X"54",X"10",X"08",X"18",X"0A",X"80",X"00",X"AA",
		X"52",X"41",X"08",X"40",X"62",X"80",X"00",X"00",X"41",X"42",X"20",X"10",X"22",X"88",X"00",X"00",
		X"09",X"08",X"00",X"44",X"2A",X"22",X"00",X"00",X"09",X"22",X"01",X"11",X"02",X"2A",X"00",X"00",
		X"20",X"22",X"00",X"10",X"44",X"00",X"00",X"02",X"24",X"20",X"00",X"00",X"00",X"40",X"00",X"00",
		X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"20",X"00",X"00",X"00",X"00",X"10",X"00",X"60",X"00",
		X"22",X"00",X"10",X"00",X"10",X"20",X"28",X"A8",X"28",X"00",X"80",X"00",X"00",X"08",X"A2",X"AA",
		X"A0",X"09",X"80",X"00",X"00",X"08",X"2A",X"2A",X"00",X"22",X"00",X"00",X"00",X"06",X"AA",X"2A",
		X"00",X"A0",X"00",X"00",X"00",X"02",X"AA",X"AA",X"02",X"A0",X"00",X"00",X"00",X"01",X"AA",X"8A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"28",X"AA",X"00",X"00",X"00",X"20",X"00",X"00",X"08",X"A0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"8A",X"28",X"00",X"00",X"00",X"00",X"00",X"00",X"2A",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"80",X"00",X"00",X"00",X"00",X"02",X"00",X"22",X"88",
		X"20",X"00",X"00",X"00",X"00",X"00",X"01",X"16",X"00",X"20",X"00",X"02",X"00",X"00",X"80",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"12",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"82",X"28",X"A0",X"00",X"00",X"02",X"AA",X"08",X"A2",X"AA",X"88",X"00",X"00",X"00",X"8A",X"AA",
		X"A8",X"80",X"00",X"00",X"00",X"00",X"08",X"2A",X"8A",X"00",X"00",X"00",X"00",X"00",X"08",X"0A",
		X"2A",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"A2",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"2A",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"28",X"80",X"00",X"00",X"00",X"00",X"00",
		X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A2",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"22",X"A0",X"A8",X"A8",X"00",X"00",X"02",X"28",X"2A",X"2A",X"A8",X"20",X"10",X"00",X"04",X"22",
		X"2A",X"8A",X"A8",X"20",X"00",X"00",X"00",X"20",X"AA",X"A8",X"80",X"60",X"40",X"00",X"00",X"22",
		X"2A",X"0A",X"A9",X"22",X"00",X"00",X"02",X"A2",X"02",X"2A",X"A0",X"28",X"00",X"00",X"18",X"8A",
		X"00",X"00",X"A0",X"A8",X"00",X"00",X"2A",X"8A",X"00",X"08",X"A4",X"A8",X"00",X"00",X"28",X"8A",
		X"00",X"0A",X"A4",X"A8",X"80",X"00",X"2A",X"2A",X"00",X"0A",X"A0",X"AA",X"00",X"00",X"2A",X"AA",
		X"02",X"0A",X"A2",X"A8",X"00",X"00",X"AA",X"AA",X"00",X"A8",X"62",X"A8",X"00",X"02",X"AA",X"8A",
		X"00",X"A9",X"42",X"A8",X"00",X"00",X"A0",X"8A",X"0A",X"88",X"0A",X"A0",X"00",X"00",X"A2",X"AA",
		X"00",X"14",X"42",X"80",X"00",X"00",X"0A",X"8A",X"00",X"41",X"0A",X"A0",X"00",X"00",X"0A",X"A0",
		X"28",X"89",X"22",X"AA",X"A2",X"A8",X"AA",X"AA",X"A2",X"A4",X"80",X"AA",X"AA",X"AA",X"2A",X"A2",
		X"AA",X"A4",X"AA",X"2A",X"AA",X"AA",X"A2",X"AA",X"AA",X"A2",X"28",X"2A",X"AA",X"AA",X"AA",X"8A",
		X"0A",X"80",X"22",X"AA",X"AA",X"AA",X"AA",X"AA",X"0A",X"84",X"8A",X"82",X"8A",X"AA",X"AA",X"AA",
		X"2A",X"0A",X"2A",X"A2",X"22",X"AA",X"AA",X"A8",X"AA",X"08",X"2A",X"A0",X"8A",X"8A",X"AA",X"AA",
		X"A8",X"20",X"AA",X"82",X"08",X"AA",X"AA",X"AA",X"A9",X"22",X"28",X"A2",X"00",X"AA",X"AA",X"A2",
		X"A8",X"2A",X"28",X"AA",X"82",X"AA",X"AA",X"AA",X"8A",X"22",X"A2",X"0A",X"20",X"22",X"AA",X"AA",
		X"0A",X"1A",X"A0",X"AA",X"AA",X"2A",X"A2",X"AA",X"08",X"02",X"A8",X"A2",X"2A",X"02",X"A8",X"AA",
		X"00",X"04",X"8A",X"A8",X"2A",X"82",X"2A",X"AA",X"00",X"0A",X"A2",X"8A",X"8A",X"AA",X"AA",X"A0",
		X"A8",X"AA",X"A8",X"00",X"08",X"A8",X"28",X"A0",X"AA",X"AA",X"A9",X"A0",X"80",X"22",X"A2",X"A0",
		X"AA",X"AA",X"AA",X"A8",X"A0",X"22",X"28",X"A8",X"AA",X"AA",X"AA",X"88",X"02",X"2A",X"28",X"8A",
		X"AA",X"A8",X"AA",X"A8",X"02",X"0A",X"AA",X"88",X"AA",X"AA",X"A2",X"02",X"08",X"A2",X"AA",X"08",
		X"A2",X"AA",X"AA",X"00",X"20",X"0A",X"A2",X"82",X"A8",X"AA",X"2A",X"A8",X"00",X"2A",X"AA",X"0A",
		X"AA",X"AA",X"20",X"82",X"20",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"08",X"00",X"AA",X"28",X"AA",
		X"AA",X"8A",X"AA",X"0A",X"80",X"22",X"AA",X"8A",X"AA",X"A8",X"20",X"A0",X"2A",X"18",X"AA",X"0A",
		X"AA",X"AA",X"A2",X"80",X"80",X"92",X"AA",X"A2",X"AA",X"8A",X"22",X"28",X"0A",X"2A",X"AA",X"82",
		X"AA",X"AA",X"20",X"00",X"82",X"AA",X"AA",X"A2",X"A8",X"A8",X"22",X"00",X"AA",X"8A",X"AA",X"2A",
		X"A2",X"2A",X"0A",X"AA",X"28",X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",X"2A",X"26",X"A8",X"AA",X"AA",
		X"8A",X"A2",X"2A",X"A2",X"A0",X"AA",X"A8",X"AA",X"A8",X"A0",X"28",X"AA",X"90",X"AA",X"AA",X"8A",
		X"AA",X"20",X"AA",X"2A",X"92",X"AA",X"8A",X"AA",X"A2",X"22",X"AA",X"22",X"0A",X"AA",X"AA",X"0A",
		X"AA",X"22",X"0A",X"2A",X"AA",X"AA",X"2A",X"88",X"A8",X"22",X"08",X"A8",X"9A",X"8A",X"AA",X"88",
		X"A8",X"22",X"A0",X"2A",X"A2",X"AA",X"2A",X"8A",X"A2",X"22",X"22",X"A8",X"A0",X"AA",X"A2",X"AA",
		X"A2",X"AA",X"20",X"28",X"A0",X"AA",X"82",X"AA",X"AA",X"02",X"22",X"2A",X"A4",X"A2",X"AA",X"AA",
		X"A8",X"2A",X"8A",X"28",X"A0",X"AA",X"82",X"AA",X"A2",X"A8",X"88",X"A8",X"86",X"AA",X"A2",X"AA",
		X"AA",X"A8",X"AA",X"22",X"86",X"A8",X"A2",X"AA",X"A0",X"A8",X"A8",X"82",X"9A",X"AA",X"A8",X"AA",
		X"40",X"00",X"40",X"2A",X"55",X"55",X"40",X"0A",X"41",X"00",X"10",X"2A",X"55",X"50",X"00",X"AA",
		X"11",X"00",X"00",X"2A",X"50",X"00",X"02",X"AA",X"50",X"60",X"00",X"2A",X"00",X"00",X"02",X"A2",
		X"94",X"00",X"00",X"5A",X"00",X"00",X"00",X"00",X"80",X"00",X"01",X"1A",X"80",X"00",X"00",X"00",
		X"10",X"00",X"20",X"1A",X"80",X"00",X"00",X"00",X"40",X"00",X"00",X"1A",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"1A",X"80",X"00",X"00",X"00",X"80",X"80",X"84",X"5A",X"80",X"00",X"00",X"00",
		X"00",X"00",X"90",X"62",X"80",X"00",X"00",X"00",X"08",X"00",X"40",X"2A",X"80",X"00",X"00",X"00",
		X"20",X"00",X"40",X"62",X"80",X"00",X"00",X"00",X"20",X"00",X"50",X"22",X"80",X"00",X"00",X"00",
		X"20",X"00",X"10",X"0A",X"80",X"00",X"00",X"00",X"00",X"00",X"10",X"8A",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"81",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"84",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",
		X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"80",X"00",X"00",X"02",X"08",X"00",X"40",X"88",X"00",
		X"00",X"02",X"00",X"01",X"A1",X"22",X"02",X"2A",X"00",X"00",X"00",X"02",X"00",X"02",X"08",X"00",
		X"00",X"00",X"00",X"02",X"08",X"20",X"A0",X"20",X"00",X"00",X"00",X"00",X"02",X"AA",X"82",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A1",X"60",X"00",X"00",X"00",X"00",X"00",X"00",
		X"05",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"41",X"A8",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"28",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"0A",X"00",X"00",X"02",X"00",X"00",X"00",
		X"10",X"8A",X"80",X"00",X"02",X"A0",X"00",X"00",X"44",X"08",X"A0",X"00",X"41",X"28",X"00",X"00",
		X"11",X"2A",X"20",X"04",X"14",X"A8",X"80",X"00",X"04",X"28",X"00",X"41",X"40",X"0A",X"80",X"00",
		X"00",X"A8",X"00",X"14",X"10",X"2A",X"00",X"00",X"80",X"00",X"00",X"14",X"40",X"28",X"00",X"00",
		X"00",X"00",X"00",X"40",X"00",X"A8",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"A8",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0A",X"A0",X"20",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",
		X"00",X"04",X"2A",X"40",X"00",X"00",X"00",X"80",X"00",X"12",X"21",X"10",X"00",X"00",X"00",X"80",
		X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"02",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"0A",
		X"00",X"01",X"44",X"40",X"00",X"00",X"00",X"18",X"00",X"10",X"40",X"00",X"00",X"00",X"00",X"08",
		X"00",X"04",X"40",X"00",X"00",X"00",X"00",X"4A",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"2A",
		X"00",X"14",X"00",X"00",X"00",X"00",X"00",X"2A",X"00",X"40",X"00",X"00",X"00",X"00",X"04",X"A8",
		X"00",X"10",X"88",X"00",X"00",X"00",X"02",X"A8",X"00",X"02",X"00",X"00",X"A0",X"00",X"02",X"A2",
		X"02",X"00",X"00",X"02",X"80",X"00",X"02",X"28",X"00",X"00",X"00",X"0A",X"A0",X"00",X"2A",X"20",
		X"00",X"00",X"02",X"08",X"00",X"00",X"AA",X"A0",X"00",X"00",X"02",X"00",X"00",X"00",X"80",X"08",
		X"00",X"2A",X"A8",X"A0",X"AA",X"AA",X"AA",X"8A",X"00",X"A0",X"28",X"88",X"28",X"A2",X"AA",X"A8",
		X"00",X"00",X"A2",X"2A",X"8A",X"22",X"2A",X"22",X"00",X"00",X"02",X"2A",X"88",X"A0",X"8A",X"A2",
		X"80",X"00",X"00",X"AA",X"A8",X"A8",X"88",X"AA",X"80",X"00",X"00",X"A2",X"A8",X"A8",X"8A",X"AA",
		X"00",X"00",X"00",X"20",X"88",X"28",X"82",X"A0",X"80",X"00",X"01",X"08",X"AA",X"AA",X"22",X"80",
		X"00",X"00",X"01",X"08",X"AA",X"82",X"A2",X"8A",X"00",X"00",X"01",X"08",X"A2",X"A0",X"AA",X"AA",
		X"00",X"00",X"00",X"48",X"A2",X"88",X"20",X"20",X"00",X"00",X"00",X"40",X"A0",X"AA",X"A2",X"AA",
		X"00",X"00",X"00",X"40",X"A8",X"28",X"22",X"AA",X"00",X"00",X"00",X"00",X"A8",X"8A",X"22",X"20",
		X"00",X"00",X"01",X"00",X"A8",X"A2",X"88",X"80",X"00",X"00",X"00",X"00",X"A8",X"A8",X"A2",X"00",
		X"AA",X"AA",X"80",X"8A",X"AA",X"2A",X"A2",X"AA",X"A2",X"AA",X"2A",X"AA",X"A8",X"6A",X"AA",X"A2",
		X"AA",X"AA",X"AA",X"AA",X"A6",X"AA",X"22",X"A2",X"2A",X"22",X"8A",X"AA",X"A8",X"2A",X"AA",X"A8",
		X"AA",X"A2",X"A8",X"AA",X"A8",X"AA",X"20",X"AA",X"A2",X"AA",X"AA",X"AA",X"A6",X"AA",X"AA",X"A8",
		X"8A",X"82",X"AA",X"8A",X"A6",X"AA",X"8A",X"88",X"A8",X"AA",X"AA",X"AA",X"AA",X"4A",X"AA",X"A8",
		X"A0",X"02",X"AA",X"AA",X"A8",X"AA",X"AA",X"AA",X"20",X"00",X"00",X"2A",X"AA",X"AA",X"88",X"A8",
		X"00",X"00",X"00",X"0A",X"2A",X"82",X"AA",X"A0",X"2A",X"00",X"00",X"0A",X"8A",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"0A",X"AA",X"AA",X"A8",X"00",X"00",X"00",X"00",X"14",X"AA",X"20",X"00",X"00",
		X"00",X"00",X"00",X"12",X"A8",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"2A",X"00",X"00",X"00",
		X"AA",X"A0",X"AA",X"AA",X"6A",X"AA",X"A8",X"90",X"A8",X"82",X"A2",X"AA",X"6A",X"AA",X"AA",X"91",
		X"AA",X"A8",X"80",X"2A",X"6A",X"AA",X"08",X"10",X"28",X"A2",X"A8",X"02",X"6A",X"28",X"AA",X"10",
		X"A8",X"AA",X"AA",X"09",X"AA",X"A2",X"22",X"80",X"AA",X"2A",X"A0",X"02",X"AA",X"02",X"22",X"00",
		X"20",X"2A",X"8A",X"02",X"AA",X"AA",X"AA",X"00",X"02",X"A0",X"00",X"08",X"A9",X"8A",X"A0",X"00",
		X"80",X"00",X"00",X"0A",X"AA",X"A2",X"A0",X"00",X"80",X"00",X"00",X"00",X"AA",X"AA",X"A0",X"00",
		X"20",X"00",X"00",X"2A",X"AA",X"8A",X"A0",X"00",X"A0",X"00",X"00",X"02",X"AA",X"AA",X"AA",X"00",
		X"00",X"00",X"00",X"20",X"2A",X"2A",X"A8",X"00",X"00",X"00",X"00",X"02",X"2A",X"AA",X"A0",X"00",
		X"00",X"00",X"00",X"0A",X"AA",X"AA",X"80",X"00",X"00",X"00",X"00",X"00",X"A8",X"2A",X"00",X"02",
		X"00",X"00",X"00",X"0A",X"80",X"00",X"00",X"00",X"00",X"00",X"44",X"0A",X"A0",X"00",X"00",X"00",
		X"00",X"00",X"42",X"0A",X"A5",X"00",X"00",X"00",X"00",X"00",X"10",X"0A",X"A5",X"40",X"00",X"00",
		X"00",X"00",X"02",X"0A",X"A5",X"40",X"00",X"00",X"00",X"00",X"48",X"0A",X"A5",X"4A",X"00",X"00",
		X"00",X"00",X"68",X"0A",X"A9",X"5A",X"80",X"00",X"00",X"01",X"00",X"0A",X"A9",X"56",X"00",X"00",
		X"00",X"01",X"00",X"0A",X"AA",X"54",X"00",X"00",X"00",X"05",X"00",X"0A",X"AA",X"55",X"80",X"00",
		X"00",X"05",X"80",X"0A",X"2A",X"55",X"AA",X"00",X"00",X"44",X"00",X"0A",X"2A",X"55",X"58",X"00",
		X"00",X"54",X"00",X"0A",X"2A",X"55",X"58",X"00",X"00",X"50",X"00",X"0A",X"2A",X"55",X"55",X"80",
		X"02",X"00",X"00",X"0A",X"2A",X"95",X"55",X"54",X"20",X"80",X"00",X"0A",X"28",X"95",X"55",X"55",
		X"20",X"00",X"00",X"00",X"00",X"02",X"A8",X"00",X"A8",X"00",X"00",X"00",X"02",X"80",X"A4",X"20",
		X"AA",X"16",X"A0",X"02",X"AA",X"A2",X"A8",X"4A",X"2A",X"68",X"A0",X"00",X"28",X"AA",X"A0",X"A2",
		X"0A",X"9A",X"AA",X"0A",X"8A",X"A2",X"A6",X"8A",X"0A",X"A2",X"A2",X"2A",X"AA",X"AA",X"80",X"A0",
		X"0A",X"AA",X"AA",X"0A",X"AA",X"A2",X"8A",X"08",X"00",X"AA",X"88",X"2A",X"AA",X"AA",X"A0",X"AA",
		X"0A",X"A8",X"A8",X"AA",X"A8",X"AA",X"88",X"28",X"00",X"22",X"A8",X"AA",X"AA",X"AA",X"A2",X"82",
		X"00",X"02",X"AA",X"A8",X"AA",X"AA",X"88",X"AA",X"00",X"0A",X"AA",X"AA",X"AA",X"8A",X"AA",X"AA",
		X"00",X"A8",X"AA",X"2A",X"A8",X"AA",X"82",X"AA",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"88",X"AA",
		X"08",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"0A",X"A2",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"2A",X"AA",X"10",X"00",X"00",X"00",X"28",X"02",X"22",X"AA",X"A4",X"02",X"08",X"8A",X"A0",X"02",
		X"0A",X"AA",X"A0",X"00",X"A0",X"00",X"00",X"0A",X"AA",X"8A",X"A0",X"2A",X"00",X"00",X"00",X"2A",
		X"AA",X"AA",X"A2",X"AA",X"00",X"00",X"0A",X"AA",X"8A",X"AA",X"AA",X"A0",X"00",X"00",X"22",X"AA",
		X"AA",X"8A",X"A0",X"A2",X"20",X"6A",X"AA",X"AA",X"AA",X"A8",X"AA",X"82",X"00",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"8A",X"AA",X"0A",X"AA",X"8A",X"AA",X"AA",X"AA",X"AA",X"AA",X"8A",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"0A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"2A",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"28",X"2A",X"AA",X"A8",X"AA",X"AA",X"AA",X"A8",X"AA",X"AA",X"AA",X"AA",
		X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"2A",X"80",X"00",X"00",X"00",X"AA",X"00",X"00",X"AA",X"AA",X"00",X"80",X"02",X"80",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"82",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"A2",X"A0",X"00",X"00",X"00",
		X"A8",X"AA",X"A2",X"28",X"AA",X"00",X"20",X"00",X"AA",X"8A",X"82",X"A2",X"88",X"00",X"00",X"00",
		X"A8",X"8A",X"AA",X"AA",X"A0",X"2A",X"80",X"00",X"A8",X"8A",X"A2",X"AA",X"8A",X"A8",X"A0",X"00",
		X"AA",X"8A",X"A8",X"AA",X"82",X"2A",X"28",X"20",X"AA",X"2A",X"AA",X"A2",X"0A",X"AA",X"AA",X"00",
		X"AA",X"AA",X"AA",X"AA",X"08",X"8A",X"A2",X"00",X"AA",X"2A",X"0A",X"AA",X"02",X"AA",X"AA",X"80",
		X"AA",X"2A",X"AA",X"AA",X"02",X"8A",X"2A",X"A0",X"8A",X"22",X"A0",X"AA",X"0A",X"AA",X"2A",X"A8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"82",X"A8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"A0",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"0A",X"01",X"10",X"A8",X"A2",X"28",X"80",X"00",X"00",X"04",X"00",X"8A",X"AA",X"AA",X"20",
		X"00",X"00",X"00",X"18",X"88",X"A0",X"82",X"00",X"00",X"00",X"00",X"12",X"AA",X"AA",X"00",X"00",
		X"00",X"08",X"00",X"08",X"88",X"02",X"80",X"00",X"00",X"28",X"00",X"02",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"28",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"02",X"20",X"02",
		X"00",X"00",X"00",X"00",X"28",X"00",X"00",X"2A",X"00",X"00",X"00",X"00",X"28",X"08",X"20",X"80",
		X"00",X"00",X"00",X"01",X"0A",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"0A",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"40",X"28",X"00",X"02",X"00",X"00",X"00",X"20",X"02",X"80",X"01",X"80",
		X"00",X"00",X"00",X"08",X"00",X"00",X"08",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"00",X"00",X"02",X"28",X"95",X"55",X"55",X"A2",X"00",X"00",X"00",X"68",X"95",X"55",X"55",
		X"AA",X"00",X"80",X"01",X"28",X"95",X"55",X"55",X"20",X"80",X"A0",X"00",X"28",X"95",X"55",X"55",
		X"88",X"82",X"28",X"80",X"68",X"95",X"55",X"55",X"00",X"02",X"A8",X"20",X"68",X"A1",X"55",X"55",
		X"00",X"00",X"82",X"00",X"08",X"A0",X"55",X"55",X"00",X"00",X"00",X"80",X"0A",X"A0",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"A0",X"15",X"55",X"00",X"00",X"00",X"00",X"02",X"20",X"05",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"8A",X"AA",X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",X"0A",X"AA",
		X"2A",X"AA",X"AA",X"AA",X"AA",X"A8",X"AA",X"AA",X"0A",X"AA",X"AA",X"AA",X"AA",X"A8",X"2A",X"AA",
		X"02",X"AA",X"AA",X"AA",X"AA",X"A2",X"AA",X"A8",X"00",X"AA",X"AA",X"AA",X"AA",X"A8",X"2A",X"AA",
		X"00",X"02",X"AA",X"AA",X"AA",X"A8",X"AA",X"AA",X"00",X"00",X"AA",X"AA",X"AA",X"A2",X"AA",X"AA",
		X"00",X"00",X"0A",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"0A",X"AA",X"AA",X"A2",X"AA",X"80",
		X"00",X"00",X"AA",X"A0",X"0A",X"8A",X"AA",X"80",X"00",X"00",X"28",X"00",X"2A",X"AA",X"A8",X"00",
		X"00",X"00",X"00",X"00",X"02",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"A0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"88",X"AA",X"AA",X"80",
		X"2A",X"AA",X"AA",X"AA",X"02",X"AA",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"8A",X"A8",X"80",X"00",
		X"AA",X"AA",X"AA",X"AA",X"0A",X"80",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"40",X"00",X"00",
		X"8A",X"AA",X"AA",X"AA",X"A9",X"00",X"00",X"02",X"00",X"02",X"AA",X"AA",X"A0",X"00",X"00",X"20",
		X"00",X"00",X"2A",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"A4",X"00",X"00",X"00",X"00",
		X"00",X"02",X"AA",X"96",X"00",X"00",X"00",X"00",X"00",X"08",X"2A",X"98",X"00",X"00",X"00",X"00",
		X"00",X"80",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"88",X"AA",X"AA",X"AA",X"0A",X"A2",X"AA",X"AA",X"82",X"AA",X"AA",X"A8",
		X"00",X"AA",X"AA",X"AA",X"0A",X"AA",X"2A",X"A8",X"02",X"AA",X"AA",X"A8",X"28",X"AA",X"AA",X"00",
		X"80",X"AA",X"AA",X"AA",X"8A",X"AA",X"AA",X"00",X"08",X"AA",X"AA",X"AA",X"28",X"AA",X"AA",X"00",
		X"80",X"AA",X"AA",X"AA",X"2A",X"AA",X"A8",X"00",X"0A",X"AA",X"AA",X"A8",X"8A",X"AA",X"A8",X"00",
		X"00",X"02",X"AA",X"AA",X"2A",X"AA",X"00",X"00",X"00",X"02",X"A2",X"A8",X"2A",X"00",X"00",X"00",
		X"00",X"02",X"00",X"A0",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"2A",X"A2",X"00",X"00",X"00",
		X"00",X"00",X"20",X"AA",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"80",X"00",X"00",X"00",
		X"00",X"00",X"28",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A2",X"20",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",
		X"00",X"00",X"01",X"00",X"00",X"40",X"01",X"60",X"00",X"04",X"01",X"00",X"01",X"00",X"01",X"68",
		X"00",X"04",X"04",X"00",X"00",X"0A",X"84",X"A8",X"00",X"14",X"00",X"88",X"00",X"AA",X"00",X"A2",
		X"00",X"10",X"00",X"AA",X"AA",X"88",X"04",X"A2",X"05",X"00",X"A8",X"00",X"02",X"80",X"00",X"2A",
		X"01",X"00",X"A8",X"00",X"00",X"00",X"00",X"0A",X"45",X"00",X"08",X"00",X"00",X"00",X"00",X"02",
		X"28",X"02",X"A8",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",
		X"50",X"00",X"02",X"00",X"00",X"00",X"06",X"00",X"55",X"40",X"00",X"00",X"00",X"00",X"02",X"00",
		X"80",X"55",X"55",X"50",X"00",X"00",X"02",X"00",X"20",X"09",X"55",X"55",X"55",X"50",X"02",X"80",
		X"AA",X"00",X"00",X"00",X"02",X"55",X"02",X"80",X"20",X"00",X"00",X"00",X"00",X"00",X"09",X"A8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"A9",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"98",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"40",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"11",X"80",X"00",X"60",X"00",X"00",X"00",
		X"00",X"0A",X"A8",X"20",X"20",X"00",X"00",X"00",X"01",X"22",X"02",X"00",X"48",X"00",X"00",X"00",
		X"00",X"0A",X"80",X"00",X"18",X"00",X"00",X"00",X"00",X"28",X"00",X"00",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"48",X"00",X"00",X"00",
		X"00",X"00",X"00",X"20",X"08",X"00",X"00",X"00",X"00",X"00",X"40",X"80",X"18",X"00",X"00",X"00",
		X"00",X"00",X"80",X"10",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"28",X"00",X"00",X"00",
		X"00",X"40",X"1A",X"90",X"19",X"00",X"50",X"26",X"00",X"40",X"6A",X"90",X"19",X"00",X"50",X"26",
		X"00",X"80",X"6A",X"90",X"19",X"00",X"50",X"25",X"00",X"80",X"6A",X"90",X"19",X"02",X"50",X"01",
		X"00",X"80",X"6A",X"90",X"19",X"02",X"50",X"00",X"00",X"80",X"6A",X"94",X"19",X"02",X"50",X"00",
		X"80",X"80",X"6A",X"A4",X"19",X"02",X"50",X"00",X"84",X"91",X"6A",X"A5",X"19",X"46",X"51",X"11",
		X"95",X"95",X"5A",X"A5",X"59",X"56",X"55",X"6A",X"95",X"95",X"5A",X"A5",X"59",X"56",X"55",X"6A",
		X"95",X"95",X"5A",X"A5",X"59",X"56",X"55",X"65",X"95",X"95",X"55",X"55",X"59",X"56",X"55",X"66",
		X"95",X"65",X"55",X"55",X"59",X"56",X"55",X"9A",X"95",X"69",X"55",X"55",X"55",X"56",X"55",X"9A",
		X"55",X"5A",X"55",X"55",X"55",X"55",X"55",X"9A",X"55",X"5A",X"AA",X"AA",X"A5",X"AA",X"55",X"9A",
		X"55",X"56",X"AA",X"AA",X"A5",X"AA",X"6A",X"9A",X"5A",X"A5",X"55",X"55",X"55",X"6A",X"AA",X"9A",
		X"A9",X"56",X"AA",X"AA",X"AA",X"95",X"55",X"5A",X"56",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"A8",X"00",X"00",X"00",X"00",X"00",X"2A",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"15",X"55",X"55",X"10",X"00",X"00",X"00",X"05",X"55",X"55",X"55",X"55",X"40",X"00",
		X"00",X"55",X"AA",X"AA",X"AA",X"A9",X"54",X"00",X"01",X"6A",X"AA",X"AA",X"AA",X"AA",X"95",X"00",
		X"06",X"AA",X"AA",X"AA",X"AA",X"AA",X"A9",X"40",X"0A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"40",
		X"0A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"80",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",
		X"00",X"0A",X"AA",X"AA",X"AA",X"AA",X"A0",X"A0",X"00",X"00",X"AA",X"A8",X"8A",X"80",X"00",X"00",
		X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"15",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"05",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"A5",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"95",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"15",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"A5",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"0A",X"A9",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"09",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"A5",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"29",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"60",X"88",X"00",X"02",X"00",X"00",X"00",X"54",X"15",X"55",
		X"00",X"00",X"00",X"00",X"55",X"15",X"55",X"55",X"00",X"02",X"AA",X"A9",X"55",X"55",X"55",X"55",
		X"0A",X"80",X"15",X"55",X"55",X"55",X"55",X"65",X"01",X"55",X"59",X"56",X"59",X"55",X"A6",X"59",
		X"A5",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"65",X"56",X"65",X"65",X"65",X"59",X"95",
		X"55",X"55",X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"55",X"55",X"55",X"55",X"55",
		X"56",X"55",X"56",X"55",X"95",X"56",X"55",X"40",X"95",X"65",X"55",X"59",X"55",X"55",X"55",X"50",
		X"00",X"00",X"00",X"00",X"00",X"00",X"95",X"55",X"00",X"00",X"00",X"01",X"48",X"55",X"65",X"50",
		X"02",X"95",X"55",X"55",X"56",X"56",X"55",X"40",X"09",X"55",X"5A",X"56",X"65",X"65",X"94",X"00",
		X"95",X"55",X"55",X"65",X"95",X"55",X"00",X"00",X"55",X"55",X"95",X"55",X"54",X"00",X"00",X"00",
		X"55",X"95",X"55",X"00",X"00",X"00",X"00",X"00",X"95",X"65",X"54",X"00",X"00",X"00",X"00",X"00",
		X"59",X"55",X"41",X"00",X"00",X"00",X"00",X"00",X"95",X"54",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"51",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"28",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"28",X"00",X"00",X"00",
		X"02",X"80",X"00",X"00",X"28",X"04",X"80",X"00",X"00",X"00",X"00",X"01",X"2A",X"0A",X"00",X"00",
		X"00",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"AA",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"2A",X"80",X"00",X"00",X"00",X"00",X"00",X"04",X"2A",X"20",X"00",X"00",
		X"00",X"00",X"00",X"80",X"0A",X"20",X"00",X"00",X"00",X"00",X"04",X"00",X"8A",X"A0",X"00",X"00",
		X"00",X"00",X"02",X"00",X"20",X"88",X"00",X"00",X"00",X"00",X"20",X"00",X"A8",X"80",X"00",X"00",
		X"00",X"00",X"00",X"02",X"A8",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"28",X"80",X"00",X"00",
		X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A8",X"3F",X"FA",X"AA",X"AA",X"AB",X"C0",X"AA",X"83",X"FE",X"AA",X"AA",X"AA",X"AA",X"BC",X"0A",
		X"0F",X"EA",X"A5",X"55",X"55",X"AA",X"AB",X"02",X"3E",X"A9",X"55",X"55",X"55",X"56",X"AA",X"C0",
		X"FA",X"95",X"55",X"55",X"55",X"55",X"5A",X"B0",X"E9",X"55",X"55",X"55",X"55",X"55",X"55",X"AC",
		X"E9",X"55",X"55",X"55",X"55",X"55",X"55",X"AC",X"A5",X"55",X"55",X"55",X"55",X"55",X"55",X"6B",
		X"A5",X"55",X"55",X"55",X"55",X"55",X"55",X"6B",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"6B",
		X"D5",X"55",X"55",X"55",X"55",X"55",X"55",X"5B",X"E5",X"55",X"55",X"55",X"55",X"55",X"55",X"7F",
		X"F9",X"55",X"55",X"55",X"55",X"55",X"55",X"FE",X"BF",X"95",X"55",X"55",X"55",X"55",X"57",X"FA",
		X"2F",X"F9",X"55",X"55",X"55",X"56",X"FF",X"E8",X"0A",X"FF",X"ED",X"55",X"57",X"BF",X"FE",X"A0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"11",X"55",X"55",X"10",X"00",X"00",X"00",X"05",X"55",X"55",X"55",X"55",X"40",X"00",
		X"00",X"55",X"AA",X"AA",X"AA",X"A9",X"54",X"00",X"05",X"6A",X"AA",X"AA",X"AA",X"AA",X"95",X"40",
		X"16",X"AA",X"AA",X"AA",X"AA",X"AA",X"A9",X"50",X"1A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"54",
		X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"94",X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"90",
		X"0A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"02",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",
		X"00",X"0A",X"AA",X"AA",X"AA",X"AA",X"80",X"00",X"00",X"00",X"2A",X"AA",X"AA",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"20",X"00",X"02",X"00",X"00",X"00",X"00",X"02",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"00",X"02",X"00",X"00",
		X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"A0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2A",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0A",X"AA",X"96",X"00",X"00",X"00",X"00",X"00",X"15",X"55",X"65",
		X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"00",X"00",X"00",X"00",X"08",X"02",X"01",X"56",
		X"00",X"00",X"00",X"00",X"22",X"08",X"25",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"15",X"55",
		X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"95",X"55",X"9A",X"55",X"55",X"95",X"55",X"50",X"59",X"55",X"55",X"55",X"55",X"54",X"44",X"00",
		X"55",X"59",X"55",X"55",X"55",X"55",X"64",X"00",X"59",X"65",X"95",X"56",X"55",X"55",X"58",X"00",
		X"55",X"55",X"56",X"55",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"90",
		X"55",X"55",X"55",X"55",X"55",X"50",X"00",X"00",X"15",X"55",X"40",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"C0",X"00",X"00",X"3F",
		X"00",X"00",X"0F",X"EB",X"FF",X"00",X"03",X"FF",X"00",X"00",X"FE",X"BF",X"FF",X"F0",X"3F",X"FF",
		X"00",X"0F",X"EB",X"FF",X"FF",X"AB",X"FF",X"FE",X"00",X"FE",X"BF",X"FF",X"FE",X"AF",X"FE",X"FF",
		X"0F",X"EB",X"FF",X"FF",X"FA",X"BF",X"FA",X"FF",X"3E",X"BF",X"FF",X"FF",X"EA",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E0",
		X"2F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"80",X"0B",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"00",
		X"02",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"00",X"0F",X"FE",X"AA",X"AA",X"AA",X"AB",X"FF",X"00",
		X"FF",X"BF",X"AA",X"AA",X"AA",X"AF",X"EF",X"F0",X"FF",X"EF",X"EA",X"AA",X"AA",X"BF",X"BF",X"FF",
		X"FF",X"FB",X"EA",X"AA",X"AA",X"BE",X"FF",X"FF",X"BF",X"FE",X"FF",X"FF",X"FF",X"FB",X"FF",X"FB",
		X"BF",X"FE",X"AA",X"AA",X"AA",X"AB",X"FF",X"FB",X"FF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AF",X"FF",
		X"FA",X"AA",X"AF",X"FF",X"FF",X"AA",X"AA",X"FF",X"AA",X"8B",X"FF",X"EE",X"FF",X"FE",X"0A",X"AF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"3F",X"F0",X"00",X"00",X"00",
		X"FC",X"00",X"0F",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"C0",X"FF",X"FF",X"FF",X"F0",X"00",X"00",
		X"FF",X"FE",X"BF",X"FF",X"FF",X"FF",X"00",X"00",X"FE",X"FF",X"AF",X"FF",X"FF",X"FF",X"F0",X"00",
		X"FE",X"FF",X"EB",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FA",X"FF",X"FF",X"FF",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"55",X"08",X"AA",X"95",X"00",X"00",
		X"00",X"01",X"2A",X"2A",X"AA",X"A9",X"00",X"00",X"00",X"00",X"A8",X"AA",X"AA",X"00",X"00",X"00",
		X"00",X"00",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0A",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"A8",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"20",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"20",X"00",X"00",X"00",X"80",X"00",X"00",X"04",X"20",X"00",X"00",X"00",X"00",
		X"00",X"00",X"40",X"20",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"28",X"02",X"00",X"00",X"08",
		X"00",X"00",X"00",X"AA",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"1A",X"00",X"20",X"00",X"00",
		X"00",X"00",X"00",X"12",X"20",X"80",X"00",X"00",X"00",X"A0",X"00",X"46",X"00",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"28",X"00",X"00",X"00",
		X"00",X"08",X"00",X"02",X"0A",X"80",X"00",X"00",X"00",X"0A",X"00",X"0A",X"AA",X"00",X"80",X"00",
		X"00",X"00",X"00",X"08",X"8A",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"8A",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"2A",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"20",X"40",X"00",X"00",X"00",X"00",X"00",
		X"20",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"8A",X"04",X"02",X"00",X"00",X"00",X"00",
		X"0A",X"28",X"68",X"00",X"A0",X"00",X"00",X"00",X"08",X"81",X"A8",X"22",X"80",X"00",X"00",X"00",
		X"02",X"A4",X"2A",X"2A",X"10",X"00",X"00",X"00",X"02",X"88",X"88",X"21",X"00",X"00",X"00",X"00",
		X"02",X"A0",X"AA",X"A9",X"62",X"28",X"00",X"00",X"02",X"80",X"A8",X"A5",X"20",X"A8",X"00",X"00",
		X"82",X"62",X"88",X"80",X"A2",X"AA",X"02",X"20",X"02",X"02",X"88",X"81",X"88",X"8A",X"8A",X"00",
		X"02",X"12",X"22",X"84",X"8A",X"82",X"A2",X"00",X"AA",X"0A",X"AA",X"00",X"8A",X"82",X"08",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"08",X"00",X"00",X"00",
		X"00",X"00",X"60",X"00",X"00",X"88",X"20",X"00",X"00",X"00",X"80",X"00",X"00",X"02",X"02",X"AA",
		X"04",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"18",X"00",X"00",X"00",X"00",X"2A",X"0A",X"AA",
		X"00",X"00",X"08",X"00",X"8A",X"22",X"0A",X"AA",X"00",X"00",X"00",X"02",X"22",X"A8",X"0A",X"AA",
		X"00",X"00",X"A0",X"2A",X"2A",X"0A",X"02",X"AA",X"00",X"2A",X"A2",X"A0",X"AA",X"8A",X"0A",X"AA",
		X"0A",X"A0",X"A2",X"28",X"A2",X"88",X"02",X"AA",X"AA",X"8A",X"22",X"82",X"22",X"AA",X"22",X"AA",
		X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"14",X"00",X"80",X"00",X"00",X"00",X"00",
		X"00",X"18",X"88",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"AA",X"00",X"00",X"0A",X"A0",
		X"00",X"00",X"00",X"22",X"AA",X"AA",X"AA",X"A0",X"00",X"00",X"00",X"A2",X"AA",X"AA",X"A0",X"A0",
		X"2A",X"8A",X"A2",X"A2",X"AA",X"AA",X"A2",X"A0",X"8A",X"A2",X"AA",X"80",X"AA",X"AA",X"A0",X"A0",
		X"88",X"22",X"A2",X"20",X"AA",X"AA",X"8A",X"A0",X"A2",X"82",X"AA",X"20",X"AA",X"AA",X"0A",X"A0",
		X"AA",X"80",X"AA",X"82",X"AA",X"AA",X"2A",X"A3",X"88",X"08",X"AA",X"82",X"AA",X"A8",X"2A",X"A3",
		X"A0",X"82",X"AA",X"82",X"AA",X"AA",X"2A",X"A2",X"A8",X"28",X"AA",X"A0",X"AA",X"A8",X"2A",X"A2",
		X"AA",X"A0",X"AA",X"A8",X"2A",X"AA",X"0A",X"A2",X"8A",X"A8",X"AA",X"A8",X"2A",X"AA",X"2A",X"A0",
		X"2B",X"FF",X"FF",X"FF",X"AB",X"FF",X"FF",X"FA",X"2A",X"AB",X"FF",X"FF",X"BF",X"FF",X"FF",X"EA",
		X"2A",X"AA",X"AA",X"BE",X"AA",X"AF",X"FF",X"A8",X"0A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AE",X"A0",
		X"00",X"0A",X"AA",X"AA",X"BF",X"EA",X"AA",X"80",X"00",X"00",X"00",X"2A",X"FF",X"FF",X"FA",X"03",
		X"00",X"00",X"00",X"02",X"FE",X"FF",X"EA",X"03",X"00",X"00",X"00",X"02",X"FF",X"AB",X"E8",X"0F",
		X"00",X"00",X"00",X"02",X"FA",X"FF",X"E8",X"0F",X"00",X"00",X"FF",X"FA",X"FF",X"AB",X"E8",X"0F",
		X"FF",X"FF",X"EA",X"BA",X"FE",X"FF",X"E8",X"03",X"EA",X"AA",X"BF",X"FA",X"FF",X"FA",X"BC",X"03",
		X"FF",X"FF",X"FF",X"FA",X"BE",X"AB",X"E8",X"02",X"BF",X"FF",X"FF",X"FE",X"AA",X"FE",X"AC",X"02",
		X"AF",X"FF",X"FF",X"FE",X"BF",X"AA",X"FF",X"00",X"AB",X"FF",X"FF",X"FF",X"AA",X"BF",X"FF",X"C0",
		X"A8",X"3F",X"FA",X"AA",X"AA",X"FF",X"C0",X"AA",X"83",X"FE",X"AA",X"AA",X"AA",X"AB",X"FC",X"0A",
		X"0F",X"EA",X"A0",X"00",X"00",X"AA",X"BF",X"02",X"3E",X"A8",X"00",X"00",X"00",X"02",X"AB",X"C0",
		X"FA",X"80",X"00",X"00",X"00",X"00",X"2A",X"F0",X"E8",X"00",X"00",X"00",X"00",X"00",X"02",X"BC",
		X"E8",X"00",X"00",X"00",X"00",X"00",X"02",X"BC",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"AF",
		X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"AF",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"AF",
		X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",
		X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"FA",X"BF",X"80",X"00",X"00",X"00",X"00",X"0F",X"E8",
		X"AF",X"F8",X"00",X"00",X"00",X"02",X"FF",X"A0",X"2A",X"FF",X"EC",X"00",X"03",X"BF",X"FA",X"80",
		X"FF",X"FF",X"FE",X"BF",X"FF",X"FF",X"FE",X"00",X"BF",X"FF",X"FF",X"AF",X"FF",X"FE",X"AA",X"00",
		X"AF",X"FF",X"AA",X"AF",X"EA",X"AA",X"A8",X"00",X"AB",X"AA",X"AA",X"AA",X"AA",X"A8",X"00",X"00",
		X"2A",X"AA",X"BF",X"EA",X"80",X"00",X"00",X"00",X"0A",X"FF",X"FF",X"FA",X"00",X"00",X"00",X"00",
		X"0A",X"BF",X"FF",X"FA",X"00",X"00",X"00",X"00",X"02",X"BF",X"EF",X"FA",X"00",X"00",X"00",X"00",
		X"02",X"BF",X"BB",X"FA",X"00",X"00",X"00",X"00",X"02",X"BF",X"EF",X"FA",X"FF",X"F0",X"00",X"00",
		X"02",X"AF",X"FF",X"FA",X"FF",X"FF",X"FF",X"FC",X"02",X"FA",X"FF",X"FA",X"FF",X"FF",X"FF",X"F8",
		X"02",X"AF",X"AB",X"EA",X"FF",X"FF",X"FF",X"F8",X"03",X"FA",X"FE",X"AA",X"FF",X"FF",X"FF",X"E8",
		X"0F",X"FF",X"AB",X"FB",X"FF",X"FF",X"FF",X"A0",X"3F",X"FF",X"FA",X"AB",X"FF",X"FF",X"FE",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",
		X"02",X"00",X"08",X"00",X"08",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"00",X"20",X"08",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"08",
		X"00",X"80",X"20",X"08",X"02",X"00",X"00",X"00",X"00",X"00",X"82",X"00",X"20",X"02",X"00",X"00",
		X"02",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"28",X"20",X"00",X"20",X"20",X"00",X"20",X"00",
		X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"08",X"00",X"20",
		X"00",X"00",X"80",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"20",X"2A",X"00",X"00",X"08",X"00",X"08",X"08",X"00",X"AA",X"20",X"00",X"00",
		X"00",X"20",X"20",X"0A",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A8",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"22",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"20",X"00",X"02",
		X"00",X"00",X"00",X"00",X"02",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"08",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",
		X"00",X"02",X"80",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A8",X"8A",X"2A",X"00",X"2A",X"80",X"08",X"00",X"80",X"88",X"22",X"02",X"82",X"80",X"28",X"00",
		X"88",X"2A",X"28",X"02",X"22",X"88",X"28",X"AA",X"00",X"28",X"88",X"02",X"A2",X"A8",X"20",X"2A",
		X"08",X"AA",X"A0",X"00",X"88",X"A0",X"22",X"AA",X"08",X"A8",X"A0",X"02",X"08",X"A0",X"A0",X"0A",
		X"02",X"AA",X"A0",X"08",X"28",X"00",X"82",X"2A",X"0A",X"AA",X"A0",X"01",X"20",X"02",X"92",X"0A",
		X"82",X"AA",X"80",X"04",X"AA",X"02",X"00",X"1A",X"0A",X"AA",X"00",X"06",X"A8",X"0A",X"40",X"12",
		X"2A",X"A8",X"00",X"02",X"22",X"08",X"40",X"22",X"AA",X"AA",X"00",X"08",X"A8",X"09",X"08",X"22",
		X"AA",X"AA",X"00",X"02",X"80",X"24",X"0A",X"80",X"0A",X"AA",X"00",X"AA",X"80",X"24",X"08",X"88",
		X"00",X"A8",X"00",X"02",X"20",X"20",X"28",X"AA",X"00",X"08",X"02",X"AA",X"02",X"A2",X"2A",X"AA",
		X"AA",X"82",X"A8",X"88",X"8A",X"8A",X"0A",X"AA",X"A2",X"28",X"8A",X"02",X"22",X"A8",X"A2",X"AA",
		X"A8",X"22",X"22",X"82",X"8A",X"2A",X"82",X"AA",X"AA",X"AA",X"8A",X"20",X"A2",X"2A",X"82",X"AA",
		X"A8",X"A8",X"A8",X"A0",X"AA",X"AA",X"82",X"AA",X"A2",X"22",X"A2",X"A0",X"A2",X"2A",X"0A",X"AA",
		X"A8",X"A8",X"A2",X"28",X"22",X"2A",X"02",X"AA",X"A8",X"2A",X"A2",X"A8",X"2A",X"2A",X"22",X"AA",
		X"A8",X"AA",X"A2",X"A0",X"AA",X"2A",X"0A",X"AA",X"A8",X"AA",X"2A",X"82",X"2A",X"AA",X"2A",X"AA",
		X"A0",X"AA",X"AA",X"02",X"0A",X"AA",X"88",X"00",X"A2",X"A8",X"A8",X"8A",X"8A",X"80",X"00",X"00",
		X"AA",X"AA",X"AA",X"80",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"A8",X"00",X"00",X"00",X"00",X"00",X"00",X"A2",X"80",X"80",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"A2",X"2A",X"AA",X"2A",X"A0",X"AA",X"AA",X"AA",X"A2",X"2A",X"A8",X"0A",X"A0",
		X"AA",X"AA",X"AA",X"A8",X"AA",X"A8",X"2A",X"A0",X"AA",X"AA",X"AA",X"A8",X"2A",X"AA",X"0A",X"A0",
		X"AA",X"AA",X"AA",X"AA",X"2A",X"AA",X"2A",X"A0",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"0A",X"A0",
		X"AA",X"AA",X"AA",X"AA",X"A2",X"AA",X"0A",X"A0",X"AA",X"AA",X"AA",X"AA",X"A2",X"A8",X"0A",X"A0",
		X"AA",X"AA",X"AA",X"8A",X"AA",X"AA",X"2A",X"A0",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"2A",X"A2",
		X"0A",X"AA",X"AA",X"AA",X"AA",X"A8",X"2A",X"A2",X"00",X"00",X"0A",X"A8",X"8A",X"AA",X"2A",X"08",
		X"00",X"00",X"0A",X"AA",X"22",X"AA",X"2A",X"A8",X"00",X"00",X"00",X"00",X"88",X"AA",X"2A",X"80",
		X"00",X"00",X"00",X"00",X"02",X"28",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"2B",X"FF",X"FF",X"FF",X"EB",X"FF",X"EF",X"F0",X"2A",X"FF",X"FF",X"FF",X"AB",X"FF",X"AF",X"FF",
		X"0A",X"BF",X"FF",X"EA",X"AA",X"BF",X"FF",X"FF",X"02",X"AF",X"FE",X"AA",X"AA",X"AF",X"FF",X"EF",
		X"00",X"AB",X"EA",X"AA",X"02",X"AB",X"FF",X"AF",X"00",X"2A",X"AA",X"80",X"00",X"AA",X"FF",X"FF",
		X"00",X"0A",X"A8",X"00",X"00",X"2A",X"AF",X"FF",X"00",X"02",X"80",X"00",X"00",X"0A",X"AA",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"02",X"AA",X"FB",X"00",X"00",X"00",X"00",X"00",X"00",X"2A",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"AF",X"FA",X"FF",X"FE",X"FF",X"AA",X"00",X"00",X"AA",X"AF",X"FA",X"FF",X"AA",X"A0",X"AF",
		X"FA",X"8A",X"AA",X"AA",X"AA",X"AA",X"0A",X"BF",X"FF",X"A8",X"8A",X"AA",X"AA",X"22",X"AF",X"FF",
		X"FA",X"FE",X"AA",X"AA",X"AA",X"AB",X"FA",X"FF",X"EF",X"FE",X"FF",X"FF",X"FF",X"FB",X"FF",X"BF",
		X"BF",X"FB",X"FA",X"AA",X"AA",X"FE",X"FF",X"EF",X"FF",X"EF",X"EA",X"AA",X"AA",X"BF",X"BF",X"FB",
		X"FA",X"BF",X"AF",X"FF",X"FF",X"AF",X"EA",X"FE",X"BB",X"FE",X"AA",X"AA",X"AA",X"AB",X"FE",X"FA",
		X"AF",X"FA",X"AA",X"AA",X"AA",X"AA",X"FF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"00",X"2A",X"AA",X"AA",X"AA",X"AA",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FA",X"FE",X"AF",X"FF",X"FF",X"FE",X"80",X"FF",X"FA",X"FA",X"AF",X"FF",X"FF",X"FA",X"00",
		X"FF",X"FF",X"EA",X"0A",X"FF",X"FF",X"E8",X"00",X"FA",X"FF",X"AA",X"02",X"AB",X"FF",X"A0",X"00",
		X"FA",X"FE",X"A8",X"00",X"0A",X"AE",X"80",X"00",X"FF",X"FA",X"80",X"00",X"00",X"AA",X"00",X"00",
		X"FF",X"AA",X"80",X"00",X"00",X"00",X"00",X"00",X"FA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FA",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"09",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"2A",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"2A",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"2A",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"29",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"2A",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"2A",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"AA",X"95",X"55",X"55",
		X"00",X"00",X"00",X"00",X"AA",X"95",X"55",X"55",X"00",X"00",X"00",X"02",X"AA",X"95",X"55",X"55",
		X"00",X"00",X"00",X"02",X"AA",X"A5",X"55",X"55",X"00",X"00",X"00",X"0A",X"AA",X"A5",X"55",X"55",
		X"00",X"00",X"00",X"00",X"AA",X"A5",X"55",X"55",X"00",X"00",X"00",X"2A",X"AA",X"95",X"55",X"55",
		X"00",X"00",X"00",X"AA",X"AA",X"95",X"55",X"55",X"00",X"00",X"0A",X"AA",X"AA",X"A9",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"05",X"55",X"55",X"55",X"55",X"5A",
		X"00",X"00",X"14",X"00",X"00",X"00",X"0A",X"68",X"50",X"00",X"10",X"00",X"00",X"00",X"0A",X"60",
		X"14",X"00",X"10",X"00",X"00",X"00",X"29",X"A0",X"04",X"00",X"10",X"00",X"00",X"00",X"29",X"80",
		X"A9",X"00",X"10",X"00",X"00",X"00",X"29",X"80",X"AA",X"40",X"90",X"00",X"AA",X"80",X"A6",X"00",
		X"2A",X"40",X"94",X"00",X"95",X"40",X"A6",X"00",X"2A",X"50",X"A4",X"00",X"9A",X"40",X"A6",X"00",
		X"6A",X"10",X"A5",X"00",X"26",X"40",X"98",X"00",X"AA",X"24",X"A9",X"00",X"26",X"40",X"98",X"00",
		X"A8",X"24",X"AA",X"40",X"0A",X"00",X"98",X"00",X"90",X"29",X"AA",X"40",X"0A",X"00",X"98",X"00",
		X"90",X"09",X"2A",X"90",X"02",X"00",X"98",X"00",X"A4",X"09",X"2A",X"90",X"02",X"00",X"98",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"15",X"55",X"54",
		X"55",X"40",X"00",X"15",X"05",X"00",X"24",X"05",X"01",X"00",X"00",X"50",X"05",X"00",X"24",X"00",
		X"01",X"00",X"01",X"40",X"19",X"00",X"14",X"00",X"04",X"00",X"04",X"00",X"1A",X"00",X"98",X"00",
		X"AA",X"2A",X"A2",X"AA",X"9A",X"8A",X"AA",X"AA",X"AA",X"2A",X"AA",X"AA",X"9A",X"8A",X"AA",X"8A",
		X"AA",X"2A",X"AA",X"A0",X"2A",X"8A",X"AA",X"80",X"AA",X"2A",X"A8",X"A0",X"AA",X"8A",X"AA",X"88",
		X"AA",X"2A",X"A8",X"A0",X"AA",X"8A",X"AA",X"89",X"0A",X"2A",X"A8",X"A2",X"AA",X"A8",X"66",X"AA",
		X"0A",X"5A",X"A8",X"A2",X"98",X"A8",X"64",X"8A",X"00",X"40",X"05",X"90",X"19",X"00",X"64",X"09",
		X"00",X"40",X"06",X"90",X"19",X"00",X"50",X"09",X"00",X"40",X"1A",X"90",X"19",X"00",X"50",X"26",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"94",X"00",X"00",X"00",X"04",X"00",X"00",
		X"0A",X"50",X"00",X"00",X"00",X"18",X"00",X"00",X"29",X"80",X"00",X"00",X"00",X"18",X"00",X"00",
		X"26",X"80",X"00",X"00",X"00",X"18",X"00",X"2A",X"26",X"80",X"00",X"00",X"00",X"1A",X"00",X"2A",
		X"26",X"80",X"00",X"00",X"00",X"1A",X"AA",X"AA",X"26",X"80",X"02",X"AA",X"80",X"16",X"55",X"2A",
		X"26",X"A0",X"01",X"55",X"A0",X"06",X"00",X"2A",X"26",X"A0",X"00",X"1A",X"60",X"06",X"00",X"A8",
		X"09",X"A8",X"00",X"1A",X"60",X"06",X"00",X"A8",X"02",X"6A",X"00",X"05",X"60",X"06",X"80",X"00",
		X"00",X"9A",X"80",X"00",X"68",X"06",X"80",X"00",X"00",X"26",X"A0",X"00",X"68",X"05",X"80",X"2A",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"80",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"80",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"80",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A2",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"00",
		X"0A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"80",X"2A",X"A8",X"0A",X"AA",X"00",X"8A",X"00",X"00",
		X"A0",X"82",X"A0",X"00",X"0A",X"88",X"20",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"12",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"20",X"28",X"48",X"00",X"00",X"00",X"00",X"00",X"A0",X"28",X"18",X"00",X"00",X"00",X"00",
		X"00",X"80",X"A8",X"18",X"00",X"00",X"00",X"00",X"02",X"A0",X"A8",X"4A",X"00",X"00",X"00",X"00",
		X"00",X"A0",X"28",X"1A",X"00",X"00",X"00",X"00",X"02",X"20",X"20",X"02",X"00",X"00",X"00",X"00",
		X"00",X"2A",X"28",X"46",X"00",X"00",X"00",X"00",X"00",X"20",X"25",X"01",X"80",X"00",X"00",X"00",
		X"00",X"2A",X"21",X"10",X"80",X"00",X"00",X"00",X"00",X"2A",X"A4",X"40",X"80",X"00",X"00",X"00",
		X"08",X"8A",X"15",X"00",X"80",X"00",X"00",X"00",X"A2",X"2A",X"11",X"00",X"20",X"00",X"00",X"00",
		X"22",X"0A",X"04",X"10",X"20",X"00",X"00",X"00",X"08",X"22",X"00",X"40",X"20",X"00",X"00",X"00",
		X"00",X"08",X"80",X"40",X"20",X"00",X"00",X"00",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"52",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"1A",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"A8",X"00",X"00",X"00",X"00",X"02",X"00",X"18",X"A8",X"00",
		X"00",X"00",X"00",X"00",X"00",X"08",X"A8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1A",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"A0",X"00",X"00",X"00",X"00",X"20",X"80",X"00",X"A0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"40",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"60",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"60",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"60",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"60",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"A8",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"28",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"2A",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"A8",X"00",X"00",X"00",X"00",X"55",X"55",X"54",X"A8",X"00",X"00",X"00",X"00",
		X"55",X"55",X"56",X"AA",X"00",X"00",X"00",X"00",X"55",X"55",X"58",X"AA",X"80",X"00",X"00",X"00",
		X"55",X"55",X"5A",X"AA",X"A0",X"00",X"00",X"00",X"55",X"55",X"5A",X"AA",X"80",X"00",X"00",X"00",
		X"55",X"55",X"5A",X"AA",X"A8",X"00",X"00",X"00",X"55",X"55",X"6A",X"AA",X"AA",X"80",X"00",X"00",
		X"55",X"55",X"55",X"55",X"5A",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"5A",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"5A",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"6A",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"68",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"68",X"80",X"00",X"00",
		X"55",X"55",X"55",X"55",X"42",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"4A",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"2A",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"A8",X"00",X"00",X"00",
		X"55",X"55",X"55",X"56",X"20",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"80",X"00",X"00",X"00",
		X"55",X"55",X"55",X"56",X"80",X"00",X"00",X"00",X"55",X"55",X"55",X"50",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"50",X"00",X"00",X"00",X"00",X"55",X"55",X"58",X"00",X"00",X"00",X"00",X"00",
		X"55",X"68",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"60",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"68",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"56",X"28",X"00",X"00",X"00",X"00",X"00",X"00",
		X"54",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"56",X"A2",X"00",X"00",X"00",X"00",X"00",X"00",
		X"58",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"5A",X"A8",X"00",X"00",X"00",X"00",X"00",X"00",
		X"5A",X"28",X"00",X"00",X"00",X"00",X"00",X"00",X"5A",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"A8",X"00",X"28",X"01",X"AA",X"AA",X"00",X"02",X"6A",X"00",X"08",X"01",X"95",X"56",
		X"00",X"00",X"9A",X"80",X"00",X"01",X"AA",X"A6",X"00",X"00",X"26",X"A8",X"00",X"01",X"AA",X"A6",
		X"00",X"00",X"09",X"A8",X"00",X"01",X"AA",X"A6",X"00",X"00",X"02",X"68",X"00",X"01",X"AA",X"A6",
		X"00",X"00",X"02",X"60",X"00",X"01",X"AA",X"A9",X"00",X"00",X"02",X"64",X"44",X"44",X"6A",X"A9",
		X"00",X"00",X"02",X"65",X"55",X"55",X"6A",X"A9",X"00",X"00",X"02",X"65",X"56",X"95",X"6A",X"A9",
		X"00",X"00",X"09",X"95",X"5A",X"95",X"6A",X"A9",X"00",X"00",X"09",X"95",X"55",X"95",X"6A",X"A9",
		X"00",X"00",X"09",X"95",X"59",X"95",X"6A",X"A9",X"00",X"00",X"09",X"95",X"59",X"95",X"55",X"55",
		X"00",X"00",X"09",X"95",X"69",X"A5",X"55",X"55",X"00",X"00",X"09",X"95",X"6A",X"65",X"55",X"55",
		X"A4",X"09",X"0A",X"A4",X"0A",X"02",X"98",X"00",X"A4",X"09",X"2A",X"94",X"00",X"02",X"98",X"00",
		X"A4",X"09",X"AA",X"50",X"00",X"02",X"98",X"00",X"54",X"09",X"AA",X"40",X"00",X"02",X"98",X"00",
		X"00",X"09",X"A9",X"40",X"00",X"02",X"60",X"00",X"00",X"09",X"A9",X"00",X"00",X"02",X"60",X"00",
		X"00",X"26",X"A5",X"00",X"00",X"0A",X"60",X"00",X"44",X"66",X"A4",X"44",X"A1",X"1A",X"60",X"00",
		X"55",X"66",X"95",X"56",X"A5",X"5A",X"60",X"00",X"A5",X"66",X"95",X"5A",X"95",X"5A",X"60",X"00",
		X"55",X"66",X"55",X"6A",X"55",X"5A",X"60",X"00",X"95",X"66",X"55",X"A9",X"95",X"5A",X"60",X"00",
		X"95",X"65",X"56",X"A6",X"95",X"5A",X"60",X"00",X"95",X"65",X"5A",X"9A",X"55",X"59",X"A0",X"00",
		X"55",X"65",X"6A",X"6A",X"55",X"69",X"80",X"00",X"55",X"A5",X"69",X"82",X"55",X"69",X"80",X"00",
		X"00",X"20",X"01",X"01",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"20",X"00",X"00",X"00",
		X"00",X"00",X"01",X"01",X"20",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"28",X"00",X"00",X"00",
		X"00",X"00",X"00",X"04",X"A8",X"02",X"00",X"00",X"00",X"00",X"00",X"02",X"A8",X"80",X"00",X"00",
		X"00",X"00",X"04",X"00",X"A8",X"08",X"20",X"00",X"00",X"00",X"10",X"28",X"0A",X"00",X"00",X"00",
		X"00",X"01",X"10",X"28",X"82",X"08",X"00",X"00",X"00",X"00",X"40",X"28",X"AA",X"80",X"00",X"00",
		X"00",X"00",X"02",X"0A",X"AA",X"20",X"00",X"00",X"00",X"00",X"28",X"02",X"A8",X"A0",X"00",X"00",
		X"00",X"00",X"8A",X"02",X"A2",X"00",X"00",X"00",X"00",X"21",X"00",X"00",X"A0",X"80",X"00",X"20",
		X"00",X"00",X"84",X"00",X"08",X"00",X"00",X"80",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"29",X"00",X"00",X"00",X"00",X"00",X"20",X"0A",X"A0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"28",X"00",X"00",X"00",X"00",X"00",X"00",X"28",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"A6",X"00",X"00",X"00",X"00",X"00",X"29",X"5A",X"55",
		X"00",X"00",X"00",X"00",X"2A",X"A9",X"55",X"55",X"00",X"00",X"00",X"00",X"55",X"55",X"95",X"59",
		X"55",X"55",X"6A",X"00",X"00",X"00",X"00",X"00",X"00",X"59",X"56",X"55",X"48",X"80",X"08",X"00",
		X"0A",X"55",X"95",X"56",X"55",X"52",X"00",X"00",X"00",X"A0",X"00",X"05",X"55",X"55",X"68",X"00",
		X"00",X"00",X"00",X"29",X"55",X"55",X"55",X"55",X"00",X"02",X"02",X"85",X"65",X"55",X"55",X"40",
		X"00",X"00",X"2A",X"55",X"55",X"95",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"80",
		X"00",X"05",X"55",X"65",X"55",X"54",X"00",X"00",X"02",X"15",X"55",X"55",X"65",X"55",X"5A",X"80",
		X"0A",X"55",X"55",X"95",X"55",X"55",X"55",X"50",X"95",X"55",X"59",X"56",X"55",X"55",X"40",X"00",
		X"95",X"65",X"55",X"95",X"55",X"55",X"80",X"00",X"55",X"55",X"95",X"56",X"00",X"00",X"00",X"00",
		X"65",X"55",X"55",X"58",X"02",X"00",X"00",X"00",X"55",X"54",X"00",X"00",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"08",X"00",X"02",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"40",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"60",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"40",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"8A",X"80",X"00",X"00",X"00",X"00",
		X"55",X"55",X"2A",X"80",X"00",X"00",X"00",X"00",X"55",X"55",X"AA",X"80",X"00",X"00",X"00",X"00",
		X"55",X"55",X"2A",X"A0",X"00",X"00",X"00",X"00",X"55",X"56",X"AA",X"A8",X"00",X"00",X"00",X"00",
		X"55",X"54",X"AA",X"A8",X"00",X"00",X"00",X"00",X"55",X"56",X"AA",X"A0",X"00",X"00",X"00",X"00",
		X"55",X"56",X"AA",X"00",X"00",X"00",X"00",X"00",X"55",X"56",X"A8",X"80",X"00",X"00",X"00",X"00",
		X"55",X"56",X"A2",X"00",X"00",X"00",X"00",X"00",X"55",X"5A",X"8A",X"00",X"00",X"00",X"00",X"00",
		X"55",X"5A",X"AA",X"00",X"00",X"00",X"00",X"00",X"55",X"5A",X"A2",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"A5",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"2A",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"02",X"85",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"02",X"95",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"09",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"01",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"15",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"A9",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"02",X"95",X"55",X"00",X"00",X"08",X"00",X"00",X"00",X"01",X"55",
		X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"95",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A5",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"05",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"01",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"01",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"08",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"21",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"2A",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"2A",X"55",
		X"00",X"00",X"00",X"00",X"00",X"02",X"AA",X"55",X"00",X"00",X"00",X"00",X"00",X"0A",X"AA",X"55",
		X"00",X"00",X"00",X"00",X"00",X"0A",X"AA",X"55",X"00",X"00",X"00",X"00",X"00",X"2A",X"AA",X"55",
		X"2A",X"95",X"A6",X"02",X"55",X"69",X"80",X"00",X"2A",X"96",X"A6",X"02",X"55",X"69",X"80",X"00",
		X"5A",X"5A",X"98",X"09",X"55",X"69",X"80",X"00",X"05",X"5A",X"60",X"09",X"55",X"69",X"80",X"00",
		X"02",X"5A",X"60",X"09",X"55",X"69",X"80",X"00",X"02",X"69",X"80",X"09",X"55",X"69",X"80",X"00",
		X"0A",X"69",X"80",X"26",X"55",X"69",X"80",X"00",X"0A",X"59",X"80",X"26",X"95",X"69",X"80",X"00",
		X"09",X"56",X"00",X"09",X"6A",X"59",X"80",X"00",X"09",X"58",X"00",X"0A",X"5A",X"A9",X"80",X"00",
		X"09",X"58",X"00",X"02",X"A5",X"A9",X"80",X"00",X"09",X"60",X"00",X"00",X"2A",X"55",X"60",X"00",
		X"0A",X"60",X"00",X"00",X"02",X"A9",X"60",X"00",X"02",X"A0",X"00",X"00",X"00",X"0A",X"A0",X"00",
		X"02",X"80",X"00",X"00",X"00",X"00",X"A8",X"00",X"02",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"80",X"00",
		X"00",X"00",X"00",X"00",X"28",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"20",X"00",X"55",X"55",X"95",X"00",X"00",X"00",X"00",X"00",X"11",X"59",X"55",
		X"00",X"00",X"08",X"00",X"8A",X"89",X"55",X"65",X"00",X"00",X"00",X"00",X"AA",X"95",X"65",X"11",
		X"00",X"00",X"00",X"25",X"55",X"55",X"55",X"50",X"00",X"00",X"2A",X"85",X"55",X"55",X"55",X"22",
		X"00",X"08",X"02",X"95",X"55",X"56",X"51",X"0A",X"00",X"00",X"09",X"55",X"55",X"55",X"55",X"45",
		X"08",X"20",X"20",X"55",X"56",X"59",X"55",X"55",X"00",X"00",X"15",X"55",X"55",X"55",X"55",X"55",
		X"00",X"89",X"55",X"55",X"55",X"55",X"55",X"55",X"22",X"95",X"55",X"59",X"59",X"55",X"55",X"55",
		X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"01",X"55",X"55",X"56",X"55",X"55",X"55",X"55",
		X"02",X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"2A",X"95",X"59",X"55",X"55",X"55",X"55",X"65",
		X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"56",X"A0",X"00",X"00",X"00",X"00",X"02",X"00",
		X"55",X"5A",X"00",X"00",X"00",X"00",X"00",X"00",X"65",X"55",X"54",X"40",X"80",X"00",X"00",X"00",
		X"65",X"65",X"55",X"56",X"28",X"00",X"00",X"00",X"59",X"95",X"55",X"55",X"55",X"56",X"80",X"00",
		X"66",X"55",X"55",X"55",X"55",X"55",X"50",X"00",X"55",X"65",X"95",X"55",X"55",X"55",X"54",X"80",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"55",X"55",X"65",X"65",X"55",X"55",X"55",X"10",
		X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"50",X"55",X"59",X"55",X"55",X"65",X"55",X"55",X"54",
		X"55",X"55",X"95",X"55",X"55",X"55",X"54",X"54",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"50",
		X"55",X"59",X"95",X"65",X"59",X"55",X"55",X"55",X"55",X"55",X"65",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"2A",X"08",
		X"02",X"00",X"00",X"00",X"00",X"80",X"95",X"55",X"08",X"00",X"00",X"02",X"A8",X"95",X"55",X"55",
		X"00",X"00",X"00",X"01",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"05",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"29",X"55",X"55",X"55",X"55",X"55",
		X"02",X"AA",X"55",X"55",X"55",X"55",X"55",X"55",X"02",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"05",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"29",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"54",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"5A",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"5A",X"02",
		X"55",X"55",X"55",X"55",X"55",X"55",X"48",X"08",X"55",X"55",X"55",X"55",X"54",X"00",X"20",X"0A",
		X"55",X"55",X"55",X"55",X"00",X"00",X"28",X"00",X"55",X"55",X"55",X"54",X"00",X"02",X"00",X"08",
		X"55",X"55",X"55",X"54",X"88",X"00",X"00",X"00",X"55",X"55",X"55",X"52",X"80",X"00",X"00",X"00",
		X"55",X"55",X"55",X"40",X"00",X"00",X"00",X"00",X"55",X"55",X"54",X"00",X"00",X"00",X"00",X"28",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"0A",X"95",X"55",X"55",X"55",X"55",X"55",X"00",X"02",X"95",X"55",X"55",X"55",X"55",X"55",
		X"00",X"0A",X"A5",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"02",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"A5",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"2A",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"25",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"29",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"15",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"05",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"01",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"09",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"09",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"04",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"95",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"25",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"25",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"09",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"0A",X"95",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A5",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",
		X"00",X"00",X"26",X"55",X"AA",X"65",X"55",X"55",X"00",X"00",X"26",X"55",X"82",X"65",X"55",X"55",
		X"00",X"00",X"26",X"55",X"82",X"69",X"59",X"6A",X"00",X"00",X"26",X"56",X"00",X"99",X"6A",X"AA",
		X"00",X"00",X"26",X"56",X"00",X"9A",X"AA",X"95",X"00",X"00",X"26",X"56",X"00",X"9A",X"A5",X"6A",
		X"00",X"00",X"26",X"56",X"00",X"9A",X"5A",X"80",X"00",X"00",X"26",X"58",X"02",X"55",X"A0",X"00",
		X"00",X"00",X"26",X"58",X"02",X"6A",X"00",X"00",X"00",X"00",X"25",X"58",X"02",X"A0",X"00",X"00",
		X"00",X"00",X"25",X"58",X"00",X"00",X"00",X"00",X"00",X"00",X"29",X"68",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"60",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"2A",X"00",X"00",X"00",X"00",X"00",X"02",X"8A",X"A5",
		X"00",X"00",X"00",X"00",X"01",X"01",X"5A",X"95",X"00",X"00",X"00",X"00",X"00",X"89",X"55",X"55",
		X"00",X"00",X"00",X"28",X"80",X"01",X"55",X"55",X"00",X"00",X"00",X"02",X"00",X"15",X"55",X"55",
		X"00",X"00",X"20",X"00",X"15",X"55",X"56",X"55",X"00",X"02",X"A0",X"09",X"55",X"55",X"55",X"55",
		X"00",X"00",X"80",X"29",X"55",X"55",X"95",X"55",X"0A",X"00",X"00",X"65",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"15",X"55",X"55",X"55",X"00",X"02",X"00",X"00",X"85",X"55",X"55",X"55",
		X"02",X"00",X"00",X"00",X"00",X"15",X"55",X"55",X"00",X"00",X"00",X"00",X"2A",X"95",X"55",X"56",
		X"00",X"00",X"02",X"02",X"00",X"14",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"80",X"01",X"55",
		X"69",X"55",X"55",X"59",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"65",X"55",
		X"55",X"65",X"96",X"55",X"55",X"55",X"55",X"55",X"59",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"55",X"55",
		X"65",X"65",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"59",X"55",X"95",X"55",X"55",X"55",X"55",X"59",X"55",X"56",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"95",X"59",
		X"55",X"56",X"55",X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"A5",X"59",X"55",
		X"56",X"55",X"55",X"95",X"55",X"59",X"55",X"55",X"55",X"55",X"55",X"65",X"55",X"55",X"55",X"55",
		X"55",X"55",X"65",X"55",X"55",X"55",X"55",X"54",X"55",X"51",X"95",X"56",X"55",X"55",X"55",X"56",
		X"55",X"85",X"56",X"55",X"55",X"55",X"55",X"50",X"59",X"12",X"65",X"55",X"55",X"55",X"50",X"00",
		X"55",X"02",X"55",X"55",X"55",X"55",X"55",X"00",X"60",X"00",X"AA",X"55",X"55",X"55",X"56",X"00",
		X"95",X"08",X"99",X"A5",X"55",X"55",X"00",X"00",X"64",X"A0",X"99",X"95",X"54",X"00",X"00",X"00",
		X"54",X"12",X"15",X"55",X"55",X"28",X"00",X"00",X"55",X"55",X"55",X"54",X"05",X"56",X"00",X"00",
		X"55",X"55",X"55",X"40",X"00",X"00",X"00",X"80",X"55",X"54",X"00",X"00",X"00",X"00",X"00",X"00",
		X"54",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"56",X"80",X"00",X"02",X"00",X"00",X"00",X"00",
		X"45",X"00",X"02",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"54",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"54",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"40",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"50",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"00",X"22",X"00",X"00",X"00",X"00",X"55",X"55",X"6A",X"20",X"00",X"00",X"00",X"00",
		X"55",X"54",X"AA",X"00",X"00",X"00",X"00",X"00",X"55",X"56",X"AA",X"00",X"00",X"00",X"00",X"00",
		X"55",X"54",X"A8",X"00",X"00",X"00",X"00",X"00",X"55",X"59",X"A0",X"00",X"00",X"00",X"00",X"00",
		X"55",X"61",X"A0",X"00",X"00",X"00",X"00",X"00",X"55",X"4A",X"80",X"00",X"00",X"00",X"00",X"00",
		X"55",X"8A",X"20",X"00",X"00",X"00",X"00",X"00",X"55",X"2A",X"A0",X"00",X"00",X"00",X"00",X"00",
		X"55",X"2A",X"28",X"00",X"00",X"00",X"00",X"00",X"55",X"A8",X"A8",X"20",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"50",X"A0",X"00",X"00",X"00",X"55",X"55",X"55",X"50",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"40",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"20",X"00",X"00",X"00",X"00",
		X"55",X"55",X"54",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"50",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"40",X"08",X"00",X"00",X"00",X"00",X"55",X"55",X"6A",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"68",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"48",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"28",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"68",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"48",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"A8",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"A0",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"A0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"01",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"02",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"02",X"95",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"15",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"29",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"02",X"95",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"95",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"85",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"A5",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"29",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"95",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"95",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",
		X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"80",X"00",X"00",X"00",
		X"00",X"02",X"8A",X"80",X"0A",X"A0",X"08",X"08",X"00",X"00",X"22",X"25",X"50",X"2A",X"A0",X"02",
		X"00",X"00",X"25",X"55",X"55",X"5A",X"AA",X"89",X"00",X"00",X"02",X"55",X"55",X"55",X"56",X"25",
		X"00",X"00",X"02",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"95",X"55",X"55",X"55",X"55",
		X"00",X"00",X"09",X"55",X"55",X"55",X"55",X"A0",X"00",X"00",X"00",X"AA",X"25",X"54",X"00",X"00",
		X"00",X"00",X"02",X"00",X"08",X"80",X"80",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"28",X"55",X"00",X"00",X"08",X"82",X"AA",X"AA",X"95",X"55",
		X"00",X"02",X"A9",X"55",X"55",X"55",X"55",X"54",X"01",X"55",X"55",X"55",X"55",X"55",X"54",X"00",
		X"00",X"15",X"55",X"55",X"55",X"54",X"00",X"00",X"00",X"05",X"55",X"55",X"55",X"56",X"20",X"00",
		X"80",X"80",X"95",X"55",X"55",X"55",X"00",X"20",X"AA",X"AA",X"15",X"55",X"55",X"54",X"00",X"80",
		X"6A",X"55",X"55",X"55",X"51",X"00",X"00",X"00",X"55",X"55",X"55",X"50",X"00",X"00",X"00",X"00",
		X"55",X"55",X"9A",X"A8",X"00",X"00",X"00",X"00",X"55",X"58",X"00",X"10",X"00",X"00",X"00",X"00",
		X"54",X"2A",X"80",X"00",X"00",X"00",X"00",X"00",X"95",X"55",X"68",X"80",X"10",X"00",X"00",X"00",
		X"80",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"54",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"54",X"00",X"00",X"00",X"00",X"09",X"55",X"00",X"00",X"00",X"00",
		X"00",X"08",X"08",X"80",X"08",X"80",X"80",X"00",X"00",X"00",X"22",X"00",X"00",X"02",X"00",X"00",
		X"00",X"08",X"80",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"2A",X"AA",X"AA",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"A8",X"00",
		X"00",X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"02",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",
		X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"00",X"0A",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",
		X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"0A",X"AA",X"AA",X"AA",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"2A",X"AA",X"AA",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"A8",X"00",
		X"00",X"2A",X"AB",X"EA",X"BE",X"AF",X"FA",X"A0",X"02",X"AA",X"AE",X"BA",X"EB",X"AA",X"EA",X"A8",
		X"00",X"AA",X"AE",X"BA",X"EB",X"AB",X"AA",X"AA",X"00",X"AA",X"AE",X"BA",X"EB",X"AF",X"AA",X"AA",
		X"00",X"2A",X"AE",X"BA",X"EB",X"AC",X"BA",X"A8",X"00",X"0A",X"AB",X"EA",X"BE",X"AB",X"EA",X"A0",
		X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"0A",X"AA",X"AA",X"AA",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"2A",X"AA",X"AA",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"A8",X"00",
		X"00",X"2A",X"AB",X"EA",X"BE",X"AB",X"FA",X"A0",X"02",X"AA",X"AE",X"BA",X"EB",X"AE",X"AA",X"A8",
		X"00",X"AA",X"AE",X"BA",X"EB",X"AE",X"AA",X"AA",X"00",X"AA",X"AE",X"BA",X"EB",X"AB",X"EA",X"AA",
		X"00",X"2A",X"AE",X"BA",X"EB",X"AE",X"AA",X"A8",X"00",X"0A",X"AB",X"EA",X"BE",X"AF",X"FA",X"A0",
		X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"0A",X"AA",X"AA",X"AA",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"2A",X"AA",X"AA",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"A8",X"00",
		X"00",X"2A",X"AB",X"EA",X"BE",X"AE",X"AA",X"A0",X"02",X"AA",X"AE",X"BA",X"EB",X"AE",X"AA",X"A8",
		X"00",X"AA",X"AE",X"BA",X"EB",X"AF",X"FA",X"AA",X"00",X"AA",X"AE",X"BA",X"EB",X"AE",X"EA",X"AA",
		X"00",X"2A",X"AE",X"BA",X"EB",X"AF",X"AA",X"A8",X"00",X"0A",X"AB",X"EA",X"BE",X"AE",X"AA",X"A0",
		X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"0A",X"AA",X"AA",X"AA",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"2A",X"AA",X"AA",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"A8",X"00",
		X"00",X"2A",X"AB",X"EA",X"BE",X"AB",X"EA",X"A0",X"02",X"AA",X"AE",X"BA",X"EB",X"AE",X"BA",X"A8",
		X"00",X"AA",X"AE",X"BA",X"EB",X"AE",X"BA",X"AA",X"00",X"AA",X"AE",X"BA",X"EB",X"AB",X"FA",X"AA",
		X"00",X"2A",X"AE",X"BA",X"EB",X"AA",X"BA",X"A8",X"00",X"0A",X"AB",X"EA",X"BE",X"AF",X"EA",X"A0",
		X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"0A",X"AA",X"AA",X"AA",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"2A",X"AA",X"AA",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"A8",X"00",
		X"00",X"2A",X"AB",X"EA",X"BE",X"AB",X"EA",X"A0",X"02",X"AA",X"AE",X"BA",X"EB",X"AE",X"BA",X"A8",
		X"00",X"AA",X"AE",X"BA",X"EB",X"AE",X"BA",X"AA",X"00",X"AA",X"AE",X"BA",X"EB",X"AB",X"EA",X"AA",
		X"00",X"2A",X"AE",X"BA",X"EB",X"AE",X"BA",X"A8",X"00",X"0A",X"AB",X"EA",X"BE",X"AB",X"EA",X"A0",
		X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"0A",X"AA",X"AA",X"AA",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"2A",X"AA",X"AA",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"A8",X"00",
		X"00",X"2A",X"BE",X"AB",X"EA",X"FF",X"AE",X"A0",X"02",X"AA",X"EB",X"AE",X"BA",X"AE",X"AE",X"A8",
		X"00",X"AA",X"EB",X"AE",X"BA",X"BA",X"AE",X"AA",X"00",X"AA",X"EB",X"AE",X"BA",X"FA",X"AF",X"AA",
		X"00",X"2A",X"EB",X"AE",X"BA",X"EB",X"AE",X"A8",X"00",X"0A",X"BE",X"AB",X"EA",X"BE",X"AE",X"A0",
		X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"0A",X"AA",X"AA",X"AA",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"2A",X"AA",X"AA",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"A8",X"00",
		X"00",X"2A",X"BE",X"AB",X"EA",X"BE",X"AE",X"A0",X"02",X"AA",X"EB",X"AE",X"BA",X"EB",X"AE",X"A8",
		X"00",X"AA",X"EB",X"AE",X"BA",X"EB",X"AE",X"AA",X"00",X"AA",X"EB",X"AE",X"BA",X"BF",X"AF",X"AA",
		X"00",X"2A",X"EB",X"AE",X"BA",X"AB",X"AE",X"A8",X"00",X"0A",X"BE",X"AB",X"EA",X"FE",X"AE",X"A0",
		X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"0A",X"AA",X"AA",X"AA",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
