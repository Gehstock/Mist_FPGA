library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity tropical_spr_bit6 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of tropical_spr_bit6 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"0F",X"1F",X"13",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"F0",X"F8",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"F0",X"E0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"0F",X"07",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"1F",X"1F",X"1F",X"1F",X"3C",X"3C",X"3C",X"78",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"F8",X"F0",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"1F",X"0F",X"07",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F8",X"F8",X"F8",X"F8",X"1C",X"0C",X"0C",X"0E",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"03",X"03",X"03",X"02",X"04",X"00",
		X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"F0",X"E0",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"F8",X"F0",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"1F",X"0F",X"07",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"07",X"07",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"C0",X"C0",X"C0",X"40",X"20",X"00",
		X"70",X"F8",X"FC",X"FC",X"FE",X"FE",X"7F",X"73",X"21",X"21",X"00",X"01",X"03",X"07",X"07",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"E0",X"E0",X"F0",X"30",
		X"0C",X"1E",X"1E",X"1E",X"1E",X"1F",X"1C",X"08",X"08",X"0C",X"04",X"06",X"03",X"03",X"03",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"1A",X"3C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",
		X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"80",X"80",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"02",X"00",X"00",
		X"52",X"38",X"0D",X"2A",X"1B",X"0B",X"03",X"0B",X"07",X"02",X"00",X"03",X"07",X"27",X"17",X"1F",
		X"00",X"44",X"01",X"24",X"42",X"E7",X"D3",X"87",X"ED",X"D1",X"87",X"E3",X"F8",X"F5",X"F7",X"BF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"02",X"08",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"20",X"00",X"04",X"00",X"80",X"20",X"01",X"28",X"80",
		X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"04",X"00",X"00",
		X"80",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"80",X"08",X"00",X"00",X"02",X"40",X"00",X"00",
		X"02",X"04",X"02",X"01",X"01",X"00",X"01",X"00",X"00",X"04",X"0F",X"1D",X"39",X"27",X"47",X"01",
		X"FC",X"7C",X"54",X"2C",X"F8",X"F8",X"F0",X"D0",X"10",X"33",X"CF",X"F9",X"FC",X"FF",X"F7",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"60",X"20",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"03",X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"06",
		X"C3",X"C2",X"C2",X"C2",X"C2",X"C2",X"40",X"C0",X"C0",X"60",X"70",X"70",X"30",X"30",X"60",X"60",
		X"00",X"03",X"07",X"0F",X"0F",X"0F",X"07",X"07",X"07",X"07",X"03",X"01",X"00",X"11",X"3F",X"3F",
		X"00",X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"C0",X"C0",X"C0",X"F8",X"FC",X"FE",
		X"00",X"00",X"00",X"10",X"01",X"01",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"58",X"18",X"00",X"80",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"03",X"01",X"01",X"00",X"00",X"01",X"03",X"00",X"00",X"01",X"01",X"01",X"01",X"04",X"04",
		X"E0",X"70",X"70",X"F0",X"F0",X"F0",X"F0",X"B0",X"90",X"90",X"90",X"B0",X"B0",X"F0",X"E0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",
		X"01",X"03",X"07",X"07",X"03",X"03",X"07",X"05",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"E4",X"F8",X"E2",X"FC",X"F8",X"E4",X"B8",X"48",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"07",X"0B",X"0B",X"17",X"07",X"07",X"05",X"04",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"C0",X"E0",X"F0",X"E8",X"F6",X"F8",X"C0",X"A0",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"03",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"05",X"07",X"07",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"C0",X"C0",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"06",X"05",X"07",X"07",X"07",X"07",X"07",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"03",X"05",X"0B",X"0B",X"0F",X"0F",X"0F",X"0F",X"07",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"C0",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"03",X"06",X"05",X"0D",X"0F",X"0F",X"0F",X"07",X"07",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",X"E0",X"E0",X"C0",X"00",
		X"00",X"00",X"00",X"03",X"06",X"0D",X"0B",X"1B",X"1F",X"1F",X"1F",X"0F",X"0F",X"07",X"03",X"00",
		X"00",X"00",X"00",X"C0",X"E0",X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",X"F0",X"F0",X"E0",X"C0",X"00",
		X"0F",X"09",X"1B",X"17",X"37",X"3F",X"3F",X"3F",X"3F",X"1F",X"1F",X"0F",X"0F",X"03",X"00",X"00",
		X"F0",X"F0",X"F8",X"F8",X"FC",X"FC",X"FC",X"FC",X"FC",X"F8",X"F8",X"F0",X"F0",X"C0",X"00",X"00",
		X"37",X"3F",X"77",X"67",X"67",X"6F",X"7F",X"7F",X"3F",X"3F",X"1F",X"1F",X"0F",X"03",X"00",X"00",
		X"FC",X"FC",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FC",X"FC",X"F8",X"F8",X"F0",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"04",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"20",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"0C",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"30",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"04",X"00",X"1C",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"20",X"00",X"38",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0E",X"18",X"00",X"38",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"30",X"08",X"00",X"1C",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"1C",X"30",X"00",X"68",X"F0",X"F3",X"7E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"78",X"38",X"0C",X"00",X"0E",X"0E",X"0F",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"78",X"C0",X"80",X"00",X"80",X"C0",X"8C",X"9B",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"7E",X"1E",X"03",X"01",X"00",X"03",X"03",X"01",X"CF",X"7C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"03",X"02",X"03",X"03",X"0F",X"07",X"03",
		X"00",X"00",X"FF",X"FE",X"F8",X"F0",X"C0",X"80",X"00",X"80",X"80",X"00",X"C0",X"80",X"F1",X"EF",
		X"00",X"00",X"7F",X"3F",X"0F",X"07",X"01",X"00",X"00",X"00",X"03",X"01",X"03",X"61",X"DF",X"F3",
		X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"00",X"C0",X"C0",X"C0",X"C0",X"F0",X"F0",X"C0",
		X"01",X"03",X"03",X"03",X"03",X"07",X"06",X"04",X"00",X"0C",X"0E",X"0F",X"0E",X"3E",X"3C",X"1F",
		X"FC",X"F8",X"F0",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"78",X"DF",
		X"1F",X"0F",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"F9",
		X"80",X"C0",X"C0",X"C0",X"40",X"60",X"60",X"20",X"00",X"70",X"70",X"F0",X"70",X"7C",X"BC",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",
		X"0F",X"1E",X"1E",X"1C",X"38",X"30",X"20",X"00",X"64",X"70",X"7C",X"FC",X"FC",X"F9",X"FF",X"1F",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"F3",X"3F",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"F3",X"01",
		X"F0",X"18",X"08",X"08",X"0C",X"0C",X"04",X"00",X"1E",X"1E",X"3E",X"3F",X"3F",X"1F",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"03",X"03",X"07",X"0F",X"0F",X"03",X"00",
		X"40",X"00",X"E8",X"C8",X"C8",X"E0",X"FC",X"FC",X"F8",X"F8",X"F8",X"F0",X"F3",X"FF",X"FF",X"3E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C1",X"FF",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"FF",X"71",X"82",
		X"02",X"00",X"1F",X"1F",X"0F",X"0F",X"3F",X"3F",X"1F",X"1F",X"1F",X"0F",X"8F",X"FF",X"FF",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"C0",X"E0",X"F0",X"E0",X"C0",X"A0",X"00",
		X"07",X"0E",X"0E",X"0E",X"0F",X"1F",X"1F",X"1F",X"3F",X"7F",X"FF",X"FF",X"FF",X"3F",X"0F",X"01",
		X"40",X"40",X"40",X"40",X"00",X"F0",X"F0",X"E0",X"E0",X"E0",X"E0",X"C0",X"F0",X"FC",X"FF",X"F3",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"1F",X"FB",X"E7",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"8F",X"FB",X"0C",
		X"07",X"1F",X"1F",X"0F",X"0F",X"0F",X"0F",X"07",X"07",X"07",X"07",X"03",X"0F",X"FF",X"F8",X"E0",
		X"E0",X"F0",X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",X"FC",X"FE",X"FF",X"FF",X"FF",X"FC",X"F0",X"08",
		X"02",X"02",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"18",X"08",X"0C",X"04",X"0E",X"1E",X"3F",X"7F",X"3F",X"3F",X"1F",X"1F",X"0F",X"0F",X"07",X"07",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"80",X"80",X"80",X"44",X"7C",X"3E",X"3E",X"3E",X"1F",X"1F",X"0F",X"0F",X"0F",X"07",X"07",
		X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"40",X"1A",X"30",X"85",X"11",X"45",X"18",X"27",X"FF",
		X"00",X"00",X"00",X"18",X"38",X"50",X"98",X"38",X"14",X"88",X"D5",X"94",X"42",X"E8",X"C6",X"B4",
		X"00",X"00",X"02",X"00",X"01",X"10",X"06",X"0C",X"31",X"07",X"34",X"8F",X"AA",X"45",X"BA",X"75",
		X"18",X"38",X"70",X"58",X"B8",X"EC",X"D8",X"15",X"EC",X"B6",X"62",X"8E",X"ED",X"D4",X"49",X"AB",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0E",X"1F",X"35",X"8A",X"3D",X"02",X"EE",
		X"00",X"00",X"00",X"06",X"0C",X"0B",X"1C",X"1E",X"15",X"0A",X"0B",X"02",X"85",X"23",X"09",X"84",
		X"00",X"00",X"00",X"81",X"44",X"08",X"C0",X"12",X"88",X"6E",X"48",X"F5",X"74",X"93",X"1F",X"B6",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"04",X"B0",X"90",X"19",X"A0",X"F0",X"DB",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"0C",X"1E",X"17",X"3D",X"0B",X"59",X"F5",X"06",X"EC",X"B5",
		X"0E",X"1D",X"17",X"1A",X"0F",X"0D",X"1A",X"0D",X"09",X"12",X"05",X"87",X"41",X"00",X"C2",X"61",
		X"90",X"20",X"D8",X"40",X"B8",X"DC",X"F8",X"6D",X"E7",X"D3",X"EE",X"AF",X"D0",X"94",X"C3",X"79",
		X"00",X"00",X"00",X"00",X"00",X"80",X"20",X"10",X"80",X"20",X"32",X"04",X"64",X"02",X"1D",X"8F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"07",X"09",X"0C",X"86",X"25",X"29",X"5C",X"77",
		X"00",X"08",X"1E",X"0F",X"0A",X"04",X"06",X"09",X"0C",X"86",X"44",X"82",X"C5",X"21",X"48",X"59",
		X"00",X"00",X"00",X"34",X"A0",X"43",X"11",X"58",X"5A",X"43",X"6F",X"E9",X"6D",X"3D",X"F8",X"5A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"D0",X"0A",X"C1",X"C5",X"AA",X"FE",
		X"00",X"00",X"00",X"00",X"04",X"06",X"0B",X"0D",X"25",X"0B",X"17",X"1D",X"6A",X"13",X"15",X"EB",
		X"17",X"1D",X"0E",X"0D",X"16",X"19",X"0C",X"8A",X"44",X"95",X"42",X"11",X"B1",X"D0",X"88",X"A0",
		X"80",X"1A",X"A8",X"D1",X"5C",X"1C",X"CE",X"BF",X"B5",X"F6",X"BD",X"46",X"1E",X"5D",X"0B",X"06",
		X"00",X"00",X"00",X"00",X"80",X"80",X"20",X"40",X"D0",X"E0",X"24",X"F8",X"C4",X"B0",X"76",X"94",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"04",X"00",X"01",X"00",X"00",
		X"00",X"00",X"20",X"00",X"80",X"20",X"50",X"38",X"78",X"BC",X"12",X"34",X"18",X"20",X"00",X"00",
		X"00",X"02",X"01",X"04",X"23",X"01",X"04",X"01",X"0B",X"01",X"40",X"05",X"00",X"00",X"00",X"09",
		X"80",X"40",X"C0",X"E0",X"E0",X"70",X"B0",X"F0",X"D8",X"44",X"91",X"C7",X"F2",X"5D",X"36",X"C1",
		X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"04",X"00",X"01",X"00",X"00",X"04",X"00",
		X"00",X"00",X"00",X"50",X"00",X"50",X"88",X"68",X"30",X"78",X"F4",X"62",X"30",X"00",X"40",X"00",
		X"01",X"14",X"03",X"01",X"03",X"05",X"01",X"2B",X"01",X"04",X"01",X"00",X"00",X"04",X"40",X"00",
		X"C0",X"C0",X"C0",X"E0",X"A0",X"E0",X"E0",X"70",X"F2",X"F9",X"AF",X"72",X"E5",X"70",X"DC",X"16",
		X"80",X"00",X"00",X"00",X"02",X"00",X"20",X"00",X"00",X"09",X"06",X"C3",X"FF",X"BF",X"EF",X"6D",
		X"00",X"10",X"04",X"28",X"18",X"12",X"3C",X"1E",X"1A",X"3F",X"EE",X"F6",X"F0",X"F8",X"E5",X"93",
		X"07",X"8E",X"0C",X"4E",X"26",X"BE",X"1F",X"0F",X"0F",X"5F",X"1F",X"3B",X"9F",X"3D",X"5F",X"F3",
		X"1B",X"B1",X"73",X"6F",X"C1",X"20",X"C9",X"92",X"E1",X"A5",X"9B",X"4F",X"9F",X"AB",X"DD",X"99",
		X"11",X"11",X"12",X"00",X"48",X"30",X"25",X"38",X"7D",X"71",X"A4",X"89",X"D8",X"92",X"A4",X"00",
		X"00",X"A1",X"C8",X"42",X"86",X"34",X"60",X"20",X"92",X"20",X"09",X"40",X"A0",X"B2",X"00",X"00",
		X"00",X"20",X"00",X"00",X"08",X"00",X"00",X"82",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"40",
		X"10",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"40",X"00",X"00",
		X"01",X"10",X"30",X"00",X"00",X"00",X"01",X"01",X"01",X"04",X"0C",X"00",X"01",X"07",X"07",X"07",
		X"C6",X"C0",X"00",X"18",X"F4",X"FE",X"DA",X"FB",X"F9",X"F1",X"07",X"7D",X"79",X"39",X"B1",X"83",
		X"00",X"90",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"06",X"07",X"07",X"07",X"07",X"07",X"07",X"07",
		X"60",X"60",X"60",X"60",X"20",X"20",X"20",X"20",X"60",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"3F",X"1F",X"0F",X"17",X"17",X"13",X"20",X"61",X"00",X"00",X"08",X"0C",X"0F",X"07",X"07",X"03",
		X"FE",X"7E",X"7B",X"79",X"78",X"78",X"04",X"36",X"B0",X"B8",X"98",X"18",X"3C",X"BC",X"9C",X"DC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"06",X"06",X"06",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",
		X"A0",X"A0",X"A0",X"A0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"DF",X"FC",X"FF",X"79",X"7E",X"19",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"80",X"60",X"80",X"60",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FD",X"FF",X"FF",X"7E",X"0D",X"06",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"90",X"60",X"90",X"60",X"80",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"02",X"05",X"0D",X"0F",X"0F",X"07",X"03",X"07",X"07",
		X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"A0",X"A0",X"40",X"40",X"E0",X"E0",X"C0",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"05",X"02",X"0A",X"05",X"07",X"03",X"07",X"07",X"0F",X"0F",X"07",X"07",
		X"00",X"00",X"00",X"00",X"00",X"80",X"A0",X"40",X"50",X"A0",X"E0",X"C0",X"80",X"80",X"80",X"00",
		X"01",X"03",X"07",X"07",X"07",X"07",X"07",X"07",X"03",X"01",X"01",X"03",X"07",X"0F",X"0F",X"1F",
		X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",X"F8",X"F0",X"F0",X"F8",X"FC",X"FE",X"FF",X"FF",X"C7",X"E9",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"03",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"18",X"F8",X"D0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"80",X"E0",X"F0",X"F0",X"F8",X"38",X"7C",X"DC",X"8E",X"8E",X"C7",X"F3",X"79",X"FC",X"B8",X"1C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"40",
		X"0F",X"0F",X"1F",X"1F",X"1F",X"1F",X"1F",X"0F",X"0F",X"1F",X"3F",X"7F",X"FF",X"FF",X"E3",X"97",
		X"80",X"C0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"C0",X"80",X"80",X"C0",X"E0",X"F0",X"F0",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"18",X"1F",X"0B",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"C0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"02",
		X"01",X"07",X"0F",X"0F",X"1F",X"1F",X"3F",X"26",X"68",X"4A",X"DB",X"B0",X"B0",X"60",X"40",X"C8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"07",X"07",X"07",X"07",X"07",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"01",X"03",X"03",X"03",X"03",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"7C",X"00",X"07",X"03",X"07",X"07",X"03",X"01",
		X"80",X"80",X"C0",X"E0",X"F0",X"F0",X"38",X"08",X"18",X"64",X"04",X"80",X"C0",X"C0",X"E0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"15",X"1E",X"1A",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"1F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"1F",
		X"FF",X"FF",X"FE",X"FE",X"F8",X"E0",X"E0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"03",X"03",X"07",X"07",X"0F",X"0F",X"1F",X"1F",X"1F",X"3E",X"3C",X"30",X"70",X"58",
		X"00",X"10",X"2C",X"78",X"78",X"70",X"18",X"1E",X"07",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E1",X"FF",X"7F",X"1E",X"00",X"00",X"00",X"00",
		X"3E",X"3F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"7F",X"3F",X"1F",X"0F",X"01",X"00",X"00",X"00",
		X"00",X"00",X"80",X"80",X"80",X"00",X"00",X"E0",X"F8",X"EC",X"F6",X"F7",X"FB",X"FB",X"7D",X"7F",
		X"00",X"00",X"00",X"28",X"14",X"1C",X"0E",X"0E",X"06",X"04",X"0C",X"5C",X"B8",X"D0",X"C0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"08",X"18",X"18",X"50",X"D0",X"D0",X"B0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"06",X"1F",X"37",X"6F",X"EF",X"DF",X"BF",X"BC",X"7E",
		X"7C",X"FC",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FE",X"FC",X"F0",X"F8",X"9C",X"7C",X"FC",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"14",X"28",X"38",X"70",X"70",X"60",X"20",X"30",X"3A",X"1D",X"09",X"01",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"06",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"81",X"C3",X"67",X"71",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"41",X"A8",X"7B",X"E7",X"1E",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CF",X"3F",X"FF",X"F7",X"83",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",
		X"F0",X"FE",X"F7",X"F9",X"FE",X"FF",X"EF",X"1F",X"1F",X"3F",X"3F",X"3F",X"7C",X"FC",X"FC",X"F8",
		X"00",X"00",X"80",X"C0",X"E0",X"70",X"F0",X"F8",X"F8",X"E8",X"E8",X"D0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"01",X"00",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"E0",X"60",X"50",X"58",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"38",X"FC",X"3F",X"E7",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",
		X"00",X"00",X"00",X"FF",X"FF",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"3E",X"FC",
		X"07",X"07",X"C3",X"C1",X"E1",X"10",X"08",X"04",X"00",X"02",X"03",X"1F",X"FF",X"FF",X"FF",X"3F",
		X"FC",X"FC",X"FE",X"F4",X"F0",X"F0",X"60",X"00",X"01",X"00",X"00",X"00",X"80",X"C0",X"E0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"60",X"60",X"C0",X"70",X"30",X"00",X"00",X"10",X"18",X"18",X"08",X"0C",X"0C",X"0C",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"E0",X"F8",X"7C",X"1F",X"03",X"03",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"0E",X"0C",X"00",X"00",X"01",X"03",X"F3",X"F8",X"7F",X"1F",X"1F",X"07",X"03",X"10",X"1C",
		X"13",X"31",X"71",X"61",X"ED",X"DD",X"FF",X"FF",X"3F",X"FE",X"FE",X"FF",X"FC",X"FE",X"FE",X"3E",
		X"E0",X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",X"E0",X"E0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"40",X"E0",X"E0",X"30",X"38",X"2C",X"06",X"03",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"D0",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"1C",X"0E",X"06",X"03",X"00",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"E0",X"70",X"38",X"3D",X"1E",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F8",X"FC",X"7C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"30",X"38",X"38",X"0C",X"1C",X"1A",X"02",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"01",X"01",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",
		X"6C",X"CC",X"CE",X"9E",X"DE",X"3E",X"9E",X"BE",X"BE",X"FE",X"FE",X"FC",X"BC",X"9C",X"9C",X"98",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"C7",X"0F",X"1F",X"BF",X"DF",X"FF",X"FE",X"FE",X"FC",X"FC",X"FA",X"F2",X"E3",X"C1",X"81",
		X"F8",X"38",X"F8",X"98",X"88",X"08",X"08",X"18",X"18",X"30",X"30",X"70",X"70",X"F0",X"F0",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"00",
		X"07",X"0F",X"1F",X"1F",X"1F",X"1F",X"3F",X"3F",X"47",X"3B",X"77",X"77",X"EF",X"FF",X"DF",X"DF",
		X"00",X"00",X"84",X"8C",X"0C",X"18",X"7E",X"FF",X"BF",X"BC",X"B8",X"7C",X"F8",X"78",X"78",X"70",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"E0",X"F8",X"3C",X"04",X"00",X"00",X"00",X"00",
		X"01",X"01",X"01",X"00",X"00",X"02",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"02",
		X"18",X"18",X"08",X"88",X"88",X"88",X"98",X"98",X"F8",X"F8",X"B0",X"B0",X"90",X"90",X"50",X"50",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"03",X"03",X"03",X"03",X"03",X"01",X"01",X"03",X"03",X"07",X"07",X"0F",X"0B",X"0B",
		X"00",X"00",X"00",X"C0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F8",X"FC",X"FF",X"F7",X"E1",X"C0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"60",X"30",
		X"00",X"00",X"00",X"00",X"01",X"03",X"00",X"00",X"03",X"03",X"03",X"03",X"03",X"00",X"00",X"00",
		X"60",X"00",X"00",X"00",X"00",X"00",X"50",X"50",X"78",X"58",X"58",X"58",X"58",X"78",X"78",X"38",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"0E",X"18",X"11",
		X"00",X"00",X"00",X"03",X"07",X"0F",X"0F",X"0F",X"0F",X"1F",X"7D",X"FD",X"9F",X"1B",X"1B",X"1B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"60",X"04",X"0E",X"FE",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"22",X"21",X"01",X"01",X"00",X"00",X"00",X"00",X"01",X"03",X"00",X"02",X"07",X"07",X"07",X"07",
		X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"00",X"00",X"60",X"60",X"60",X"60",X"60",X"40",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"FD",X"3F",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"02",X"01",X"18",X"23",X"03",X"4F",X"27",X"0F",X"1E",X"AF",X"1B",X"64",X"91",X"06",X"21",
		X"D6",X"FF",X"2D",X"34",X"0E",X"3E",X"9D",X"FF",X"EF",X"FF",X"FD",X"BF",X"F7",X"FF",X"BB",X"1D",
		X"00",X"02",X"80",X"80",X"40",X"40",X"89",X"E1",X"F0",X"F8",X"FE",X"FF",X"3F",X"AF",X"B7",X"D7",
		X"05",X"05",X"00",X"02",X"02",X"01",X"01",X"04",X"00",X"10",X"40",X"00",X"90",X"82",X"A8",X"80",
		X"84",X"86",X"84",X"02",X"00",X"01",X"03",X"06",X"06",X"00",X"16",X"84",X"05",X"27",X"C6",X"97",
		X"20",X"02",X"10",X"44",X"00",X"90",X"04",X"10",X"80",X"08",X"30",X"60",X"30",X"12",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"41",X"00",
		X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"08",X"80",X"00",X"00",X"12",X"0D",X"07",X"05",
		X"00",X"00",X"00",X"04",X"00",X"00",X"20",X"00",X"04",X"02",X"86",X"0B",X"03",X"11",X"0D",X"A4",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"02",X"11",X"05",X"53",X"61",X"69",X"3D",X"3B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"08",X"20",X"A0",X"80",X"80",X"C0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"13",X"20",X"04",X"0C",X"13",X"01",X"00",X"02",X"07",X"01",X"00",X"00",X"01",X"00",X"00",X"00",
		X"AE",X"58",X"21",X"9B",X"7F",X"FF",X"3E",X"1C",X"FC",X"EE",X"C7",X"83",X"03",X"04",X"01",X"18",
		X"44",X"36",X"9E",X"2F",X"BD",X"FC",X"9E",X"5F",X"BD",X"6E",X"B7",X"83",X"57",X"AD",X"CD",X"5E",
		X"F4",X"FD",X"7E",X"FE",X"7D",X"7F",X"3F",X"DD",X"BF",X"0F",X"A7",X"93",X"7B",X"FF",X"BE",X"1F",
		X"21",X"90",X"2B",X"73",X"91",X"0D",X"8C",X"A6",X"BB",X"FB",X"FD",X"FF",X"FF",X"FF",X"FF",X"EF",
		X"DE",X"CF",X"A7",X"93",X"D9",X"F3",X"FB",X"FB",X"FD",X"FF",X"FE",X"7F",X"BE",X"5F",X"8F",X"CE",
		X"F9",X"6C",X"6C",X"91",X"9D",X"D3",X"EE",X"F4",X"F2",X"F0",X"FD",X"FC",X"FE",X"FE",X"F5",X"F6",
		X"C0",X"20",X"80",X"00",X"C0",X"20",X"80",X"00",X"C8",X"40",X"22",X"40",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1B",X"3B",X"3B",X"2D",X"2D",X"60",X"40",X"41",X"81",X"00",X"04",X"0A",X"05",X"06",X"08",X"04",
		X"FC",X"EC",X"F4",X"F0",X"EE",X"FF",X"FF",X"FF",X"DF",X"DF",X"CF",X"4F",X"07",X"03",X"01",X"10",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"00",X"00",X"40",X"01",X"00",X"00",X"00",X"00",
		X"01",X"FF",X"FF",X"FF",X"FF",X"F8",X"C0",X"01",X"00",X"1F",X"6F",X"9F",X"3E",X"38",X"01",X"00",
		X"1E",X"07",X"01",X"04",X"03",X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"60",X"E0",X"F0",X"F0",X"38",X"B8",X"FC",X"FC",X"FE",X"FE",X"7F",X"7F",X"3F",X"3F",X"1F",X"1F",
		X"3F",X"37",X"2F",X"0F",X"77",X"FF",X"FF",X"FB",X"F9",X"FB",X"F3",X"E2",X"C0",X"80",X"04",X"0C",
		X"D8",X"DC",X"DC",X"B4",X"B4",X"06",X"02",X"82",X"81",X"00",X"20",X"50",X"A0",X"60",X"10",X"20",
		X"81",X"F7",X"CF",X"BF",X"7F",X"FF",X"FF",X"03",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",
		X"06",X"05",X"0C",X"08",X"18",X"19",X"3F",X"3F",X"7F",X"7F",X"FE",X"FE",X"FC",X"FC",X"F8",X"F8",
		X"90",X"30",X"60",X"60",X"C0",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"54",X"2C",X"40",X"04",X"04",X"06",X"05",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"03",X"0F",X"1F",X"3D",X"7D",X"DB",X"DF",X"9F",X"37",X"2F",X"2F",X"3F",X"7E",X"7F",X"FF",
		X"C0",X"E0",X"F0",X"F8",X"FC",X"FE",X"FE",X"CF",X"C7",X"C3",X"C1",X"80",X"80",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"70",X"60",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"78",X"3C",X"06",X"0F",X"1B",X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"18",X"9C",X"C8",X"C8",X"70",X"30",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"70",X"FF",X"FF",X"FE",X"F0",X"70",X"78",X"B8",X"DC",X"DC",X"EE",X"F7",X"FB",X"FF",X"FF",
		X"30",X"E0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"0E",X"06",X"07",X"03",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"08",X"0F",X"1F",X"3F",X"7F",X"7F",X"FF",X"FF",X"E1",X"83",X"03",X"01",X"00",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"09",X"0D",X"1B",X"1A",X"1E",X"14",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"C0",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"C1",X"F1",X"E7",X"4F",X"1F",X"3F",X"3F",X"7F",X"7C",X"F0",X"80",X"C0",X"60",X"00",
		X"FF",X"FF",X"FF",X"FE",X"FE",X"F1",X"F0",X"F0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"E0",X"E0",X"E0",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"60",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"01",X"3F",X"01",X"00",
		X"73",X"73",X"67",X"E7",X"EF",X"EF",X"C6",X"C6",X"C0",X"80",X"00",X"80",X"C0",X"A0",X"F0",X"78",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"03",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"03",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"06",X"06",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"51",X"AB",X"7B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"F0",X"F8",X"FC",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"30",X"39",X"3F",X"1E",X"14",X"00",X"00",X"00",
		X"07",X"0F",X"0F",X"1F",X"3C",X"30",X"58",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"F0",X"C0",X"03",X"06",X"0F",X"CC",X"E8",X"D8",X"70",X"60",X"40",X"00",X"00",X"00",X"00",
		X"00",X"20",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"20",X"30",X"38",X"1C",X"17",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"68",
		X"0E",X"07",X"03",X"01",X"00",X"00",X"00",X"C0",X"F8",X"3E",X"1F",X"0D",X"00",X"01",X"01",X"00",
		X"00",X"80",X"C0",X"E0",X"70",X"3C",X"1E",X"0F",X"03",X"31",X"F8",X"FC",X"FD",X"3F",X"1F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"60",X"30",X"F8",X"84",X"78",X"FC",
		X"F7",X"3F",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F1",X"E1",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"3F",X"06",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"FF",X"3F",X"03",X"00",X"00",X"00",X"00",X"00",X"07",X"0F",X"0F",X"1F",X"1F",X"1F",X"19",
		X"06",X"86",X"86",X"C4",X"44",X"E0",X"63",X"62",X"32",X"B3",X"FB",X"FB",X"7B",X"7B",X"33",X"B3",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"E0",
		X"00",X"00",X"87",X"FF",X"FF",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"38",X"70",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"01",X"04",X"03",X"04",X"01",
		X"B8",X"00",X"6C",X"06",X"03",X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"85",
		X"00",X"0C",X"0C",X"0C",X"18",X"18",X"98",X"B8",X"B0",X"70",X"60",X"60",X"C0",X"C0",X"E0",X"80",
		X"01",X"03",X"07",X"00",X"00",X"00",X"00",X"02",X"06",X"0E",X"1F",X"39",X"F0",X"C0",X"00",X"00",
		X"7E",X"B6",X"AF",X"C7",X"FF",X"FF",X"F8",X"FB",X"FB",X"FD",X"7F",X"7F",X"7F",X"3E",X"3E",X"1E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"01",X"0F",X"02",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"60",X"FC",X"1F",X"03",X"00",X"00",
		X"38",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"C1",X"C1",X"E1",X"E1",X"E1",X"DF",X"CF",X"EB",X"F1",X"FC",X"FF",X"CF",
		X"00",X"00",X"E0",X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"03",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",
		X"30",X"10",X"10",X"10",X"10",X"10",X"10",X"30",X"20",X"20",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",
		X"5F",X"BF",X"BF",X"BF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"C0",X"C0",X"00",
		X"78",X"7E",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3C",X"00",X"10",X"09",X"01",
		X"00",X"00",X"00",X"80",X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"60",X"20",X"50",X"D0",X"18",
		X"02",X"03",X"03",X"03",X"03",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"03",X"03",X"03",X"01",
		X"70",X"30",X"30",X"F0",X"F0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"C0",X"C0",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"19",X"11",X"13",X"03",X"03",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"02",X"00",X"00",X"00",
		X"80",X"00",X"81",X"82",X"84",X"C1",X"C0",X"C0",X"E0",X"E0",X"E0",X"E0",X"C0",X"00",X"00",X"20",
		X"18",X"08",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"02",X"02",X"02",X"03",X"03",X"03",X"03",X"07",X"07",X"07",X"07",X"07",X"07",X"03",X"01",
		X"10",X"10",X"10",X"10",X"30",X"30",X"F0",X"F0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"C0",X"80",
		X"02",X"03",X"06",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"9B",X"17",X"3F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",X"FB",X"F3",X"72",X"62",X"01",
		X"F0",X"E0",X"C0",X"E0",X"E0",X"E0",X"F0",X"F0",X"F0",X"F1",X"F0",X"E0",X"80",X"80",X"00",X"00",
		X"C0",X"40",X"60",X"20",X"30",X"10",X"10",X"08",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"07",X"07",X"06",X"07",X"07",X"07",X"03",X"01",
		X"40",X"40",X"40",X"60",X"70",X"70",X"70",X"70",X"30",X"20",X"60",X"E0",X"E0",X"E0",X"C0",X"80",
		X"06",X"04",X"04",X"14",X"24",X"18",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"07",X"0F",X"1F",X"3F",X"3F",X"7F",X"7F",X"7F",X"7D",X"79",X"71",X"62",X"42",X"62",X"22",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"25",X"1C",X"09",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"01",X"01",X"04",X"20",X"C0",X"70",X"D0",X"68",X"DC",
		X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"01",X"08",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"02",X"00",X"22",X"15",X"1F",X"0B",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"40",X"00",X"00",X"40",X"80",X"02",X"85",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"40",X"00",X"00",X"20",X"00",X"00",X"00",
		X"02",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"97",X"0B",X"21",X"11",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"DF",X"EF",X"E7",X"7B",X"91",X"CB",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EA",X"F4",X"BF",X"9F",X"BF",X"F5",X"F3",X"45",X"01",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"4E",X"9C",X"AF",X"3E",X"F4",X"7B",X"7F",X"ED",X"90",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"80",X"00",X"20",X"C0",X"80",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"08",X"00",X"01",X"00",X"0E",
		X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"04",X"20",X"00",X"00",X"00",X"04",X"22",X"1B",
		X"00",X"02",X"01",X"85",X"00",X"20",X"0C",X"06",X"28",X"02",X"10",X"89",X"5C",X"70",X"63",X"28",
		X"83",X"43",X"13",X"4D",X"AD",X"7F",X"7F",X"67",X"3B",X"BF",X"79",X"34",X"F8",X"FD",X"EB",X"E8",
		X"33",X"79",X"7F",X"A7",X"B6",X"FF",X"FF",X"6B",X"91",X"C3",X"DB",X"A7",X"F3",X"F9",X"69",X"F5",
		X"E8",X"C0",X"C0",X"E1",X"F5",X"F8",X"F1",X"B9",X"EB",X"EA",X"B7",X"C7",X"CB",X"E9",X"FD",X"FF",
		X"00",X"00",X"40",X"00",X"44",X"80",X"90",X"02",X"00",X"20",X"40",X"69",X"B2",X"A6",X"F1",X"F5",
		X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"10",X"02",X"00",X"40",X"80",X"40",X"90",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"31",X"D7",X"C2",X"86",X"24",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",
		X"66",X"F7",X"7E",X"FF",X"FF",X"FF",X"EF",X"6D",X"7E",X"36",X"01",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FB",X"ED",X"F5",X"F0",X"F9",X"E4",X"90",X"80",X"00",X"60",X"00",X"00",X"00",X"00",X"00",
		X"EF",X"E7",X"F7",X"F3",X"DB",X"CF",X"5D",X"18",X"0E",X"1F",X"1D",X"28",X"05",X"00",X"00",X"00",
		X"EF",X"FF",X"FB",X"FF",X"FF",X"EB",X"DD",X"99",X"4F",X"00",X"80",X"40",X"00",X"00",X"00",X"00",
		X"F2",X"E8",X"CC",X"EA",X"C0",X"20",X"80",X"80",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
