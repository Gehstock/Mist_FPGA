----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    21:49:44 12/03/2009 
-- Design Name: 
-- Module Name:    BMP - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

---- Uncomment the following library declaration if instantiating
---- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity BMP is
end BMP;

architecture Behavioral of BMP is

begin

-- Header
-- MAGIC NUMBER   : 2 octets 'BM'
-- Size of bitmap : 4 octets
-- Reserved       : 2 octets
-- Reserved       : 2 octets
-- Offset         : 4 octets



end Behavioral;

