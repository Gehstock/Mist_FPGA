library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity tropical_chr_bit2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of tropical_chr_bit2 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"61",X"35",X"72",X"F1",X"96",X"D9",X"DB",X"6A",X"FF",X"FF",X"FF",X"FE",X"F5",X"E8",X"73",X"E6",
		X"FF",X"FF",X"FF",X"BF",X"5F",X"1F",X"7F",X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FB",X"FF",X"FE",
		X"7C",X"BE",X"FE",X"FD",X"ED",X"BF",X"FF",X"FF",X"3D",X"9C",X"98",X"6C",X"74",X"E0",X"FB",X"F8",
		X"6F",X"FF",X"FF",X"BF",X"BF",X"3F",X"3F",X"1F",X"FF",X"FF",X"FF",X"FF",X"FC",X"FF",X"FD",X"FF",
		X"FD",X"E3",X"FA",X"77",X"FD",X"F2",X"FF",X"FF",X"DF",X"BF",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"03",X"03",X"03",X"01",X"01",
		X"FE",X"FF",X"FF",X"FB",X"FC",X"FF",X"FC",X"FE",X"9B",X"53",X"85",X"D3",X"E3",X"C9",X"D1",X"6D",
		X"FF",X"FF",X"EF",X"CF",X"DF",X"BF",X"BF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"F5",X"FB",
		X"3C",X"F0",X"E8",X"C0",X"80",X"90",X"F8",X"F8",X"01",X"01",X"01",X"03",X"03",X"07",X"07",X"0F",
		X"F8",X"D0",X"80",X"80",X"C0",X"C0",X"C0",X"E0",X"0F",X"0F",X"17",X"17",X"1A",X"1B",X"39",X"33",
		X"C0",X"C8",X"80",X"A0",X"40",X"80",X"40",X"80",X"3F",X"1F",X"1F",X"0E",X"1F",X"1D",X"1F",X"1F",
		X"98",X"38",X"7C",X"FC",X"FC",X"E0",X"04",X"0C",X"1F",X"1D",X"1D",X"1E",X"1E",X"0F",X"0F",X"0F",
		X"0C",X"9C",X"FE",X"7E",X"7E",X"7E",X"3E",X"3E",X"2F",X"0F",X"4F",X"AF",X"9F",X"07",X"07",X"07",
		X"BE",X"9F",X"FE",X"9E",X"9E",X"8E",X"8E",X"0E",X"07",X"07",X"07",X"07",X"07",X"03",X"03",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"1E",X"1C",X"1C",X"1C",X"1C",X"18",X"38",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"01",X"01",X"0E",X"1A",X"01",X"00",X"00",
		X"30",X"F0",X"F0",X"90",X"90",X"88",X"04",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"A7",X"00",X"00",X"00",X"00",X"00",X"0E",X"FB",X"4D",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"06",X"BF",X"11",X"00",
		X"00",X"00",X"00",X"6C",X"97",X"C2",X"00",X"00",X"00",X"00",X"00",X"0C",X"BF",X"09",X"50",X"00",
		X"00",X"00",X"01",X"1E",X"F4",X"40",X"10",X"00",X"01",X"00",X"00",X"A1",X"14",X"BB",X"CD",X"87",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"02",X"07",X"04",X"00",
		X"00",X"00",X"00",X"40",X"40",X"80",X"00",X"01",X"11",X"1A",X"07",X"8E",X"04",X"02",X"11",X"31",
		X"00",X"00",X"00",X"80",X"41",X"62",X"C0",X"A0",X"40",X"02",X"04",X"0B",X"19",X"20",X"00",X"81",
		X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"48",X"48",X"5C",X"BC",X"F9",X"F3",X"E7",X"FF",X"FF",
		X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"10",X"08",X"01",X"02",X"0A",X"15",X"1B",X"00",X"00",
		X"00",X"80",X"00",X"C0",X"72",X"A6",X"6C",X"C0",X"C2",X"98",X"B4",X"FC",X"58",X"BC",X"66",X"00",
		X"01",X"0F",X"02",X"01",X"00",X"00",X"00",X"00",X"43",X"73",X"AE",X"4C",X"9D",X"9F",X"08",X"00",
		X"43",X"87",X"12",X"6D",X"D8",X"01",X"00",X"00",X"E9",X"D2",X"A2",X"E5",X"CF",X"CF",X"00",X"00",
		X"00",X"00",X"42",X"8C",X"1E",X"0C",X"A0",X"00",X"84",X"46",X"CF",X"BC",X"F9",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"12",X"21",X"06",X"0C",X"F8",X"DC",X"8D",X"2E",X"15",X"15",X"2B",X"09",
		X"00",X"40",X"20",X"41",X"02",X"0C",X"10",X"60",X"40",X"02",X"04",X"0B",X"19",X"20",X"00",X"81",
		X"00",X"08",X"04",X"16",X"0C",X"04",X"08",X"00",X"01",X"00",X"08",X"14",X"0E",X"1E",X"00",X"00",
		X"00",X"01",X"40",X"28",X"30",X"40",X"40",X"A0",X"B0",X"10",X"0D",X"9E",X"7C",X"1B",X"06",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"08",X"00",X"00",X"00",X"00",X"40",X"40",X"81",
		X"00",X"00",X"00",X"00",X"10",X"20",X"70",X"20",X"1A",X"0F",X"0E",X"04",X"1D",X"B8",X"70",X"78",
		X"00",X"20",X"68",X"F0",X"40",X"00",X"00",X"01",X"C3",X"E7",X"C7",X"D7",X"AF",X"FF",X"FD",X"E3",
		X"00",X"00",X"00",X"80",X"00",X"00",X"80",X"00",X"80",X"02",X"86",X"CE",X"CC",X"80",X"C0",X"F1",
		X"48",X"5C",X"BC",X"F8",X"FE",X"FD",X"DE",X"EF",X"DF",X"8E",X"57",X"FE",X"D8",X"28",X"42",X"87",
		X"01",X"0F",X"02",X"01",X"00",X"00",X"C3",X"F1",X"E8",X"94",X"00",X"80",X"04",X"10",X"25",X"FF",
		X"43",X"87",X"12",X"6D",X"F9",X"CB",X"B1",X"E2",X"44",X"1E",X"0D",X"00",X"40",X"84",X"6C",X"FB",
		X"43",X"73",X"BC",X"79",X"F3",X"E2",X"07",X"88",X"00",X"00",X"02",X"80",X"44",X"48",X"84",X"FD",
		X"E9",X"D2",X"A2",X"E5",X"CF",X"8F",X"00",X"04",X"1D",X"23",X"76",X"FC",X"00",X"04",X"89",X"7F",
		X"48",X"5C",X"BC",X"F8",X"FE",X"FD",X"DE",X"EF",X"1D",X"23",X"76",X"FC",X"00",X"04",X"89",X"7F",
		X"00",X"00",X"00",X"40",X"88",X"51",X"E3",X"FF",X"43",X"87",X"12",X"6D",X"D3",X"1E",X"7C",X"FF",
		X"00",X"00",X"00",X"00",X"40",X"00",X"80",X"FF",X"43",X"76",X"BF",X"7D",X"4F",X"22",X"74",X"FF",
		X"00",X"00",X"00",X"00",X"04",X"09",X"1E",X"FF",X"00",X"00",X"00",X"00",X"82",X"1D",X"7F",X"FF",
		X"00",X"00",X"00",X"00",X"82",X"1D",X"7B",X"FF",X"00",X"00",X"00",X"00",X"41",X"B8",X"DE",X"FF",
		X"00",X"00",X"00",X"00",X"20",X"90",X"38",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"C3",X"F1",
		X"01",X"0F",X"02",X"01",X"04",X"09",X"1C",X"FF",X"00",X"00",X"00",X"00",X"01",X"C3",X"B1",X"E2",
		X"00",X"00",X"1C",X"79",X"F3",X"E2",X"07",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"C3",X"F1",
		X"00",X"00",X"00",X"80",X"C0",X"80",X"00",X"04",X"00",X"00",X"00",X"00",X"01",X"C3",X"B1",X"E2",
		X"5F",X"33",X"E7",X"76",X"DF",X"7E",X"ED",X"DF",X"FB",X"F2",X"63",X"A7",X"EE",X"77",X"AC",X"F9",
		X"C3",X"C7",X"9B",X"DF",X"FF",X"CF",X"DB",X"EE",X"00",X"18",X"20",X"F4",X"D9",X"5B",X"FD",X"EF",
		X"00",X"00",X"00",X"80",X"00",X"80",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"A0",X"B0",X"E8",X"78",X"E8",X"DF",X"7F",X"00",X"05",X"0D",X"17",X"1E",X"17",X"FB",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"5C",X"EC",X"7F",X"FA",X"67",X"F7",X"9D",X"03",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"87",X"CC",X"BE",X"F7",X"FF",X"7A",X"30",X"DC",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"11",X"7A",X"F3",X"EF",X"FF",X"FF",X"6E",X"B8",X"F7",
		X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"83",X"87",X"C7",X"6F",X"CD",X"EB",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"07",X"0F",X"1F",X"37",X"FF",X"FE",X"FF",X"F3",X"D8",X"B2",X"FD",X"FB",X"FF",
		X"1D",X"39",X"7C",X"7E",X"FC",X"FB",X"DF",X"FF",X"B6",X"E1",X"F6",X"3F",X"F3",X"7C",X"EB",X"FF",
		X"F4",X"FE",X"FF",X"7F",X"FD",X"FC",X"F9",X"F2",X"FB",X"77",X"F6",X"F4",X"E2",X"0D",X"03",X"FF",
		X"80",X"D0",X"DA",X"D7",X"DF",X"BE",X"FC",X"DC",X"E9",X"69",X"DB",X"4F",X"7F",X"BB",X"F7",X"E7",
		X"02",X"01",X"40",X"28",X"70",X"38",X"5C",X"38",X"83",X"C7",X"1F",X"AF",X"F7",X"E7",X"BD",X"7E",
		X"F8",X"DC",X"8D",X"2E",X"15",X"15",X"FB",X"79",X"FF",X"F5",X"FE",X"FD",X"F6",X"D9",X"BD",X"0F",
		X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"FF",X"00",X"01",X"01",X"03",X"07",X"07",X"07",X"0F",
		X"01",X"03",X"07",X"E3",X"F7",X"CF",X"FE",X"FF",X"80",X"80",X"B0",X"DC",X"B8",X"5C",X"F8",X"F0",
		X"C3",X"C7",X"CA",X"60",X"F8",X"F4",X"FA",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FB",X"72",X"63",X"47",X"02",X"00",X"20",X"40",X"00",X"18",X"20",X"80",X"40",X"00",X"00",X"00",
		X"87",X"CF",X"FD",X"6E",X"BF",X"77",X"21",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",X"EF",X"EF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"26",X"9B",X"34",X"A0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"21",X"09",X"42",X"09",
		X"00",X"00",X"00",X"00",X"00",X"00",X"12",X"40",X"3E",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"90",X"66",X"19",X"00",X"00",X"00",X"00",X"01",X"11",X"44",X"19",X"C6",X"6C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"AE",X"5B",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"AC",X"00",
		X"00",X"08",X"40",X"12",X"AD",X"EB",X"BF",X"6A",X"00",X"04",X"51",X"A4",X"E8",X"B8",X"5E",X"0A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"41",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"43",X"10",X"04",X"93",X"20",X"35",X"6F",X"BE",X"05",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"20",X"84",X"D1",X"00",X"00",X"00",X"00",X"00",X"10",X"02",X"4C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"4B",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"7F",X"3F",X"BF",X"BF",X"BF",X"BF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"F0",X"FC",X"FE",X"FC",X"F0",X"C0",
		X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"18",X"63",X"04",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"78",X"F1",X"EE",X"FC",X"68",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"1C",X"36",X"71",X"F8",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1B",X"3F",X"66",X"0C",X"0F",X"1C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"43",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"E0",X"04",X"03",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"04",X"03",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1E",X"F8",X"44",X"80",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"18",X"7C",X"3F",X"3F",X"7B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7C",X"08",X"FC",X"F8",X"9C",X"2E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"A9",X"67",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"FC",X"68",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7E",X"2C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EC",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"F1",X"C3",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"E9",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",
		X"00",X"00",X"01",X"67",X"CB",X"FF",X"FF",X"73",X"00",X"00",X"00",X"00",X"00",X"00",X"DB",X"FF",
		X"00",X"00",X"C6",X"7C",X"FF",X"EE",X"77",X"C3",X"00",X"00",X"00",X"00",X"00",X"01",X"EF",X"FE",
		X"00",X"00",X"0C",X"F9",X"F0",X"C0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"04",X"ED",X"07",
		X"00",X"00",X"A0",X"79",X"03",X"03",X"21",X"C3",X"00",X"00",X"00",X"00",X"00",X"00",X"27",X"DF",
		X"00",X"10",X"58",X"E7",X"DF",X"9F",X"C7",X"EF",X"00",X"00",X"00",X"00",X"26",X"73",X"C3",X"1C",
		X"00",X"40",X"98",X"3C",X"FC",X"FC",X"98",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",
		X"00",X"00",X"00",X"12",X"66",X"FF",X"AF",X"F9",X"04",X"08",X"FC",X"CC",X"F8",X"7C",X"10",X"F8",
		X"00",X"00",X"00",X"00",X"C0",X"E0",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"05",X"03",X"07",X"0E",X"18",X"06",X"1F",X"3B",X"17",X"32",X"7F",X"7C",
		X"00",X"29",X"42",X"EF",X"FF",X"FF",X"FF",X"FF",X"06",X"1B",X"FF",X"FF",X"E7",X"F3",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"02",X"40",X"00",X"10",X"00",X"80",
		X"00",X"00",X"0C",X"1B",X"1E",X"BC",X"64",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"01",X"07",X"07",X"03",X"00",
		X"00",X"00",X"00",X"00",X"03",X"07",X"03",X"00",X"00",X"01",X"79",X"B7",X"FF",X"FA",X"9F",X"DF",
		X"00",X"00",X"00",X"00",X"00",X"04",X"3A",X"71",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"24",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"74",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3D",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"28",
		X"00",X"00",X"00",X"00",X"60",X"58",X"F1",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"18",X"5E",X"07",X"9E",X"27",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"12",X"E6",X"C1",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"87",X"C7",X"29",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"23",X"88",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"72",X"2C",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"09",X"07",X"04",X"1E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"18",X"C0",X"26",X"8F",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"7F",X"06",X"BE",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"E7",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C3",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"9F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C7",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"0C",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"13",X"FE",X"CE",X"97",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"08",X"1C",X"7C",X"F9",X"FF",X"DD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",
		X"00",X"00",X"00",X"10",X"F3",X"E4",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",
		X"00",X"00",X"00",X"00",X"C1",X"FB",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"11",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C3",X"EF",X"FF",X"FF",
		X"00",X"00",X"00",X"C0",X"FC",X"3C",X"FC",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"03",X"0F",X"0F",X"07",
		X"00",X"00",X"00",X"00",X"00",X"06",X"0F",X"07",X"00",X"00",X"02",X"F3",X"2F",X"FF",X"F4",X"9F",
		X"00",X"00",X"00",X"00",X"24",X"CD",X"FF",X"5E",X"00",X"08",X"10",X"FC",X"CC",X"F8",X"7C",X"10",
		X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"0B",X"07",X"0F",X"00",X"00",X"00",X"3F",X"77",X"2F",X"65",X"FF",
		X"00",X"00",X"00",X"52",X"AF",X"FF",X"FF",X"FF",X"00",X"0C",X"06",X"FF",X"FF",X"E7",X"F3",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"04",X"80",X"00",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"1F",X"1F",X"17",X"04",X"00",X"00",X"00",X"00",X"C0",X"F0",X"7C",X"3E",X"1E",X"0F",
		X"02",X"2F",X"3F",X"1D",X"1F",X"0F",X"08",X"1C",X"79",X"FF",X"FF",X"FF",X"FF",X"FC",X"FF",X"3B",
		X"FF",X"FB",X"AE",X"58",X"14",X"40",X"A0",X"F5",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"7E",X"7C",
		X"7E",X"FB",X"F4",X"F8",X"F8",X"F0",X"E0",X"E1",X"00",X"93",X"6F",X"1F",X"3F",X"7F",X"FF",X"FE",
		X"D3",X"E0",X"F5",X"FF",X"DE",X"3D",X"7C",X"3C",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",
		X"72",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"73",X"FB",X"FD",X"FD",X"FC",X"FC",X"F8",X"F8",
		X"FC",X"F8",X"F8",X"F0",X"E1",X"C3",X"C3",X"81",X"1E",X"0F",X"17",X"7B",X"FB",X"F0",X"C0",X"80",
		X"00",X"00",X"F0",X"F8",X"F8",X"70",X"00",X"00",X"03",X"03",X"03",X"2F",X"5E",X"38",X"4C",X"18",
		X"81",X"81",X"00",X"00",X"00",X"00",X"00",X"00",X"F3",X"F7",X"E7",X"0F",X"9F",X"DF",X"FF",X"FF",
		X"E3",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"00",X"C0",X"C0",X"E0",X"E0",X"E0",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"07",X"0F",X"1A",X"06",X"1C",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"30",X"9F",X"3F",X"9F",X"7B",X"17",X"41",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0E",X"DF",X"E3",X"41",X"88",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"7F",X"9E",X"FB",X"78",X"FC",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"8E",X"37",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"B3",X"0F",X"07",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"06",X"FE",X"F0",X"E3",X"87",X"E4",X"C8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"07",X"C1",X"FF",X"EF",X"39",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"80",X"C0",X"E0",X"E4",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"03",X"03",X"07",X"06",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"58",X"EB",X"C7",X"93",X"3D",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"6F",X"FF",X"F3",X"EB",X"F9",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"04",X"BF",X"F8",X"60",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"10",X"BC",X"1F",X"00",X"00",X"04",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"BF",X"7E",X"38",X"0C",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"26",X"72",X"C3",X"1C",X"7F",X"9F",X"06",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"26",X"FC",X"9D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"38",X"79",X"F3",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"A0",X"E7",X"DC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"E3",X"F7",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"11",X"30",X"FC",X"E7",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"0F",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"1F",X"00",X"00",X"00",X"00",X"00",X"6F",X"FF",X"EF",
		X"00",X"00",X"00",X"00",X"00",X"48",X"9B",X"FF",X"00",X"00",X"00",X"20",X"60",X"CC",X"F8",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"02",X"00",X"00",X"01",X"17",X"0E",X"00",X"00",X"00",X"00",X"00",X"6F",X"DF",X"CB",
		X"20",X"00",X"00",X"40",X"02",X"2F",X"FF",X"FF",X"80",X"00",X"00",X"00",X"00",X"FF",X"FF",X"E7",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"05",X"80",X"19",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"71",X"EE",X"7C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"2C",X"62",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"7C",X"72",X"B0",X"98",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"18",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"27",X"1C",X"12",X"78",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"0C",X"1F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"7F",X"06",X"7E",X"FD",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"0F",X"1F",X"36",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"1E",X"3C",X"6A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"7C",X"FF",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"3C",X"7F",X"8E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"FF",X"3C",X"F6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"1C",X"6E",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"67",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"06",X"FC",X"E0",X"C3",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"00",X"07",X"C1",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"07",X"0F",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"A0",X"CE",X"AF",X"3E",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"DF",X"FF",X"CF",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"08",X"7F",X"F4",X"F0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"20",X"BA",X"1D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"0F",X"BF",X"7E",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"86",X"C3",X"C1",X"18",X"7F",X"F6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"00",X"C0",X"E0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"3B",X"00",X"00",X"00",X"00",X"00",X"00",X"DF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"39",X"00",X"00",X"00",X"00",X"20",X"60",X"CC",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"7C",
		X"00",X"28",X"42",X"42",X"34",X"00",X"49",X"7F",X"06",X"02",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"02",X"40",X"00",X"10",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"7C",X"7E",X"3E",X"0C",X"04",X"00",X"00",X"7C",X"FC",X"F8",X"78",X"70",X"10",X"00",X"00",
		X"0F",X"0F",X"1F",X"1F",X"1F",X"3E",X"3E",X"7C",X"00",X"01",X"01",X"03",X"03",X"03",X"07",X"07",
		X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"80",X"E0",X"F0",X"F8",X"FE",X"FE",X"FF",
		X"FF",X"FF",X"F2",X"F0",X"E0",X"E0",X"C0",X"C0",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"03",X"03",X"07",X"07",X"0F",X"0F",X"1F",X"1F",
		X"1F",X"3F",X"3F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",X"6F",X"07",X"06",X"02",X"00",
		X"00",X"40",X"70",X"F8",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"FC",X"FC",X"F8",
		X"F8",X"F0",X"E0",X"E0",X"E0",X"E0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"03",
		X"03",X"07",X"07",X"0F",X"0F",X"1F",X"1F",X"1F",X"3F",X"3F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"7F",X"7F",X"3E",X"1C",X"00",X"00",X"00",X"78",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",
		X"FF",X"FE",X"FE",X"FE",X"FC",X"FC",X"F8",X"F8",X"F0",X"F0",X"F0",X"E0",X"E0",X"C0",X"C0",X"80",
		X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"3F",X"3F",X"7C",X"7C",X"FC",X"F8",X"F8",
		X"F0",X"F0",X"E0",X"E0",X"C0",X"40",X"00",X"00",X"F8",X"F0",X"F0",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"20",X"38",X"78",X"7C",X"7C",X"F8",X"F8",X"F0",X"F0",X"F0",X"E0",X"E0",X"C0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"40",X"9D",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"3A",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"20",X"30",X"FC",X"F7",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"74",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"03",X"0F",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"06",X"93",X"EF",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"80",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"36",X"7F",X"9F",X"FC",X"F7",X"3C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"A7",X"CF",X"FF",X"F4",X"7E",X"3C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"86",X"F6",X"03",X"00",X"00",X"01",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"93",X"EF",X"0E",X"0F",X"86",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"38",X"F0",X"C7",X"1F",X"3F",X"07",X"8E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"F0",X"38",X"FC",X"FC",X"38",X"0C",
		X"00",X"01",X"06",X"06",X"0C",X"0B",X"0F",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"52",X"82",X"84",X"02",X"49",X"00",X"0C",X"06",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"04",X"80",X"00",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"60",X"C1",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0A",X"07",X"87",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"03",X"83",X"12",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"07",X"87",X"C7",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"20",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"38",X"70",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"1E",X"F8",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"40",X"80",X"00",X"18",X"78",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"F6",X"7C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"03",X"67",X"C7",X"83",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C3",X"E1",X"DC",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B6",X"C1",X"F6",X"A6",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"F0",X"F8",X"E4",X"B0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"DC",X"0E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"03",X"02",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"E0",X"93",X"47",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"1F",X"03",X"DF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"1E",X"0C",X"7A",X"33",X"E0",X"C4",X"BF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"74",X"FD",X"7F",X"F6",X"78",X"FE",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F5",X"CF",X"F3",X"7F",X"3F",X"9D",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"F9",X"EE",X"C0",X"C0",X"00",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"C0",X"E8",X"74",X"03",X"01",X"00",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"3F",X"7C",X"F9",X"E3",X"F2",X"E0",X"78",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"07",X"61",X"FF",X"F6",X"3F",X"0F",X"19",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"E0",X"E4",X"F8",X"E0",
		X"00",X"19",X"33",X"7F",X"7F",X"79",X"3D",X"0F",X"00",X"00",X"00",X"00",X"6D",X"FF",X"3F",X"FC",
		X"40",X"DF",X"FF",X"F7",X"BB",X"E1",X"F8",X"FF",X"00",X"00",X"00",X"00",X"4F",X"97",X"FF",X"EC",
		X"80",X"38",X"F8",X"60",X"F0",X"E0",X"F0",X"F0",X"00",X"00",X"00",X"84",X"ED",X"07",X"00",X"00",
		X"00",X"01",X"03",X"03",X"01",X"63",X"07",X"03",X"00",X"00",X"00",X"00",X"27",X"DF",X"3C",X"1E",
		X"58",X"EF",X"DF",X"9F",X"C7",X"EF",X"FF",X"F8",X"00",X"00",X"13",X"39",X"C3",X"1C",X"7F",X"9F",
		X"0C",X"7E",X"FE",X"FE",X"CC",X"86",X"FE",X"FC",X"00",X"00",X"00",X"80",X"E0",X"F0",X"F8",X"F8",
		X"00",X"00",X"00",X"02",X"1C",X"1C",X"39",X"17",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"6C",X"FF",X"FE",X"E7",X"37",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"F2",X"FF",X"9E",X"C7",X"FE",X"FE",X"B4",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"0C",X"1E",X"78",
		X"00",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"02",X"3B",X"77",X"3E",X"FF",X"6F",X"DF",X"CB",
		X"20",X"00",X"00",X"00",X"02",X"22",X"84",X"85",X"9B",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E7",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"08",X"00",X"00",X"00",
		X"3E",X"3E",X"7E",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"9E",X"9C",X"84",X"00",X"00",
		X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"80",X"01",X"01",X"03",X"03",X"07",X"07",X"0F",X"0F",
		X"1F",X"1F",X"3F",X"3F",X"7F",X"7F",X"FF",X"FF",X"7F",X"77",X"37",X"03",X"03",X"01",X"00",X"00",
		X"00",X"10",X"3C",X"3E",X"7E",X"7F",X"FF",X"FE",X"FE",X"FE",X"FC",X"FC",X"FC",X"F8",X"F8",X"F8",
		X"F0",X"F0",X"F0",X"E0",X"E0",X"E0",X"C0",X"C0",X"C0",X"80",X"80",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"03",X"03",X"07",X"07",X"0F",X"0F",
		X"0F",X"1F",X"1F",X"3E",X"3E",X"7E",X"7C",X"FC",X"00",X"20",X"38",X"78",X"7C",X"FC",X"F8",X"F8",
		X"F0",X"F0",X"E0",X"E0",X"C0",X"C0",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"07",X"0F",X"0F",X"1F",X"1F",X"1F",X"3F",X"3F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"80",X"E0",X"E0",X"FC",X"FE",X"FE",X"FF",X"FF",X"FE",X"FE",X"FC",X"FC",X"F8",X"F8",X"F8",
		X"F0",X"F0",X"E0",X"E0",X"C0",X"C0",X"C0",X"80",X"03",X"07",X"07",X"0F",X"0F",X"1F",X"1F",X"1F",
		X"FF",X"FF",X"7F",X"7F",X"3E",X"1E",X"04",X"00",X"FF",X"FE",X"FE",X"9E",X"9C",X"84",X"C0",X"E0",
		X"E0",X"F0",X"F0",X"E0",X"E0",X"C0",X"C0",X"80",X"FF",X"FF",X"7F",X"0E",X"0E",X"02",X"00",X"00",
		X"00",X"20",X"38",X"7C",X"7E",X"FE",X"FF",X"FF",X"F6",X"F2",X"E0",X"E0",X"C0",X"C0",X"E0",X"E0",
		X"F0",X"F0",X"60",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"01",X"01",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"1E",X"1F",X"7C",X"F8",X"FB",X"E7",X"4F",X"5E",X"1C",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
