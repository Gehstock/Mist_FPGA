library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_PGM_0 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_PGM_0 is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"C3",X"C8",X"B1",X"C3",X"67",X"32",X"FE",X"00",X"C3",X"24",X"31",X"00",X"C3",X"C7",X"17",X"00",
		X"C3",X"1B",X"16",X"00",X"C3",X"2D",X"1A",X"00",X"C3",X"DF",X"19",X"00",X"C3",X"82",X"0F",X"00",
		X"C3",X"A6",X"0E",X"00",X"C3",X"A3",X"32",X"00",X"C3",X"91",X"34",X"00",X"C3",X"8C",X"19",X"00",
		X"C3",X"97",X"31",X"00",X"C3",X"C2",X"19",X"00",X"C3",X"45",X"0B",X"1A",X"BE",X"D8",X"C0",X"13",
		X"23",X"1A",X"BE",X"D8",X"C0",X"13",X"23",X"1A",X"BE",X"C9",X"21",X"00",X"40",X"11",X"00",X"04",
		X"06",X"0F",X"18",X"33",X"21",X"00",X"44",X"11",X"00",X"04",X"18",X"29",X"21",X"F0",X"4F",X"11",
		X"40",X"50",X"06",X"40",X"3E",X"00",X"77",X"12",X"23",X"13",X"10",X"FA",X"C9",X"21",X"00",X"4C",
		X"11",X"20",X"00",X"18",X"10",X"21",X"80",X"40",X"11",X"00",X"03",X"06",X"0F",X"18",X"08",X"21",
		X"00",X"4C",X"11",X"D0",X"03",X"06",X"00",X"70",X"23",X"1B",X"7A",X"B3",X"20",X"F9",X"C9",X"DD",
		X"21",X"21",X"4C",X"11",X"26",X"4C",X"DD",X"7E",X"00",X"A7",X"28",X"08",X"DD",X"35",X"00",X"20",
		X"03",X"3E",X"01",X"12",X"DD",X"23",X"13",X"DD",X"7E",X"00",X"A7",X"28",X"11",X"DD",X"35",X"01",
		X"20",X"0C",X"DD",X"36",X"01",X"3C",X"DD",X"35",X"00",X"20",X"03",X"3E",X"01",X"12",X"2A",X"24",
		X"4C",X"13",X"7C",X"B5",X"C8",X"01",X"FF",X"FF",X"3F",X"ED",X"5A",X"20",X"06",X"3E",X"01",X"12",
		X"21",X"00",X"00",X"22",X"24",X"4C",X"C9",X"DD",X"21",X"00",X"04",X"EB",X"DD",X"19",X"EB",X"23",
		X"DD",X"23",X"77",X"DD",X"70",X"00",X"C6",X"02",X"2B",X"DD",X"2B",X"77",X"DD",X"70",X"00",X"3D",
		X"11",X"21",X"00",X"19",X"DD",X"19",X"77",X"DD",X"70",X"00",X"C6",X"02",X"2B",X"DD",X"2B",X"77",
		X"DD",X"70",X"00",X"C9",X"21",X"31",X"01",X"87",X"16",X"00",X"5F",X"19",X"5E",X"23",X"56",X"EB",
		X"5E",X"23",X"56",X"23",X"4E",X"23",X"DD",X"21",X"00",X"04",X"DD",X"19",X"7E",X"FE",X"00",X"C8",
		X"D6",X"30",X"FE",X"0A",X"38",X"01",X"3D",X"12",X"DD",X"71",X"00",X"13",X"23",X"DD",X"23",X"18",
		X"EB",X"6B",X"01",X"88",X"01",X"A6",X"01",X"BA",X"01",X"CE",X"01",X"E6",X"01",X"FE",X"01",X"0B",
		X"02",X"13",X"02",X"1B",X"02",X"28",X"02",X"32",X"02",X"3F",X"02",X"4E",X"02",X"5D",X"02",X"72",
		X"02",X"82",X"02",X"9A",X"02",X"AD",X"02",X"C2",X"02",X"DA",X"02",X"F1",X"02",X"07",X"03",X"1E",
		X"03",X"29",X"03",X"3D",X"03",X"52",X"03",X"6D",X"03",X"82",X"03",X"A2",X"41",X"03",X"50",X"55",
		X"53",X"48",X"40",X"4F",X"4E",X"4C",X"59",X"40",X"31",X"40",X"50",X"4C",X"41",X"59",X"45",X"52",
		X"40",X"42",X"55",X"54",X"54",X"4F",X"4E",X"00",X"A2",X"41",X"03",X"50",X"55",X"53",X"48",X"40",
		X"31",X"40",X"4F",X"52",X"40",X"32",X"40",X"50",X"4C",X"41",X"59",X"45",X"52",X"53",X"40",X"42",
		X"55",X"54",X"54",X"4F",X"4E",X"00",X"A8",X"41",X"0F",X"50",X"4C",X"41",X"59",X"45",X"52",X"40",
		X"4F",X"4E",X"45",X"40",X"53",X"54",X"41",X"52",X"54",X"00",X"A8",X"41",X"0F",X"50",X"4C",X"41",
		X"59",X"45",X"52",X"40",X"54",X"57",X"4F",X"40",X"53",X"54",X"41",X"52",X"54",X"00",X"A6",X"41",
		X"01",X"50",X"4C",X"41",X"59",X"45",X"52",X"40",X"4F",X"4E",X"45",X"40",X"47",X"41",X"4D",X"45",
		X"40",X"4F",X"56",X"45",X"52",X"00",X"A6",X"41",X"01",X"50",X"4C",X"41",X"59",X"45",X"52",X"40",
		X"54",X"57",X"4F",X"40",X"47",X"41",X"4D",X"45",X"40",X"4F",X"56",X"45",X"52",X"00",X"AA",X"41",
		X"01",X"47",X"41",X"4D",X"45",X"40",X"4F",X"56",X"45",X"52",X"00",X"41",X"40",X"0F",X"31",X"40",
		X"55",X"50",X"00",X"5A",X"40",X"0F",X"32",X"40",X"55",X"50",X"00",X"4B",X"40",X"0F",X"54",X"4F",
		X"50",X"40",X"53",X"43",X"4F",X"52",X"45",X"00",X"B8",X"43",X"01",X"43",X"52",X"45",X"44",X"49",
		X"54",X"00",X"B7",X"43",X"05",X"46",X"52",X"45",X"45",X"40",X"50",X"4C",X"41",X"59",X"00",X"1A",
		X"41",X"01",X"49",X"4E",X"53",X"45",X"52",X"54",X"40",X"43",X"4F",X"49",X"4E",X"00",X"AA",X"41",
		X"07",X"49",X"4E",X"53",X"45",X"52",X"54",X"40",X"43",X"4F",X"49",X"4E",X"00",X"89",X"41",X"05",
		X"42",X"4F",X"4E",X"55",X"53",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",
		X"40",X"00",X"E9",X"41",X"07",X"4E",X"45",X"58",X"54",X"40",X"50",X"41",X"54",X"54",X"45",X"52",
		X"4E",X"00",X"E6",X"40",X"01",X"3D",X"3D",X"4C",X"45",X"54",X"53",X"40",X"53",X"49",X"4E",X"47",
		X"40",X"41",X"40",X"53",X"4F",X"4E",X"47",X"3D",X"3D",X"00",X"48",X"41",X"07",X"52",X"55",X"4E",
		X"40",X"52",X"55",X"4E",X"40",X"50",X"4F",X"4E",X"50",X"4F",X"4B",X"4F",X"00",X"87",X"41",X"07",
		X"54",X"4F",X"40",X"45",X"41",X"54",X"40",X"54",X"48",X"45",X"40",X"46",X"52",X"55",X"49",X"54",
		X"53",X"00",X"47",X"43",X"0F",X"53",X"49",X"47",X"4D",X"41",X"40",X"45",X"4E",X"54",X"3B",X"49",
		X"4E",X"43",X"3B",X"3E",X"40",X"31",X"39",X"38",X"32",X"00",X"A6",X"41",X"0F",X"50",X"40",X"40",
		X"4F",X"40",X"40",X"4E",X"40",X"40",X"50",X"40",X"40",X"4F",X"40",X"40",X"4B",X"40",X"40",X"4F",
		X"00",X"87",X"41",X"07",X"31",X"40",X"50",X"4C",X"41",X"59",X"40",X"4F",X"4E",X"4C",X"59",X"40",
		X"31",X"30",X"30",X"59",X"45",X"4E",X"00",X"C7",X"41",X"01",X"32",X"40",X"50",X"4C",X"41",X"59",
		X"53",X"40",X"4A",X"55",X"53",X"54",X"40",X"32",X"30",X"30",X"59",X"45",X"4E",X"00",X"CD",X"40",
		X"0F",X"52",X"41",X"4E",X"4B",X"49",X"4E",X"47",X"00",X"09",X"41",X"0F",X"52",X"41",X"4E",X"4B",
		X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"53",X"43",X"4F",X"52",X"45",X"00",X"C7",X"41",X"07",
		X"4A",X"55",X"4D",X"50",X"40",X"42",X"4F",X"55",X"4E",X"44",X"40",X"41",X"52",X"4F",X"55",X"4E",
		X"44",X"00",X"05",X"42",X"07",X"57",X"49",X"54",X"48",X"40",X"59",X"4F",X"55",X"52",X"40",X"42",
		X"49",X"47",X"40",X"42",X"45",X"4C",X"4C",X"59",X"40",X"4F",X"55",X"54",X"00",X"E8",X"42",X"0F",
		X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",
		X"40",X"00",X"27",X"43",X"0F",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",
		X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"00",X"1A",X"47",X"0E",X"0F",X"07",X"07",X"07",
		X"07",X"A1",X"20",X"2F",X"36",X"0F",X"23",X"78",X"A1",X"20",X"2C",X"36",X"0F",X"23",X"13",X"1A",
		X"47",X"07",X"07",X"07",X"07",X"A1",X"20",X"29",X"36",X"0F",X"23",X"78",X"A1",X"20",X"26",X"36",
		X"0F",X"23",X"13",X"1A",X"47",X"07",X"07",X"07",X"07",X"A1",X"20",X"23",X"36",X"0F",X"23",X"78",
		X"A1",X"77",X"C9",X"77",X"23",X"78",X"A1",X"77",X"23",X"13",X"1A",X"47",X"07",X"07",X"07",X"07",
		X"A1",X"77",X"23",X"78",X"A1",X"77",X"23",X"13",X"1A",X"47",X"07",X"07",X"07",X"07",X"A1",X"77",
		X"18",X"DC",X"AF",X"06",X"06",X"21",X"3A",X"4C",X"77",X"23",X"10",X"FC",X"C9",X"3A",X"2D",X"4C",
		X"32",X"2E",X"4C",X"3A",X"2B",X"4C",X"32",X"2D",X"4C",X"2A",X"29",X"4C",X"22",X"2B",X"4C",X"21",
		X"2B",X"4C",X"3A",X"29",X"4C",X"A6",X"32",X"2F",X"4C",X"23",X"3A",X"2A",X"4C",X"A6",X"32",X"30",
		X"4C",X"3A",X"00",X"50",X"32",X"29",X"4C",X"3A",X"40",X"50",X"32",X"2A",X"4C",X"C9",X"3A",X"C0",
		X"50",X"47",X"E6",X"40",X"07",X"32",X"53",X"4E",X"78",X"06",X"00",X"E6",X"0F",X"26",X"00",X"6F",
		X"29",X"29",X"11",X"71",X"04",X"19",X"0E",X"02",X"11",X"6F",X"4E",X"7E",X"B7",X"28",X"18",X"3E",
		X"01",X"12",X"11",X"72",X"4E",X"ED",X"B0",X"11",X"76",X"4E",X"0E",X"02",X"ED",X"B0",X"3E",X"01",
		X"32",X"7A",X"4E",X"32",X"7B",X"4E",X"C9",X"3E",X"FF",X"32",X"6E",X"4E",X"3E",X"0B",X"C3",X"04",
		X"01",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"02",X"01",X"02",X"01",X"01",X"02",X"01",
		X"02",X"03",X"01",X"03",X"01",X"01",X"01",X"02",X"03",X"01",X"01",X"04",X"05",X"02",X"01",X"01",
		X"03",X"01",X"01",X"01",X"05",X"01",X"01",X"01",X"06",X"01",X"01",X"01",X"03",X"02",X"01",X"01",
		X"05",X"02",X"01",X"01",X"06",X"02",X"01",X"01",X"01",X"03",X"01",X"01",X"02",X"03",X"01",X"01",
		X"04",X"3A",X"80",X"50",X"47",X"E6",X"03",X"32",X"31",X"4C",X"78",X"E6",X"0C",X"0F",X"0F",X"32",
		X"32",X"4C",X"78",X"E6",X"30",X"0F",X"0F",X"0F",X"0F",X"32",X"33",X"4C",X"78",X"E6",X"40",X"07",
		X"07",X"32",X"52",X"4E",X"78",X"E6",X"3F",X"32",X"35",X"4C",X"78",X"07",X"07",X"E6",X"01",X"3E",
		X"01",X"32",X"34",X"4C",X"C9",X"3A",X"31",X"4C",X"21",X"FF",X"1A",X"87",X"16",X"00",X"5F",X"19",
		X"5E",X"23",X"56",X"21",X"36",X"4C",X"72",X"23",X"73",X"23",X"36",X"00",X"C9",X"3A",X"6E",X"4E",
		X"FE",X"FF",X"C8",X"FE",X"64",X"D0",X"3E",X"20",X"21",X"70",X"4E",X"11",X"00",X"50",X"ED",X"4B",
		X"72",X"4E",X"CD",X"34",X"05",X"3E",X"40",X"21",X"74",X"4E",X"11",X"00",X"50",X"ED",X"4B",X"76",
		X"4E",X"CD",X"34",X"05",X"3E",X"80",X"21",X"78",X"4E",X"11",X"00",X"50",X"ED",X"4B",X"7A",X"4E",
		X"CD",X"34",X"05",X"C9",X"EB",X"A6",X"EB",X"20",X"1A",X"7E",X"B7",X"C8",X"36",X"00",X"23",X"34",
		X"7E",X"91",X"D8",X"77",X"21",X"6E",X"4E",X"7E",X"80",X"77",X"CD",X"56",X"05",X"3E",X"0A",X"32",
		X"45",X"4E",X"C9",X"36",X"01",X"C9",X"0E",X"00",X"3A",X"6E",X"4E",X"B7",X"28",X"0F",X"FE",X"64",
		X"38",X"02",X"3E",X"63",X"D6",X"0A",X"38",X"03",X"0C",X"18",X"F9",X"C6",X"0A",X"11",X"00",X"04",
		X"21",X"BE",X"43",X"71",X"19",X"36",X"05",X"21",X"BF",X"43",X"77",X"19",X"36",X"05",X"C9",X"3A",
		X"33",X"4C",X"C6",X"01",X"32",X"39",X"4C",X"C9",X"3A",X"39",X"4C",X"47",X"3A",X"46",X"4C",X"3D",
		X"21",X"48",X"4C",X"70",X"20",X"02",X"06",X"00",X"23",X"70",X"C9",X"3E",X"08",X"CD",X"04",X"01",
		X"3E",X"00",X"32",X"7E",X"40",X"3E",X"05",X"32",X"7E",X"44",X"C9",X"3E",X"0F",X"32",X"7E",X"40",
		X"21",X"5A",X"40",X"06",X"04",X"77",X"23",X"10",X"FC",X"C9",X"AF",X"21",X"3A",X"4C",X"06",X"06",
		X"77",X"23",X"10",X"FC",X"21",X"60",X"40",X"11",X"79",X"40",X"3E",X"0F",X"06",X"06",X"77",X"12",
		X"23",X"13",X"10",X"FA",X"AF",X"2B",X"1B",X"77",X"12",X"C9",X"3A",X"47",X"4C",X"FE",X"01",X"20",
		X"05",X"21",X"3A",X"4C",X"18",X"03",X"21",X"3D",X"4C",X"11",X"40",X"4C",X"CD",X"3B",X"00",X"21",
		X"45",X"4C",X"36",X"00",X"D0",X"34",X"C9",X"21",X"44",X"4C",X"7E",X"2B",X"B6",X"C8",X"5E",X"23",
		X"56",X"21",X"00",X"00",X"22",X"43",X"4C",X"3A",X"47",X"4C",X"3D",X"20",X"05",X"21",X"3C",X"4C",
		X"18",X"03",X"21",X"3F",X"4C",X"AF",X"7B",X"86",X"27",X"77",X"2B",X"7A",X"8E",X"27",X"77",X"2B",
		X"3E",X"00",X"8E",X"27",X"77",X"3A",X"47",X"4C",X"3D",X"20",X"05",X"3A",X"4A",X"4C",X"18",X"03",
		X"3A",X"4B",X"4C",X"A7",X"20",X"33",X"11",X"36",X"4C",X"EB",X"7E",X"23",X"B6",X"23",X"B6",X"28",
		X"28",X"2B",X"2B",X"CD",X"3B",X"00",X"38",X"21",X"3A",X"47",X"4C",X"3D",X"20",X"0A",X"21",X"48",
		X"4C",X"3E",X"01",X"32",X"4A",X"4C",X"18",X"08",X"21",X"49",X"4C",X"3E",X"01",X"32",X"4B",X"4C",
		X"34",X"CD",X"51",X"34",X"3E",X"01",X"32",X"45",X"4E",X"3A",X"45",X"4C",X"A7",X"CC",X"DA",X"05",
		X"3A",X"47",X"4C",X"3D",X"20",X"08",X"11",X"3A",X"4C",X"21",X"60",X"40",X"18",X"06",X"11",X"3D",
		X"4C",X"21",X"79",X"40",X"CD",X"99",X"03",X"3A",X"45",X"4C",X"A7",X"C8",X"1B",X"1B",X"21",X"40",
		X"4C",X"1A",X"77",X"13",X"23",X"1A",X"77",X"13",X"23",X"1A",X"77",X"21",X"6C",X"40",X"1B",X"1B",
		X"CD",X"99",X"03",X"C9",X"31",X"F0",X"4F",X"AF",X"32",X"00",X"50",X"F3",X"ED",X"56",X"AF",X"32",
		X"03",X"50",X"32",X"45",X"4E",X"CD",X"B4",X"0A",X"3E",X"0C",X"32",X"46",X"4E",X"3E",X"01",X"32",
		X"20",X"4C",X"FB",X"3E",X"01",X"32",X"00",X"50",X"3A",X"20",X"4C",X"87",X"16",X"00",X"5F",X"21",
		X"31",X"0A",X"E5",X"21",X"DC",X"06",X"19",X"5E",X"23",X"56",X"EB",X"E9",X"E4",X"06",X"E7",X"06",
		X"EF",X"07",X"09",X"08",X"C3",X"00",X"00",X"21",X"CA",X"07",X"E5",X"21",X"FB",X"06",X"3A",X"40",
		X"4E",X"87",X"5F",X"16",X"00",X"19",X"5E",X"23",X"56",X"EB",X"E9",X"05",X"07",X"46",X"07",X"5D",
		X"07",X"5E",X"07",X"C9",X"07",X"CD",X"75",X"00",X"CD",X"D0",X"0D",X"3E",X"13",X"CD",X"04",X"01",
		X"3E",X"14",X"CD",X"04",X"01",X"21",X"26",X"07",X"11",X"00",X"4C",X"01",X"20",X"00",X"ED",X"B0",
		X"3E",X"01",X"32",X"47",X"4C",X"C9",X"98",X"14",X"98",X"14",X"98",X"14",X"98",X"14",X"98",X"14",
		X"98",X"14",X"98",X"14",X"98",X"0C",X"78",X"2C",X"78",X"43",X"78",X"5C",X"78",X"73",X"78",X"8C",
		X"78",X"A3",X"78",X"BC",X"78",X"CC",X"3A",X"0B",X"4E",X"FE",X"00",X"C8",X"CD",X"75",X"00",X"CD",
		X"FE",X"0D",X"3E",X"01",X"32",X"47",X"4C",X"3E",X"02",X"32",X"40",X"4E",X"C9",X"C9",X"3A",X"4D",
		X"4E",X"A7",X"C0",X"CD",X"75",X"00",X"CD",X"D0",X"0D",X"CD",X"F3",X"12",X"CD",X"34",X"34",X"AF",
		X"32",X"4C",X"4C",X"32",X"46",X"4C",X"3E",X"0A",X"32",X"4E",X"4C",X"32",X"66",X"4C",X"CF",X"CD",
		X"21",X"32",X"CD",X"FB",X"31",X"CD",X"F6",X"33",X"CD",X"96",X"33",X"3E",X"9F",X"32",X"64",X"4C",
		X"3E",X"26",X"32",X"65",X"4C",X"3E",X"F0",X"32",X"11",X"4C",X"3E",X"28",X"32",X"10",X"4C",X"3E",
		X"98",X"32",X"00",X"4C",X"3E",X"14",X"32",X"01",X"4C",X"AF",X"32",X"58",X"4C",X"32",X"57",X"4C",
		X"32",X"56",X"4C",X"32",X"4F",X"4C",X"32",X"3E",X"4E",X"3E",X"01",X"32",X"5A",X"4C",X"3E",X"08",
		X"32",X"4D",X"4C",X"3E",X"04",X"32",X"40",X"4E",X"C9",X"C9",X"3A",X"6E",X"4E",X"A7",X"28",X"13",
		X"3E",X"02",X"32",X"20",X"4C",X"AF",X"32",X"40",X"4E",X"32",X"41",X"4E",X"CD",X"75",X"00",X"CD",
		X"D0",X"0D",X"C9",X"3A",X"41",X"4E",X"A7",X"20",X"FA",X"3E",X"FF",X"32",X"41",X"4E",X"C9",X"3A",
		X"46",X"4C",X"A7",X"C8",X"3E",X"03",X"32",X"20",X"4C",X"32",X"C0",X"50",X"AF",X"32",X"3F",X"4E",
		X"32",X"50",X"4C",X"3E",X"03",X"32",X"45",X"4E",X"C9",X"AF",X"32",X"4A",X"4C",X"32",X"4B",X"4C",
		X"3E",X"01",X"32",X"4C",X"4C",X"AF",X"32",X"3F",X"4E",X"CD",X"F3",X"12",X"CD",X"88",X"05",X"CD",
		X"BA",X"05",X"3E",X"01",X"32",X"51",X"4C",X"32",X"52",X"4C",X"32",X"4E",X"4C",X"3A",X"46",X"4C",
		X"FE",X"01",X"CC",X"AB",X"05",X"3A",X"46",X"4C",X"FE",X"01",X"28",X"22",X"3A",X"47",X"4C",X"FE",
		X"01",X"20",X"04",X"3E",X"02",X"18",X"02",X"3E",X"03",X"CD",X"04",X"01",X"3E",X"60",X"32",X"21",
		X"4C",X"AF",X"32",X"26",X"4C",X"3A",X"26",X"4C",X"A7",X"28",X"FA",X"CD",X"75",X"00",X"3A",X"4E",
		X"4C",X"3D",X"CF",X"CD",X"21",X"32",X"CD",X"FB",X"31",X"CD",X"7E",X"34",X"CD",X"51",X"34",X"CD",
		X"96",X"33",X"CD",X"F6",X"33",X"3E",X"9F",X"32",X"64",X"4C",X"3E",X"26",X"32",X"65",X"4C",X"3E",
		X"F0",X"32",X"11",X"4C",X"3E",X"28",X"32",X"10",X"4C",X"3E",X"98",X"32",X"00",X"4C",X"3E",X"14",
		X"32",X"01",X"4C",X"AF",X"32",X"58",X"4C",X"32",X"57",X"4C",X"32",X"56",X"4C",X"32",X"4F",X"4C",
		X"3C",X"32",X"5A",X"4C",X"3E",X"08",X"32",X"4D",X"4C",X"AF",X"32",X"4C",X"4C",X"3C",X"32",X"66",
		X"4C",X"CD",X"F7",X"05",X"3A",X"4F",X"4C",X"A7",X"C2",X"34",X"0A",X"21",X"50",X"4C",X"7E",X"A7",
		X"28",X"E7",X"3E",X"64",X"32",X"50",X"4E",X"3E",X"02",X"32",X"45",X"4E",X"3E",X"01",X"32",X"4F",
		X"4E",X"AF",X"32",X"3F",X"4E",X"32",X"50",X"4C",X"3A",X"50",X"4E",X"A7",X"20",X"FA",X"AF",X"32",
		X"4F",X"4E",X"21",X"50",X"4C",X"36",X"00",X"3E",X"01",X"32",X"4C",X"4C",X"32",X"66",X"4C",X"CD",
		X"34",X"34",X"21",X"48",X"4C",X"3A",X"46",X"4C",X"FE",X"01",X"20",X"60",X"7E",X"A7",X"20",X"49",
		X"3E",X"0B",X"32",X"45",X"4E",X"CD",X"75",X"00",X"CD",X"6D",X"00",X"3E",X"06",X"CD",X"04",X"01",
		X"AF",X"32",X"45",X"4C",X"32",X"03",X"50",X"CD",X"9B",X"05",X"3E",X"02",X"32",X"22",X"4C",X"AF",
		X"32",X"27",X"4C",X"3A",X"27",X"4C",X"A7",X"28",X"FA",X"3A",X"46",X"4C",X"3D",X"20",X"06",X"CD",
		X"14",X"13",X"CD",X"75",X"00",X"3A",X"6E",X"4E",X"A7",X"20",X"04",X"3E",X"01",X"18",X"02",X"3E",
		X"02",X"32",X"20",X"4C",X"AF",X"32",X"46",X"4C",X"C9",X"35",X"3E",X"01",X"32",X"22",X"4C",X"AF",
		X"32",X"27",X"4C",X"3A",X"27",X"4C",X"A7",X"28",X"FA",X"C3",X"5E",X"08",X"3A",X"47",X"4C",X"FE",
		X"01",X"C2",X"CE",X"09",X"7E",X"35",X"FE",X"00",X"CA",X"9C",X"09",X"23",X"7E",X"FE",X"FF",X"28",
		X"22",X"CD",X"75",X"00",X"CD",X"6D",X"00",X"3E",X"02",X"32",X"47",X"4C",X"3A",X"52",X"4E",X"A7",
		X"20",X"05",X"3E",X"01",X"32",X"03",X"50",X"3A",X"52",X"4C",X"32",X"4E",X"4C",X"CD",X"DA",X"05",
		X"C3",X"35",X"08",X"CD",X"75",X"00",X"CD",X"6D",X"00",X"C3",X"35",X"08",X"E5",X"3E",X"0B",X"32",
		X"45",X"4E",X"CD",X"75",X"00",X"CD",X"6D",X"00",X"3E",X"04",X"CD",X"04",X"01",X"E1",X"3E",X"60",
		X"32",X"21",X"4C",X"AF",X"32",X"26",X"4C",X"3A",X"26",X"4C",X"A7",X"28",X"FA",X"E5",X"CD",X"14",
		X"13",X"CD",X"75",X"00",X"E1",X"23",X"7E",X"FE",X"FF",X"CA",X"05",X"09",X"20",X"A3",X"23",X"7E",
		X"35",X"FE",X"00",X"28",X"2A",X"2B",X"7E",X"FE",X"FF",X"28",X"1B",X"CD",X"75",X"00",X"CD",X"6D",
		X"00",X"AF",X"32",X"03",X"50",X"3A",X"51",X"4C",X"32",X"4E",X"4C",X"3E",X"01",X"32",X"47",X"4C",
		X"CD",X"DA",X"05",X"C3",X"35",X"08",X"CD",X"75",X"00",X"CD",X"6D",X"00",X"C3",X"35",X"08",X"E5",
		X"3E",X"0B",X"32",X"45",X"4E",X"CD",X"75",X"00",X"CD",X"6D",X"00",X"3E",X"05",X"CD",X"04",X"01",
		X"E1",X"3E",X"60",X"32",X"21",X"4C",X"AF",X"32",X"26",X"4C",X"3A",X"26",X"4C",X"A7",X"28",X"FA",
		X"E5",X"CD",X"14",X"13",X"CD",X"75",X"00",X"E1",X"2B",X"7E",X"FE",X"FF",X"20",X"AD",X"CA",X"05",
		X"09",X"C3",X"C8",X"06",X"AF",X"32",X"50",X"4C",X"32",X"3F",X"4E",X"3E",X"46",X"32",X"50",X"4E",
		X"3E",X"01",X"32",X"4F",X"4E",X"3A",X"50",X"4E",X"A7",X"20",X"FA",X"AF",X"32",X"4F",X"4E",X"3E",
		X"01",X"32",X"4C",X"4C",X"32",X"66",X"4C",X"AF",X"32",X"4F",X"4C",X"CD",X"34",X"34",X"CD",X"6D",
		X"00",X"CD",X"75",X"00",X"3E",X"0E",X"CD",X"04",X"01",X"CD",X"4B",X"33",X"3E",X"0C",X"32",X"45",
		X"4E",X"3E",X"60",X"32",X"21",X"4C",X"AF",X"21",X"26",X"4C",X"77",X"7E",X"A7",X"28",X"FC",X"3E",
		X"0F",X"CD",X"04",X"01",X"3E",X"60",X"32",X"21",X"4C",X"AF",X"21",X"26",X"4C",X"77",X"7E",X"A7",
		X"28",X"FC",X"CD",X"75",X"00",X"21",X"4E",X"4C",X"7E",X"FE",X"14",X"28",X"10",X"34",X"21",X"51",
		X"4C",X"3A",X"47",X"4C",X"FE",X"01",X"28",X"01",X"23",X"3A",X"4E",X"4C",X"77",X"CF",X"CD",X"FB",
		X"31",X"C3",X"6F",X"08",X"CD",X"5C",X"00",X"CD",X"4A",X"00",X"CD",X"7F",X"00",X"CD",X"F2",X"03",
		X"CD",X"B1",X"04",X"CD",X"2E",X"04",X"CD",X"E5",X"04",X"CD",X"7F",X"05",X"CD",X"BA",X"05",X"AF",
		X"32",X"70",X"50",X"32",X"0A",X"4E",X"32",X"3F",X"4E",X"DD",X"21",X"02",X"4E",X"DD",X"36",X"00",
		X"88",X"DD",X"36",X"01",X"A0",X"DD",X"36",X"02",X"A8",X"DD",X"36",X"03",X"AC",X"DD",X"36",X"04",
		X"8A",X"DD",X"36",X"05",X"A2",X"DD",X"36",X"06",X"AB",X"DD",X"36",X"07",X"AD",X"16",X"01",X"21",
		X"00",X"44",X"01",X"00",X"04",X"72",X"23",X"0B",X"78",X"B1",X"20",X"F9",X"0E",X"07",X"06",X"03",
		X"C5",X"79",X"CD",X"04",X"01",X"C1",X"0C",X"10",X"F7",X"3A",X"6E",X"4E",X"FE",X"FF",X"28",X"05",
		X"3E",X"0A",X"CD",X"04",X"01",X"3E",X"3C",X"32",X"23",X"4C",X"AF",X"32",X"65",X"40",X"32",X"71",
		X"40",X"32",X"7E",X"40",X"3E",X"05",X"06",X"20",X"21",X"60",X"44",X"77",X"23",X"10",X"FC",X"3A",
		X"32",X"4C",X"FE",X"03",X"C9",X"F3",X"F5",X"AF",X"32",X"C0",X"50",X"32",X"00",X"50",X"C5",X"D5",
		X"E5",X"DD",X"E5",X"FD",X"E5",X"DD",X"21",X"00",X"4C",X"21",X"F0",X"4F",X"11",X"60",X"50",X"06",
		X"08",X"3A",X"47",X"4C",X"FE",X"01",X"28",X"28",X"3A",X"52",X"4E",X"A7",X"20",X"22",X"DD",X"7E",
		X"00",X"EE",X"03",X"77",X"23",X"DD",X"7E",X"01",X"77",X"DD",X"7E",X"10",X"C6",X"0F",X"12",X"13",
		X"DD",X"7E",X"11",X"C6",X"0F",X"12",X"13",X"23",X"DD",X"23",X"DD",X"23",X"10",X"DA",X"18",X"13",
		X"06",X"10",X"DD",X"7E",X"00",X"77",X"DD",X"7E",X"10",X"ED",X"44",X"3D",X"12",X"13",X"23",X"DD",
		X"23",X"10",X"EF",X"21",X"53",X"4C",X"34",X"CD",X"FD",X"03",X"CD",X"FD",X"04",X"CD",X"8F",X"00",
		X"EF",X"CD",X"05",X"13",X"3A",X"4F",X"4E",X"A7",X"C2",X"19",X"0D",X"21",X"19",X"0D",X"E5",X"3A",
		X"20",X"4C",X"87",X"16",X"00",X"5F",X"21",X"CF",X"0B",X"19",X"5E",X"23",X"56",X"EB",X"E9",X"D7",
		X"0B",X"D8",X"0B",X"9A",X"0C",X"F5",X"0C",X"C9",X"3A",X"41",X"4E",X"FE",X"FF",X"C0",X"AF",X"32",
		X"41",X"4E",X"21",X"F2",X"0B",X"3A",X"40",X"4E",X"87",X"5F",X"16",X"00",X"19",X"5E",X"23",X"56",
		X"EB",X"E9",X"FC",X"0B",X"10",X"0C",X"14",X"0C",X"57",X"0C",X"83",X"0C",X"3E",X"01",X"32",X"40",
		X"4E",X"AF",X"32",X"0B",X"4E",X"3E",X"01",X"32",X"0C",X"4E",X"3E",X"43",X"32",X"0D",X"4E",X"C9",
		X"CD",X"DC",X"0D",X"C9",X"E7",X"FE",X"FF",X"C0",X"3E",X"10",X"CD",X"04",X"01",X"3E",X"11",X"CD",
		X"04",X"01",X"3E",X"12",X"CD",X"04",X"01",X"3E",X"19",X"CD",X"04",X"01",X"3E",X"1A",X"CD",X"04",
		X"01",X"3E",X"1B",X"CD",X"04",X"01",X"3E",X"1C",X"CD",X"04",X"01",X"3E",X"03",X"32",X"40",X"4E",
		X"3E",X"09",X"32",X"45",X"4E",X"32",X"4D",X"4E",X"3E",X"02",X"32",X"7C",X"4E",X"3E",X"FF",X"32",
		X"7D",X"4E",X"AF",X"32",X"0E",X"4E",X"C9",X"CD",X"A9",X"0D",X"3A",X"20",X"4C",X"3D",X"C0",X"3A",
		X"53",X"4E",X"A7",X"C8",X"3A",X"7D",X"4E",X"A7",X"28",X"05",X"3D",X"32",X"7D",X"4E",X"C9",X"3A",
		X"7C",X"4E",X"A7",X"28",X"0A",X"3D",X"32",X"7C",X"4E",X"3E",X"FF",X"32",X"7D",X"4E",X"C9",X"32",
		X"4D",X"4E",X"C9",X"3A",X"3F",X"4E",X"FE",X"00",X"C2",X"2B",X"0D",X"CD",X"5E",X"10",X"D7",X"DF",
		X"CD",X"D3",X"32",X"CD",X"50",X"36",X"CD",X"57",X"37",X"C9",X"3A",X"6E",X"4E",X"FE",X"01",X"28",
		X"07",X"3E",X"01",X"CD",X"04",X"01",X"18",X"05",X"3E",X"00",X"CD",X"04",X"01",X"3A",X"30",X"4C",
		X"07",X"07",X"07",X"E6",X"03",X"C8",X"21",X"6E",X"4E",X"CB",X"47",X"20",X"17",X"7E",X"FE",X"02",
		X"D8",X"FE",X"FF",X"28",X"05",X"35",X"35",X"CD",X"56",X"05",X"3E",X"02",X"32",X"46",X"4C",X"CD",
		X"0F",X"16",X"18",X"0E",X"7E",X"FE",X"FF",X"28",X"04",X"35",X"CD",X"56",X"05",X"3E",X"01",X"32",
		X"46",X"4C",X"CD",X"03",X"16",X"3A",X"32",X"4C",X"FE",X"03",X"28",X"00",X"CD",X"75",X"00",X"3E",
		X"01",X"32",X"47",X"4C",X"C9",X"3A",X"3F",X"4E",X"FE",X"00",X"20",X"2F",X"3A",X"4C",X"4C",X"A7",
		X"C0",X"CD",X"D4",X"1A",X"3A",X"50",X"4C",X"A7",X"28",X"0B",X"DF",X"CD",X"D3",X"32",X"CD",X"50",
		X"36",X"CD",X"57",X"37",X"C9",X"D7",X"C3",X"0A",X"0D",X"FD",X"E1",X"DD",X"E1",X"E1",X"D1",X"C1",
		X"3E",X"01",X"32",X"00",X"50",X"32",X"C0",X"50",X"F1",X"FB",X"C9",X"CD",X"45",X"0D",X"3A",X"00",
		X"4E",X"FE",X"01",X"C0",X"3E",X"01",X"32",X"50",X"4C",X"3E",X"00",X"32",X"3F",X"4E",X"32",X"40",
		X"4E",X"32",X"01",X"50",X"C9",X"21",X"10",X"4C",X"CB",X"46",X"20",X"3A",X"3A",X"01",X"4E",X"A7",
		X"20",X"37",X"3A",X"10",X"4C",X"FE",X"2A",X"28",X"35",X"FE",X"28",X"28",X"41",X"21",X"10",X"4C",
		X"35",X"35",X"21",X"02",X"4E",X"16",X"00",X"3A",X"0A",X"4E",X"5F",X"19",X"7E",X"32",X"00",X"4C",
		X"3E",X"03",X"32",X"01",X"4E",X"3A",X"0A",X"4E",X"FE",X"07",X"28",X"05",X"3C",X"32",X"0A",X"4E",
		X"C9",X"AF",X"32",X"0A",X"4E",X"C9",X"CB",X"86",X"C9",X"21",X"01",X"4E",X"35",X"C9",X"21",X"10",
		X"4C",X"35",X"35",X"3E",X"8A",X"32",X"00",X"4C",X"3E",X"03",X"32",X"01",X"4E",X"C9",X"3E",X"01",
		X"32",X"00",X"4E",X"3E",X"8A",X"32",X"00",X"4C",X"C9",X"3A",X"0E",X"4E",X"A7",X"20",X"1C",X"21",
		X"00",X"4C",X"06",X"08",X"7E",X"FE",X"98",X"20",X"0D",X"3E",X"99",X"77",X"23",X"23",X"10",X"FB",
		X"3E",X"20",X"32",X"0E",X"4E",X"C9",X"3E",X"98",X"C3",X"BB",X"0D",X"21",X"0E",X"4E",X"35",X"C9",
		X"21",X"01",X"4C",X"AF",X"06",X"08",X"77",X"23",X"23",X"10",X"FB",X"C9",X"3A",X"0D",X"4E",X"FE",
		X"00",X"20",X"10",X"3A",X"0C",X"4E",X"FE",X"00",X"28",X"0E",X"21",X"0D",X"4E",X"35",X"21",X"0C",
		X"4E",X"35",X"C9",X"21",X"0D",X"4E",X"35",X"C9",X"3E",X"FF",X"32",X"0B",X"4E",X"C9",X"DD",X"21",
		X"0E",X"4E",X"DD",X"36",X"00",X"00",X"3E",X"FF",X"DD",X"77",X"06",X"DD",X"77",X"0C",X"DD",X"77",
		X"12",X"DD",X"77",X"18",X"DD",X"77",X"1E",X"DD",X"77",X"24",X"DD",X"77",X"2A",X"3E",X"80",X"DD",
		X"77",X"01",X"DD",X"77",X"07",X"DD",X"77",X"0D",X"DD",X"77",X"13",X"DD",X"77",X"19",X"DD",X"77",
		X"1F",X"DD",X"77",X"25",X"DD",X"77",X"2B",X"3E",X"14",X"DD",X"77",X"02",X"DD",X"77",X"08",X"DD",
		X"77",X"0E",X"DD",X"77",X"14",X"DD",X"77",X"1A",X"DD",X"77",X"20",X"DD",X"77",X"26",X"DD",X"77",
		X"2C",X"3E",X"58",X"DD",X"77",X"03",X"DD",X"77",X"09",X"DD",X"77",X"0F",X"DD",X"77",X"15",X"DD",
		X"77",X"1B",X"DD",X"77",X"21",X"DD",X"77",X"27",X"DD",X"77",X"2D",X"3E",X"EE",X"DD",X"77",X"04",
		X"DD",X"77",X"0A",X"DD",X"77",X"10",X"DD",X"77",X"16",X"DD",X"77",X"1C",X"DD",X"77",X"22",X"DD",
		X"77",X"28",X"DD",X"77",X"2E",X"DD",X"36",X"05",X"20",X"DD",X"36",X"0B",X"38",X"DD",X"36",X"11",
		X"50",X"DD",X"36",X"17",X"68",X"DD",X"36",X"1D",X"88",X"DD",X"36",X"23",X"A0",X"DD",X"36",X"29",
		X"B8",X"DD",X"36",X"2F",X"D0",X"C9",X"CD",X"AD",X"0F",X"DD",X"21",X"0E",X"4E",X"DD",X"7E",X"00",
		X"FE",X"FF",X"28",X"3F",X"DD",X"7E",X"01",X"FE",X"98",X"CA",X"7B",X"0F",X"DD",X"7E",X"04",X"FE",
		X"E0",X"CA",X"74",X"0F",X"FE",X"D0",X"CA",X"6D",X"0F",X"FE",X"C0",X"CA",X"66",X"0F",X"FE",X"B0",
		X"CA",X"5F",X"0F",X"FE",X"A0",X"CA",X"58",X"0F",X"FE",X"90",X"28",X"75",X"FE",X"80",X"CA",X"43",
		X"0F",X"FE",X"20",X"28",X"65",X"DD",X"35",X"04",X"DD",X"7E",X"01",X"FE",X"80",X"28",X"4D",X"DD",
		X"36",X"01",X"80",X"DD",X"21",X"14",X"4E",X"CD",X"1C",X"00",X"DD",X"21",X"1A",X"4E",X"CD",X"1C",
		X"00",X"DD",X"21",X"20",X"4E",X"CD",X"1C",X"00",X"DD",X"21",X"26",X"4E",X"CD",X"1C",X"00",X"DD",
		X"21",X"2C",X"4E",X"CD",X"1C",X"00",X"DD",X"21",X"32",X"4E",X"CD",X"1C",X"00",X"DD",X"21",X"38",
		X"4E",X"CD",X"1C",X"00",X"3A",X"0E",X"4E",X"FE",X"FF",X"20",X"0F",X"3A",X"38",X"4E",X"FE",X"FF",
		X"20",X"08",X"3E",X"98",X"32",X"0E",X"4C",X"3E",X"FF",X"C9",X"AF",X"C9",X"DD",X"36",X"01",X"84",
		X"C3",X"F3",X"0E",X"AF",X"32",X"38",X"4E",X"C3",X"E5",X"0E",X"DD",X"36",X"01",X"98",X"C3",X"F3",
		X"0E",X"AF",X"32",X"32",X"4E",X"C3",X"E5",X"0E",X"AF",X"32",X"2C",X"4E",X"C3",X"E5",X"0E",X"AF",
		X"32",X"26",X"4E",X"C3",X"E5",X"0E",X"AF",X"32",X"20",X"4E",X"C3",X"E5",X"0E",X"AF",X"32",X"1A",
		X"4E",X"C3",X"E5",X"0E",X"AF",X"32",X"14",X"4E",X"C3",X"E5",X"0E",X"DD",X"36",X"00",X"FF",X"C3",
		X"F3",X"0E",X"DD",X"7E",X"00",X"FE",X"FF",X"C8",X"DD",X"7E",X"04",X"DD",X"BE",X"05",X"28",X"14",
		X"DD",X"35",X"04",X"DD",X"7E",X"01",X"FE",X"80",X"20",X"05",X"DD",X"36",X"01",X"84",X"C9",X"DD",
		X"36",X"01",X"80",X"C9",X"DD",X"36",X"01",X"98",X"DD",X"36",X"00",X"FF",X"C9",X"21",X"0F",X"4E",
		X"11",X"00",X"4C",X"01",X"02",X"00",X"ED",X"B0",X"21",X"11",X"4E",X"11",X"10",X"4C",X"01",X"02",
		X"00",X"ED",X"B0",X"21",X"15",X"4E",X"11",X"02",X"4C",X"01",X"02",X"00",X"ED",X"B0",X"21",X"17",
		X"4E",X"11",X"12",X"4C",X"01",X"02",X"00",X"ED",X"B0",X"21",X"1B",X"4E",X"11",X"04",X"4C",X"01",
		X"02",X"00",X"ED",X"B0",X"21",X"1D",X"4E",X"11",X"14",X"4C",X"01",X"02",X"00",X"ED",X"B0",X"21",
		X"21",X"4E",X"11",X"06",X"4C",X"01",X"02",X"00",X"ED",X"B0",X"21",X"23",X"4E",X"11",X"16",X"4C",
		X"01",X"02",X"00",X"ED",X"B0",X"21",X"27",X"4E",X"11",X"08",X"4C",X"01",X"02",X"00",X"ED",X"B0",
		X"21",X"29",X"4E",X"11",X"18",X"4C",X"01",X"02",X"00",X"ED",X"B0",X"21",X"2D",X"4E",X"11",X"0A",
		X"4C",X"01",X"02",X"00",X"ED",X"B0",X"21",X"2F",X"4E",X"11",X"1A",X"4C",X"01",X"02",X"00",X"ED",
		X"B0",X"21",X"33",X"4E",X"11",X"0C",X"4C",X"01",X"02",X"00",X"ED",X"B0",X"21",X"35",X"4E",X"11",
		X"1C",X"4C",X"01",X"02",X"00",X"ED",X"B0",X"21",X"39",X"4E",X"11",X"0E",X"4C",X"01",X"02",X"00",
		X"ED",X"B0",X"21",X"3B",X"4E",X"11",X"1E",X"4C",X"01",X"02",X"00",X"ED",X"B0",X"C9",X"21",X"6F",
		X"10",X"3A",X"3E",X"4E",X"87",X"5F",X"16",X"00",X"19",X"5E",X"23",X"56",X"EB",X"E9",X"35",X"97",
		X"10",X"AE",X"10",X"F0",X"10",X"0D",X"11",X"2A",X"11",X"47",X"11",X"64",X"11",X"81",X"11",X"9E",
		X"11",X"BB",X"11",X"D9",X"11",X"F1",X"11",X"09",X"12",X"20",X"12",X"3E",X"12",X"56",X"12",X"6D",
		X"12",X"B0",X"12",X"C8",X"12",X"E0",X"12",X"3A",X"11",X"4C",X"FE",X"94",X"28",X"06",X"3E",X"02",
		X"32",X"60",X"4C",X"C9",X"AF",X"32",X"60",X"4C",X"3E",X"01",X"32",X"3E",X"4E",X"C9",X"3A",X"60",
		X"4C",X"A7",X"28",X"17",X"3A",X"10",X"4C",X"FE",X"48",X"28",X"06",X"3E",X"01",X"32",X"60",X"4C",
		X"C9",X"AF",X"32",X"60",X"4C",X"3E",X"02",X"32",X"3E",X"4E",X"C9",X"3A",X"1D",X"4C",X"47",X"3A",
		X"CD",X"4C",X"A7",X"28",X"10",X"3E",X"88",X"B8",X"38",X"06",X"3E",X"01",X"32",X"60",X"4C",X"C9",
		X"AF",X"32",X"60",X"4C",X"C9",X"3E",X"20",X"B8",X"38",X"F6",X"3E",X"01",X"32",X"60",X"4C",X"C9",
		X"3A",X"60",X"4C",X"A7",X"28",X"07",X"3A",X"11",X"4C",X"FE",X"B0",X"28",X"06",X"3E",X"04",X"32",
		X"60",X"4C",X"C9",X"AF",X"32",X"60",X"4C",X"3E",X"03",X"32",X"3E",X"4E",X"C9",X"3A",X"60",X"4C",
		X"A7",X"28",X"07",X"3A",X"10",X"4C",X"FE",X"48",X"28",X"06",X"3E",X"10",X"32",X"60",X"4C",X"C9",
		X"AF",X"32",X"60",X"4C",X"3E",X"04",X"32",X"3E",X"4E",X"C9",X"3A",X"60",X"4C",X"A7",X"28",X"07",
		X"3A",X"11",X"4C",X"FE",X"C8",X"28",X"06",X"3E",X"04",X"32",X"60",X"4C",X"C9",X"AF",X"32",X"60",
		X"4C",X"3E",X"05",X"32",X"3E",X"4E",X"C9",X"3A",X"60",X"4C",X"A7",X"28",X"07",X"3A",X"10",X"4C",
		X"FE",X"68",X"28",X"06",X"3E",X"01",X"32",X"60",X"4C",X"C9",X"AF",X"32",X"60",X"4C",X"3E",X"06",
		X"32",X"3E",X"4E",X"C9",X"3A",X"60",X"4C",X"A7",X"28",X"07",X"3A",X"11",X"4C",X"FE",X"C4",X"28",
		X"06",X"3E",X"02",X"32",X"60",X"4C",X"C9",X"AF",X"32",X"60",X"4C",X"3E",X"07",X"32",X"3E",X"4E",
		X"C9",X"3A",X"60",X"4C",X"A7",X"28",X"07",X"3A",X"10",X"4C",X"FE",X"68",X"28",X"06",X"3E",X"10",
		X"32",X"60",X"4C",X"C9",X"AF",X"32",X"60",X"4C",X"3E",X"08",X"32",X"3E",X"4E",X"C9",X"3A",X"60",
		X"4C",X"A7",X"28",X"07",X"3A",X"11",X"4C",X"FE",X"A0",X"28",X"06",X"3E",X"02",X"32",X"60",X"4C",
		X"C9",X"AF",X"32",X"60",X"4C",X"3E",X"09",X"32",X"3E",X"4E",X"C9",X"3A",X"60",X"4C",X"A7",X"28",
		X"07",X"3A",X"10",X"4C",X"FE",X"68",X"28",X"06",X"3E",X"12",X"32",X"60",X"4C",X"C9",X"3E",X"02",
		X"32",X"60",X"4C",X"3E",X"0A",X"32",X"3E",X"4E",X"C9",X"3A",X"11",X"4C",X"FE",X"64",X"28",X"06",
		X"3E",X"02",X"32",X"60",X"4C",X"C9",X"3E",X"01",X"32",X"60",X"4C",X"3E",X"0B",X"32",X"3E",X"4E",
		X"C9",X"3A",X"10",X"4C",X"FE",X"88",X"28",X"06",X"3E",X"01",X"32",X"60",X"4C",X"C9",X"3E",X"02",
		X"32",X"60",X"4C",X"3E",X"0C",X"32",X"3E",X"4E",X"C9",X"3A",X"11",X"4C",X"FE",X"44",X"28",X"06",
		X"3E",X"02",X"32",X"60",X"4C",X"C9",X"AF",X"32",X"60",X"4C",X"3E",X"0D",X"32",X"3E",X"4E",X"C9",
		X"3A",X"60",X"4C",X"A7",X"28",X"07",X"3A",X"10",X"4C",X"FE",X"88",X"28",X"06",X"3E",X"12",X"32",
		X"60",X"4C",X"C9",X"3E",X"02",X"32",X"60",X"4C",X"3E",X"0E",X"32",X"3E",X"4E",X"C9",X"3A",X"11",
		X"4C",X"FE",X"02",X"28",X"06",X"3E",X"02",X"32",X"60",X"4C",X"C9",X"3E",X"04",X"32",X"60",X"4C",
		X"3E",X"0F",X"32",X"3E",X"4E",X"C9",X"3A",X"11",X"4C",X"FE",X"18",X"28",X"06",X"3E",X"04",X"32",
		X"60",X"4C",X"C9",X"AF",X"32",X"60",X"4C",X"3E",X"10",X"32",X"3E",X"4E",X"C9",X"3A",X"60",X"4C",
		X"FE",X"00",X"28",X"18",X"3A",X"10",X"4C",X"FE",X"A8",X"28",X"06",X"3E",X"01",X"32",X"60",X"4C",
		X"C9",X"3E",X"02",X"32",X"60",X"4C",X"3E",X"11",X"32",X"3E",X"4E",X"C9",X"3A",X"1B",X"4C",X"47",
		X"3A",X"C6",X"4C",X"A7",X"20",X"10",X"3E",X"30",X"B8",X"38",X"05",X"AF",X"32",X"60",X"4C",X"C9",
		X"3E",X"01",X"32",X"60",X"4C",X"C9",X"3E",X"B0",X"B8",X"38",X"F5",X"AF",X"32",X"60",X"4C",X"C9",
		X"3A",X"11",X"4C",X"FE",X"02",X"28",X"06",X"3E",X"02",X"32",X"60",X"4C",X"C9",X"3E",X"04",X"32",
		X"60",X"4C",X"3E",X"12",X"32",X"3E",X"4E",X"C9",X"3A",X"11",X"4C",X"FE",X"18",X"28",X"06",X"3E",
		X"04",X"32",X"60",X"4C",X"C9",X"3E",X"08",X"32",X"60",X"4C",X"3E",X"13",X"32",X"3E",X"4E",X"C9",
		X"3A",X"10",X"4C",X"FE",X"88",X"28",X"06",X"3E",X"08",X"32",X"60",X"4C",X"C9",X"3E",X"04",X"32",
		X"60",X"4C",X"C9",X"DD",X"21",X"A5",X"4C",X"11",X"08",X"00",X"06",X"04",X"AF",X"DD",X"77",X"00",
		X"DD",X"19",X"10",X"F9",X"C9",X"3A",X"4F",X"4E",X"A7",X"C8",X"3A",X"50",X"4E",X"A7",X"C8",X"3D",
		X"32",X"50",X"4E",X"C9",X"F5",X"AF",X"32",X"00",X"50",X"C5",X"D5",X"E5",X"DD",X"E5",X"FD",X"E5",
		X"CD",X"75",X"00",X"3E",X"0F",X"32",X"5D",X"4E",X"32",X"61",X"4E",X"32",X"65",X"4E",X"32",X"69",
		X"4E",X"32",X"6D",X"4E",X"3E",X"17",X"CD",X"04",X"01",X"3E",X"18",X"CD",X"04",X"01",X"CD",X"66",
		X"14",X"11",X"4A",X"41",X"3A",X"5D",X"4E",X"4F",X"21",X"E9",X"15",X"CD",X"CE",X"15",X"11",X"8A",
		X"41",X"21",X"EC",X"15",X"3A",X"61",X"4E",X"4F",X"CD",X"CE",X"15",X"11",X"CA",X"41",X"21",X"EF",
		X"15",X"3A",X"65",X"4E",X"4F",X"CD",X"CE",X"15",X"11",X"0A",X"42",X"21",X"F2",X"15",X"3A",X"69",
		X"4E",X"4F",X"CD",X"CE",X"15",X"11",X"4A",X"42",X"21",X"F5",X"15",X"3A",X"6D",X"4E",X"4F",X"CD",
		X"CE",X"15",X"11",X"53",X"41",X"21",X"5A",X"4E",X"3A",X"5D",X"4E",X"4F",X"CD",X"AA",X"15",X"11",
		X"93",X"41",X"21",X"5E",X"4E",X"3A",X"61",X"4E",X"4F",X"CD",X"AA",X"15",X"11",X"D3",X"41",X"21",
		X"62",X"4E",X"3A",X"65",X"4E",X"4F",X"CD",X"AA",X"15",X"11",X"13",X"42",X"21",X"66",X"4E",X"3A",
		X"69",X"4E",X"4F",X"CD",X"AA",X"15",X"11",X"53",X"42",X"21",X"6A",X"4E",X"3A",X"6D",X"4E",X"4F",
		X"CD",X"AA",X"15",X"3E",X"06",X"32",X"22",X"4C",X"3E",X"1F",X"32",X"21",X"4C",X"AF",X"32",X"27",
		X"4C",X"32",X"26",X"4C",X"3C",X"32",X"00",X"50",X"3A",X"26",X"4C",X"A7",X"20",X"0F",X"3A",X"27",
		X"4C",X"A7",X"28",X"F4",X"FD",X"E1",X"DD",X"E1",X"E1",X"D1",X"C1",X"F1",X"C9",X"3E",X"1F",X"32",
		X"21",X"4C",X"AF",X"32",X"26",X"4C",X"3E",X"18",X"21",X"5D",X"4E",X"BE",X"28",X"1B",X"21",X"61",
		X"4E",X"BE",X"28",X"19",X"21",X"65",X"4E",X"BE",X"28",X"18",X"21",X"69",X"4E",X"BE",X"28",X"17",
		X"21",X"6D",X"4E",X"BE",X"28",X"16",X"C3",X"DE",X"13",X"AF",X"C3",X"31",X"14",X"3E",X"01",X"C3",
		X"31",X"14",X"3E",X"02",X"C3",X"31",X"14",X"3E",X"03",X"C3",X"31",X"14",X"3E",X"04",X"C3",X"31",
		X"14",X"87",X"21",X"5C",X"14",X"16",X"00",X"5F",X"19",X"5E",X"23",X"56",X"DD",X"21",X"00",X"04",
		X"DD",X"19",X"DD",X"7E",X"00",X"FE",X"18",X"20",X"0E",X"3E",X"0F",X"06",X"0F",X"DD",X"77",X"00",
		X"DD",X"23",X"10",X"F9",X"C3",X"DE",X"13",X"3E",X"18",X"C3",X"4B",X"14",X"4A",X"41",X"8A",X"41",
		X"CA",X"41",X"0A",X"42",X"4A",X"42",X"3A",X"47",X"4C",X"3D",X"20",X"39",X"21",X"3A",X"4C",X"E5",
		X"11",X"5A",X"4E",X"CD",X"F8",X"15",X"38",X"33",X"E1",X"E5",X"11",X"5E",X"4E",X"CD",X"F8",X"15",
		X"38",X"72",X"E1",X"E5",X"11",X"62",X"4E",X"CD",X"F8",X"15",X"DA",X"32",X"15",X"E1",X"E5",X"11",
		X"66",X"4E",X"CD",X"F8",X"15",X"DA",X"65",X"15",X"E1",X"E5",X"11",X"6A",X"4E",X"CD",X"F8",X"15",
		X"DA",X"8D",X"15",X"E1",X"C9",X"21",X"3D",X"4C",X"C3",X"6F",X"14",X"21",X"5D",X"4E",X"36",X"18",
		X"3E",X"0F",X"32",X"61",X"4E",X"32",X"65",X"4E",X"32",X"69",X"4E",X"32",X"6D",X"4E",X"21",X"66",
		X"4E",X"11",X"6A",X"4E",X"01",X"03",X"00",X"ED",X"B0",X"21",X"62",X"4E",X"11",X"66",X"4E",X"01",
		X"03",X"00",X"ED",X"B0",X"21",X"5E",X"4E",X"11",X"62",X"4E",X"01",X"03",X"00",X"ED",X"B0",X"21",
		X"5A",X"4E",X"11",X"5E",X"4E",X"01",X"03",X"00",X"ED",X"B0",X"E1",X"11",X"5A",X"4E",X"01",X"03",
		X"00",X"ED",X"B0",X"C9",X"21",X"61",X"4E",X"36",X"18",X"3E",X"0F",X"32",X"5D",X"4E",X"32",X"65",
		X"4E",X"32",X"69",X"4E",X"32",X"6D",X"4E",X"21",X"66",X"4E",X"11",X"6A",X"4E",X"01",X"03",X"00",
		X"ED",X"B0",X"21",X"62",X"4E",X"11",X"66",X"4E",X"01",X"03",X"00",X"ED",X"B0",X"21",X"5E",X"4E",
		X"11",X"62",X"4E",X"01",X"03",X"00",X"ED",X"B0",X"E1",X"11",X"5E",X"4E",X"01",X"03",X"00",X"ED",
		X"B0",X"C9",X"21",X"65",X"4E",X"36",X"18",X"3E",X"0F",X"32",X"5D",X"4E",X"32",X"61",X"4E",X"32",
		X"69",X"4E",X"32",X"6D",X"4E",X"21",X"66",X"4E",X"11",X"6A",X"4E",X"01",X"03",X"00",X"ED",X"B0",
		X"21",X"62",X"4E",X"11",X"66",X"4E",X"01",X"03",X"00",X"ED",X"B0",X"E1",X"11",X"62",X"4E",X"01",
		X"03",X"00",X"ED",X"B0",X"C9",X"21",X"69",X"4E",X"36",X"18",X"3E",X"0F",X"32",X"5D",X"4E",X"32",
		X"61",X"4E",X"32",X"65",X"4E",X"32",X"6D",X"4E",X"21",X"66",X"4E",X"11",X"6A",X"4E",X"01",X"03",
		X"00",X"ED",X"B0",X"E1",X"11",X"66",X"4E",X"01",X"03",X"00",X"ED",X"B0",X"C9",X"21",X"6D",X"4E",
		X"36",X"18",X"3E",X"0F",X"32",X"5D",X"4E",X"32",X"61",X"4E",X"32",X"65",X"4E",X"32",X"69",X"4E",
		X"E1",X"11",X"6A",X"4E",X"01",X"03",X"00",X"ED",X"B0",X"C9",X"DD",X"21",X"00",X"04",X"DD",X"19",
		X"06",X"03",X"7E",X"E6",X"F0",X"0F",X"0F",X"0F",X"0F",X"12",X"DD",X"71",X"00",X"13",X"DD",X"23",
		X"7E",X"E6",X"0F",X"12",X"DD",X"71",X"00",X"13",X"DD",X"23",X"23",X"10",X"E5",X"C9",X"06",X"03",
		X"DD",X"21",X"00",X"04",X"DD",X"19",X"7E",X"D6",X"30",X"FE",X"0A",X"38",X"01",X"3D",X"12",X"DD",
		X"71",X"00",X"23",X"13",X"DD",X"23",X"10",X"EE",X"C9",X"54",X"4F",X"50",X"32",X"4E",X"44",X"33",
		X"52",X"44",X"34",X"54",X"48",X"35",X"54",X"48",X"06",X"03",X"1A",X"96",X"C0",X"23",X"13",X"10",
		X"F9",X"A7",X"C9",X"3A",X"31",X"4C",X"A7",X"20",X"05",X"3E",X"01",X"32",X"4A",X"4C",X"C9",X"3A",
		X"31",X"4C",X"A7",X"20",X"05",X"3E",X"01",X"32",X"4B",X"4C",X"C9",X"21",X"60",X"4C",X"CB",X"66",
		X"20",X"04",X"AF",X"32",X"5E",X"4C",X"3A",X"5E",X"4C",X"A7",X"20",X"06",X"CB",X"66",X"C4",X"0C",
		X"00",X"D8",X"3A",X"58",X"4C",X"A7",X"C2",X"13",X"18",X"3A",X"57",X"4C",X"A7",X"C2",X"36",X"17",
		X"7E",X"FE",X"00",X"CA",X"95",X"16",X"CB",X"47",X"C2",X"02",X"17",X"CB",X"5F",X"C2",X"1B",X"17",
		X"CB",X"4F",X"20",X"6A",X"CB",X"57",X"C8",X"21",X"56",X"4C",X"7E",X"FE",X"02",X"20",X"49",X"3A",
		X"5A",X"4C",X"FE",X"01",X"20",X"0D",X"3A",X"11",X"4C",X"FE",X"ED",X"CA",X"95",X"16",X"D2",X"95",
		X"16",X"18",X"07",X"3A",X"11",X"4C",X"FE",X"CD",X"C8",X"D0",X"CB",X"4F",X"28",X"04",X"3E",X"88",
		X"18",X"02",X"3E",X"8C",X"32",X"00",X"4C",X"3A",X"11",X"4C",X"C6",X"01",X"32",X"11",X"4C",X"3E",
		X"08",X"32",X"45",X"4E",X"C9",X"3A",X"46",X"4E",X"FE",X"07",X"C0",X"AF",X"32",X"01",X"50",X"32",
		X"45",X"4E",X"3E",X"0C",X"32",X"46",X"4E",X"C9",X"3A",X"11",X"4C",X"CB",X"4F",X"28",X"04",X"3E",
		X"88",X"18",X"02",X"3E",X"8C",X"32",X"00",X"4C",X"3E",X"02",X"32",X"56",X"4C",X"C9",X"21",X"56",
		X"4C",X"7E",X"FE",X"01",X"20",X"26",X"3A",X"11",X"4C",X"FE",X"02",X"CA",X"95",X"16",X"DA",X"95",
		X"16",X"CB",X"4F",X"28",X"04",X"3E",X"80",X"18",X"02",X"3E",X"84",X"32",X"00",X"4C",X"3A",X"11",
		X"4C",X"D6",X"01",X"32",X"11",X"4C",X"3E",X"08",X"32",X"45",X"4E",X"C9",X"3A",X"11",X"4C",X"CB",
		X"4F",X"28",X"04",X"3E",X"80",X"18",X"02",X"3E",X"84",X"32",X"00",X"4C",X"3E",X"01",X"32",X"56",
		X"4C",X"C9",X"CD",X"2C",X"00",X"D2",X"95",X"16",X"AF",X"32",X"59",X"4C",X"3C",X"32",X"57",X"4C",
		X"3E",X"90",X"32",X"00",X"4C",X"3E",X"08",X"32",X"45",X"4E",X"C9",X"CD",X"34",X"00",X"D2",X"95",
		X"16",X"3E",X"20",X"32",X"59",X"4C",X"3E",X"01",X"32",X"57",X"4C",X"3E",X"90",X"32",X"00",X"4C",
		X"3E",X"08",X"32",X"45",X"4E",X"C9",X"CB",X"46",X"20",X"05",X"CB",X"5E",X"20",X"44",X"C9",X"3A",
		X"59",X"4C",X"3C",X"32",X"59",X"4C",X"21",X"10",X"4C",X"34",X"FE",X"20",X"30",X"12",X"CB",X"4E",
		X"28",X"07",X"21",X"00",X"4C",X"3E",X"90",X"77",X"C9",X"21",X"00",X"4C",X"3E",X"94",X"77",X"C9",
		X"7E",X"E6",X"F8",X"77",X"3E",X"98",X"32",X"00",X"4C",X"21",X"10",X"4C",X"7E",X"CB",X"3F",X"CB",
		X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"32",X"5A",X"4C",X"AF",X"32",X"57",X"4C",X"32",X"56",
		X"4C",X"C9",X"3A",X"59",X"4C",X"3D",X"32",X"59",X"4C",X"21",X"10",X"4C",X"35",X"FE",X"01",X"FA",
		X"A4",X"17",X"CB",X"4E",X"28",X"07",X"21",X"00",X"4C",X"3E",X"90",X"77",X"C9",X"21",X"00",X"4C",
		X"3E",X"94",X"77",X"C9",X"7E",X"3C",X"E6",X"F8",X"77",X"3E",X"98",X"32",X"00",X"4C",X"21",X"10",
		X"4C",X"7E",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"32",X"5A",X"4C",X"AF",
		X"32",X"57",X"4C",X"32",X"56",X"4C",X"C9",X"3A",X"57",X"4C",X"A7",X"C0",X"3A",X"58",X"4C",X"A7",
		X"C0",X"3E",X"01",X"32",X"5E",X"4C",X"32",X"58",X"4C",X"3E",X"07",X"32",X"45",X"4E",X"AF",X"32",
		X"5B",X"4C",X"3A",X"60",X"4C",X"CB",X"4F",X"20",X"13",X"CB",X"57",X"20",X"1E",X"3A",X"56",X"4C",
		X"A7",X"28",X"0E",X"CB",X"4F",X"20",X"0F",X"21",X"E9",X"18",X"18",X"12",X"21",X"4B",X"19",X"18",
		X"0D",X"21",X"A7",X"18",X"18",X"08",X"21",X"C8",X"18",X"18",X"03",X"21",X"0A",X"19",X"22",X"5C",
		X"4C",X"37",X"C9",X"21",X"5B",X"4C",X"7E",X"FE",X"00",X"28",X"02",X"35",X"C9",X"3A",X"5F",X"4C",
		X"A7",X"20",X"59",X"2A",X"5C",X"4C",X"7E",X"FE",X"10",X"28",X"46",X"3A",X"11",X"4C",X"FE",X"02",
		X"28",X"44",X"38",X"42",X"3A",X"5A",X"4C",X"FE",X"01",X"20",X"0B",X"3A",X"11",X"4C",X"FE",X"ED",
		X"28",X"34",X"30",X"32",X"18",X"09",X"3A",X"11",X"4C",X"FE",X"CD",X"28",X"29",X"30",X"27",X"DD",
		X"21",X"00",X"4C",X"7E",X"DD",X"86",X"10",X"DD",X"77",X"10",X"23",X"7E",X"DD",X"86",X"11",X"DD",
		X"77",X"11",X"23",X"7E",X"DD",X"77",X"00",X"23",X"7E",X"32",X"5B",X"4C",X"23",X"22",X"5C",X"4C",
		X"C9",X"AF",X"32",X"58",X"4C",X"C9",X"3E",X"01",X"32",X"5F",X"4C",X"C9",X"2A",X"5C",X"4C",X"7E",
		X"FE",X"10",X"28",X"1B",X"DD",X"21",X"00",X"4C",X"7E",X"DD",X"86",X"10",X"DD",X"77",X"10",X"23",
		X"23",X"7E",X"DD",X"77",X"00",X"23",X"7E",X"32",X"5B",X"4C",X"23",X"22",X"5C",X"4C",X"C9",X"AF",
		X"32",X"58",X"4C",X"32",X"5F",X"4C",X"C9",X"03",X"00",X"98",X"02",X"02",X"00",X"98",X"02",X"02",
		X"00",X"99",X"02",X"01",X"00",X"99",X"02",X"FF",X"00",X"98",X"02",X"FE",X"00",X"98",X"02",X"FE",
		X"00",X"99",X"02",X"FD",X"00",X"99",X"02",X"10",X"02",X"03",X"A1",X"02",X"02",X"02",X"A5",X"02",
		X"01",X"02",X"A9",X"02",X"01",X"02",X"A9",X"02",X"FF",X"02",X"A9",X"02",X"FF",X"02",X"AD",X"02",
		X"FE",X"02",X"B1",X"02",X"FE",X"03",X"B5",X"02",X"10",X"02",X"FD",X"A0",X"02",X"02",X"FE",X"A4",
		X"02",X"01",X"FE",X"A8",X"02",X"01",X"FE",X"A8",X"02",X"FF",X"FE",X"A8",X"02",X"FF",X"FE",X"AC",
		X"02",X"FE",X"FE",X"B0",X"02",X"FE",X"FD",X"B4",X"02",X"10",X"02",X"03",X"A1",X"02",X"02",X"03",
		X"A1",X"02",X"02",X"03",X"A5",X"02",X"01",X"02",X"A5",X"02",X"01",X"02",X"A9",X"02",X"01",X"01",
		X"A9",X"02",X"01",X"01",X"A9",X"02",X"00",X"01",X"A9",X"02",X"00",X"01",X"A9",X"02",X"FF",X"01",
		X"A9",X"02",X"FF",X"01",X"AD",X"02",X"FF",X"02",X"AD",X"02",X"FF",X"02",X"B1",X"02",X"FE",X"03",
		X"B1",X"02",X"FE",X"03",X"B5",X"02",X"FE",X"03",X"B5",X"02",X"10",X"02",X"FD",X"A0",X"02",X"02",
		X"FD",X"A0",X"02",X"02",X"FE",X"A4",X"02",X"01",X"FE",X"A4",X"02",X"01",X"FE",X"A8",X"02",X"01",
		X"FF",X"A8",X"02",X"01",X"FF",X"A8",X"02",X"00",X"FF",X"A8",X"02",X"00",X"FF",X"A8",X"02",X"FF",
		X"FF",X"A8",X"02",X"FF",X"FF",X"AC",X"02",X"FF",X"FE",X"AC",X"02",X"FF",X"FE",X"B0",X"02",X"FE",
		X"FE",X"B0",X"02",X"FE",X"FD",X"B4",X"02",X"FE",X"FD",X"B4",X"02",X"10",X"3A",X"5A",X"4C",X"FE",
		X"05",X"28",X"2C",X"21",X"07",X"1B",X"3A",X"4E",X"4C",X"3D",X"87",X"5F",X"16",X"00",X"19",X"5E",
		X"23",X"56",X"EB",X"3A",X"5A",X"4C",X"3D",X"87",X"5F",X"16",X"00",X"19",X"5E",X"23",X"56",X"EB",
		X"3A",X"11",X"4C",X"47",X"7E",X"23",X"FE",X"00",X"28",X"05",X"B8",X"20",X"F7",X"37",X"C9",X"37",
		X"3F",X"C9",X"3A",X"5A",X"4C",X"FE",X"01",X"28",X"F6",X"21",X"07",X"1B",X"3A",X"4E",X"4C",X"3D",
		X"87",X"5F",X"16",X"00",X"19",X"5E",X"23",X"56",X"EB",X"3A",X"5A",X"4C",X"3D",X"18",X"C7",X"CD",
		X"14",X"00",X"3A",X"3F",X"4E",X"FE",X"04",X"C8",X"3A",X"58",X"4C",X"A7",X"C0",X"3A",X"4E",X"4C",
		X"3D",X"87",X"16",X"00",X"5F",X"21",X"5B",X"1F",X"19",X"5E",X"23",X"56",X"EB",X"3A",X"5A",X"4C",
		X"A7",X"C8",X"3D",X"87",X"16",X"00",X"5F",X"19",X"5E",X"23",X"56",X"EB",X"3A",X"11",X"4C",X"47",
		X"7E",X"A7",X"C8",X"D6",X"08",X"B8",X"28",X"03",X"23",X"18",X"F5",X"3E",X"04",X"32",X"3F",X"4E",
		X"AF",X"32",X"00",X"4E",X"32",X"0A",X"4E",X"3E",X"04",X"32",X"45",X"4E",X"C9",X"DD",X"21",X"A5",
		X"4C",X"FD",X"21",X"00",X"4C",X"06",X"04",X"DD",X"7E",X"00",X"A7",X"28",X"3F",X"DD",X"7E",X"04",
		X"A7",X"20",X"39",X"DD",X"6E",X"05",X"DD",X"66",X"06",X"11",X"10",X"00",X"19",X"7E",X"4F",X"FD",
		X"7E",X"10",X"91",X"F2",X"58",X"1A",X"ED",X"44",X"FE",X"0C",X"30",X"20",X"23",X"7E",X"FD",X"96",
		X"11",X"F2",X"66",X"1A",X"ED",X"44",X"FE",X"0A",X"30",X"12",X"3E",X"04",X"32",X"3F",X"4E",X"AF",
		X"32",X"00",X"4E",X"32",X"0A",X"4E",X"3E",X"04",X"32",X"45",X"4E",X"C9",X"11",X"08",X"00",X"DD",
		X"19",X"10",X"B4",X"DD",X"21",X"C5",X"4C",X"FD",X"21",X"00",X"4C",X"06",X"03",X"DD",X"7E",X"00",
		X"A7",X"28",X"39",X"DD",X"6E",X"04",X"DD",X"66",X"05",X"11",X"10",X"00",X"19",X"7E",X"4F",X"FD",
		X"7E",X"10",X"91",X"F2",X"A8",X"1A",X"ED",X"44",X"FE",X"0C",X"30",X"20",X"23",X"7E",X"FD",X"96",
		X"11",X"F2",X"B6",X"1A",X"ED",X"44",X"FE",X"0A",X"30",X"12",X"3E",X"04",X"32",X"3F",X"4E",X"AF",
		X"32",X"00",X"4E",X"32",X"0A",X"4E",X"3E",X"04",X"32",X"45",X"4E",X"C9",X"11",X"07",X"00",X"DD",
		X"19",X"10",X"BA",X"C9",X"3A",X"20",X"4C",X"FE",X"01",X"28",X"1D",X"3A",X"47",X"4C",X"FE",X"01",
		X"28",X"0A",X"3A",X"30",X"4C",X"E6",X"1F",X"32",X"62",X"4C",X"18",X"08",X"3A",X"2F",X"4C",X"E6",
		X"1F",X"32",X"61",X"4C",X"32",X"60",X"4C",X"C9",X"3A",X"63",X"4C",X"E6",X"1F",X"18",X"F5",X"00",
		X"00",X"00",X"01",X"00",X"03",X"00",X"05",X"2F",X"1C",X"BF",X"1B",X"2F",X"1B",X"73",X"1B",X"EB",
		X"1B",X"A7",X"1C",X"5B",X"1C",X"EB",X"1C",X"1F",X"1D",X"6B",X"1D",X"FB",X"1D",X"AF",X"1D",X"47",
		X"1E",X"AF",X"1E",X"83",X"1E",X"1F",X"1D",X"FB",X"1D",X"DB",X"1E",X"AF",X"1D",X"1F",X"1F",X"37",
		X"1B",X"48",X"1B",X"51",X"1B",X"62",X"1B",X"28",X"29",X"2A",X"2B",X"2C",X"2D",X"2E",X"2F",X"B0",
		X"B1",X"B2",X"B3",X"B4",X"B5",X"B6",X"B7",X"00",X"10",X"11",X"12",X"13",X"14",X"15",X"16",X"17",
		X"00",X"38",X"39",X"3A",X"3B",X"3C",X"3D",X"3E",X"3F",X"B0",X"B1",X"B2",X"B3",X"B4",X"B5",X"B6",
		X"B7",X"00",X"20",X"21",X"22",X"23",X"24",X"25",X"26",X"27",X"C8",X"C9",X"CA",X"CB",X"CC",X"CD",
		X"CE",X"CF",X"00",X"7B",X"1B",X"8C",X"1B",X"9D",X"1B",X"AE",X"1B",X"38",X"39",X"3A",X"3B",X"3C",
		X"3D",X"3E",X"3F",X"90",X"91",X"92",X"93",X"94",X"95",X"96",X"97",X"00",X"08",X"09",X"0A",X"0B",
		X"0C",X"0D",X"0E",X"0F",X"B8",X"B9",X"BA",X"BB",X"BC",X"BD",X"BE",X"BF",X"00",X"28",X"29",X"2A",
		X"2B",X"2C",X"2D",X"2E",X"2F",X"A0",X"A1",X"A2",X"A3",X"A4",X"A5",X"A6",X"A7",X"00",X"08",X"09",
		X"0A",X"0B",X"0C",X"0D",X"0E",X"0F",X"C8",X"C9",X"CA",X"CB",X"CC",X"CD",X"CE",X"CF",X"00",X"C7",
		X"1B",X"D0",X"1B",X"D9",X"1B",X"E2",X"1B",X"70",X"71",X"72",X"73",X"74",X"75",X"76",X"77",X"00",
		X"28",X"29",X"2A",X"2B",X"2C",X"2D",X"2E",X"2F",X"00",X"80",X"81",X"82",X"83",X"84",X"85",X"86",
		X"87",X"00",X"28",X"29",X"2A",X"2B",X"2C",X"2D",X"2E",X"2F",X"00",X"F3",X"1B",X"04",X"1C",X"0D",
		X"1C",X"1E",X"1C",X"40",X"41",X"42",X"43",X"44",X"45",X"46",X"47",X"B0",X"B1",X"B2",X"B3",X"B4",
		X"B5",X"B6",X"B7",X"00",X"08",X"09",X"0A",X"0B",X"0C",X"0D",X"0E",X"0F",X"00",X"18",X"19",X"1A",
		X"1B",X"1C",X"1D",X"1E",X"1F",X"A0",X"A1",X"A2",X"A3",X"A4",X"A5",X"A6",X"A7",X"00",X"08",X"09",
		X"0A",X"0B",X"0C",X"0D",X"0E",X"0F",X"B0",X"B1",X"B2",X"B3",X"B4",X"B5",X"B6",X"B7",X"00",X"37",
		X"1C",X"40",X"1C",X"49",X"1C",X"52",X"1C",X"70",X"71",X"72",X"73",X"74",X"75",X"76",X"77",X"00",
		X"A8",X"A9",X"AA",X"AB",X"AC",X"AD",X"AE",X"AF",X"00",X"80",X"81",X"82",X"83",X"84",X"85",X"86",
		X"87",X"00",X"50",X"51",X"52",X"53",X"54",X"55",X"56",X"57",X"00",X"63",X"1C",X"74",X"1C",X"85",
		X"1C",X"96",X"1C",X"08",X"09",X"0A",X"0B",X"0C",X"0D",X"0E",X"0F",X"90",X"91",X"92",X"93",X"94",
		X"95",X"96",X"97",X"00",X"40",X"41",X"42",X"43",X"44",X"45",X"46",X"47",X"B8",X"B9",X"BA",X"BB",
		X"BC",X"BD",X"BE",X"BF",X"00",X"08",X"09",X"0A",X"0B",X"0C",X"0D",X"0E",X"0F",X"90",X"91",X"92",
		X"93",X"94",X"95",X"96",X"97",X"00",X"38",X"39",X"3A",X"3B",X"3C",X"3D",X"3E",X"3F",X"C8",X"C9",
		X"CA",X"CB",X"CC",X"CD",X"CE",X"CF",X"00",X"AF",X"1C",X"B8",X"1C",X"C9",X"1C",X"DA",X"1C",X"40",
		X"41",X"42",X"43",X"44",X"45",X"46",X"47",X"00",X"08",X"09",X"0A",X"0B",X"0C",X"0D",X"0E",X"0F",
		X"80",X"81",X"82",X"83",X"84",X"85",X"86",X"87",X"00",X"58",X"59",X"5A",X"5B",X"5C",X"5D",X"5E",
		X"5F",X"C8",X"C9",X"CA",X"CB",X"CC",X"CD",X"CE",X"CF",X"00",X"18",X"19",X"1A",X"1B",X"1C",X"1D",
		X"1E",X"1F",X"88",X"89",X"8A",X"8B",X"8C",X"8D",X"8E",X"8F",X"00",X"F3",X"1C",X"FC",X"1C",X"05",
		X"1D",X"16",X"1D",X"60",X"61",X"62",X"63",X"64",X"65",X"66",X"67",X"00",X"88",X"89",X"8A",X"8B",
		X"8C",X"8D",X"8E",X"8F",X"00",X"08",X"09",X"0A",X"0B",X"0C",X"0D",X"0E",X"0F",X"C8",X"C9",X"CA",
		X"CB",X"CC",X"CD",X"CE",X"CF",X"00",X"40",X"41",X"42",X"43",X"44",X"45",X"46",X"47",X"00",X"27",
		X"1D",X"38",X"1D",X"49",X"1D",X"5A",X"1D",X"38",X"39",X"3A",X"3B",X"3C",X"3D",X"3E",X"3F",X"A0",
		X"A1",X"A2",X"A3",X"A4",X"A5",X"A6",X"A7",X"00",X"10",X"11",X"12",X"13",X"14",X"15",X"16",X"17",
		X"C8",X"C9",X"CA",X"CB",X"CC",X"CD",X"CE",X"CF",X"00",X"08",X"09",X"0A",X"0B",X"0C",X"0D",X"0E",
		X"0F",X"78",X"79",X"7A",X"7B",X"7C",X"7D",X"7E",X"7F",X"00",X"40",X"41",X"42",X"43",X"44",X"45",
		X"46",X"47",X"C8",X"C9",X"CA",X"CB",X"CC",X"CD",X"CE",X"CF",X"00",X"73",X"1D",X"84",X"1D",X"95",
		X"1D",X"9E",X"1D",X"28",X"29",X"2A",X"2B",X"2C",X"2D",X"2E",X"2F",X"90",X"91",X"92",X"93",X"94",
		X"95",X"96",X"97",X"00",X"08",X"09",X"0A",X"0B",X"0C",X"0D",X"0E",X"0F",X"C8",X"C9",X"CA",X"CB",
		X"CC",X"CD",X"CE",X"CF",X"00",X"60",X"61",X"62",X"63",X"64",X"65",X"66",X"67",X"00",X"18",X"19",
		X"1A",X"1B",X"1C",X"1D",X"1E",X"1F",X"C8",X"C9",X"CA",X"CB",X"CC",X"CD",X"CE",X"CF",X"00",X"B7",
		X"1D",X"C8",X"1D",X"D9",X"1D",X"EA",X"1D",X"08",X"09",X"0A",X"0B",X"0C",X"0D",X"0E",X"0F",X"C0",
		X"C1",X"C2",X"C3",X"C4",X"C5",X"C6",X"C7",X"00",X"40",X"41",X"42",X"43",X"44",X"45",X"46",X"47",
		X"90",X"91",X"92",X"93",X"94",X"95",X"96",X"97",X"00",X"48",X"49",X"4A",X"4B",X"4C",X"4D",X"4E",
		X"4F",X"C8",X"C9",X"CA",X"CB",X"CC",X"CD",X"CE",X"CF",X"00",X"08",X"09",X"0A",X"0B",X"0C",X"0D",
		X"0E",X"0F",X"88",X"89",X"8A",X"8B",X"8C",X"8D",X"8E",X"8F",X"00",X"03",X"1E",X"14",X"1E",X"25",
		X"1E",X"36",X"1E",X"40",X"41",X"42",X"43",X"44",X"45",X"46",X"47",X"80",X"81",X"82",X"83",X"84",
		X"85",X"86",X"87",X"00",X"08",X"09",X"0A",X"0B",X"0C",X"0D",X"0E",X"0F",X"B8",X"B9",X"BA",X"BB",
		X"BC",X"BD",X"BE",X"BF",X"00",X"38",X"39",X"3A",X"3B",X"3C",X"3D",X"3E",X"3F",X"C8",X"C9",X"CA",
		X"CB",X"CC",X"CD",X"CE",X"CF",X"00",X"08",X"09",X"0A",X"0B",X"0C",X"0D",X"0E",X"0F",X"B8",X"B9",
		X"BA",X"BB",X"BC",X"BD",X"BE",X"BF",X"00",X"4F",X"1E",X"60",X"1E",X"69",X"1E",X"7A",X"1E",X"08",
		X"09",X"0A",X"0B",X"0C",X"0D",X"0E",X"0F",X"C0",X"C1",X"C2",X"C3",X"C4",X"C5",X"C6",X"C7",X"00",
		X"C8",X"C9",X"CA",X"CB",X"CC",X"CD",X"CE",X"CF",X"00",X"50",X"51",X"52",X"53",X"54",X"55",X"56",
		X"57",X"98",X"99",X"9A",X"9B",X"9C",X"9D",X"9E",X"9F",X"00",X"10",X"11",X"12",X"13",X"14",X"15",
		X"16",X"17",X"00",X"8B",X"1E",X"94",X"1E",X"9D",X"1E",X"A6",X"1E",X"40",X"41",X"42",X"43",X"44",
		X"45",X"46",X"47",X"00",X"08",X"09",X"0A",X"0B",X"0C",X"0D",X"0E",X"0F",X"00",X"60",X"61",X"62",
		X"63",X"64",X"65",X"66",X"67",X"00",X"88",X"89",X"8A",X"8B",X"8C",X"8D",X"8E",X"8F",X"00",X"B7",
		X"1E",X"C0",X"1E",X"C9",X"1E",X"D2",X"1E",X"38",X"39",X"3A",X"3B",X"3C",X"3D",X"3E",X"3F",X"00",
		X"10",X"11",X"12",X"13",X"14",X"15",X"16",X"17",X"00",X"08",X"09",X"0A",X"0B",X"0C",X"0D",X"0E",
		X"0F",X"00",X"40",X"41",X"42",X"43",X"44",X"45",X"46",X"47",X"00",X"E3",X"1E",X"EC",X"1E",X"FD",
		X"1E",X"0E",X"1F",X"70",X"71",X"72",X"73",X"74",X"75",X"76",X"77",X"00",X"08",X"09",X"0A",X"0B",
		X"0C",X"0D",X"0E",X"0F",X"C8",X"C9",X"CA",X"CB",X"CC",X"CD",X"CE",X"CF",X"00",X"30",X"31",X"32",
		X"33",X"34",X"35",X"36",X"37",X"90",X"91",X"92",X"93",X"94",X"95",X"96",X"97",X"00",X"08",X"09",
		X"0A",X"0B",X"0C",X"0D",X"0E",X"0F",X"C8",X"C9",X"CA",X"CB",X"CC",X"CD",X"CE",X"CF",X"00",X"27",
		X"1F",X"38",X"1F",X"41",X"1F",X"52",X"1F",X"10",X"11",X"12",X"13",X"14",X"15",X"16",X"17",X"C0",
		X"C1",X"C2",X"C3",X"C4",X"C5",X"C6",X"C7",X"00",X"A8",X"A9",X"AA",X"AB",X"AC",X"AD",X"AE",X"AF",
		X"00",X"48",X"49",X"4A",X"4B",X"4C",X"4D",X"4E",X"4F",X"88",X"89",X"8A",X"8B",X"8C",X"8D",X"8E",
		X"8F",X"00",X"68",X"69",X"6A",X"6B",X"6C",X"6D",X"6E",X"6F",X"00",X"E8",X"22",X"4A",X"21",X"83",
		X"1F",X"6A",X"20",X"F9",X"21",X"7E",X"24",X"57",X"23",X"7D",X"25",X"84",X"26",X"AB",X"27",X"D1",
		X"29",X"8A",X"28",X"10",X"2B",X"96",X"2D",X"5F",X"2C",X"84",X"26",X"D1",X"29",X"BD",X"2E",X"8A",
		X"28",X"04",X"30",X"8D",X"1F",X"A6",X"1F",X"DF",X"1F",X"F8",X"1F",X"41",X"20",X"70",X"71",X"72",
		X"73",X"74",X"75",X"76",X"77",X"88",X"89",X"8A",X"8B",X"8C",X"8D",X"8E",X"8F",X"A0",X"A1",X"A2",
		X"A3",X"A4",X"A5",X"A6",X"A7",X"00",X"50",X"51",X"52",X"53",X"54",X"55",X"56",X"57",X"58",X"59",
		X"5A",X"5B",X"5C",X"5D",X"5E",X"5F",X"60",X"61",X"62",X"63",X"64",X"65",X"66",X"67",X"68",X"69",
		X"6A",X"6B",X"6C",X"6D",X"6E",X"6F",X"70",X"71",X"72",X"73",X"74",X"75",X"76",X"77",X"78",X"79",
		X"7A",X"7B",X"7C",X"7D",X"7E",X"7F",X"80",X"81",X"82",X"83",X"84",X"85",X"86",X"87",X"00",X"50",
		X"51",X"52",X"53",X"54",X"55",X"56",X"57",X"88",X"89",X"8A",X"8B",X"8C",X"8D",X"8E",X"8F",X"A0",
		X"A1",X"A2",X"A3",X"A4",X"A5",X"A6",X"A7",X"00",X"18",X"19",X"1A",X"1B",X"1C",X"1D",X"1E",X"1F",
		X"50",X"51",X"52",X"53",X"54",X"55",X"56",X"57",X"58",X"59",X"5A",X"5B",X"5C",X"5D",X"5E",X"5F",
		X"60",X"61",X"62",X"63",X"64",X"65",X"66",X"67",X"68",X"69",X"6A",X"6B",X"6C",X"6D",X"6E",X"6F",
		X"70",X"71",X"72",X"73",X"74",X"75",X"76",X"77",X"78",X"79",X"7A",X"7B",X"7C",X"7D",X"7E",X"7F",
		X"80",X"81",X"82",X"83",X"84",X"85",X"86",X"87",X"A0",X"A1",X"A2",X"A3",X"A4",X"A5",X"A6",X"A7",
		X"00",X"40",X"41",X"42",X"43",X"44",X"45",X"46",X"47",X"68",X"69",X"6A",X"6B",X"6C",X"6D",X"6E",
		X"6F",X"70",X"71",X"72",X"73",X"74",X"75",X"76",X"77",X"A8",X"A9",X"AA",X"AB",X"AC",X"AD",X"AE",
		X"AF",X"C0",X"C1",X"C2",X"C3",X"C4",X"C5",X"C6",X"C7",X"00",X"74",X"20",X"8D",X"20",X"B6",X"20",
		X"DF",X"20",X"08",X"21",X"80",X"81",X"82",X"83",X"84",X"85",X"86",X"87",X"A8",X"A9",X"AA",X"AB",
		X"AC",X"AD",X"AE",X"AF",X"C0",X"C1",X"C2",X"C3",X"C4",X"C5",X"C6",X"C7",X"00",X"28",X"29",X"2A",
		X"2B",X"2C",X"2D",X"2E",X"2F",X"68",X"69",X"6A",X"6B",X"6C",X"6D",X"6E",X"6F",X"70",X"71",X"72",
		X"73",X"74",X"75",X"76",X"77",X"78",X"79",X"7A",X"7B",X"7C",X"7D",X"7E",X"7F",X"B0",X"B1",X"B2",
		X"B3",X"B4",X"B5",X"B6",X"B7",X"00",X"20",X"21",X"22",X"23",X"24",X"25",X"26",X"27",X"68",X"69",
		X"6A",X"6B",X"6C",X"6D",X"6E",X"6F",X"70",X"71",X"72",X"73",X"74",X"75",X"76",X"77",X"78",X"79",
		X"7A",X"7B",X"7C",X"7D",X"7E",X"7F",X"80",X"81",X"82",X"83",X"84",X"85",X"86",X"87",X"00",X"58",
		X"59",X"5A",X"5B",X"5C",X"5D",X"5E",X"5F",X"78",X"79",X"7A",X"7B",X"7C",X"7D",X"7E",X"7F",X"80",
		X"81",X"82",X"83",X"84",X"85",X"86",X"87",X"88",X"89",X"8A",X"8B",X"8C",X"8D",X"8E",X"8F",X"B8",
		X"B9",X"BA",X"BB",X"BC",X"BD",X"BE",X"BF",X"00",X"20",X"21",X"22",X"23",X"24",X"25",X"26",X"27",
		X"40",X"41",X"42",X"43",X"44",X"45",X"46",X"47",X"60",X"61",X"62",X"63",X"64",X"65",X"66",X"67",
		X"68",X"69",X"6A",X"6B",X"6C",X"6D",X"6E",X"6F",X"70",X"71",X"72",X"73",X"74",X"75",X"76",X"77",
		X"78",X"79",X"7A",X"7B",X"7C",X"7D",X"7E",X"7F",X"A0",X"A1",X"A2",X"A3",X"A4",X"A5",X"A6",X"A7",
		X"C0",X"C1",X"C2",X"C3",X"C4",X"C5",X"C6",X"C7",X"00",X"D3",X"54",X"21",X"65",X"21",X"8E",X"21",
		X"A7",X"21",X"C8",X"21",X"60",X"61",X"62",X"63",X"64",X"65",X"66",X"67",X"A8",X"A9",X"AA",X"AB",
		X"AC",X"AD",X"AE",X"AF",X"00",X"18",X"19",X"1A",X"1B",X"1C",X"1D",X"1E",X"1F",X"50",X"51",X"52",
		X"53",X"54",X"55",X"56",X"57",X"68",X"69",X"6A",X"6B",X"6C",X"6D",X"6E",X"6F",X"90",X"91",X"92",
		X"93",X"94",X"95",X"96",X"97",X"C0",X"C1",X"C2",X"C3",X"C4",X"C5",X"C6",X"C7",X"00",X"58",X"59",
		X"5A",X"5B",X"5C",X"5D",X"5E",X"5F",X"A0",X"A1",X"A2",X"A3",X"A4",X"A5",X"A6",X"A7",X"B8",X"B9",
		X"BA",X"BB",X"BC",X"BD",X"BE",X"BF",X"00",X"48",X"49",X"4A",X"4B",X"4C",X"4D",X"4E",X"4F",X"70",
		X"71",X"72",X"73",X"74",X"75",X"76",X"77",X"98",X"99",X"9A",X"9B",X"9C",X"9D",X"9E",X"9F",X"C0",
		X"C1",X"C2",X"C3",X"C4",X"C5",X"C6",X"C7",X"00",X"18",X"19",X"1A",X"1B",X"1C",X"1D",X"1E",X"1F",
		X"48",X"49",X"4A",X"4B",X"4C",X"4D",X"4E",X"4F",X"50",X"51",X"52",X"53",X"54",X"55",X"56",X"57",
		X"68",X"69",X"6A",X"6B",X"6C",X"6D",X"6E",X"6F",X"70",X"71",X"72",X"73",X"74",X"75",X"76",X"77",
		X"88",X"89",X"8A",X"8B",X"8C",X"8D",X"8E",X"8F",X"00",X"03",X"22",X"14",X"22",X"45",X"22",X"6E",
		X"22",X"AF",X"22",X"60",X"61",X"62",X"63",X"64",X"65",X"66",X"67",X"98",X"99",X"9A",X"9B",X"9C",
		X"9D",X"9E",X"9F",X"00",X"60",X"61",X"62",X"63",X"64",X"65",X"66",X"67",X"68",X"69",X"6A",X"6B",
		X"6C",X"6D",X"6E",X"6F",X"70",X"71",X"72",X"73",X"74",X"75",X"76",X"77",X"78",X"79",X"7A",X"7B",
		X"7C",X"7D",X"7E",X"7F",X"80",X"81",X"82",X"83",X"84",X"85",X"86",X"87",X"A0",X"A1",X"A2",X"A3",
		X"A4",X"A5",X"A6",X"A7",X"00",X"30",X"31",X"32",X"33",X"34",X"35",X"36",X"37",X"48",X"49",X"4A",
		X"4B",X"4C",X"4D",X"4E",X"4F",X"60",X"61",X"62",X"63",X"64",X"65",X"66",X"67",X"90",X"91",X"92",
		X"93",X"94",X"95",X"96",X"97",X"C0",X"C1",X"C2",X"C3",X"C4",X"C5",X"C6",X"C7",X"00",X"30",X"31",
		X"32",X"33",X"34",X"35",X"36",X"37",X"50",X"51",X"52",X"53",X"54",X"55",X"56",X"57",X"58",X"59",
		X"5A",X"5B",X"5C",X"5D",X"5E",X"5F",X"60",X"61",X"62",X"63",X"64",X"65",X"66",X"67",X"68",X"69",
		X"6A",X"6B",X"6C",X"6D",X"6E",X"6F",X"70",X"71",X"72",X"73",X"74",X"75",X"76",X"77",X"78",X"79",
		X"7A",X"7B",X"7C",X"7D",X"7E",X"7F",X"80",X"81",X"82",X"83",X"84",X"85",X"86",X"87",X"00",X"28",
		X"29",X"2A",X"2B",X"2C",X"2D",X"2E",X"2F",X"40",X"41",X"42",X"43",X"44",X"45",X"46",X"47",X"60",
		X"61",X"62",X"63",X"64",X"65",X"66",X"67",X"68",X"69",X"6A",X"6B",X"6C",X"6D",X"6E",X"6F",X"70",
		X"71",X"72",X"73",X"74",X"75",X"76",X"77",X"88",X"89",X"8A",X"8B",X"8C",X"8D",X"8E",X"8F",X"90",
		X"91",X"92",X"93",X"94",X"95",X"96",X"97",X"00",X"F2",X"22",X"FB",X"22",X"04",X"23",X"1D",X"23",
		X"36",X"23",X"B8",X"B9",X"BA",X"BB",X"BC",X"BD",X"BE",X"BF",X"00",X"48",X"49",X"4A",X"4B",X"4C",
		X"4D",X"4E",X"4F",X"00",X"30",X"31",X"32",X"33",X"34",X"35",X"36",X"37",X"70",X"71",X"72",X"73",
		X"74",X"75",X"76",X"77",X"A0",X"A1",X"A2",X"A3",X"A4",X"A5",X"A6",X"A7",X"00",X"38",X"39",X"3A",
		X"3B",X"3C",X"3D",X"3E",X"3F",X"70",X"71",X"72",X"73",X"74",X"75",X"76",X"77",X"C0",X"C1",X"C2",
		X"C3",X"C4",X"C5",X"C6",X"C7",X"00",X"18",X"19",X"1A",X"1B",X"1C",X"1D",X"1E",X"1F",X"40",X"41",
		X"42",X"43",X"44",X"45",X"46",X"47",X"70",X"71",X"72",X"73",X"74",X"75",X"76",X"77",X"C0",X"C1",
		X"C2",X"C3",X"C4",X"C5",X"C6",X"C7",X"00",X"61",X"23",X"82",X"23",X"B3",X"23",X"EC",X"23",X"25",
		X"24",X"38",X"39",X"3A",X"3B",X"3C",X"3D",X"3E",X"3F",X"68",X"69",X"6A",X"6B",X"6C",X"6D",X"6E",
		X"6F",X"80",X"81",X"82",X"83",X"84",X"85",X"86",X"87",X"B0",X"B1",X"B2",X"B3",X"B4",X"B5",X"B6",
		X"B7",X"00",X"20",X"21",X"22",X"23",X"24",X"25",X"26",X"27",X"38",X"39",X"3A",X"3B",X"3C",X"3D",
		X"3E",X"3F",X"68",X"69",X"6A",X"6B",X"6C",X"6D",X"6E",X"6F",X"70",X"71",X"72",X"73",X"74",X"75",
		X"76",X"77",X"78",X"79",X"7A",X"7B",X"7C",X"7D",X"7E",X"7F",X"B0",X"B1",X"B2",X"B3",X"B4",X"B5",
		X"B6",X"B7",X"00",X"58",X"59",X"5A",X"5B",X"5C",X"5D",X"5E",X"5E",X"60",X"61",X"62",X"63",X"64",
		X"65",X"66",X"67",X"68",X"69",X"6A",X"6B",X"6C",X"6D",X"6E",X"6F",X"70",X"71",X"72",X"73",X"74",
		X"75",X"76",X"77",X"78",X"79",X"7A",X"7B",X"7C",X"7D",X"7E",X"7F",X"80",X"81",X"82",X"83",X"84",
		X"85",X"86",X"87",X"88",X"89",X"8A",X"8B",X"8C",X"8D",X"8E",X"8F",X"00",X"20",X"21",X"22",X"23",
		X"24",X"25",X"26",X"27",X"50",X"51",X"52",X"53",X"54",X"55",X"56",X"57",X"70",X"71",X"72",X"73",
		X"74",X"75",X"76",X"77",X"78",X"79",X"7A",X"7B",X"7C",X"7D",X"7E",X"7F",X"80",X"81",X"82",X"83",
		X"84",X"85",X"86",X"87",X"88",X"89",X"8A",X"8B",X"8C",X"8D",X"8E",X"8F",X"B8",X"B9",X"BA",X"BB",
		X"BC",X"BD",X"BE",X"BF",X"00",X"28",X"29",X"2A",X"2B",X"2C",X"2D",X"2E",X"2F",X"50",X"51",X"52",
		X"53",X"54",X"55",X"56",X"57",X"58",X"59",X"5A",X"5B",X"5C",X"5D",X"5E",X"5F",X"60",X"61",X"62",
		X"63",X"64",X"65",X"66",X"67",X"68",X"69",X"6A",X"6B",X"6C",X"6D",X"6E",X"6F",X"70",X"71",X"72",
		X"73",X"74",X"75",X"76",X"77",X"78",X"79",X"7A",X"7B",X"7C",X"7D",X"7E",X"7F",X"80",X"81",X"82",
		X"83",X"84",X"85",X"86",X"87",X"88",X"89",X"8A",X"8B",X"8C",X"8D",X"8E",X"8F",X"A8",X"A9",X"AA",
		X"AB",X"AC",X"AD",X"AE",X"AF",X"C0",X"C1",X"C2",X"C3",X"C4",X"C5",X"C6",X"C7",X"00",X"88",X"24",
		X"B1",X"24",X"EA",X"24",X"1B",X"25",X"54",X"25",X"60",X"61",X"62",X"63",X"64",X"65",X"66",X"67",
		X"78",X"79",X"7A",X"7B",X"7C",X"7D",X"7E",X"7F",X"80",X"81",X"82",X"83",X"84",X"85",X"86",X"87",
		X"98",X"99",X"9A",X"9B",X"9C",X"9D",X"9E",X"9F",X"B0",X"B1",X"B2",X"B3",X"B4",X"B5",X"B6",X"B7",
		X"00",X"28",X"29",X"2A",X"2B",X"2C",X"2D",X"2E",X"2F",X"68",X"69",X"6A",X"6B",X"6C",X"6D",X"6E",
		X"6F",X"70",X"71",X"72",X"73",X"74",X"75",X"76",X"77",X"78",X"79",X"7A",X"7B",X"7C",X"7D",X"7E",
		X"7F",X"98",X"99",X"9A",X"9B",X"9C",X"9D",X"9E",X"9F",X"B0",X"B1",X"B2",X"B3",X"B4",X"B5",X"B6",
		X"B7",X"B8",X"B9",X"BA",X"BB",X"BC",X"BD",X"BE",X"BF",X"00",X"28",X"29",X"2A",X"2B",X"2C",X"2D",
		X"2E",X"2F",X"30",X"31",X"32",X"33",X"34",X"35",X"36",X"37",X"70",X"71",X"72",X"73",X"74",X"75",
		X"76",X"77",X"78",X"79",X"7A",X"7B",X"7C",X"7D",X"7E",X"7F",X"A8",X"A9",X"AA",X"AB",X"AC",X"AD",
		X"AE",X"AF",X"C0",X"C1",X"C2",X"C3",X"C4",X"C5",X"C6",X"C7",X"00",X"30",X"31",X"32",X"33",X"34",
		X"35",X"36",X"37",X"50",X"51",X"52",X"53",X"54",X"55",X"56",X"57",X"70",X"71",X"72",X"73",X"74",
		X"75",X"76",X"77",X"78",X"79",X"7A",X"7B",X"7C",X"7D",X"7E",X"7F",X"80",X"81",X"82",X"83",X"84",
		X"85",X"86",X"87",X"A8",X"A9",X"AA",X"AB",X"AC",X"AD",X"AE",X"AF",X"C0",X"C1",X"C2",X"C3",X"C4",
		X"C5",X"C6",X"C7",X"00",X"40",X"41",X"42",X"43",X"44",X"45",X"46",X"47",X"60",X"61",X"62",X"63",
		X"64",X"65",X"66",X"67",X"68",X"69",X"6A",X"6B",X"6C",X"6D",X"6E",X"6F",X"70",X"71",X"72",X"73",
		X"74",X"75",X"76",X"77",X"78",X"79",X"7A",X"7B",X"7C",X"7D",X"7E",X"7F",X"00",X"87",X"25",X"A8",
		X"25",X"F1",X"25",X"1A",X"26",X"53",X"26",X"58",X"59",X"5A",X"5B",X"5C",X"5D",X"5E",X"5F",X"80",
		X"81",X"82",X"83",X"84",X"85",X"86",X"87",X"B0",X"B1",X"B2",X"B3",X"B4",X"B5",X"B6",X"B7",X"C8",
		X"C9",X"CA",X"CB",X"CC",X"CD",X"CE",X"CF",X"00",X"18",X"19",X"1A",X"1B",X"1C",X"1D",X"1E",X"1F",
		X"20",X"21",X"22",X"23",X"24",X"25",X"26",X"27",X"38",X"39",X"3A",X"3B",X"3C",X"3D",X"3E",X"3F",
		X"50",X"51",X"52",X"53",X"54",X"55",X"56",X"57",X"58",X"59",X"5A",X"5B",X"5C",X"5D",X"5E",X"5F",
		X"80",X"81",X"82",X"83",X"84",X"85",X"86",X"87",X"A0",X"A1",X"A2",X"A3",X"A4",X"A5",X"A6",X"A7",
		X"A8",X"A9",X"AA",X"AB",X"AC",X"AD",X"AE",X"AF",X"C0",X"C1",X"C2",X"C3",X"C4",X"C5",X"C6",X"C7",
		X"00",X"20",X"21",X"22",X"23",X"24",X"25",X"26",X"27",X"38",X"39",X"3A",X"3B",X"3C",X"3D",X"3E",
		X"3F",X"48",X"49",X"4A",X"4B",X"4C",X"4D",X"4E",X"4F",X"60",X"61",X"62",X"63",X"64",X"65",X"66",
		X"67",X"78",X"79",X"7A",X"7B",X"7C",X"7D",X"7E",X"7F",X"00",X"38",X"39",X"3A",X"3B",X"3C",X"3D",
		X"3E",X"3F",X"58",X"59",X"5A",X"5B",X"5C",X"5D",X"5E",X"5F",X"70",X"71",X"72",X"73",X"74",X"75",
		X"76",X"77",X"88",X"89",X"8A",X"8B",X"8C",X"8D",X"8E",X"8F",X"90",X"91",X"92",X"93",X"94",X"95",
		X"96",X"97",X"B0",X"B1",X"B2",X"B3",X"B4",X"B5",X"B6",X"B7",X"B8",X"B9",X"BA",X"BB",X"BC",X"BD",
		X"BE",X"BF",X"00",X"18",X"19",X"1A",X"1B",X"1C",X"1D",X"1E",X"1F",X"30",X"31",X"32",X"33",X"34",
		X"35",X"36",X"37",X"60",X"61",X"62",X"63",X"64",X"65",X"66",X"67",X"78",X"79",X"7A",X"7B",X"7C",
		X"7D",X"7E",X"7F",X"80",X"81",X"82",X"83",X"84",X"85",X"86",X"87",X"98",X"99",X"9A",X"9B",X"9C",
		X"9D",X"9E",X"9F",X"00",X"8E",X"26",X"B7",X"26",X"E8",X"26",X"29",X"27",X"62",X"27",X"20",X"21",
		X"22",X"23",X"24",X"25",X"26",X"27",X"50",X"51",X"52",X"53",X"54",X"55",X"56",X"57",X"68",X"69",
		X"6A",X"6B",X"6C",X"6D",X"6E",X"6F",X"80",X"81",X"82",X"83",X"84",X"85",X"86",X"87",X"98",X"99",
		X"9A",X"9B",X"9C",X"9D",X"9E",X"9F",X"00",X"50",X"51",X"52",X"53",X"54",X"55",X"56",X"57",X"58",
		X"59",X"5A",X"5B",X"5C",X"5D",X"5E",X"5F",X"60",X"61",X"62",X"63",X"64",X"65",X"66",X"67",X"68",
		X"69",X"6A",X"6B",X"6C",X"6D",X"6E",X"6F",X"70",X"71",X"72",X"73",X"74",X"75",X"76",X"77",X"98",
		X"99",X"9A",X"9B",X"9C",X"9D",X"9E",X"9F",X"00",X"28",X"29",X"2A",X"2B",X"2C",X"2D",X"2E",X"2F",
		X"48",X"49",X"4A",X"4B",X"4C",X"4D",X"4E",X"4F",X"60",X"61",X"62",X"63",X"64",X"65",X"66",X"67",
		X"68",X"69",X"6A",X"6B",X"6C",X"6D",X"6E",X"6F",X"70",X"71",X"72",X"73",X"74",X"75",X"76",X"77",
		X"90",X"91",X"92",X"93",X"94",X"95",X"96",X"97",X"A8",X"A9",X"AA",X"AB",X"AC",X"AD",X"AE",X"AF",
		X"C0",X"C1",X"C2",X"C3",X"C4",X"C5",X"C6",X"C7",X"00",X"20",X"21",X"22",X"23",X"24",X"25",X"26",
		X"27",X"38",X"39",X"3A",X"3B",X"3C",X"3D",X"3E",X"3F",X"58",X"59",X"5A",X"5B",X"5C",X"5D",X"5E",
		X"5F",X"70",X"71",X"72",X"73",X"74",X"75",X"76",X"77",X"90",X"91",X"92",X"93",X"94",X"95",X"96",
		X"97",X"A8",X"A9",X"AA",X"AB",X"AC",X"AD",X"AE",X"AF",X"C0",X"C1",X"C2",X"C3",X"C4",X"C5",X"C6",
		X"C7",X"00",X"18",X"19",X"1A",X"1B",X"1C",X"1D",X"1E",X"1F",X"20",X"21",X"22",X"23",X"24",X"25",
		X"26",X"27",X"38",X"39",X"3A",X"3B",X"3C",X"3D",X"3E",X"3F",X"58",X"59",X"5A",X"5B",X"5C",X"5D",
		X"5E",X"5F",X"60",X"61",X"62",X"63",X"64",X"65",X"66",X"67",X"68",X"69",X"6A",X"6B",X"6C",X"6D",
		X"6E",X"6F",X"70",X"71",X"72",X"73",X"74",X"75",X"76",X"77",X"A8",X"A9",X"AA",X"AB",X"AC",X"AD",
		X"AE",X"AF",X"C0",X"C1",X"C2",X"C3",X"C4",X"C5",X"C6",X"C7",X"00",X"B5",X"27",X"B6",X"27",X"E7",
		X"27",X"18",X"28",X"59",X"28",X"00",X"20",X"21",X"22",X"23",X"24",X"25",X"26",X"27",X"40",X"41",
		X"42",X"43",X"44",X"45",X"46",X"47",X"68",X"69",X"6A",X"6B",X"6C",X"6D",X"6E",X"6F",X"70",X"71",
		X"72",X"73",X"74",X"75",X"76",X"77",X"88",X"89",X"8A",X"8B",X"8C",X"8D",X"8E",X"8F",X"C0",X"C1",
		X"C2",X"C3",X"C4",X"C5",X"C6",X"C7",X"00",X"20",X"21",X"22",X"23",X"24",X"25",X"26",X"27",X"38",
		X"39",X"3A",X"3B",X"3C",X"3D",X"3E",X"3F",X"58",X"59",X"5A",X"5B",X"5C",X"5D",X"5E",X"5F",X"90",
		X"91",X"92",X"93",X"94",X"95",X"96",X"97",X"98",X"99",X"9A",X"9B",X"9C",X"9D",X"9E",X"9F",X"C0",
		X"C1",X"C2",X"C3",X"C4",X"C5",X"C6",X"C7",X"00",X"30",X"31",X"32",X"33",X"34",X"35",X"36",X"37",
		X"38",X"39",X"3A",X"3B",X"3C",X"3D",X"3E",X"3F",X"40",X"41",X"42",X"43",X"44",X"45",X"46",X"47",
		X"78",X"79",X"7A",X"7B",X"7C",X"7D",X"7E",X"7F",X"80",X"81",X"82",X"83",X"84",X"85",X"86",X"87",
		X"A0",X"A1",X"A2",X"A3",X"A4",X"A5",X"A6",X"A7",X"A8",X"A9",X"AA",X"AB",X"AC",X"AD",X"AE",X"AF",
		X"C0",X"C1",X"C2",X"C3",X"C4",X"C5",X"C6",X"C7",X"00",X"30",X"31",X"32",X"33",X"34",X"35",X"36",
		X"37",X"48",X"49",X"4A",X"4B",X"4C",X"4D",X"4E",X"4F",X"68",X"69",X"6A",X"6B",X"6C",X"6D",X"6E",
		X"6F",X"80",X"81",X"82",X"83",X"84",X"85",X"86",X"87",X"A8",X"A9",X"AA",X"AB",X"AC",X"AD",X"AE",
		X"AF",X"C0",X"C1",X"C2",X"C3",X"C4",X"C5",X"C6",X"C7",X"00",X"94",X"28",X"C5",X"28",X"FE",X"28",
		X"3F",X"29",X"88",X"29",X"20",X"21",X"22",X"23",X"24",X"25",X"26",X"27",X"38",X"39",X"3A",X"3B",
		X"3C",X"3D",X"3E",X"3F",X"50",X"51",X"52",X"53",X"54",X"55",X"56",X"57",X"68",X"69",X"6A",X"6B",
		X"6C",X"6D",X"6E",X"6F",X"80",X"81",X"82",X"83",X"84",X"85",X"86",X"87",X"98",X"99",X"9A",X"9B",
		X"9C",X"9D",X"9E",X"9F",X"00",X"20",X"21",X"22",X"23",X"24",X"25",X"26",X"27",X"38",X"39",X"3A",
		X"3B",X"3C",X"3D",X"3E",X"3F",X"58",X"59",X"5A",X"5B",X"5C",X"5D",X"5E",X"5F",X"68",X"69",X"6A",
		X"6B",X"6C",X"6D",X"6E",X"6F",X"78",X"79",X"7A",X"7B",X"7C",X"7D",X"7E",X"7F",X"88",X"89",X"8A",
		X"8B",X"8C",X"8D",X"8E",X"8F",X"A8",X"A9",X"AA",X"AB",X"AC",X"AD",X"8E",X"8F",X"00",X"18",X"19",
		X"1A",X"1B",X"1C",X"1D",X"1E",X"1F",X"38",X"39",X"3A",X"3B",X"3C",X"3D",X"3E",X"3F",X"60",X"61",
		X"62",X"63",X"64",X"65",X"66",X"67",X"68",X"69",X"6A",X"6B",X"6C",X"6D",X"6E",X"6F",X"70",X"71",
		X"72",X"73",X"74",X"75",X"76",X"77",X"78",X"79",X"7A",X"7B",X"7C",X"7D",X"7E",X"7F",X"A8",X"A9",
		X"AA",X"AB",X"AC",X"AD",X"AE",X"AF",X"C0",X"C1",X"C2",X"C3",X"C4",X"C5",X"C6",X"C7",X"00",X"20",
		X"21",X"22",X"23",X"24",X"25",X"26",X"27",X"38",X"39",X"3A",X"3B",X"3C",X"3D",X"3E",X"3F",X"40",
		X"41",X"42",X"43",X"44",X"45",X"46",X"47",X"60",X"61",X"62",X"63",X"64",X"65",X"66",X"67",X"68",
		X"69",X"6A",X"6B",X"6C",X"6D",X"6E",X"6F",X"70",X"71",X"72",X"73",X"74",X"75",X"76",X"77",X"A0",
		X"A1",X"A2",X"A3",X"A4",X"A5",X"A6",X"A7",X"A8",X"A9",X"AA",X"AB",X"AC",X"AD",X"AE",X"AF",X"C0",
		X"C1",X"C2",X"C3",X"C4",X"C5",X"C6",X"C7",X"00",X"20",X"21",X"22",X"23",X"24",X"25",X"26",X"27",
		X"38",X"39",X"3A",X"3B",X"3C",X"3D",X"3E",X"3F",X"50",X"51",X"52",X"53",X"54",X"55",X"56",X"57",
		X"68",X"69",X"6A",X"6B",X"6C",X"6D",X"6E",X"6F",X"70",X"71",X"72",X"73",X"74",X"75",X"76",X"77",
		X"78",X"79",X"7A",X"7B",X"7C",X"7D",X"7E",X"7F",X"80",X"81",X"82",X"83",X"84",X"85",X"86",X"87",
		X"A0",X"A1",X"A2",X"A3",X"A4",X"A5",X"A6",X"A7",X"B8",X"B9",X"BA",X"BB",X"BC",X"BD",X"BE",X"BF",
		X"00",X"DB",X"29",X"FC",X"29",X"45",X"2A",X"7E",X"2A",X"C7",X"2A",X"20",X"21",X"22",X"23",X"24",
		X"25",X"26",X"27",X"38",X"39",X"3A",X"3B",X"3C",X"3D",X"3E",X"3F",X"58",X"59",X"5A",X"5B",X"5C",
		X"5D",X"5E",X"5F",X"78",X"79",X"7A",X"7B",X"7C",X"7D",X"7E",X"7F",X"00",X"20",X"21",X"22",X"23",
		X"24",X"25",X"26",X"27",X"38",X"39",X"3A",X"3B",X"3C",X"3D",X"3E",X"3F",X"58",X"59",X"5A",X"5B",
		X"5C",X"5D",X"5E",X"5F",X"60",X"61",X"62",X"63",X"64",X"65",X"66",X"67",X"68",X"69",X"6A",X"6B",
		X"6C",X"6D",X"6E",X"6F",X"70",X"71",X"72",X"73",X"74",X"75",X"76",X"77",X"78",X"79",X"7A",X"7B",
		X"7C",X"7D",X"7E",X"7F",X"98",X"99",X"9A",X"9B",X"9C",X"9D",X"9E",X"9F",X"B0",X"B1",X"B2",X"B3",
		X"B4",X"B5",X"B6",X"B7",X"00",X"30",X"31",X"32",X"33",X"34",X"35",X"36",X"37",X"60",X"61",X"62",
		X"63",X"64",X"65",X"66",X"67",X"68",X"69",X"6A",X"6B",X"6C",X"6D",X"6E",X"6F",X"70",X"71",X"72",
		X"73",X"74",X"75",X"76",X"77",X"90",X"91",X"92",X"93",X"94",X"95",X"96",X"97",X"A8",X"A9",X"AA",
		X"AB",X"AC",X"AD",X"AE",X"AF",X"B0",X"B1",X"B2",X"B3",X"B4",X"B5",X"B6",X"B7",X"00",X"30",X"31",
		X"32",X"33",X"34",X"35",X"36",X"37",X"50",X"51",X"52",X"53",X"54",X"55",X"56",X"57",X"58",X"59",
		X"5A",X"5B",X"5C",X"5D",X"5E",X"5F",X"60",X"61",X"62",X"63",X"64",X"65",X"66",X"67",X"70",X"71",
		X"72",X"73",X"74",X"75",X"76",X"77",X"78",X"79",X"7A",X"7B",X"7C",X"7D",X"7E",X"7F",X"80",X"81",
		X"82",X"83",X"84",X"85",X"86",X"87",X"98",X"99",X"9A",X"9B",X"9C",X"9D",X"9E",X"9F",X"B0",X"B1",
		X"B2",X"B3",X"B4",X"B5",X"B6",X"B7",X"00",X"28",X"29",X"2A",X"2B",X"2C",X"2D",X"2E",X"2F",X"30",
		X"31",X"32",X"33",X"34",X"35",X"36",X"37",X"50",X"51",X"52",X"53",X"54",X"55",X"56",X"57",X"60",
		X"61",X"62",X"63",X"64",X"65",X"66",X"67",X"68",X"69",X"6A",X"6B",X"6C",X"6D",X"6E",X"6F",X"70",
		X"71",X"72",X"73",X"74",X"75",X"76",X"77",X"80",X"81",X"82",X"83",X"84",X"85",X"86",X"87",X"98",
		X"99",X"9A",X"9B",X"9C",X"9D",X"9E",X"9F",X"B0",X"B1",X"B2",X"B3",X"B4",X"B5",X"B6",X"B7",X"00",
		X"1A",X"2B",X"3B",X"2B",X"8C",X"2B",X"DD",X"2B",X"1E",X"2C",X"60",X"61",X"62",X"63",X"64",X"65",
		X"66",X"67",X"70",X"71",X"72",X"73",X"74",X"75",X"76",X"77",X"80",X"81",X"82",X"83",X"84",X"85",
		X"86",X"87",X"90",X"91",X"92",X"93",X"94",X"95",X"96",X"97",X"00",X"20",X"21",X"22",X"23",X"24",
		X"25",X"26",X"27",X"38",X"39",X"3A",X"3B",X"3C",X"3D",X"3E",X"3F",X"40",X"41",X"42",X"43",X"44",
		X"45",X"46",X"47",X"50",X"51",X"52",X"53",X"54",X"55",X"56",X"57",X"60",X"61",X"62",X"63",X"64",
		X"65",X"66",X"67",X"68",X"69",X"6A",X"6B",X"6C",X"6D",X"6E",X"6F",X"80",X"81",X"82",X"83",X"84",
		X"85",X"86",X"87",X"90",X"91",X"92",X"93",X"94",X"95",X"96",X"97",X"A8",X"A9",X"AA",X"AB",X"AC",
		X"AD",X"AE",X"AF",X"B8",X"B9",X"BA",X"BB",X"BC",X"BD",X"BE",X"BF",X"00",X"18",X"19",X"1A",X"1B",
		X"1C",X"1D",X"1E",X"1F",X"38",X"39",X"3A",X"3B",X"3C",X"3D",X"3E",X"3F",X"48",X"49",X"4A",X"4B",
		X"4C",X"4D",X"4E",X"4F",X"70",X"71",X"72",X"73",X"74",X"75",X"76",X"77",X"78",X"79",X"7A",X"7B",
		X"7C",X"7D",X"7E",X"7F",X"80",X"81",X"82",X"83",X"84",X"85",X"86",X"87",X"88",X"89",X"8A",X"8B",
		X"8C",X"8D",X"8E",X"8F",X"90",X"91",X"92",X"93",X"94",X"95",X"96",X"97",X"B8",X"B9",X"BA",X"BB",
		X"BC",X"BD",X"BE",X"BF",X"C0",X"C1",X"C2",X"C3",X"C4",X"C5",X"C6",X"C7",X"00",X"28",X"29",X"2A",
		X"2B",X"2C",X"2D",X"2E",X"2F",X"38",X"39",X"3A",X"3B",X"3C",X"3D",X"3E",X"3F",X"50",X"51",X"52",
		X"53",X"54",X"55",X"56",X"57",X"68",X"69",X"6A",X"6B",X"6C",X"6D",X"6E",X"6F",X"70",X"71",X"72",
		X"73",X"74",X"75",X"76",X"77",X"78",X"79",X"7A",X"7B",X"7C",X"7D",X"7E",X"7F",X"90",X"91",X"92",
		X"93",X"94",X"95",X"96",X"97",X"C0",X"C1",X"C2",X"C3",X"C4",X"C5",X"C6",X"C7",X"00",X"30",X"31",
		X"32",X"33",X"34",X"35",X"36",X"37",X"40",X"41",X"42",X"43",X"44",X"45",X"46",X"47",X"50",X"51",
		X"52",X"53",X"54",X"55",X"56",X"57",X"60",X"61",X"62",X"63",X"64",X"65",X"66",X"67",X"80",X"81",
		X"82",X"83",X"84",X"85",X"86",X"87",X"90",X"91",X"92",X"93",X"94",X"95",X"96",X"97",X"A8",X"A9",
		X"AA",X"AB",X"AC",X"AD",X"AE",X"AF",X"B8",X"B9",X"BA",X"BB",X"BC",X"BD",X"BE",X"BF",X"00",X"69",
		X"2C",X"8A",X"2C",X"CB",X"2C",X"14",X"2D",X"55",X"2D",X"60",X"61",X"62",X"63",X"64",X"65",X"66",
		X"67",X"78",X"79",X"7A",X"7B",X"7C",X"7D",X"7E",X"7F",X"98",X"99",X"9A",X"9B",X"9C",X"9D",X"9E",
		X"9F",X"B0",X"B1",X"B2",X"B3",X"B4",X"B5",X"B6",X"B7",X"00",X"28",X"29",X"2A",X"2B",X"2C",X"2D",
		X"2E",X"2F",X"68",X"69",X"6A",X"6B",X"6C",X"6D",X"6E",X"6F",X"70",X"71",X"72",X"73",X"74",X"75",
		X"76",X"77",X"78",X"79",X"7A",X"7B",X"7C",X"7D",X"7E",X"7F",X"90",X"91",X"92",X"93",X"94",X"95",
		X"96",X"97",X"98",X"99",X"9A",X"9B",X"9C",X"9D",X"9E",X"9F",X"B0",X"B1",X"B2",X"B3",X"B4",X"B5",
		X"B6",X"B7",X"B8",X"B9",X"BA",X"BB",X"BC",X"BD",X"BE",X"BF",X"00",X"20",X"21",X"22",X"23",X"24",
		X"25",X"26",X"27",X"28",X"29",X"2A",X"2B",X"2C",X"2D",X"2E",X"2F",X"30",X"31",X"32",X"33",X"34",
		X"35",X"36",X"37",X"48",X"49",X"4A",X"4B",X"4C",X"4D",X"4E",X"4F",X"50",X"51",X"52",X"53",X"54",
		X"55",X"56",X"57",X"78",X"79",X"7A",X"7B",X"7C",X"7D",X"7E",X"7F",X"90",X"91",X"92",X"93",X"94",
		X"95",X"96",X"97",X"98",X"99",X"9A",X"9B",X"9C",X"9D",X"9E",X"9F",X"A0",X"A1",X"A2",X"A3",X"A4",
		X"A5",X"A6",X"A7",X"00",X"18",X"19",X"1A",X"1B",X"1C",X"1D",X"1E",X"1F",X"28",X"29",X"2A",X"2B",
		X"2C",X"2D",X"2E",X"2F",X"38",X"39",X"3A",X"3B",X"3C",X"3D",X"3E",X"3F",X"78",X"79",X"7A",X"7B",
		X"7C",X"7D",X"7E",X"7F",X"80",X"81",X"82",X"83",X"84",X"85",X"86",X"87",X"A0",X"A1",X"A2",X"A3",
		X"A4",X"A5",X"A6",X"A7",X"B0",X"B1",X"B2",X"B3",X"B4",X"B5",X"B6",X"B7",X"C0",X"C1",X"C2",X"C3",
		X"C4",X"C5",X"C6",X"C7",X"00",X"38",X"39",X"3A",X"3B",X"3C",X"3D",X"3E",X"3F",X"48",X"49",X"4A",
		X"4B",X"4C",X"4D",X"4E",X"4F",X"50",X"51",X"52",X"53",X"54",X"55",X"56",X"57",X"58",X"59",X"5A",
		X"5B",X"5C",X"5D",X"5E",X"5F",X"68",X"69",X"6A",X"6B",X"6C",X"6D",X"6E",X"6F",X"78",X"79",X"7A",
		X"7B",X"7C",X"7D",X"7E",X"7F",X"B0",X"B1",X"B2",X"B3",X"B4",X"B5",X"B6",X"B7",X"C0",X"C1",X"C2",
		X"C3",X"C4",X"C5",X"C6",X"C7",X"00",X"A0",X"2D",X"C1",X"2D",X"DA",X"2D",X"3B",X"2E",X"74",X"2E",
		X"20",X"21",X"22",X"23",X"24",X"25",X"26",X"27",X"60",X"61",X"62",X"63",X"64",X"65",X"66",X"67",
		X"78",X"79",X"7A",X"7B",X"7C",X"7D",X"7E",X"7F",X"88",X"89",X"8A",X"8B",X"8C",X"8D",X"8E",X"8F",
		X"00",X"58",X"59",X"5A",X"5B",X"5C",X"5D",X"5E",X"5F",X"98",X"99",X"9A",X"9B",X"9C",X"9D",X"9E",
		X"9F",X"B8",X"B9",X"BA",X"BB",X"BC",X"BD",X"BE",X"BF",X"00",X"28",X"29",X"2A",X"2B",X"2C",X"2D",
		X"2E",X"2F",X"38",X"39",X"3A",X"3B",X"3C",X"3D",X"3E",X"3F",X"48",X"49",X"4A",X"4B",X"4C",X"4D",
		X"4E",X"4F",X"50",X"51",X"52",X"53",X"54",X"55",X"56",X"57",X"58",X"59",X"5A",X"5B",X"5C",X"5D",
		X"5E",X"5F",X"68",X"69",X"6A",X"6B",X"6C",X"6D",X"6E",X"6F",X"80",X"81",X"82",X"83",X"84",X"85",
		X"86",X"87",X"90",X"91",X"92",X"93",X"94",X"95",X"96",X"97",X"98",X"99",X"9A",X"9B",X"9C",X"9D",
		X"9E",X"9F",X"B0",X"B1",X"B2",X"B3",X"B4",X"B5",X"B6",X"B7",X"B8",X"B9",X"BA",X"BB",X"BC",X"BD",
		X"BE",X"BF",X"C0",X"C1",X"C2",X"C3",X"C4",X"C5",X"C6",X"C7",X"00",X"20",X"21",X"22",X"23",X"24",
		X"25",X"26",X"27",X"38",X"39",X"3A",X"3B",X"3C",X"3D",X"3E",X"3F",X"58",X"59",X"5A",X"5B",X"5C",
		X"5D",X"5E",X"5F",X"70",X"71",X"72",X"73",X"74",X"75",X"76",X"77",X"90",X"91",X"92",X"93",X"94",
		X"95",X"96",X"97",X"A8",X"A9",X"AA",X"AB",X"AC",X"AD",X"AE",X"AF",X"C0",X"C1",X"C2",X"C3",X"C4",
		X"C5",X"C6",X"C7",X"00",X"18",X"19",X"1A",X"1B",X"1C",X"1D",X"1E",X"1F",X"20",X"21",X"22",X"23",
		X"24",X"25",X"26",X"27",X"38",X"39",X"3A",X"3B",X"3C",X"3D",X"3E",X"3F",X"58",X"59",X"5A",X"5B",
		X"5C",X"5D",X"5E",X"5F",X"68",X"69",X"6A",X"6B",X"6C",X"6D",X"6E",X"6F",X"78",X"79",X"7A",X"7B",
		X"7C",X"7D",X"7E",X"7F",X"80",X"81",X"82",X"83",X"84",X"85",X"86",X"87",X"A8",X"A9",X"AA",X"AB",
		X"AC",X"AD",X"AE",X"AF",X"B0",X"B1",X"B2",X"B3",X"B4",X"B5",X"B6",X"B7",X"00",X"C7",X"2E",X"00",
		X"2F",X"39",X"2F",X"8A",X"2F",X"BB",X"2F",X"30",X"31",X"32",X"33",X"34",X"35",X"36",X"37",X"48",
		X"49",X"4A",X"4B",X"4C",X"4D",X"4E",X"4F",X"88",X"89",X"8A",X"8B",X"8C",X"8D",X"8E",X"8F",X"90",
		X"91",X"92",X"93",X"94",X"95",X"96",X"97",X"A8",X"A9",X"AA",X"AB",X"AC",X"AD",X"AE",X"AF",X"C0",
		X"C1",X"C2",X"C3",X"C4",X"C5",X"C6",X"C7",X"C8",X"C9",X"CA",X"CB",X"CC",X"CD",X"CE",X"CF",X"00",
		X"20",X"21",X"22",X"23",X"24",X"25",X"26",X"27",X"38",X"39",X"3A",X"3B",X"3C",X"3D",X"3E",X"3F",
		X"48",X"49",X"4A",X"4B",X"4C",X"4D",X"4E",X"4F",X"88",X"89",X"8A",X"8B",X"8C",X"8D",X"8E",X"8F",
		X"98",X"99",X"9A",X"9B",X"9C",X"9D",X"9E",X"9F",X"B0",X"B1",X"B2",X"B3",X"B4",X"B5",X"B6",X"B7",
		X"C0",X"C1",X"C2",X"C3",X"C4",X"C5",X"C6",X"C7",X"00",X"20",X"21",X"22",X"23",X"24",X"25",X"26",
		X"27",X"28",X"29",X"2A",X"2B",X"2C",X"2D",X"2E",X"2F",X"48",X"49",X"4A",X"4B",X"4C",X"4D",X"4E",
		X"4F",X"50",X"51",X"52",X"53",X"54",X"55",X"56",X"57",X"68",X"69",X"6A",X"6B",X"6C",X"6D",X"6E",
		X"6F",X"80",X"81",X"82",X"83",X"84",X"85",X"86",X"87",X"88",X"89",X"8A",X"8B",X"8C",X"8D",X"8E",
		X"8F",X"A8",X"A9",X"AA",X"AB",X"AC",X"AD",X"AE",X"AF",X"B0",X"B1",X"B2",X"B3",X"B4",X"B5",X"B6",
		X"B7",X"B8",X"B9",X"BA",X"BB",X"BC",X"BD",X"BE",X"BF",X"00",X"48",X"49",X"4A",X"4B",X"4C",X"4D",
		X"4E",X"4F",X"58",X"59",X"5A",X"5B",X"5C",X"5D",X"5E",X"5F",X"60",X"61",X"62",X"63",X"64",X"65",
		X"66",X"67",X"78",X"79",X"7A",X"7B",X"7C",X"7D",X"7E",X"7F",X"80",X"81",X"82",X"83",X"84",X"85",
		X"86",X"87",X"B0",X"B1",X"B2",X"B3",X"B4",X"B5",X"B6",X"B7",X"00",X"20",X"21",X"22",X"23",X"24",
		X"25",X"26",X"27",X"28",X"29",X"2A",X"2B",X"2C",X"2D",X"2E",X"2F",X"50",X"51",X"52",X"53",X"54",
		X"55",X"56",X"57",X"60",X"61",X"62",X"63",X"64",X"65",X"66",X"67",X"70",X"71",X"72",X"73",X"74",
		X"75",X"76",X"77",X"80",X"81",X"82",X"83",X"84",X"85",X"86",X"87",X"88",X"89",X"8A",X"8B",X"8C",
		X"8D",X"8E",X"8F",X"B0",X"B1",X"B2",X"B3",X"B4",X"B5",X"B6",X"B7",X"C0",X"C1",X"C2",X"C3",X"C4",
		X"C5",X"C6",X"C7",X"00",X"0E",X"30",X"37",X"30",X"78",X"30",X"99",X"30",X"DA",X"30",X"58",X"59",
		X"5A",X"5B",X"5C",X"5D",X"5E",X"5F",X"60",X"61",X"62",X"63",X"64",X"65",X"66",X"67",X"78",X"79",
		X"7A",X"7B",X"7C",X"7D",X"7E",X"7F",X"80",X"81",X"82",X"83",X"84",X"85",X"86",X"87",X"88",X"89",
		X"8A",X"8B",X"8C",X"8D",X"8E",X"8F",X"00",X"28",X"29",X"2A",X"2B",X"2C",X"2D",X"2E",X"2F",X"40",
		X"41",X"42",X"43",X"44",X"45",X"46",X"47",X"48",X"49",X"4A",X"4B",X"4C",X"4D",X"4E",X"4F",X"50",
		X"51",X"52",X"53",X"54",X"55",X"56",X"57",X"60",X"61",X"62",X"63",X"64",X"65",X"66",X"67",X"88",
		X"89",X"8A",X"8B",X"8C",X"8D",X"8E",X"8F",X"98",X"99",X"9A",X"9B",X"9C",X"9D",X"9E",X"9F",X"A0",
		X"A1",X"A2",X"A3",X"A4",X"A5",X"A6",X"A7",X"00",X"68",X"69",X"6A",X"6B",X"6C",X"6D",X"6E",X"6F",
		X"70",X"71",X"72",X"73",X"74",X"75",X"76",X"77",X"78",X"79",X"7A",X"7B",X"7C",X"7D",X"7E",X"7F",
		X"C0",X"C1",X"C2",X"C3",X"C4",X"C5",X"C6",X"C7",X"00",X"30",X"31",X"32",X"33",X"34",X"35",X"36",
		X"37",X"38",X"39",X"3A",X"3B",X"3C",X"3D",X"3E",X"3F",X"40",X"41",X"42",X"43",X"44",X"45",X"46",
		X"47",X"60",X"61",X"62",X"63",X"64",X"65",X"66",X"67",X"80",X"81",X"82",X"83",X"84",X"85",X"86",
		X"87",X"A0",X"A1",X"A2",X"A3",X"A4",X"A5",X"A6",X"A7",X"A8",X"A9",X"AA",X"AB",X"AC",X"AD",X"AE",
		X"AF",X"B8",X"B9",X"BA",X"BB",X"BC",X"BD",X"BE",X"BF",X"00",X"18",X"19",X"1A",X"1B",X"1C",X"1D",
		X"1E",X"1F",X"28",X"29",X"2A",X"2B",X"2C",X"2D",X"2E",X"2F",X"38",X"39",X"3A",X"3B",X"3C",X"3D",
		X"3E",X"3F",X"50",X"51",X"52",X"53",X"54",X"55",X"56",X"57",X"60",X"61",X"62",X"63",X"64",X"65",
		X"66",X"67",X"88",X"89",X"8A",X"8B",X"8C",X"8D",X"8E",X"8F",X"98",X"99",X"9A",X"9B",X"9C",X"9D",
		X"9E",X"9F",X"B0",X"B1",X"B2",X"B3",X"B4",X"B5",X"B6",X"B7",X"C0",X"C1",X"C2",X"C3",X"C4",X"C5",
		X"C6",X"C7",X"00",X"46",X"3A",X"4E",X"4C",X"3D",X"21",X"00",X"80",X"16",X"00",X"5F",X"19",X"7E",
		X"21",X"14",X"80",X"E6",X"1F",X"87",X"16",X"00",X"5F",X"19",X"5E",X"23",X"56",X"1A",X"4F",X"21",
		X"40",X"41",X"DD",X"21",X"00",X"04",X"EB",X"DD",X"19",X"EB",X"1A",X"FE",X"FF",X"28",X"40",X"FE",
		X"00",X"28",X"11",X"FE",X"01",X"28",X"22",X"77",X"13",X"1A",X"4F",X"DD",X"71",X"00",X"13",X"23",
		X"DD",X"23",X"18",X"E6",X"7D",X"E6",X"E0",X"C6",X"20",X"6F",X"3E",X"00",X"8C",X"67",X"DD",X"21",
		X"00",X"04",X"EB",X"DD",X"19",X"EB",X"13",X"18",X"D1",X"13",X"1A",X"47",X"13",X"1A",X"08",X"13",
		X"1A",X"4F",X"08",X"13",X"77",X"DD",X"71",X"00",X"23",X"DD",X"23",X"10",X"F7",X"18",X"BB",X"F7",
		X"CD",X"03",X"00",X"CD",X"24",X"00",X"C9",X"21",X"E0",X"40",X"DD",X"21",X"00",X"04",X"EB",X"DD",
		X"19",X"EB",X"3E",X"3D",X"0E",X"05",X"06",X"1C",X"77",X"DD",X"71",X"00",X"23",X"DD",X"23",X"10",
		X"F7",X"21",X"60",X"43",X"DD",X"21",X"00",X"04",X"EB",X"DD",X"19",X"EB",X"3E",X"3E",X"06",X"20",
		X"77",X"DD",X"71",X"00",X"23",X"DD",X"23",X"10",X"F7",X"21",X"9C",X"40",X"DD",X"21",X"00",X"04",
		X"EB",X"DD",X"19",X"EB",X"11",X"20",X"00",X"3E",X"3F",X"06",X"14",X"77",X"DD",X"71",X"00",X"19",
		X"DD",X"19",X"10",X"F7",X"21",X"96",X"40",X"DD",X"21",X"96",X"44",X"3E",X"1B",X"0E",X"E0",X"06",
		X"14",X"71",X"DD",X"77",X"00",X"2B",X"DD",X"2B",X"10",X"F7",X"C9",X"3A",X"4E",X"4C",X"3D",X"87",
		X"21",X"B4",X"94",X"16",X"00",X"5F",X"19",X"EB",X"21",X"A8",X"40",X"0E",X"0A",X"1A",X"47",X"13",
		X"1A",X"13",X"C5",X"D5",X"E5",X"CD",X"D7",X"00",X"E1",X"D1",X"C1",X"23",X"23",X"0D",X"20",X"ED",
		X"C9",X"21",X"DD",X"40",X"11",X"40",X"00",X"3E",X"0F",X"06",X"00",X"0E",X"08",X"F5",X"C5",X"D5",
		X"E5",X"CD",X"D7",X"00",X"E1",X"D1",X"C1",X"F1",X"19",X"0D",X"20",X"F1",X"C9",X"21",X"DD",X"40",
		X"3A",X"4D",X"4C",X"A7",X"28",X"07",X"47",X"11",X"40",X"00",X"19",X"10",X"FD",X"E5",X"3A",X"4E",
		X"4C",X"3D",X"87",X"4F",X"87",X"47",X"3E",X"70",X"80",X"47",X"16",X"00",X"59",X"21",X"C6",X"94",
		X"19",X"78",X"46",X"E1",X"C3",X"D7",X"00",X"3A",X"4E",X"4C",X"3D",X"87",X"21",X"26",X"96",X"5F",
		X"16",X"00",X"19",X"5E",X"23",X"56",X"1A",X"FE",X"FF",X"C8",X"EB",X"23",X"5E",X"23",X"56",X"23",
		X"EB",X"A7",X"28",X"0C",X"1A",X"47",X"13",X"1A",X"13",X"D5",X"CD",X"D7",X"00",X"D1",X"18",X"E6",
		X"1A",X"4F",X"DD",X"21",X"00",X"04",X"EB",X"DD",X"19",X"EB",X"DD",X"71",X"00",X"13",X"1A",X"77",
		X"13",X"18",X"D3",X"3A",X"4E",X"4C",X"3D",X"87",X"21",X"EE",X"94",X"16",X"00",X"5F",X"19",X"5E",
		X"23",X"56",X"DD",X"21",X"02",X"4C",X"06",X"04",X"1A",X"DD",X"77",X"00",X"13",X"1A",X"DD",X"77",
		X"01",X"13",X"1A",X"DD",X"77",X"11",X"13",X"1A",X"DD",X"77",X"10",X"13",X"DD",X"23",X"DD",X"23",
		X"10",X"E6",X"C9",X"3A",X"4C",X"4C",X"A7",X"C0",X"3A",X"34",X"4C",X"A7",X"C8",X"3A",X"66",X"4C",
		X"A7",X"C8",X"21",X"65",X"4C",X"35",X"C0",X"36",X"26",X"2B",X"35",X"28",X"4C",X"7E",X"FE",X"0F",
		X"38",X"41",X"FE",X"32",X"38",X"39",X"0E",X"1B",X"7E",X"47",X"E6",X"07",X"57",X"78",X"0F",X"0F",
		X"0F",X"E6",X"1F",X"47",X"FE",X"00",X"21",X"96",X"40",X"DD",X"21",X"96",X"44",X"3E",X"E0",X"28",
		X"09",X"77",X"DD",X"71",X"00",X"2B",X"DD",X"2B",X"10",X"F7",X"7A",X"A7",X"28",X"09",X"3E",X"01",
		X"82",X"3D",X"77",X"DD",X"71",X"00",X"C9",X"3E",X"0A",X"77",X"DD",X"36",X"00",X"00",X"C9",X"0E",
		X"18",X"18",X"02",X"0E",X"1D",X"3E",X"01",X"18",X"BF",X"3E",X"04",X"32",X"3F",X"4E",X"AF",X"32",
		X"00",X"4E",X"32",X"0A",X"4E",X"3E",X"04",X"32",X"45",X"4E",X"C9",X"CD",X"F7",X"05",X"3A",X"64",
		X"4C",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"21",X"82",X"33",X"87",X"16",X"00",X"5F",X"19",X"5E",
		X"23",X"56",X"21",X"43",X"4C",X"73",X"23",X"72",X"D5",X"F5",X"CD",X"F7",X"05",X"F1",X"D1",X"21",
		X"67",X"4C",X"36",X"00",X"23",X"72",X"23",X"73",X"11",X"67",X"4C",X"21",X"90",X"41",X"CD",X"99",
		X"03",X"C9",X"05",X"00",X"10",X"00",X"50",X"00",X"00",X"01",X"00",X"05",X"00",X"10",X"00",X"50",
		X"00",X"70",X"00",X"80",X"00",X"90",X"3A",X"4E",X"4C",X"3D",X"87",X"21",X"70",X"9C",X"16",X"00",
		X"5F",X"19",X"5E",X"23",X"56",X"21",X"6A",X"4C",X"EB",X"01",X"25",X"00",X"ED",X"B0",X"21",X"00",
		X"00",X"22",X"43",X"4C",X"AF",X"32",X"DA",X"4C",X"32",X"A9",X"4C",X"32",X"B1",X"4C",X"32",X"B9",
		X"4C",X"32",X"C1",X"4C",X"3A",X"4E",X"4C",X"3D",X"87",X"21",X"0D",X"9F",X"16",X"00",X"5F",X"19",
		X"5E",X"23",X"56",X"21",X"8F",X"4C",X"EB",X"01",X"15",X"00",X"ED",X"B0",X"AF",X"32",X"A4",X"4C",
		X"C9",X"3A",X"A4",X"4C",X"87",X"21",X"9A",X"A0",X"16",X"00",X"5F",X"19",X"11",X"43",X"4C",X"7E",
		X"12",X"23",X"13",X"7E",X"12",X"C9",X"3A",X"4E",X"4C",X"3D",X"21",X"B2",X"A0",X"87",X"16",X"00",
		X"5F",X"19",X"5E",X"23",X"56",X"21",X"C5",X"4C",X"DD",X"21",X"0A",X"4C",X"1A",X"FE",X"FF",X"C8",
		X"DD",X"77",X"00",X"13",X"1A",X"DD",X"77",X"01",X"13",X"1A",X"DD",X"77",X"10",X"13",X"1A",X"DD",
		X"77",X"11",X"36",X"01",X"13",X"23",X"06",X"06",X"1A",X"77",X"13",X"23",X"10",X"FA",X"DD",X"23",
		X"DD",X"23",X"18",X"D8",X"21",X"DA",X"4C",X"06",X"24",X"AF",X"77",X"23",X"10",X"FC",X"21",X"C5",
		X"4C",X"06",X"15",X"77",X"23",X"10",X"FC",X"21",X"A5",X"4C",X"06",X"20",X"77",X"23",X"10",X"FC",
		X"C9",X"CD",X"7E",X"34",X"3A",X"47",X"4C",X"FE",X"01",X"20",X"05",X"21",X"48",X"4C",X"18",X"03",
		X"21",X"49",X"4C",X"7E",X"FE",X"00",X"C8",X"4F",X"21",X"81",X"43",X"06",X"14",X"3E",X"FC",X"F5",
		X"C5",X"E5",X"CD",X"D7",X"00",X"E1",X"C1",X"F1",X"23",X"23",X"0D",X"20",X"F2",X"C9",X"DD",X"21",
		X"81",X"43",X"3E",X"0F",X"06",X"10",X"DD",X"77",X"00",X"DD",X"77",X"20",X"DD",X"23",X"10",X"F6",
		X"C9",X"3A",X"20",X"4C",X"3D",X"20",X"10",X"3A",X"53",X"4E",X"A7",X"28",X"0A",X"AF",X"32",X"45",
		X"4E",X"3E",X"0C",X"32",X"46",X"4E",X"C9",X"AF",X"32",X"C0",X"50",X"3A",X"45",X"4E",X"A7",X"28",
		X"28",X"3D",X"47",X"3A",X"46",X"4E",X"FE",X"0C",X"28",X"05",X"B8",X"28",X"29",X"38",X"20",X"78",
		X"32",X"46",X"4E",X"CD",X"7E",X"35",X"CD",X"9B",X"35",X"CD",X"C2",X"35",X"CD",X"F0",X"35",X"3E",
		X"01",X"32",X"01",X"50",X"AF",X"32",X"45",X"4E",X"C9",X"3A",X"46",X"4E",X"FE",X"0C",X"C8",X"CD",
		X"ED",X"34",X"CD",X"27",X"35",X"C9",X"FE",X"07",X"28",X"F5",X"C3",X"BD",X"34",X"3A",X"42",X"4E",
		X"A7",X"CA",X"00",X"35",X"3A",X"42",X"4E",X"FE",X"FF",X"CA",X"00",X"35",X"3D",X"32",X"42",X"4E",
		X"3A",X"43",X"4E",X"A7",X"CA",X"13",X"35",X"3A",X"43",X"4E",X"FE",X"FF",X"CA",X"13",X"35",X"3D",
		X"32",X"43",X"4E",X"3A",X"44",X"4E",X"A7",X"CA",X"26",X"35",X"3A",X"44",X"4E",X"FE",X"FF",X"CA",
		X"26",X"35",X"3D",X"32",X"44",X"4E",X"C9",X"3A",X"42",X"4E",X"FE",X"00",X"CA",X"3A",X"35",X"3A",
		X"42",X"4E",X"FE",X"FF",X"CA",X"71",X"35",X"C3",X"40",X"35",X"CD",X"CC",X"35",X"CD",X"FA",X"35",
		X"3A",X"43",X"4E",X"FE",X"00",X"CA",X"53",X"35",X"3A",X"43",X"4E",X"FE",X"FF",X"CA",X"71",X"35",
		X"C3",X"59",X"35",X"CD",X"D8",X"35",X"CD",X"1A",X"36",X"3A",X"44",X"4E",X"FE",X"00",X"CA",X"6A",
		X"35",X"3A",X"44",X"4E",X"FE",X"FF",X"CA",X"71",X"35",X"C9",X"CD",X"E4",X"35",X"CD",X"35",X"36",
		X"C9",X"3E",X"0B",X"32",X"46",X"4E",X"AF",X"32",X"4D",X"4E",X"32",X"01",X"50",X"C9",X"21",X"1C",
		X"A3",X"3A",X"46",X"4E",X"87",X"16",X"00",X"5F",X"19",X"5E",X"23",X"56",X"1A",X"32",X"45",X"50",
		X"13",X"1A",X"32",X"4A",X"50",X"13",X"1A",X"32",X"4F",X"50",X"C9",X"21",X"58",X"A3",X"3A",X"46",
		X"4E",X"87",X"16",X"00",X"5F",X"19",X"5E",X"23",X"56",X"EB",X"5E",X"23",X"56",X"ED",X"53",X"47",
		X"4E",X"23",X"5E",X"23",X"56",X"ED",X"53",X"49",X"4E",X"23",X"5E",X"23",X"56",X"ED",X"53",X"4B",
		X"4E",X"C9",X"CD",X"CC",X"35",X"CD",X"D8",X"35",X"CD",X"E4",X"35",X"C9",X"2A",X"47",X"4E",X"7E",
		X"32",X"42",X"4E",X"23",X"22",X"47",X"4E",X"C9",X"2A",X"49",X"4E",X"7E",X"32",X"43",X"4E",X"23",
		X"22",X"49",X"4E",X"C9",X"2A",X"4B",X"4E",X"7E",X"32",X"44",X"4E",X"23",X"22",X"4B",X"4E",X"C9",
		X"CD",X"FA",X"35",X"CD",X"1A",X"36",X"CD",X"35",X"36",X"C9",X"2A",X"47",X"4E",X"7E",X"32",X"55",
		X"50",X"23",X"7E",X"32",X"50",X"50",X"23",X"7E",X"32",X"51",X"50",X"23",X"7E",X"32",X"52",X"50",
		X"23",X"7E",X"32",X"53",X"50",X"23",X"22",X"47",X"4E",X"C9",X"2A",X"49",X"4E",X"7E",X"32",X"5A",
		X"50",X"23",X"7E",X"32",X"56",X"50",X"23",X"7E",X"32",X"57",X"50",X"23",X"7E",X"32",X"58",X"50",
		X"23",X"22",X"49",X"4E",X"C9",X"2A",X"4B",X"4E",X"7E",X"32",X"5F",X"50",X"23",X"7E",X"32",X"5B",
		X"50",X"23",X"7E",X"32",X"5C",X"50",X"23",X"7E",X"32",X"5D",X"50",X"23",X"22",X"4B",X"4E",X"C9",
		X"CD",X"57",X"36",X"CD",X"ED",X"36",X"C9",X"DD",X"21",X"A5",X"4C",X"06",X"04",X"DD",X"7E",X"04",
		X"A7",X"C2",X"C8",X"36",X"DD",X"7E",X"00",X"A7",X"CA",X"BF",X"36",X"DD",X"35",X"03",X"C2",X"BF",
		X"36",X"DD",X"7E",X"07",X"DD",X"77",X"03",X"DD",X"6E",X"05",X"DD",X"66",X"06",X"11",X"11",X"00",
		X"19",X"7E",X"FE",X"00",X"28",X"2F",X"38",X"2D",X"FE",X"CF",X"28",X"29",X"30",X"27",X"DD",X"CB",
		X"01",X"46",X"28",X"07",X"7E",X"DD",X"96",X"02",X"77",X"18",X"05",X"7E",X"DD",X"86",X"02",X"77",
		X"DD",X"7E",X"02",X"DD",X"4E",X"01",X"DD",X"6E",X"05",X"DD",X"66",X"06",X"7E",X"E6",X"FE",X"B1",
		X"EE",X"05",X"77",X"18",X"0A",X"DD",X"7E",X"01",X"EE",X"01",X"DD",X"77",X"01",X"18",X"CF",X"11",
		X"08",X"00",X"DD",X"19",X"05",X"20",X"96",X"C9",X"DD",X"35",X"04",X"28",X"15",X"DD",X"6E",X"05",
		X"DD",X"66",X"06",X"23",X"DD",X"CB",X"04",X"4E",X"28",X"04",X"36",X"15",X"18",X"E1",X"36",X"00",
		X"18",X"DD",X"DD",X"6E",X"05",X"DD",X"66",X"06",X"23",X"36",X"15",X"18",X"D2",X"DD",X"21",X"C5",
		X"4C",X"06",X"03",X"DD",X"7E",X"00",X"A7",X"CA",X"4E",X"37",X"DD",X"35",X"03",X"C2",X"4E",X"37",
		X"DD",X"7E",X"06",X"DD",X"77",X"03",X"DD",X"6E",X"04",X"DD",X"66",X"05",X"11",X"11",X"00",X"19",
		X"7E",X"FE",X"00",X"28",X"2F",X"38",X"2D",X"FE",X"D0",X"28",X"29",X"30",X"27",X"DD",X"CB",X"01",
		X"46",X"28",X"07",X"7E",X"DD",X"96",X"02",X"77",X"18",X"05",X"7E",X"DD",X"86",X"02",X"77",X"DD",
		X"7E",X"02",X"DD",X"4E",X"01",X"DD",X"6E",X"04",X"DD",X"66",X"05",X"7E",X"E6",X"FE",X"B1",X"EE",
		X"05",X"77",X"18",X"0A",X"DD",X"7E",X"01",X"EE",X"01",X"DD",X"77",X"01",X"18",X"CF",X"11",X"07",
		X"00",X"DD",X"19",X"05",X"20",X"9D",X"C9",X"CD",X"64",X"37",X"CD",X"D3",X"37",X"CD",X"9D",X"38",
		X"CD",X"C9",X"38",X"C9",X"21",X"6A",X"4C",X"3A",X"5A",X"4C",X"3D",X"47",X"28",X"08",X"7E",X"23",
		X"FE",X"FF",X"20",X"FA",X"10",X"F8",X"06",X"08",X"11",X"04",X"00",X"3A",X"11",X"4C",X"E6",X"FC",
		X"4F",X"7E",X"FE",X"FF",X"C8",X"B9",X"28",X"04",X"19",X"10",X"F6",X"C9",X"36",X"F8",X"23",X"23",
		X"5E",X"23",X"56",X"21",X"DA",X"4C",X"06",X"08",X"7E",X"A7",X"28",X"06",X"23",X"23",X"23",X"10",
		X"F7",X"C9",X"36",X"50",X"23",X"73",X"23",X"72",X"3A",X"A4",X"4C",X"87",X"87",X"C6",X"40",X"EB",
		X"06",X"05",X"CD",X"D7",X"00",X"CD",X"E1",X"33",X"21",X"4D",X"4C",X"35",X"21",X"A4",X"4C",X"34",
		X"CD",X"3D",X"32",X"3E",X"06",X"32",X"45",X"4E",X"3A",X"4D",X"4C",X"A7",X"C0",X"3E",X"01",X"32",
		X"4F",X"4C",X"C9",X"21",X"8F",X"4C",X"3A",X"5A",X"4C",X"3D",X"47",X"28",X"08",X"7E",X"23",X"FE",
		X"FF",X"20",X"FA",X"10",X"F8",X"06",X"08",X"11",X"04",X"00",X"3A",X"11",X"4C",X"4F",X"7E",X"FE",
		X"FF",X"C8",X"E6",X"FC",X"B9",X"28",X"04",X"19",X"10",X"F4",X"C9",X"36",X"F8",X"23",X"7E",X"23",
		X"5E",X"23",X"56",X"4F",X"08",X"79",X"E6",X"0F",X"FE",X"03",X"CA",X"39",X"38",X"21",X"F2",X"4C",
		X"06",X"04",X"7E",X"A7",X"28",X"06",X"23",X"23",X"23",X"10",X"F7",X"C9",X"36",X"50",X"23",X"73",
		X"23",X"72",X"21",X"A4",X"4C",X"7E",X"34",X"87",X"87",X"C6",X"40",X"12",X"13",X"3E",X"05",X"12",
		X"CD",X"E1",X"33",X"3E",X"06",X"32",X"45",X"4E",X"C9",X"3E",X"05",X"32",X"45",X"4E",X"EB",X"E5",
		X"DD",X"E1",X"0E",X"F0",X"3A",X"53",X"4C",X"CB",X"47",X"28",X"04",X"79",X"EE",X"01",X"4F",X"71",
		X"23",X"36",X"14",X"21",X"A5",X"4C",X"11",X"08",X"00",X"06",X"04",X"7E",X"A7",X"28",X"04",X"19",
		X"10",X"F9",X"C9",X"36",X"01",X"23",X"3A",X"53",X"4C",X"CB",X"47",X"28",X"03",X"AF",X"18",X"02",
		X"3E",X"01",X"77",X"23",X"E5",X"21",X"C1",X"A2",X"08",X"07",X"07",X"07",X"07",X"E6",X"0F",X"87",
		X"16",X"00",X"5F",X"19",X"5E",X"23",X"56",X"E1",X"1A",X"77",X"13",X"23",X"1A",X"77",X"4F",X"13",
		X"23",X"1A",X"77",X"23",X"DD",X"E5",X"D1",X"73",X"23",X"72",X"23",X"71",X"C9",X"DD",X"21",X"DA",
		X"4C",X"06",X"08",X"DD",X"7E",X"00",X"A7",X"28",X"18",X"DD",X"35",X"00",X"20",X"13",X"DD",X"6E",
		X"01",X"DD",X"66",X"02",X"3E",X"0F",X"C5",X"06",X"00",X"DD",X"E5",X"CD",X"D7",X"00",X"DD",X"E1",
		X"C1",X"11",X"03",X"00",X"DD",X"19",X"10",X"DB",X"C9",X"DD",X"21",X"F2",X"4C",X"06",X"04",X"DD",
		X"7E",X"00",X"A7",X"28",X"10",X"DD",X"35",X"00",X"20",X"0B",X"DD",X"6E",X"01",X"DD",X"66",X"02",
		X"36",X"0F",X"23",X"36",X"00",X"11",X"03",X"00",X"DD",X"19",X"10",X"E3",X"C9",X"0F",X"30",X"00",
		X"56",X"43",X"0F",X"30",X"FF",X"01",X"20",X"41",X"15",X"94",X"01",X"32",X"41",X"15",X"94",X"01",
		X"A1",X"41",X"15",X"94",X"01",X"AA",X"41",X"15",X"94",X"01",X"28",X"42",X"15",X"94",X"01",X"35",
		X"42",X"15",X"94",X"01",X"A0",X"42",X"15",X"94",X"01",X"B5",X"42",X"15",X"94",X"00",X"46",X"41",
		X"0F",X"30",X"00",X"49",X"41",X"0F",X"30",X"00",X"50",X"41",X"0F",X"30",X"00",X"55",X"41",X"0F",
		X"30",X"00",X"D8",X"41",X"0F",X"30",X"00",X"44",X"42",X"0F",X"30",X"00",X"4B",X"42",X"0F",X"30",
		X"00",X"C8",X"42",X"0F",X"30",X"FF",X"01",X"21",X"41",X"17",X"90",X"01",X"32",X"41",X"17",X"90",
		X"01",X"26",X"42",X"17",X"90",X"01",X"36",X"42",X"17",X"90",X"01",X"A0",X"42",X"17",X"90",X"01",
		X"B0",X"42",X"17",X"90",X"01",X"21",X"43",X"17",X"90",X"01",X"31",X"43",X"17",X"90",X"00",X"55",
		X"41",X"0F",X"30",X"00",X"58",X"41",X"0F",X"30",X"00",X"55",X"42",X"0F",X"30",X"00",X"44",X"43",
		X"0F",X"30",X"00",X"4A",X"43",X"0F",X"30",X"00",X"4D",X"43",X"0F",X"30",X"00",X"50",X"43",X"0F",
		X"30",X"00",X"53",X"43",X"0F",X"30",X"FF",X"01",X"2B",X"41",X"0F",X"9C",X"01",X"39",X"41",X"0F",
		X"9C",X"01",X"A5",X"41",X"0F",X"9C",X"01",X"AF",X"41",X"0F",X"9C",X"01",X"20",X"42",X"0F",X"9C",
		X"01",X"36",X"42",X"0F",X"9C",X"01",X"A5",X"42",X"0F",X"9C",X"01",X"2B",X"43",X"0F",X"9C",X"00",
		X"54",X"41",X"0F",X"30",X"00",X"57",X"41",X"0F",X"30",X"00",X"44",X"43",X"0F",X"30",X"00",X"47",
		X"43",X"0F",X"30",X"00",X"4A",X"43",X"0F",X"30",X"00",X"4D",X"43",X"0F",X"30",X"00",X"50",X"43",
		X"0F",X"30",X"00",X"53",X"43",X"0F",X"30",X"FF",X"01",X"24",X"41",X"07",X"A0",X"01",X"33",X"41",
		X"07",X"A0",X"01",X"39",X"41",X"07",X"A0",X"01",X"A8",X"41",X"07",X"A0",X"01",X"B9",X"41",X"07",
		X"FF",X"01",X"20",X"42",X"07",X"A0",X"01",X"AE",X"42",X"07",X"A0",X"01",X"24",X"43",X"07",X"A0",
		X"00",X"55",X"41",X"0F",X"30",X"00",X"CA",X"41",X"0F",X"30",X"00",X"43",X"42",X"0F",X"30",X"00",
		X"C7",X"42",X"0F",X"30",X"00",X"4C",X"43",X"0F",X"30",X"00",X"4E",X"43",X"0F",X"30",X"00",X"50",
		X"43",X"0F",X"30",X"00",X"52",X"43",X"0F",X"30",X"FF",X"01",X"25",X"41",X"0F",X"A8",X"01",X"39",
		X"41",X"0F",X"A8",X"01",X"A0",X"41",X"0F",X"A8",X"01",X"B9",X"41",X"0F",X"A8",X"01",X"38",X"42",
		X"0F",X"A8",X"01",X"AB",X"42",X"0F",X"A8",X"01",X"B8",X"42",X"0F",X"A8",X"01",X"22",X"43",X"0F",
		X"A8",X"00",X"C7",X"41",X"0F",X"30",X"00",X"D8",X"41",X"0F",X"30",X"00",X"49",X"42",X"0F",X"30",
		X"00",X"D2",X"42",X"0F",X"30",X"00",X"4C",X"43",X"0F",X"30",X"00",X"4F",X"43",X"0F",X"30",X"00",
		X"53",X"43",X"0F",X"30",X"00",X"56",X"43",X"0F",X"30",X"FF",X"01",X"39",X"41",X"17",X"A4",X"01",
		X"B6",X"41",X"17",X"A4",X"01",X"2E",X"42",X"17",X"A4",X"01",X"39",X"42",X"17",X"A4",X"01",X"A0",
		X"42",X"17",X"A4",X"01",X"B0",X"42",X"17",X"A4",X"01",X"B9",X"42",X"17",X"A4",X"01",X"21",X"43",
		X"17",X"A4",X"00",X"4F",X"41",X"0F",X"30",X"00",X"50",X"41",X"0F",X"30",X"00",X"55",X"41",X"0F",
		X"30",X"00",X"CE",X"41",X"0F",X"30",X"00",X"44",X"43",X"0F",X"30",X"00",X"4C",X"43",X"0F",X"30",
		X"00",X"4F",X"43",X"0F",X"30",X"00",X"51",X"43",X"0F",X"30",X"FF",X"01",X"28",X"41",X"18",X"B4",
		X"01",X"32",X"41",X"18",X"B4",X"01",X"AD",X"41",X"18",X"B4",X"01",X"2B",X"42",X"18",X"B4",X"01",
		X"2E",X"42",X"18",X"B4",X"01",X"A5",X"42",X"18",X"B4",X"01",X"B4",X"42",X"18",X"B4",X"01",X"22",
		X"43",X"18",X"B4",X"00",X"D6",X"41",X"0F",X"30",X"00",X"46",X"43",X"0F",X"30",X"00",X"49",X"43",
		X"0F",X"30",X"00",X"51",X"43",X"0F",X"30",X"00",X"52",X"43",X"0F",X"30",X"00",X"55",X"43",X"0F",
		X"30",X"00",X"58",X"43",X"0F",X"30",X"00",X"59",X"43",X"0F",X"30",X"FF",X"01",X"21",X"41",X"16",
		X"BC",X"01",X"39",X"41",X"16",X"BC",X"01",X"A4",X"41",X"16",X"BC",X"01",X"B8",X"41",X"16",X"BC",
		X"01",X"21",X"42",X"16",X"BC",X"01",X"39",X"42",X"16",X"BC",X"01",X"AD",X"42",X"16",X"BC",X"01",
		X"2D",X"43",X"16",X"BC",X"00",X"C8",X"41",X"0F",X"30",X"00",X"D7",X"41",X"0F",X"30",X"00",X"CC",
		X"42",X"0F",X"30",X"00",X"4B",X"43",X"0F",X"30",X"00",X"4C",X"43",X"0F",X"30",X"00",X"4F",X"43",
		X"0F",X"30",X"00",X"50",X"43",X"0F",X"30",X"00",X"51",X"43",X"0F",X"30",X"FF",X"01",X"21",X"41",
		X"03",X"AC",X"01",X"32",X"41",X"03",X"AC",X"01",X"26",X"42",X"03",X"AC",X"01",X"36",X"42",X"03",
		X"AC",X"01",X"A0",X"42",X"03",X"AC",X"01",X"B0",X"42",X"03",X"AC",X"01",X"21",X"43",X"03",X"AC",
		X"01",X"31",X"43",X"03",X"AC",X"00",X"55",X"41",X"0F",X"30",X"00",X"58",X"41",X"0F",X"30",X"00",
		X"55",X"42",X"0F",X"30",X"00",X"44",X"43",X"0F",X"30",X"00",X"4A",X"43",X"0F",X"30",X"00",X"4D",
		X"43",X"0F",X"30",X"00",X"50",X"43",X"0F",X"30",X"00",X"53",X"43",X"0F",X"30",X"FF",X"01",X"28",
		X"41",X"15",X"B0",X"01",X"31",X"41",X"15",X"B0",X"01",X"B1",X"41",X"15",X"B0",X"01",X"2A",X"42",
		X"15",X"B0",X"01",X"2F",X"42",X"15",X"B0",X"01",X"A5",X"42",X"15",X"B0",X"01",X"B9",X"42",X"15",
		X"B0",X"01",X"21",X"43",X"15",X"B0",X"00",X"C4",X"42",X"0F",X"30",X"00",X"C7",X"42",X"0F",X"30",
		X"FF",X"D3",X"42",X"0F",X"30",X"00",X"D6",X"42",X"0F",X"30",X"00",X"44",X"43",X"0F",X"30",X"00",
		X"47",X"43",X"0F",X"30",X"00",X"4B",X"43",X"0F",X"30",X"00",X"4F",X"43",X"0F",X"30",X"FF",X"01",
		X"2B",X"41",X"17",X"B8",X"01",X"39",X"41",X"17",X"B8",X"01",X"A5",X"41",X"17",X"B8",X"01",X"AF",
		X"41",X"17",X"B8",X"01",X"20",X"42",X"17",X"B8",X"01",X"36",X"42",X"17",X"B8",X"01",X"A5",X"42",
		X"17",X"B8",X"01",X"2B",X"43",X"17",X"B8",X"00",X"54",X"41",X"0F",X"30",X"00",X"57",X"41",X"0F",
		X"30",X"00",X"44",X"43",X"0F",X"30",X"00",X"47",X"43",X"0F",X"30",X"00",X"4A",X"43",X"0F",X"30",
		X"00",X"4D",X"43",X"0F",X"30",X"00",X"50",X"43",X"0F",X"30",X"00",X"53",X"43",X"0F",X"30",X"FF",
		X"2C",X"9D",X"E2",X"9C",X"98",X"9C",X"BD",X"9C",X"07",X"9D",X"76",X"9D",X"51",X"9D",X"9B",X"9D",
		X"C0",X"9D",X"E5",X"9D",X"2F",X"9E",X"0A",X"9E",X"54",X"9E",X"9E",X"9E",X"79",X"9E",X"C0",X"9D",
		X"2F",X"9E",X"C3",X"9E",X"0A",X"9E",X"E8",X"9E",X"08",X"00",X"21",X"43",X"FF",X"40",X"00",X"A8",
		X"42",X"98",X"00",X"B3",X"42",X"FF",X"68",X"00",X"2D",X"42",X"FF",X"00",X"00",X"A0",X"41",X"FF",
		X"00",X"00",X"20",X"41",X"50",X"00",X"2A",X"41",X"78",X"00",X"2F",X"41",X"FF",X"FF",X"50",X"00",
		X"AA",X"42",X"80",X"00",X"B0",X"42",X"FF",X"50",X"00",X"2A",X"42",X"FF",X"18",X"00",X"A3",X"41",
		X"68",X"00",X"AD",X"41",X"90",X"00",X"B2",X"41",X"FF",X"28",X"00",X"25",X"41",X"88",X"00",X"31",
		X"41",X"FF",X"48",X"00",X"29",X"43",X"FF",X"08",X"00",X"A1",X"42",X"C8",X"00",X"B9",X"42",X"FF",
		X"40",X"00",X"28",X"42",X"FF",X"18",X"00",X"A3",X"41",X"58",X"00",X"AB",X"41",X"C8",X"00",X"B9",
		X"41",X"FF",X"08",X"00",X"21",X"41",X"FF",X"78",X"00",X"2F",X"43",X"FF",X"20",X"00",X"A4",X"42",
		X"FF",X"68",X"00",X"2D",X"42",X"C8",X"00",X"39",X"42",X"FF",X"88",X"00",X"B1",X"41",X"FF",X"50",
		X"00",X"2A",X"41",X"78",X"00",X"2F",X"41",X"98",X"00",X"33",X"41",X"FF",X"48",X"00",X"29",X"43",
		X"FF",X"08",X"00",X"A1",X"42",X"C8",X"00",X"B9",X"42",X"FF",X"40",X"00",X"28",X"42",X"C8",X"00",
		X"39",X"42",X"FF",X"C8",X"00",X"B9",X"41",X"FF",X"28",X"00",X"25",X"41",X"A8",X"00",X"35",X"41",
		X"FF",X"20",X"00",X"24",X"43",X"FF",X"58",X"00",X"AB",X"42",X"80",X"00",X"B0",X"42",X"FF",X"A8",
		X"00",X"35",X"42",X"FF",X"28",X"00",X"A5",X"41",X"A8",X"00",X"B5",X"41",X"FF",X"08",X"00",X"21",
		X"41",X"98",X"00",X"33",X"41",X"FF",X"30",X"00",X"26",X"43",X"FF",X"58",X"00",X"AB",X"42",X"C0",
		X"00",X"B8",X"42",X"FF",X"48",X"00",X"29",X"42",X"FF",X"08",X"00",X"A1",X"41",X"B0",X"00",X"B6",
		X"41",X"FF",X"50",X"00",X"2A",X"41",X"A0",X"00",X"34",X"41",X"FF",X"40",X"00",X"28",X"43",X"FF",
		X"08",X"00",X"A1",X"42",X"C8",X"00",X"B9",X"42",X"FF",X"A0",X"00",X"34",X"42",X"FF",X"20",X"00",
		X"A4",X"41",X"78",X"00",X"AF",X"41",X"FF",X"08",X"00",X"21",X"41",X"A8",X"00",X"35",X"41",X"FF",
		X"08",X"00",X"21",X"43",X"88",X"00",X"31",X"43",X"FF",X"00",X"00",X"A0",X"42",X"80",X"00",X"B0",
		X"42",X"FF",X"30",X"00",X"26",X"42",X"B0",X"00",X"36",X"42",X"FF",X"FF",X"08",X"00",X"21",X"41",
		X"90",X"00",X"32",X"41",X"FF",X"FF",X"00",X"00",X"A0",X"42",X"A8",X"00",X"B5",X"42",X"FF",X"40",
		X"00",X"28",X"42",X"A8",X"00",X"35",X"42",X"FF",X"08",X"00",X"A1",X"41",X"50",X"00",X"AA",X"41",
		X"FF",X"00",X"00",X"20",X"41",X"90",X"00",X"32",X"41",X"FF",X"58",X"00",X"2B",X"43",X"FF",X"28",
		X"00",X"A5",X"42",X"FF",X"00",X"00",X"20",X"42",X"B0",X"00",X"36",X"42",X"FF",X"28",X"00",X"A5",
		X"41",X"78",X"00",X"AF",X"41",X"FF",X"58",X"00",X"2B",X"41",X"C8",X"00",X"39",X"41",X"FF",X"08",
		X"00",X"21",X"43",X"FF",X"28",X"00",X"A5",X"42",X"C8",X"00",X"B9",X"42",X"FF",X"50",X"00",X"2A",
		X"42",X"78",X"00",X"2F",X"42",X"FF",X"88",X"00",X"B1",X"41",X"FF",X"40",X"00",X"28",X"41",X"88",
		X"00",X"31",X"41",X"FF",X"20",X"00",X"24",X"43",X"FF",X"70",X"00",X"AE",X"42",X"FF",X"00",X"00",
		X"20",X"42",X"FF",X"40",X"00",X"A8",X"41",X"C8",X"00",X"B9",X"41",X"FF",X"20",X"00",X"24",X"41",
		X"98",X"00",X"33",X"41",X"C8",X"00",X"39",X"41",X"FF",X"10",X"00",X"22",X"43",X"FF",X"58",X"00",
		X"AB",X"42",X"C0",X"00",X"B8",X"42",X"FF",X"C0",X"00",X"38",X"42",X"FF",X"00",X"00",X"A0",X"41",
		X"C8",X"00",X"B9",X"41",X"FF",X"28",X"00",X"25",X"41",X"C8",X"00",X"39",X"41",X"FF",X"08",X"00",
		X"21",X"43",X"FF",X"00",X"00",X"A0",X"42",X"80",X"00",X"B0",X"42",X"C8",X"00",X"B9",X"42",X"FF",
		X"70",X"00",X"2E",X"42",X"C8",X"00",X"39",X"42",X"FF",X"B0",X"00",X"B6",X"41",X"FF",X"C8",X"00",
		X"39",X"41",X"FF",X"10",X"00",X"22",X"43",X"FF",X"28",X"00",X"A5",X"42",X"A0",X"00",X"B4",X"42",
		X"FF",X"58",X"00",X"2B",X"42",X"70",X"00",X"2E",X"42",X"FF",X"68",X"00",X"AD",X"41",X"FF",X"40",
		X"00",X"28",X"41",X"90",X"00",X"32",X"41",X"FF",X"68",X"00",X"2D",X"43",X"FF",X"68",X"00",X"AD",
		X"42",X"FF",X"08",X"00",X"21",X"42",X"C8",X"00",X"39",X"42",X"FF",X"20",X"00",X"A4",X"41",X"C0",
		X"00",X"B8",X"41",X"FF",X"08",X"00",X"21",X"41",X"C8",X"00",X"39",X"41",X"FF",X"89",X"9F",X"5F",
		X"9F",X"35",X"9F",X"4A",X"9F",X"74",X"9F",X"B3",X"9F",X"9E",X"9F",X"C8",X"9F",X"DD",X"9F",X"F2",
		X"9F",X"1C",X"A0",X"07",X"A0",X"31",X"A0",X"5B",X"A0",X"46",X"A0",X"DD",X"9F",X"1C",X"A0",X"70",
		X"A0",X"07",X"A0",X"85",X"A0",X"FF",X"07",X"33",X"08",X"4C",X"FF",X"27",X"43",X"06",X"4C",X"FF",
		X"8F",X"02",X"04",X"4C",X"FF",X"8F",X"53",X"02",X"4C",X"FF",X"67",X"02",X"08",X"4C",X"FF",X"FF",
		X"87",X"02",X"06",X"4C",X"FF",X"40",X"63",X"04",X"4C",X"FF",X"AF",X"02",X"02",X"4C",X"FF",X"FF",
		X"3F",X"02",X"08",X"4C",X"FF",X"C7",X"53",X"06",X"4C",X"FF",X"08",X"63",X"04",X"4C",X"FF",X"97",
		X"02",X"02",X"4C",X"FF",X"FF",X"87",X"02",X"08",X"4C",X"FF",X"4F",X"33",X"06",X"4C",X"FF",X"3F",
		X"02",X"04",X"4C",X"FF",X"C7",X"43",X"02",X"4C",X"FF",X"FF",X"8F",X"02",X"08",X"4C",X"FF",X"FF",
		X"07",X"53",X"06",X"4C",X"FF",X"87",X"02",X"04",X"4C",X"07",X"63",X"02",X"4C",X"FF",X"FF",X"27",
		X"02",X"08",X"4C",X"CF",X"33",X"06",X"4C",X"FF",X"27",X"43",X"04",X"4C",X"FF",X"5F",X"02",X"02",
		X"4C",X"FF",X"FF",X"FF",X"2F",X"43",X"08",X"4C",X"FF",X"97",X"02",X"06",X"4C",X"FF",X"3F",X"53",
		X"04",X"4C",X"FF",X"B7",X"02",X"02",X"4C",X"FF",X"97",X"02",X"08",X"4C",X"FF",X"6F",X"02",X"06",
		X"4C",X"FF",X"B7",X"33",X"04",X"4C",X"FF",X"97",X"43",X"02",X"4C",X"FF",X"FF",X"FF",X"27",X"43",
		X"08",X"4C",X"B7",X"02",X"06",X"4C",X"FF",X"FF",X"27",X"33",X"04",X"4C",X"AF",X"63",X"02",X"4C",
		X"FF",X"FF",X"FF",X"4F",X"02",X"08",X"4C",X"FF",X"77",X"63",X"06",X"4C",X"FF",X"8F",X"33",X"04");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
