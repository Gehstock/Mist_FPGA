library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity basic is
    generic(
        AddrWidth   : integer := 14
    );
    port (
        clk  : in std_logic;
        addr : in std_logic_vector(AddrWidth-1 downto 0);
        data : out std_logic_vector(7 downto 0)
    );
end basic;

architecture rtl of basic is
    signal romAddr : integer range 0 to 2**AddrWidth-1;
    type rom16384x8 is array (0 to 2**AddrWidth-1) of std_logic_vector(7 downto 0); 
    constant romData : rom16384x8 := (
         x"18",  x"0b",  x"c3",  x"8c",  x"c0",  x"7f",  x"7f",  x"42", -- 0000
         x"41",  x"53",  x"49",  x"43",  x"00",  x"21",  x"bd",  x"c0", -- 0008
         x"11",  x"00",  x"03",  x"01",  x"67",  x"00",  x"ed",  x"b0", -- 0010
         x"eb",  x"f9",  x"cd",  x"69",  x"c6",  x"32",  x"ab",  x"03", -- 0018
         x"32",  x"00",  x"04",  x"21",  x"92",  x"c0",  x"cd",  x"c9", -- 0020
         x"d1",  x"21",  x"ae",  x"c0",  x"cd",  x"c9",  x"d1",  x"cd", -- 0028
         x"ae",  x"c5",  x"21",  x"62",  x"03",  x"cd",  x"86",  x"c9", -- 0030
         x"7a",  x"d6",  x"06",  x"21",  x"00",  x"03",  x"2b",  x"30", -- 0038
         x"03",  x"11",  x"ff",  x"bf",  x"23",  x"cd",  x"89",  x"c6", -- 0040
         x"28",  x"09",  x"7e",  x"47",  x"2f",  x"77",  x"be",  x"70", -- 0048
         x"28",  x"f2",  x"2b",  x"11",  x"00",  x"ff",  x"22",  x"b0", -- 0050
         x"03",  x"19",  x"22",  x"56",  x"03",  x"cd",  x"41",  x"c6", -- 0058
         x"2a",  x"56",  x"03",  x"11",  x"ef",  x"fb",  x"19",  x"cd", -- 0060
         x"29",  x"d8",  x"21",  x"a0",  x"c0",  x"cd",  x"c9",  x"d1", -- 0068
         x"2a",  x"04",  x"e0",  x"7e",  x"fe",  x"78",  x"20",  x"01", -- 0070
         x"3e",  x"af",  x"32",  x"fc",  x"03",  x"31",  x"67",  x"03", -- 0078
         x"18",  x"0a",  x"7f",  x"7f",  x"52",  x"45",  x"42",  x"41", -- 0080
         x"53",  x"49",  x"43",  x"00",  x"cd",  x"69",  x"c6",  x"c3", -- 0088
         x"88",  x"c3",  x"0c",  x"0a",  x"0d",  x"48",  x"43",  x"2d", -- 0090
         x"42",  x"41",  x"53",  x"49",  x"43",  x"0a",  x"0d",  x"00", -- 0098
         x"20",  x"42",  x"59",  x"54",  x"45",  x"53",  x"20",  x"46", -- 00A0
         x"52",  x"45",  x"45",  x"0a",  x"0d",  x"00",  x"4d",  x"45", -- 00A8
         x"4d",  x"4f",  x"52",  x"59",  x"20",  x"45",  x"4e",  x"44", -- 00B0
         x"20",  x"3f",  x"20",  x"3a",  x"00",  x"c3",  x"89",  x"c0", -- 00B8
         x"c3",  x"67",  x"c9",  x"00",  x"00",  x"00",  x"00",  x"00", -- 00C0
         x"d6",  x"00",  x"6f",  x"7c",  x"de",  x"00",  x"67",  x"78", -- 00C8
         x"de",  x"00",  x"47",  x"3e",  x"00",  x"c9",  x"00",  x"00", -- 00D0
         x"00",  x"35",  x"4a",  x"ca",  x"99",  x"39",  x"1c",  x"76", -- 00D8
         x"98",  x"22",  x"95",  x"b3",  x"98",  x"0a",  x"dd",  x"47", -- 00E0
         x"98",  x"53",  x"d1",  x"99",  x"99",  x"0a",  x"1a",  x"9f", -- 00E8
         x"98",  x"65",  x"bc",  x"cd",  x"98",  x"d6",  x"77",  x"3e", -- 00F0
         x"98",  x"52",  x"c7",  x"4f",  x"80",  x"0b",  x"ff",  x"1b", -- 00F8
         x"00",  x"0a",  x"00",  x"0a",  x"00",  x"00",  x"00",  x"c3", -- 0100
         x"ae",  x"c5",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0108
         x"00",  x"00",  x"00",  x"65",  x"04",  x"fe",  x"ff",  x"00", -- 0110
         x"00",  x"c9",  x"00",  x"00",  x"01",  x"04",  x"00",  x"00", -- 0118
         x"00",  x"c5",  x"4e",  x"44",  x"c6",  x"4f",  x"52",  x"ce", -- 0120
         x"45",  x"58",  x"54",  x"c4",  x"41",  x"54",  x"41",  x"c9", -- 0128
         x"4e",  x"50",  x"55",  x"54",  x"c4",  x"49",  x"4d",  x"d2", -- 0130
         x"45",  x"41",  x"44",  x"cc",  x"45",  x"54",  x"c7",  x"4f", -- 0138
         x"54",  x"4f",  x"d2",  x"55",  x"4e",  x"c9",  x"46",  x"d2", -- 0140
         x"45",  x"53",  x"54",  x"4f",  x"52",  x"45",  x"c7",  x"4f", -- 0148
         x"53",  x"55",  x"42",  x"d2",  x"45",  x"54",  x"55",  x"52", -- 0150
         x"4e",  x"d2",  x"45",  x"4d",  x"d3",  x"54",  x"4f",  x"50", -- 0158
         x"cf",  x"55",  x"54",  x"cf",  x"4e",  x"ce",  x"55",  x"4c", -- 0160
         x"4c",  x"d7",  x"41",  x"49",  x"54",  x"c4",  x"45",  x"46", -- 0168
         x"d0",  x"4f",  x"4b",  x"45",  x"c4",  x"4f",  x"4b",  x"45", -- 0170
         x"c1",  x"55",  x"54",  x"4f",  x"cc",  x"49",  x"4e",  x"45", -- 0178
         x"53",  x"c3",  x"4c",  x"53",  x"d7",  x"49",  x"44",  x"54", -- 0180
         x"48",  x"c2",  x"59",  x"45",  x"a1",  x"c3",  x"41",  x"4c", -- 0188
         x"4c",  x"d0",  x"52",  x"49",  x"4e",  x"54",  x"c3",  x"4f", -- 0190
         x"4e",  x"54",  x"cc",  x"49",  x"53",  x"54",  x"c3",  x"4c", -- 0198
         x"45",  x"41",  x"52",  x"c3",  x"4c",  x"4f",  x"41",  x"44", -- 01A0
         x"c3",  x"53",  x"41",  x"56",  x"45",  x"ce",  x"45",  x"57", -- 01A8
         x"d4",  x"41",  x"42",  x"28",  x"d4",  x"4f",  x"c6",  x"4e", -- 01B0
         x"d3",  x"50",  x"43",  x"28",  x"d4",  x"48",  x"45",  x"4e", -- 01B8
         x"ce",  x"4f",  x"54",  x"d3",  x"54",  x"45",  x"50",  x"ab", -- 01C0
         x"ad",  x"aa",  x"af",  x"de",  x"c1",  x"4e",  x"44",  x"cf", -- 01C8
         x"52",  x"be",  x"bd",  x"bc",  x"d3",  x"47",  x"4e",  x"c9", -- 01D0
         x"4e",  x"54",  x"c1",  x"42",  x"53",  x"d5",  x"53",  x"52", -- 01D8
         x"c6",  x"52",  x"45",  x"c9",  x"4e",  x"50",  x"d0",  x"4f", -- 01E0
         x"53",  x"d3",  x"51",  x"52",  x"d2",  x"4e",  x"44",  x"cc", -- 01E8
         x"4e",  x"c5",  x"58",  x"50",  x"c3",  x"4f",  x"53",  x"d3", -- 01F0
         x"49",  x"4e",  x"d4",  x"41",  x"4e",  x"c1",  x"54",  x"4e", -- 01F8
         x"d0",  x"45",  x"45",  x"4b",  x"c4",  x"45",  x"45",  x"4b", -- 0200
         x"d0",  x"49",  x"cc",  x"45",  x"4e",  x"d3",  x"54",  x"52", -- 0208
         x"24",  x"d6",  x"41",  x"4c",  x"c1",  x"53",  x"43",  x"c3", -- 0210
         x"48",  x"52",  x"24",  x"cc",  x"45",  x"46",  x"54",  x"24", -- 0218
         x"d2",  x"49",  x"47",  x"48",  x"54",  x"24",  x"cd",  x"49", -- 0220
         x"44",  x"24",  x"cc",  x"4f",  x"41",  x"44",  x"d4",  x"52", -- 0228
         x"4f",  x"4e",  x"d4",  x"52",  x"4f",  x"46",  x"46",  x"c5", -- 0230
         x"44",  x"49",  x"54",  x"c5",  x"4c",  x"53",  x"45",  x"80", -- 0238
         x"1a",  x"c9",  x"de",  x"c7",  x"dc",  x"cc",  x"48",  x"ca", -- 0240
         x"ec",  x"cb",  x"01",  x"cf",  x"1f",  x"cc",  x"5d",  x"ca", -- 0248
         x"07",  x"ca",  x"eb",  x"c9",  x"cf",  x"ca",  x"df",  x"c8", -- 0250
         x"f6",  x"c9",  x"25",  x"ca",  x"4a",  x"ca",  x"18",  x"c9", -- 0258
         x"ec",  x"d3",  x"b3",  x"ca",  x"c0",  x"cb",  x"f7",  x"d3", -- 0260
         x"c4",  x"d0",  x"37",  x"d4",  x"4e",  x"d4",  x"fa",  x"c5", -- 0268
         x"ea",  x"c6",  x"d0",  x"dd",  x"b9",  x"cb",  x"f4",  x"df", -- 0270
         x"4a",  x"ca",  x"38",  x"db",  x"fa",  x"ca",  x"48",  x"c9", -- 0278
         x"f2",  x"c6",  x"aa",  x"c9",  x"43",  x"dc",  x"41",  x"dd", -- 0280
         x"40",  x"c6",  x"2d",  x"c6",  x"b7",  x"c7",  x"b8",  x"c7", -- 0288
         x"e7",  x"c3",  x"4a",  x"ca",  x"a6",  x"d6",  x"70",  x"d7", -- 0290
         x"bc",  x"d6",  x"03",  x"03",  x"90",  x"d0",  x"e3",  x"d3", -- 0298
         x"bd",  x"d0",  x"1f",  x"d9",  x"fd",  x"d9",  x"59",  x"d5", -- 02A0
         x"6d",  x"d9",  x"70",  x"da",  x"76",  x"da",  x"d7",  x"da", -- 02A8
         x"ec",  x"da",  x"31",  x"d4",  x"44",  x"d4",  x"d5",  x"d6", -- 02B0
         x"2c",  x"d3",  x"56",  x"d1",  x"bf",  x"d3",  x"3b",  x"d3", -- 02B8
         x"4b",  x"d3",  x"5b",  x"d3",  x"89",  x"d3",  x"92",  x"d3", -- 02C0
         x"79",  x"11",  x"d8",  x"79",  x"6a",  x"d4",  x"7c",  x"98", -- 02C8
         x"d5",  x"7c",  x"f3",  x"d5",  x"7f",  x"28",  x"d9",  x"50", -- 02D0
         x"5e",  x"ce",  x"46",  x"5d",  x"ce",  x"4e",  x"46",  x"53", -- 02D8
         x"4e",  x"52",  x"47",  x"4f",  x"44",  x"46",  x"43",  x"4f", -- 02E0
         x"56",  x"4f",  x"4d",  x"55",  x"4c",  x"42",  x"53",  x"44", -- 02E8
         x"44",  x"2f",  x"30",  x"49",  x"44",  x"54",  x"4d",  x"4f", -- 02F0
         x"53",  x"4c",  x"53",  x"53",  x"54",  x"43",  x"4e",  x"55", -- 02F8
         x"46",  x"4d",  x"4f",  x"49",  x"4f",  x"20",  x"45",  x"52", -- 0300
         x"52",  x"4f",  x"52",  x"07",  x"00",  x"20",  x"49",  x"4e", -- 0308
         x"20",  x"00",  x"46",  x"49",  x"4c",  x"45",  x"20",  x"46", -- 0310
         x"4f",  x"55",  x"4e",  x"44",  x"0d",  x"4f",  x"4b",  x"0d", -- 0318
         x"00",  x"42",  x"52",  x"45",  x"41",  x"4b",  x"00",  x"e5", -- 0320
         x"2a",  x"db",  x"03",  x"06",  x"00",  x"09",  x"09",  x"3e", -- 0328
         x"e5",  x"3e",  x"d0",  x"95",  x"6f",  x"3e",  x"ff",  x"9c", -- 0330
         x"38",  x"04",  x"67",  x"39",  x"e1",  x"d8",  x"1e",  x"0c", -- 0338
         x"18",  x"14",  x"2a",  x"ca",  x"03",  x"22",  x"58",  x"03", -- 0340
         x"1e",  x"02",  x"01",  x"1e",  x"14",  x"01",  x"1e",  x"00", -- 0348
         x"01",  x"1e",  x"12",  x"01",  x"1e",  x"22",  x"cd",  x"69", -- 0350
         x"c6",  x"32",  x"43",  x"03",  x"cd",  x"55",  x"cb",  x"21", -- 0358
         x"dd",  x"c2",  x"57",  x"19",  x"44",  x"4d",  x"0b",  x"3e", -- 0360
         x"3f",  x"1e",  x"03",  x"cd",  x"d6",  x"d1",  x"21",  x"05", -- 0368
         x"c3",  x"cd",  x"c9",  x"d1",  x"2a",  x"58",  x"03",  x"11", -- 0370
         x"fe",  x"ff",  x"cd",  x"89",  x"c6",  x"ca",  x"0d",  x"c0", -- 0378
         x"7c",  x"a5",  x"3c",  x"c4",  x"21",  x"d8",  x"3e",  x"c1", -- 0380
         x"af",  x"32",  x"43",  x"03",  x"cd",  x"55",  x"cb",  x"21", -- 0388
         x"1d",  x"c3",  x"cd",  x"c9",  x"d1",  x"37",  x"dc",  x"fd", -- 0390
         x"dd",  x"cd",  x"df",  x"c6",  x"2b",  x"22",  x"58",  x"03", -- 0398
         x"21",  x"ea",  x"03",  x"3a",  x"4d",  x"03",  x"b7",  x"28", -- 03A0
         x"6b",  x"ed",  x"5b",  x"4e",  x"03",  x"f2",  x"f0",  x"c3", -- 03A8
         x"d5",  x"cd",  x"2a",  x"d8",  x"d1",  x"d5",  x"cd",  x"bb", -- 03B0
         x"c4",  x"3e",  x"2a",  x"38",  x"02",  x"3e",  x"20",  x"cd", -- 03B8
         x"ae",  x"c6",  x"cd",  x"ae",  x"c5",  x"d1",  x"30",  x"06", -- 03C0
         x"af",  x"32",  x"4d",  x"03",  x"18",  x"ba",  x"2a",  x"50", -- 03C8
         x"03",  x"19",  x"38",  x"f4",  x"d5",  x"11",  x"f9",  x"ff", -- 03D0
         x"cd",  x"89",  x"c6",  x"d1",  x"30",  x"ea",  x"22",  x"4e", -- 03D8
         x"03",  x"21",  x"62",  x"03",  x"f5",  x"18",  x"47",  x"c8", -- 03E0
         x"cd",  x"97",  x"c6",  x"cd",  x"86",  x"c9",  x"c0",  x"c1", -- 03E8
         x"cd",  x"bb",  x"c4",  x"30",  x"58",  x"d5",  x"7e",  x"23", -- 03F0
         x"b6",  x"23",  x"28",  x"02",  x"3e",  x"7f",  x"32",  x"4d", -- 03F8
         x"03",  x"7e",  x"23",  x"66",  x"6f",  x"22",  x"4e",  x"03", -- 0400
         x"cd",  x"98",  x"de",  x"d1",  x"c2",  x"96",  x"c3",  x"38", -- 0408
         x"b7",  x"3f",  x"18",  x"cd",  x"3e",  x"3e",  x"cd",  x"ae", -- 0410
         x"c6",  x"cd",  x"ae",  x"c5",  x"da",  x"96",  x"c3",  x"21", -- 0418
         x"61",  x"03",  x"cd",  x"bd",  x"c8",  x"3c",  x"3d",  x"ca", -- 0420
         x"96",  x"c3",  x"f5",  x"cd",  x"86",  x"c9",  x"d5",  x"cd", -- 0428
         x"da",  x"c4",  x"47",  x"d1",  x"f1",  x"d2",  x"8a",  x"c8", -- 0430
         x"d5",  x"c5",  x"af",  x"32",  x"cd",  x"03",  x"cd",  x"bd", -- 0438
         x"c8",  x"b7",  x"f5",  x"cd",  x"bb",  x"c4",  x"38",  x"08", -- 0440
         x"f1",  x"f5",  x"b7",  x"20",  x"03",  x"c3",  x"20",  x"ca", -- 0448
         x"c5",  x"30",  x"11",  x"eb",  x"2a",  x"d7",  x"03",  x"1a", -- 0450
         x"02",  x"03",  x"13",  x"cd",  x"89",  x"c6",  x"20",  x"f7", -- 0458
         x"ed",  x"43",  x"d7",  x"03",  x"d1",  x"f1",  x"28",  x"22", -- 0460
         x"2a",  x"d7",  x"03",  x"e3",  x"c1",  x"09",  x"e5",  x"cd", -- 0468
         x"ab",  x"c4",  x"e1",  x"22",  x"d7",  x"03",  x"eb",  x"36", -- 0470
         x"ff",  x"d1",  x"23",  x"23",  x"73",  x"23",  x"72",  x"23", -- 0478
         x"11",  x"62",  x"03",  x"1a",  x"77",  x"23",  x"13",  x"b7", -- 0480
         x"20",  x"f9",  x"cd",  x"4f",  x"c6",  x"23",  x"eb",  x"21", -- 0488
         x"96",  x"c3",  x"e5",  x"62",  x"6b",  x"7e",  x"23",  x"b6", -- 0490
         x"c8",  x"23",  x"7e",  x"23",  x"a6",  x"3c",  x"c8",  x"23", -- 0498
         x"af",  x"be",  x"23",  x"20",  x"fc",  x"eb",  x"73",  x"23", -- 04A0
         x"72",  x"18",  x"e8",  x"cd",  x"30",  x"c3",  x"c5",  x"e3", -- 04A8
         x"c1",  x"cd",  x"89",  x"c6",  x"7e",  x"02",  x"c8",  x"0b", -- 04B0
         x"2b",  x"18",  x"f6",  x"2a",  x"5f",  x"03",  x"44",  x"4d", -- 04B8
         x"7e",  x"23",  x"b6",  x"2b",  x"c8",  x"23",  x"23",  x"7e", -- 04C0
         x"23",  x"66",  x"6f",  x"cd",  x"89",  x"c6",  x"60",  x"69", -- 04C8
         x"7e",  x"23",  x"66",  x"6f",  x"3f",  x"c8",  x"3f",  x"d0", -- 04D0
         x"18",  x"e4",  x"af",  x"32",  x"af",  x"03",  x"0e",  x"05", -- 04D8
         x"11",  x"62",  x"03",  x"af",  x"32",  x"fb",  x"03",  x"7e", -- 04E0
         x"fe",  x"20",  x"ca",  x"71",  x"c5",  x"47",  x"fe",  x"22", -- 04E8
         x"ca",  x"91",  x"c5",  x"b7",  x"ca",  x"97",  x"c5",  x"3a", -- 04F0
         x"af",  x"03",  x"b7",  x"7e",  x"20",  x"73",  x"fe",  x"3f", -- 04F8
         x"3e",  x"9e",  x"28",  x"6d",  x"7e",  x"fe",  x"30",  x"38", -- 0500
         x"04",  x"fe",  x"3c",  x"38",  x"64",  x"d5",  x"11",  x"20", -- 0508
         x"c1",  x"c5",  x"01",  x"6d",  x"c5",  x"c5",  x"06",  x"7f", -- 0510
         x"7e",  x"fe",  x"61",  x"38",  x"07",  x"fe",  x"7b",  x"30", -- 0518
         x"03",  x"e6",  x"5f",  x"77",  x"4e",  x"eb",  x"23",  x"b6", -- 0520
         x"f2",  x"26",  x"c5",  x"04",  x"7e",  x"e6",  x"7f",  x"20", -- 0528
         x"15",  x"3a",  x"fc",  x"03",  x"a7",  x"c8",  x"3a",  x"fb", -- 0530
         x"03",  x"a7",  x"c0",  x"3c",  x"32",  x"fb",  x"03",  x"2a", -- 0538
         x"0c",  x"e0",  x"7e",  x"e6",  x"7f",  x"c8",  x"b9",  x"20", -- 0540
         x"dd",  x"eb",  x"e5",  x"13",  x"1a",  x"b7",  x"fa",  x"69", -- 0548
         x"c5",  x"4f",  x"78",  x"fe",  x"88",  x"20",  x"04",  x"cd", -- 0550
         x"bd",  x"c8",  x"2b",  x"23",  x"7e",  x"fe",  x"61",  x"38", -- 0558
         x"02",  x"e6",  x"5f",  x"b9",  x"28",  x"e5",  x"e1",  x"18", -- 0560
         x"bb",  x"48",  x"f1",  x"eb",  x"c9",  x"eb",  x"79",  x"c1", -- 0568
         x"d1",  x"23",  x"12",  x"13",  x"0c",  x"d6",  x"3a",  x"28", -- 0570
         x"04",  x"fe",  x"49",  x"20",  x"03",  x"32",  x"af",  x"03", -- 0578
         x"d6",  x"54",  x"28",  x"05",  x"d6",  x"0e",  x"c2",  x"e3", -- 0580
         x"c4",  x"47",  x"7e",  x"b7",  x"28",  x"09",  x"b8",  x"28", -- 0588
         x"e0",  x"23",  x"12",  x"0c",  x"13",  x"18",  x"f3",  x"21", -- 0590
         x"61",  x"03",  x"12",  x"13",  x"12",  x"13",  x"12",  x"c9", -- 0598
         x"4c",  x"49",  x"53",  x"54",  x"00",  x"52",  x"55",  x"4e", -- 05A0
         x"00",  x"43",  x"4f",  x"4e",  x"54",  x"00",  x"e5",  x"21", -- 05A8
         x"62",  x"03",  x"e3",  x"cd",  x"e4",  x"dd",  x"e3",  x"fe", -- 05B0
         x"1c",  x"11",  x"9f",  x"c5",  x"28",  x"0e",  x"fe",  x"1d", -- 05B8
         x"11",  x"a4",  x"c5",  x"28",  x"07",  x"fe",  x"1e",  x"11", -- 05C0
         x"a8",  x"c5",  x"20",  x"14",  x"21",  x"61",  x"03",  x"23", -- 05C8
         x"13",  x"1a",  x"77",  x"a7",  x"20",  x"f9",  x"21",  x"62", -- 05D0
         x"03",  x"cd",  x"f1",  x"c5",  x"e1",  x"c3",  x"5e",  x"cb", -- 05D8
         x"cd",  x"0f",  x"df",  x"20",  x"02",  x"e1",  x"c9",  x"cd", -- 05E0
         x"27",  x"df",  x"38",  x"f9",  x"cd",  x"32",  x"df",  x"18", -- 05E8
         x"c1",  x"7e",  x"b7",  x"c8",  x"cd",  x"d5",  x"dd",  x"23", -- 05F0
         x"18",  x"f7",  x"11",  x"0a",  x"00",  x"d5",  x"28",  x"17", -- 05F8
         x"cd",  x"86",  x"c9",  x"eb",  x"e3",  x"28",  x"11",  x"eb", -- 0600
         x"cd",  x"d6",  x"c8",  x"ed",  x"5b",  x"50",  x"03",  x"28", -- 0608
         x"06",  x"cd",  x"86",  x"c9",  x"c2",  x"48",  x"c3",  x"eb", -- 0610
         x"7d",  x"b4",  x"ca",  x"67",  x"c9",  x"22",  x"50",  x"03", -- 0618
         x"cb",  x"ff",  x"32",  x"4d",  x"03",  x"e1",  x"22",  x"4e", -- 0620
         x"03",  x"c1",  x"c3",  x"96",  x"c3",  x"cd",  x"5f",  x"de", -- 0628
         x"3a",  x"09",  x"03",  x"e6",  x"03",  x"28",  x"f3",  x"3e", -- 0630
         x"d5",  x"cd",  x"b2",  x"dc",  x"f1",  x"af",  x"18",  x"ea", -- 0638
         x"c0",  x"2a",  x"5f",  x"03",  x"af",  x"32",  x"5e",  x"03", -- 0640
         x"77",  x"23",  x"77",  x"23",  x"22",  x"d7",  x"03",  x"2a", -- 0648
         x"5f",  x"03",  x"2b",  x"22",  x"cf",  x"03",  x"2a",  x"b0", -- 0650
         x"03",  x"22",  x"c4",  x"03",  x"af",  x"cd",  x"df",  x"c8", -- 0658
         x"2a",  x"d7",  x"03",  x"22",  x"d9",  x"03",  x"22",  x"db", -- 0660
         x"03",  x"c1",  x"2a",  x"56",  x"03",  x"f9",  x"21",  x"b4", -- 0668
         x"03",  x"22",  x"b2",  x"03",  x"cd",  x"1d",  x"de",  x"af", -- 0670
         x"6f",  x"67",  x"22",  x"d5",  x"03",  x"32",  x"cc",  x"03", -- 0678
         x"22",  x"df",  x"03",  x"e5",  x"c5",  x"2a",  x"cf",  x"03", -- 0680
         x"c9",  x"7c",  x"92",  x"c0",  x"7d",  x"93",  x"c9",  x"7e", -- 0688
         x"fe",  x"41",  x"d8",  x"fe",  x"5b",  x"3f",  x"c9",  x"3a", -- 0690
         x"5e",  x"03",  x"a7",  x"c8",  x"cd",  x"69",  x"c6",  x"c3", -- 0698
         x"6e",  x"c3",  x"cd",  x"89",  x"c6",  x"3e",  x"08",  x"18", -- 06A0
         x"02",  x"3e",  x"20",  x"c3",  x"d5",  x"dd",  x"f5",  x"c5", -- 06A8
         x"4f",  x"fe",  x"20",  x"38",  x"13",  x"3a",  x"41",  x"03", -- 06B0
         x"47",  x"3a",  x"ac",  x"03",  x"04",  x"28",  x"05",  x"05", -- 06B8
         x"b8",  x"cc",  x"61",  x"cb",  x"3c",  x"32",  x"ac",  x"03", -- 06C0
         x"79",  x"cd",  x"d5",  x"dd",  x"c1",  x"f1",  x"c9",  x"3e", -- 06C8
         x"3f",  x"cd",  x"ae",  x"c6",  x"3e",  x"09",  x"cd",  x"ae", -- 06D0
         x"c6",  x"cd",  x"df",  x"c6",  x"c3",  x"4a",  x"03",  x"21", -- 06D8
         x"00",  x"20",  x"22",  x"61",  x"03",  x"22",  x"63",  x"03", -- 06E0
         x"65",  x"c9",  x"cd",  x"6c",  x"c9",  x"ed",  x"53",  x"46", -- 06E8
         x"03",  x"c9",  x"cd",  x"97",  x"c6",  x"cd",  x"25",  x"de", -- 06F0
         x"cd",  x"c8",  x"dd",  x"28",  x"12",  x"3e",  x"d5",  x"cd", -- 06F8
         x"b2",  x"dc",  x"2a",  x"46",  x"03",  x"22",  x"4e",  x"03", -- 0700
         x"21",  x"ff",  x"ff",  x"22",  x"46",  x"03",  x"e1",  x"cd", -- 0708
         x"86",  x"c9",  x"c0",  x"c1",  x"cd",  x"bb",  x"c4",  x"c5", -- 0710
         x"cd",  x"91",  x"c7",  x"e1",  x"4e",  x"23",  x"46",  x"23", -- 0718
         x"78",  x"b1",  x"28",  x"59",  x"cd",  x"67",  x"c7",  x"cd", -- 0720
         x"f9",  x"c8",  x"c5",  x"5e",  x"23",  x"56",  x"23",  x"e5", -- 0728
         x"21",  x"ea",  x"03",  x"cd",  x"61",  x"cb",  x"cd",  x"2a", -- 0730
         x"d8",  x"3e",  x"20",  x"e1",  x"cd",  x"ae",  x"c6",  x"7e", -- 0738
         x"23",  x"fe",  x"22",  x"28",  x"14",  x"b7",  x"28",  x"d3", -- 0740
         x"f2",  x"3c",  x"c7",  x"cd",  x"9a",  x"c7",  x"cd",  x"ae", -- 0748
         x"c6",  x"1a",  x"13",  x"b7",  x"f2",  x"4e",  x"c7",  x"18", -- 0750
         x"e6",  x"cd",  x"ae",  x"c6",  x"7e",  x"23",  x"b7",  x"28", -- 0758
         x"ba",  x"fe",  x"22",  x"28",  x"d7",  x"18",  x"f2",  x"e5", -- 0760
         x"2a",  x"44",  x"03",  x"7d",  x"b4",  x"2b",  x"22",  x"44", -- 0768
         x"03",  x"e1",  x"c0",  x"cd",  x"91",  x"c7",  x"cd",  x"e4", -- 0770
         x"dd",  x"fe",  x"03",  x"20",  x"ea",  x"cd",  x"c8",  x"dd", -- 0778
         x"28",  x"0c",  x"cd",  x"61",  x"cb",  x"cd",  x"fd",  x"dd", -- 0780
         x"2a",  x"4e",  x"03",  x"22",  x"46",  x"03",  x"c3",  x"8c", -- 0788
         x"c0",  x"e5",  x"2a",  x"46",  x"03",  x"22",  x"44",  x"03", -- 0790
         x"e1",  x"c9",  x"d6",  x"7f",  x"fe",  x"56",  x"38",  x"08", -- 0798
         x"d6",  x"55",  x"ed",  x"5b",  x"0c",  x"e0",  x"18",  x"03", -- 07A0
         x"11",  x"21",  x"c1",  x"47",  x"1a",  x"13",  x"b7",  x"f2", -- 07A8
         x"ac",  x"c7",  x"10",  x"f8",  x"e6",  x"7f",  x"c9",  x"3e", -- 07B0
         x"af",  x"32",  x"0a",  x"03",  x"c9",  x"21",  x"04",  x"00", -- 07B8
         x"39",  x"7e",  x"23",  x"fe",  x"81",  x"c0",  x"4e",  x"23", -- 07C0
         x"46",  x"23",  x"e5",  x"69",  x"60",  x"7a",  x"b3",  x"eb", -- 07C8
         x"28",  x"04",  x"eb",  x"cd",  x"89",  x"c6",  x"01",  x"0d", -- 07D0
         x"00",  x"e1",  x"c8",  x"09",  x"18",  x"e3",  x"3e",  x"64", -- 07D8
         x"32",  x"cc",  x"03",  x"cd",  x"5d",  x"ca",  x"c1",  x"e5", -- 07E0
         x"cd",  x"48",  x"ca",  x"22",  x"c8",  x"03",  x"21",  x"02", -- 07E8
         x"00",  x"39",  x"cd",  x"c1",  x"c7",  x"d1",  x"20",  x"14", -- 07F0
         x"09",  x"d5",  x"2b",  x"56",  x"2b",  x"5e",  x"23",  x"23", -- 07F8
         x"e5",  x"2a",  x"c8",  x"03",  x"cd",  x"89",  x"c6",  x"e1", -- 0800
         x"20",  x"e8",  x"d1",  x"f9",  x"eb",  x"0e",  x"08",  x"cd", -- 0808
         x"27",  x"c3",  x"e5",  x"2a",  x"c8",  x"03",  x"e3",  x"e5", -- 0810
         x"2a",  x"58",  x"03",  x"e3",  x"cd",  x"29",  x"cd",  x"cd", -- 0818
         x"cc",  x"c8",  x"a6",  x"cd",  x"26",  x"cd",  x"e5",  x"cd", -- 0820
         x"eb",  x"d6",  x"e1",  x"c5",  x"d5",  x"01",  x"00",  x"81", -- 0828
         x"51",  x"5a",  x"7e",  x"fe",  x"ab",  x"3e",  x"01",  x"20", -- 0830
         x"0e",  x"cd",  x"bd",  x"c8",  x"cd",  x"26",  x"cd",  x"e5", -- 0838
         x"cd",  x"eb",  x"d6",  x"cd",  x"97",  x"d6",  x"e1",  x"c5", -- 0840
         x"d5",  x"f5",  x"33",  x"e5",  x"2a",  x"cf",  x"03",  x"e3", -- 0848
         x"06",  x"81",  x"c5",  x"33",  x"cd",  x"16",  x"de",  x"cd", -- 0850
         x"f9",  x"c8",  x"22",  x"cf",  x"03",  x"7e",  x"fe",  x"3a", -- 0858
         x"28",  x"28",  x"b7",  x"c2",  x"48",  x"c3",  x"23",  x"7e", -- 0860
         x"23",  x"b6",  x"ca",  x"22",  x"c9",  x"23",  x"5e",  x"23", -- 0868
         x"56",  x"ed",  x"53",  x"58",  x"03",  x"3a",  x"0a",  x"03", -- 0870
         x"b7",  x"28",  x"0f",  x"e5",  x"3e",  x"3c",  x"cd",  x"ae", -- 0878
         x"c6",  x"cd",  x"2a",  x"d8",  x"3e",  x"3e",  x"cd",  x"ae", -- 0880
         x"c6",  x"e1",  x"cd",  x"bd",  x"c8",  x"11",  x"54",  x"c8", -- 0888
         x"d5",  x"c8",  x"d6",  x"80",  x"da",  x"5d",  x"ca",  x"fe", -- 0890
         x"25",  x"38",  x"14",  x"d6",  x"50",  x"38",  x"34",  x"fe", -- 0898
         x"05",  x"38",  x"0a",  x"47",  x"3a",  x"fc",  x"03",  x"a7", -- 08A0
         x"28",  x"29",  x"c3",  x"03",  x"e0",  x"c6",  x"25",  x"07", -- 08A8
         x"4f",  x"06",  x"00",  x"eb",  x"21",  x"40",  x"c2",  x"09", -- 08B0
         x"4e",  x"23",  x"46",  x"c5",  x"eb",  x"23",  x"7e",  x"fe", -- 08B8
         x"3a",  x"d0",  x"fe",  x"20",  x"28",  x"f7",  x"fe",  x"30", -- 08C0
         x"3f",  x"3c",  x"3d",  x"c9",  x"7e",  x"e3",  x"be",  x"23", -- 08C8
         x"e3",  x"28",  x"ea",  x"c3",  x"48",  x"c3",  x"3e",  x"2c", -- 08D0
         x"be",  x"18",  x"f6",  x"3e",  x"29",  x"18",  x"f9",  x"eb", -- 08D8
         x"2a",  x"5f",  x"03",  x"28",  x"0e",  x"eb",  x"cd",  x"86", -- 08E0
         x"c9",  x"e5",  x"cd",  x"bb",  x"c4",  x"60",  x"69",  x"d1", -- 08E8
         x"d2",  x"20",  x"ca",  x"2b",  x"22",  x"dd",  x"03",  x"eb", -- 08F0
         x"c9",  x"cd",  x"f3",  x"dd",  x"c0",  x"fe",  x"13",  x"28", -- 08F8
         x"08",  x"fe",  x"03",  x"c0",  x"cd",  x"e4",  x"dd",  x"18", -- 0900
         x"0f",  x"cd",  x"e4",  x"dd",  x"fe",  x"1e",  x"c8",  x"fe", -- 0908
         x"0a",  x"c8",  x"fe",  x"03",  x"28",  x"02",  x"18",  x"f1", -- 0910
         x"c0",  x"f6",  x"c0",  x"22",  x"cf",  x"03",  x"21",  x"f6", -- 0918
         x"ff",  x"c1",  x"2a",  x"58",  x"03",  x"f5",  x"7d",  x"a4", -- 0920
         x"3c",  x"28",  x"09",  x"22",  x"d3",  x"03",  x"2a",  x"cf", -- 0928
         x"03",  x"22",  x"d5",  x"03",  x"af",  x"32",  x"43",  x"03", -- 0930
         x"cd",  x"1d",  x"de",  x"cd",  x"55",  x"cb",  x"f1",  x"21", -- 0938
         x"21",  x"c3",  x"c2",  x"71",  x"c3",  x"c3",  x"88",  x"c3", -- 0940
         x"2a",  x"d5",  x"03",  x"7c",  x"b5",  x"1e",  x"20",  x"ca", -- 0948
         x"56",  x"c3",  x"eb",  x"2a",  x"d3",  x"03",  x"22",  x"58", -- 0950
         x"03",  x"eb",  x"c9",  x"cd",  x"bd",  x"c8",  x"cd",  x"26", -- 0958
         x"cd",  x"cd",  x"97",  x"d6",  x"f2",  x"6f",  x"c9",  x"1e", -- 0960
         x"08",  x"c3",  x"56",  x"c3",  x"cd",  x"26",  x"cd",  x"3a", -- 0968
         x"e8",  x"03",  x"fe",  x"90",  x"da",  x"45",  x"d7",  x"01", -- 0970
         x"80",  x"90",  x"11",  x"00",  x"00",  x"e5",  x"cd",  x"18", -- 0978
         x"d7",  x"e1",  x"51",  x"c8",  x"18",  x"e1",  x"2b",  x"11", -- 0980
         x"00",  x"00",  x"cd",  x"bd",  x"c8",  x"d0",  x"e5",  x"f5", -- 0988
         x"21",  x"98",  x"19",  x"cd",  x"89",  x"c6",  x"da",  x"48", -- 0990
         x"c3",  x"62",  x"6b",  x"19",  x"29",  x"19",  x"29",  x"f1", -- 0998
         x"d6",  x"30",  x"5f",  x"16",  x"00",  x"19",  x"eb",  x"e1", -- 09A0
         x"18",  x"e0",  x"28",  x"3c",  x"cd",  x"5e",  x"c9",  x"cd", -- 09A8
         x"be",  x"c8",  x"e5",  x"2a",  x"b0",  x"03",  x"28",  x"10", -- 09B0
         x"e1",  x"cd",  x"d6",  x"c8",  x"d5",  x"cd",  x"6c",  x"c9", -- 09B8
         x"cd",  x"be",  x"c8",  x"c2",  x"48",  x"c3",  x"e3",  x"eb", -- 09C0
         x"7d",  x"93",  x"5f",  x"7c",  x"9a",  x"57",  x"da",  x"3e", -- 09C8
         x"c3",  x"e5",  x"2a",  x"d7",  x"03",  x"01",  x"28",  x"00", -- 09D0
         x"09",  x"cd",  x"89",  x"c6",  x"d2",  x"3e",  x"c3",  x"eb", -- 09D8
         x"22",  x"56",  x"03",  x"e1",  x"22",  x"b0",  x"03",  x"e1", -- 09E0
         x"c3",  x"53",  x"c6",  x"ca",  x"4f",  x"c6",  x"cd",  x"53", -- 09E8
         x"c6",  x"01",  x"54",  x"c8",  x"18",  x"10",  x"0e",  x"03", -- 09F0
         x"cd",  x"27",  x"c3",  x"c1",  x"e5",  x"e5",  x"2a",  x"58", -- 09F8
         x"03",  x"e3",  x"3e",  x"8c",  x"f5",  x"33",  x"c5",  x"cd", -- 0A00
         x"86",  x"c9",  x"cd",  x"4a",  x"ca",  x"e5",  x"2a",  x"58", -- 0A08
         x"03",  x"cd",  x"89",  x"c6",  x"e1",  x"23",  x"dc",  x"be", -- 0A10
         x"c4",  x"d4",  x"bb",  x"c4",  x"60",  x"69",  x"2b",  x"d8", -- 0A18
         x"1e",  x"0e",  x"c3",  x"56",  x"c3",  x"c0",  x"16",  x"ff", -- 0A20
         x"cd",  x"bd",  x"c7",  x"f9",  x"fe",  x"8c",  x"1e",  x"04", -- 0A28
         x"20",  x"f0",  x"e1",  x"22",  x"58",  x"03",  x"23",  x"7c", -- 0A30
         x"b5",  x"20",  x"07",  x"3a",  x"cd",  x"03",  x"b7",  x"c2", -- 0A38
         x"87",  x"c3",  x"21",  x"54",  x"c8",  x"e3",  x"3e",  x"e1", -- 0A40
         x"01",  x"3a",  x"0e",  x"00",  x"06",  x"00",  x"79",  x"48", -- 0A48
         x"47",  x"7e",  x"b7",  x"c8",  x"b8",  x"c8",  x"23",  x"fe", -- 0A50
         x"22",  x"28",  x"f3",  x"18",  x"f4",  x"cd",  x"06",  x"cf", -- 0A58
         x"cd",  x"cc",  x"c8",  x"b4",  x"d5",  x"3a",  x"ae",  x"03", -- 0A60
         x"f5",  x"cd",  x"3a",  x"cd",  x"f1",  x"e3",  x"22",  x"cf", -- 0A68
         x"03",  x"1f",  x"cd",  x"2b",  x"cd",  x"28",  x"35",  x"e5", -- 0A70
         x"2a",  x"e5",  x"03",  x"e5",  x"23",  x"23",  x"5e",  x"23", -- 0A78
         x"56",  x"2a",  x"5f",  x"03",  x"cd",  x"89",  x"c6",  x"30", -- 0A80
         x"12",  x"2a",  x"56",  x"03",  x"cd",  x"89",  x"c6",  x"d1", -- 0A88
         x"30",  x"11",  x"21",  x"c0",  x"03",  x"cd",  x"89",  x"c6", -- 0A90
         x"30",  x"09",  x"3e",  x"d1",  x"cd",  x"1b",  x"d3",  x"eb", -- 0A98
         x"cd",  x"66",  x"d1",  x"cd",  x"1b",  x"d3",  x"e1",  x"cd", -- 0AA0
         x"fa",  x"d6",  x"e1",  x"c9",  x"e5",  x"cd",  x"f7",  x"d6", -- 0AA8
         x"d1",  x"e1",  x"c9",  x"cd",  x"21",  x"d4",  x"7e",  x"47", -- 0AB0
         x"fe",  x"8c",  x"28",  x"05",  x"cd",  x"cc",  x"c8",  x"88", -- 0AB8
         x"2b",  x"4b",  x"0d",  x"78",  x"ca",  x"92",  x"c8",  x"cd", -- 0AC0
         x"87",  x"c9",  x"fe",  x"2c",  x"c0",  x"18",  x"f3",  x"cd", -- 0AC8
         x"3a",  x"cd",  x"7e",  x"fe",  x"88",  x"28",  x"05",  x"cd", -- 0AD0
         x"cc",  x"c8",  x"a9",  x"2b",  x"cd",  x"29",  x"cd",  x"cd", -- 0AD8
         x"97",  x"d6",  x"20",  x"08",  x"23",  x"7e",  x"b7",  x"c8", -- 0AE0
         x"fe",  x"d4",  x"20",  x"f8",  x"cd",  x"bd",  x"c8",  x"da", -- 0AE8
         x"07",  x"ca",  x"c3",  x"91",  x"c8",  x"cd",  x"be",  x"c8", -- 0AF0
         x"18",  x"07",  x"af",  x"32",  x"fd",  x"03",  x"cd",  x"25", -- 0AF8
         x"de",  x"28",  x"5e",  x"c8",  x"fe",  x"d5",  x"38",  x"09", -- 0B00
         x"3a",  x"fc",  x"03",  x"a7",  x"28",  x"03",  x"cd",  x"06", -- 0B08
         x"e0",  x"fe",  x"a5",  x"ca",  x"92",  x"cb",  x"fe",  x"a8", -- 0B10
         x"28",  x"78",  x"e5",  x"fe",  x"2c",  x"28",  x"5d",  x"fe", -- 0B18
         x"3b",  x"ca",  x"b2",  x"cb",  x"c1",  x"cd",  x"3a",  x"cd", -- 0B20
         x"e5",  x"3a",  x"ae",  x"03",  x"b7",  x"20",  x"20",  x"cd", -- 0B28
         x"34",  x"d8",  x"cd",  x"8a",  x"d1",  x"36",  x"20",  x"2a", -- 0B30
         x"e5",  x"03",  x"34",  x"2a",  x"e5",  x"03",  x"3a",  x"41", -- 0B38
         x"03",  x"47",  x"04",  x"28",  x"0a",  x"04",  x"3a",  x"ac", -- 0B40
         x"03",  x"86",  x"3d",  x"b8",  x"d4",  x"61",  x"cb",  x"cd", -- 0B48
         x"cc",  x"d1",  x"e1",  x"18",  x"a0",  x"3a",  x"ac",  x"03", -- 0B50
         x"b7",  x"c8",  x"18",  x"05",  x"36",  x"00",  x"21",  x"61", -- 0B58
         x"03",  x"3e",  x"0d",  x"cd",  x"ae",  x"c6",  x"3e",  x"0a", -- 0B60
         x"cd",  x"ae",  x"c6",  x"af",  x"32",  x"ac",  x"03",  x"3a", -- 0B68
         x"40",  x"03",  x"3d",  x"c8",  x"f5",  x"af",  x"cd",  x"ae", -- 0B70
         x"c6",  x"f1",  x"18",  x"f6",  x"3a",  x"42",  x"03",  x"47", -- 0B78
         x"3a",  x"ac",  x"03",  x"b8",  x"d4",  x"61",  x"cb",  x"30", -- 0B80
         x"29",  x"d6",  x"0d",  x"38",  x"02",  x"20",  x"fa",  x"2f", -- 0B88
         x"18",  x"15",  x"f5",  x"cd",  x"1e",  x"d4",  x"cd",  x"db", -- 0B90
         x"c8",  x"2b",  x"f1",  x"d6",  x"a8",  x"e5",  x"28",  x"03", -- 0B98
         x"3a",  x"ac",  x"03",  x"2f",  x"83",  x"30",  x"0b",  x"3c", -- 0BA0
         x"28",  x"08",  x"47",  x"3e",  x"20",  x"cd",  x"ae",  x"c6", -- 0BA8
         x"10",  x"fb",  x"e1",  x"cd",  x"bd",  x"c8",  x"c3",  x"03", -- 0BB0
         x"cb",  x"cd",  x"21",  x"d4",  x"32",  x"41",  x"03",  x"c9", -- 0BB8
         x"cd",  x"21",  x"d4",  x"c0",  x"3c",  x"32",  x"40",  x"03", -- 0BC0
         x"c9",  x"3f",  x"52",  x"45",  x"44",  x"4f",  x"20",  x"46", -- 0BC8
         x"52",  x"4f",  x"4d",  x"20",  x"53",  x"54",  x"41",  x"52", -- 0BD0
         x"54",  x"0d",  x"00",  x"3a",  x"ce",  x"03",  x"b7",  x"c2", -- 0BD8
         x"42",  x"c3",  x"c1",  x"21",  x"c9",  x"cb",  x"cd",  x"c9", -- 0BE0
         x"d1",  x"c3",  x"85",  x"c6",  x"cd",  x"37",  x"d1",  x"cd", -- 0BE8
         x"5f",  x"de",  x"af",  x"32",  x"43",  x"03",  x"7e",  x"fe", -- 0BF0
         x"22",  x"20",  x"10",  x"cd",  x"8b",  x"d1",  x"cd",  x"cc", -- 0BF8
         x"c8",  x"3b",  x"e5",  x"cd",  x"cc",  x"d1",  x"cd",  x"d4", -- 0C00
         x"c6",  x"18",  x"04",  x"e5",  x"cd",  x"cf",  x"c6",  x"c1", -- 0C08
         x"38",  x"36",  x"21",  x"62",  x"03",  x"7e",  x"b7",  x"2b", -- 0C10
         x"c5",  x"28",  x"37",  x"36",  x"2c",  x"18",  x"05",  x"e5", -- 0C18
         x"2a",  x"dd",  x"03",  x"f6",  x"af",  x"32",  x"ce",  x"03", -- 0C20
         x"e3",  x"18",  x"03",  x"cd",  x"d6",  x"c8",  x"cd",  x"06", -- 0C28
         x"cf",  x"e3",  x"d5",  x"7e",  x"fe",  x"2c",  x"28",  x"1e", -- 0C30
         x"3a",  x"ce",  x"03",  x"b7",  x"20",  x"7d",  x"3e",  x"3f", -- 0C38
         x"cd",  x"ae",  x"c6",  x"cd",  x"cf",  x"c6",  x"d1",  x"c1", -- 0C40
         x"da",  x"1f",  x"c9",  x"21",  x"62",  x"03",  x"7e",  x"b7", -- 0C48
         x"2b",  x"c5",  x"ca",  x"47",  x"ca",  x"d5",  x"3a",  x"ae", -- 0C50
         x"03",  x"b7",  x"28",  x"21",  x"cd",  x"bd",  x"c8",  x"57", -- 0C58
         x"47",  x"fe",  x"22",  x"28",  x"0c",  x"3a",  x"ce",  x"03", -- 0C60
         x"b7",  x"57",  x"28",  x"02",  x"16",  x"3a",  x"06",  x"2c", -- 0C68
         x"2b",  x"cd",  x"8e",  x"d1",  x"eb",  x"21",  x"88",  x"cc", -- 0C70
         x"e3",  x"d5",  x"c3",  x"77",  x"ca",  x"cd",  x"bd",  x"c8", -- 0C78
         x"cd",  x"a1",  x"d7",  x"e3",  x"cd",  x"f7",  x"d6",  x"e1", -- 0C80
         x"cd",  x"be",  x"c8",  x"28",  x"05",  x"fe",  x"2c",  x"c2", -- 0C88
         x"db",  x"cb",  x"e3",  x"cd",  x"be",  x"c8",  x"20",  x"93", -- 0C90
         x"d1",  x"3a",  x"ce",  x"03",  x"b7",  x"eb",  x"c2",  x"f4", -- 0C98
         x"c8",  x"d5",  x"b6",  x"21",  x"ab",  x"cc",  x"c4",  x"c9", -- 0CA0
         x"d1",  x"e1",  x"c9",  x"3f",  x"45",  x"58",  x"54",  x"52", -- 0CA8
         x"41",  x"20",  x"49",  x"47",  x"4e",  x"4f",  x"52",  x"45", -- 0CB0
         x"44",  x"0d",  x"00",  x"cd",  x"48",  x"ca",  x"b7",  x"20", -- 0CB8
         x"11",  x"23",  x"7e",  x"23",  x"b6",  x"1e",  x"06",  x"ca", -- 0CC0
         x"56",  x"c3",  x"23",  x"5e",  x"23",  x"56",  x"ed",  x"53", -- 0CC8
         x"ca",  x"03",  x"cd",  x"bd",  x"c8",  x"fe",  x"83",  x"20", -- 0CD0
         x"e2",  x"c3",  x"56",  x"cc",  x"11",  x"00",  x"00",  x"c4", -- 0CD8
         x"06",  x"cf",  x"22",  x"cf",  x"03",  x"cd",  x"bd",  x"c7", -- 0CE0
         x"c2",  x"4e",  x"c3",  x"f9",  x"d5",  x"7e",  x"23",  x"f5", -- 0CE8
         x"d5",  x"cd",  x"dd",  x"d6",  x"e3",  x"e5",  x"cd",  x"61", -- 0CF0
         x"d4",  x"e1",  x"cd",  x"f7",  x"d6",  x"e1",  x"cd",  x"ee", -- 0CF8
         x"d6",  x"e5",  x"cd",  x"18",  x"d7",  x"e1",  x"c1",  x"90", -- 0D00
         x"cd",  x"ee",  x"d6",  x"28",  x"09",  x"ed",  x"53",  x"58", -- 0D08
         x"03",  x"69",  x"60",  x"c3",  x"50",  x"c8",  x"f9",  x"2a", -- 0D10
         x"cf",  x"03",  x"7e",  x"fe",  x"2c",  x"c2",  x"54",  x"c8", -- 0D18
         x"cd",  x"bd",  x"c8",  x"cd",  x"df",  x"cc",  x"cd",  x"3a", -- 0D20
         x"cd",  x"f6",  x"37",  x"3a",  x"ae",  x"03",  x"8f",  x"b7", -- 0D28
         x"e8",  x"1e",  x"18",  x"c3",  x"56",  x"c3",  x"cd",  x"cc", -- 0D30
         x"c8",  x"28",  x"2b",  x"16",  x"00",  x"d5",  x"0e",  x"01", -- 0D38
         x"cd",  x"27",  x"c3",  x"cd",  x"ad",  x"cd",  x"22",  x"d1", -- 0D40
         x"03",  x"2a",  x"d1",  x"03",  x"c1",  x"78",  x"fe",  x"78", -- 0D48
         x"d4",  x"29",  x"cd",  x"7e",  x"16",  x"00",  x"d6",  x"b3", -- 0D50
         x"38",  x"15",  x"fe",  x"03",  x"30",  x"11",  x"fe",  x"01", -- 0D58
         x"17",  x"aa",  x"ba",  x"57",  x"da",  x"48",  x"c3",  x"22", -- 0D60
         x"c6",  x"03",  x"cd",  x"bd",  x"c8",  x"18",  x"e7",  x"7a", -- 0D68
         x"b7",  x"c2",  x"84",  x"ce",  x"7e",  x"22",  x"c6",  x"03", -- 0D70
         x"d6",  x"ac",  x"d8",  x"fe",  x"07",  x"d0",  x"5f",  x"3a", -- 0D78
         x"ae",  x"03",  x"3d",  x"b3",  x"7b",  x"ca",  x"b3",  x"d2", -- 0D80
         x"07",  x"83",  x"5f",  x"21",  x"c8",  x"c2",  x"19",  x"78", -- 0D88
         x"56",  x"ba",  x"d0",  x"23",  x"cd",  x"29",  x"cd",  x"c5", -- 0D90
         x"01",  x"49",  x"cd",  x"c5",  x"43",  x"4a",  x"cd",  x"c8", -- 0D98
         x"d6",  x"58",  x"51",  x"4e",  x"23",  x"46",  x"23",  x"c5", -- 0DA0
         x"2a",  x"c6",  x"03",  x"18",  x"90",  x"af",  x"32",  x"ae", -- 0DA8
         x"03",  x"cd",  x"bd",  x"c8",  x"1e",  x"24",  x"ca",  x"56", -- 0DB0
         x"c3",  x"da",  x"a1",  x"d7",  x"cd",  x"8f",  x"c6",  x"30", -- 0DB8
         x"37",  x"fe",  x"ac",  x"28",  x"e8",  x"fe",  x"2e",  x"ca", -- 0DC0
         x"a1",  x"d7",  x"fe",  x"ad",  x"28",  x"19",  x"fe",  x"22", -- 0DC8
         x"ca",  x"8b",  x"d1",  x"fe",  x"aa",  x"ca",  x"e3",  x"ce", -- 0DD0
         x"fe",  x"a7",  x"ca",  x"f0",  x"d0",  x"d6",  x"b6",  x"30", -- 0DD8
         x"28",  x"cd",  x"36",  x"cd",  x"c3",  x"db",  x"c8",  x"16", -- 0DE0
         x"7d",  x"cd",  x"3d",  x"cd",  x"2a",  x"d1",  x"03",  x"e5", -- 0DE8
         x"cd",  x"c0",  x"d6",  x"cd",  x"29",  x"cd",  x"e1",  x"c9", -- 0DF0
         x"cd",  x"06",  x"cf",  x"e5",  x"eb",  x"22",  x"e5",  x"03", -- 0DF8
         x"3a",  x"ae",  x"03",  x"b7",  x"cc",  x"dd",  x"d6",  x"e1", -- 0E00
         x"c9",  x"06",  x"00",  x"07",  x"4f",  x"c5",  x"cd",  x"bd", -- 0E08
         x"c8",  x"79",  x"fe",  x"33",  x"38",  x"07",  x"3a",  x"fc", -- 0E10
         x"03",  x"a7",  x"c2",  x"09",  x"e0",  x"fe",  x"22",  x"28", -- 0E18
         x"1e",  x"fe",  x"2d",  x"38",  x"17",  x"cd",  x"36",  x"cd", -- 0E20
         x"cd",  x"d6",  x"c8",  x"cd",  x"2a",  x"cd",  x"eb",  x"2a", -- 0E28
         x"e5",  x"03",  x"e3",  x"e5",  x"eb",  x"cd",  x"21",  x"d4", -- 0E30
         x"eb",  x"e3",  x"18",  x"08",  x"cd",  x"e1",  x"cd",  x"e3", -- 0E38
         x"11",  x"f3",  x"cd",  x"d5",  x"01",  x"94",  x"c2",  x"09", -- 0E40
         x"4e",  x"23",  x"66",  x"69",  x"e9",  x"15",  x"fe",  x"ad", -- 0E48
         x"c8",  x"fe",  x"2d",  x"c8",  x"14",  x"fe",  x"2b",  x"c8", -- 0E50
         x"fe",  x"ac",  x"c8",  x"2b",  x"c9",  x"f6",  x"af",  x"f5", -- 0E58
         x"cd",  x"29",  x"cd",  x"cd",  x"6f",  x"c9",  x"f1",  x"eb", -- 0E60
         x"c1",  x"e3",  x"eb",  x"cd",  x"e0",  x"d6",  x"f5",  x"cd", -- 0E68
         x"6f",  x"c9",  x"f1",  x"c1",  x"79",  x"21",  x"b0",  x"d0", -- 0E70
         x"20",  x"05",  x"a3",  x"4f",  x"78",  x"a2",  x"e9",  x"b3", -- 0E78
         x"4f",  x"78",  x"b2",  x"e9",  x"21",  x"96",  x"ce",  x"3a", -- 0E80
         x"ae",  x"03",  x"1f",  x"7a",  x"17",  x"5f",  x"16",  x"64", -- 0E88
         x"78",  x"ba",  x"d0",  x"c3",  x"97",  x"cd",  x"98",  x"ce", -- 0E90
         x"79",  x"b7",  x"1f",  x"c1",  x"d1",  x"f5",  x"cd",  x"2b", -- 0E98
         x"cd",  x"21",  x"d9",  x"ce",  x"e5",  x"ca",  x"18",  x"d7", -- 0EA0
         x"af",  x"32",  x"ae",  x"03",  x"d5",  x"cd",  x"fe",  x"d2", -- 0EA8
         x"7e",  x"23",  x"23",  x"4e",  x"23",  x"46",  x"d1",  x"c5", -- 0EB0
         x"f5",  x"cd",  x"02",  x"d3",  x"cd",  x"ee",  x"d6",  x"f1", -- 0EB8
         x"57",  x"e1",  x"7b",  x"b2",  x"c8",  x"7a",  x"d6",  x"01", -- 0EC0
         x"d8",  x"af",  x"bb",  x"3c",  x"d0",  x"15",  x"1d",  x"0a", -- 0EC8
         x"be",  x"23",  x"03",  x"28",  x"ed",  x"3f",  x"c3",  x"a2", -- 0ED0
         x"d6",  x"3c",  x"8f",  x"c1",  x"a0",  x"c6",  x"ff",  x"9f", -- 0ED8
         x"c3",  x"a9",  x"d6",  x"16",  x"5a",  x"cd",  x"3d",  x"cd", -- 0EE0
         x"cd",  x"29",  x"cd",  x"cd",  x"6f",  x"c9",  x"7b",  x"2f", -- 0EE8
         x"4f",  x"7a",  x"2f",  x"cd",  x"b0",  x"d0",  x"c1",  x"c3", -- 0EF0
         x"49",  x"cd",  x"cd",  x"be",  x"c8",  x"c8",  x"cd",  x"d6", -- 0EF8
         x"c8",  x"01",  x"fa",  x"ce",  x"c5",  x"f6",  x"af",  x"32", -- 0F00
         x"ad",  x"03",  x"46",  x"cd",  x"8f",  x"c6",  x"da",  x"48", -- 0F08
         x"c3",  x"af",  x"4f",  x"32",  x"ae",  x"03",  x"cd",  x"bd", -- 0F10
         x"c8",  x"38",  x"05",  x"cd",  x"8f",  x"c6",  x"38",  x"0b", -- 0F18
         x"4f",  x"cd",  x"bd",  x"c8",  x"38",  x"fb",  x"cd",  x"8f", -- 0F20
         x"c6",  x"30",  x"f6",  x"d6",  x"24",  x"20",  x"0a",  x"3c", -- 0F28
         x"32",  x"ae",  x"03",  x"0f",  x"81",  x"4f",  x"cd",  x"bd", -- 0F30
         x"c8",  x"3a",  x"cc",  x"03",  x"3d",  x"ca",  x"dd",  x"cf", -- 0F38
         x"f2",  x"48",  x"cf",  x"7e",  x"d6",  x"28",  x"28",  x"6f", -- 0F40
         x"af",  x"32",  x"cc",  x"03",  x"e5",  x"50",  x"59",  x"2a", -- 0F48
         x"df",  x"03",  x"cd",  x"89",  x"c6",  x"11",  x"e1",  x"03", -- 0F50
         x"ca",  x"e0",  x"d5",  x"2a",  x"d9",  x"03",  x"eb",  x"2a", -- 0F58
         x"d7",  x"03",  x"cd",  x"89",  x"c6",  x"28",  x"10",  x"79", -- 0F60
         x"96",  x"23",  x"20",  x"02",  x"78",  x"96",  x"23",  x"28", -- 0F68
         x"38",  x"23",  x"23",  x"23",  x"23",  x"18",  x"eb",  x"e1", -- 0F70
         x"e3",  x"d5",  x"11",  x"fb",  x"cd",  x"cd",  x"89",  x"c6", -- 0F78
         x"d1",  x"28",  x"29",  x"e3",  x"e5",  x"c5",  x"01",  x"06", -- 0F80
         x"00",  x"2a",  x"db",  x"03",  x"e5",  x"09",  x"c1",  x"e5", -- 0F88
         x"cd",  x"ab",  x"c4",  x"e1",  x"22",  x"db",  x"03",  x"60", -- 0F90
         x"69",  x"22",  x"d9",  x"03",  x"2b",  x"36",  x"00",  x"cd", -- 0F98
         x"89",  x"c6",  x"20",  x"f8",  x"d1",  x"73",  x"23",  x"72", -- 0FA0
         x"23",  x"eb",  x"e1",  x"c9",  x"32",  x"e8",  x"03",  x"21", -- 0FA8
         x"20",  x"c3",  x"22",  x"e5",  x"03",  x"e1",  x"c9",  x"e5", -- 0FB0
         x"2a",  x"ad",  x"03",  x"e3",  x"57",  x"d5",  x"c5",  x"cd", -- 0FB8
         x"5b",  x"c9",  x"c1",  x"f1",  x"eb",  x"e3",  x"e5",  x"eb", -- 0FC0
         x"3c",  x"57",  x"7e",  x"fe",  x"2c",  x"28",  x"ee",  x"cd", -- 0FC8
         x"db",  x"c8",  x"22",  x"d1",  x"03",  x"e1",  x"22",  x"ad", -- 0FD0
         x"03",  x"1e",  x"00",  x"d5",  x"11",  x"e5",  x"f5",  x"2a", -- 0FD8
         x"d9",  x"03",  x"3e",  x"19",  x"ed",  x"5b",  x"db",  x"03", -- 0FE0
         x"cd",  x"89",  x"c6",  x"28",  x"23",  x"7e",  x"b9",  x"23", -- 0FE8
         x"20",  x"02",  x"7e",  x"b8",  x"23",  x"5e",  x"23",  x"56", -- 0FF0
         x"23",  x"20",  x"e8",  x"3a",  x"ad",  x"03",  x"b7",  x"c2", -- 0FF8
         x"51",  x"c3",  x"f1",  x"44",  x"4d",  x"ca",  x"aa",  x"cf", -- 1000
         x"96",  x"28",  x"5f",  x"1e",  x"10",  x"c3",  x"56",  x"c3", -- 1008
         x"11",  x"04",  x"00",  x"f1",  x"ca",  x"67",  x"c9",  x"71", -- 1010
         x"23",  x"70",  x"23",  x"4f",  x"cd",  x"27",  x"c3",  x"23", -- 1018
         x"23",  x"22",  x"c6",  x"03",  x"71",  x"23",  x"3a",  x"ad", -- 1020
         x"03",  x"17",  x"79",  x"01",  x"0b",  x"00",  x"30",  x"02", -- 1028
         x"c1",  x"03",  x"71",  x"23",  x"70",  x"23",  x"f5",  x"e5", -- 1030
         x"cd",  x"89",  x"d7",  x"eb",  x"e1",  x"f1",  x"3d",  x"20", -- 1038
         x"ea",  x"f5",  x"42",  x"4b",  x"eb",  x"19",  x"da",  x"3e", -- 1040
         x"c3",  x"cd",  x"30",  x"c3",  x"22",  x"db",  x"03",  x"2b", -- 1048
         x"36",  x"00",  x"cd",  x"89",  x"c6",  x"20",  x"f8",  x"03", -- 1050
         x"57",  x"2a",  x"c6",  x"03",  x"5e",  x"eb",  x"29",  x"09", -- 1058
         x"eb",  x"2b",  x"2b",  x"73",  x"23",  x"72",  x"23",  x"f1", -- 1060
         x"38",  x"22",  x"47",  x"4f",  x"7e",  x"23",  x"16",  x"e1", -- 1068
         x"5e",  x"23",  x"56",  x"23",  x"e3",  x"f5",  x"cd",  x"89", -- 1070
         x"c6",  x"30",  x"90",  x"e5",  x"cd",  x"89",  x"d7",  x"d1", -- 1078
         x"19",  x"f1",  x"3d",  x"44",  x"4d",  x"20",  x"e8",  x"29", -- 1080
         x"29",  x"c1",  x"09",  x"eb",  x"2a",  x"d1",  x"03",  x"c9", -- 1088
         x"ed",  x"5b",  x"db",  x"03",  x"21",  x"00",  x"00",  x"39", -- 1090
         x"3a",  x"ae",  x"03",  x"b7",  x"28",  x"0d",  x"cd",  x"fe", -- 1098
         x"d2",  x"cd",  x"09",  x"d2",  x"ed",  x"5b",  x"56",  x"03", -- 10A0
         x"2a",  x"c4",  x"03",  x"7d",  x"93",  x"4f",  x"7c",  x"9a", -- 10A8
         x"41",  x"50",  x"1e",  x"00",  x"21",  x"ae",  x"03",  x"73", -- 10B0
         x"06",  x"90",  x"c3",  x"ae",  x"d6",  x"3a",  x"ac",  x"03", -- 10B8
         x"47",  x"af",  x"18",  x"ed",  x"cd",  x"45",  x"d1",  x"cd", -- 10C0
         x"37",  x"d1",  x"01",  x"48",  x"ca",  x"c5",  x"d5",  x"cd", -- 10C8
         x"cc",  x"c8",  x"28",  x"cd",  x"06",  x"cf",  x"e5",  x"eb", -- 10D0
         x"2b",  x"56",  x"2b",  x"5e",  x"e1",  x"cd",  x"29",  x"cd", -- 10D8
         x"cd",  x"db",  x"c8",  x"cd",  x"cc",  x"c8",  x"b4",  x"44", -- 10E0
         x"4d",  x"e3",  x"71",  x"23",  x"70",  x"c3",  x"84",  x"d1", -- 10E8
         x"cd",  x"45",  x"d1",  x"d5",  x"cd",  x"e1",  x"cd",  x"cd", -- 10F0
         x"29",  x"cd",  x"e3",  x"5e",  x"23",  x"56",  x"23",  x"7a", -- 10F8
         x"b3",  x"ca",  x"54",  x"c3",  x"7e",  x"23",  x"66",  x"6f", -- 1100
         x"e5",  x"2a",  x"df",  x"03",  x"e3",  x"22",  x"df",  x"03", -- 1108
         x"2a",  x"e3",  x"03",  x"e5",  x"2a",  x"e1",  x"03",  x"e5", -- 1110
         x"21",  x"e1",  x"03",  x"d5",  x"cd",  x"f7",  x"d6",  x"e1", -- 1118
         x"cd",  x"26",  x"cd",  x"cd",  x"be",  x"c8",  x"c2",  x"48", -- 1120
         x"c3",  x"e1",  x"22",  x"e1",  x"03",  x"e1",  x"22",  x"e3", -- 1128
         x"03",  x"e1",  x"22",  x"df",  x"03",  x"e1",  x"c9",  x"e5", -- 1130
         x"2a",  x"58",  x"03",  x"23",  x"7c",  x"b5",  x"e1",  x"c0", -- 1138
         x"1e",  x"16",  x"c3",  x"56",  x"c3",  x"cd",  x"cc",  x"c8", -- 1140
         x"a7",  x"3e",  x"80",  x"32",  x"cc",  x"03",  x"b6",  x"47", -- 1148
         x"cd",  x"0b",  x"cf",  x"c3",  x"29",  x"cd",  x"cd",  x"29", -- 1150
         x"cd",  x"cd",  x"34",  x"d8",  x"cd",  x"8a",  x"d1",  x"cd", -- 1158
         x"fe",  x"d2",  x"01",  x"57",  x"d3",  x"c5",  x"7e",  x"23", -- 1160
         x"23",  x"e5",  x"cd",  x"e1",  x"d1",  x"e1",  x"4e",  x"23", -- 1168
         x"46",  x"cd",  x"7e",  x"d1",  x"e5",  x"6f",  x"cd",  x"f2", -- 1170
         x"d2",  x"d1",  x"c9",  x"cd",  x"e1",  x"d1",  x"21",  x"c0", -- 1178
         x"03",  x"e5",  x"77",  x"23",  x"23",  x"73",  x"23",  x"72", -- 1180
         x"e1",  x"c9",  x"2b",  x"06",  x"22",  x"50",  x"e5",  x"0e", -- 1188
         x"ff",  x"23",  x"7e",  x"0c",  x"b7",  x"28",  x"06",  x"ba", -- 1190
         x"28",  x"03",  x"b8",  x"20",  x"f4",  x"fe",  x"22",  x"cc", -- 1198
         x"bd",  x"c8",  x"e3",  x"23",  x"eb",  x"79",  x"cd",  x"7e", -- 11A0
         x"d1",  x"11",  x"c0",  x"03",  x"2a",  x"b2",  x"03",  x"22", -- 11A8
         x"e5",  x"03",  x"3e",  x"01",  x"32",  x"ae",  x"03",  x"cd", -- 11B0
         x"fa",  x"d6",  x"cd",  x"89",  x"c6",  x"22",  x"b2",  x"03", -- 11B8
         x"e1",  x"7e",  x"c0",  x"1e",  x"1e",  x"c3",  x"56",  x"c3", -- 11C0
         x"23",  x"cd",  x"8a",  x"d1",  x"cd",  x"fe",  x"d2",  x"cd", -- 11C8
         x"ee",  x"d6",  x"1c",  x"1d",  x"c8",  x"0a",  x"cd",  x"ae", -- 11D0
         x"c6",  x"fe",  x"0d",  x"cc",  x"66",  x"cb",  x"03",  x"18", -- 11D8
         x"f2",  x"b7",  x"0e",  x"f1",  x"f5",  x"ed",  x"5b",  x"56", -- 11E0
         x"03",  x"2a",  x"c4",  x"03",  x"2f",  x"4f",  x"06",  x"ff", -- 11E8
         x"09",  x"23",  x"cd",  x"89",  x"c6",  x"38",  x"07",  x"22", -- 11F0
         x"c4",  x"03",  x"23",  x"eb",  x"f1",  x"c9",  x"f1",  x"1e", -- 11F8
         x"1a",  x"28",  x"c2",  x"bf",  x"f5",  x"01",  x"e3",  x"d1", -- 1200
         x"c5",  x"2a",  x"b0",  x"03",  x"22",  x"c4",  x"03",  x"21", -- 1208
         x"00",  x"00",  x"e5",  x"2a",  x"56",  x"03",  x"e5",  x"21", -- 1210
         x"b4",  x"03",  x"ed",  x"5b",  x"b2",  x"03",  x"cd",  x"89", -- 1218
         x"c6",  x"01",  x"1a",  x"d2",  x"20",  x"3f",  x"2a",  x"d7", -- 1220
         x"03",  x"ed",  x"5b",  x"d9",  x"03",  x"cd",  x"89",  x"c6", -- 1228
         x"28",  x"0a",  x"7e",  x"23",  x"23",  x"b7",  x"cd",  x"68", -- 1230
         x"d2",  x"18",  x"ee",  x"c1",  x"ed",  x"5b",  x"db",  x"03", -- 1238
         x"cd",  x"89",  x"c6",  x"28",  x"49",  x"cd",  x"ee",  x"d6", -- 1240
         x"7b",  x"e5",  x"09",  x"b7",  x"f2",  x"3b",  x"d2",  x"22", -- 1248
         x"c6",  x"03",  x"e1",  x"4e",  x"06",  x"00",  x"09",  x"09", -- 1250
         x"23",  x"ed",  x"5b",  x"c6",  x"03",  x"cd",  x"89",  x"c6", -- 1258
         x"28",  x"da",  x"01",  x"59",  x"d2",  x"c5",  x"f6",  x"80", -- 1260
         x"7e",  x"23",  x"23",  x"5e",  x"23",  x"56",  x"23",  x"f0", -- 1268
         x"b7",  x"c8",  x"44",  x"4d",  x"2a",  x"c4",  x"03",  x"cd", -- 1270
         x"89",  x"c6",  x"60",  x"69",  x"d8",  x"e1",  x"e3",  x"cd", -- 1278
         x"89",  x"c6",  x"e3",  x"e5",  x"60",  x"69",  x"d0",  x"c1", -- 1280
         x"f1",  x"f1",  x"e5",  x"d5",  x"c5",  x"c9",  x"d1",  x"e1", -- 1288
         x"7d",  x"b4",  x"c8",  x"2b",  x"46",  x"2b",  x"4e",  x"e5", -- 1290
         x"2b",  x"2b",  x"6e",  x"26",  x"00",  x"09",  x"50",  x"59", -- 1298
         x"2b",  x"44",  x"4d",  x"2a",  x"c4",  x"03",  x"cd",  x"ae", -- 12A0
         x"c4",  x"e1",  x"71",  x"23",  x"70",  x"69",  x"60",  x"2b", -- 12A8
         x"c3",  x"0c",  x"d2",  x"c5",  x"e5",  x"2a",  x"e5",  x"03", -- 12B0
         x"e3",  x"cd",  x"ad",  x"cd",  x"e3",  x"cd",  x"2a",  x"cd", -- 12B8
         x"7e",  x"e5",  x"2a",  x"e5",  x"03",  x"e5",  x"86",  x"1e", -- 12C0
         x"1c",  x"da",  x"56",  x"c3",  x"cd",  x"7b",  x"d1",  x"d1", -- 12C8
         x"cd",  x"02",  x"d3",  x"e3",  x"cd",  x"01",  x"d3",  x"e5", -- 12D0
         x"2a",  x"c2",  x"03",  x"eb",  x"cd",  x"e9",  x"d2",  x"cd", -- 12D8
         x"e9",  x"d2",  x"21",  x"46",  x"cd",  x"e3",  x"e5",  x"18", -- 12E0
         x"6f",  x"e1",  x"e3",  x"7e",  x"23",  x"23",  x"4e",  x"23", -- 12E8
         x"46",  x"6f",  x"2c",  x"2d",  x"c8",  x"0a",  x"12",  x"03", -- 12F0
         x"13",  x"18",  x"f8",  x"cd",  x"2a",  x"cd",  x"2a",  x"e5", -- 12F8
         x"03",  x"eb",  x"cd",  x"1b",  x"d3",  x"eb",  x"c0",  x"d5", -- 1300
         x"50",  x"59",  x"1b",  x"4e",  x"2a",  x"c4",  x"03",  x"cd", -- 1308
         x"89",  x"c6",  x"20",  x"05",  x"47",  x"09",  x"22",  x"c4", -- 1310
         x"03",  x"e1",  x"c9",  x"2a",  x"b2",  x"03",  x"2b",  x"46", -- 1318
         x"2b",  x"4e",  x"2b",  x"2b",  x"cd",  x"89",  x"c6",  x"c0", -- 1320
         x"22",  x"b2",  x"03",  x"c9",  x"01",  x"c0",  x"d0",  x"c5", -- 1328
         x"cd",  x"fb",  x"d2",  x"af",  x"57",  x"32",  x"ae",  x"03", -- 1330
         x"7e",  x"b7",  x"c9",  x"01",  x"c0",  x"d0",  x"c5",  x"cd", -- 1338
         x"30",  x"d3",  x"28",  x"55",  x"23",  x"23",  x"5e",  x"23", -- 1340
         x"56",  x"1a",  x"c9",  x"3e",  x"01",  x"cd",  x"7b",  x"d1", -- 1348
         x"cd",  x"24",  x"d4",  x"2a",  x"c2",  x"03",  x"73",  x"c1", -- 1350
         x"c3",  x"a9",  x"d1",  x"cd",  x"da",  x"d3",  x"af",  x"e3", -- 1358
         x"4f",  x"e5",  x"7e",  x"b8",  x"38",  x"02",  x"78",  x"11", -- 1360
         x"0e",  x"00",  x"c5",  x"cd",  x"e1",  x"d1",  x"c1",  x"e1", -- 1368
         x"e5",  x"23",  x"23",  x"46",  x"23",  x"66",  x"68",  x"06", -- 1370
         x"00",  x"09",  x"44",  x"4d",  x"cd",  x"7e",  x"d1",  x"6f", -- 1378
         x"cd",  x"f2",  x"d2",  x"d1",  x"cd",  x"02",  x"d3",  x"18", -- 1380
         x"cf",  x"cd",  x"da",  x"d3",  x"d1",  x"d5",  x"1a",  x"90", -- 1388
         x"18",  x"cd",  x"eb",  x"7e",  x"cd",  x"de",  x"d3",  x"04", -- 1390
         x"05",  x"ca",  x"67",  x"c9",  x"c5",  x"1e",  x"ff",  x"fe", -- 1398
         x"29",  x"28",  x"06",  x"cd",  x"d6",  x"c8",  x"cd",  x"21", -- 13A0
         x"d4",  x"cd",  x"db",  x"c8",  x"f1",  x"e3",  x"01",  x"61", -- 13A8
         x"d3",  x"c5",  x"3d",  x"be",  x"06",  x"00",  x"d0",  x"4f", -- 13B0
         x"7e",  x"91",  x"bb",  x"47",  x"d8",  x"43",  x"c9",  x"cd", -- 13B8
         x"30",  x"d3",  x"ca",  x"cf",  x"d4",  x"5f",  x"23",  x"23", -- 13C0
         x"7e",  x"23",  x"66",  x"6f",  x"e5",  x"19",  x"46",  x"72", -- 13C8
         x"e3",  x"c5",  x"7e",  x"cd",  x"a1",  x"d7",  x"c1",  x"e1", -- 13D0
         x"70",  x"c9",  x"eb",  x"cd",  x"db",  x"c8",  x"c1",  x"d1", -- 13D8
         x"c5",  x"43",  x"c9",  x"cd",  x"24",  x"d4",  x"4f",  x"ed", -- 13E0
         x"78",  x"c3",  x"c0",  x"d0",  x"cd",  x"14",  x"d4",  x"3a", -- 13E8
         x"06",  x"03",  x"4f",  x"7b",  x"ed",  x"79",  x"c9",  x"cd", -- 13F0
         x"14",  x"d4",  x"f5",  x"1e",  x"00",  x"cd",  x"be",  x"c8", -- 13F8
         x"28",  x"06",  x"cd",  x"d6",  x"c8",  x"cd",  x"21",  x"d4", -- 1400
         x"c1",  x"3a",  x"06",  x"03",  x"4f",  x"ed",  x"78",  x"ab", -- 1408
         x"a0",  x"28",  x"fa",  x"c9",  x"cd",  x"21",  x"d4",  x"32", -- 1410
         x"06",  x"03",  x"cd",  x"d6",  x"c8",  x"2b",  x"cd",  x"bd", -- 1418
         x"c8",  x"cd",  x"26",  x"cd",  x"cd",  x"61",  x"c9",  x"7a", -- 1420
         x"b7",  x"c2",  x"67",  x"c9",  x"cd",  x"be",  x"c8",  x"7b", -- 1428
         x"c9",  x"cd",  x"6f",  x"c9",  x"1a",  x"18",  x"b2",  x"cd", -- 1430
         x"6c",  x"c9",  x"d5",  x"cd",  x"d6",  x"c8",  x"cd",  x"21", -- 1438
         x"d4",  x"d1",  x"12",  x"c9",  x"cd",  x"6f",  x"c9",  x"eb", -- 1440
         x"46",  x"23",  x"7e",  x"c3",  x"b1",  x"d0",  x"cd",  x"6c", -- 1448
         x"c9",  x"d5",  x"cd",  x"d6",  x"c8",  x"cd",  x"6c",  x"c9", -- 1450
         x"e3",  x"73",  x"23",  x"72",  x"e1",  x"c9",  x"21",  x"04", -- 1458
         x"d9",  x"cd",  x"ee",  x"d6",  x"18",  x"09",  x"cd",  x"ee", -- 1460
         x"d6",  x"21",  x"c1",  x"d1",  x"cd",  x"c0",  x"d6",  x"78", -- 1468
         x"b7",  x"c8",  x"3a",  x"e8",  x"03",  x"b7",  x"ca",  x"e0", -- 1470
         x"d6",  x"90",  x"30",  x"0c",  x"2f",  x"3c",  x"eb",  x"cd", -- 1478
         x"c8",  x"d6",  x"eb",  x"cd",  x"e0",  x"d6",  x"c1",  x"d1", -- 1480
         x"fe",  x"19",  x"d0",  x"f5",  x"cd",  x"03",  x"d7",  x"67", -- 1488
         x"f1",  x"cd",  x"2a",  x"d5",  x"b4",  x"21",  x"e5",  x"03", -- 1490
         x"f2",  x"ab",  x"d4",  x"cd",  x"0a",  x"d5",  x"30",  x"4b", -- 1498
         x"23",  x"34",  x"28",  x"63",  x"2e",  x"01",  x"cd",  x"3e", -- 14A0
         x"d5",  x"18",  x"40",  x"af",  x"90",  x"47",  x"7e",  x"9b", -- 14A8
         x"5f",  x"23",  x"7e",  x"9a",  x"57",  x"23",  x"7e",  x"99", -- 14B0
         x"4f",  x"dc",  x"16",  x"d5",  x"68",  x"63",  x"af",  x"47", -- 14B8
         x"79",  x"b7",  x"20",  x"16",  x"4a",  x"54",  x"65",  x"6f", -- 14C0
         x"78",  x"d6",  x"08",  x"fe",  x"e0",  x"20",  x"f0",  x"af", -- 14C8
         x"32",  x"e8",  x"03",  x"c9",  x"05",  x"29",  x"cb",  x"12", -- 14D0
         x"cb",  x"11",  x"f2",  x"d4",  x"d4",  x"78",  x"5c",  x"45", -- 14D8
         x"b7",  x"28",  x"08",  x"21",  x"e8",  x"03",  x"86",  x"77", -- 14E0
         x"30",  x"e5",  x"c8",  x"78",  x"21",  x"e8",  x"03",  x"b7", -- 14E8
         x"fc",  x"fd",  x"d4",  x"46",  x"23",  x"7e",  x"e6",  x"80", -- 14F0
         x"a9",  x"4f",  x"c3",  x"e0",  x"d6",  x"1c",  x"c0",  x"14", -- 14F8
         x"c0",  x"0c",  x"c0",  x"0e",  x"80",  x"34",  x"c0",  x"c3", -- 1500
         x"53",  x"d6",  x"7e",  x"83",  x"5f",  x"23",  x"7e",  x"8a", -- 1508
         x"57",  x"23",  x"7e",  x"89",  x"4f",  x"c9",  x"21",  x"e9", -- 1510
         x"03",  x"7e",  x"2f",  x"77",  x"af",  x"6f",  x"90",  x"47", -- 1518
         x"7d",  x"9b",  x"5f",  x"7d",  x"9a",  x"57",  x"7d",  x"99", -- 1520
         x"4f",  x"c9",  x"06",  x"00",  x"d6",  x"08",  x"38",  x"07", -- 1528
         x"43",  x"5a",  x"51",  x"0e",  x"00",  x"18",  x"f5",  x"c6", -- 1530
         x"09",  x"6f",  x"af",  x"2d",  x"c8",  x"79",  x"1f",  x"4f", -- 1538
         x"cb",  x"1a",  x"cb",  x"1b",  x"cb",  x"18",  x"18",  x"f2", -- 1540
         x"00",  x"00",  x"00",  x"81",  x"03",  x"aa",  x"56",  x"19", -- 1548
         x"80",  x"f1",  x"22",  x"76",  x"80",  x"45",  x"aa",  x"38", -- 1550
         x"82",  x"cd",  x"97",  x"d6",  x"b7",  x"ea",  x"67",  x"c9", -- 1558
         x"21",  x"e8",  x"03",  x"7e",  x"01",  x"35",  x"80",  x"11", -- 1560
         x"f3",  x"04",  x"90",  x"f5",  x"70",  x"d5",  x"c5",  x"cd", -- 1568
         x"6f",  x"d4",  x"c1",  x"d1",  x"04",  x"cd",  x"f5",  x"d5", -- 1570
         x"21",  x"48",  x"d5",  x"cd",  x"66",  x"d4",  x"21",  x"4c", -- 1578
         x"d5",  x"cd",  x"ce",  x"d9",  x"01",  x"80",  x"80",  x"11", -- 1580
         x"00",  x"00",  x"cd",  x"6f",  x"d4",  x"f1",  x"cd",  x"0b", -- 1588
         x"d8",  x"01",  x"31",  x"80",  x"11",  x"18",  x"72",  x"21", -- 1590
         x"c1",  x"d1",  x"cd",  x"97",  x"d6",  x"c8",  x"2e",  x"00", -- 1598
         x"cd",  x"58",  x"d6",  x"79",  x"32",  x"f7",  x"03",  x"eb", -- 15A0
         x"22",  x"f8",  x"03",  x"01",  x"00",  x"00",  x"50",  x"58", -- 15A8
         x"21",  x"bc",  x"d4",  x"e5",  x"21",  x"bc",  x"d5",  x"e5", -- 15B0
         x"e5",  x"21",  x"e5",  x"03",  x"7e",  x"23",  x"b7",  x"28", -- 15B8
         x"21",  x"e5",  x"2e",  x"08",  x"1f",  x"67",  x"79",  x"30", -- 15C0
         x"0b",  x"e5",  x"2a",  x"f8",  x"03",  x"19",  x"eb",  x"e1", -- 15C8
         x"3a",  x"f7",  x"03",  x"89",  x"1f",  x"4f",  x"cb",  x"1a", -- 15D0
         x"cb",  x"1b",  x"cb",  x"18",  x"2d",  x"7c",  x"20",  x"e4", -- 15D8
         x"e1",  x"c9",  x"43",  x"5a",  x"51",  x"4f",  x"c9",  x"cd", -- 15E0
         x"c8",  x"d6",  x"01",  x"20",  x"84",  x"11",  x"00",  x"00", -- 15E8
         x"cd",  x"e0",  x"d6",  x"c1",  x"d1",  x"cd",  x"97",  x"d6", -- 15F0
         x"ca",  x"4b",  x"c3",  x"2e",  x"ff",  x"cd",  x"58",  x"d6", -- 15F8
         x"34",  x"34",  x"2b",  x"7e",  x"32",  x"14",  x"03",  x"2b", -- 1600
         x"7e",  x"32",  x"10",  x"03",  x"2b",  x"7e",  x"32",  x"0c", -- 1608
         x"03",  x"41",  x"eb",  x"af",  x"4f",  x"57",  x"5f",  x"32", -- 1610
         x"17",  x"03",  x"e5",  x"c5",  x"7d",  x"cd",  x"0b",  x"03", -- 1618
         x"de",  x"00",  x"3f",  x"30",  x"07",  x"32",  x"17",  x"03", -- 1620
         x"f1",  x"f1",  x"37",  x"d2",  x"c1",  x"e1",  x"79",  x"3c", -- 1628
         x"3d",  x"1f",  x"fa",  x"ec",  x"d4",  x"17",  x"cb",  x"13", -- 1630
         x"cb",  x"12",  x"cb",  x"11",  x"29",  x"cb",  x"10",  x"3a", -- 1638
         x"17",  x"03",  x"17",  x"32",  x"17",  x"03",  x"79",  x"b2", -- 1640
         x"b3",  x"20",  x"cf",  x"e5",  x"21",  x"e8",  x"03",  x"35", -- 1648
         x"e1",  x"20",  x"c7",  x"1e",  x"0a",  x"c3",  x"56",  x"c3", -- 1650
         x"78",  x"b7",  x"ca",  x"7c",  x"d6",  x"7d",  x"21",  x"e8", -- 1658
         x"03",  x"ae",  x"80",  x"47",  x"1f",  x"a8",  x"78",  x"f2", -- 1660
         x"7b",  x"d6",  x"c6",  x"80",  x"77",  x"ca",  x"e0",  x"d5", -- 1668
         x"cd",  x"03",  x"d7",  x"77",  x"2b",  x"c9",  x"cd",  x"97", -- 1670
         x"d6",  x"2f",  x"e1",  x"b7",  x"e1",  x"f2",  x"cf",  x"d4", -- 1678
         x"18",  x"d1",  x"cd",  x"eb",  x"d6",  x"78",  x"b7",  x"c8", -- 1680
         x"c6",  x"02",  x"38",  x"c7",  x"47",  x"cd",  x"6f",  x"d4", -- 1688
         x"21",  x"e8",  x"03",  x"34",  x"c0",  x"18",  x"bc",  x"3a", -- 1690
         x"e8",  x"03",  x"b7",  x"c8",  x"3a",  x"e7",  x"03",  x"fe", -- 1698
         x"2f",  x"17",  x"9f",  x"c0",  x"3c",  x"c9",  x"cd",  x"97", -- 16A0
         x"d6",  x"06",  x"88",  x"11",  x"00",  x"00",  x"21",  x"e8", -- 16A8
         x"03",  x"4f",  x"70",  x"06",  x"00",  x"23",  x"36",  x"80", -- 16B0
         x"17",  x"c3",  x"b9",  x"d4",  x"cd",  x"97",  x"d6",  x"f0", -- 16B8
         x"21",  x"e7",  x"03",  x"7e",  x"ee",  x"80",  x"77",  x"c9", -- 16C0
         x"eb",  x"2a",  x"e5",  x"03",  x"e3",  x"e5",  x"2a",  x"e7", -- 16C8
         x"03",  x"e3",  x"e5",  x"eb",  x"c9",  x"01",  x"49",  x"82", -- 16D0
         x"11",  x"db",  x"0f",  x"18",  x"03",  x"cd",  x"ee",  x"d6", -- 16D8
         x"ed",  x"53",  x"e5",  x"03",  x"ed",  x"43",  x"e7",  x"03", -- 16E0
         x"50",  x"59",  x"c9",  x"21",  x"e5",  x"03",  x"5e",  x"23", -- 16E8
         x"56",  x"23",  x"4e",  x"23",  x"46",  x"23",  x"c9",  x"11", -- 16F0
         x"e5",  x"03",  x"06",  x"04",  x"1a",  x"77",  x"13",  x"23", -- 16F8
         x"10",  x"fa",  x"c9",  x"21",  x"e7",  x"03",  x"7e",  x"07", -- 1700
         x"37",  x"1f",  x"77",  x"3f",  x"1f",  x"23",  x"23",  x"77", -- 1708
         x"79",  x"07",  x"37",  x"1f",  x"4f",  x"1f",  x"ae",  x"c9", -- 1710
         x"78",  x"b7",  x"ca",  x"97",  x"d6",  x"21",  x"a0",  x"d6", -- 1718
         x"e5",  x"cd",  x"97",  x"d6",  x"79",  x"c8",  x"21",  x"e7", -- 1720
         x"03",  x"ae",  x"79",  x"f8",  x"cd",  x"32",  x"d7",  x"1f", -- 1728
         x"a9",  x"c9",  x"23",  x"78",  x"be",  x"c0",  x"2b",  x"79", -- 1730
         x"be",  x"c0",  x"2b",  x"7a",  x"be",  x"c0",  x"2b",  x"7b", -- 1738
         x"96",  x"c0",  x"e1",  x"e1",  x"c9",  x"47",  x"4f",  x"57", -- 1740
         x"5f",  x"b7",  x"c8",  x"e5",  x"cd",  x"eb",  x"d6",  x"cd", -- 1748
         x"03",  x"d7",  x"ae",  x"67",  x"fc",  x"69",  x"d7",  x"3e", -- 1750
         x"98",  x"90",  x"cd",  x"2a",  x"d5",  x"7c",  x"17",  x"dc", -- 1758
         x"fd",  x"d4",  x"06",  x"00",  x"dc",  x"16",  x"d5",  x"e1", -- 1760
         x"c9",  x"1b",  x"7a",  x"a3",  x"3c",  x"c0",  x"0b",  x"c9", -- 1768
         x"21",  x"e8",  x"03",  x"7e",  x"fe",  x"98",  x"3a",  x"e5", -- 1770
         x"03",  x"d0",  x"7e",  x"cd",  x"45",  x"d7",  x"36",  x"98", -- 1778
         x"7b",  x"f5",  x"79",  x"17",  x"cd",  x"b9",  x"d4",  x"f1", -- 1780
         x"c9",  x"21",  x"00",  x"00",  x"78",  x"b1",  x"c8",  x"3e", -- 1788
         x"10",  x"29",  x"38",  x"06",  x"eb",  x"29",  x"eb",  x"30", -- 1790
         x"04",  x"09",  x"da",  x"0b",  x"d0",  x"3d",  x"20",  x"f1", -- 1798
         x"c9",  x"fe",  x"2d",  x"f5",  x"28",  x"05",  x"fe",  x"2b", -- 17A0
         x"28",  x"01",  x"2b",  x"cd",  x"cf",  x"d4",  x"47",  x"57", -- 17A8
         x"5f",  x"2f",  x"4f",  x"cd",  x"bd",  x"c8",  x"38",  x"3d", -- 17B0
         x"fe",  x"2e",  x"28",  x"16",  x"fe",  x"45",  x"20",  x"15", -- 17B8
         x"cd",  x"bd",  x"c8",  x"cd",  x"4d",  x"ce",  x"cd",  x"bd", -- 17C0
         x"c8",  x"38",  x"4b",  x"14",  x"20",  x"07",  x"af",  x"93", -- 17C8
         x"5f",  x"0c",  x"0c",  x"28",  x"de",  x"e5",  x"7b",  x"90", -- 17D0
         x"f4",  x"ed",  x"d7",  x"f2",  x"e4",  x"d7",  x"f5",  x"cd", -- 17D8
         x"e7",  x"d5",  x"f1",  x"3c",  x"20",  x"f2",  x"d1",  x"f1", -- 17E0
         x"cc",  x"c0",  x"d6",  x"eb",  x"c9",  x"c8",  x"f5",  x"cd", -- 17E8
         x"82",  x"d6",  x"f1",  x"3d",  x"c9",  x"d5",  x"57",  x"78", -- 17F0
         x"89",  x"47",  x"c5",  x"e5",  x"d5",  x"cd",  x"82",  x"d6", -- 17F8
         x"f1",  x"d6",  x"30",  x"cd",  x"0b",  x"d8",  x"e1",  x"c1", -- 1800
         x"d1",  x"18",  x"a8",  x"cd",  x"c8",  x"d6",  x"cd",  x"a9", -- 1808
         x"d6",  x"c1",  x"d1",  x"c3",  x"6f",  x"d4",  x"7b",  x"07", -- 1810
         x"07",  x"83",  x"07",  x"86",  x"d6",  x"30",  x"5f",  x"18", -- 1818
         x"a5",  x"e5",  x"21",  x"0d",  x"c3",  x"cd",  x"c9",  x"d1", -- 1820
         x"e1",  x"eb",  x"af",  x"06",  x"98",  x"cd",  x"ae",  x"d6", -- 1828
         x"21",  x"c8",  x"d1",  x"e5",  x"21",  x"ea",  x"03",  x"e5", -- 1830
         x"cd",  x"97",  x"d6",  x"36",  x"20",  x"f2",  x"42",  x"d8", -- 1838
         x"36",  x"2d",  x"23",  x"36",  x"30",  x"ca",  x"ef",  x"d8", -- 1840
         x"e5",  x"fc",  x"c0",  x"d6",  x"af",  x"f5",  x"cd",  x"f5", -- 1848
         x"d8",  x"01",  x"43",  x"91",  x"11",  x"f8",  x"4f",  x"cd", -- 1850
         x"18",  x"d7",  x"b7",  x"e2",  x"6e",  x"d8",  x"f1",  x"cd", -- 1858
         x"ee",  x"d7",  x"f5",  x"18",  x"ec",  x"cd",  x"e7",  x"d5", -- 1860
         x"f1",  x"3c",  x"f5",  x"cd",  x"f5",  x"d8",  x"cd",  x"5e", -- 1868
         x"d4",  x"3c",  x"cd",  x"45",  x"d7",  x"cd",  x"e0",  x"d6", -- 1870
         x"01",  x"06",  x"03",  x"f1",  x"81",  x"3c",  x"fa",  x"89", -- 1878
         x"d8",  x"fe",  x"08",  x"30",  x"04",  x"3c",  x"47",  x"3e", -- 1880
         x"02",  x"3d",  x"3d",  x"e1",  x"f5",  x"11",  x"08",  x"d9", -- 1888
         x"05",  x"20",  x"06",  x"36",  x"2e",  x"23",  x"36",  x"30", -- 1890
         x"23",  x"05",  x"36",  x"2e",  x"cc",  x"f5",  x"d6",  x"c5", -- 1898
         x"e5",  x"d5",  x"cd",  x"eb",  x"d6",  x"e1",  x"06",  x"2f", -- 18A0
         x"04",  x"7b",  x"96",  x"5f",  x"23",  x"7a",  x"9e",  x"57", -- 18A8
         x"23",  x"79",  x"9e",  x"4f",  x"2b",  x"2b",  x"30",  x"f0", -- 18B0
         x"cd",  x"0a",  x"d5",  x"23",  x"cd",  x"e0",  x"d6",  x"eb", -- 18B8
         x"e1",  x"70",  x"23",  x"c1",  x"0d",  x"20",  x"d2",  x"05", -- 18C0
         x"28",  x"0b",  x"2b",  x"7e",  x"fe",  x"30",  x"28",  x"fa", -- 18C8
         x"fe",  x"2e",  x"c4",  x"f5",  x"d6",  x"f1",  x"28",  x"1a", -- 18D0
         x"36",  x"45",  x"23",  x"36",  x"2b",  x"f2",  x"e4",  x"d8", -- 18D8
         x"36",  x"2d",  x"2f",  x"3c",  x"06",  x"2f",  x"04",  x"d6", -- 18E0
         x"0a",  x"30",  x"fb",  x"c6",  x"3a",  x"23",  x"70",  x"23", -- 18E8
         x"77",  x"23",  x"71",  x"e1",  x"c9",  x"01",  x"74",  x"94", -- 18F0
         x"11",  x"f7",  x"23",  x"cd",  x"18",  x"d7",  x"b7",  x"e1", -- 18F8
         x"e2",  x"65",  x"d8",  x"e9",  x"00",  x"00",  x"00",  x"80", -- 1900
         x"a0",  x"86",  x"01",  x"10",  x"27",  x"00",  x"e8",  x"03", -- 1908
         x"00",  x"64",  x"00",  x"00",  x"0a",  x"00",  x"00",  x"01", -- 1910
         x"00",  x"00",  x"21",  x"c0",  x"d6",  x"e3",  x"e9",  x"cd", -- 1918
         x"c8",  x"d6",  x"21",  x"04",  x"d9",  x"cd",  x"dd",  x"d6", -- 1920
         x"c1",  x"d1",  x"cd",  x"97",  x"d6",  x"78",  x"ca",  x"6d", -- 1928
         x"d9",  x"f2",  x"38",  x"d9",  x"b7",  x"ca",  x"4b",  x"c3", -- 1930
         x"b7",  x"ca",  x"d0",  x"d4",  x"d5",  x"c5",  x"79",  x"f6", -- 1938
         x"7f",  x"cd",  x"eb",  x"d6",  x"f2",  x"55",  x"d9",  x"d5", -- 1940
         x"c5",  x"cd",  x"70",  x"d7",  x"c1",  x"d1",  x"f5",  x"cd", -- 1948
         x"18",  x"d7",  x"e1",  x"7c",  x"1f",  x"e1",  x"22",  x"e7", -- 1950
         x"03",  x"e1",  x"22",  x"e5",  x"03",  x"dc",  x"1a",  x"d9", -- 1958
         x"cc",  x"c0",  x"d6",  x"d5",  x"c5",  x"cd",  x"59",  x"d5", -- 1960
         x"c1",  x"d1",  x"cd",  x"9a",  x"d5",  x"cd",  x"c8",  x"d6", -- 1968
         x"01",  x"38",  x"81",  x"11",  x"3b",  x"aa",  x"cd",  x"9a", -- 1970
         x"d5",  x"3a",  x"e8",  x"03",  x"fe",  x"88",  x"d2",  x"76", -- 1978
         x"d6",  x"cd",  x"70",  x"d7",  x"c6",  x"80",  x"c6",  x"02", -- 1980
         x"da",  x"76",  x"d6",  x"f5",  x"21",  x"48",  x"d5",  x"cd", -- 1988
         x"61",  x"d4",  x"cd",  x"91",  x"d5",  x"f1",  x"c1",  x"d1", -- 1990
         x"f5",  x"cd",  x"6c",  x"d4",  x"cd",  x"c0",  x"d6",  x"21", -- 1998
         x"ad",  x"d9",  x"cd",  x"dd",  x"d9",  x"11",  x"00",  x"00", -- 19A0
         x"c1",  x"4a",  x"c3",  x"9a",  x"d5",  x"08",  x"40",  x"2e", -- 19A8
         x"94",  x"74",  x"70",  x"4f",  x"2e",  x"77",  x"6e",  x"02", -- 19B0
         x"88",  x"7a",  x"e6",  x"a0",  x"2a",  x"7c",  x"50",  x"aa", -- 19B8
         x"aa",  x"7e",  x"ff",  x"ff",  x"7f",  x"7f",  x"00",  x"00", -- 19C0
         x"80",  x"81",  x"00",  x"00",  x"00",  x"81",  x"cd",  x"c8", -- 19C8
         x"d6",  x"11",  x"98",  x"d5",  x"d5",  x"e5",  x"cd",  x"eb", -- 19D0
         x"d6",  x"cd",  x"9a",  x"d5",  x"e1",  x"cd",  x"c8",  x"d6", -- 19D8
         x"7e",  x"23",  x"cd",  x"dd",  x"d6",  x"06",  x"f1",  x"c1", -- 19E0
         x"d1",  x"3d",  x"c8",  x"d5",  x"c5",  x"f5",  x"e5",  x"cd", -- 19E8
         x"9a",  x"d5",  x"e1",  x"cd",  x"ee",  x"d6",  x"e5",  x"cd", -- 19F0
         x"6f",  x"d4",  x"e1",  x"18",  x"e9",  x"cd",  x"97",  x"d6", -- 19F8
         x"21",  x"1b",  x"03",  x"fa",  x"5d",  x"da",  x"21",  x"3c", -- 1A00
         x"03",  x"cd",  x"dd",  x"d6",  x"21",  x"1b",  x"03",  x"c8", -- 1A08
         x"86",  x"e6",  x"07",  x"06",  x"00",  x"77",  x"23",  x"87", -- 1A10
         x"87",  x"4f",  x"09",  x"cd",  x"ee",  x"d6",  x"cd",  x"9a", -- 1A18
         x"d5",  x"3a",  x"1a",  x"03",  x"3c",  x"e6",  x"03",  x"06", -- 1A20
         x"00",  x"fe",  x"01",  x"88",  x"32",  x"1a",  x"03",  x"21", -- 1A28
         x"60",  x"da",  x"87",  x"87",  x"4f",  x"09",  x"cd",  x"61", -- 1A30
         x"d4",  x"cd",  x"eb",  x"d6",  x"7b",  x"59",  x"ee",  x"4f", -- 1A38
         x"4f",  x"36",  x"80",  x"2b",  x"46",  x"36",  x"80",  x"21", -- 1A40
         x"19",  x"03",  x"34",  x"7e",  x"d6",  x"ab",  x"20",  x"04", -- 1A48
         x"77",  x"0c",  x"15",  x"1c",  x"cd",  x"bc",  x"d4",  x"21", -- 1A50
         x"3c",  x"03",  x"c3",  x"f7",  x"d6",  x"77",  x"2b",  x"77", -- 1A58
         x"2b",  x"77",  x"18",  x"d5",  x"68",  x"b1",  x"46",  x"68", -- 1A60
         x"99",  x"e9",  x"92",  x"69",  x"10",  x"d1",  x"75",  x"68", -- 1A68
         x"21",  x"ba",  x"da",  x"cd",  x"61",  x"d4",  x"cd",  x"c8", -- 1A70
         x"d6",  x"01",  x"49",  x"83",  x"11",  x"db",  x"0f",  x"cd", -- 1A78
         x"e0",  x"d6",  x"c1",  x"d1",  x"cd",  x"f5",  x"d5",  x"cd", -- 1A80
         x"c8",  x"d6",  x"cd",  x"70",  x"d7",  x"c1",  x"d1",  x"cd", -- 1A88
         x"6c",  x"d4",  x"21",  x"be",  x"da",  x"cd",  x"66",  x"d4", -- 1A90
         x"cd",  x"97",  x"d6",  x"37",  x"f2",  x"a6",  x"da",  x"cd", -- 1A98
         x"5e",  x"d4",  x"cd",  x"97",  x"d6",  x"b7",  x"f5",  x"f4", -- 1AA0
         x"c0",  x"d6",  x"21",  x"be",  x"da",  x"cd",  x"61",  x"d4", -- 1AA8
         x"f1",  x"d4",  x"c0",  x"d6",  x"21",  x"c2",  x"da",  x"c3", -- 1AB0
         x"ce",  x"d9",  x"db",  x"0f",  x"49",  x"81",  x"00",  x"00", -- 1AB8
         x"00",  x"7f",  x"05",  x"ba",  x"d7",  x"1e",  x"86",  x"64", -- 1AC0
         x"26",  x"99",  x"87",  x"58",  x"34",  x"23",  x"87",  x"e0", -- 1AC8
         x"5d",  x"a5",  x"86",  x"da",  x"0f",  x"49",  x"83",  x"cd", -- 1AD0
         x"c8",  x"d6",  x"cd",  x"76",  x"da",  x"c1",  x"e1",  x"cd", -- 1AD8
         x"c8",  x"d6",  x"eb",  x"cd",  x"e0",  x"d6",  x"cd",  x"70", -- 1AE0
         x"da",  x"c3",  x"f3",  x"d5",  x"cd",  x"97",  x"d6",  x"fc", -- 1AE8
         x"1a",  x"d9",  x"fc",  x"c0",  x"d6",  x"3a",  x"e8",  x"03", -- 1AF0
         x"fe",  x"81",  x"da",  x"09",  x"db",  x"01",  x"00",  x"81", -- 1AF8
         x"51",  x"59",  x"cd",  x"f5",  x"d5",  x"21",  x"66",  x"d4", -- 1B00
         x"e5",  x"21",  x"13",  x"db",  x"cd",  x"ce",  x"d9",  x"21", -- 1B08
         x"ba",  x"da",  x"c9",  x"09",  x"4a",  x"d7",  x"3b",  x"78", -- 1B10
         x"02",  x"6e",  x"84",  x"7b",  x"fe",  x"c1",  x"2f",  x"7c", -- 1B18
         x"74",  x"31",  x"9a",  x"7d",  x"84",  x"3d",  x"5a",  x"7d", -- 1B20
         x"c8",  x"7f",  x"91",  x"7e",  x"e4",  x"bb",  x"4c",  x"7e", -- 1B28
         x"6c",  x"aa",  x"aa",  x"7f",  x"00",  x"00",  x"00",  x"81", -- 1B30
         x"cd",  x"49",  x"db",  x"28",  x"03",  x"cd",  x"6c",  x"c9", -- 1B38
         x"e5",  x"21",  x"47",  x"db",  x"e5",  x"eb",  x"e9",  x"e1", -- 1B40
         x"c9",  x"fe",  x"ae",  x"c0",  x"11",  x"00",  x"00",  x"cd", -- 1B48
         x"bd",  x"c8",  x"c8",  x"38",  x"0b",  x"fe",  x"94",  x"28", -- 1B50
         x"16",  x"fe",  x"47",  x"d2",  x"48",  x"c3",  x"d6",  x"07", -- 1B58
         x"d6",  x"30",  x"da",  x"48",  x"c3",  x"eb",  x"29",  x"29", -- 1B60
         x"29",  x"29",  x"b5",  x"6f",  x"eb",  x"18",  x"e0",  x"7b", -- 1B68
         x"87",  x"87",  x"87",  x"87",  x"f6",  x"0d",  x"57",  x"1e", -- 1B70
         x"ef",  x"18",  x"d4",  x"d5",  x"e5",  x"36",  x"00",  x"23", -- 1B78
         x"cd",  x"89",  x"c6",  x"20",  x"f8",  x"e3",  x"e5",  x"cd", -- 1B80
         x"fe",  x"d2",  x"cd",  x"09",  x"d2",  x"2a",  x"c4",  x"03", -- 1B88
         x"ed",  x"5b",  x"56",  x"03",  x"af",  x"ed",  x"52",  x"d1", -- 1B90
         x"e3",  x"ed",  x"52",  x"e5",  x"cd",  x"28",  x"dd",  x"4f", -- 1B98
         x"cd",  x"e4",  x"dd",  x"47",  x"e1",  x"cd",  x"e4",  x"dd", -- 1BA0
         x"12",  x"13",  x"2b",  x"7d",  x"b4",  x"20",  x"f6",  x"e1", -- 1BA8
         x"cd",  x"e4",  x"dd",  x"5f",  x"cd",  x"e4",  x"dd",  x"57", -- 1BB0
         x"af",  x"ed",  x"52",  x"38",  x"44",  x"2a",  x"56",  x"03", -- 1BB8
         x"23",  x"cd",  x"e4",  x"dd",  x"77",  x"23",  x"1b",  x"7b", -- 1BC0
         x"b2",  x"20",  x"f6",  x"d1",  x"e3",  x"c5",  x"cd",  x"f8", -- 1BC8
         x"dc",  x"e3",  x"ed",  x"42",  x"20",  x"2d",  x"e1",  x"cd", -- 1BD0
         x"77",  x"dd",  x"e3",  x"2b",  x"d5",  x"ed",  x"5b",  x"c4", -- 1BD8
         x"03",  x"ed",  x"b8",  x"ed",  x"53",  x"c4",  x"03",  x"e1", -- 1BE0
         x"42",  x"4b",  x"03",  x"d1",  x"2b",  x"70",  x"2b",  x"71", -- 1BE8
         x"2b",  x"35",  x"03",  x"20",  x"fc",  x"0b",  x"2b",  x"cd", -- 1BF0
         x"89",  x"c6",  x"20",  x"f0",  x"e1",  x"cd",  x"fd",  x"dd", -- 1BF8
         x"c9",  x"d1",  x"e1",  x"36",  x"00",  x"23",  x"cd",  x"89", -- 1C00
         x"c6",  x"20",  x"f8",  x"18",  x"29",  x"cd",  x"87",  x"dc", -- 1C08
         x"e5",  x"e2",  x"7b",  x"db",  x"eb",  x"ed",  x"52",  x"e5", -- 1C10
         x"cd",  x"28",  x"dd",  x"4f",  x"cd",  x"e4",  x"dd",  x"47", -- 1C18
         x"e1",  x"cd",  x"e4",  x"dd",  x"12",  x"13",  x"2b",  x"7d", -- 1C20
         x"b4",  x"20",  x"f6",  x"e1",  x"c5",  x"cd",  x"f8",  x"dc", -- 1C28
         x"e1",  x"ed",  x"42",  x"e1",  x"28",  x"c7",  x"cd",  x"1d", -- 1C30
         x"de",  x"21",  x"3f",  x"dc",  x"c3",  x"71",  x"c3",  x"42", -- 1C38
         x"41",  x"44",  x"00",  x"fe",  x"ae",  x"28",  x"c6",  x"cd", -- 1C40
         x"b0",  x"dc",  x"ed",  x"5b",  x"d7",  x"03",  x"1b",  x"1b", -- 1C48
         x"21",  x"00",  x"00",  x"39",  x"01",  x"d1",  x"ff",  x"ed", -- 1C50
         x"52",  x"09",  x"44",  x"4d",  x"cd",  x"28",  x"dd",  x"6f", -- 1C58
         x"cd",  x"e4",  x"dd",  x"67",  x"e5",  x"ed",  x"42",  x"e1", -- 1C60
         x"d2",  x"3e",  x"c3",  x"cd",  x"e4",  x"dd",  x"12",  x"13", -- 1C68
         x"2b",  x"7d",  x"b4",  x"20",  x"f6",  x"ed",  x"53",  x"d7", -- 1C70
         x"03",  x"21",  x"12",  x"c3",  x"cd",  x"c9",  x"d1",  x"c3", -- 1C78
         x"8a",  x"c4",  x"1e",  x"26",  x"c3",  x"56",  x"c3",  x"cd", -- 1C80
         x"ac",  x"dc",  x"e1",  x"cd",  x"cc",  x"c8",  x"3b",  x"3e", -- 1C88
         x"01",  x"32",  x"cc",  x"03",  x"cd",  x"06",  x"cf",  x"32", -- 1C90
         x"cc",  x"03",  x"e3",  x"e5",  x"60",  x"69",  x"eb",  x"19", -- 1C98
         x"eb",  x"4e",  x"06",  x"00",  x"09",  x"09",  x"23",  x"3a", -- 1CA0
         x"ae",  x"03",  x"b7",  x"c9",  x"3e",  x"d4",  x"23",  x"01", -- 1CA8
         x"3e",  x"d3",  x"f5",  x"3a",  x"5d",  x"03",  x"a7",  x"3e", -- 1CB0
         x"00",  x"32",  x"5d",  x"03",  x"28",  x"04",  x"f1",  x"c6", -- 1CB8
         x"04",  x"f5",  x"cd",  x"be",  x"c8",  x"cd",  x"3a",  x"cd", -- 1CC0
         x"f1",  x"e3",  x"e5",  x"f5",  x"cd",  x"3f",  x"d3",  x"21", -- 1CC8
         x"f7",  x"03",  x"06",  x"0d",  x"2b",  x"36",  x"20",  x"10", -- 1CD0
         x"fb",  x"d5",  x"11",  x"82",  x"dc",  x"73",  x"23",  x"72", -- 1CD8
         x"d1",  x"23",  x"f1",  x"77",  x"23",  x"77",  x"23",  x"77", -- 1CE0
         x"23",  x"eb",  x"06",  x"00",  x"79",  x"fe",  x"09",  x"38", -- 1CE8
         x"04",  x"0d",  x"23",  x"18",  x"f7",  x"ed",  x"b0",  x"c9", -- 1CF0
         x"e5",  x"af",  x"47",  x"86",  x"cd",  x"03",  x"dd",  x"20", -- 1CF8
         x"fa",  x"e1",  x"c9",  x"4f",  x"30",  x"01",  x"04",  x"23", -- 1D00
         x"cd",  x"89",  x"c6",  x"79",  x"c9",  x"f5",  x"3a",  x"07", -- 1D08
         x"03",  x"cb",  x"4f",  x"cb",  x"cf",  x"32",  x"07",  x"03", -- 1D10
         x"3e",  x"13",  x"20",  x"02",  x"c6",  x"08",  x"32",  x"08", -- 1D18
         x"03",  x"21",  x"ea",  x"03",  x"f1",  x"c3",  x"d5",  x"dd", -- 1D20
         x"3a",  x"07",  x"03",  x"cb",  x"47",  x"cb",  x"c7",  x"32", -- 1D28
         x"07",  x"03",  x"3e",  x"12",  x"20",  x"02",  x"c6",  x"08", -- 1D30
         x"32",  x"09",  x"03",  x"21",  x"ea",  x"03",  x"c3",  x"e4", -- 1D38
         x"dd",  x"fe",  x"ae",  x"28",  x"24",  x"cd",  x"97",  x"c6", -- 1D40
         x"cd",  x"b0",  x"dc",  x"2a",  x"d7",  x"03",  x"11",  x"ff", -- 1D48
         x"fb",  x"19",  x"44",  x"4d",  x"11",  x"01",  x"04",  x"cd", -- 1D50
         x"b5",  x"dd",  x"e1",  x"e5",  x"21",  x"07",  x"03",  x"cb", -- 1D58
         x"8e",  x"11",  x"43",  x"03",  x"cd",  x"f6",  x"df",  x"e1", -- 1D60
         x"c9",  x"cd",  x"87",  x"dc",  x"e2",  x"89",  x"dd",  x"cd", -- 1D68
         x"f8",  x"dc",  x"eb",  x"ed",  x"52",  x"18",  x"e0",  x"e5", -- 1D70
         x"01",  x"00",  x"00",  x"7e",  x"23",  x"77",  x"34",  x"81", -- 1D78
         x"23",  x"23",  x"cd",  x"03",  x"dd",  x"20",  x"f4",  x"e1", -- 1D80
         x"c9",  x"cd",  x"77",  x"dd",  x"c5",  x"cd",  x"f8",  x"dc", -- 1D88
         x"eb",  x"ed",  x"52",  x"cd",  x"b5",  x"dd",  x"c1",  x"79", -- 1D90
         x"cd",  x"d5",  x"dd",  x"78",  x"eb",  x"cd",  x"d5",  x"dd", -- 1D98
         x"2b",  x"2b",  x"78",  x"b1",  x"28",  x"b4",  x"56",  x"2b", -- 1DA0
         x"5e",  x"2b",  x"35",  x"28",  x"f3",  x"1a",  x"cd",  x"d5", -- 1DA8
         x"dd",  x"13",  x"0b",  x"18",  x"f5",  x"23",  x"e5",  x"79", -- 1DB0
         x"cd",  x"0d",  x"dd",  x"78",  x"e1",  x"cd",  x"d5",  x"dd", -- 1DB8
         x"2b",  x"7d",  x"b4",  x"1a",  x"13",  x"20",  x"f6",  x"c9", -- 1DC0
         x"3a",  x"08",  x"03",  x"e6",  x"07",  x"d6",  x"01",  x"c9", -- 1DC8
         x"cd",  x"1d",  x"de",  x"3e",  x"0c",  x"f5",  x"d5",  x"57", -- 1DD0
         x"3a",  x"08",  x"03",  x"5f",  x"7a",  x"cd",  x"f6",  x"df", -- 1DD8
         x"7b",  x"d1",  x"18",  x"3c",  x"d5",  x"3a",  x"09",  x"03", -- 1DE0
         x"5f",  x"cd",  x"f6",  x"df",  x"7b",  x"32",  x"09",  x"03", -- 1DE8
         x"7a",  x"18",  x"06",  x"d5",  x"1e",  x"80",  x"cd",  x"f6", -- 1DF0
         x"df",  x"cb",  x"7b",  x"d1",  x"c9",  x"f5",  x"e5",  x"d5", -- 1DF8
         x"c5",  x"11",  x"42",  x"03",  x"06",  x"06",  x"7a",  x"21", -- 1E00
         x"07",  x"03",  x"cb",  x"3e",  x"dc",  x"f6",  x"df",  x"1c", -- 1E08
         x"10",  x"f8",  x"c1",  x"d1",  x"e1",  x"3e",  x"f5",  x"3e", -- 1E10
         x"00",  x"32",  x"09",  x"03",  x"3e",  x"f5",  x"3e",  x"01", -- 1E18
         x"32",  x"08",  x"03",  x"f1",  x"c9",  x"7e",  x"fe",  x"23", -- 1E20
         x"20",  x"31",  x"cd",  x"bd",  x"c8",  x"30",  x"38",  x"23", -- 1E28
         x"e5",  x"e6",  x"03",  x"28",  x"12",  x"21",  x"07",  x"03", -- 1E30
         x"87",  x"fe",  x"04",  x"28",  x"12",  x"30",  x"16",  x"cb", -- 1E38
         x"4e",  x"cb",  x"ce",  x"20",  x"02",  x"c6",  x"08",  x"3c", -- 1E40
         x"32",  x"08",  x"03",  x"e1",  x"c3",  x"be",  x"c8",  x"cb", -- 1E48
         x"5e",  x"cb",  x"de",  x"18",  x"ee",  x"cb",  x"6e",  x"cb", -- 1E50
         x"ee",  x"18",  x"e8",  x"e5",  x"af",  x"18",  x"e8",  x"7e", -- 1E58
         x"fe",  x"23",  x"20",  x"30",  x"cd",  x"bd",  x"c8",  x"d2", -- 1E60
         x"48",  x"c3",  x"23",  x"e5",  x"e6",  x"03",  x"28",  x"12", -- 1E68
         x"21",  x"07",  x"03",  x"87",  x"fe",  x"04",  x"28",  x"10", -- 1E70
         x"38",  x"14",  x"cb",  x"66",  x"cb",  x"e6",  x"20",  x"02", -- 1E78
         x"c6",  x"08",  x"32",  x"09",  x"03",  x"e1",  x"18",  x"c4", -- 1E80
         x"cb",  x"56",  x"cb",  x"d6",  x"18",  x"f0",  x"cb",  x"46", -- 1E88
         x"cb",  x"c6",  x"18",  x"ea",  x"e5",  x"af",  x"18",  x"ea", -- 1E90
         x"c5",  x"cd",  x"2a",  x"d8",  x"e1",  x"23",  x"23",  x"23", -- 1E98
         x"23",  x"01",  x"61",  x"03",  x"c5",  x"18",  x"03",  x"cd", -- 1EA0
         x"d7",  x"de",  x"7e",  x"23",  x"fe",  x"22",  x"28",  x"16", -- 1EA8
         x"b7",  x"28",  x"1f",  x"f2",  x"a7",  x"de",  x"c5",  x"cd", -- 1EB0
         x"9a",  x"c7",  x"c1",  x"cd",  x"d7",  x"de",  x"1a",  x"13", -- 1EB8
         x"b7",  x"f2",  x"bb",  x"de",  x"18",  x"e4",  x"cd",  x"d7", -- 1EC0
         x"de",  x"7e",  x"23",  x"fe",  x"22",  x"28",  x"d8",  x"b7", -- 1EC8
         x"20",  x"f4",  x"3e",  x"20",  x"03",  x"18",  x"0c",  x"03", -- 1ED0
         x"02",  x"e5",  x"21",  x"56",  x"fc",  x"09",  x"e1",  x"d0", -- 1ED8
         x"e1",  x"3e",  x"2a",  x"cd",  x"d5",  x"dd",  x"af",  x"02", -- 1EE0
         x"e1",  x"77",  x"23",  x"e5",  x"cd",  x"f1",  x"c5",  x"d1", -- 1EE8
         x"23",  x"36",  x"00",  x"2b",  x"36",  x"20",  x"cd",  x"e4", -- 1EF0
         x"dd",  x"fe",  x"0a",  x"20",  x"05",  x"cd",  x"12",  x"df", -- 1EF8
         x"3c",  x"c9",  x"cd",  x"0f",  x"df",  x"c8",  x"cd",  x"27", -- 1F00
         x"df",  x"d8",  x"cd",  x"32",  x"df",  x"18",  x"e7",  x"fe", -- 1F08
         x"0d",  x"c0",  x"3e",  x"09",  x"cd",  x"d5",  x"dd",  x"23", -- 1F10
         x"7e",  x"b7",  x"20",  x"f6",  x"2b",  x"7e",  x"fe",  x"20", -- 1F18
         x"20",  x"02",  x"36",  x"00",  x"c3",  x"5e",  x"cb",  x"fe", -- 1F20
         x"03",  x"28",  x"02",  x"a7",  x"c9",  x"cd",  x"12",  x"df", -- 1F28
         x"37",  x"c9",  x"fe",  x"08",  x"28",  x"44",  x"fe",  x"09", -- 1F30
         x"28",  x"2a",  x"fe",  x"1f",  x"28",  x"47",  x"fe",  x"19", -- 1F38
         x"ca",  x"c5",  x"df",  x"fe",  x"18",  x"ca",  x"cf",  x"df", -- 1F40
         x"fe",  x"02",  x"ca",  x"db",  x"df",  x"fe",  x"1a",  x"28", -- 1F48
         x"48",  x"fe",  x"0b",  x"c8",  x"fe",  x"0a",  x"c8",  x"fe", -- 1F50
         x"01",  x"c8",  x"fe",  x"20",  x"30",  x"05",  x"3f",  x"cd", -- 1F58
         x"d5",  x"dd",  x"c9",  x"77",  x"cd",  x"d5",  x"dd",  x"23", -- 1F60
         x"7e",  x"b7",  x"c0",  x"11",  x"ab",  x"03",  x"cd",  x"89", -- 1F68
         x"c6",  x"28",  x"07",  x"36",  x"20",  x"23",  x"36",  x"00", -- 1F70
         x"18",  x"03",  x"cd",  x"a2",  x"c6",  x"2b",  x"7e",  x"b7", -- 1F78
         x"c0",  x"3e",  x"09",  x"18",  x"df",  x"e5",  x"23",  x"cd", -- 1F80
         x"f1",  x"c5",  x"cd",  x"a9",  x"c6",  x"d1",  x"af",  x"2b", -- 1F88
         x"46",  x"77",  x"cd",  x"a2",  x"c6",  x"78",  x"20",  x"f7", -- 1F90
         x"c9",  x"cd",  x"a9",  x"c6",  x"e5",  x"cd",  x"f1",  x"c5", -- 1F98
         x"11",  x"ab",  x"03",  x"cd",  x"89",  x"c6",  x"20",  x"0c", -- 1FA0
         x"cd",  x"a2",  x"c6",  x"cd",  x"a9",  x"c6",  x"cd",  x"a2", -- 1FA8
         x"c6",  x"2b",  x"36",  x"00",  x"d1",  x"44",  x"4d",  x"03", -- 1FB0
         x"7e",  x"02",  x"0b",  x"cd",  x"a2",  x"c6",  x"2b",  x"20", -- 1FB8
         x"f7",  x"23",  x"36",  x"20",  x"c9",  x"cd",  x"a2",  x"c6", -- 1FC0
         x"2b",  x"7e",  x"b7",  x"20",  x"f8",  x"18",  x"b2",  x"3e", -- 1FC8
         x"09",  x"cd",  x"d5",  x"dd",  x"23",  x"7e",  x"b7",  x"20", -- 1FD0
         x"f6",  x"18",  x"90",  x"cd",  x"c5",  x"df",  x"e5",  x"7e", -- 1FD8
         x"b7",  x"28",  x"05",  x"36",  x"20",  x"23",  x"18",  x"f7", -- 1FE0
         x"e1",  x"cd",  x"f1",  x"c5",  x"cd",  x"c5",  x"df",  x"23", -- 1FE8
         x"36",  x"00",  x"2b",  x"c9",  x"1e",  x"ff",  x"c3",  x"0e", -- 1FF0
         x"e0",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1FF8
         x"ff",  x"ff",  x"ff",  x"c3",  x"d2",  x"e0",  x"c3",  x"f3", -- 2000
         x"e0",  x"c3",  x"57",  x"e1",  x"11",  x"e0",  x"c3",  x"00", -- 2008
         x"e6",  x"c9",  x"4e",  x"4b",  x"45",  x"59",  x"24",  x"ca", -- 2010
         x"4f",  x"59",  x"53",  x"54",  x"d3",  x"54",  x"52",  x"49", -- 2018
         x"4e",  x"47",  x"24",  x"c9",  x"4e",  x"53",  x"54",  x"52", -- 2020
         x"d2",  x"45",  x"4e",  x"55",  x"4d",  x"c4",  x"45",  x"4c", -- 2028
         x"45",  x"54",  x"45",  x"d0",  x"41",  x"55",  x"53",  x"45", -- 2030
         x"c2",  x"45",  x"45",  x"50",  x"d7",  x"49",  x"4e",  x"44", -- 2038
         x"4f",  x"57",  x"c2",  x"4f",  x"52",  x"44",  x"45",  x"52", -- 2040
         x"c9",  x"4e",  x"4b",  x"d0",  x"41",  x"50",  x"45",  x"52", -- 2048
         x"c1",  x"54",  x"d0",  x"53",  x"45",  x"54",  x"cc",  x"49", -- 2050
         x"4e",  x"45",  x"c3",  x"49",  x"52",  x"43",  x"4c",  x"45", -- 2058
         x"a1",  x"d0",  x"41",  x"49",  x"4e",  x"54",  x"cc",  x"41", -- 2060
         x"42",  x"45",  x"4c",  x"d3",  x"49",  x"5a",  x"45",  x"da", -- 2068
         x"45",  x"52",  x"4f",  x"c8",  x"4f",  x"4d",  x"45",  x"a1", -- 2070
         x"c7",  x"43",  x"4c",  x"53",  x"d3",  x"43",  x"41",  x"4c", -- 2078
         x"45",  x"d3",  x"43",  x"52",  x"45",  x"45",  x"4e",  x"d0", -- 2080
         x"4f",  x"49",  x"4e",  x"54",  x"d8",  x"50",  x"4f",  x"53", -- 2088
         x"a1",  x"d9",  x"50",  x"4f",  x"53",  x"80",  x"19",  x"e4", -- 2090
         x"f5",  x"e4",  x"3c",  x"e4",  x"c1",  x"e4",  x"f8",  x"e1", -- 2098
         x"cd",  x"e5",  x"a7",  x"e3",  x"34",  x"e4",  x"b5",  x"e1", -- 20A0
         x"79",  x"e1",  x"7d",  x"e1",  x"7e",  x"e1",  x"17",  x"e5", -- 20A8
         x"d6",  x"a7",  x"d9",  x"a7",  x"dc",  x"a7",  x"4a",  x"ca", -- 20B0
         x"df",  x"a7",  x"e2",  x"a7",  x"e5",  x"a7",  x"e8",  x"a7", -- 20B8
         x"eb",  x"a7",  x"4a",  x"ca",  x"ee",  x"a7",  x"f1",  x"a7", -- 20C0
         x"f4",  x"a7",  x"f7",  x"a7",  x"fa",  x"a7",  x"4a",  x"ca", -- 20C8
         x"fd",  x"a7",  x"78",  x"d6",  x"09",  x"38",  x"6d",  x"fe", -- 20D0
         x"09",  x"38",  x"07",  x"cd",  x"f1",  x"e5",  x"fe",  x"16", -- 20D8
         x"30",  x"62",  x"07",  x"4f",  x"06",  x"00",  x"eb",  x"21", -- 20E0
         x"9e",  x"e0",  x"09",  x"4e",  x"23",  x"46",  x"c5",  x"eb", -- 20E8
         x"c3",  x"bd",  x"c8",  x"7e",  x"fe",  x"df",  x"d8",  x"fe", -- 20F0
         x"e2",  x"d0",  x"fe",  x"e1",  x"ca",  x"17",  x"e5",  x"3a", -- 20F8
         x"fd",  x"03",  x"a7",  x"20",  x"3f",  x"3c",  x"32",  x"fd", -- 2100
         x"03",  x"3a",  x"27",  x"00",  x"f5",  x"7e",  x"fe",  x"df", -- 2108
         x"28",  x"0d",  x"cd",  x"bd",  x"c8",  x"cd",  x"7e",  x"e1", -- 2110
         x"7e",  x"fe",  x"3b",  x"28",  x"35",  x"18",  x"25",  x"cd", -- 2118
         x"bd",  x"c8",  x"cd",  x"7d",  x"e1",  x"7e",  x"fe",  x"3b", -- 2120
         x"28",  x"28",  x"cd",  x"d6",  x"c8",  x"fe",  x"e0",  x"20", -- 2128
         x"13",  x"cd",  x"bd",  x"c8",  x"cd",  x"7e",  x"e1",  x"cd", -- 2130
         x"cc",  x"c8",  x"3b",  x"cd",  x"03",  x"cb",  x"f1",  x"32", -- 2138
         x"27",  x"00",  x"c1",  x"c9",  x"3e",  x"e2",  x"d3",  x"b8", -- 2140
         x"c3",  x"48",  x"c3",  x"3e",  x"e2",  x"d3",  x"b8",  x"c3", -- 2148
         x"67",  x"c9",  x"cd",  x"bd",  x"c8",  x"18",  x"e4",  x"79", -- 2150
         x"d6",  x"3e",  x"38",  x"e8",  x"fe",  x"07",  x"38",  x"0b", -- 2158
         x"cd",  x"f1",  x"e5",  x"fe",  x"32",  x"38",  x"dd",  x"fe", -- 2160
         x"3b",  x"30",  x"d9",  x"eb",  x"01",  x"96",  x"e0",  x"e1", -- 2168
         x"6f",  x"09",  x"4e",  x"23",  x"66",  x"69",  x"e5",  x"eb", -- 2170
         x"c9",  x"3e",  x"01",  x"18",  x"02",  x"f6",  x"af",  x"f5", -- 2178
         x"cd",  x"21",  x"d4",  x"fe",  x"01",  x"38",  x"6e",  x"fe", -- 2180
         x"09",  x"30",  x"6a",  x"3d",  x"4f",  x"f1",  x"b7",  x"28", -- 2188
         x"0b",  x"cb",  x"21",  x"cb",  x"21",  x"cb",  x"21",  x"3d", -- 2190
         x"28",  x"17",  x"cb",  x"21",  x"41",  x"b7",  x"3a",  x"27", -- 2198
         x"00",  x"28",  x"0a",  x"e6",  x"07",  x"b0",  x"32",  x"27", -- 21A0
         x"00",  x"32",  x"28",  x"00",  x"c9",  x"e6",  x"70",  x"18", -- 21A8
         x"f4",  x"79",  x"d3",  x"88",  x"c9",  x"0e",  x"1d",  x"cd", -- 21B0
         x"05",  x"00",  x"cd",  x"be",  x"c8",  x"28",  x"2d",  x"cd", -- 21B8
         x"f7",  x"e7",  x"f5",  x"cd",  x"f7",  x"e7",  x"f5",  x"cd", -- 21C0
         x"f7",  x"e7",  x"f5",  x"cd",  x"21",  x"d4",  x"3c",  x"3c", -- 21C8
         x"57",  x"fe",  x"2a",  x"30",  x"20",  x"f1",  x"5f",  x"f1", -- 21D0
         x"3c",  x"3c",  x"47",  x"fe",  x"1a",  x"30",  x"16",  x"f1", -- 21D8
         x"4f",  x"3c",  x"b8",  x"30",  x"10",  x"7b",  x"3c",  x"ba", -- 21E0
         x"30",  x"0b",  x"18",  x"06",  x"01",  x"00",  x"19",  x"11", -- 21E8
         x"00",  x"29",  x"c3",  x"e6",  x"e7",  x"c3",  x"4b",  x"e1", -- 21F0
         x"01",  x"0a",  x"00",  x"c5",  x"50",  x"58",  x"28",  x"27", -- 21F8
         x"fe",  x"2c",  x"28",  x"09",  x"d5",  x"cd",  x"86",  x"c9", -- 2200
         x"42",  x"4b",  x"d1",  x"28",  x"1a",  x"cd",  x"d6",  x"c8", -- 2208
         x"cd",  x"86",  x"c9",  x"28",  x"12",  x"f1",  x"cd",  x"d6", -- 2210
         x"c8",  x"d5",  x"cd",  x"86",  x"c9",  x"c2",  x"44",  x"e1", -- 2218
         x"7a",  x"b3",  x"28",  x"d1",  x"eb",  x"e3",  x"eb",  x"d5", -- 2220
         x"c5",  x"cd",  x"bb",  x"c4",  x"d1",  x"d5",  x"c5",  x"cd", -- 2228
         x"bb",  x"c4",  x"60",  x"69",  x"d1",  x"cd",  x"89",  x"c6", -- 2230
         x"eb",  x"38",  x"ba",  x"d1",  x"f1",  x"c1",  x"d5",  x"f5", -- 2238
         x"18",  x"0e",  x"09",  x"38",  x"f4",  x"eb",  x"e5",  x"21", -- 2240
         x"f9",  x"ff",  x"cd",  x"89",  x"c6",  x"e1",  x"38",  x"e9", -- 2248
         x"d5",  x"5e",  x"23",  x"56",  x"7a",  x"b3",  x"eb",  x"d1", -- 2250
         x"28",  x"07",  x"7e",  x"23",  x"b6",  x"2b",  x"eb",  x"20", -- 2258
         x"e1",  x"c5",  x"0e",  x"80",  x"cd",  x"27",  x"c3",  x"af", -- 2260
         x"cd",  x"9a",  x"e2",  x"af",  x"3c",  x"cd",  x"9a",  x"e2", -- 2268
         x"c1",  x"d1",  x"c5",  x"cd",  x"bb",  x"c4",  x"60",  x"69", -- 2270
         x"c1",  x"d1",  x"f1",  x"d5",  x"5e",  x"23",  x"56",  x"7a", -- 2278
         x"b3",  x"28",  x"0d",  x"eb",  x"e3",  x"eb",  x"23",  x"73", -- 2280
         x"23",  x"72",  x"eb",  x"09",  x"eb",  x"e1",  x"18",  x"eb", -- 2288
         x"3d",  x"cd",  x"9a",  x"e2",  x"01",  x"8a",  x"c4",  x"c5", -- 2290
         x"3e",  x"02",  x"32",  x"4e",  x"03",  x"2a",  x"5f",  x"03", -- 2298
         x"2b",  x"c5",  x"c5",  x"23",  x"c1",  x"c1",  x"44",  x"4d", -- 22A0
         x"5e",  x"23",  x"56",  x"7a",  x"b3",  x"c8",  x"c5",  x"d5", -- 22A8
         x"23",  x"23",  x"cd",  x"bd",  x"c8",  x"b7",  x"28",  x"eb", -- 22B0
         x"4f",  x"3a",  x"4e",  x"03",  x"b7",  x"79",  x"28",  x"5f", -- 22B8
         x"fe",  x"0d",  x"20",  x"ee",  x"e5",  x"e5",  x"23",  x"5e", -- 22C0
         x"23",  x"56",  x"3a",  x"4e",  x"03",  x"3d",  x"28",  x"7e", -- 22C8
         x"3d",  x"28",  x"0e",  x"eb",  x"23",  x"23",  x"1b",  x"ed", -- 22D0
         x"a0",  x"ed",  x"a0",  x"eb",  x"d1",  x"d1",  x"2b",  x"18", -- 22D8
         x"d1",  x"d5",  x"eb",  x"13",  x"2a",  x"d7",  x"03",  x"ed", -- 22E0
         x"52",  x"44",  x"4d",  x"e1",  x"e3",  x"eb",  x"c5",  x"ed", -- 22E8
         x"b0",  x"c1",  x"d1",  x"e1",  x"e5",  x"c5",  x"af",  x"06", -- 22F0
         x"98",  x"cd",  x"ae",  x"d6",  x"cd",  x"34",  x"d8",  x"c1", -- 22F8
         x"d1",  x"23",  x"7e",  x"eb",  x"2b",  x"b7",  x"28",  x"aa", -- 2300
         x"23",  x"eb",  x"c5",  x"e5",  x"eb",  x"09",  x"54",  x"5d", -- 2308
         x"13",  x"ed",  x"53",  x"d7",  x"03",  x"1b",  x"2b",  x"ed", -- 2310
         x"b8",  x"e1",  x"ed",  x"a0",  x"c1",  x"18",  x"e3",  x"fe", -- 2318
         x"88",  x"28",  x"19",  x"fe",  x"8c",  x"28",  x"15",  x"fe", -- 2320
         x"8b",  x"28",  x"11",  x"fe",  x"d4",  x"28",  x"0d",  x"fe", -- 2328
         x"da",  x"28",  x"09",  x"fe",  x"d3",  x"28",  x"05",  x"fe", -- 2330
         x"a9",  x"c2",  x"b2",  x"e2",  x"cd",  x"87",  x"c9",  x"e5", -- 2338
         x"cd",  x"bb",  x"c4",  x"e1",  x"38",  x"14",  x"7e",  x"fe", -- 2340
         x"2c",  x"28",  x"f1",  x"2b",  x"18",  x"eb",  x"cd",  x"bb", -- 2348
         x"c4",  x"e1",  x"23",  x"71",  x"23",  x"70",  x"d1",  x"c3", -- 2350
         x"b2",  x"e2",  x"d5",  x"eb",  x"2a",  x"d7",  x"03",  x"ed", -- 2358
         x"52",  x"23",  x"e5",  x"c1",  x"62",  x"6b",  x"1b",  x"1a", -- 2360
         x"fe",  x"2c",  x"28",  x"10",  x"fe",  x"3a",  x"30",  x"0c", -- 2368
         x"f1",  x"e3",  x"2b",  x"e3",  x"f5",  x"c5",  x"d5",  x"ed", -- 2370
         x"b0",  x"d1",  x"18",  x"e7",  x"eb",  x"09",  x"54",  x"5d", -- 2378
         x"13",  x"13",  x"13",  x"13",  x"ed",  x"53",  x"d7",  x"03", -- 2380
         x"1b",  x"ed",  x"b8",  x"3e",  x"0d",  x"23",  x"77",  x"23", -- 2388
         x"d1",  x"73",  x"23",  x"72",  x"d1",  x"e3",  x"13",  x"13", -- 2390
         x"13",  x"73",  x"23",  x"72",  x"2b",  x"e3",  x"d5",  x"e5", -- 2398
         x"cd",  x"93",  x"c4",  x"e1",  x"23",  x"18",  x"9f",  x"cd", -- 23A0
         x"be",  x"c8",  x"20",  x"11",  x"cd",  x"f3",  x"dd",  x"20", -- 23A8
         x"fb",  x"fe",  x"03",  x"28",  x"07",  x"fe",  x"1e",  x"20", -- 23B0
         x"f3",  x"cd",  x"e4",  x"dd",  x"c9",  x"cd",  x"5e",  x"c9", -- 23B8
         x"7a",  x"b3",  x"c8",  x"e5",  x"21",  x"01",  x"00",  x"dd", -- 23C0
         x"21",  x"0b",  x"e4",  x"3e",  x"05",  x"0e",  x"8d",  x"06", -- 23C8
         x"0a",  x"dd",  x"86",  x"00",  x"10",  x"fb",  x"0d",  x"20", -- 23D0
         x"f6",  x"3d",  x"20",  x"f1",  x"a7",  x"eb",  x"ed",  x"52", -- 23D8
         x"eb",  x"28",  x"1b",  x"f5",  x"c5",  x"d5",  x"cd",  x"f3", -- 23E0
         x"dd",  x"20",  x"08",  x"fe",  x"1e",  x"28",  x"09",  x"fe", -- 23E8
         x"03",  x"28",  x"08",  x"d1",  x"c1",  x"f1",  x"18",  x"cf", -- 23F0
         x"cd",  x"e4",  x"dd",  x"d1",  x"c1",  x"f1",  x"e1",  x"c9", -- 23F8
         x"c3",  x"0d",  x"c0",  x"42",  x"41",  x"53",  x"49",  x"43", -- 2400
         x"20",  x"20",  x"20",  x"00",  x"c3",  x"8c",  x"c0",  x"57", -- 2408
         x"42",  x"41",  x"53",  x"49",  x"43",  x"20",  x"20",  x"00", -- 2410
         x"00",  x"e5",  x"cd",  x"f3",  x"dd",  x"20",  x"0f",  x"3e", -- 2418
         x"01",  x"cd",  x"7b",  x"d1",  x"cd",  x"e4",  x"dd",  x"2a", -- 2420
         x"c2",  x"03",  x"77",  x"c3",  x"a9",  x"d1",  x"af",  x"cd", -- 2428
         x"7b",  x"d1",  x"18",  x"f7",  x"0e",  x"02",  x"1e",  x"07", -- 2430
         x"cd",  x"05",  x"00",  x"c9",  x"cd",  x"cc",  x"c8",  x"28", -- 2438
         x"cd",  x"f7",  x"e7",  x"f5",  x"cd",  x"8e",  x"e4",  x"f5", -- 2440
         x"cd",  x"db",  x"c8",  x"f1",  x"e3",  x"44",  x"e5",  x"f5", -- 2448
         x"d5",  x"4f",  x"af",  x"b9",  x"28",  x"0c",  x"b8",  x"28", -- 2450
         x"09",  x"79",  x"05",  x"28",  x"05",  x"81",  x"38",  x"29", -- 2458
         x"10",  x"fb",  x"47",  x"0e",  x"00",  x"cd",  x"e1",  x"d1", -- 2460
         x"c1",  x"c5",  x"cd",  x"7e",  x"d1",  x"e1",  x"e3",  x"7c", -- 2468
         x"e1",  x"e3",  x"6f",  x"24",  x"25",  x"e5",  x"c5",  x"28", -- 2470
         x"07",  x"cd",  x"f2",  x"d2",  x"c1",  x"e1",  x"18",  x"f4", -- 2478
         x"c1",  x"e1",  x"d1",  x"cd",  x"02",  x"d3",  x"c3",  x"a9", -- 2480
         x"d1",  x"1e",  x"1c",  x"c3",  x"56",  x"c3",  x"cd",  x"3a", -- 2488
         x"cd",  x"e5",  x"cd",  x"30",  x"d3",  x"23",  x"23",  x"5e", -- 2490
         x"23",  x"56",  x"e1",  x"c9",  x"23",  x"e5",  x"2b",  x"0d", -- 2498
         x"c5",  x"0c",  x"13",  x"05",  x"28",  x"11",  x"23",  x"0d", -- 24A0
         x"28",  x"09",  x"1a",  x"be",  x"28",  x"f4",  x"c1",  x"e1", -- 24A8
         x"d1",  x"18",  x"2c",  x"e1",  x"e1",  x"18",  x"31",  x"d1", -- 24B0
         x"e1",  x"d1",  x"d1",  x"a7",  x"ed",  x"52",  x"7d",  x"18", -- 24B8
         x"2a",  x"cd",  x"cc",  x"c8",  x"28",  x"cd",  x"8e",  x"e4", -- 24C0
         x"d5",  x"f5",  x"cd",  x"d6",  x"c8",  x"cd",  x"8e",  x"e4", -- 24C8
         x"f5",  x"cd",  x"db",  x"c8",  x"f1",  x"28",  x"1a",  x"4f", -- 24D0
         x"f1",  x"28",  x"6d",  x"47",  x"e3",  x"eb",  x"e5",  x"d5", -- 24D8
         x"1a",  x"be",  x"28",  x"b8",  x"23",  x"0d",  x"20",  x"f9", -- 24E0
         x"af",  x"e1",  x"e1",  x"11",  x"f3",  x"cd",  x"d5",  x"18", -- 24E8
         x"23",  x"d1",  x"e3",  x"18",  x"f6",  x"cd",  x"e1",  x"cd", -- 24F0
         x"e5",  x"11",  x"f3",  x"cd",  x"d5",  x"cd",  x"24",  x"d4", -- 24F8
         x"a7",  x"28",  x"45",  x"fe",  x"03",  x"30",  x"41",  x"0e", -- 2500
         x"06",  x"cd",  x"05",  x"00",  x"38",  x"3a",  x"fe",  x"01", -- 2508
         x"28",  x"01",  x"48",  x"79",  x"c3",  x"c0",  x"d0",  x"3a", -- 2510
         x"fd",  x"03",  x"cb",  x"4f",  x"cb",  x"cf",  x"32",  x"fd", -- 2518
         x"03",  x"20",  x"25",  x"cd",  x"bd",  x"c8",  x"cd",  x"cc", -- 2520
         x"c8",  x"28",  x"cd",  x"f7",  x"e7",  x"f5",  x"cd",  x"21", -- 2528
         x"d4",  x"f5",  x"cd",  x"db",  x"c8",  x"cd",  x"cc",  x"c8", -- 2530
         x"3b",  x"f1",  x"4f",  x"f1",  x"e5",  x"47",  x"78",  x"fe", -- 2538
         x"18",  x"30",  x"05",  x"79",  x"fe",  x"28",  x"38",  x"03", -- 2540
         x"c3",  x"4b",  x"e1",  x"2e",  x"00",  x"65",  x"55",  x"1e", -- 2548
         x"28",  x"04",  x"05",  x"28",  x"03",  x"19",  x"10",  x"fd", -- 2550
         x"59",  x"19",  x"11",  x"00",  x"ec",  x"19",  x"54",  x"5d", -- 2558
         x"01",  x"00",  x"fc",  x"09",  x"e3",  x"d5",  x"fe",  x"d5", -- 2560
         x"38",  x"09",  x"3a",  x"fc",  x"03",  x"a7",  x"28",  x"03", -- 2568
         x"cd",  x"06",  x"e0",  x"cd",  x"3a",  x"cd",  x"e5",  x"3a", -- 2570
         x"ae",  x"03",  x"b7",  x"20",  x"0c",  x"cd",  x"34",  x"d8", -- 2578
         x"cd",  x"8a",  x"d1",  x"36",  x"20",  x"2a",  x"e5",  x"03", -- 2580
         x"34",  x"cd",  x"fe",  x"d2",  x"cd",  x"ee",  x"d6",  x"e1", -- 2588
         x"dd",  x"e1",  x"fd",  x"e1",  x"3a",  x"27",  x"00",  x"57", -- 2590
         x"1c",  x"1d",  x"28",  x"13",  x"0a",  x"cd",  x"bf",  x"e5", -- 2598
         x"30",  x"0d",  x"dd",  x"77",  x"00",  x"fd",  x"72",  x"00", -- 25A0
         x"dd",  x"23",  x"fd",  x"23",  x"03",  x"18",  x"ea",  x"cd", -- 25A8
         x"be",  x"c8",  x"20",  x"02",  x"c1",  x"c9",  x"cd",  x"d6", -- 25B0
         x"c8",  x"fd",  x"e5",  x"dd",  x"e5",  x"18",  x"a7",  x"e5", -- 25B8
         x"dd",  x"e5",  x"e1",  x"d5",  x"11",  x"c0",  x"ef",  x"a7", -- 25C0
         x"ed",  x"52",  x"d1",  x"e1",  x"c9",  x"c8",  x"cd",  x"86", -- 25C8
         x"c9",  x"ca",  x"42",  x"c4",  x"cd",  x"d6",  x"c8",  x"d5", -- 25D0
         x"cd",  x"86",  x"c9",  x"e1",  x"c0",  x"eb",  x"e5",  x"cd", -- 25D8
         x"bb",  x"c4",  x"d2",  x"4d",  x"c4",  x"d1",  x"f5",  x"c5", -- 25E0
         x"cd",  x"be",  x"c4",  x"30",  x"f5",  x"c1",  x"c3",  x"50", -- 25E8
         x"c4",  x"47",  x"e5",  x"2a",  x"b0",  x"e0",  x"3e",  x"c3", -- 25F0
         x"be",  x"78",  x"e1",  x"c8",  x"c3",  x"44",  x"e1",  x"ff", -- 25F8
         x"cb",  x"6b",  x"c2",  x"00",  x"00",  x"22",  x"77",  x"00", -- 2600
         x"e5",  x"c5",  x"21",  x"1e",  x"e6",  x"e5",  x"7b",  x"e6", -- 2608
         x"07",  x"17",  x"4f",  x"06",  x"00",  x"21",  x"42",  x"e6", -- 2610
         x"09",  x"7e",  x"23",  x"66",  x"6f",  x"e9",  x"c1",  x"e1", -- 2618
         x"c9",  x"0a",  x"0d",  x"56",  x"65",  x"72",  x"69",  x"66", -- 2620
         x"79",  x"20",  x"28",  x"28",  x"59",  x"29",  x"2f",  x"4e", -- 2628
         x"29",  x"3f",  x"3a",  x"00",  x"0a",  x"52",  x"65",  x"77", -- 2630
         x"69",  x"6e",  x"64",  x"20",  x"3c",  x"3d",  x"3d",  x"0a", -- 2638
         x"0d",  x"00",  x"52",  x"e6",  x"72",  x"e6",  x"34",  x"e7", -- 2640
         x"85",  x"e6",  x"82",  x"dc",  x"6e",  x"e6",  x"82",  x"dc", -- 2648
         x"82",  x"dc",  x"cb",  x"7b",  x"28",  x"11",  x"0e",  x"0b", -- 2650
         x"cd",  x"05",  x"00",  x"b7",  x"28",  x"0e",  x"cb",  x"bb", -- 2658
         x"18",  x"0a",  x"0e",  x"09",  x"cd",  x"05",  x"00",  x"0e", -- 2660
         x"01",  x"cd",  x"05",  x"00",  x"57",  x"c9",  x"0e",  x"05", -- 2668
         x"18",  x"02",  x"0e",  x"02",  x"d5",  x"5a",  x"cd",  x"05", -- 2670
         x"00",  x"d1",  x"cb",  x"bb",  x"c9",  x"16",  x"0a",  x"18", -- 2678
         x"f1",  x"16",  x"0d",  x"18",  x"ed",  x"d5",  x"cb",  x"5b", -- 2680
         x"28",  x"22",  x"d5",  x"0e",  x"0f",  x"cd",  x"05",  x"00", -- 2688
         x"16",  x"20",  x"cd",  x"72",  x"e6",  x"01",  x"0b",  x"00", -- 2690
         x"2a",  x"77",  x"00",  x"23",  x"23",  x"7e",  x"32",  x"75", -- 2698
         x"00",  x"11",  x"80",  x"00",  x"ed",  x"b0",  x"d1",  x"21", -- 26A0
         x"6e",  x"00",  x"36",  x"0b",  x"21",  x"80",  x"00",  x"3a", -- 26A8
         x"6e",  x"00",  x"4f",  x"06",  x"00",  x"09",  x"72",  x"3c", -- 26B0
         x"32",  x"6e",  x"00",  x"cb",  x"73",  x"20",  x"08",  x"3a", -- 26B8
         x"6e",  x"00",  x"fe",  x"80",  x"c2",  x"7d",  x"e7",  x"3a", -- 26C0
         x"75",  x"00",  x"fe",  x"d5",  x"20",  x"1a",  x"21",  x"80", -- 26C8
         x"00",  x"3a",  x"6e",  x"00",  x"47",  x"56",  x"cd",  x"72", -- 26D0
         x"e6",  x"23",  x"10",  x"f9",  x"21",  x"00",  x"00",  x"06", -- 26D8
         x"00",  x"0e",  x"01",  x"a7",  x"ed",  x"42",  x"20",  x"f7", -- 26E0
         x"21",  x"80",  x"00",  x"22",  x"1b",  x"00",  x"0e",  x"15", -- 26E8
         x"cd",  x"05",  x"00",  x"af",  x"32",  x"6e",  x"00",  x"16", -- 26F0
         x"20",  x"cd",  x"72",  x"e6",  x"cb",  x"73",  x"28",  x"74", -- 26F8
         x"af",  x"32",  x"5a",  x"00",  x"11",  x"21",  x"e6",  x"cd", -- 2700
         x"62",  x"e6",  x"cd",  x"72",  x"e6",  x"cd",  x"7d",  x"e6", -- 2708
         x"cd",  x"81",  x"e6",  x"fe",  x"4e",  x"28",  x"66",  x"11", -- 2710
         x"34",  x"e6",  x"cd",  x"62",  x"e6",  x"cd",  x"7d",  x"e6", -- 2718
         x"cd",  x"81",  x"e6",  x"3a",  x"6b",  x"00",  x"47",  x"af", -- 2720
         x"32",  x"6c",  x"00",  x"c5",  x"cd",  x"83",  x"e7",  x"c1", -- 2728
         x"10",  x"f9",  x"18",  x"49",  x"d5",  x"cb",  x"73",  x"20", -- 2730
         x"44",  x"cb",  x"5b",  x"28",  x"1b",  x"cd",  x"7d",  x"e6", -- 2738
         x"3e",  x"01",  x"32",  x"6c",  x"00",  x"cd",  x"83",  x"e7", -- 2740
         x"cd",  x"9d",  x"e7",  x"d1",  x"21",  x"8b",  x"00",  x"56", -- 2748
         x"d5",  x"21",  x"6e",  x"00",  x"36",  x"0c",  x"18",  x"1c", -- 2750
         x"21",  x"80",  x"00",  x"3a",  x"6e",  x"00",  x"4f",  x"06", -- 2758
         x"00",  x"09",  x"d1",  x"56",  x"d5",  x"3c",  x"32",  x"6e", -- 2760
         x"00",  x"fe",  x"80",  x"20",  x"10",  x"cd",  x"83",  x"e7", -- 2768
         x"af",  x"32",  x"6e",  x"00",  x"0e",  x"0b",  x"cd",  x"05", -- 2770
         x"00",  x"fe",  x"03",  x"28",  x"1d",  x"d1",  x"cb",  x"bb", -- 2778
         x"cb",  x"9b",  x"c9",  x"21",  x"80",  x"00",  x"22",  x"1b", -- 2780
         x"00",  x"0e",  x"14",  x"cd",  x"05",  x"00",  x"d0",  x"cd", -- 2788
         x"67",  x"e6",  x"fe",  x"0d",  x"28",  x"ed",  x"fe",  x"03", -- 2790
         x"20",  x"f5",  x"c3",  x"82",  x"dc",  x"21",  x"80",  x"00", -- 2798
         x"06",  x"0b",  x"56",  x"cd",  x"72",  x"e6",  x"23",  x"10", -- 27A0
         x"f9",  x"2a",  x"77",  x"00",  x"0e",  x"0c",  x"09",  x"06", -- 27A8
         x"0b",  x"11",  x"8a",  x"00",  x"1a",  x"be",  x"1b",  x"20", -- 27B0
         x"04",  x"2b",  x"10",  x"f8",  x"c9",  x"d6",  x"04",  x"be", -- 27B8
         x"20",  x"d8",  x"3e",  x"ff",  x"32",  x"5e",  x"03",  x"18", -- 27C0
         x"f0",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 27C8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 27D0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 27D8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ed",  x"53", -- 27E0
         x"3d",  x"00",  x"ed",  x"43",  x"3b",  x"00",  x"51",  x"14", -- 27E8
         x"1c",  x"0e",  x"12",  x"cd",  x"05",  x"00",  x"c9",  x"cd", -- 27F0
         x"21",  x"d4",  x"f5",  x"cd",  x"d6",  x"c8",  x"f1",  x"c9", -- 27F8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2800
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2808
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2810
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2818
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2820
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2828
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2830
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2838
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2840
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2848
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2850
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2858
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2860
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2868
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2870
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2878
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2880
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2888
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2890
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2898
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 28A0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 28A8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 28B0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 28B8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 28C0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 28C8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 28D0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 28D8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 28E0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 28E8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 28F0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 28F8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2900
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2908
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2910
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2918
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2920
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2928
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2930
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2938
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2940
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2948
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2950
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2958
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2960
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2968
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2970
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2978
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2980
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2988
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2990
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2998
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 29A0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 29A8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 29B0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 29B8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 29C0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 29C8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 29D0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 29D8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 29E0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 29E8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 29F0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 29F8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2A00
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2A08
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2A10
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2A18
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2A20
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2A28
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2A30
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2A38
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2A40
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2A48
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2A50
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2A58
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2A60
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2A68
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2A70
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2A78
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2A80
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2A88
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2A90
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2A98
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2AA0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2AA8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2AB0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2AB8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2AC0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2AC8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2AD0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2AD8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2AE0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2AE8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2AF0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2AF8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2B00
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2B08
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2B10
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2B18
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2B20
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2B28
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2B30
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2B38
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2B40
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2B48
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2B50
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2B58
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2B60
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2B68
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2B70
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2B78
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2B80
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2B88
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2B90
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2B98
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2BA0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2BA8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2BB0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2BB8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2BC0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2BC8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2BD0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2BD8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2BE0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2BE8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2BF0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2BF8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2C00
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2C08
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2C10
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2C18
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2C20
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2C28
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2C30
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2C38
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2C40
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2C48
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2C50
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2C58
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2C60
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2C68
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2C70
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2C78
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2C80
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2C88
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2C90
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2C98
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2CA0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2CA8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2CB0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2CB8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2CC0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2CC8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2CD0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2CD8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2CE0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2CE8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2CF0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2CF8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2D00
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2D08
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2D10
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2D18
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2D20
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2D28
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2D30
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2D38
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2D40
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2D48
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2D50
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2D58
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2D60
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2D68
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2D70
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2D78
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2D80
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2D88
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2D90
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2D98
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2DA0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2DA8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2DB0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2DB8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2DC0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2DC8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2DD0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2DD8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2DE0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2DE8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2DF0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2DF8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2E00
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2E08
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2E10
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2E18
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2E20
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2E28
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2E30
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2E38
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2E40
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2E48
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2E50
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2E58
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2E60
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2E68
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2E70
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2E78
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2E80
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2E88
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2E90
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2E98
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2EA0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2EA8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2EB0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2EB8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2EC0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2EC8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2ED0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2ED8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2EE0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2EE8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2EF0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2EF8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2F00
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2F08
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2F10
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2F18
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2F20
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2F28
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2F30
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2F38
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2F40
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2F48
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2F50
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2F58
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2F60
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2F68
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2F70
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2F78
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2F80
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2F88
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2F90
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2F98
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2FA0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2FA8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2FB0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2FB8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2FC0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2FC8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2FD0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2FD8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2FE0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2FE8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2FF0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 2FF8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3000
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3008
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3010
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3018
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3020
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3028
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3030
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3038
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3040
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3048
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3050
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3058
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3060
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3068
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3070
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3078
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3080
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3088
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3090
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3098
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 30A0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 30A8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 30B0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 30B8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 30C0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 30C8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 30D0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 30D8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 30E0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 30E8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 30F0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 30F8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3100
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3108
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3110
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3118
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3120
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3128
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3130
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3138
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3140
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3148
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3150
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3158
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3160
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3168
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3170
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3178
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3180
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3188
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3190
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3198
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 31A0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 31A8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 31B0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 31B8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 31C0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 31C8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 31D0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 31D8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 31E0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 31E8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 31F0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 31F8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3200
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3208
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3210
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3218
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3220
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3228
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3230
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3238
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3240
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3248
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3250
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3258
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3260
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3268
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3270
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3278
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3280
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3288
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3290
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3298
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 32A0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 32A8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 32B0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 32B8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 32C0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 32C8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 32D0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 32D8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 32E0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 32E8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 32F0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 32F8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3300
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3308
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3310
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3318
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3320
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3328
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3330
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3338
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3340
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3348
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3350
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3358
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3360
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3368
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3370
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3378
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3380
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3388
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3390
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3398
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 33A0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 33A8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 33B0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 33B8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 33C0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 33C8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 33D0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 33D8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 33E0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 33E8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 33F0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 33F8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3400
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3408
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3410
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3418
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3420
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3428
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3430
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3438
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3440
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3448
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3450
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3458
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3460
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3468
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3470
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3478
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3480
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3488
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3490
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3498
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 34A0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 34A8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 34B0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 34B8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 34C0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 34C8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 34D0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 34D8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 34E0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 34E8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 34F0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 34F8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3500
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3508
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3510
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3518
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3520
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3528
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3530
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3538
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3540
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3548
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3550
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3558
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3560
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3568
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3570
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3578
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3580
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3588
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3590
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3598
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 35A0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 35A8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 35B0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 35B8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 35C0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 35C8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 35D0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 35D8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 35E0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 35E8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 35F0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 35F8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3600
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3608
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3610
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3618
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3620
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3628
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3630
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3638
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3640
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3648
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3650
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3658
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3660
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3668
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3670
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3678
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3680
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3688
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3690
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3698
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 36A0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 36A8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 36B0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 36B8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 36C0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 36C8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 36D0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 36D8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 36E0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 36E8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 36F0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 36F8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3700
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3708
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3710
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3718
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3720
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3728
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3730
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3738
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3740
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3748
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3750
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3758
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3760
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3768
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3770
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3778
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3780
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3788
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3790
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3798
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 37A0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 37A8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 37B0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 37B8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 37C0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 37C8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 37D0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 37D8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 37E0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 37E8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 37F0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 37F8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3800
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3808
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3810
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3818
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3820
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3828
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3830
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3838
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3840
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3848
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3850
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3858
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3860
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3868
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3870
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3878
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3880
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3888
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3890
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3898
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 38A0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 38A8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 38B0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 38B8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 38C0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 38C8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 38D0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 38D8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 38E0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 38E8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 38F0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 38F8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3900
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3908
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3910
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3918
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3920
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3928
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3930
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3938
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3940
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3948
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3950
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3958
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3960
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3968
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3970
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3978
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3980
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3988
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3990
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3998
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 39A0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 39A8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 39B0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 39B8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 39C0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 39C8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 39D0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 39D8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 39E0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 39E8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 39F0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 39F8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A00
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A08
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A10
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A18
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A20
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A28
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A30
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A38
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A40
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A48
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A50
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A58
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A60
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A68
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A70
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A78
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A80
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A88
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A90
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3A98
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3AA0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3AA8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3AB0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3AB8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3AC0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3AC8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3AD0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3AD8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3AE0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3AE8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3AF0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3AF8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B00
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B08
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B10
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B18
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B20
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B28
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B30
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B38
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B40
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B48
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B50
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B58
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B60
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B68
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B70
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B78
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B80
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B88
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B90
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3B98
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3BA0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3BA8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3BB0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3BB8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3BC0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3BC8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3BD0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3BD8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3BE0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3BE8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3BF0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3BF8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C00
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C08
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C10
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C18
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C20
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C28
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C30
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C38
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C40
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C48
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C50
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C58
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C60
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C68
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C70
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C78
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C80
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C88
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C90
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3C98
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3CA0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3CA8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3CB0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3CB8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3CC0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3CC8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3CD0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3CD8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3CE0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3CE8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3CF0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3CF8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D00
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D08
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D10
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D18
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D20
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D28
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D30
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D38
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D40
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D48
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D50
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D58
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D60
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D68
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D70
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D78
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D80
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D88
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D90
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3D98
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3DA0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3DA8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3DB0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3DB8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3DC0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3DC8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3DD0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3DD8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3DE0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3DE8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3DF0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3DF8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E00
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E08
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E10
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E18
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E20
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E28
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E30
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E38
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E40
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E48
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E50
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E58
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E60
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E68
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E70
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E78
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E80
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E88
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E90
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3E98
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3EA0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3EA8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3EB0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3EB8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3EC0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3EC8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3ED0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3ED8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3EE0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3EE8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3EF0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3EF8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F00
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F08
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F10
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F18
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F20
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F28
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F30
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F38
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F40
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F48
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F50
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F58
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F60
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F68
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F70
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F78
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F80
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F88
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F90
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3F98
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3FA0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3FA8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3FB0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3FB8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3FC0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3FC8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3FD0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3FD8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3FE0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3FE8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3FF0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00"  -- 3FF8
        );
    
begin
    process begin
        wait until rising_edge(clk);
        data <= romData(to_integer(unsigned(addr)));
    end process;
end;
