library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity bwidow_vec_rom2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of bwidow_vec_rom2 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"32",X"00",X"00",X"00",X"25",X"45",X"00",X"00",X"28",X"20",X"25",X"5B",X"20",X"5B",X"16",X"56",
		X"2A",X"40",X"20",X"5B",X"3B",X"5B",X"1B",X"45",X"36",X"40",X"28",X"00",X"00",X"20",X"CE",X"1F",
		X"28",X"00",X"0A",X"40",X"5A",X"00",X"00",X"00",X"2A",X"40",X"CE",X"1F",X"00",X"20",X"2A",X"4A",
		X"2A",X"40",X"11",X"51",X"2F",X"51",X"00",X"00",X"D8",X"1F",X"20",X"4A",X"EC",X"1F",X"28",X"00",
		X"0A",X"40",X"00",X"C0",X"5A",X"00",X"00",X"00",X"2A",X"40",X"25",X"56",X"05",X"4A",X"2A",X"40",
		X"25",X"56",X"05",X"4A",X"2A",X"40",X"A6",X"1F",X"EC",X"3F",X"32",X"00",X"E2",X"1F",X"CE",X"1F",
		X"EC",X"3F",X"00",X"00",X"46",X"00",X"0A",X"40",X"3C",X"00",X"00",X"00",X"2A",X"40",X"C4",X"1F",
		X"00",X"20",X"46",X"00",X"00",X"00",X"20",X"4A",X"36",X"40",X"A6",X"1F",X"14",X"00",X"0A",X"40",
		X"5A",X"00",X"28",X"00",X"2A",X"40",X"A6",X"1F",X"00",X"20",X"32",X"00",X"EC",X"1F",X"3B",X"45",
		X"36",X"40",X"3B",X"5B",X"D8",X"1F",X"28",X"00",X"3B",X"5B",X"28",X"00",X"EC",X"1F",X"20",X"51",
		X"25",X"40",X"F6",X"1F",X"28",X"00",X"0A",X"40",X"32",X"00",X"00",X"00",X"25",X"45",X"00",X"00",
		X"28",X"20",X"25",X"5B",X"D8",X"1F",X"00",X"20",X"3B",X"5B",X"1B",X"45",X"36",X"40",X"28",X"00",
		X"00",X"20",X"CE",X"1F",X"28",X"00",X"0A",X"40",X"3C",X"00",X"00",X"00",X"2A",X"40",X"25",X"56",
		X"05",X"4A",X"2A",X"40",X"25",X"56",X"05",X"4A",X"2A",X"40",X"C4",X"1F",X"EC",X"3F",X"11",X"4F",
		X"3B",X"51",X"00",X"00",X"3C",X"00",X"0A",X"40",X"00",X"C0",X"00",X"49",X"3E",X"5B",X"3B",X"43",
		X"23",X"5B",X"3B",X"5E",X"25",X"5E",X"3D",X"5B",X"25",X"43",X"22",X"5B",X"22",X"45",X"25",X"5D",
		X"3D",X"45",X"25",X"42",X"3B",X"42",X"23",X"45",X"3B",X"5D",X"3E",X"45",X"00",X"57",X"00",X"C0",
		X"02",X"49",X"3D",X"5B",X"3C",X"45",X"22",X"5A",X"3A",X"5F",X"25",X"5F",X"3B",X"5A",X"26",X"42",
		X"21",X"5A",X"21",X"45",X"26",X"5B",X"3E",X"46",X"26",X"41",X"3B",X"43",X"25",X"44",X"3A",X"5E",
		X"3F",X"46",X"1E",X"57",X"00",X"C0",X"04",X"48",X"3C",X"5C",X"3D",X"46",X"21",X"5A",X"3A",X"40",
		X"24",X"5C",X"3A",X"5D",X"26",X"41",X"20",X"5A",X"24",X"44",X"23",X"5A",X"3F",X"46",X"26",X"40",
		X"3C",X"44",X"26",X"43",X"3A",X"5F",X"20",X"46",X"1C",X"58",X"00",X"C0",X"1E",X"43",X"3E",X"5D",
		X"21",X"5D",X"23",X"54",X"23",X"4C",X"21",X"43",X"3E",X"43",X"3E",X"48",X"3E",X"58",X"02",X"5D",
		X"00",X"C0",X"1F",X"44",X"3D",X"5E",X"20",X"5C",X"3E",X"54",X"28",X"4A",X"22",X"42",X"3F",X"44",
		X"21",X"48",X"3B",X"5A",X"01",X"5C",X"00",X"C0",X"1F",X"44",X"3E",X"5F",X"3F",X"5D",X"39",X"55",
		X"2B",X"47",X"23",X"41",X"21",X"44",X"24",X"47",X"37",X"5C",X"01",X"5C",X"00",X"C0",X"02",X"43",
		X"3C",X"41",X"3E",X"5E",X"36",X"58",X"2C",X"42",X"24",X"40",X"22",X"45",X"26",X"43",X"38",X"5F",
		X"1E",X"5D",X"00",X"C0",X"03",X"42",X"3D",X"42",X"3D",X"5F",X"34",X"5D",X"2C",X"5D",X"23",X"5F",
		X"23",X"42",X"28",X"42",X"38",X"42",X"1D",X"5E",X"00",X"C0",X"04",X"41",X"3E",X"43",X"3C",X"40",
		X"34",X"42",X"2A",X"58",X"22",X"5E",X"24",X"41",X"28",X"5F",X"3A",X"45",X"1C",X"5F",X"00",X"C0",
		X"04",X"41",X"3F",X"42",X"3D",X"41",X"35",X"47",X"27",X"55",X"21",X"5D",X"22",X"5F",X"29",X"5C",
		X"3C",X"49",X"1C",X"5F",X"00",X"C0",X"03",X"5E",X"21",X"44",X"3E",X"42",X"38",X"4A",X"22",X"54",
		X"20",X"5C",X"23",X"5E",X"25",X"5A",X"3F",X"48",X"1D",X"42",X"00",X"C0",X"02",X"5D",X"22",X"43",
		X"3F",X"43",X"3D",X"4C",X"3D",X"54",X"3F",X"5D",X"22",X"5D",X"22",X"58",X"22",X"48",X"1E",X"43",
		X"00",X"C0",X"1F",X"5C",X"25",X"42",X"20",X"44",X"22",X"4C",X"38",X"56",X"3E",X"5E",X"21",X"5C",
		X"3F",X"58",X"23",X"46",X"01",X"44",X"00",X"C0",X"1F",X"5C",X"24",X"41",X"21",X"43",X"27",X"4B",
		X"35",X"59",X"3D",X"5F",X"3F",X"5E",X"3C",X"57",X"27",X"44",X"01",X"44",X"00",X"C0",X"1E",X"5D",
		X"24",X"5F",X"22",X"42",X"2A",X"48",X"34",X"5E",X"3C",X"40",X"3E",X"5D",X"3A",X"5B",X"28",X"41",
		X"02",X"43",X"00",X"C0",X"1D",X"5E",X"23",X"5E",X"23",X"41",X"2C",X"43",X"34",X"43",X"3D",X"41",
		X"3D",X"5E",X"38",X"5E",X"28",X"5E",X"03",X"42",X"00",X"C0",X"1C",X"41",X"22",X"5B",X"24",X"40",
		X"2C",X"5E",X"36",X"48",X"3E",X"42",X"3C",X"5F",X"38",X"41",X"26",X"5D",X"04",X"5F",X"00",X"C0",
		X"1C",X"41",X"21",X"5C",X"23",X"5F",X"2B",X"59",X"39",X"4B",X"3F",X"43",X"3C",X"41",X"39",X"44",
		X"24",X"59",X"04",X"5F",X"00",X"C0",X"1D",X"42",X"3F",X"5C",X"22",X"5E",X"28",X"56",X"3E",X"4C",
		X"20",X"44",X"3B",X"42",X"3D",X"46",X"21",X"58",X"03",X"5E",X"00",X"C0",X"1E",X"43",X"3E",X"5D",
		X"21",X"5D",X"22",X"5F",X"3B",X"5C",X"20",X"5B",X"24",X"5C",X"24",X"40",X"24",X"44",X"20",X"45",
		X"3B",X"44",X"22",X"41",X"21",X"43",X"3E",X"43",X"3C",X"40",X"02",X"5D",X"00",X"C0",X"1F",X"44",
		X"3D",X"5E",X"20",X"5C",X"22",X"5F",X"39",X"5E",X"3E",X"5B",X"23",X"5B",X"23",X"5F",X"24",X"42",
		X"23",X"44",X"3D",X"46",X"23",X"40",X"22",X"42",X"3F",X"44",X"3C",X"42",X"01",X"5C",X"00",X"C0",
		X"1F",X"44",X"3E",X"5F",X"3F",X"5D",X"20",X"5E",X"3A",X"41",X"3D",X"5C",X"20",X"5A",X"22",X"5E",
		X"26",X"40",X"24",X"43",X"3F",X"46",X"22",X"40",X"23",X"41",X"21",X"44",X"3B",X"43",X"01",X"5C",
		X"00",X"C0",X"02",X"43",X"3C",X"41",X"3E",X"5E",X"20",X"5F",X"3A",X"41",X"3C",X"5F",X"3E",X"5A",
		X"21",X"5D",X"25",X"5D",X"25",X"42",X"22",X"47",X"21",X"5E",X"24",X"40",X"22",X"45",X"3E",X"42",
		X"1E",X"5D",X"00",X"C0",X"03",X"42",X"3D",X"42",X"3D",X"5F",X"3F",X"5E",X"3C",X"45",X"3B",X"40",
		X"3C",X"5C",X"20",X"5C",X"24",X"5C",X"25",X"40",X"24",X"45",X"21",X"5E",X"23",X"5F",X"23",X"42",
		X"20",X"44",X"1D",X"5E",X"00",X"C0",X"04",X"41",X"3E",X"43",X"3C",X"40",X"3F",X"5E",X"3E",X"47",
		X"3B",X"42",X"3B",X"5D",X"3F",X"5D",X"22",X"5C",X"24",X"5D",X"26",X"43",X"20",X"5D",X"22",X"5E",
		X"24",X"41",X"22",X"44",X"1C",X"5F",X"00",X"C0",X"04",X"41",X"3F",X"42",X"3D",X"41",X"3E",X"40",
		X"21",X"46",X"3C",X"43",X"3A",X"40",X"3E",X"5E",X"20",X"5A",X"23",X"5C",X"26",X"41",X"20",X"5E",
		X"21",X"5D",X"22",X"5F",X"25",X"45",X"1C",X"5F",X"00",X"C0",X"03",X"5E",X"21",X"44",X"3E",X"42",
		X"3D",X"40",X"23",X"46",X"3D",X"44",X"3C",X"42",X"3D",X"5F",X"3D",X"5B",X"22",X"5B",X"27",X"5E",
		X"3E",X"5F",X"20",X"5C",X"23",X"5E",X"24",X"42",X"1D",X"42",X"00",X"C0",X"02",X"5D",X"22",X"43",
		X"3F",X"43",X"3C",X"41",X"27",X"44",X"20",X"45",X"3C",X"44",X"3C",X"40",X"3C",X"5C",X"20",X"5B",
		X"25",X"5C",X"3E",X"5F",X"3F",X"5D",X"22",X"5D",X"24",X"40",X"1E",X"43",X"00",X"C0",X"1F",X"5C",
		X"25",X"42",X"20",X"44",X"3E",X"41",X"27",X"42",X"22",X"45",X"3D",X"45",X"3D",X"41",X"3A",X"5E",
		X"3F",X"5C",X"21",X"5A",X"3F",X"40",X"3E",X"5E",X"21",X"5C",X"22",X"5E",X"01",X"44",X"00",X"C0",
		X"1F",X"5C",X"24",X"41",X"21",X"43",X"20",X"42",X"26",X"5F",X"23",X"44",X"20",X"46",X"3E",X"42",
		X"3A",X"40",X"3C",X"5D",X"21",X"5A",X"3E",X"40",X"3D",X"5F",X"3F",X"5E",X"23",X"5B",X"01",X"44",
		X"00",X"C0",X"1E",X"5D",X"24",X"5F",X"22",X"42",X"20",X"43",X"26",X"5D",X"24",X"43",X"22",X"44",
		X"3F",X"43",X"3B",X"43",X"3B",X"5E",X"3E",X"59",X"3F",X"42",X"3C",X"40",X"3E",X"5D",X"22",X"5C",
		X"02",X"43",X"00",X"C0",X"1D",X"5E",X"23",X"5E",X"23",X"41",X"21",X"42",X"24",X"5B",X"25",X"40",
		X"24",X"44",X"20",X"44",X"3C",X"44",X"3B",X"40",X"3C",X"5B",X"3F",X"42",X"3D",X"41",X"3D",X"5E",
		X"20",X"5C",X"03",X"42",X"00",X"C0",X"1C",X"41",X"22",X"5B",X"24",X"40",X"21",X"42",X"22",X"59",
		X"25",X"5E",X"25",X"43",X"21",X"43",X"3E",X"46",X"3C",X"41",X"3A",X"5F",X"20",X"41",X"3E",X"42",
		X"3C",X"5F",X"3E",X"5E",X"04",X"5F",X"00",X"C0",X"1C",X"41",X"21",X"5C",X"23",X"5F",X"22",X"40",
		X"3F",X"5A",X"24",X"5D",X"26",X"40",X"22",X"42",X"20",X"46",X"3D",X"44",X"3A",X"5F",X"20",X"42",
		X"3F",X"43",X"3C",X"41",X"3D",X"5D",X"04",X"5F",X"00",X"C0",X"1D",X"42",X"3F",X"5C",X"22",X"5E",
		X"21",X"40",X"3F",X"5A",X"21",X"5C",X"26",X"5E",X"23",X"41",X"23",X"45",X"3E",X"45",X"39",X"42",
		X"22",X"41",X"20",X"44",X"3B",X"42",X"3E",X"5E",X"03",X"5E",X"00",X"C0",X"1E",X"43",X"3E",X"5D",
		X"21",X"5D",X"3F",X"5D",X"20",X"5C",X"24",X"5D",X"24",X"43",X"20",X"44",X"3F",X"43",X"21",X"43",
		X"3E",X"43",X"21",X"43",X"20",X"43",X"3D",X"42",X"3D",X"5E",X"20",X"5D",X"21",X"5D",X"1E",X"57",
		X"28",X"40",X"00",X"5E",X"38",X"40",X"00",X"5E",X"28",X"40",X"1C",X"4A",X"00",X"C0",X"1F",X"44",
		X"3D",X"5E",X"20",X"5C",X"3E",X"5E",X"3E",X"5C",X"23",X"5C",X"25",X"41",X"21",X"44",X"21",X"43",
		X"22",X"42",X"3F",X"44",X"22",X"42",X"21",X"43",X"3E",X"43",X"3B",X"5F",X"21",X"5E",X"3F",X"5D",
		X"1B",X"58",X"27",X"5D",X"1E",X"5E",X"3A",X"43",X"1F",X"5E",X"28",X"5D",X"00",X"4B",X"00",X"C0",
		X"1F",X"44",X"3E",X"5F",X"3F",X"5D",X"3D",X"5F",X"3D",X"5D",X"21",X"5B",X"25",X"5F",X"23",X"43",
		X"21",X"43",X"23",X"41",X"21",X"44",X"22",X"41",X"22",X"42",X"20",X"44",X"3C",X"40",X"3E",X"5E",
		X"3D",X"5E",X"1A",X"5B",X"26",X"5A",X"1E",X"5F",X"3B",X"45",X"1E",X"5F",X"26",X"5A",X"04",X"4A",
		X"00",X"C0",X"E7",X"00",X"02",X"43",X"3C",X"41",X"3E",X"5E",X"3D",X"5F",X"3C",X"5F",X"3F",X"5B",
		X"24",X"5D",X"24",X"42",X"22",X"42",X"24",X"40",X"22",X"45",X"23",X"5F",X"22",X"41",X"21",X"43",
		X"3D",X"42",X"3D",X"5F",X"3E",X"5E",X"17",X"5E",X"23",X"59",X"1E",X"5F",X"3D",X"48",X"1E",X"5F",
		X"23",X"58",X"08",X"48",X"00",X"C0",X"03",X"42",X"3D",X"42",X"3D",X"5F",X"3D",X"41",X"3C",X"40",
		X"3D",X"5C",X"23",X"5C",X"24",X"40",X"23",X"41",X"23",X"5F",X"23",X"42",X"23",X"5F",X"23",X"40",
		X"22",X"43",X"3E",X"43",X"3D",X"40",X"3D",X"5F",X"17",X"42",X"20",X"58",X"1E",X"40",X"20",X"48",
		X"1E",X"40",X"20",X"58",X"0A",X"44",X"00",X"C0",X"04",X"41",X"3E",X"43",X"3C",X"40",X"3E",X"42",
		X"3C",X"42",X"3C",X"5D",X"21",X"5B",X"24",X"5F",X"23",X"5F",X"22",X"5E",X"24",X"41",X"22",X"5E",
		X"23",X"5F",X"23",X"42",X"3F",X"45",X"3E",X"5F",X"3D",X"41",X"18",X"45",X"3D",X"59",X"1E",X"42",
		X"23",X"46",X"1E",X"41",X"3D",X"58",X"0B",X"40",X"00",X"C0",X"04",X"41",X"3F",X"42",X"3D",X"41",
		X"3F",X"43",X"3D",X"43",X"3B",X"5F",X"3F",X"5B",X"23",X"5D",X"23",X"5F",X"21",X"5D",X"22",X"5F",
		X"23",X"5E",X"22",X"5E",X"24",X"40",X"20",X"44",X"3E",X"42",X"3E",X"43",X"1B",X"46",X"3A",X"5A",
		X"1F",X"42",X"25",X"45",X"1F",X"42",X"3A",X"5A",X"0A",X"5C",X"00",X"C0",X"03",X"5E",X"21",X"44",
		X"3E",X"42",X"3F",X"43",X"3F",X"44",X"3B",X"41",X"3D",X"5C",X"22",X"5C",X"22",X"5E",X"20",X"5C",
		X"23",X"5E",X"21",X"5D",X"3F",X"5E",X"25",X"5F",X"22",X"43",X"3F",X"43",X"3E",X"42",X"1E",X"49",
		X"39",X"5D",X"1F",X"42",X"26",X"43",X"01",X"42",X"38",X"5D",X"08",X"58",X"00",X"C0",X"02",X"5D",
		X"22",X"43",X"3F",X"43",X"21",X"43",X"20",X"44",X"3C",X"43",X"3C",X"5D",X"20",X"5C",X"21",X"5D",
		X"3F",X"5D",X"22",X"5D",X"3F",X"5D",X"20",X"5D",X"23",X"5E",X"23",X"42",X"20",X"43",X"3F",X"43",
		X"02",X"49",X"38",X"40",X"00",X"42",X"28",X"40",X"00",X"42",X"38",X"40",X"04",X"56",X"00",X"C0",
		X"1F",X"5C",X"25",X"42",X"20",X"44",X"22",X"42",X"22",X"44",X"3D",X"44",X"3B",X"5F",X"3F",X"5C",
		X"3F",X"5D",X"3E",X"5E",X"21",X"5C",X"3E",X"5E",X"3F",X"5D",X"22",X"5D",X"23",X"41",X"21",X"42",
		X"3F",X"43",X"07",X"48",X"39",X"43",X"00",X"42",X"28",X"5D",X"01",X"42",X"38",X"43",X"00",X"55",
		X"00",X"C0",X"1F",X"5C",X"24",X"41",X"21",X"43",X"23",X"41",X"23",X"43",X"3F",X"45",X"3B",X"41",
		X"3D",X"5D",X"3F",X"5D",X"3D",X"5F",X"3F",X"5E",X"3E",X"5D",X"3E",X"5E",X"20",X"5C",X"24",X"40",
		X"22",X"42",X"21",X"42",X"08",X"45",X"3A",X"46",X"02",X"41",X"25",X"5B",X"02",X"41",X"3A",X"46",
		X"1C",X"56",X"00",X"C0",X"1E",X"5D",X"24",X"5F",X"22",X"42",X"23",X"41",X"24",X"41",X"21",X"45",
		X"3C",X"43",X"3C",X"5E",X"3E",X"5E",X"3C",X"40",X"3E",X"5D",X"3D",X"5F",X"3E",X"41",X"3F",X"5B",
		X"23",X"5E",X"23",X"41",X"22",X"42",X"09",X"42",X"3D",X"47",X"02",X"41",X"23",X"5A",X"02",X"5F",
		X"3D",X"48",X"18",X"58",X"00",X"C0",X"1D",X"5E",X"23",X"5E",X"23",X"41",X"23",X"5F",X"24",X"40",
		X"23",X"44",X"3D",X"44",X"3C",X"40",X"3D",X"5F",X"3D",X"41",X"3D",X"5E",X"3D",X"41",X"3D",X"40",
		X"3E",X"5D",X"22",X"5D",X"23",X"40",X"23",X"41",X"09",X"5E",X"20",X"48",X"02",X"40",X"20",X"58",
		X"02",X"40",X"20",X"48",X"16",X"5C",X"00",X"C0",X"1C",X"41",X"22",X"5B",X"24",X"40",X"22",X"5E",
		X"24",X"5E",X"24",X"43",X"3F",X"45",X"3C",X"41",X"3D",X"41",X"3E",X"42",X"3C",X"5F",X"3E",X"42",
		X"3D",X"41",X"3D",X"5E",X"21",X"5D",X"22",X"5F",X"23",X"41",X"08",X"59",X"23",X"47",X"02",X"40",
		X"3D",X"58",X"02",X"5F",X"23",X"48",X"15",X"40",X"00",X"C0",X"1C",X"41",X"21",X"5C",X"23",X"5F",
		X"21",X"5D",X"23",X"5D",X"25",X"41",X"21",X"45",X"3D",X"43",X"3D",X"41",X"3F",X"43",X"3C",X"41",
		X"3F",X"42",X"3E",X"42",X"3C",X"40",X"20",X"5C",X"22",X"5E",X"22",X"5F",X"05",X"58",X"26",X"46",
		X"01",X"5E",X"3B",X"5B",X"01",X"5E",X"26",X"46",X"16",X"44",X"00",X"C0",X"1D",X"42",X"3F",X"5C",
		X"22",X"5E",X"21",X"5D",X"21",X"5C",X"25",X"5F",X"23",X"44",X"3E",X"44",X"3E",X"42",X"20",X"44",
		X"3B",X"42",X"21",X"43",X"3F",X"42",X"3D",X"41",X"3E",X"5D",X"21",X"5D",X"22",X"5E",X"02",X"57",
		X"27",X"43",X"01",X"5E",X"38",X"5D",X"01",X"5E",X"28",X"43",X"18",X"48",X"00",X"C0",X"24",X"40",
		X"23",X"43",X"20",X"44",X"3D",X"43",X"38",X"40",X"3D",X"5D",X"07",X"59",X"3C",X"40",X"3D",X"5D",
		X"20",X"5C",X"23",X"5D",X"28",X"40",X"23",X"43",X"1B",X"5A",X"20",X"4D",X"20",X"4D",X"1C",X"40",
		X"20",X"53",X"20",X"53",X"02",X"4D",X"00",X"C0",X"24",X"5E",X"24",X"42",X"21",X"44",X"3F",X"44",
		X"38",X"43",X"3C",X"5E",X"04",X"57",X"3C",X"42",X"3C",X"5E",X"3F",X"5C",X"21",X"5C",X"28",X"5D",
		X"24",X"42",X"19",X"5C",X"25",X"4E",X"25",X"4A",X"1C",X"42",X"3B",X"54",X"3B",X"54",X"07",X"4B",
		X"00",X"C0",X"23",X"5D",X"24",X"40",X"23",X"43",X"20",X"44",X"3A",X"46",X"3C",X"40",X"00",X"56",
		X"3D",X"43",X"3C",X"40",X"3D",X"5D",X"20",X"5C",X"26",X"5A",X"24",X"40",X"18",X"5F",X"29",X"4A",
		X"2A",X"49",X"1D",X"43",X"37",X"56",X"36",X"57",X"0B",X"48",X"00",X"C0",X"22",X"5C",X"23",X"5F",
		X"24",X"41",X"22",X"44",X"3D",X"48",X"3C",X"41",X"1C",X"57",X"3E",X"44",X"3D",X"41",X"3C",X"5F",
		X"3E",X"5C",X"23",X"58",X"24",X"5F",X"19",X"42",X"2A",X"45",X"2E",X"45",X"1E",X"44",X"34",X"5B",
		X"34",X"5B",X"0D",X"43",X"00",X"C0",X"20",X"5C",X"23",X"5D",X"24",X"40",X"23",X"43",X"20",X"48",
		X"3D",X"43",X"19",X"59",X"20",X"44",X"3D",X"43",X"3C",X"40",X"3D",X"5D",X"20",X"58",X"23",X"5D",
		X"1A",X"45",X"2D",X"40",X"2D",X"40",X"00",X"44",X"33",X"40",X"33",X"40",X"0D",X"5E",X"00",X"C0",
		X"3E",X"5C",X"22",X"5C",X"24",X"5F",X"24",X"41",X"23",X"48",X"3E",X"44",X"17",X"5C",X"22",X"44",
		X"3E",X"44",X"3C",X"41",X"3C",X"5F",X"3D",X"58",X"22",X"5C",X"1C",X"47",X"2C",X"5B",X"2C",X"5B",
		X"02",X"44",X"32",X"45",X"36",X"45",X"0B",X"59",X"00",X"C0",X"3D",X"5D",X"20",X"5C",X"23",X"5D",
		X"24",X"40",X"26",X"46",X"20",X"44",X"16",X"40",X"23",X"43",X"20",X"44",X"3D",X"43",X"3C",X"40",
		X"3A",X"5A",X"20",X"5C",X"1F",X"48",X"2A",X"57",X"29",X"56",X"03",X"43",X"36",X"49",X"37",X"4A",
		X"08",X"55",X"00",X"C0",X"3C",X"5E",X"3F",X"5D",X"21",X"5C",X"24",X"5E",X"28",X"43",X"21",X"44",
		X"17",X"44",X"24",X"42",X"21",X"43",X"3F",X"44",X"3C",X"42",X"38",X"5D",X"3F",X"5C",X"02",X"47",
		X"25",X"56",X"25",X"52",X"04",X"42",X"3B",X"4C",X"3B",X"4C",X"03",X"53",X"00",X"C0",X"3C",X"40",
		X"3D",X"5D",X"20",X"5C",X"23",X"5D",X"28",X"40",X"23",X"43",X"19",X"47",X"24",X"40",X"23",X"43",
		X"20",X"44",X"3D",X"43",X"38",X"40",X"3D",X"5D",X"05",X"46",X"20",X"53",X"20",X"53",X"04",X"40",
		X"20",X"4D",X"20",X"4D",X"1E",X"53",X"00",X"C0",X"3C",X"42",X"3C",X"5E",X"3F",X"5C",X"21",X"5C",
		X"28",X"5D",X"24",X"42",X"1C",X"49",X"24",X"5E",X"24",X"42",X"21",X"44",X"3F",X"44",X"38",X"43",
		X"3C",X"5E",X"07",X"44",X"3B",X"54",X"3B",X"54",X"04",X"5E",X"25",X"4E",X"25",X"4A",X"19",X"55",
		X"00",X"C0",X"3D",X"43",X"3C",X"40",X"3D",X"5D",X"20",X"5C",X"26",X"5A",X"24",X"40",X"00",X"4A",
		X"23",X"5D",X"24",X"40",X"23",X"43",X"20",X"44",X"3A",X"46",X"3C",X"40",X"08",X"41",X"37",X"56",
		X"36",X"57",X"03",X"5D",X"29",X"4A",X"2A",X"49",X"15",X"58",X"00",X"C0",X"3E",X"44",X"3D",X"41",
		X"3C",X"5F",X"3E",X"5C",X"23",X"58",X"24",X"5F",X"04",X"49",X"22",X"5C",X"23",X"5F",X"24",X"41",
		X"22",X"44",X"3D",X"48",X"3C",X"41",X"07",X"5E",X"34",X"5B",X"34",X"5B",X"02",X"5C",X"2A",X"45",
		X"2E",X"45",X"13",X"5D",X"00",X"C0",X"20",X"44",X"3D",X"43",X"3C",X"40",X"3D",X"5D",X"20",X"58",
		X"23",X"5D",X"07",X"47",X"20",X"5C",X"23",X"5D",X"24",X"40",X"23",X"43",X"20",X"48",X"3D",X"43",
		X"06",X"5B",X"33",X"40",X"33",X"40",X"00",X"5C",X"2D",X"40",X"2D",X"40",X"13",X"42",X"00",X"C0",
		X"22",X"44",X"3E",X"44",X"3C",X"41",X"3C",X"5F",X"3D",X"58",X"22",X"5C",X"09",X"44",X"3E",X"5C",
		X"22",X"5C",X"24",X"5F",X"24",X"41",X"23",X"48",X"3E",X"44",X"04",X"59",X"32",X"45",X"36",X"45",
		X"1E",X"5C",X"2C",X"5B",X"2C",X"5B",X"15",X"47",X"00",X"C0",X"23",X"43",X"20",X"44",X"3D",X"43",
		X"3C",X"40",X"3A",X"5A",X"20",X"5C",X"0A",X"40",X"3D",X"5D",X"20",X"5C",X"23",X"5D",X"24",X"40",
		X"26",X"46",X"20",X"44",X"01",X"58",X"36",X"49",X"37",X"4A",X"1D",X"5D",X"2A",X"57",X"29",X"56",
		X"18",X"4B",X"00",X"C0",X"24",X"42",X"21",X"43",X"3F",X"44",X"3C",X"42",X"38",X"5D",X"3F",X"5C",
		X"09",X"5C",X"3C",X"5E",X"3F",X"5D",X"21",X"5C",X"24",X"5E",X"28",X"43",X"21",X"44",X"1E",X"59",
		X"3B",X"4C",X"3B",X"4C",X"1C",X"5E",X"25",X"56",X"25",X"52",X"1D",X"4D",X"00",X"C0",X"1C",X"40",
		X"21",X"5D",X"3F",X"5D",X"22",X"58",X"22",X"48",X"22",X"58",X"22",X"48",X"3F",X"43",X"21",X"43",
		X"3C",X"46",X"3C",X"5A",X"03",X"56",X"21",X"5C",X"21",X"44",X"1F",X"4A",X"00",X"C0",X"1C",X"42",
		X"20",X"5C",X"3E",X"5E",X"3F",X"58",X"25",X"46",X"3E",X"58",X"25",X"47",X"21",X"43",X"22",X"42",
		X"3E",X"48",X"3A",X"5C",X"1F",X"55",X"20",X"5C",X"22",X"43",X"03",X"4A",X"00",X"C0",X"1D",X"43",
		X"3F",X"5D",X"3D",X"5F",X"3C",X"59",X"27",X"44",X"3C",X"59",X"27",X"44",X"21",X"43",X"23",X"41",
		X"21",X"47",X"39",X"5F",X"1B",X"57",X"3E",X"5C",X"24",X"42",X"06",X"48",X"00",X"C0",X"1E",X"44",
		X"3E",X"5E",X"3D",X"5F",X"39",X"5B",X"28",X"42",X"3A",X"5B",X"28",X"41",X"22",X"42",X"24",X"40",
		X"24",X"46",X"38",X"42",X"18",X"59",X"3D",X"5E",X"24",X"40",X"09",X"45",X"00",X"C0",X"00",X"44",
		X"3D",X"5F",X"3D",X"41",X"38",X"5E",X"28",X"5E",X"38",X"5E",X"28",X"5E",X"23",X"41",X"23",X"5F",
		X"26",X"44",X"3A",X"44",X"16",X"5D",X"3C",X"5F",X"24",X"5F",X"0A",X"41",X"00",X"C0",X"02",X"44",
		X"3C",X"40",X"3E",X"42",X"38",X"41",X"26",X"5B",X"38",X"42",X"27",X"5B",X"23",X"5F",X"22",X"5E",
		X"28",X"42",X"3C",X"46",X"15",X"41",X"3C",X"40",X"23",X"5E",X"0A",X"5D",X"00",X"C0",X"03",X"43",
		X"3D",X"41",X"3F",X"43",X"39",X"44",X"24",X"59",X"39",X"44",X"24",X"59",X"23",X"5F",X"21",X"5D",
		X"27",X"5F",X"3F",X"47",X"17",X"45",X"3C",X"42",X"22",X"5C",X"08",X"5A",X"00",X"C0",X"04",X"42",
		X"3E",X"42",X"3F",X"43",X"3B",X"47",X"22",X"58",X"3B",X"46",X"21",X"58",X"22",X"5E",X"20",X"5C",
		X"26",X"5C",X"22",X"48",X"19",X"48",X"3E",X"43",X"20",X"5C",X"05",X"57",X"00",X"C0",X"04",X"40",
		X"3F",X"43",X"21",X"43",X"3E",X"48",X"3E",X"58",X"3E",X"48",X"3E",X"58",X"21",X"5D",X"3F",X"5D",
		X"24",X"5A",X"24",X"46",X"1B",X"4A",X"21",X"44",X"3F",X"5C",X"01",X"56",X"00",X"C0",X"04",X"5E",
		X"20",X"44",X"22",X"42",X"21",X"48",X"3B",X"5A",X"22",X"48",X"3B",X"59",X"3F",X"5D",X"3E",X"5E",
		X"22",X"58",X"26",X"44",X"01",X"4B",X"20",X"44",X"3E",X"5D",X"1D",X"56",X"00",X"C0",X"03",X"5D",
		X"21",X"43",X"23",X"41",X"24",X"47",X"39",X"5C",X"24",X"47",X"39",X"5C",X"3F",X"5D",X"3D",X"5F",
		X"3F",X"59",X"27",X"41",X"05",X"49",X"22",X"44",X"3C",X"5E",X"1A",X"58",X"00",X"C0",X"02",X"5C",
		X"22",X"42",X"23",X"41",X"27",X"45",X"38",X"5E",X"26",X"45",X"38",X"5F",X"3E",X"5E",X"3C",X"40",
		X"3C",X"5A",X"28",X"5E",X"08",X"47",X"23",X"42",X"3C",X"40",X"17",X"5B",X"00",X"C0",X"00",X"5C",
		X"23",X"41",X"23",X"5F",X"28",X"42",X"38",X"42",X"28",X"42",X"38",X"42",X"3D",X"5F",X"3D",X"41",
		X"3A",X"5C",X"26",X"5C",X"0A",X"43",X"24",X"41",X"3C",X"41",X"16",X"5F",X"00",X"C0",X"1E",X"5C",
		X"24",X"40",X"22",X"5E",X"28",X"5F",X"3A",X"45",X"28",X"5E",X"39",X"45",X"3D",X"41",X"3E",X"42",
		X"38",X"5E",X"24",X"5A",X"0B",X"5F",X"24",X"40",X"3D",X"42",X"16",X"43",X"00",X"C0",X"1D",X"5D",
		X"23",X"5F",X"21",X"5D",X"27",X"5C",X"3C",X"47",X"27",X"5C",X"3C",X"47",X"3D",X"41",X"3F",X"43",
		X"39",X"41",X"21",X"59",X"09",X"5B",X"24",X"5E",X"3E",X"44",X"18",X"46",X"00",X"C0",X"1C",X"5E",
		X"22",X"5E",X"21",X"5D",X"25",X"59",X"3E",X"48",X"25",X"5A",X"3F",X"48",X"3E",X"42",X"20",X"44",
		X"3A",X"44",X"3E",X"58",X"07",X"58",X"22",X"5D",X"20",X"44",X"1B",X"49",X"00",X"C0",X"1E",X"43",
		X"3E",X"5D",X"21",X"5D",X"3D",X"5B",X"20",X"5A",X"23",X"5E",X"26",X"40",X"23",X"42",X"20",X"46",
		X"3D",X"45",X"21",X"43",X"3E",X"43",X"01",X"5A",X"3A",X"40",X"03",X"53",X"20",X"4D",X"00",X"43",
		X"00",X"C0",X"1F",X"44",X"3D",X"5E",X"20",X"5C",X"3B",X"5D",X"3E",X"5A",X"22",X"5D",X"26",X"5E",
		X"23",X"41",X"22",X"45",X"20",X"46",X"22",X"42",X"3F",X"44",X"1F",X"5A",X"3A",X"42",X"1E",X"53",
		X"25",X"4C",X"01",X"43",X"00",X"C0",X"1F",X"44",X"3E",X"5F",X"3F",X"5D",X"3A",X"5F",X"3C",X"5B",
		X"21",X"5D",X"24",X"5C",X"23",X"5F",X"25",X"44",X"21",X"46",X"23",X"41",X"21",X"44",X"1C",X"5B",
		X"3C",X"44",X"19",X"55",X"29",X"49",X"02",X"42",X"00",X"C0",X"02",X"43",X"3C",X"41",X"3E",X"5E",
		X"3A",X"40",X"3B",X"5E",X"3F",X"5D",X"22",X"5A",X"23",X"5E",X"26",X"42",X"23",X"45",X"24",X"40",
		X"22",X"45",X"1A",X"5B",X"3E",X"46",X"15",X"58",X"2C",X"45",X"03",X"41",X"00",X"C0",X"03",X"42",
		X"3D",X"42",X"3D",X"5F",X"3B",X"43",X"3A",X"40",X"3E",X"5D",X"20",X"5A",X"22",X"5D",X"26",X"40",
		X"25",X"43",X"23",X"5F",X"23",X"42",X"1A",X"5F",X"20",X"46",X"13",X"5D",X"2D",X"40",X"03",X"40",
		X"00",X"C0",X"04",X"41",X"3E",X"43",X"3C",X"40",X"3D",X"45",X"3A",X"42",X"3D",X"5E",X"3E",X"5A",
		X"21",X"5D",X"25",X"5E",X"26",X"40",X"22",X"5E",X"24",X"41",X"1A",X"41",X"22",X"46",X"13",X"42",
		X"2C",X"5B",X"03",X"5F",X"00",X"C0",X"04",X"41",X"3F",X"42",X"3D",X"41",X"3F",X"46",X"3B",X"44",
		X"3D",X"5F",X"3C",X"5C",X"3F",X"5D",X"24",X"5B",X"26",X"5F",X"21",X"5D",X"22",X"5F",X"1D",X"44",
		X"24",X"44",X"15",X"47",X"29",X"57",X"02",X"5E",X"00",X"C0",X"03",X"5E",X"21",X"44",X"3E",X"42",
		X"20",X"46",X"3E",X"45",X"3D",X"41",X"3A",X"5E",X"3E",X"5D",X"22",X"5A",X"25",X"5D",X"20",X"5C",
		X"23",X"5E",X"1D",X"46",X"26",X"42",X"18",X"4B",X"25",X"54",X"01",X"5D",X"00",X"C0",X"02",X"5D",
		X"22",X"43",X"3F",X"43",X"23",X"45",X"20",X"46",X"3D",X"42",X"3A",X"40",X"3D",X"5E",X"20",X"5A",
		X"23",X"5B",X"3F",X"5D",X"22",X"5D",X"1F",X"46",X"26",X"40",X"1D",X"4D",X"20",X"53",X"00",X"5D",
		X"00",X"C0",X"1F",X"5C",X"25",X"42",X"20",X"44",X"25",X"43",X"22",X"46",X"3E",X"43",X"3A",X"42",
		X"3D",X"5F",X"3E",X"5B",X"20",X"5A",X"3E",X"5E",X"21",X"5C",X"01",X"46",X"26",X"5E",X"02",X"4D",
		X"3B",X"54",X"1F",X"5D",X"00",X"C0",X"1F",X"5C",X"24",X"41",X"21",X"43",X"26",X"41",X"24",X"45",
		X"3F",X"43",X"3C",X"44",X"3D",X"41",X"3B",X"5C",X"3F",X"5A",X"3D",X"5F",X"3F",X"5E",X"04",X"43",
		X"24",X"5C",X"07",X"4B",X"37",X"57",X"1E",X"5E",X"00",X"C0",X"1E",X"5D",X"24",X"5F",X"22",X"42",
		X"26",X"40",X"25",X"42",X"21",X"43",X"3E",X"46",X"3D",X"42",X"3A",X"5E",X"3D",X"5B",X"3C",X"40",
		X"3E",X"5D",X"06",X"43",X"22",X"5A",X"0B",X"48",X"34",X"5B",X"1D",X"5F",X"00",X"C0",X"1D",X"5E",
		X"23",X"5E",X"23",X"41",X"25",X"5D",X"26",X"40",X"22",X"43",X"20",X"46",X"3E",X"43",X"3A",X"40",
		X"3B",X"5D",X"3D",X"41",X"3D",X"5E",X"06",X"41",X"20",X"5A",X"0D",X"43",X"33",X"40",X"1D",X"40",
		X"00",X"C0",X"1C",X"41",X"22",X"5B",X"24",X"40",X"23",X"5B",X"26",X"5E",X"23",X"42",X"22",X"46",
		X"3F",X"43",X"3B",X"42",X"3A",X"40",X"3E",X"42",X"3C",X"5F",X"06",X"5F",X"3E",X"5A",X"0D",X"5E",
		X"34",X"45",X"1D",X"41",X"00",X"C0",X"1C",X"41",X"21",X"5C",X"23",X"5F",X"21",X"5A",X"25",X"5C",
		X"23",X"41",X"24",X"44",X"21",X"43",X"3C",X"45",X"3A",X"41",X"3F",X"43",X"3C",X"41",X"05",X"5C",
		X"3C",X"5C",X"0B",X"59",X"37",X"49",X"1E",X"42",X"00",X"C0",X"1D",X"42",X"3F",X"5C",X"22",X"5E",
		X"20",X"5A",X"22",X"5B",X"23",X"5F",X"26",X"42",X"22",X"43",X"3E",X"46",X"3B",X"43",X"20",X"44",
		X"3B",X"42",X"05",X"5A",X"3A",X"5E",X"08",X"55",X"3B",X"4C",X"1F",X"43",X"00",X"C0",X"00",X"4A",
		X"3A",X"56",X"24",X"40",X"20",X"5A",X"24",X"40",X"20",X"46",X"24",X"40",X"3A",X"4A",X"00",X"56",
		X"00",X"C0",X"04",X"49",X"36",X"59",X"24",X"5F",X"3E",X"5A",X"24",X"5F",X"22",X"47",X"24",X"5D",
		X"3E",X"4B",X"1C",X"57",X"00",X"C0",X"07",X"47",X"35",X"5D",X"23",X"5D",X"3B",X"5C",X"23",X"5D",
		X"24",X"45",X"23",X"5D",X"23",X"4B",X"19",X"59",X"00",X"C0",X"09",X"44",X"35",X"42",X"21",X"5C",
		X"3B",X"5E",X"21",X"5C",X"24",X"42",X"23",X"5C",X"27",X"4A",X"17",X"5C",X"00",X"C0",X"0A",X"40",
		X"36",X"46",X"20",X"5C",X"3A",X"40",X"20",X"5C",X"26",X"40",X"20",X"5C",X"2A",X"46",X"16",X"40",
		X"00",X"C0",X"09",X"5C",X"39",X"4A",X"3D",X"5C",X"3C",X"42",X"3F",X"5C",X"25",X"5E",X"3F",X"5C",
		X"2B",X"42",X"17",X"44",X"00",X"C0",X"07",X"59",X"3D",X"4B",X"3D",X"5D",X"3C",X"45",X"3D",X"5D",
		X"25",X"5C",X"3D",X"5D",X"2B",X"5D",X"19",X"47",X"00",X"C0",X"04",X"57",X"22",X"4B",X"3C",X"5F",
		X"3E",X"45",X"3C",X"5F",X"22",X"5C",X"3C",X"5D",X"2A",X"59",X"1C",X"49",X"00",X"C0",X"00",X"56",
		X"26",X"4A",X"3C",X"40",X"20",X"46",X"3C",X"40",X"20",X"5A",X"3C",X"40",X"26",X"56",X"00",X"4A",
		X"00",X"C0",X"1C",X"57",X"2A",X"47",X"3C",X"43",X"22",X"44",X"3C",X"41",X"3E",X"5B",X"3C",X"41",
		X"22",X"55",X"04",X"49",X"00",X"C0",X"19",X"59",X"2B",X"43",X"3D",X"43",X"25",X"44",X"3D",X"43",
		X"3C",X"5B",X"3D",X"43",X"3D",X"55",X"07",X"47",X"00",X"C0",X"17",X"5C",X"2B",X"5E",X"3D",X"44",
		X"27",X"42",X"3F",X"44",X"3A",X"5E",X"3F",X"44",X"39",X"56",X"09",X"44",X"00",X"C0",X"16",X"40",
		X"2A",X"5A",X"20",X"44",X"26",X"40",X"20",X"44",X"3A",X"40",X"20",X"44",X"36",X"5A",X"0A",X"40",
		X"00",X"C0",X"17",X"44",X"27",X"56",X"21",X"44",X"26",X"5E",X"21",X"44",X"39",X"42",X"23",X"44",
		X"35",X"5E",X"09",X"5C",X"00",X"C0",X"19",X"47",X"23",X"55",X"23",X"43",X"24",X"5B",X"23",X"43");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
