`define BUILD_DATE "180204"
`define BUILD_TIME "164559"
