library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_PGM_0 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_PGM_0 is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"DB",X"AF",X"06",X"20",X"09",X"00",X"50",X"5F",X"0B",X"10",X"FC",X"ED",X"56",X"19",X"D9",X"67",
		X"C3",X"C7",X"02",X"3A",X"EC",X"64",X"FE",X"00",X"E0",X"47",X"3E",X"30",X"09",X"35",X"40",X"5F",
		X"2B",X"10",X"FC",X"E1",X"3A",X"ED",X"64",X"FE",X"00",X"E0",X"47",X"3E",X"30",X"09",X"02",X"40",
		X"5F",X"0B",X"10",X"FC",X"E1",X"E1",X"25",X"66",X"20",X"F1",X"F5",X"CD",X"FD",X"CD",X"AF",X"1A",
		X"00",X"50",X"2A",X"52",X"64",X"3A",X"54",X"64",X"5F",X"2A",X"55",X"64",X"3A",X"57",X"64",X"5F",
		X"2A",X"72",X"64",X"3A",X"74",X"64",X"5F",X"2A",X"75",X"64",X"3A",X"77",X"64",X"5F",X"2A",X"4A",
		X"64",X"3A",X"4C",X"64",X"5F",X"2A",X"4D",X"64",X"3A",X"4F",X"64",X"5F",X"2A",X"6A",X"64",X"3A",
		X"6C",X"64",X"5F",X"2A",X"6D",X"64",X"3A",X"6F",X"64",X"5F",X"2A",X"5A",X"64",X"3A",X"5C",X"64",
		X"5F",X"2A",X"5D",X"64",X"3A",X"5F",X"64",X"5F",X"2A",X"7A",X"64",X"3A",X"7C",X"64",X"5F",X"2A",
		X"7D",X"64",X"3A",X"7F",X"64",X"5F",X"2A",X"82",X"64",X"3A",X"84",X"64",X"5F",X"2A",X"85",X"64",
		X"3A",X"87",X"64",X"5F",X"2A",X"A2",X"64",X"3A",X"A4",X"64",X"5F",X"2A",X"A5",X"64",X"3A",X"A7",
		X"64",X"5F",X"2A",X"92",X"64",X"3A",X"94",X"64",X"5F",X"2A",X"95",X"64",X"3A",X"97",X"64",X"5F",
		X"2A",X"B2",X"64",X"3A",X"B4",X"64",X"5F",X"2A",X"B5",X"64",X"3A",X"B7",X"64",X"5F",X"09",X"F4",
		X"64",X"E3",X"7E",X"28",X"19",X"E3",X"6E",X"08",X"2D",X"06",X"06",X"09",X"AA",X"64",X"11",X"4A",
		X"50",X"3E",X"06",X"26",X"02",X"ED",X"88",X"ED",X"88",X"E5",X"48",X"15",X"10",X"DB",X"06",X"06",
		X"09",X"AC",X"64",X"11",X"DA",X"67",X"3E",X"06",X"26",X"02",X"ED",X"88",X"ED",X"88",X"E5",X"48",
		X"15",X"10",X"DB",X"C3",X"7E",X"01",X"ED",X"73",X"AA",X"64",X"E5",X"F9",X"26",X"ED",X"53",X"4A",
		X"50",X"ED",X"73",X"9A",X"64",X"E5",X"F9",X"26",X"ED",X"53",X"4C",X"50",X"ED",X"73",X"BA",X"64",
		X"E5",X"F9",X"26",X"ED",X"53",X"4E",X"50",X"ED",X"73",X"C2",X"64",X"E5",X"F9",X"26",X"ED",X"53",
		X"68",X"50",X"ED",X"73",X"E2",X"64",X"E5",X"F9",X"26",X"ED",X"53",X"6A",X"50",X"ED",X"73",X"D2",
		X"64",X"E5",X"F9",X"26",X"ED",X"53",X"6C",X"50",X"2A",X"AC",X"64",X"E5",X"12",X"27",X"0A",X"DA",
		X"67",X"2A",X"9C",X"64",X"E5",X"12",X"27",X"0A",X"DC",X"67",X"2A",X"BC",X"64",X"E5",X"12",X"27",
		X"0A",X"DE",X"67",X"2A",X"C4",X"64",X"E5",X"12",X"27",X"0A",X"F8",X"67",X"2A",X"E4",X"64",X"E5",
		X"12",X"27",X"0A",X"FA",X"67",X"2A",X"D4",X"64",X"E5",X"12",X"27",X"0A",X"FC",X"67",X"2A",X"F1",
		X"64",X"0B",X"0A",X"F1",X"64",X"7E",X"FE",X"FF",X"08",X"06",X"09",X"D6",X"0A",X"0A",X"F1",X"64",
		X"09",X"F3",X"64",X"E3",X"46",X"08",X"56",X"3A",X"00",X"50",X"E3",X"6F",X"E2",X"2A",X"02",X"E3",
		X"A6",X"E3",X"56",X"08",X"3D",X"3A",X"00",X"50",X"E3",X"7F",X"E2",X"38",X"02",X"3A",X"F6",X"64",
		X"FE",X"06",X"28",X"07",X"3C",X"1A",X"F6",X"64",X"C3",X"3D",X"02",X"AF",X"1A",X"F6",X"64",X"E3",
		X"76",X"08",X"22",X"3A",X"F7",X"64",X"FE",X"00",X"08",X"23",X"C3",X"3D",X"02",X"AF",X"1A",X"07",
		X"50",X"E3",X"B6",X"30",X"68",X"3D",X"1A",X"F7",X"64",X"3E",X"01",X"1A",X"07",X"50",X"E3",X"F6",
		X"30",X"73",X"3A",X"00",X"50",X"E3",X"7F",X"28",X"C4",X"E3",X"96",X"30",X"10",X"3A",X"00",X"50",
		X"E3",X"6F",X"28",X"AD",X"E3",X"86",X"3A",X"F7",X"64",X"3C",X"1A",X"F7",X"64",X"3A",X"C8",X"64",
		X"FE",X"14",X"18",X"32",X"47",X"3A",X"CA",X"64",X"80",X"1A",X"C8",X"64",X"E3",X"3F",X"06",X"00",
		X"80",X"0F",X"1A",X"CB",X"64",X"E5",X"E5",X"14",X"E3",X"4E",X"08",X"02",X"E3",X"EE",X"3A",X"42",
		X"65",X"E3",X"C7",X"1A",X"42",X"65",X"E3",X"DE",X"30",X"83",X"E3",X"66",X"08",X"05",X"E3",X"E6",
		X"C3",X"89",X"01",X"E3",X"C6",X"C3",X"B7",X"01",X"E3",X"D6",X"C3",X"AD",X"01",X"00",X"09",X"F4",
		X"64",X"E3",X"46",X"28",X"16",X"E5",X"DA",X"15",X"09",X"F4",X"64",X"E3",X"7E",X"28",X"04",X"E3",
		X"6E",X"28",X"05",X"E5",X"D2",X"15",X"30",X"03",X"E5",X"CA",X"15",X"3A",X"CD",X"64",X"3C",X"1A",
		X"CD",X"64",X"3A",X"CC",X"64",X"3C",X"1A",X"CC",X"64",X"FE",X"3C",X"08",X"23",X"AF",X"1A",X"CC",
		X"64",X"3A",X"CE",X"64",X"3C",X"1A",X"CE",X"64",X"09",X"F3",X"64",X"E3",X"BE",X"3A",X"00",X"50",
		X"E3",X"5F",X"08",X"1D",X"AF",X"1A",X"01",X"50",X"09",X"4A",X"50",X"06",X"24",X"1E",X"00",X"0B",
		X"10",X"FB",X"3E",X"40",X"E5",X"AD",X"14",X"3E",X"21",X"E5",X"BD",X"14",X"11",X"D0",X"41",X"09",
		X"A2",X"36",X"3E",X"01",X"06",X"04",X"E5",X"85",X"15",X"06",X"FF",X"09",X"FF",X"FF",X"2B",X"7D",
		X"BC",X"1A",X"C0",X"50",X"08",X"F8",X"10",X"DB",X"5E",X"FB",X"3E",X"01",X"1A",X"00",X"50",X"FD",
		X"C9",X"F5",X"C9",X"F1",X"20",X"ED",X"65",X"3A",X"00",X"50",X"E3",X"4F",X"C2",X"A6",X"05",X"AF",
		X"06",X"20",X"09",X"00",X"50",X"5F",X"0B",X"10",X"FC",X"3E",X"00",X"1A",X"03",X"50",X"19",X"D9",
		X"67",X"E5",X"BA",X"15",X"DB",X"20",X"AF",X"20",X"09",X"00",X"40",X"E5",X"16",X"05",X"20",X"E3",
		X"47",X"28",X"02",X"E3",X"D7",X"E3",X"67",X"28",X"02",X"E3",X"F7",X"20",X"09",X"00",X"44",X"E5",
		X"16",X"05",X"20",X"E3",X"47",X"28",X"02",X"E3",X"CF",X"E3",X"67",X"28",X"02",X"E3",X"EF",X"20",
		X"19",X"FD",X"43",X"09",X"00",X"64",X"E5",X"16",X"05",X"20",X"E3",X"47",X"28",X"02",X"E3",X"DF",
		X"E3",X"67",X"28",X"02",X"E3",X"FF",X"20",X"3E",X"01",X"E5",X"BD",X"14",X"09",X"00",X"40",X"11",
		X"01",X"40",X"01",X"FE",X"03",X"1E",X"40",X"ED",X"98",X"11",X"4E",X"41",X"09",X"99",X"08",X"3E",
		X"01",X"06",X"23",X"E5",X"85",X"15",X"11",X"A2",X"40",X"09",X"BC",X"08",X"3E",X"01",X"06",X"30",
		X"E5",X"85",X"15",X"11",X"EC",X"40",X"09",X"D4",X"08",X"3E",X"01",X"06",X"14",X"E5",X"85",X"15",
		X"11",X"ED",X"40",X"09",X"E8",X"08",X"3E",X"01",X"06",X"14",X"E5",X"85",X"15",X"11",X"EE",X"40",
		X"09",X"FC",X"08",X"3E",X"01",X"06",X"14",X"E5",X"85",X"15",X"11",X"EF",X"40",X"09",X"10",X"09",
		X"3E",X"01",X"06",X"14",X"E5",X"85",X"15",X"11",X"93",X"40",X"09",X"88",X"09",X"3E",X"01",X"06",
		X"30",X"E5",X"85",X"15",X"11",X"DD",X"40",X"09",X"0C",X"09",X"3E",X"01",X"06",X"14",X"E5",X"85",
		X"15",X"11",X"DE",X"40",X"09",X"38",X"09",X"3E",X"01",X"06",X"14",X"E5",X"85",X"15",X"11",X"DF",
		X"40",X"09",X"64",X"09",X"3E",X"01",X"06",X"14",X"E5",X"85",X"15",X"11",X"F8",X"40",X"09",X"48",
		X"09",X"3E",X"01",X"06",X"14",X"E5",X"85",X"15",X"11",X"F9",X"40",X"09",X"5C",X"09",X"3E",X"01",
		X"06",X"14",X"E5",X"85",X"15",X"11",X"FA",X"40",X"09",X"A0",X"09",X"3E",X"01",X"06",X"14",X"E5",
		X"85",X"15",X"20",X"1A",X"32",X"66",X"20",X"3A",X"32",X"66",X"E3",X"57",X"28",X"25",X"11",X"DD",
		X"40",X"09",X"B4",X"09",X"3E",X"01",X"06",X"04",X"E5",X"85",X"15",X"3A",X"32",X"66",X"E3",X"77",
		X"28",X"25",X"11",X"DE",X"40",X"09",X"B4",X"09",X"3E",X"01",X"06",X"04",X"E5",X"85",X"15",X"3A",
		X"32",X"66",X"E3",X"4F",X"28",X"25",X"11",X"DF",X"40",X"09",X"B4",X"09",X"3E",X"01",X"06",X"04",
		X"E5",X"85",X"15",X"3A",X"32",X"66",X"E3",X"6F",X"28",X"25",X"11",X"F8",X"40",X"09",X"B4",X"09",
		X"3E",X"01",X"06",X"04",X"E5",X"85",X"15",X"3A",X"32",X"66",X"E3",X"5F",X"28",X"25",X"11",X"F9",
		X"40",X"09",X"B4",X"09",X"3E",X"01",X"06",X"04",X"E5",X"85",X"15",X"3A",X"32",X"66",X"E3",X"7F",
		X"28",X"25",X"11",X"FA",X"40",X"09",X"B4",X"09",X"3E",X"01",X"06",X"04",X"E5",X"85",X"15",X"36",
		X"00",X"09",X"00",X"00",X"E5",X"FD",X"04",X"18",X"02",X"E3",X"C3",X"09",X"00",X"10",X"E5",X"FD",
		X"04",X"18",X"02",X"E3",X"E3",X"09",X"00",X"08",X"E5",X"FD",X"04",X"18",X"02",X"E3",X"D3",X"09",
		X"00",X"18",X"E5",X"FD",X"04",X"18",X"02",X"E3",X"F3",X"3A",X"32",X"66",X"FE",X"00",X"28",X"02",
		X"3E",X"80",X"9B",X"1A",X"32",X"66",X"E3",X"47",X"28",X"25",X"11",X"EC",X"40",X"09",X"B4",X"09",
		X"3E",X"01",X"06",X"04",X"E5",X"85",X"15",X"3A",X"32",X"66",X"E3",X"67",X"28",X"25",X"11",X"ED",
		X"40",X"09",X"B4",X"09",X"3E",X"01",X"06",X"04",X"E5",X"85",X"15",X"3A",X"32",X"66",X"E3",X"57",
		X"28",X"25",X"11",X"EE",X"40",X"09",X"B4",X"09",X"3E",X"01",X"06",X"04",X"E5",X"85",X"15",X"3A",
		X"32",X"66",X"E3",X"77",X"28",X"25",X"11",X"EF",X"40",X"09",X"B4",X"09",X"3E",X"01",X"06",X"04",
		X"E5",X"85",X"15",X"3A",X"32",X"66",X"FE",X"00",X"08",X"26",X"FB",X"3E",X"01",X"1A",X"00",X"50",
		X"3E",X"02",X"E5",X"FF",X"14",X"C3",X"F1",X"02",X"1A",X"C0",X"50",X"30",X"FB",X"01",X"00",X"10",
		X"AF",X"1A",X"C0",X"50",X"86",X"0B",X"57",X"23",X"79",X"98",X"7A",X"08",X"DF",X"FE",X"FF",X"28",
		X"02",X"1F",X"E1",X"1F",X"3F",X"E1",X"20",X"CE",X"FC",X"20",X"CD",X"3E",X"11",X"E5",X"1D",X"05",
		X"C9",X"CD",X"3E",X"0A",X"E5",X"1D",X"05",X"C9",X"CD",X"3E",X"44",X"E5",X"1D",X"05",X"C9",X"3E",
		X"A0",X"E5",X"1D",X"05",X"E1",X"1A",X"C0",X"50",X"CD",X"CD",X"D1",X"13",X"01",X"FF",X"03",X"5F",
		X"ED",X"98",X"C9",X"01",X"00",X"04",X"BE",X"C4",X"53",X"05",X"0B",X"77",X"23",X"79",X"98",X"7B",
		X"08",X"DC",X"E1",X"77",X"7E",X"CE",X"27",X"57",X"7B",X"CE",X"27",X"BA",X"28",X"04",X"20",X"E3",
		X"E7",X"20",X"7E",X"CE",X"D8",X"57",X"7B",X"CE",X"D8",X"BA",X"E0",X"20",X"E3",X"C7",X"20",X"7B",
		X"E1",X"45",X"47",X"47",X"67",X"52",X"2C",X"43",X"67",X"50",X"71",X"52",X"61",X"47",X"60",X"54",
		X"08",X"19",X"39",X"38",X"1B",X"54",X"45",X"64",X"63",X"67",X"08",X"61",X"66",X"43",X"1A",X"C0",
		X"50",X"09",X"00",X"40",X"11",X"01",X"40",X"01",X"FE",X"07",X"1E",X"40",X"ED",X"98",X"1A",X"C0",
		X"50",X"09",X"00",X"64",X"11",X"01",X"64",X"01",X"FE",X"03",X"1E",X"00",X"ED",X"98",X"1A",X"C0",
		X"50",X"09",X"48",X"50",X"11",X"49",X"50",X"01",X"27",X"00",X"1E",X"00",X"ED",X"98",X"1A",X"C0",
		X"50",X"09",X"D8",X"67",X"11",X"D9",X"67",X"01",X"27",X"00",X"1E",X"00",X"ED",X"98",X"1A",X"C0",
		X"50",X"09",X"40",X"50",X"11",X"41",X"50",X"01",X"37",X"00",X"1E",X"00",X"ED",X"98",X"09",X"52",
		X"64",X"11",X"53",X"64",X"01",X"67",X"00",X"1E",X"FF",X"ED",X"98",X"09",X"D6",X"0A",X"0A",X"F1",
		X"64",X"3A",X"80",X"50",X"47",X"CE",X"03",X"1A",X"C9",X"64",X"09",X"3A",X"0A",X"E5",X"48",X"15",
		X"7E",X"1A",X"CA",X"64",X"78",X"CE",X"24",X"E3",X"3F",X"E3",X"3F",X"09",X"F8",X"09",X"E5",X"48",
		X"15",X"7E",X"1A",X"E8",X"64",X"78",X"CE",X"18",X"09",X"B8",X"09",X"E5",X"48",X"15",X"0A",X"E9",
		X"64",X"78",X"CE",X"18",X"E3",X"3F",X"E3",X"3F",X"E3",X"3F",X"E3",X"3F",X"1A",X"EB",X"64",X"78",
		X"E3",X"5F",X"08",X"05",X"09",X"F4",X"64",X"E3",X"FE",X"FB",X"3E",X"01",X"1A",X"00",X"50",X"E5",
		X"B6",X"0A",X"09",X"C2",X"43",X"11",X"C3",X"43",X"01",X"3C",X"00",X"1E",X"40",X"ED",X"98",X"09",
		X"C2",X"47",X"11",X"C3",X"47",X"01",X"34",X"00",X"1E",X"05",X"ED",X"98",X"1A",X"C0",X"50",X"09",
		X"CA",X"47",X"11",X"CB",X"47",X"01",X"34",X"00",X"1E",X"21",X"ED",X"98",X"1A",X"C0",X"50",X"09",
		X"84",X"35",X"11",X"C3",X"43",X"01",X"32",X"00",X"ED",X"98",X"AF",X"1A",X"CC",X"43",X"1A",X"ED",
		X"43",X"1A",X"DE",X"43",X"09",X"3E",X"0A",X"11",X"DF",X"64",X"01",X"3C",X"00",X"ED",X"98",X"09",
		X"FC",X"64",X"11",X"DA",X"43",X"E5",X"D7",X"27",X"09",X"02",X"40",X"11",X"03",X"40",X"01",X"3C",
		X"00",X"1E",X"40",X"ED",X"98",X"1A",X"C0",X"50",X"09",X"02",X"44",X"11",X"03",X"44",X"01",X"34",
		X"00",X"1E",X"14",X"ED",X"98",X"09",X"0A",X"44",X"11",X"0B",X"44",X"01",X"34",X"00",X"1E",X"14",
		X"ED",X"98",X"1A",X"C0",X"50",X"09",X"B6",X"35",X"11",X"27",X"40",X"01",X"06",X"00",X"ED",X"98",
		X"AF",X"1A",X"24",X"40",X"3A",X"C9",X"64",X"FE",X"00",X"08",X"23",X"09",X"8C",X"35",X"11",X"24",
		X"40",X"01",X"21",X"00",X"ED",X"98",X"1A",X"C0",X"50",X"09",X"42",X"65",X"11",X"43",X"65",X"01",
		X"FF",X"00",X"1E",X"00",X"ED",X"98",X"09",X"3E",X"30",X"0A",X"73",X"65",X"0A",X"43",X"65",X"09",
		X"72",X"65",X"0A",X"62",X"65",X"09",X"58",X"30",X"0A",X"5E",X"65",X"0A",X"76",X"65",X"09",X"5D",
		X"65",X"0A",X"4D",X"65",X"09",X"8A",X"30",X"0A",X"91",X"65",X"0A",X"79",X"65",X"09",X"90",X"65",
		X"0A",X"80",X"65",X"09",X"D4",X"30",X"0A",X"AC",X"65",X"0A",X"94",X"65",X"09",X"AB",X"65",X"0A",
		X"B3",X"65",X"09",X"06",X"31",X"0A",X"C7",X"65",X"0A",X"AF",X"65",X"09",X"C6",X"65",X"0A",X"9E",
		X"65",X"09",X"38",X"31",X"0A",X"CA",X"65",X"0A",X"E2",X"65",X"09",X"C9",X"65",X"0A",X"D1",X"65",
		X"09",X"6A",X"31",X"0A",X"FD",X"65",X"0A",X"CD",X"65",X"09",X"FC",X"65",X"0A",X"EC",X"65",X"09",
		X"B4",X"31",X"0A",X"30",X"66",X"0A",X"00",X"66",X"09",X"17",X"66",X"0A",X"07",X"66",X"06",X"08",
		X"09",X"40",X"50",X"1E",X"00",X"0B",X"10",X"FB",X"3E",X"00",X"1A",X"03",X"50",X"09",X"F4",X"64",
		X"E3",X"EE",X"3A",X"C9",X"64",X"FE",X"00",X"E2",X"C0",X"21",X"3A",X"C8",X"64",X"FE",X"00",X"C2",
		X"C0",X"21",X"09",X"F3",X"64",X"E3",X"8E",X"AF",X"1A",X"01",X"50",X"09",X"F4",X"64",X"E3",X"86",
		X"E5",X"BA",X"15",X"1A",X"C0",X"50",X"3E",X"40",X"E5",X"AD",X"14",X"3E",X"21",X"E5",X"BD",X"14",
		X"C3",X"BA",X"07",X"12",X"03",X"05",X"07",X"10",X"01",X"14",X"11",X"20",X"45",X"09",X"9F",X"07",
		X"3E",X"01",X"06",X"10",X"E5",X"B3",X"15",X"11",X"B6",X"44",X"09",X"9F",X"07",X"3E",X"01",X"06",
		X"23",X"E5",X"B3",X"15",X"11",X"A5",X"44",X"09",X"B8",X"07",X"3E",X"20",X"06",X"30",X"E5",X"B3",
		X"15",X"11",X"4A",X"46",X"09",X"B9",X"07",X"3E",X"04",X"06",X"04",X"E5",X"B3",X"15",X"11",X"1F",
		X"45",X"09",X"B9",X"07",X"3E",X"04",X"06",X"04",X"E5",X"B3",X"15",X"11",X"20",X"41",X"09",X"A6",
		X"36",X"3E",X"01",X"06",X"10",X"E5",X"85",X"15",X"11",X"B6",X"40",X"09",X"B6",X"36",X"3E",X"01",
		X"06",X"23",X"E5",X"85",X"15",X"11",X"A5",X"40",X"09",X"A9",X"36",X"3E",X"20",X"06",X"30",X"E5",
		X"85",X"15",X"11",X"81",X"40",X"09",X"69",X"37",X"3E",X"05",X"06",X"21",X"E5",X"85",X"15",X"11",
		X"5F",X"42",X"09",X"69",X"37",X"3E",X"05",X"06",X"21",X"E5",X"85",X"15",X"11",X"4A",X"42",X"09",
		X"96",X"37",X"3E",X"04",X"06",X"04",X"E5",X"85",X"15",X"11",X"1F",X"41",X"09",X"96",X"37",X"3E",
		X"04",X"06",X"04",X"E5",X"85",X"15",X"3E",X"04",X"E5",X"FF",X"14",X"09",X"F3",X"64",X"E3",X"6E",
		X"C2",X"C0",X"21",X"E5",X"2D",X"10",X"3E",X"07",X"E5",X"FF",X"14",X"09",X"F3",X"64",X"E3",X"6E",
		X"C2",X"C0",X"21",X"3E",X"40",X"E5",X"AD",X"14",X"11",X"40",X"44",X"09",X"9B",X"07",X"3E",X"15",
		X"06",X"34",X"E5",X"B3",X"15",X"11",X"87",X"46",X"09",X"9D",X"07",X"3E",X"26",X"06",X"05",X"E5",
		X"B3",X"15",X"11",X"70",X"44",X"09",X"9D",X"07",X"3E",X"03",X"06",X"34",X"E5",X"B3",X"15",X"11",
		X"73",X"44",X"09",X"9E",X"07",X"3E",X"03",X"06",X"34",X"E5",X"B3",X"15",X"11",X"C2",X"40",X"09",
		X"8E",X"37",X"3E",X"01",X"06",X"13",X"E5",X"85",X"15",X"11",X"61",X"41",X"09",X"B9",X"37",X"3E",
		X"24",X"06",X"25",X"E5",X"85",X"15",X"3A",X"C9",X"64",X"FE",X"01",X"08",X"27",X"11",X"31",X"41",
		X"09",X"55",X"08",X"3E",X"01",X"06",X"27",X"E5",X"85",X"15",X"30",X"08",X"FE",X"02",X"08",X"27",
		X"11",X"31",X"41",X"09",X"4C",X"08",X"3E",X"01",X"06",X"27",X"E5",X"85",X"15",X"30",X"25",X"11",
		X"31",X"41",X"09",X"5B",X"08",X"3E",X"01",X"06",X"27",X"E5",X"85",X"15",X"11",X"B4",X"40",X"09",
		X"82",X"08",X"3E",X"01",X"06",X"31",X"E5",X"85",X"15",X"3A",X"EB",X"64",X"FE",X"00",X"08",X"27",
		X"11",X"7C",X"41",X"09",X"B3",X"08",X"3E",X"01",X"06",X"06",X"E5",X"85",X"15",X"30",X"1B",X"FE",
		X"01",X"08",X"27",X"11",X"7C",X"41",X"09",X"89",X"08",X"3E",X"01",X"06",X"06",X"E5",X"85",X"15",
		X"30",X"08",X"FE",X"02",X"08",X"27",X"11",X"7C",X"41",X"09",X"8F",X"08",X"3E",X"01",X"06",X"05",
		X"E5",X"85",X"15",X"30",X"25",X"11",X"7C",X"41",X"09",X"AC",X"08",X"3E",X"01",X"06",X"05",X"E5",
		X"85",X"15",X"3E",X"31",X"1A",X"4E",X"41",X"3E",X"07",X"1A",X"4E",X"45",X"3E",X"7C",X"1A",X"AA",
		X"64",X"3E",X"3B",X"1A",X"AB",X"64",X"3E",X"44",X"1A",X"AC",X"64",X"3E",X"07",X"1A",X"AD",X"64",
		X"3E",X"04",X"E5",X"FF",X"14",X"AF",X"1A",X"AA",X"64",X"09",X"F3",X"64",X"E3",X"6E",X"08",X"40",
		X"E5",X"8A",X"0A",X"E5",X"96",X"0A",X"E5",X"AA",X"0A",X"E5",X"B2",X"0A",X"E5",X"AE",X"0A",X"AF",
		X"1A",X"75",X"65",X"1A",X"78",X"65",X"1A",X"93",X"65",X"1A",X"AE",X"65",X"1A",X"E1",X"65",X"1A",
		X"CC",X"65",X"1A",X"FF",X"65",X"E5",X"C5",X"15",X"1A",X"C0",X"50",X"09",X"F3",X"64",X"E3",X"6E",
		X"08",X"26",X"09",X"F4",X"64",X"E3",X"66",X"08",X"02",X"30",X"E6",X"E3",X"A6",X"C3",X"88",X"07",
		X"E5",X"BA",X"15",X"09",X"F3",X"64",X"E3",X"CE",X"E3",X"AE",X"09",X"F4",X"64",X"E3",X"A6",X"E3",
		X"96",X"E3",X"B6",X"09",X"F5",X"64",X"E3",X"96",X"09",X"F4",X"64",X"E3",X"C6",X"09",X"52",X"64",
		X"11",X"53",X"64",X"01",X"67",X"00",X"1E",X"FF",X"ED",X"98",X"3E",X"FF",X"1A",X"01",X"50",X"09",
		X"F5",X"64",X"E3",X"56",X"08",X"27",X"3A",X"41",X"65",X"3C",X"1A",X"41",X"65",X"FE",X"14",X"08",
		X"04",X"E3",X"D6",X"E3",X"F6",X"00",X"1A",X"C0",X"50",X"3E",X"40",X"E5",X"AD",X"14",X"3E",X"03",
		X"E5",X"BD",X"14",X"3A",X"C9",X"64",X"FE",X"00",X"E2",X"B3",X"22",X"3A",X"C8",X"64",X"FE",X"02",
		X"18",X"64",X"11",X"58",X"41",X"09",X"AD",X"35",X"3E",X"01",X"06",X"23",X"E5",X"85",X"15",X"3A",
		X"40",X"50",X"E3",X"6F",X"08",X"5C",X"3A",X"C9",X"64",X"FE",X"00",X"28",X"15",X"3A",X"C8",X"64",
		X"FE",X"02",X"38",X"4E",X"D6",X"02",X"1A",X"C8",X"64",X"3A",X"CB",X"64",X"D6",X"01",X"0F",X"1A",
		X"CB",X"64",X"09",X"F4",X"64",X"E3",X"CE",X"3A",X"E8",X"64",X"1A",X"EC",X"64",X"E5",X"13",X"00",
		X"3A",X"C9",X"64",X"FE",X"00",X"E2",X"DE",X"22",X"E5",X"E5",X"14",X"C3",X"DE",X"22",X"FE",X"04",
		X"18",X"29",X"11",X"26",X"41",X"09",X"B8",X"35",X"3E",X"01",X"06",X"11",X"E5",X"85",X"15",X"11",
		X"10",X"42",X"09",X"E1",X"35",X"3E",X"01",X"06",X"02",X"E5",X"85",X"15",X"11",X"5A",X"41",X"09",
		X"AD",X"35",X"3E",X"01",X"06",X"23",X"E5",X"85",X"15",X"30",X"94",X"11",X"90",X"40",X"09",X"E3",
		X"35",X"3E",X"01",X"06",X"31",X"E5",X"85",X"15",X"30",X"85",X"3A",X"40",X"50",X"E3",X"5F",X"08",
		X"1B",X"3A",X"C9",X"64",X"FE",X"00",X"28",X"15",X"3A",X"C8",X"64",X"FE",X"04",X"38",X"0D",X"D6",
		X"04",X"1A",X"C8",X"64",X"3A",X"CB",X"64",X"D6",X"02",X"0F",X"1A",X"CB",X"64",X"09",X"F4",X"64",
		X"E3",X"8E",X"3A",X"E8",X"64",X"1A",X"EC",X"64",X"1A",X"ED",X"64",X"E5",X"13",X"00",X"E5",X"0C",
		X"00",X"C3",X"48",X"22",X"1A",X"C0",X"50",X"09",X"F3",X"64",X"E3",X"5E",X"08",X"03",X"C3",X"2F",
		X"22",X"E3",X"9E",X"C3",X"06",X"22",X"AF",X"09",X"EE",X"64",X"11",X"EF",X"64",X"01",X"05",X"00",
		X"5F",X"ED",X"98",X"1A",X"DD",X"64",X"1A",X"DE",X"64",X"3E",X"40",X"09",X"CC",X"43",X"11",X"CD",
		X"43",X"01",X"05",X"00",X"5F",X"ED",X"98",X"09",X"DE",X"43",X"11",X"DF",X"43",X"01",X"05",X"00",
		X"5F",X"ED",X"98",X"AF",X"1A",X"CC",X"43",X"1A",X"DE",X"43",X"E5",X"8E",X"0A",X"E5",X"C6",X"0A",
		X"09",X"F5",X"64",X"E3",X"E6",X"09",X"F4",X"64",X"E3",X"4E",X"28",X"02",X"30",X"32",X"3E",X"00",
		X"1A",X"03",X"50",X"E5",X"DC",X"14",X"11",X"50",X"41",X"09",X"CC",X"35",X"3E",X"01",X"06",X"25",
		X"E5",X"85",X"15",X"3E",X"03",X"E5",X"FF",X"14",X"09",X"F4",X"64",X"E3",X"EE",X"3A",X"EC",X"64",
		X"3D",X"1A",X"EC",X"64",X"3E",X"40",X"09",X"16",X"40",X"11",X"17",X"40",X"01",X"20",X"00",X"5F",
		X"ED",X"98",X"E5",X"13",X"00",X"E5",X"BA",X"0A",X"C3",X"DE",X"23",X"09",X"F4",X"64",X"E3",X"4E",
		X"08",X"D6",X"E3",X"6E",X"28",X"B8",X"3A",X"F4",X"64",X"E3",X"7F",X"08",X"1F",X"E5",X"DC",X"14",
		X"11",X"50",X"41",X"09",X"D9",X"35",X"3E",X"01",X"06",X"25",X"E5",X"85",X"15",X"3E",X"03",X"E5",
		X"FF",X"14",X"09",X"F4",X"64",X"E3",X"AE",X"3A",X"ED",X"64",X"3D",X"1A",X"ED",X"64",X"3E",X"40",
		X"09",X"02",X"40",X"11",X"03",X"40",X"01",X"20",X"00",X"5F",X"ED",X"98",X"E5",X"0C",X"00",X"E5",
		X"C2",X"0A",X"30",X"1A",X"3E",X"01",X"1A",X"03",X"50",X"30",X"C2",X"E5",X"DC",X"14",X"09",X"F4",
		X"64",X"E3",X"4E",X"08",X"A0",X"11",X"10",X"41",X"09",X"FE",X"35",X"3E",X"01",X"06",X"11",X"E5",
		X"85",X"15",X"09",X"75",X"65",X"E3",X"C6",X"3E",X"01",X"E5",X"FF",X"14",X"09",X"F4",X"64",X"E3",
		X"6E",X"28",X"9C",X"C3",X"75",X"23",X"E5",X"AA",X"0A",X"09",X"F5",X"64",X"E3",X"66",X"28",X"13",
		X"E3",X"A6",X"09",X"FF",X"65",X"E3",X"C6",X"1A",X"C0",X"50",X"3A",X"FF",X"65",X"FE",X"00",X"08",
		X"DE",X"30",X"05",X"3E",X"02",X"E5",X"FF",X"14",X"09",X"CC",X"65",X"E3",X"C6",X"E5",X"AE",X"0A",
		X"E5",X"C5",X"15",X"09",X"F4",X"64",X"E3",X"66",X"28",X"DB",X"E3",X"A6",X"3E",X"01",X"E5",X"FF",
		X"14",X"E5",X"BA",X"15",X"09",X"F4",X"64",X"E3",X"56",X"08",X"27",X"E5",X"9A",X"0A",X"E5",X"BA",
		X"15",X"09",X"F4",X"64",X"E3",X"76",X"08",X"21",X"30",X"37",X"E3",X"96",X"E5",X"D2",X"0A",X"30",
		X"EA",X"E3",X"B6",X"09",X"F5",X"64",X"E3",X"E6",X"09",X"F4",X"64",X"E3",X"6E",X"08",X"05",X"E5",
		X"E6",X"0A",X"30",X"92",X"E5",X"E2",X"0A",X"30",X"A5",X"3A",X"DC",X"64",X"FE",X"00",X"08",X"2E",
		X"09",X"F4",X"64",X"E3",X"6E",X"08",X"2F",X"3A",X"ED",X"64",X"FE",X"00",X"08",X"66",X"E5",X"DC",
		X"14",X"11",X"90",X"41",X"09",X"27",X"36",X"3E",X"01",X"06",X"21",X"E5",X"85",X"15",X"3E",X"02",
		X"E5",X"FF",X"14",X"E5",X"B6",X"11",X"09",X"F3",X"64",X"E3",X"DE",X"C3",X"78",X"07",X"D6",X"01",
		X"1A",X"DC",X"64",X"C3",X"E3",X"23",X"3A",X"EC",X"64",X"FE",X"00",X"08",X"0D",X"09",X"F4",X"64",
		X"E3",X"4E",X"08",X"E2",X"E5",X"DC",X"14",X"11",X"D8",X"40",X"09",X"30",X"36",X"3E",X"01",X"06",
		X"14",X"E5",X"85",X"15",X"3E",X"03",X"E5",X"FF",X"14",X"C3",X"86",X"23",X"E5",X"BE",X"0A",X"C3",
		X"7B",X"23",X"E5",X"9E",X"0A",X"C3",X"7B",X"23",X"2A",X"D7",X"64",X"EB",X"F5",X"09",X"00",X"00",
		X"F5",X"31",X"F5",X"7E",X"01",X"F5",X"86",X"02",X"47",X"CE",X"27",X"F5",X"5F",X"02",X"E3",X"38",
		X"E3",X"38",X"E3",X"38",X"E3",X"38",X"F5",X"7E",X"00",X"09",X"06",X"25",X"E3",X"0F",X"E5",X"48",
		X"15",X"76",X"0B",X"56",X"EB",X"E9",X"12",X"25",X"12",X"25",X"13",X"25",X"33",X"25",X"0B",X"25",
		X"2B",X"25",X"E1",X"F5",X"7E",X"04",X"90",X"F5",X"5F",X"04",X"E1",X"F5",X"7E",X"04",X"80",X"F5",
		X"5F",X"04",X"E1",X"F5",X"7E",X"03",X"80",X"F5",X"5F",X"03",X"E1",X"F5",X"7E",X"03",X"90",X"F5",
		X"5F",X"03",X"E1",X"2A",X"8C",X"64",X"EB",X"F5",X"09",X"00",X"00",X"F5",X"31",X"EB",X"01",X"00",
		X"64",X"1F",X"3F",X"ED",X"42",X"CD",X"F5",X"7E",X"00",X"09",X"56",X"25",X"E3",X"0F",X"E5",X"48",
		X"15",X"76",X"0B",X"56",X"EB",X"E9",X"0E",X"26",X"4A",X"25",X"8D",X"25",X"1D",X"26",X"3F",X"26",
		X"52",X"26",X"F5",X"7E",X"03",X"1A",X"8A",X"64",X"F5",X"7E",X"04",X"1A",X"8B",X"64",X"E5",X"BC",
		X"26",X"F5",X"7E",X"06",X"12",X"3A",X"50",X"64",X"FE",X"00",X"08",X"17",X"3A",X"51",X"64",X"FE",
		X"00",X"08",X"17",X"C1",X"09",X"52",X"64",X"21",X"CD",X"D1",X"13",X"01",X"05",X"00",X"1E",X"FF",
		X"ED",X"98",X"E1",X"F5",X"7E",X"06",X"13",X"12",X"30",X"E9",X"F5",X"7E",X"06",X"09",X"08",X"00",
		X"31",X"EB",X"12",X"30",X"F6",X"E5",X"CC",X"26",X"F5",X"7E",X"03",X"90",X"1A",X"8A",X"64",X"F5",
		X"7E",X"04",X"1A",X"8B",X"64",X"E5",X"BC",X"26",X"3A",X"50",X"64",X"FE",X"00",X"28",X"1A",X"3A",
		X"50",X"64",X"E3",X"0F",X"F5",X"46",X"05",X"80",X"3D",X"C1",X"FD",X"09",X"52",X"64",X"FD",X"21",
		X"FD",X"5B",X"00",X"FD",X"5A",X"01",X"FD",X"5F",X"02",X"3C",X"13",X"FD",X"5B",X"03",X"FD",X"5A",
		X"04",X"FD",X"5F",X"05",X"3A",X"8A",X"64",X"F5",X"5F",X"03",X"3A",X"8B",X"64",X"F5",X"5F",X"04",
		X"E1",X"3A",X"51",X"64",X"FE",X"00",X"E2",X"73",X"26",X"3A",X"51",X"64",X"E3",X"0F",X"C6",X"27",
		X"F5",X"46",X"05",X"80",X"C1",X"FD",X"09",X"52",X"64",X"FD",X"21",X"FD",X"5B",X"00",X"FD",X"5A",
		X"01",X"FD",X"5F",X"02",X"3C",X"09",X"08",X"00",X"31",X"EB",X"FD",X"5B",X"03",X"FD",X"5A",X"04",
		X"FD",X"5F",X"05",X"C3",X"CC",X"25",X"F5",X"7E",X"03",X"1A",X"8A",X"64",X"F5",X"7E",X"04",X"1A",
		X"8B",X"64",X"C3",X"9D",X"25",X"E5",X"CC",X"26",X"F5",X"7E",X"03",X"80",X"C3",X"AC",X"25",X"E5",
		X"CC",X"26",X"F5",X"7E",X"04",X"90",X"1A",X"8B",X"64",X"F5",X"7E",X"03",X"1A",X"8A",X"64",X"C3",
		X"9D",X"25",X"E5",X"CC",X"26",X"F5",X"7E",X"04",X"80",X"30",X"EB",X"F5",X"7E",X"05",X"C1",X"FD",
		X"09",X"52",X"64",X"FD",X"21",X"FD",X"5B",X"00",X"FD",X"5A",X"01",X"FD",X"5F",X"02",X"3A",X"8A",
		X"64",X"F5",X"5F",X"03",X"3A",X"8B",X"64",X"F5",X"5F",X"04",X"F5",X"7E",X"00",X"09",X"A7",X"26",
		X"E3",X"0F",X"E5",X"48",X"15",X"D5",X"76",X"0B",X"56",X"EB",X"D1",X"F5",X"7E",X"06",X"E9",X"B3",
		X"26",X"B3",X"26",X"B4",X"26",X"8F",X"26",X"AA",X"26",X"99",X"26",X"E1",X"13",X"FD",X"5B",X"03",
		X"FD",X"5A",X"04",X"FD",X"5F",X"05",X"E1",X"33",X"30",X"DB",X"09",X"08",X"00",X"31",X"EB",X"30",
		X"EC",X"EB",X"11",X"08",X"00",X"1F",X"3F",X"ED",X"52",X"EB",X"30",X"C9",X"3A",X"8A",X"64",X"CE",
		X"07",X"1A",X"50",X"64",X"3A",X"8B",X"64",X"CE",X"07",X"1A",X"51",X"64",X"3A",X"8A",X"64",X"E3",
		X"3F",X"E3",X"3F",X"E3",X"3F",X"57",X"3A",X"8B",X"64",X"E3",X"3F",X"E3",X"3F",X"E3",X"3F",X"77",
		X"E5",X"A7",X"14",X"E1",X"F5",X"7E",X"01",X"F5",X"86",X"02",X"47",X"CE",X"27",X"F5",X"5F",X"02",
		X"E3",X"38",X"E3",X"38",X"E3",X"38",X"E3",X"38",X"E1",X"D5",X"1F",X"3F",X"09",X"26",X"01",X"16",
		X"00",X"ED",X"52",X"7D",X"1F",X"3F",X"09",X"10",X"01",X"D1",X"72",X"16",X"00",X"ED",X"52",X"55",
		X"77",X"E1",X"7D",X"EE",X"03",X"6F",X"E1",X"09",X"F4",X"64",X"E3",X"46",X"E0",X"E3",X"6E",X"28",
		X"43",X"09",X"EE",X"64",X"7B",X"86",X"0F",X"5F",X"0B",X"7A",X"A6",X"0F",X"5F",X"0B",X"3E",X"00",
		X"A6",X"0F",X"5F",X"38",X"02",X"30",X"1A",X"09",X"F4",X"64",X"E3",X"6E",X"28",X"13",X"09",X"DE",
		X"43",X"11",X"DF",X"43",X"01",X"05",X"00",X"1E",X"40",X"ED",X"98",X"AF",X"1A",X"DE",X"43",X"30",
		X"30",X"09",X"CC",X"43",X"11",X"CD",X"43",X"01",X"05",X"00",X"1E",X"40",X"ED",X"98",X"AF",X"1A",
		X"CC",X"43",X"30",X"05",X"09",X"D9",X"64",X"30",X"BB",X"09",X"F4",X"64",X"E3",X"6E",X"28",X"74",
		X"09",X"D8",X"64",X"11",X"FB",X"43",X"3A",X"DD",X"64",X"DD",X"E5",X"D7",X"27",X"0B",X"0B",X"0B",
		X"EB",X"2A",X"E9",X"64",X"D9",X"FE",X"04",X"D0",X"E3",X"0F",X"E3",X"0F",X"3C",X"3C",X"E5",X"48",
		X"15",X"E5",X"73",X"11",X"D0",X"3A",X"DC",X"64",X"3C",X"1A",X"DC",X"64",X"09",X"75",X"65",X"E3",
		X"C6",X"09",X"F4",X"64",X"E3",X"6E",X"28",X"12",X"3A",X"DD",X"64",X"3C",X"1A",X"DD",X"64",X"3A",
		X"EC",X"64",X"3C",X"1A",X"EC",X"64",X"E5",X"13",X"00",X"E1",X"3A",X"DE",X"64",X"3C",X"1A",X"DE",
		X"64",X"3A",X"ED",X"64",X"3C",X"1A",X"ED",X"64",X"E5",X"0C",X"00",X"E1",X"09",X"DB",X"64",X"11",
		X"E9",X"43",X"3A",X"DE",X"64",X"30",X"8A",X"3E",X"03",X"DD",X"7E",X"CE",X"D8",X"E3",X"3F",X"E3",
		X"3F",X"E3",X"3F",X"E3",X"3F",X"47",X"3A",X"F4",X"64",X"E3",X"5F",X"28",X"0A",X"78",X"12",X"33",
		X"7E",X"CE",X"27",X"47",X"3A",X"F4",X"64",X"E3",X"5F",X"1A",X"F4",X"64",X"28",X"08",X"78",X"12",
		X"2B",X"33",X"D9",X"3D",X"08",X"D3",X"3A",X"F4",X"64",X"E3",X"9F",X"1A",X"F4",X"64",X"E1",X"78",
		X"FE",X"00",X"28",X"F3",X"3A",X"F4",X"64",X"E3",X"DF",X"1A",X"F4",X"64",X"30",X"E7",X"78",X"FE",
		X"00",X"28",X"F5",X"3A",X"F4",X"64",X"E3",X"DF",X"1A",X"F4",X"64",X"30",X"D1",X"09",X"F5",X"64",
		X"E3",X"76",X"28",X"2C",X"E3",X"B6",X"09",X"40",X"40",X"E5",X"52",X"10",X"FE",X"B3",X"08",X"24",
		X"09",X"40",X"44",X"E5",X"52",X"10",X"FE",X"B5",X"08",X"02",X"30",X"14",X"AF",X"1A",X"C9",X"64",
		X"30",X"26",X"AF",X"11",X"80",X"03",X"86",X"0B",X"33",X"47",X"7A",X"9B",X"78",X"08",X"DF",X"E1",
		X"00",X"3E",X"40",X"E5",X"AD",X"14",X"3E",X"21",X"E5",X"BD",X"14",X"11",X"29",X"45",X"09",X"B7",
		X"10",X"3E",X"15",X"06",X"23",X"E5",X"B3",X"15",X"11",X"45",X"41",X"09",X"2C",X"36",X"3E",X"01",
		X"06",X"24",X"E5",X"85",X"15",X"09",X"FD",X"09",X"11",X"E2",X"42",X"01",X"FF",X"21",X"ED",X"88",
		X"13",X"10",X"FB",X"AF",X"12",X"E5",X"9A",X"15",X"3E",X"01",X"12",X"E5",X"88",X"10",X"E1",X"03",
		X"09",X"DF",X"64",X"11",X"6A",X"42",X"E5",X"C8",X"10",X"11",X"6C",X"42",X"E5",X"C8",X"10",X"11",
		X"6E",X"42",X"E5",X"C8",X"10",X"11",X"58",X"42",X"E5",X"C8",X"10",X"11",X"5A",X"42",X"E5",X"C8",
		X"10",X"11",X"5C",X"42",X"E5",X"C8",X"10",X"11",X"5E",X"42",X"E5",X"C8",X"10",X"11",X"78",X"42",
		X"E5",X"C8",X"10",X"11",X"7A",X"42",X"E5",X"C8",X"10",X"11",X"7C",X"42",X"E5",X"C8",X"10",X"E1",
		X"06",X"03",X"26",X"27",X"3E",X"09",X"ED",X"88",X"E5",X"79",X"15",X"10",X"DF",X"0B",X"0B",X"3E",
		X"40",X"E5",X"79",X"15",X"E5",X"FD",X"10",X"3E",X"04",X"E5",X"48",X"15",X"E1",X"3E",X"03",X"DD",
		X"7E",X"CE",X"D8",X"E3",X"3F",X"E3",X"3F",X"E3",X"3F",X"E3",X"3F",X"47",X"3A",X"F4",X"64",X"E3",
		X"5F",X"28",X"2A",X"78",X"12",X"3E",X"08",X"E5",X"79",X"15",X"7E",X"CE",X"27",X"47",X"3A",X"F4",
		X"64",X"E3",X"5F",X"1A",X"F4",X"64",X"28",X"0C",X"78",X"12",X"2B",X"3E",X"08",X"E5",X"79",X"15",
		X"D9",X"3D",X"08",X"E3",X"3A",X"F4",X"64",X"E3",X"9F",X"1A",X"F4",X"64",X"E1",X"78",X"FE",X"00",
		X"28",X"D3",X"3A",X"F4",X"64",X"E3",X"DF",X"1A",X"F4",X"64",X"30",X"C7",X"78",X"FE",X"00",X"28",
		X"F1",X"3A",X"F4",X"64",X"E3",X"DF",X"1A",X"F4",X"64",X"30",X"E5",X"06",X"03",X"32",X"BE",X"38",
		X"20",X"08",X"26",X"2B",X"33",X"10",X"DE",X"30",X"06",X"E5",X"5E",X"11",X"1F",X"3F",X"E1",X"1F",
		X"E1",X"E5",X"5E",X"11",X"1F",X"E1",X"78",X"FE",X"00",X"E0",X"2B",X"33",X"3D",X"08",X"FB",X"E1",
		X"5C",X"45",X"47",X"47",X"67",X"52",X"2C",X"43",X"67",X"50",X"71",X"52",X"61",X"47",X"60",X"54",
		X"08",X"19",X"39",X"38",X"1B",X"54",X"45",X"64",X"63",X"67",X"08",X"61",X"66",X"43",X"09",X"F4",
		X"64",X"E3",X"EE",X"09",X"EE",X"64",X"11",X"39",X"65",X"01",X"03",X"00",X"ED",X"98",X"E5",X"E0",
		X"11",X"09",X"F4",X"64",X"E3",X"4E",X"C0",X"E3",X"AE",X"09",X"D9",X"64",X"11",X"39",X"65",X"01",
		X"03",X"00",X"ED",X"98",X"E5",X"E0",X"11",X"E1",X"01",X"00",X"22",X"09",X"1D",X"65",X"11",X"3B",
		X"65",X"2B",X"2B",X"2B",X"C5",X"E5",X"73",X"11",X"C1",X"18",X"22",X"3E",X"06",X"81",X"67",X"10",
		X"ED",X"2B",X"2B",X"30",X"20",X"79",X"FE",X"00",X"E0",X"0B",X"0B",X"0B",X"0B",X"C5",X"CD",X"06",
		X"00",X"09",X"1A",X"65",X"11",X"38",X"65",X"ED",X"B8",X"3E",X"40",X"E5",X"AD",X"14",X"09",X"F4",
		X"64",X"E3",X"6E",X"08",X"33",X"11",X"4A",X"41",X"09",X"DC",X"35",X"3E",X"01",X"06",X"22",X"E5",
		X"85",X"15",X"09",X"F4",X"64",X"E3",X"7E",X"28",X"31",X"3E",X"01",X"1A",X"03",X"50",X"30",X"12",
		X"11",X"4A",X"41",X"09",X"CF",X"35",X"3E",X"01",X"06",X"22",X"E5",X"85",X"15",X"3E",X"00",X"1A",
		X"03",X"50",X"11",X"40",X"44",X"09",X"A3",X"14",X"3E",X"23",X"06",X"34",X"E5",X"B3",X"15",X"11",
		X"64",X"44",X"09",X"A4",X"14",X"3E",X"03",X"06",X"34",X"E5",X"B3",X"15",X"11",X"51",X"44",X"09",
		X"A5",X"14",X"3E",X"10",X"06",X"34",X"E5",X"B3",X"15",X"11",X"50",X"44",X"09",X"A6",X"14",X"3E",
		X"02",X"06",X"34",X"E5",X"B3",X"15",X"D1",X"D5",X"3E",X"40",X"D5",X"C9",X"13",X"01",X"03",X"00",
		X"5F",X"ED",X"98",X"1E",X"00",X"01",X"02",X"00",X"ED",X"98",X"D1",X"C1",X"D5",X"78",X"09",X"7A",
		X"0A",X"E3",X"0F",X"E5",X"48",X"15",X"66",X"0B",X"46",X"C5",X"09",X"80",X"04",X"21",X"26",X"01",
		X"06",X"27",X"59",X"3E",X"08",X"E5",X"6F",X"15",X"10",X"F8",X"11",X"C3",X"40",X"09",X"38",X"36",
		X"3E",X"01",X"06",X"14",X"E5",X"85",X"15",X"11",X"8D",X"41",X"09",X"64",X"36",X"3E",X"01",X"06",
		X"07",X"E5",X"85",X"15",X"11",X"8F",X"40",X"09",X"53",X"36",X"3E",X"01",X"06",X"16",X"E5",X"85",
		X"15",X"11",X"A8",X"40",X"09",X"69",X"36",X"3E",X"01",X"06",X"16",X"E5",X"85",X"15",X"11",X"69",
		X"42",X"09",X"7F",X"36",X"3E",X"01",X"06",X"20",X"E5",X"85",X"15",X"11",X"64",X"40",X"09",X"87",
		X"36",X"3E",X"03",X"06",X"01",X"E5",X"85",X"15",X"11",X"A5",X"40",X"09",X"08",X"0A",X"3E",X"01",
		X"06",X"32",X"E5",X"85",X"15",X"3E",X"01",X"11",X"AD",X"47",X"12",X"AF",X"1A",X"3D",X"65",X"1A",
		X"3E",X"65",X"09",X"AD",X"47",X"0A",X"3F",X"65",X"11",X"59",X"41",X"09",X"2C",X"36",X"3E",X"01",
		X"06",X"24",X"E5",X"85",X"15",X"09",X"FD",X"09",X"11",X"DC",X"42",X"01",X"21",X"00",X"ED",X"98",
		X"AF",X"12",X"E5",X"9A",X"15",X"3E",X"01",X"12",X"09",X"DF",X"64",X"11",X"94",X"42",X"E5",X"C8",
		X"10",X"11",X"95",X"42",X"E5",X"C8",X"10",X"11",X"96",X"42",X"E5",X"C8",X"10",X"11",X"97",X"42",
		X"E5",X"C8",X"10",X"11",X"B0",X"42",X"E5",X"C8",X"10",X"11",X"B1",X"42",X"E5",X"C8",X"10",X"11",
		X"B2",X"42",X"E5",X"C8",X"10",X"11",X"B3",X"42",X"E5",X"C8",X"10",X"11",X"B4",X"42",X"E5",X"C8",
		X"10",X"11",X"B5",X"42",X"E5",X"C8",X"10",X"3A",X"3C",X"65",X"E3",X"67",X"E2",X"DB",X"13",X"E3",
		X"57",X"E2",X"2B",X"14",X"3A",X"3C",X"65",X"E3",X"4F",X"C2",X"6C",X"14",X"3A",X"3D",X"65",X"FE",
		X"33",X"28",X"37",X"09",X"06",X"0A",X"E5",X"48",X"15",X"7E",X"C9",X"D1",X"12",X"13",X"5F",X"3E",
		X"08",X"E5",X"6F",X"15",X"D5",X"CD",X"3A",X"3E",X"65",X"3C",X"1A",X"3E",X"65",X"FE",X"03",X"C2",
		X"7F",X"14",X"09",X"A6",X"0A",X"3A",X"3E",X"65",X"E5",X"48",X"15",X"7E",X"C9",X"D1",X"CD",X"E5",
		X"4D",X"15",X"09",X"39",X"65",X"01",X"03",X"00",X"ED",X"98",X"3A",X"3E",X"65",X"FE",X"00",X"28",
		X"0D",X"09",X"92",X"0A",X"E5",X"48",X"15",X"7E",X"D1",X"E5",X"79",X"15",X"09",X"3B",X"65",X"E5",
		X"FD",X"10",X"09",X"FC",X"64",X"11",X"DA",X"43",X"E5",X"D7",X"27",X"09",X"F5",X"64",X"E3",X"86",
		X"3E",X"01",X"E5",X"FF",X"14",X"E1",X"D1",X"3E",X"80",X"E5",X"79",X"15",X"3E",X"08",X"E5",X"79",
		X"15",X"30",X"F1",X"3A",X"3D",X"65",X"FE",X"00",X"E2",X"5C",X"13",X"3D",X"1A",X"3D",X"65",X"FE",
		X"32",X"28",X"14",X"3E",X"05",X"2A",X"3F",X"65",X"5F",X"3E",X"08",X"E5",X"48",X"15",X"0A",X"3F",
		X"65",X"3E",X"01",X"5F",X"C3",X"5C",X"13",X"3D",X"1A",X"3D",X"65",X"3E",X"05",X"2A",X"3F",X"65",
		X"2B",X"5F",X"0B",X"5F",X"0B",X"5F",X"2B",X"3E",X"40",X"30",X"C8",X"3A",X"3D",X"65",X"FE",X"33",
		X"E2",X"5C",X"13",X"3C",X"1A",X"3D",X"65",X"FE",X"32",X"28",X"14",X"3E",X"05",X"2A",X"3F",X"65",
		X"5F",X"3E",X"08",X"E5",X"6F",X"15",X"0A",X"3F",X"65",X"3E",X"01",X"5F",X"C3",X"5C",X"13",X"3C",
		X"1A",X"3D",X"65",X"3E",X"05",X"2A",X"3F",X"65",X"5F",X"3E",X"40",X"E5",X"6F",X"15",X"0A",X"3F",
		X"65",X"3E",X"01",X"2B",X"5F",X"0B",X"5F",X"0B",X"5F",X"C3",X"5C",X"13",X"3E",X"20",X"E5",X"63",
		X"15",X"1A",X"C0",X"50",X"06",X"14",X"E5",X"17",X"15",X"F2",X"8A",X"13",X"C3",X"4F",X"13",X"3A",
		X"3C",X"65",X"E3",X"4F",X"1A",X"C0",X"50",X"28",X"DE",X"30",X"CE",X"21",X"05",X"10",X"01",X"D5",
		X"AF",X"E3",X"0B",X"17",X"E3",X"0B",X"17",X"E3",X"0B",X"17",X"E3",X"0B",X"17",X"E3",X"0B",X"17",
		X"57",X"EB",X"01",X"40",X"40",X"21",X"06",X"00",X"D1",X"62",X"21",X"EB",X"E1",X"09",X"40",X"40",
		X"11",X"41",X"40",X"01",X"7F",X"03",X"5F",X"ED",X"98",X"1A",X"C0",X"50",X"E1",X"09",X"40",X"44",
		X"11",X"41",X"44",X"01",X"7F",X"03",X"5F",X"ED",X"98",X"1A",X"C0",X"50",X"E1",X"3A",X"C9",X"64",
		X"FE",X"00",X"E0",X"3A",X"CB",X"64",X"CE",X"D8",X"E3",X"3F",X"E3",X"3F",X"E3",X"3F",X"E3",X"3F",
		X"FE",X"00",X"28",X"24",X"1A",X"25",X"40",X"3A",X"CB",X"64",X"CE",X"27",X"1A",X"24",X"40",X"E1",
		X"3E",X"40",X"30",X"D8",X"3E",X"21",X"E5",X"BD",X"14",X"3E",X"40",X"E5",X"AD",X"14",X"E1",X"47",
		X"AF",X"1A",X"CC",X"64",X"1A",X"CE",X"64",X"3A",X"CE",X"64",X"B8",X"E0",X"09",X"F3",X"64",X"E3",
		X"6E",X"C0",X"1A",X"C0",X"50",X"30",X"D8",X"3A",X"F5",X"64",X"E3",X"47",X"28",X"25",X"3A",X"CF",
		X"64",X"47",X"3A",X"CE",X"64",X"B8",X"18",X"31",X"1F",X"3F",X"E1",X"78",X"1A",X"CF",X"64",X"3A",
		X"F5",X"64",X"E3",X"C7",X"1A",X"F5",X"64",X"AF",X"1A",X"CE",X"64",X"1A",X"CC",X"64",X"1F",X"3F",
		X"E1",X"3A",X"F5",X"64",X"E3",X"87",X"1A",X"F5",X"64",X"1F",X"E1",X"47",X"AF",X"1A",X"CD",X"64",
		X"3A",X"CD",X"64",X"B8",X"E0",X"09",X"F3",X"64",X"E3",X"6E",X"C0",X"1A",X"C0",X"50",X"30",X"D8",
		X"85",X"6F",X"D0",X"0C",X"E1",X"83",X"77",X"D0",X"14",X"E1",X"81",X"67",X"D0",X"04",X"E1",X"D5",
		X"16",X"00",X"77",X"1F",X"3F",X"ED",X"52",X"D1",X"E1",X"CD",X"EB",X"16",X"00",X"77",X"1F",X"3F",
		X"ED",X"52",X"EB",X"C9",X"E1",X"1A",X"8E",X"64",X"D5",X"3A",X"8E",X"64",X"67",X"ED",X"88",X"79",
		X"FE",X"00",X"08",X"F9",X"D1",X"E5",X"9A",X"15",X"10",X"EE",X"E1",X"1A",X"8E",X"64",X"D5",X"3A",
		X"8E",X"64",X"67",X"ED",X"88",X"2B",X"79",X"FE",X"00",X"08",X"F8",X"D1",X"E5",X"9A",X"15",X"10",
		X"ED",X"E1",X"CD",X"09",X"08",X"00",X"31",X"EB",X"C9",X"E1",X"09",X"8F",X"64",X"06",X"2F",X"1E",
		X"00",X"0B",X"10",X"FB",X"E1",X"09",X"F3",X"64",X"E3",X"FE",X"E3",X"7E",X"E0",X"1A",X"C0",X"50",
		X"30",X"F8",X"3A",X"00",X"50",X"CE",X"27",X"47",X"3A",X"40",X"50",X"CE",X"D8",X"98",X"1A",X"3C",
		X"65",X"E1",X"3A",X"40",X"50",X"47",X"CE",X"27",X"E3",X"78",X"28",X"02",X"E3",X"CF",X"1A",X"3C",
		X"65",X"E1",X"F5",X"09",X"42",X"65",X"F5",X"E3",X"00",X"46",X"C4",X"0B",X"17",X"F5",X"E3",X"00",
		X"56",X"28",X"10",X"E5",X"2B",X"17",X"FD",X"09",X"51",X"50",X"E5",X"FA",X"16",X"F5",X"7E",X"06",
		X"1A",X"45",X"50",X"F5",X"09",X"75",X"65",X"F5",X"E3",X"00",X"46",X"C4",X"0B",X"17",X"F5",X"E3",
		X"00",X"56",X"28",X"10",X"E5",X"2B",X"17",X"FD",X"09",X"51",X"50",X"E5",X"FA",X"16",X"F5",X"7E",
		X"06",X"1A",X"45",X"50",X"F5",X"09",X"78",X"65",X"F5",X"E3",X"00",X"46",X"C4",X"0B",X"17",X"F5",
		X"E3",X"00",X"56",X"28",X"10",X"E5",X"2B",X"17",X"FD",X"09",X"51",X"50",X"E5",X"FA",X"16",X"F5",
		X"7E",X"06",X"1A",X"45",X"50",X"F5",X"09",X"93",X"65",X"F5",X"E3",X"00",X"46",X"C4",X"0B",X"17",
		X"F5",X"E3",X"00",X"56",X"28",X"10",X"E5",X"2B",X"17",X"FD",X"09",X"56",X"50",X"E5",X"FA",X"16",
		X"F5",X"7E",X"06",X"1A",X"62",X"50",X"F5",X"09",X"AE",X"65",X"F5",X"E3",X"00",X"46",X"C4",X"0B",
		X"17",X"F5",X"E3",X"00",X"56",X"28",X"10",X"E5",X"2B",X"17",X"FD",X"09",X"56",X"50",X"E5",X"FA",
		X"16",X"F5",X"7E",X"06",X"1A",X"62",X"50",X"F5",X"09",X"E1",X"65",X"F5",X"E3",X"00",X"46",X"C4",
		X"0B",X"17",X"F5",X"E3",X"00",X"56",X"28",X"10",X"E5",X"2B",X"17",X"FD",X"09",X"56",X"50",X"E5",
		X"FA",X"16",X"F5",X"7E",X"06",X"1A",X"62",X"50",X"F5",X"09",X"CC",X"65",X"F5",X"E3",X"00",X"46",
		X"C4",X"0B",X"17",X"F5",X"E3",X"00",X"56",X"28",X"10",X"E5",X"2B",X"17",X"FD",X"09",X"73",X"50",
		X"E5",X"FA",X"16",X"F5",X"7E",X"06",X"1A",X"67",X"50",X"F5",X"09",X"FF",X"65",X"F5",X"E3",X"00",
		X"46",X"C4",X"0B",X"17",X"F5",X"E3",X"00",X"56",X"E0",X"E5",X"2B",X"17",X"FD",X"09",X"73",X"50",
		X"E5",X"FA",X"16",X"F5",X"7E",X"06",X"1A",X"67",X"50",X"E1",X"F5",X"7E",X"03",X"FD",X"5F",X"00",
		X"E3",X"3F",X"E3",X"3F",X"E3",X"3F",X"E3",X"3F",X"FD",X"5F",X"01",X"F5",X"7E",X"04",X"FD",X"5F",
		X"02",X"E3",X"3F",X"E3",X"3F",X"E3",X"3F",X"E3",X"3F",X"FD",X"5F",X"03",X"F5",X"7E",X"05",X"FD",
		X"5F",X"04",X"E1",X"E5",X"FF",X"17",X"F5",X"E3",X"00",X"D6",X"E1",X"F5",X"E3",X"00",X"66",X"C2",
		X"FF",X"17",X"F5",X"6E",X"01",X"F5",X"4E",X"02",X"7E",X"E3",X"0F",X"11",X"61",X"17",X"E5",X"4D",
		X"15",X"0B",X"CD",X"32",X"6F",X"13",X"32",X"4F",X"E9",X"4B",X"17",X"4F",X"17",X"5D",X"17",X"7E",
		X"17",X"94",X"17",X"89",X"17",X"BB",X"17",X"D4",X"17",X"DE",X"17",X"FE",X"17",X"35",X"30",X"29",
		X"30",X"1D",X"30",X"C9",X"C3",X"38",X"17",X"C9",X"7E",X"F5",X"5F",X"03",X"0B",X"7E",X"0B",X"F5",
		X"5F",X"04",X"C3",X"38",X"17",X"C9",X"7E",X"F5",X"5F",X"05",X"0B",X"C3",X"38",X"17",X"C9",X"7E",
		X"F5",X"46",X"03",X"80",X"F5",X"5F",X"03",X"0B",X"7E",X"0B",X"F5",X"46",X"04",X"A0",X"F5",X"5F",
		X"04",X"C3",X"38",X"17",X"C9",X"7E",X"F5",X"46",X"05",X"80",X"F5",X"5F",X"05",X"0B",X"C3",X"38",
		X"17",X"C9",X"7E",X"F5",X"BE",X"07",X"28",X"23",X"F5",X"1C",X"07",X"2B",X"F5",X"5D",X"01",X"F5",
		X"5C",X"02",X"E1",X"F5",X"1E",X"07",X"00",X"0B",X"C3",X"38",X"17",X"F5",X"6E",X"20",X"F5",X"4E",
		X"21",X"D1",X"D5",X"2B",X"5A",X"2B",X"5B",X"2B",X"1E",X"00",X"F5",X"5D",X"20",X"F5",X"5C",X"21",
		X"C9",X"C3",X"38",X"17",X"D1",X"32",X"F5",X"6E",X"20",X"F5",X"4E",X"21",X"BE",X"28",X"21",X"1C",
		X"0B",X"76",X"0B",X"56",X"EB",X"C3",X"38",X"17",X"0B",X"0B",X"0B",X"F5",X"5D",X"20",X"F5",X"5C",
		X"21",X"13",X"EB",X"C3",X"38",X"17",X"C9",X"76",X"0B",X"56",X"EB",X"C3",X"38",X"17",X"C9",X"F5",
		X"CD",X"F5",X"CD",X"C9",X"D1",X"13",X"1E",X"00",X"01",X"30",X"00",X"ED",X"98",X"32",X"F5",X"5F",
		X"01",X"13",X"32",X"F5",X"5F",X"02",X"F5",X"5D",X"20",X"F5",X"5C",X"21",X"E1",X"C9",X"F5",X"5D",
		X"01",X"F5",X"5C",X"02",X"F5",X"1E",X"00",X"00",X"E1",X"C9",X"76",X"0B",X"56",X"EB",X"1E",X"06",
		X"13",X"EB",X"C3",X"38",X"17",X"C9",X"7E",X"F5",X"5F",X"06",X"0B",X"C3",X"38",X"17",X"23",X"75",
		X"65",X"23",X"78",X"65",X"24",X"02",X"01",X"43",X"00",X"02",X"20",X"05",X"04",X"01",X"54",X"00",
		X"05",X"04",X"01",X"1A",X"00",X"05",X"04",X"01",X"85",X"00",X"05",X"04",X"01",X"8F",X"00",X"05",
		X"04",X"01",X"4C",X"00",X"05",X"04",X"01",X"23",X"01",X"05",X"04",X"21",X"00",X"E2",X"7B",X"30",
		X"23",X"42",X"65",X"23",X"78",X"65",X"01",X"D8",X"00",X"24",X"02",X"06",X"02",X"20",X"05",X"03",
		X"02",X"00",X"05",X"03",X"07",X"20",X"21",X"E5",X"0B",X"14",X"E5",X"DD",X"23",X"44",X"65",X"E5",
		X"94",X"15",X"26",X"29",X"E5",X"0B",X"14",X"C3",X"F2",X"30",X"E5",X"E6",X"23",X"CE",X"40",X"FE",
		X"00",X"C2",X"23",X"42",X"65",X"23",X"75",X"65",X"24",X"02",X"02",X"22",X"06",X"01",X"80",X"00",
		X"06",X"03",X"18",X"00",X"05",X"01",X"07",X"20",X"04",X"FE",X"07",X"04",X"21",X"07",X"01",X"56",
		X"13",X"E5",X"99",X"15",X"C3",X"F2",X"30",X"26",X"28",X"E5",X"0B",X"14",X"E5",X"DD",X"23",X"0B",
		X"44",X"65",X"E5",X"94",X"23",X"AE",X"65",X"06",X"24",X"04",X"06",X"01",X"90",X"00",X"06",X"03",
		X"20",X"00",X"04",X"05",X"05",X"02",X"07",X"02",X"02",X"00",X"07",X"02",X"24",X"03",X"02",X"06",
		X"06",X"03",X"20",X"00",X"04",X"05",X"05",X"02",X"07",X"02",X"05",X"07",X"02",X"00",X"07",X"02",
		X"21",X"36",X"9D",X"E2",X"21",X"31",X"23",X"93",X"65",X"24",X"06",X"01",X"80",X"00",X"02",X"27",
		X"06",X"03",X"08",X"00",X"05",X"02",X"07",X"20",X"21",X"4B",X"31",X"2A",X"25",X"00",X"EB",X"2A",
		X"A4",X"20",X"31",X"0A",X"BA",X"23",X"2A",X"BA",X"23",X"76",X"0B",X"56",X"EB",X"0A",X"A4",X"20",
		X"E5",X"D6",X"23",X"D6",X"01",X"C6",X"FF",X"B7",X"23",X"93",X"65",X"23",X"AE",X"65",X"23",X"CC",
		X"65",X"24",X"02",X"02",X"27",X"06",X"01",X"00",X"01",X"06",X"03",X"30",X"00",X"05",X"01",X"07",
		X"24",X"05",X"02",X"04",X"FF",X"07",X"26",X"21",X"29",X"21",X"66",X"0B",X"46",X"E5",X"DB",X"14",
		X"C3",X"27",X"31",X"2A",X"4A",X"07",X"0A",X"91",X"20",X"3E",X"24",X"02",X"01",X"00",X"D8",X"02",
		X"07",X"06",X"03",X"68",X"00",X"05",X"01",X"07",X"20",X"03",X"00",X"07",X"20",X"59",X"31",X"23",
		X"2A",X"BA",X"23",X"76",X"0B",X"56",X"EB",X"0A",X"91",X"20",X"E5",X"D6",X"23",X"6F",X"0E",X"00",
		X"0A",X"A6",X"20",X"2A",X"A6",X"20",X"01",X"48",X"05",X"29",X"21",X"66",X"23",X"CC",X"65",X"24",
		X"02",X"01",X"95",X"00",X"02",X"26",X"06",X"04",X"FE",X"05",X"02",X"07",X"04",X"01",X"C7",X"00",
		X"02",X"26",X"06",X"04",X"FE",X"05",X"02",X"07",X"04",X"01",X"C7",X"00",X"02",X"26",X"06",X"04",
		X"FE",X"05",X"02",X"07",X"04",X"01",X"FA",X"00",X"02",X"26",X"06",X"04",X"FE",X"05",X"02",X"07",
		X"02",X"01",X"C7",X"00",X"02",X"26",X"06",X"04",X"FE",X"05",X"02",X"07",X"02",X"01",X"FA",X"00",
		X"02",X"26",X"06",X"04",X"FE",X"05",X"02",X"07",X"02",X"01",X"2A",X"01",X"02",X"26",X"06",X"04",
		X"FE",X"05",X"02",X"07",X"06",X"01",X"FA",X"00",X"02",X"26",X"06",X"04",X"FE",X"05",X"02",X"07",
		X"04",X"01",X"C7",X"00",X"02",X"26",X"06",X"04",X"FE",X"05",X"02",X"07",X"04",X"01",X"95",X"00",
		X"02",X"26",X"06",X"04",X"FE",X"05",X"02",X"07",X"02",X"01",X"95",X"00",X"02",X"26",X"06",X"04",
		X"FE",X"05",X"02",X"07",X"02",X"01",X"C7",X"00",X"02",X"26",X"06",X"04",X"FE",X"05",X"02",X"07",
		X"04",X"01",X"C7",X"00",X"02",X"26",X"06",X"04",X"FE",X"05",X"02",X"07",X"04",X"01",X"FA",X"00",
		X"02",X"26",X"06",X"04",X"FE",X"05",X"02",X"07",X"02",X"01",X"C7",X"00",X"02",X"26",X"06",X"04",
		X"FE",X"05",X"02",X"07",X"02",X"01",X"FA",X"00",X"02",X"26",X"06",X"04",X"FE",X"05",X"02",X"07",
		X"04",X"01",X"C8",X"00",X"02",X"26",X"06",X"04",X"FE",X"05",X"02",X"07",X"20",X"05",X"20",X"01",
		X"95",X"00",X"02",X"26",X"06",X"04",X"FE",X"05",X"02",X"07",X"02",X"01",X"95",X"00",X"02",X"26",
		X"06",X"04",X"FE",X"05",X"02",X"07",X"02",X"01",X"C7",X"00",X"02",X"26",X"06",X"04",X"FE",X"05",
		X"02",X"07",X"04",X"01",X"C7",X"00",X"02",X"26",X"06",X"04",X"FE",X"05",X"02",X"07",X"04",X"01",
		X"FA",X"00",X"02",X"26",X"06",X"04",X"FE",X"05",X"02",X"07",X"02",X"01",X"C7",X"00",X"02",X"26",
		X"06",X"04",X"FE",X"05",X"02",X"07",X"02",X"01",X"FA",X"00",X"02",X"26",X"06",X"04",X"FE",X"05",
		X"02",X"07",X"02",X"01",X"2A",X"01",X"02",X"26",X"06",X"04",X"FE",X"05",X"02",X"07",X"06",X"01",
		X"FA",X"00",X"02",X"26",X"06",X"04",X"FE",X"05",X"02",X"07",X"04",X"01",X"C7",X"00",X"02",X"26",
		X"06",X"04",X"FE",X"05",X"02",X"07",X"04",X"01",X"95",X"00",X"02",X"26",X"06",X"04",X"FE",X"05",
		X"02",X"07",X"02",X"01",X"95",X"00",X"02",X"26",X"06",X"04",X"FE",X"05",X"02",X"07",X"02",X"01",
		X"95",X"00",X"02",X"26",X"06",X"04",X"FE",X"05",X"02",X"07",X"04",X"01",X"95",X"00",X"02",X"26",
		X"06",X"04",X"FE",X"05",X"02",X"07",X"04",X"01",X"95",X"00",X"02",X"26",X"06",X"04",X"FE",X"05",
		X"02",X"07",X"04",X"01",X"8F",X"00",X"02",X"26",X"06",X"04",X"FE",X"05",X"02",X"07",X"02",X"01",
		X"BC",X"00",X"02",X"26",X"06",X"04",X"FE",X"05",X"02",X"07",X"02",X"01",X"C7",X"00",X"02",X"26",
		X"06",X"04",X"FE",X"05",X"02",X"07",X"06",X"21",X"67",X"33",X"09",X"B5",X"07",X"1E",X"00",X"3A",
		X"41",X"04",X"FE",X"1A",X"F2",X"75",X"33",X"E5",X"16",X"27",X"C3",X"4E",X"33",X"E5",X"F6",X"15",
		X"E5",X"F6",X"15",X"E5",X"F6",X"15",X"01",X"4E",X"07",X"E5",X"03",X"27",X"01",X"4E",X"07",X"E5",
		X"23",X"21",X"3E",X"00",X"11",X"23",X"00",X"E5",X"18",X"36",X"9D",X"C2",X"90",X"33",X"E5",X"F6",
		X"15",X"01",X"D6",X"07",X"E5",X"03",X"27",X"01",X"D6",X"07",X"E5",X"23",X"21",X"C3",X"CB",X"33",
		X"E5",X"F6",X"15",X"2A",X"23",X"00",X"44",X"65",X"11",X"A9",X"07",X"E5",X"FF",X"25",X"3E",X"01",
		X"11",X"23",X"00",X"E5",X"18",X"36",X"9D",X"C2",X"AF",X"33",X"09",X"9C",X"07",X"1E",X"08",X"3E",
		X"00",X"11",X"D4",X"04",X"E5",X"18",X"36",X"9D",X"E2",X"C6",X"33",X"2A",X"D4",X"04",X"44",X"65",
		X"11",X"BE",X"07",X"E5",X"FF",X"25",X"3E",X"01",X"11",X"D4",X"04",X"E5",X"18",X"36",X"9D",X"C2",
		X"D7",X"33",X"09",X"D4",X"07",X"1E",X"08",X"01",X"A9",X"07",X"E5",X"03",X"27",X"01",X"A9",X"07",
		X"E5",X"23",X"21",X"E1",X"09",X"94",X"20",X"58",X"2B",X"59",X"3E",X"FF",X"37",X"D2",X"7E",X"34",
		X"2A",X"93",X"20",X"3E",X"00",X"E5",X"3B",X"36",X"9D",X"C2",X"17",X"34",X"01",X"25",X"00",X"11",
		X"BA",X"23",X"E5",X"0B",X"36",X"CD",X"2A",X"93",X"20",X"C1",X"59",X"0B",X"58",X"2A",X"BA",X"23",
		X"3E",X"00",X"5F",X"0B",X"1E",X"00",X"E1",X"2A",X"93",X"20",X"11",X"25",X"00",X"E5",X"AC",X"35",
		X"2B",X"CD",X"E5",X"D8",X"23",X"44",X"65",X"36",X"00",X"E5",X"CE",X"22",X"67",X"06",X"00",X"09",
		X"5D",X"34",X"21",X"21",X"76",X"0B",X"56",X"EB",X"E9",X"2A",X"93",X"20",X"11",X"25",X"00",X"E5",
		X"AC",X"35",X"0A",X"93",X"20",X"C3",X"7B",X"34",X"01",X"5F",X"13",X"E5",X"23",X"21",X"C3",X"7B",
		X"34",X"2A",X"93",X"20",X"CD",X"2A",X"BA",X"23",X"CB",X"66",X"0B",X"46",X"C9",X"59",X"0B",X"58",
		X"01",X"25",X"00",X"11",X"BA",X"23",X"E5",X"0B",X"36",X"CD",X"2A",X"93",X"20",X"C1",X"59",X"0B",
		X"58",X"E1",X"C3",X"7B",X"34",X"39",X"34",X"60",X"34",X"51",X"34",X"C3",X"EA",X"33",X"E1",X"2A",
		X"25",X"00",X"0B",X"0B",X"76",X"0B",X"56",X"EB",X"0A",X"76",X"05",X"09",X"95",X"20",X"1E",X"00",
		X"3E",X"27",X"09",X"95",X"20",X"BE",X"F2",X"FE",X"34",X"2A",X"95",X"20",X"0E",X"00",X"01",X"02",
		X"00",X"29",X"21",X"EB",X"2A",X"25",X"00",X"31",X"11",X"25",X"00",X"E5",X"AC",X"35",X"0A",X"BA",
		X"23",X"09",X"01",X"00",X"0A",X"96",X"20",X"2A",X"BA",X"23",X"3E",X"00",X"E5",X"3B",X"36",X"9D",
		X"E2",X"F1",X"34",X"2A",X"BA",X"23",X"11",X"25",X"00",X"E5",X"AC",X"35",X"0A",X"BA",X"23",X"2A",
		X"96",X"20",X"0B",X"0A",X"96",X"20",X"C3",X"9F",X"34",X"2A",X"95",X"20",X"0E",X"00",X"01",X"04",
		X"00",X"29",X"21",X"EB",X"2A",X"25",X"00",X"31",X"CD",X"2A",X"BA",X"23",X"CB",X"66",X"0B",X"46",
		X"C9",X"59",X"0B",X"58",X"3A",X"95",X"20",X"3C",X"1A",X"95",X"20",X"C2",X"90",X"34",X"2A",X"BA",
		X"23",X"3E",X"00",X"5F",X"0B",X"1E",X"00",X"3E",X"00",X"11",X"76",X"05",X"E5",X"18",X"36",X"9D",
		X"E2",X"A9",X"35",X"2A",X"25",X"00",X"EB",X"2A",X"76",X"05",X"31",X"0A",X"BA",X"23",X"2A",X"BA",
		X"23",X"76",X"0B",X"56",X"EB",X"0A",X"76",X"05",X"E5",X"E2",X"23",X"D6",X"05",X"D6",X"01",X"B7",
		X"DD",X"E5",X"E2",X"23",X"D6",X"06",X"D6",X"01",X"B7",X"C1",X"60",X"99",X"37",X"D2",X"61",X"35",
		X"01",X"48",X"07",X"E5",X"CC",X"33",X"C3",X"8E",X"35",X"E5",X"E2",X"23",X"D6",X"01",X"D6",X"01",
		X"B7",X"DD",X"E5",X"E2",X"23",X"D6",X"07",X"D6",X"01",X"B7",X"C1",X"60",X"99",X"37",X"D2",X"B0",
		X"35",X"E5",X"D2",X"23",X"CE",X"03",X"FE",X"03",X"C2",X"5C",X"35",X"01",X"4A",X"07",X"E5",X"CC",
		X"33",X"C3",X"95",X"35",X"E5",X"D2",X"23",X"CE",X"80",X"FE",X"00",X"E2",X"85",X"35",X"2A",X"D4",
		X"04",X"0B",X"0A",X"D4",X"1A",X"40",X"52",X"45",X"71",X"41",X"64",X"50",X"40",X"45",X"52",X"67",
		X"43",X"53",X"50",X"67",X"54",X"40",X"19",X"40",X"52",X"45",X"71",X"41",X"64",X"50",X"54",X"61",
		X"44",X"45",X"52",X"43",X"71",X"41",X"64",X"50",X"45",X"45",X"52",X"46",X"40",X"66",X"61",X"67",
		X"43",X"40",X"54",X"52",X"45",X"53",X"66",X"61",X"52",X"45",X"71",X"41",X"64",X"50",X"40",X"45",
		X"66",X"67",X"40",X"54",X"43",X"45",X"64",X"45",X"53",X"52",X"67",X"53",X"52",X"45",X"71",X"41",
		X"64",X"50",X"40",X"67",X"57",X"54",X"40",X"52",X"67",X"40",X"45",X"66",X"67",X"40",X"54",X"43",
		X"45",X"64",X"45",X"53",X"50",X"55",X"40",X"45",X"66",X"67",X"40",X"52",X"45",X"71",X"41",X"64",
		X"50",X"50",X"55",X"40",X"67",X"57",X"54",X"40",X"52",X"45",X"71",X"41",X"64",X"50",X"66",X"61",
		X"41",X"47",X"41",X"40",X"52",X"45",X"71",X"41",X"64",X"50",X"40",X"45",X"65",X"41",X"53",X"52",
		X"45",X"56",X"67",X"40",X"45",X"65",X"41",X"47",X"52",X"45",X"56",X"67",X"40",X"45",X"65",X"41",
		X"47",X"40",X"45",X"66",X"67",X"40",X"52",X"45",X"71",X"41",X"64",X"50",X"45",X"65",X"41",X"46",
		X"40",X"46",X"67",X"40",X"64",X"64",X"41",X"60",X"45",X"60",X"54",X"40",X"66",X"61",X"40",X"53",
		X"61",X"40",X"45",X"52",X"67",X"43",X"53",X"40",X"52",X"55",X"67",X"71",X"66",X"45",X"54",X"40",
		X"50",X"67",X"54",X"54",X"43",X"45",X"64",X"45",X"53",X"40",X"67",X"54",X"40",X"63",X"43",X"61",
		X"54",X"53",X"71",X"67",X"62",X"40",X"45",X"53",X"55",X"66",X"67",X"54",X"54",X"55",X"42",X"40",
		X"45",X"52",X"61",X"46",X"40",X"44",X"66",X"41",X"40",X"52",X"45",X"54",X"54",X"45",X"64",X"54",
		X"66",X"61",X"52",X"50",X"40",X"67",X"54",X"45",X"66",X"44",X"65",X"41",X"64",X"53",X"53",X"54",
		X"66",X"45",X"53",X"45",X"52",X"50",X"40",X"72",X"45",X"60",X"43",X"66",X"41",X"53",X"67",X"63",
		X"64",X"45",X"54",X"40",X"1B",X"38",X"39",X"19",X"2F",X"E0",X"40",X"40",X"40",X"40",X"40",X"40",
		X"40",X"C6",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"C7",X"E1",X"40",X"40",X"40",X"40",X"40",
		X"40",X"C7",X"C6",X"C6",X"C6",X"C6",X"C6",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",
		X"40",X"E0",X"C6",X"C6",X"C6",X"C6",X"E1",X"40",X"40",X"C6",X"40",X"40",X"40",X"40",X"C6",X"40",
		X"40",X"C6",X"40",X"40",X"40",X"40",X"C6",X"40",X"40",X"C7",X"C6",X"C6",X"C6",X"C6",X"E2",X"40",
		X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"E0",X"C6",X"C6",X"C6",X"C6",X"C6",X"C6",
		X"C6",X"C6",X"40",X"40",X"40",X"C6",X"40",X"40",X"C6",X"C6",X"E1",X"40",X"40",X"C6",X"40",X"C7",
		X"E2",X"C7",X"C6",X"C6",X"C6",X"E2",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",
		X"40",X"E0",X"C6",X"C6",X"C6",X"C6",X"C6",X"C6",X"C6",X"C6",X"40",X"40",X"40",X"C6",X"40",X"40",
		X"C6",X"C6",X"E1",X"40",X"40",X"C6",X"40",X"C7",X"E2",X"C7",X"C6",X"C6",X"C6",X"E2",X"40",X"40",
		X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"E0",X"C6",X"E1",X"40",X"E0",X"E1",X"40",
		X"40",X"C6",X"40",X"C6",X"40",X"40",X"C6",X"40",X"40",X"C6",X"40",X"C6",X"40",X"40",X"C6",X"40",
		X"40",X"C7",X"C6",X"C6",X"C6",X"C6",X"E2",X"40",X"40",X"E1",X"40",X"40",X"40",X"40",X"C6",X"40",
		X"40",X"40",X"40",X"C6",X"40",X"E1",X"40",X"40",X"C6",X"40",X"C6",X"40",X"40",X"C7",X"40",X"C6",
		X"40",X"E1",X"40",X"40",X"C6",X"40",X"C6",X"40",X"40",X"C7",X"40",X"C6",X"40",X"40",X"40",X"40",
		X"C6",X"40",X"40",X"40",X"40",X"C7",X"E3",X"E4",X"E5",X"E6",X"E7",X"D0",X"D1",X"D2",X"D3",X"D4",
		X"D5",X"D6",X"D7",X"F0",X"F1",X"F2",X"45",X"64",X"42",X"41",X"54",X"40",X"45",X"43",X"66",X"41",
		X"56",X"44",X"41",X"40",X"45",X"52",X"67",X"43",X"53",X"18",X"18",X"18",X"18",X"18",X"18",X"18",
		X"18",X"18",X"18",X"18",X"18",X"18",X"1D",X"18",X"1D",X"18",X"1D",X"18",X"1D",X"18",X"1D",X"18",
		X"1D",X"18",X"1A",X"1D",X"1F",X"18",X"1A",X"1D",X"1F",X"18",X"1A",X"1D",X"1F",X"19",X"19",X"19",
		X"19",X"1A",X"1A",X"1A",X"1A",X"1B",X"1B",X"1B",X"1B",X"40",X"40",X"40",X"40",X"40",X"40",X"40",
		X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",
		X"40",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",
		X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"19",X"1A",X"1B",X"1C",X"1D",X"1E",X"1F",
		X"38",X"39",X"18",X"19",X"1A",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"19",X"19",
		X"19",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"19",X"1A",X"1B",
		X"1C",X"1D",X"1E",X"1F",X"38",X"39",X"18",X"19",X"1A",X"40",X"40",X"40",X"40",X"40",X"40",X"40",
		X"40",X"40",X"19",X"19",X"19",X"40",X"71",X"41",X"64",X"50",X"40",X"19",X"40",X"53",X"66",X"61",
		X"67",X"43",X"40",X"1A",X"53",X"71",X"41",X"64",X"50",X"40",X"1A",X"40",X"40",X"66",X"61",X"67",
		X"43",X"40",X"19",X"40",X"71",X"41",X"64",X"50",X"40",X"19",X"40",X"40",X"66",X"61",X"67",X"43",
		X"40",X"19",X"53",X"54",X"66",X"61",X"67",X"50",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",
		X"71",X"52",X"45",X"56",X"45",X"40",X"53",X"55",X"66",X"67",X"42",X"18",X"18",X"18",X"1D",X"1A",
		X"19",X"18",X"18",X"18",X"18",X"18",X"19",X"18",X"18",X"18",X"1D",X"1F",X"18",X"18",X"18",X"18",
		X"1D",X"53",X"43",X"61",X"54",X"53",X"67",X"66",X"47",X"41",X"61",X"44",X"66",X"67",X"61",X"54",
		X"61",X"44",X"66",X"67",X"43",X"40",X"40",X"66",X"67",X"61",X"54",X"41",X"43",X"67",X"64",X"40",
		X"40",X"65",X"67",X"52",X"44",X"67",X"67",X"47",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"44",
		X"1F",X"40",X"40",X"40",X"40",X"40",X"40",X"19",X"44",X"67",X"67",X"47",X"40",X"40",X"40",X"40",
		X"40",X"40",X"40",X"46",X"1F",X"40",X"40",X"40",X"40",X"40",X"40",X"1A",X"44",X"67",X"67",X"47",
		X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"60",X"1F",X"40",X"40",X"40",X"40",X"40",X"40",X"1B",
		X"44",X"67",X"67",X"47",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"62",X"1F",X"40",X"40",X"40",
		X"40",X"40",X"40",X"1C",X"44",X"67",X"67",X"47",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"60",
		X"1C",X"40",X"40",X"40",X"40",X"40",X"40",X"19",X"44",X"67",X"67",X"47",X"40",X"40",X"40",X"40",
		X"40",X"40",X"40",X"64",X"1C",X"40",X"40",X"40",X"40",X"40",X"40",X"1A",X"44",X"67",X"67",X"47",
		X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"62",X"1C",X"40",X"40",X"40",X"40",X"40",X"40",X"1B",
		X"44",X"67",X"67",X"47",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"65",X"1C",X"40",X"40",X"40",
		X"40",X"40",X"40",X"1C",X"44",X"67",X"67",X"47",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"63",
		X"1C",X"40",X"40",X"40",X"40",X"40",X"40",X"1D",X"44",X"67",X"67",X"47",X"40",X"40",X"40",X"40",
		X"40",X"40",X"40",X"66",X"1C",X"40",X"40",X"40",X"40",X"40",X"40",X"1E",X"44",X"41",X"42",X"40",
		X"66",X"67",X"61",X"54",X"61",X"44",X"66",X"67",X"43",X"40",X"40",X"66",X"67",X"61",X"54",X"41",
		X"43",X"67",X"64",X"40",X"40",X"65",X"41",X"52",X"00",X"50",X"12",X"00",X"00",X"00",X"0D",X"00",
		X"00",X"50",X"1F",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"08",X"00",
		X"00",X"00",X"18",X"00",X"00",X"00",X"40",X"00",X"00",X"50",X"07",X"00",X"00",X"00",X"15",X"00",
		X"00",X"50",X"0A",X"00",X"00",X"00",X"18",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"10",X"00",
		X"00",X"00",X"15",X"00",X"00",X"00",X"08",X"00",X"05",X"04",X"03",X"02",X"00",X"01",X"02",X"03",
		X"04",X"05",X"06",X"07",X"20",X"21",X"41",X"42",X"43",X"44",X"45",X"46",X"47",X"60",X"61",X"62",
		X"63",X"64",X"65",X"66",X"67",X"50",X"51",X"52",X"53",X"54",X"55",X"56",X"57",X"70",X"71",X"72",
		X"72",X"71",X"70",X"57",X"56",X"55",X"54",X"53",X"52",X"51",X"50",X"67",X"66",X"65",X"64",X"63",
		X"62",X"61",X"60",X"47",X"46",X"45",X"44",X"43",X"42",X"41",X"00",X"01",X"04",X"02",X"64",X"52",
		X"53",X"40",X"4D",X"02",X"65",X"43",X"53",X"80",X"11",X"02",X"62",X"65",X"53",X"08",X"4B",X"01",
		X"42",X"67",X"40",X"80",X"31",X"01",X"62",X"53",X"40",X"18",X"96",X"00",X"62",X"46",X"53",X"48",
		X"82",X"00",X"46",X"53",X"65",X"50",X"5F",X"00",X"43",X"53",X"65",X"10",X"5C",X"00",X"43",X"44",
		X"40",X"58",X"68",X"00",X"60",X"44",X"43",X"90",X"52",X"00",X"94",X"42",X"95",X"42",X"96",X"42",
		X"97",X"42",X"B0",X"42",X"B1",X"42",X"B2",X"42",X"B3",X"42",X"B4",X"42",X"B5",X"42",X"03",X"02",
		X"01",X"00",X"00",X"80",X"48",X"40",X"E5",X"F0",X"0A",X"E1",X"E5",X"F7",X"0A",X"E1",X"E5",X"5C",
		X"0B",X"E1",X"E5",X"5D",X"0B",X"E1",X"E5",X"81",X"0B",X"E1",X"E5",X"F3",X"0B",X"E1",X"E5",X"F1",
		X"2C",X"E1",X"E5",X"65",X"3D",X"E1",X"E5",X"66",X"3D",X"E1",X"E5",X"67",X"3D",X"E1",X"E5",X"4A",
		X"3D",X"E1",X"E5",X"4B",X"3D",X"E1",X"E5",X"5E",X"3D",X"E1",X"E5",X"5F",X"3D",X"E1",X"E5",X"89",
		X"3D",X"E1",X"E5",X"E3",X"3D",X"E1",X"00",X"FF",X"09",X"2B",X"0B",X"0A",X"50",X"67",X"E1",X"3E",
		X"10",X"1A",X"D0",X"64",X"3E",X"08",X"1A",X"66",X"67",X"3A",X"67",X"67",X"FE",X"07",X"C2",X"6D",
		X"0B",X"AF",X"1A",X"67",X"67",X"3A",X"3C",X"65",X"EE",X"10",X"1A",X"3C",X"65",X"2A",X"50",X"67",
		X"7E",X"FE",X"00",X"28",X"26",X"0B",X"46",X"3A",X"D2",X"64",X"B8",X"28",X"14",X"2B",X"0A",X"50",
		X"67",X"30",X"17",X"0B",X"46",X"3A",X"D3",X"64",X"B8",X"28",X"06",X"2B",X"0A",X"50",X"67",X"30",
		X"21",X"0B",X"7E",X"1A",X"3C",X"65",X"0B",X"0A",X"50",X"67",X"E1",X"01",X"6B",X"26",X"00",X"14",
		X"23",X"01",X"EB",X"07",X"00",X"C4",X"25",X"01",X"D3",X"07",X"00",X"CC",X"25",X"01",X"BB",X"07",
		X"00",X"FC",X"25",X"01",X"53",X"26",X"00",X"CC",X"25",X"01",X"3B",X"26",X"00",X"AC",X"25",X"01",
		X"0B",X"26",X"00",X"64",X"23",X"01",X"53",X"26",X"00",X"14",X"23",X"01",X"BB",X"07",X"00",X"64",
		X"23",X"01",X"D3",X"07",X"00",X"CC",X"25",X"01",X"8B",X"26",X"00",X"14",X"25",X"3C",X"1A",X"67",
		X"67",X"C3",X"FD",X"0A",X"E1",X"09",X"57",X"66",X"0A",X"CF",X"66",X"09",X"EC",X"66",X"0A",X"3C",
		X"67",X"09",X"7D",X"3A",X"11",X"57",X"66",X"01",X"60",X"00",X"ED",X"98",X"09",X"7D",X"3A",X"11",
		X"B7",X"66",X"01",X"60",X"00",X"ED",X"98",X"AF",X"1A",X"42",X"67",X"1A",X"43",X"67",X"1A",X"44",
		X"67",X"3A",X"34",X"66",X"E3",X"A7",X"1A",X"34",X"66",X"3E",X"31",X"1A",X"3E",X"67",X"1A",X"3F",
		X"67",X"1A",X"40",X"67",X"1A",X"41",X"67",X"AF",X"1A",X"45",X"67",X"1A",X"E9",X"66",X"09",X"A7",
		X"3B",X"11",X"EC",X"66",X"01",X"28",X"00",X"ED",X"98",X"09",X"A7",X"3B",X"11",X"14",X"67",X"01",
		X"28",X"00",X"ED",X"98",X"09",X"57",X"66",X"0A",X"CF",X"66",X"E1",X"09",X"A5",X"0C",X"11",X"8F",
		X"64",X"01",X"18",X"00",X"ED",X"98",X"09",X"2F",X"66",X"11",X"18",X"66",X"01",X"35",X"00",X"1E",
		X"00",X"ED",X"98",X"09",X"9F",X"3B",X"0A",X"37",X"66",X"09",X"56",X"3C",X"0A",X"09",X"66",X"09",
		X"15",X"3D",X"0A",X"0B",X"66",X"09",X"19",X"3D",X"0A",X"0D",X"66",X"3E",X"80",X"1A",X"2D",X"66",
		X"3E",X"08",X"1A",X"55",X"66",X"3E",X"40",X"1A",X"06",X"64",X"1A",X"26",X"64",X"1A",X"16",X"64",
		X"1A",X"36",X"64",X"1A",X"0E",X"64",X"1A",X"2E",X"64",X"1A",X"1E",X"64",X"1A",X"3E",X"64",X"1A",
		X"46",X"64",X"1A",X"66",X"64",X"3E",X"48",X"1A",X"05",X"64",X"1A",X"25",X"64",X"1A",X"15",X"64",
		X"1A",X"35",X"64",X"1A",X"0D",X"64",X"1A",X"2D",X"64",X"1A",X"1D",X"64",X"1A",X"3D",X"64",X"1A",
		X"45",X"64",X"1A",X"65",X"64",X"09",X"2C",X"01",X"0A",X"64",X"67",X"30",X"48",X"03",X"00",X"00",
		X"0B",X"1C",X"28",X"07",X"25",X"03",X"00",X"00",X"0B",X"CC",X"28",X"07",X"25",X"04",X"00",X"00",
		X"87",X"14",X"28",X"07",X"FD",X"03",X"00",X"00",X"EB",X"1C",X"28",X"07",X"00",X"03",X"00",X"00",
		X"EB",X"CC",X"28",X"07",X"00",X"05",X"10",X"00",X"87",X"7C",X"0E",X"14",X"DF",X"03",X"00",X"00",
		X"00",X"1C",X"28",X"07",X"25",X"03",X"00",X"00",X"00",X"CC",X"28",X"07",X"25",X"04",X"00",X"00",
		X"00",X"14",X"28",X"07",X"FD",X"03",X"00",X"00",X"00",X"1C",X"28",X"07",X"00",X"03",X"00",X"00",
		X"00",X"CC",X"28",X"07",X"00",X"05",X"10",X"00",X"87",X"7C",X"0E",X"14",X"DF",X"3E",X"40",X"E5",
		X"AD",X"14",X"11",X"82",X"40",X"09",X"13",X"2B",X"3E",X"34",X"06",X"02",X"E5",X"85",X"15",X"3E",
		X"26",X"1A",X"C2",X"40",X"1A",X"F4",X"40",X"3E",X"27",X"1A",X"C3",X"40",X"1A",X"F5",X"40",X"11",
		X"CA",X"40",X"09",X"63",X"2B",X"3E",X"34",X"06",X"02",X"E5",X"85",X"15",X"3E",X"26",X"1A",X"29",
		X"41",X"1A",X"2F",X"41",X"1A",X"1D",X"41",X"3E",X"27",X"1A",X"2A",X"41",X"1A",X"18",X"41",X"1A",
		X"1E",X"41",X"11",X"42",X"41",X"09",X"83",X"2B",X"3E",X"34",X"06",X"02",X"E5",X"85",X"15",X"11",
		X"8A",X"41",X"09",X"BB",X"2B",X"3E",X"34",X"06",X"01",X"E5",X"85",X"15",X"11",X"C2",X"41",X"09",
		X"D7",X"2B",X"3E",X"34",X"06",X"01",X"E5",X"85",X"15",X"11",X"CA",X"41",X"09",X"D7",X"2B",X"3E",
		X"34",X"06",X"01",X"E5",X"85",X"15",X"11",X"02",X"42",X"09",X"D7",X"2B",X"3E",X"34",X"06",X"01",
		X"E5",X"85",X"15",X"11",X"0A",X"42",X"09",X"D7",X"2B",X"3E",X"34",X"06",X"01",X"E5",X"85",X"15",
		X"11",X"42",X"42",X"09",X"DB",X"2B",X"3E",X"34",X"06",X"01",X"E5",X"85",X"15",X"11",X"82",X"42",
		X"09",X"27",X"2C",X"3E",X"34",X"06",X"02",X"E5",X"85",X"15",X"3E",X"26",X"1A",X"E1",X"42",X"1A",
		X"E7",X"42",X"1A",X"D5",X"42",X"3E",X"27",X"1A",X"E2",X"42",X"1A",X"D0",X"42",X"1A",X"D6",X"42",
		X"11",X"CA",X"42",X"09",X"47",X"2C",X"3E",X"34",X"06",X"02",X"E5",X"85",X"15",X"3E",X"26",X"1A",
		X"0A",X"43",X"1A",X"3C",X"43",X"3E",X"27",X"1A",X"0B",X"43",X"1A",X"3D",X"43",X"11",X"42",X"43",
		X"09",X"7F",X"2C",X"3E",X"34",X"06",X"02",X"E5",X"85",X"15",X"11",X"40",X"40",X"09",X"9F",X"2C",
		X"3E",X"08",X"06",X"01",X"E5",X"B3",X"15",X"11",X"88",X"43",X"09",X"B8",X"2C",X"3E",X"08",X"06",
		X"01",X"E5",X"B3",X"15",X"11",X"40",X"40",X"09",X"B9",X"2C",X"3E",X"01",X"06",X"34",X"E5",X"B3",
		X"15",X"11",X"77",X"40",X"09",X"BA",X"2C",X"3E",X"01",X"06",X"34",X"E5",X"B3",X"15",X"3E",X"C4",
		X"1A",X"40",X"40",X"3E",X"C5",X"1A",X"88",X"43",X"3E",X"C2",X"1A",X"77",X"40",X"3E",X"C3",X"1A",
		X"BF",X"43",X"AF",X"1A",X"45",X"67",X"1A",X"E9",X"66",X"1A",X"56",X"66",X"1A",X"4A",X"67",X"3A",
		X"44",X"67",X"09",X"27",X"0E",X"E3",X"0F",X"E5",X"48",X"15",X"76",X"0B",X"56",X"EB",X"E9",X"0F",
		X"0E",X"6F",X"0E",X"9F",X"0E",X"FF",X"0E",X"47",X"0F",X"A7",X"0F",X"D7",X"0F",X"37",X"28",X"4F",
		X"28",X"AF",X"28",X"DF",X"28",X"3F",X"29",X"09",X"00",X"01",X"0A",X"65",X"66",X"09",X"00",X"05",
		X"0A",X"53",X"66",X"3E",X"01",X"E5",X"BD",X"14",X"3E",X"07",X"1A",X"EB",X"66",X"3E",X"31",X"1A",
		X"EA",X"66",X"3E",X"01",X"1A",X"A8",X"64",X"3E",X"03",X"1A",X"98",X"64",X"3E",X"05",X"1A",X"B8",
		X"64",X"3E",X"07",X"1A",X"C0",X"64",X"3E",X"21",X"1A",X"E0",X"64",X"3E",X"FF",X"1A",X"63",X"67",
		X"3E",X"18",X"1A",X"66",X"67",X"06",X"40",X"3E",X"01",X"E5",X"03",X"2B",X"C3",X"84",X"29",X"09",
		X"00",X"02",X"0A",X"65",X"66",X"09",X"50",X"07",X"0A",X"53",X"66",X"3E",X"10",X"E5",X"BD",X"14",
		X"3E",X"07",X"1A",X"EB",X"66",X"3E",X"31",X"1A",X"EA",X"66",X"3E",X"02",X"1A",X"A8",X"64",X"3E",
		X"04",X"1A",X"98",X"64",X"3E",X"06",X"1A",X"B8",X"64",X"3E",X"20",X"1A",X"C0",X"64",X"3E",X"22",
		X"1A",X"E0",X"64",X"3E",X"EF",X"1A",X"63",X"67",X"3E",X"15",X"1A",X"66",X"67",X"06",X"40",X"3E",
		X"02",X"E5",X"03",X"2B",X"C3",X"84",X"29",X"09",X"00",X"03",X"0A",X"65",X"66",X"09",X"00",X"10",
		X"0A",X"53",X"66",X"3E",X"05",X"E5",X"BD",X"14",X"3E",X"07",X"1A",X"EB",X"66",X"3E",X"31",X"1A",
		X"EA",X"66",X"3E",X"03",X"1A",X"A8",X"64",X"3E",X"05",X"1A",X"98",X"64",X"3E",X"07",X"1A",X"B8",
		X"64",X"3E",X"21",X"1A",X"C0",X"64",X"3E",X"23",X"1A",X"E0",X"64",X"3E",X"F7",X"1A",X"63",X"67",
		X"3E",X"08",X"1A",X"66",X"67",X"06",X"40",X"3E",X"03",X"E5",X"03",X"2B",X"C3",X"84",X"29",X"09",
		X"00",X"04",X"0A",X"65",X"66",X"09",X"50",X"12",X"0A",X"53",X"66",X"3E",X"35",X"E5",X"BD",X"14",
		X"3E",X"07",X"1A",X"EB",X"66",X"3E",X"31",X"1A",X"EA",X"66",X"3E",X"04",X"1A",X"A8",X"64",X"3E",
		X"06",X"1A",X"98",X"64",X"3E",X"20",X"1A",X"B8",X"64",X"3E",X"22",X"1A",X"C0",X"64",X"3E",X"24",
		X"1A",X"E0",X"64",X"3E",X"E7",X"1A",X"63",X"67",X"3E",X"10",X"1A",X"66",X"67",X"06",X"40",X"3E",
		X"04",X"E5",X"03",X"2B",X"C3",X"84",X"29",X"09",X"00",X"05",X"0A",X"65",X"66",X"09",X"00",X"15",
		X"0A",X"53",X"66",X"3E",X"21",X"E5",X"BD",X"14",X"3E",X"07",X"1A",X"EB",X"66",X"3E",X"31",X"1A",
		X"EA",X"66",X"3E",X"05",X"1A",X"A8",X"64",X"3E",X"07",X"1A",X"98",X"64",X"3E",X"21",X"1A",X"B8",
		X"64",X"3E",X"23",X"1A",X"C0",X"64",X"3E",X"25",X"1A",X"E0",X"64",X"3E",X"BF",X"1A",X"63",X"67",
		X"3E",X"06",X"1A",X"66",X"67",X"06",X"40",X"3E",X"05",X"E5",X"03",X"2B",X"C3",X"84",X"29",X"09",
		X"00",X"06",X"0A",X"65",X"66",X"09",X"50",X"17",X"0A",X"53",X"66",X"3E",X"01",X"E5",X"BD",X"14",
		X"3E",X"07",X"1A",X"EB",X"66",X"3E",X"31",X"1A",X"EA",X"66",X"3E",X"06",X"1A",X"A8",X"64",X"3E",
		X"20",X"1A",X"98",X"64",X"3E",X"22",X"1A",X"B8",X"64",X"3E",X"24",X"1A",X"C0",X"64",X"3E",X"26",
		X"1A",X"E0",X"64",X"3E",X"BF",X"1A",X"63",X"67",X"3E",X"01",X"1A",X"66",X"67",X"06",X"40",X"3E",
		X"06",X"E5",X"03",X"2B",X"C3",X"84",X"29",X"09",X"00",X"07",X"0A",X"65",X"66",X"09",X"00",X"08",
		X"0A",X"53",X"66",X"3E",X"10",X"E5",X"BD",X"14",X"3E",X"07",X"1A",X"EB",X"66",X"3E",X"31",X"1A",
		X"EA",X"66",X"3E",X"07",X"1A",X"A8",X"64",X"3E",X"21",X"1A",X"98",X"64",X"3E",X"23",X"1A",X"B8",
		X"64",X"3E",X"25",X"1A",X"C0",X"64",X"3E",X"27",X"1A",X"E0",X"64",X"3E",X"BF",X"1A",X"63",X"67",
		X"3E",X"01",X"1A",X"66",X"67",X"06",X"40",X"3E",X"07",X"E5",X"03",X"2B",X"C3",X"84",X"29",X"09",
		X"00",X"20",X"0A",X"65",X"66",X"09",X"50",X"0A",X"0A",X"53",X"66",X"3E",X"05",X"E5",X"BD",X"14",
		X"3E",X"07",X"1A",X"EB",X"66",X"3E",X"31",X"1A",X"EA",X"66",X"3E",X"20",X"1A",X"A8",X"64",X"3E",
		X"22",X"1A",X"98",X"64",X"3E",X"24",X"1A",X"B8",X"64",X"3E",X"26",X"1A",X"C0",X"64",X"3E",X"10",
		X"1A",X"E0",X"64",X"3E",X"BF",X"1A",X"63",X"67",X"3E",X"01",X"1A",X"66",X"67",X"06",X"40",X"3E",
		X"20",X"E5",X"03",X"2B",X"C3",X"84",X"29",X"09",X"00",X"21",X"0A",X"65",X"66",X"09",X"00",X"0D",
		X"0A",X"53",X"66",X"3E",X"35",X"E5",X"BD",X"14",X"3E",X"07",X"1A",X"EB",X"66",X"3E",X"31",X"1A",
		X"EA",X"66",X"3E",X"20",X"1A",X"A8",X"64",X"3E",X"22",X"1A",X"98",X"64",X"3E",X"24",X"1A",X"B8",
		X"64",X"3E",X"26",X"1A",X"C0",X"64",X"3E",X"10",X"1A",X"E0",X"64",X"3E",X"BF",X"1A",X"63",X"67",
		X"3E",X"01",X"1A",X"66",X"67",X"06",X"40",X"3E",X"21",X"E5",X"03",X"2B",X"C3",X"84",X"29",X"09",
		X"00",X"10",X"0A",X"65",X"66",X"09",X"50",X"0F",X"0A",X"53",X"66",X"3E",X"21",X"E5",X"BD",X"14",
		X"3E",X"07",X"1A",X"EB",X"66",X"3E",X"31",X"1A",X"EA",X"66",X"3E",X"20",X"1A",X"A8",X"64",X"3E",
		X"22",X"1A",X"98",X"64",X"3E",X"24",X"1A",X"B8",X"64",X"3E",X"26",X"1A",X"C0",X"64",X"3E",X"10",
		X"1A",X"E0",X"64",X"3E",X"BF",X"1A",X"63",X"67",X"3E",X"01",X"1A",X"66",X"67",X"06",X"01",X"3E",
		X"00",X"E5",X"03",X"2B",X"C3",X"84",X"29",X"09",X"00",X"11",X"0A",X"65",X"66",X"09",X"00",X"18",
		X"0A",X"53",X"66",X"3E",X"01",X"E5",X"BD",X"14",X"3E",X"07",X"1A",X"EB",X"66",X"3E",X"31",X"1A",
		X"EA",X"66",X"3E",X"20",X"1A",X"A8",X"64",X"3E",X"22",X"1A",X"98",X"64",X"3E",X"24",X"1A",X"B8",
		X"64",X"3E",X"26",X"1A",X"C0",X"64",X"3E",X"10",X"1A",X"E0",X"64",X"3E",X"BF",X"1A",X"63",X"67",
		X"3E",X"01",X"1A",X"66",X"67",X"06",X"01",X"3E",X"01",X"E5",X"03",X"2B",X"C3",X"84",X"29",X"09",
		X"00",X"12",X"0A",X"65",X"66",X"09",X"50",X"1A",X"0A",X"53",X"66",X"3E",X"10",X"E5",X"BD",X"14",
		X"3E",X"07",X"1A",X"EB",X"66",X"3E",X"31",X"1A",X"EA",X"66",X"3E",X"20",X"1A",X"A8",X"64",X"3E",
		X"22",X"1A",X"98",X"64",X"3E",X"24",X"1A",X"B8",X"64",X"3E",X"26",X"1A",X"C0",X"64",X"3E",X"10",
		X"1A",X"E0",X"64",X"3E",X"BF",X"1A",X"63",X"67",X"3E",X"01",X"1A",X"66",X"67",X"06",X"01",X"3E",
		X"02",X"E5",X"03",X"2B",X"11",X"49",X"44",X"09",X"EB",X"66",X"3E",X"36",X"06",X"01",X"E5",X"B3",
		X"15",X"11",X"C4",X"44",X"09",X"EB",X"66",X"3E",X"30",X"06",X"01",X"E5",X"B3",X"15",X"11",X"1F",
		X"45",X"09",X"EB",X"66",X"3E",X"20",X"06",X"01",X"E5",X"B3",X"15",X"11",X"19",X"45",X"09",X"EB",
		X"66",X"3E",X"04",X"06",X"01",X"E5",X"B3",X"15",X"11",X"2B",X"45",X"09",X"EB",X"66",X"3E",X"04",
		X"06",X"01",X"E5",X"B3",X"15",X"11",X"09",X"45",X"09",X"EB",X"66",X"3E",X"20",X"06",X"01",X"E5",
		X"B3",X"15",X"11",X"81",X"45",X"09",X"EB",X"66",X"3E",X"36",X"06",X"01",X"E5",X"B3",X"15",X"11",
		X"49",X"46",X"09",X"EB",X"66",X"3E",X"36",X"06",X"01",X"E5",X"B3",X"15",X"11",X"D7",X"46",X"09",
		X"EB",X"66",X"3E",X"05",X"06",X"01",X"E5",X"B3",X"15",X"11",X"D1",X"46",X"09",X"EB",X"66",X"3E",
		X"04",X"06",X"01",X"E5",X"B3",X"15",X"11",X"E3",X"46",X"09",X"EB",X"66",X"3E",X"04",X"06",X"01",
		X"E5",X"B3",X"15",X"11",X"C1",X"46",X"09",X"EB",X"66",X"3E",X"20",X"06",X"01",X"E5",X"B3",X"15",
		X"11",X"0C",X"47",X"09",X"EB",X"66",X"3E",X"30",X"06",X"01",X"E5",X"B3",X"15",X"11",X"81",X"47",
		X"09",X"EB",X"66",X"3E",X"36",X"06",X"01",X"E5",X"B3",X"15",X"11",X"49",X"44",X"09",X"EB",X"66",
		X"3E",X"01",X"06",X"32",X"E5",X"B3",X"15",X"11",X"C4",X"44",X"09",X"EB",X"66",X"3E",X"01",X"06",
		X"14",X"E5",X"B3",X"15",X"11",X"68",X"44",X"09",X"EB",X"66",X"3E",X"01",X"06",X"32",X"E5",X"B3",
		X"15",X"11",X"E3",X"46",X"09",X"EB",X"66",X"3E",X"01",X"06",X"07",X"E5",X"B3",X"15",X"11",X"A3",
		X"45",X"09",X"EB",X"66",X"3E",X"01",X"06",X"20",X"E5",X"B3",X"15",X"11",X"6B",X"44",X"09",X"EB",
		X"66",X"3E",X"01",X"06",X"07",X"E5",X"B3",X"15",X"11",X"E6",X"44",X"09",X"EB",X"66",X"3E",X"01",
		X"06",X"14",X"E5",X"B3",X"15",X"11",X"D1",X"44",X"09",X"EB",X"66",X"3E",X"01",X"06",X"14",X"E5",
		X"B3",X"15",X"11",X"D4",X"46",X"09",X"EB",X"66",X"3E",X"01",X"06",X"07",X"E5",X"B3",X"15",X"11",
		X"94",X"45",X"09",X"EB",X"66",X"3E",X"01",X"06",X"20",X"E5",X"B3",X"15",X"11",X"5C",X"44",X"09",
		X"EB",X"66",X"3E",X"01",X"06",X"07",X"E5",X"B3",X"15",X"11",X"5F",X"44",X"09",X"EB",X"66",X"3E",
		X"01",X"06",X"32",X"E5",X"B3",X"15",X"11",X"F3",X"44",X"09",X"EB",X"66",X"3E",X"01",X"06",X"14",
		X"E5",X"B3",X"15",X"11",X"7E",X"44",X"09",X"EB",X"66",X"3E",X"01",X"06",X"32",X"E5",X"B3",X"15",
		X"3A",X"EA",X"66",X"1A",X"3E",X"67",X"1A",X"3F",X"67",X"1A",X"40",X"67",X"1A",X"41",X"67",X"E5",
		X"BD",X"1F",X"E1",X"1A",X"F9",X"41",X"78",X"1A",X"31",X"42",X"3E",X"21",X"1A",X"F9",X"45",X"1A",
		X"31",X"46",X"E1",X"23",X"11",X"11",X"11",X"11",X"25",X"40",X"23",X"25",X"40",X"23",X"11",X"11",
		X"11",X"11",X"11",X"11",X"25",X"40",X"23",X"25",X"40",X"23",X"11",X"11",X"11",X"11",X"25",X"26",
		X"C4",X"10",X"10",X"10",X"24",X"40",X"22",X"24",X"40",X"22",X"10",X"10",X"10",X"10",X"10",X"10",
		X"24",X"40",X"22",X"24",X"40",X"22",X"10",X"10",X"10",X"C2",X"27",X"26",X"27",X"40",X"23",X"11",
		X"25",X"40",X"23",X"25",X"40",X"23",X"25",X"40",X"23",X"25",X"40",X"23",X"25",X"40",X"23",X"25",
		X"40",X"23",X"11",X"25",X"40",X"26",X"27",X"22",X"24",X"40",X"22",X"10",X"24",X"40",X"26",X"27",
		X"40",X"22",X"24",X"40",X"26",X"27",X"40",X"22",X"24",X"40",X"26",X"27",X"40",X"22",X"10",X"24",
		X"40",X"22",X"24",X"23",X"25",X"40",X"23",X"11",X"25",X"40",X"26",X"C5",X"11",X"11",X"25",X"40",
		X"26",X"27",X"40",X"23",X"11",X"11",X"C3",X"27",X"40",X"23",X"11",X"25",X"40",X"23",X"25",X"22",
		X"24",X"40",X"22",X"10",X"24",X"40",X"22",X"10",X"10",X"10",X"24",X"40",X"22",X"24",X"40",X"22",
		X"10",X"10",X"10",X"24",X"40",X"22",X"10",X"24",X"40",X"22",X"24",X"23",X"25",X"40",X"23",X"11",
		X"25",X"40",X"23",X"25",X"40",X"23",X"25",X"40",X"23",X"25",X"40",X"23",X"25",X"40",X"23",X"25",
		X"40",X"23",X"11",X"25",X"40",X"23",X"25",X"26",X"27",X"40",X"26",X"2E",X"27",X"40",X"26",X"27",
		X"40",X"26",X"27",X"40",X"26",X"27",X"40",X"26",X"27",X"40",X"26",X"27",X"40",X"26",X"40",X"27",
		X"40",X"26",X"27",X"22",X"24",X"40",X"22",X"10",X"24",X"40",X"22",X"24",X"40",X"22",X"24",X"40",
		X"22",X"24",X"40",X"22",X"24",X"40",X"22",X"24",X"40",X"22",X"10",X"24",X"40",X"22",X"24",X"23",
		X"25",X"40",X"23",X"11",X"25",X"40",X"23",X"11",X"11",X"11",X"25",X"40",X"23",X"25",X"40",X"23",
		X"11",X"11",X"11",X"25",X"40",X"23",X"11",X"25",X"40",X"23",X"25",X"22",X"24",X"40",X"22",X"10",
		X"24",X"40",X"26",X"C4",X"10",X"10",X"24",X"40",X"26",X"27",X"40",X"22",X"10",X"10",X"C2",X"27",
		X"40",X"22",X"10",X"24",X"40",X"22",X"24",X"23",X"25",X"40",X"23",X"11",X"25",X"40",X"26",X"27",
		X"40",X"23",X"25",X"40",X"26",X"27",X"40",X"23",X"25",X"40",X"26",X"27",X"40",X"23",X"11",X"25",
		X"40",X"23",X"25",X"26",X"27",X"40",X"22",X"10",X"24",X"40",X"22",X"24",X"40",X"22",X"24",X"40",
		X"22",X"24",X"40",X"22",X"24",X"40",X"22",X"24",X"40",X"22",X"10",X"24",X"40",X"26",X"27",X"26",
		X"C5",X"11",X"11",X"11",X"25",X"40",X"23",X"25",X"40",X"23",X"11",X"11",X"11",X"11",X"11",X"11",
		X"25",X"40",X"23",X"25",X"40",X"23",X"11",X"11",X"11",X"C3",X"27",X"22",X"10",X"10",X"10",X"10",
		X"24",X"40",X"22",X"24",X"40",X"22",X"10",X"10",X"10",X"10",X"10",X"10",X"24",X"40",X"22",X"24",
		X"40",X"22",X"10",X"10",X"10",X"10",X"24",X"10",X"11",X"27",X"26",X"45",X"47",X"47",X"67",X"52",
		X"2C",X"43",X"67",X"50",X"71",X"52",X"61",X"47",X"60",X"54",X"08",X"19",X"39",X"38",X"1B",X"54",
		X"45",X"64",X"63",X"67",X"08",X"61",X"66",X"43",X"5F",X"09",X"4A",X"67",X"E3",X"46",X"C2",X"09",
		X"2D",X"3E",X"0B",X"1A",X"AA",X"64",X"1A",X"9A",X"64",X"3E",X"87",X"1A",X"BA",X"64",X"3E",X"EB",
		X"1A",X"C2",X"64",X"1A",X"E2",X"64",X"0B",X"7E",X"FE",X"20",X"08",X"0A",X"AF",X"5F",X"3A",X"AC",
		X"64",X"C6",X"04",X"1A",X"AC",X"64",X"1A",X"9C",X"64",X"1A",X"BC",X"64",X"1A",X"C4",X"64",X"1A",
		X"E4",X"64",X"FE",X"44",X"C0",X"2B",X"E3",X"C6",X"09",X"AE",X"65",X"E3",X"C6",X"E1",X"3C",X"5F",
		X"E1",X"09",X"62",X"66",X"E3",X"46",X"C2",X"2C",X"1B",X"09",X"00",X"00",X"0A",X"67",X"66",X"09",
		X"E7",X"64",X"0A",X"D7",X"64",X"F5",X"09",X"E7",X"64",X"F5",X"7E",X"07",X"FE",X"80",X"D2",X"99",
		X"2D",X"2A",X"0B",X"66",X"E3",X"0F",X"E5",X"48",X"15",X"0A",X"0F",X"66",X"3A",X"3C",X"65",X"CE",
		X"27",X"47",X"FE",X"27",X"28",X"0E",X"3E",X"10",X"1A",X"D0",X"64",X"78",X"E3",X"47",X"08",X"0D",
		X"2A",X"0F",X"66",X"46",X"F5",X"7E",X"04",X"B8",X"E2",X"54",X"2E",X"F5",X"1E",X"00",X"02",X"06",
		X"34",X"26",X"36",X"E5",X"D6",X"1C",X"E5",X"F0",X"24",X"C3",X"09",X"2E",X"F5",X"7E",X"00",X"FE",
		X"03",X"28",X"06",X"30",X"F3",X"E3",X"77",X"08",X"35",X"2A",X"0F",X"66",X"0B",X"46",X"F5",X"7E",
		X"04",X"B8",X"E2",X"54",X"2E",X"F5",X"1E",X"00",X"03",X"06",X"08",X"26",X"0A",X"E5",X"D6",X"1C",
		X"E5",X"F0",X"24",X"C3",X"09",X"2E",X"F5",X"46",X"04",X"E5",X"E6",X"1B",X"18",X"E6",X"C3",X"1D",
		X"2D",X"CE",X"27",X"2A",X"0D",X"66",X"E3",X"0F",X"E5",X"48",X"15",X"0A",X"0F",X"66",X"3A",X"3C",
		X"65",X"CE",X"27",X"47",X"FE",X"27",X"28",X"0E",X"3E",X"10",X"1A",X"D0",X"64",X"78",X"E3",X"67",
		X"08",X"0D",X"2A",X"0F",X"66",X"46",X"F5",X"7E",X"03",X"B8",X"E2",X"54",X"2E",X"F5",X"1E",X"00",
		X"05",X"06",X"16",X"26",X"32",X"E5",X"D6",X"1C",X"E5",X"F0",X"24",X"C3",X"09",X"2E",X"F5",X"7E",
		X"00",X"FE",X"04",X"28",X"06",X"30",X"F3",X"E3",X"57",X"08",X"33",X"2A",X"0F",X"66",X"0B",X"46",
		X"F5",X"7E",X"03",X"B8",X"28",X"66",X"F5",X"1E",X"00",X"04",X"06",X"14",X"26",X"30",X"E5",X"D6",
		X"1C",X"E5",X"F0",X"24",X"30",X"23",X"F5",X"46",X"03",X"E5",X"E6",X"1B",X"18",X"D0",X"C3",X"1D",
		X"2D",X"3E",X"DB",X"F5",X"46",X"03",X"90",X"1A",X"60",X"66",X"F5",X"7E",X"04",X"D6",X"24",X"1A",
		X"61",X"66",X"3A",X"74",X"67",X"FE",X"05",X"08",X"15",X"AF",X"1A",X"74",X"67",X"3A",X"D4",X"64",
		X"01",X"24",X"00",X"09",X"75",X"1C",X"ED",X"99",X"7E",X"1A",X"D4",X"64",X"30",X"22",X"3C",X"1A",
		X"74",X"67",X"30",X"04",X"F5",X"1E",X"05",X"0E",X"09",X"75",X"0C",X"F5",X"09",X"8F",X"64",X"FD",
		X"09",X"4C",X"67",X"E5",X"86",X"1C",X"FD",X"09",X"2F",X"66",X"FD",X"E3",X"02",X"46",X"28",X"25",
		X"11",X"46",X"67",X"E5",X"D9",X"1C",X"09",X"33",X"66",X"E3",X"86",X"30",X"0B",X"09",X"8F",X"64",
		X"0A",X"D7",X"64",X"E5",X"C9",X"1F",X"3A",X"75",X"67",X"E5",X"1D",X"1C",X"1A",X"75",X"67",X"3E",
		X"DB",X"F5",X"46",X"03",X"90",X"1A",X"2F",X"66",X"F5",X"7E",X"04",X"D6",X"24",X"1A",X"18",X"66",
		X"09",X"19",X"66",X"F5",X"09",X"28",X"64",X"FD",X"09",X"8F",X"64",X"E5",X"C9",X"1D",X"09",X"4D",
		X"0C",X"F5",X"09",X"AF",X"64",X"FD",X"09",X"4D",X"67",X"E5",X"86",X"1C",X"FD",X"09",X"1C",X"66",
		X"FD",X"E3",X"02",X"46",X"28",X"25",X"11",X"47",X"67",X"E5",X"D9",X"1C",X"09",X"33",X"66",X"E3",
		X"86",X"30",X"0B",X"09",X"AF",X"64",X"0A",X"D7",X"64",X"E5",X"C9",X"1F",X"3A",X"76",X"67",X"E5",
		X"1D",X"1C",X"1A",X"76",X"67",X"3E",X"DB",X"F5",X"46",X"03",X"90",X"1A",X"1C",X"66",X"F5",X"7E",
		X"04",X"D6",X"24",X"1A",X"1D",X"66",X"09",X"1E",X"66",X"F5",X"09",X"18",X"64",X"FD",X"09",X"AF",
		X"64",X"E5",X"C9",X"1D",X"09",X"6D",X"0C",X"F5",X"09",X"9F",X"64",X"FD",X"09",X"4E",X"67",X"E5",
		X"86",X"1C",X"FD",X"09",X"39",X"66",X"FD",X"E3",X"02",X"46",X"28",X"25",X"11",X"60",X"67",X"E5",
		X"D9",X"1C",X"09",X"33",X"66",X"E3",X"86",X"30",X"0B",X"09",X"9F",X"64",X"0A",X"D7",X"64",X"E5",
		X"C9",X"1F",X"3A",X"77",X"67",X"E5",X"1D",X"1C",X"1A",X"77",X"67",X"3E",X"DB",X"F5",X"46",X"03",
		X"90",X"1A",X"39",X"66",X"F5",X"7E",X"04",X"D6",X"24",X"1A",X"3A",X"66",X"09",X"3B",X"66",X"F5",
		X"09",X"38",X"64",X"FD",X"09",X"9F",X"64",X"E5",X"C9",X"1D",X"09",X"5D",X"0C",X"F5",X"09",X"BF",
		X"64",X"FD",X"09",X"4F",X"67",X"E5",X"86",X"1C",X"FD",X"09",X"3E",X"66",X"FD",X"E3",X"02",X"46",
		X"28",X"25",X"11",X"61",X"67",X"E5",X"D9",X"1C",X"09",X"33",X"66",X"E3",X"86",X"30",X"0B",X"09",
		X"BF",X"64",X"0A",X"D7",X"64",X"E5",X"C9",X"1F",X"3A",X"48",X"67",X"E5",X"1D",X"1C",X"1A",X"48",
		X"67",X"3E",X"DB",X"F5",X"46",X"03",X"90",X"1A",X"3E",X"66",X"F5",X"7E",X"04",X"D6",X"24",X"1A",
		X"3F",X"66",X"09",X"40",X"66",X"F5",X"09",X"40",X"64",X"FD",X"09",X"BF",X"64",X"E5",X"C9",X"1D",
		X"09",X"7D",X"0C",X"F5",X"09",X"C7",X"64",X"FD",X"09",X"68",X"67",X"E5",X"86",X"1C",X"FD",X"09",
		X"43",X"66",X"FD",X"E3",X"02",X"46",X"28",X"25",X"11",X"62",X"67",X"E5",X"D9",X"1C",X"09",X"33",
		X"66",X"E3",X"86",X"30",X"0B",X"09",X"C7",X"64",X"0A",X"D7",X"64",X"E5",X"C9",X"1F",X"3A",X"49",
		X"67",X"E5",X"1D",X"1C",X"1A",X"49",X"67",X"3E",X"DB",X"F5",X"46",X"03",X"90",X"1A",X"43",X"66",
		X"F5",X"7E",X"04",X"D6",X"24",X"1A",X"44",X"66",X"09",X"45",X"66",X"F5",X"09",X"60",X"64",X"FD",
		X"09",X"C7",X"64",X"E5",X"C9",X"1D",X"09",X"33",X"66",X"E3",X"56",X"C2",X"5C",X"19",X"3A",X"3C",
		X"65",X"E3",X"4F",X"C2",X"DB",X"18",X"F5",X"09",X"00",X"64",X"F5",X"E3",X"06",X"7E",X"28",X"17",
		X"F5",X"09",X"20",X"64",X"F5",X"E3",X"06",X"7E",X"28",X"25",X"F5",X"09",X"10",X"64",X"F5",X"E3",
		X"06",X"7E",X"28",X"03",X"C3",X"DB",X"18",X"F5",X"E3",X"06",X"FE",X"E3",X"D6",X"3A",X"E7",X"64",
		X"F5",X"5F",X"00",X"3A",X"2D",X"66",X"F5",X"5F",X"01",X"3A",X"E7",X"64",X"FE",X"02",X"28",X"26",
		X"FE",X"03",X"28",X"0F",X"3A",X"61",X"66",X"CE",X"F8",X"F5",X"5F",X"03",X"30",X"3B",X"3A",X"61",
		X"66",X"CE",X"F8",X"F5",X"5F",X"03",X"3A",X"D6",X"64",X"CE",X"27",X"E3",X"0F",X"2A",X"0B",X"66",
		X"E5",X"48",X"15",X"7E",X"D6",X"24",X"F5",X"5F",X"07",X"30",X"0F",X"3A",X"61",X"66",X"CE",X"F8",
		X"F5",X"5F",X"03",X"3A",X"D6",X"64",X"CE",X"27",X"E3",X"0F",X"2A",X"0B",X"66",X"E5",X"48",X"15",
		X"0B",X"7E",X"D6",X"24",X"F5",X"5F",X"07",X"30",X"21",X"3A",X"E7",X"64",X"FE",X"04",X"28",X"24",
		X"30",X"29",X"3A",X"60",X"66",X"CE",X"F8",X"F5",X"5F",X"04",X"30",X"3B",X"3A",X"60",X"66",X"CE",
		X"F8",X"F5",X"5F",X"04",X"3A",X"D6",X"64",X"CE",X"27",X"E3",X"0F",X"2A",X"0D",X"66",X"E5",X"48",
		X"15",X"0B",X"3E",X"DB",X"46",X"90",X"F5",X"5F",X"07",X"30",X"34",X"3A",X"60",X"66",X"CE",X"F8",
		X"F5",X"5F",X"04",X"3A",X"D6",X"64",X"CE",X"27",X"E3",X"0F",X"2A",X"0D",X"66",X"E5",X"48",X"15",
		X"3E",X"DB",X"46",X"90",X"F5",X"5F",X"07",X"3A",X"75",X"65",X"FE",X"00",X"08",X"05",X"09",X"78",
		X"65",X"E3",X"C6",X"F5",X"09",X"00",X"64",X"F5",X"E3",X"06",X"7E",X"28",X"27",X"E5",X"21",X"3A",
		X"E5",X"93",X"19",X"09",X"00",X"64",X"0A",X"8C",X"64",X"E5",X"1B",X"25",X"F5",X"09",X"20",X"64",
		X"F5",X"E3",X"06",X"7E",X"28",X"27",X"E5",X"21",X"3A",X"E5",X"93",X"19",X"09",X"20",X"64",X"0A",
		X"8C",X"64",X"E5",X"1B",X"25",X"F5",X"09",X"10",X"64",X"F5",X"E3",X"06",X"7E",X"28",X"27",X"E5",
		X"21",X"3A",X"E5",X"93",X"19",X"09",X"10",X"64",X"0A",X"8C",X"64",X"E5",X"1B",X"25",X"F5",X"09",
		X"30",X"64",X"F5",X"E3",X"06",X"7E",X"28",X"27",X"E5",X"21",X"3A",X"E5",X"93",X"19",X"09",X"30",
		X"64",X"0A",X"8C",X"64",X"E5",X"1B",X"25",X"F5",X"09",X"08",X"64",X"F5",X"E3",X"06",X"7E",X"E2",
		X"46",X"1A",X"E5",X"21",X"3A",X"E5",X"93",X"19",X"09",X"08",X"64",X"0A",X"8C",X"64",X"E5",X"1B",
		X"25",X"C3",X"46",X"1A",X"3A",X"2E",X"66",X"FE",X"20",X"08",X"11",X"3A",X"3C",X"65",X"E3",X"4F",
		X"E2",X"DB",X"18",X"E3",X"96",X"AF",X"1A",X"2E",X"66",X"C3",X"DB",X"18",X"3C",X"1A",X"2E",X"66",
		X"C3",X"DB",X"18",X"F5",X"7E",X"00",X"FE",X"04",X"18",X"12",X"F5",X"7E",X"03",X"F5",X"BE",X"07",
		X"08",X"27",X"F5",X"1E",X"00",X"01",X"F5",X"E3",X"06",X"BE",X"30",X"05",X"F5",X"7E",X"04",X"30",
		X"EC",X"09",X"19",X"66",X"E3",X"46",X"08",X"07",X"2B",X"E5",X"12",X"1A",X"F4",X"DF",X"19",X"09",
		X"1E",X"66",X"E3",X"46",X"08",X"07",X"2B",X"E5",X"12",X"1A",X"F4",X"DF",X"19",X"09",X"3B",X"66",
		X"E3",X"46",X"08",X"07",X"2B",X"E5",X"12",X"1A",X"F4",X"DF",X"19",X"09",X"40",X"66",X"E3",X"46",
		X"08",X"07",X"2B",X"E5",X"12",X"1A",X"F4",X"DF",X"19",X"09",X"45",X"66",X"E3",X"46",X"C0",X"2B",
		X"E5",X"12",X"1A",X"F4",X"DF",X"19",X"E1",X"E3",X"C6",X"09",X"93",X"65",X"E3",X"C6",X"F5",X"1E",
		X"00",X"01",X"F5",X"E3",X"06",X"BE",X"2A",X"65",X"66",X"ED",X"73",X"67",X"66",X"31",X"0A",X"67",
		X"66",X"E1",X"F5",X"7E",X"03",X"46",X"B8",X"38",X"31",X"90",X"FE",X"22",X"18",X"11",X"F5",X"7E",
		X"04",X"2B",X"46",X"B8",X"38",X"16",X"90",X"FE",X"22",X"18",X"04",X"0B",X"0B",X"1F",X"E1",X"1F",
		X"3F",X"E1",X"67",X"78",X"41",X"90",X"FE",X"22",X"38",X"CC",X"30",X"DB",X"67",X"78",X"41",X"90",
		X"FE",X"22",X"38",X"CF",X"30",X"E9",X"00",X"E5",X"BD",X"1F",X"2A",X"64",X"67",X"2B",X"0A",X"64",
		X"67",X"7D",X"9C",X"28",X"02",X"30",X"55",X"3A",X"66",X"67",X"FE",X"04",X"38",X"05",X"D6",X"03",
		X"1A",X"66",X"67",X"3A",X"A8",X"64",X"3C",X"FE",X"21",X"18",X"03",X"1A",X"A8",X"64",X"3A",X"98",
		X"64",X"3C",X"FE",X"22",X"18",X"03",X"1A",X"98",X"64",X"3A",X"B8",X"64",X"3C",X"FE",X"23",X"18",
		X"03",X"1A",X"B8",X"64",X"3A",X"C0",X"64",X"3C",X"FE",X"25",X"18",X"03",X"1A",X"C0",X"64",X"3A",
		X"E0",X"64",X"3C",X"FE",X"10",X"18",X"03",X"1A",X"E0",X"64",X"09",X"2C",X"01",X"0A",X"64",X"67",
		X"3A",X"63",X"67",X"D6",X"08",X"FE",X"0D",X"38",X"03",X"1A",X"63",X"67",X"00",X"09",X"55",X"3B",
		X"3A",X"44",X"67",X"E5",X"48",X"15",X"46",X"3A",X"45",X"67",X"3C",X"1A",X"45",X"67",X"B8",X"C2",
		X"E9",X"1A",X"AF",X"1A",X"45",X"67",X"3A",X"E9",X"66",X"47",X"3A",X"EA",X"66",X"80",X"1A",X"3E",
		X"67",X"1A",X"3F",X"67",X"1A",X"40",X"67",X"1A",X"41",X"67",X"78",X"FE",X"02",X"28",X"06",X"3C",
		X"1A",X"E9",X"66",X"30",X"04",X"AF",X"1A",X"E9",X"66",X"00",X"2A",X"67",X"66",X"EB",X"E5",X"17",
		X"27",X"AF",X"06",X"28",X"2A",X"3C",X"67",X"9E",X"0B",X"10",X"FC",X"FE",X"00",X"C0",X"E5",X"C5",
		X"15",X"E5",X"D8",X"1E",X"09",X"F4",X"64",X"E3",X"E6",X"E3",X"F6",X"E5",X"BD",X"1F",X"3E",X"0E",
		X"1A",X"D4",X"64",X"3E",X"44",X"1A",X"AC",X"64",X"1A",X"9C",X"64",X"1A",X"BC",X"64",X"1A",X"C4",
		X"64",X"1A",X"E4",X"64",X"09",X"CC",X"65",X"E3",X"E6",X"C3",X"5A",X"1B",X"3A",X"F4",X"64",X"E3",
		X"B7",X"1A",X"F4",X"64",X"E3",X"66",X"28",X"0E",X"3A",X"63",X"66",X"FE",X"06",X"08",X"32",X"AF",
		X"1A",X"63",X"66",X"3A",X"E7",X"64",X"FE",X"23",X"28",X"6D",X"3C",X"1A",X"E7",X"64",X"09",X"D5",
		X"1D",X"E5",X"48",X"15",X"7E",X"1A",X"D4",X"64",X"E1",X"3C",X"1A",X"63",X"66",X"E1",X"E3",X"E6",
		X"E5",X"C5",X"15",X"E5",X"D8",X"1E",X"E5",X"BD",X"1F",X"3E",X"17",X"1A",X"D4",X"64",X"AF",X"1A",
		X"E7",X"64",X"AF",X"09",X"19",X"66",X"E3",X"46",X"28",X"03",X"1A",X"AA",X"64",X"09",X"1E",X"66",
		X"E3",X"46",X"28",X"03",X"1A",X"9A",X"64",X"09",X"3B",X"66",X"E3",X"46",X"28",X"03",X"1A",X"BA",
		X"64",X"09",X"40",X"66",X"E3",X"46",X"28",X"03",X"1A",X"C2",X"64",X"09",X"45",X"66",X"E3",X"46",
		X"28",X"03",X"1A",X"E2",X"64",X"3E",X"44",X"1A",X"AC",X"64",X"1A",X"9C",X"64",X"1A",X"BC",X"64",
		X"1A",X"C4",X"64",X"1A",X"E4",X"64",X"E1",X"AF",X"1A",X"D2",X"64",X"09",X"2F",X"66",X"11",X"18",
		X"66",X"01",X"35",X"00",X"1E",X"00",X"ED",X"98",X"09",X"F4",X"64",X"E3",X"E6",X"E1",X"2A",X"37",
		X"66",X"F5",X"7E",X"07",X"FE",X"80",X"38",X"03",X"2A",X"09",X"66",X"CE",X"27",X"E3",X"0F",X"E3",
		X"0F",X"E5",X"48",X"15",X"7E",X"DD",X"0B",X"76",X"0B",X"56",X"EB",X"7E",X"B8",X"28",X"25",X"0B",
		X"0B",X"D9",X"3D",X"DD",X"28",X"02",X"30",X"DB",X"D9",X"1F",X"3F",X"E1",X"D9",X"2B",X"7E",X"DD",
		X"2A",X"0B",X"66",X"FE",X"80",X"38",X"03",X"2A",X"0D",X"66",X"CE",X"27",X"E3",X"0F",X"E5",X"48",
		X"15",X"3A",X"3C",X"65",X"E3",X"67",X"28",X"15",X"E3",X"47",X"28",X"05",X"0B",X"E3",X"57",X"28",
		X"24",X"7E",X"F5",X"BE",X"04",X"28",X"D1",X"D9",X"F5",X"5F",X"07",X"1F",X"E1",X"7E",X"F5",X"BE",
		X"03",X"28",X"C5",X"30",X"DA",X"67",X"F5",X"7E",X"05",X"FE",X"44",X"E0",X"F5",X"7E",X"01",X"09",
		X"5D",X"1C",X"E5",X"48",X"15",X"7E",X"B9",X"38",X"03",X"79",X"3C",X"E1",X"F5",X"7E",X"05",X"01",
		X"24",X"00",X"09",X"69",X"1C",X"ED",X"99",X"7E",X"F5",X"5F",X"05",X"AF",X"E1",X"34",X"36",X"34",
		X"08",X"0A",X"08",X"16",X"32",X"16",X"14",X"30",X"14",X"24",X"26",X"24",X"10",X"12",X"10",X"04",
		X"20",X"04",X"06",X"22",X"06",X"00",X"10",X"27",X"26",X"25",X"24",X"23",X"22",X"21",X"20",X"07",
		X"06",X"05",X"04",X"03",X"02",X"01",X"F5",X"E3",X"06",X"7E",X"28",X"36",X"F5",X"E3",X"06",X"5E",
		X"08",X"2A",X"3E",X"40",X"FD",X"BE",X"00",X"08",X"36",X"FD",X"1E",X"00",X"00",X"F5",X"E3",X"06",
		X"DE",X"CD",X"09",X"85",X"0C",X"0A",X"35",X"66",X"C9",X"E1",X"FD",X"1E",X"00",X"00",X"CD",X"09",
		X"E7",X"64",X"0A",X"35",X"66",X"C9",X"E1",X"FD",X"1C",X"00",X"30",X"DA",X"3E",X"40",X"FD",X"BE",
		X"00",X"08",X"26",X"FD",X"1E",X"00",X"00",X"F5",X"E3",X"06",X"9E",X"F5",X"E3",X"06",X"BE",X"30",
		X"F5",X"FD",X"1C",X"00",X"30",X"E3",X"2A",X"35",X"66",X"7D",X"FE",X"E7",X"08",X"20",X"F5",X"E3",
		X"06",X"9E",X"F5",X"E3",X"06",X"BE",X"F5",X"7E",X"05",X"B8",X"E0",X"B9",X"E0",X"F5",X"58",X"05",
		X"E1",X"FD",X"E3",X"02",X"66",X"08",X"52",X"FD",X"E3",X"02",X"56",X"28",X"0E",X"FD",X"7E",X"03",
		X"FE",X"06",X"08",X"32",X"FD",X"1E",X"03",X"00",X"F5",X"7E",X"00",X"FE",X"23",X"28",X"19",X"3C",
		X"F5",X"5F",X"00",X"09",X"E1",X"1D",X"E5",X"48",X"15",X"7E",X"F5",X"5F",X"05",X"E1",X"3C",X"FD",
		X"5F",X"03",X"E1",X"F5",X"1E",X"05",X"07",X"F5",X"7E",X"01",X"12",X"F5",X"1E",X"01",X"00",X"F5",
		X"1E",X"00",X"00",X"FD",X"1E",X"03",X"00",X"FD",X"1E",X"04",X"00",X"FD",X"E3",X"02",X"D6",X"E1",
		X"FD",X"E3",X"02",X"E6",X"F5",X"1E",X"03",X"00",X"E1",X"FD",X"46",X"03",X"3A",X"63",X"67",X"B8",
		X"38",X"05",X"04",X"FD",X"58",X"03",X"E1",X"F5",X"7E",X"03",X"FE",X"00",X"08",X"36",X"F5",X"CD",
		X"CD",X"F5",X"C9",X"F5",X"7E",X"07",X"FE",X"FD",X"28",X"18",X"3A",X"D2",X"64",X"F5",X"46",X"03",
		X"B8",X"F5",X"C9",X"E0",X"F5",X"7E",X"03",X"FE",X"00",X"E4",X"8A",X"1D",X"FD",X"7E",X"04",X"FE",
		X"20",X"08",X"12",X"AF",X"FD",X"1E",X"04",X"00",X"F5",X"7E",X"05",X"FE",X"44",X"28",X"0D",X"C6",
		X"04",X"F5",X"5F",X"05",X"E1",X"3C",X"FD",X"5F",X"04",X"E1",X"3A",X"D3",X"64",X"F5",X"46",X"04",
		X"30",X"E6",X"D5",X"F5",X"CD",X"D1",X"01",X"20",X"00",X"ED",X"98",X"D1",X"CD",X"09",X"AE",X"65",
		X"E3",X"C6",X"C9",X"E1",X"FD",X"1E",X"00",X"00",X"FD",X"1E",X"01",X"00",X"FD",X"1E",X"02",X"00",
		X"FD",X"1E",X"03",X"00",X"32",X"F5",X"5F",X"01",X"E1",X"07",X"25",X"05",X"21",X"07",X"25",X"05",
		X"21",X"07",X"25",X"05",X"21",X"17",X"35",X"15",X"31",X"17",X"35",X"15",X"31",X"17",X"35",X"15",
		X"31",X"F5",X"E3",X"06",X"7E",X"28",X"1C",X"F5",X"7E",X"00",X"FE",X"04",X"18",X"28",X"F5",X"7E",
		X"03",X"F5",X"BE",X"07",X"08",X"27",X"F5",X"1E",X"00",X"01",X"F5",X"E3",X"06",X"BE",X"3A",X"56",
		X"66",X"3D",X"1A",X"56",X"66",X"09",X"61",X"66",X"E5",X"12",X"1A",X"F2",X"E8",X"1E",X"F5",X"0A",
		X"8C",X"64",X"E5",X"1B",X"25",X"E1",X"F5",X"7E",X"04",X"30",X"D6",X"E3",X"46",X"C0",X"3A",X"33",
		X"66",X"E3",X"47",X"28",X"3A",X"0B",X"7E",X"3D",X"5F",X"FE",X"00",X"C0",X"3A",X"66",X"67",X"5F",
		X"2B",X"3A",X"56",X"66",X"FE",X"02",X"E0",X"3C",X"1A",X"56",X"66",X"F5",X"E3",X"06",X"FE",X"FD",
		X"7E",X"00",X"F5",X"5F",X"00",X"3A",X"55",X"66",X"F5",X"5F",X"01",X"2B",X"FD",X"7E",X"00",X"FE",
		X"02",X"28",X"12",X"FE",X"03",X"28",X"2A",X"7E",X"CE",X"F8",X"F5",X"5F",X"03",X"30",X"3F",X"3A",
		X"66",X"67",X"0B",X"5F",X"E1",X"CD",X"7E",X"CE",X"F8",X"F5",X"5F",X"03",X"FD",X"7E",X"07",X"CE",
		X"27",X"E3",X"0F",X"2A",X"0B",X"66",X"E5",X"48",X"15",X"7E",X"D6",X"24",X"F5",X"5F",X"07",X"30",
		X"0F",X"CD",X"7E",X"CE",X"F8",X"F5",X"5F",X"03",X"FD",X"7E",X"07",X"CE",X"27",X"E3",X"0F",X"2A",
		X"0B",X"66",X"E5",X"48",X"15",X"0B",X"7E",X"D6",X"24",X"F5",X"5F",X"07",X"30",X"22",X"2B",X"FD",
		X"7E",X"00",X"FE",X"04",X"28",X"23",X"30",X"0D",X"C9",X"2B",X"7E",X"CE",X"F8",X"F5",X"5F",X"04",
		X"E1",X"7E",X"CE",X"F8",X"F5",X"5F",X"04",X"FD",X"7E",X"07",X"CE",X"27",X"E3",X"0F",X"2A",X"0D",
		X"66",X"E5",X"48",X"15",X"0B",X"3E",X"DB",X"46",X"90",X"F5",X"5F",X"07",X"E1",X"7E",X"CE",X"F8",
		X"F5",X"5F",X"04",X"FD",X"7E",X"07",X"CE",X"27",X"E3",X"0F",X"2A",X"0D",X"66",X"E5",X"48",X"15",
		X"3E",X"DB",X"46",X"90",X"F5",X"5F",X"07",X"E1",X"E3",X"C6",X"09",X"E1",X"65",X"E3",X"C6",X"E1",
		X"F5",X"09",X"00",X"64",X"F5",X"E3",X"06",X"7E",X"28",X"27",X"F5",X"1E",X"00",X"01",X"F5",X"E3",
		X"06",X"BE",X"F5",X"0A",X"8C",X"64",X"E5",X"1B",X"25",X"F5",X"09",X"20",X"64",X"F5",X"E3",X"06",
		X"7E",X"28",X"27",X"F5",X"1E",X"00",X"01",X"F5",X"E3",X"06",X"BE",X"F5",X"0A",X"8C",X"64",X"E5",
		X"1B",X"25",X"F5",X"09",X"10",X"64",X"F5",X"E3",X"06",X"7E",X"28",X"27",X"F5",X"1E",X"00",X"01",
		X"F5",X"E3",X"06",X"BE",X"F5",X"0A",X"8C",X"64",X"E5",X"1B",X"25",X"F5",X"09",X"28",X"64",X"F5",
		X"E3",X"06",X"7E",X"28",X"27",X"F5",X"1E",X"00",X"01",X"F5",X"E3",X"06",X"BE",X"F5",X"0A",X"8C",
		X"64",X"E5",X"1B",X"25",X"F5",X"09",X"18",X"64",X"F5",X"E3",X"06",X"7E",X"28",X"27",X"F5",X"1E",
		X"00",X"01",X"F5",X"E3",X"06",X"BE",X"F5",X"0A",X"8C",X"64",X"E5",X"1B",X"25",X"F5",X"09",X"38",
		X"64",X"F5",X"E3",X"06",X"7E",X"28",X"27",X"F5",X"1E",X"00",X"01",X"F5",X"E3",X"06",X"BE",X"F5",
		X"0A",X"8C",X"64",X"E5",X"1B",X"25",X"F5",X"09",X"40",X"64",X"F5",X"E3",X"06",X"7E",X"28",X"27",
		X"F5",X"1E",X"00",X"01",X"F5",X"E3",X"06",X"BE",X"F5",X"0A",X"8C",X"64",X"E5",X"1B",X"25",X"F5",
		X"09",X"60",X"64",X"F5",X"E3",X"06",X"7E",X"28",X"27",X"F5",X"1E",X"00",X"01",X"F5",X"E3",X"06",
		X"BE",X"F5",X"0A",X"8C",X"64",X"E5",X"1B",X"25",X"AF",X"1A",X"56",X"66",X"E1",X"2A",X"CF",X"66",
		X"3A",X"3E",X"67",X"06",X"04",X"E5",X"C5",X"3A",X"3A",X"3F",X"67",X"06",X"24",X"E5",X"C5",X"3A",
		X"3A",X"40",X"67",X"06",X"10",X"E5",X"C5",X"3A",X"3A",X"41",X"67",X"06",X"04",X"E5",X"C5",X"3A",
		X"E1",X"09",X"33",X"66",X"E3",X"86",X"E3",X"A6",X"2A",X"35",X"66",X"EB",X"FD",X"09",X"00",X"00",
		X"FD",X"31",X"2A",X"D7",X"64",X"EB",X"F5",X"09",X"00",X"00",X"F5",X"31",X"F5",X"7E",X"07",X"FE",
		X"80",X"D2",X"EC",X"38",X"F5",X"46",X"04",X"FD",X"7E",X"04",X"B8",X"F2",X"9F",X"38",X"F5",X"7E",
		X"07",X"FD",X"46",X"07",X"B8",X"E2",X"5F",X"38",X"E5",X"D4",X"39",X"09",X"33",X"66",X"E3",X"66",
		X"C4",X"B7",X"38",X"2A",X"29",X"66",X"7E",X"FD",X"46",X"04",X"2A",X"2B",X"66",X"DD",X"30",X"07",
		X"0B",X"0B",X"D9",X"3D",X"DD",X"28",X"20",X"7E",X"B8",X"28",X"06",X"18",X"DB",X"30",X"02",X"2B",
		X"2B",X"D9",X"F5",X"46",X"04",X"7E",X"B8",X"28",X"08",X"38",X"27",X"F5",X"1E",X"00",X"03",X"06",
		X"10",X"26",X"12",X"E5",X"D6",X"1C",X"E5",X"F0",X"24",X"E1",X"F5",X"1E",X"00",X"02",X"06",X"24",
		X"26",X"26",X"E5",X"D6",X"1C",X"E5",X"F0",X"24",X"E1",X"2B",X"7E",X"F5",X"5F",X"07",X"F5",X"1E",
		X"05",X"44",X"F5",X"E3",X"06",X"FE",X"E1",X"09",X"33",X"66",X"E3",X"C6",X"F5",X"1E",X"00",X"03",
		X"06",X"10",X"26",X"12",X"E5",X"D6",X"1C",X"E5",X"F0",X"24",X"E1",X"09",X"33",X"66",X"E3",X"C6",
		X"F5",X"1E",X"00",X"02",X"06",X"24",X"26",X"26",X"E5",X"D6",X"1C",X"E5",X"F0",X"24",X"E1",X"FD",
		X"7E",X"03",X"F5",X"46",X"03",X"B8",X"38",X"22",X"90",X"FE",X"21",X"D0",X"09",X"33",X"66",X"E3",
		X"C6",X"E1",X"67",X"78",X"41",X"30",X"D9",X"F5",X"7E",X"07",X"FD",X"46",X"07",X"B8",X"E2",X"A3",
		X"38",X"E5",X"D4",X"39",X"09",X"33",X"66",X"E3",X"66",X"C4",X"B7",X"38",X"2A",X"29",X"66",X"7E",
		X"FD",X"46",X"04",X"2A",X"2B",X"66",X"DD",X"30",X"07",X"0B",X"0B",X"D9",X"3D",X"DD",X"28",X"07",
		X"7E",X"B8",X"E2",X"41",X"38",X"18",X"DA",X"2B",X"2B",X"C3",X"41",X"38",X"F5",X"46",X"03",X"FD",
		X"7E",X"03",X"B8",X"F2",X"B7",X"39",X"F5",X"7E",X"07",X"FD",X"46",X"07",X"B8",X"E2",X"77",X"39",
		X"E5",X"D4",X"39",X"09",X"33",X"66",X"E3",X"66",X"C4",X"87",X"39",X"2A",X"29",X"66",X"7E",X"FD",
		X"46",X"03",X"2A",X"2B",X"66",X"DD",X"30",X"07",X"0B",X"0B",X"D9",X"3D",X"DD",X"28",X"20",X"7E",
		X"B8",X"28",X"06",X"18",X"DB",X"30",X"02",X"2B",X"2B",X"D9",X"F5",X"46",X"03",X"7E",X"B8",X"28",
		X"08",X"38",X"27",X"F5",X"1E",X"00",X"04",X"06",X"04",X"26",X"20",X"E5",X"D6",X"1C",X"E5",X"F0",
		X"24",X"E1",X"F5",X"1E",X"00",X"05",X"06",X"06",X"26",X"22",X"E5",X"D6",X"1C",X"E5",X"F0",X"24",
		X"E1",X"2B",X"7E",X"F5",X"5F",X"07",X"F5",X"1E",X"05",X"44",X"F5",X"E3",X"06",X"FE",X"E1",X"09",
		X"33",X"66",X"E3",X"C6",X"F5",X"1E",X"00",X"04",X"06",X"04",X"26",X"20",X"E5",X"D6",X"1C",X"E5",
		X"F0",X"24",X"E1",X"09",X"33",X"66",X"E3",X"C6",X"F5",X"1E",X"00",X"05",X"06",X"06",X"26",X"22",
		X"E5",X"D6",X"1C",X"E5",X"F0",X"24",X"E1",X"FD",X"7E",X"04",X"F5",X"46",X"04",X"B8",X"38",X"22",
		X"90",X"FE",X"21",X"D0",X"09",X"33",X"66",X"E3",X"C6",X"E1",X"67",X"78",X"41",X"30",X"D9",X"F5",
		X"7E",X"07",X"FD",X"46",X"07",X"B8",X"E2",X"5B",X"39",X"E5",X"D4",X"39",X"09",X"33",X"66",X"E3",
		X"66",X"C4",X"87",X"39",X"2A",X"29",X"66",X"7E",X"FD",X"46",X"03",X"2A",X"2B",X"66",X"DD",X"30",
		X"07",X"0B",X"0B",X"D9",X"3D",X"DD",X"28",X"07",X"7E",X"B8",X"E2",X"29",X"39",X"18",X"DA",X"2B",
		X"2B",X"C3",X"29",X"39",X"2A",X"37",X"66",X"F5",X"7E",X"07",X"FE",X"80",X"38",X"03",X"2A",X"09",
		X"66",X"CE",X"27",X"E3",X"0F",X"E3",X"0F",X"E5",X"48",X"15",X"0A",X"29",X"66",X"46",X"FD",X"7E",
		X"07",X"0B",X"76",X"0B",X"56",X"EB",X"0A",X"2B",X"66",X"2B",X"66",X"B9",X"28",X"05",X"0B",X"0B",
		X"10",X"F8",X"E1",X"09",X"33",X"66",X"E3",X"E6",X"E1",X"06",X"22",X"F5",X"7E",X"03",X"09",X"75",
		X"3B",X"BE",X"28",X"06",X"0B",X"10",X"FA",X"C3",X"7C",X"3A",X"78",X"3E",X"22",X"90",X"2A",X"3C",
		X"67",X"E3",X"0F",X"E3",X"0F",X"E5",X"48",X"15",X"F5",X"7E",X"04",X"46",X"B8",X"28",X"12",X"0B",
		X"46",X"B8",X"28",X"25",X"0B",X"46",X"B8",X"28",X"20",X"0B",X"46",X"B8",X"28",X"03",X"C3",X"7C",
		X"3A",X"1E",X"00",X"F5",X"1E",X"00",X"01",X"F5",X"E3",X"06",X"BE",X"1F",X"3F",X"ED",X"73",X"3C",
		X"67",X"ED",X"52",X"EB",X"09",X"4F",X"3B",X"31",X"7E",X"2A",X"CF",X"66",X"E3",X"0F",X"E5",X"48",
		X"15",X"76",X"1E",X"FF",X"0B",X"56",X"1E",X"FF",X"EB",X"1E",X"40",X"2A",X"53",X"66",X"ED",X"73",
		X"67",X"66",X"31",X"0A",X"67",X"66",X"09",X"2C",X"01",X"0A",X"64",X"67",X"E1",X"A6",X"41",X"91",
		X"41",X"59",X"42",X"6E",X"42",X"A0",X"41",X"2B",X"41",X"E6",X"40",X"D1",X"40",X"1C",X"41",X"97",
		X"41",X"5F",X"42",X"D4",X"42",X"19",X"43",X"2E",X"43",X"E3",X"42",X"68",X"42",X"81",X"41",X"0C",
		X"41",X"E0",X"40",X"6B",X"40",X"5C",X"40",X"D7",X"40",X"3B",X"41",X"B6",X"41",X"7E",X"42",X"F3",
		X"42",X"1F",X"43",X"94",X"43",X"A3",X"43",X"28",X"43",X"C4",X"42",X"49",X"42",X"49",X"40",X"7E",
		X"40",X"B6",X"43",X"81",X"43",X"76",X"0B",X"56",X"12",X"0B",X"10",X"F9",X"E1",X"3E",X"21",X"1A",
		X"52",X"67",X"AF",X"1A",X"AA",X"64",X"1A",X"9A",X"64",X"1A",X"BA",X"64",X"1A",X"C2",X"64",X"1A",
		X"E2",X"64",X"1A",X"D2",X"64",X"3E",X"02",X"1A",X"53",X"67",X"3E",X"20",X"1A",X"54",X"67",X"1A",
		X"56",X"67",X"3E",X"20",X"1A",X"55",X"67",X"1A",X"71",X"67",X"3E",X"16",X"1A",X"57",X"67",X"1A",
		X"73",X"67",X"3E",X"12",X"1A",X"70",X"67",X"1A",X"72",X"67",X"ED",X"73",X"54",X"67",X"E5",X"46",
		X"3B",X"ED",X"73",X"56",X"67",X"E5",X"46",X"3B",X"ED",X"73",X"70",X"67",X"E5",X"46",X"3B",X"ED",
		X"73",X"72",X"67",X"E5",X"46",X"3B",X"3A",X"53",X"67",X"C6",X"02",X"1A",X"53",X"67",X"06",X"20",
		X"09",X"54",X"67",X"1D",X"0B",X"10",X"FC",X"3E",X"05",X"E5",X"63",X"15",X"3A",X"52",X"67",X"3D",
		X"1A",X"52",X"67",X"08",X"C5",X"E1",X"E5",X"A7",X"14",X"09",X"54",X"3B",X"3A",X"53",X"67",X"47",
		X"E5",X"B3",X"15",X"E1",X"2E",X"05",X"04",X"03",X"22",X"06",X"03",X"22",X"05",X"20",X"08",X"40",
		X"70",X"58",X"A0",X"88",X"B8",X"F0",X"D8",X"08",X"10",X"37",X"0B",X"11",X"36",X"00",X"00",X"12",
		X"04",X"27",X"35",X"13",X"05",X"26",X"34",X"06",X"00",X"03",X"25",X"07",X"01",X"02",X"24",X"14",
		X"20",X"23",X"33",X"15",X"21",X"22",X"32",X"16",X"31",X"00",X"00",X"09",X"17",X"30",X"0A",X"20",
		X"50",X"A0",X"D0",X"38",X"88",X"00",X"00",X"08",X"50",X"A0",X"B8",X"20",X"38",X"88",X"D0",X"08",
		X"50",X"A0",X"B8",X"08",X"50",X"A0",X"B8",X"20",X"38",X"88",X"D0",X"08",X"50",X"A0",X"B8",X"38",
		X"88",X"00",X"00",X"20",X"50",X"A0",X"D0",X"06",X"EF",X"3B",X"00",X"20",X"FB",X"3B",X"00",X"03",
		X"23",X"3C",X"00",X"02",X"11",X"3C",X"00",X"02",X"15",X"3C",X"00",X"03",X"31",X"3C",X"00",X"22",
		X"37",X"3C",X"00",X"22",X"37",X"3C",X"00",X"03",X"23",X"3C",X"00",X"02",X"1B",X"3C",X"00",X"02",
		X"1F",X"3C",X"00",X"03",X"31",X"3C",X"00",X"20",X"3B",X"3C",X"00",X"06",X"63",X"3C",X"D8",X"FC",
		X"DA",X"C4",X"DD",X"AC",X"FA",X"4C",X"FB",X"64",X"FD",X"14",X"D9",X"CC",X"DA",X"C4",X"DD",X"AC",
		X"DE",X"94",X"DF",X"7C",X"FA",X"4C",X"FB",X"64",X"FC",X"2C",X"D8",X"FC",X"D9",X"CC",X"DA",X"C4",
		X"DD",X"AC",X"DE",X"94",X"DF",X"7C",X"FA",X"4C",X"FB",X"64",X"FC",X"2C",X"FD",X"14",X"D8",X"FC",
		X"D9",X"CC",X"DA",X"C4",X"DC",X"AC",X"DE",X"94",X"DF",X"7C",X"F9",X"4C",X"FB",X"64",X"FC",X"2C",
		X"FD",X"14",X"DB",X"AC",X"DE",X"94",X"DF",X"7C",X"F8",X"4C",X"D9",X"CC",X"DA",X"C4",X"DB",X"AC",
		X"DE",X"94",X"DF",X"7C",X"F8",X"4C",X"FB",X"64",X"FC",X"2C",X"D8",X"FC",X"DA",X"C4",X"DB",X"AC",
		X"F8",X"4C",X"FB",X"64",X"FD",X"14",X"06",X"A6",X"3C",X"00",X"06",X"B2",X"3C",X"00",X"20",X"8E",
		X"3C",X"00",X"03",X"9E",X"3C",X"00",X"02",X"BC",X"3C",X"00",X"03",X"C0",X"3C",X"00",X"06",X"C6",
		X"3C",X"00",X"06",X"D2",X"3C",X"00",X"03",X"F6",X"3C",X"00",X"02",X"CC",X"3C",X"00",X"03",X"E8",
		X"3C",X"00",X"20",X"EE",X"3C",X"00",X"06",X"FE",X"3C",X"00",X"06",X"22",X"3D",X"00",X"EB",X"02",
		X"BB",X"06",X"8B",X"07",X"6B",X"20",X"53",X"25",X"0B",X"01",X"D3",X"02",X"BB",X"06",X"8B",X"07",
		X"6B",X"20",X"53",X"24",X"3B",X"00",X"EB",X"01",X"D3",X"02",X"BB",X"06",X"8B",X"07",X"6B",X"20",
		X"53",X"24",X"3B",X"25",X"0B",X"21",X"53",X"24",X"3B",X"25",X"0B",X"06",X"8B",X"07",X"6B",X"00",
		X"EB",X"01",X"D3",X"03",X"BB",X"01",X"D3",X"03",X"BB",X"06",X"8B",X"07",X"6B",X"21",X"53",X"24",
		X"3B",X"01",X"D3",X"04",X"BB",X"06",X"8B",X"07",X"6B",X"22",X"53",X"24",X"3B",X"22",X"53",X"24",
		X"3B",X"25",X"0B",X"06",X"8B",X"07",X"6B",X"00",X"EB",X"01",X"D3",X"04",X"BB",X"00",X"EB",X"01",
		X"D3",X"05",X"BB",X"06",X"8B",X"07",X"6B",X"23",X"53",X"24",X"3B",X"25",X"0B",X"01",X"D3",X"05",
		X"BB",X"06",X"8B",X"07",X"6B",X"23",X"53",X"24",X"3B",X"00",X"EB",X"05",X"BB",X"06",X"8B",X"07",
		X"6B",X"23",X"53",X"25",X"0B",X"14",X"FC",X"2C",X"CC",X"C4",X"FC",X"94",X"AC",X"4C",X"7C",X"14",
		X"64",X"14",X"FC",X"14",X"FC",X"C4",X"FC",X"94",X"AC",X"4C",X"7C",X"14",X"64",X"2C",X"CC",X"14",
		X"FC",X"0B",X"EB",X"3B",X"D3",X"0B",X"EB",X"0B",X"53",X"6B",X"8B",X"BB",X"EB",X"3B",X"D3",X"3B",
		X"D3",X"0B",X"53",X"6B",X"8B",X"BB",X"EB",X"0B",X"EB",X"3B",X"D3",X"0B",X"EB",X"E1",X"E1",X"09",
		X"57",X"66",X"0A",X"CF",X"66",X"09",X"EC",X"66",X"0A",X"3C",X"67",X"3A",X"42",X"67",X"1A",X"44",
		X"67",X"E1",X"E1",X"09",X"B7",X"66",X"0A",X"CF",X"66",X"09",X"14",X"67",X"0A",X"3C",X"67",X"3A",
		X"43",X"67",X"1A",X"44",X"67",X"E1",X"E1",X"09",X"7D",X"3A",X"11",X"57",X"66",X"01",X"60",X"00",
		X"ED",X"98",X"09",X"A7",X"3B",X"11",X"EC",X"66",X"01",X"28",X"00",X"ED",X"98",X"3A",X"42",X"67",
		X"3C",X"FE",X"24",X"08",X"02",X"3E",X"23",X"1A",X"42",X"67",X"1A",X"44",X"67",X"E5",X"E5",X"3A",
		X"E1",X"09",X"7D",X"3A",X"11",X"B7",X"66",X"01",X"60",X"00",X"ED",X"98",X"09",X"A7",X"3B",X"11",
		X"14",X"67",X"01",X"28",X"00",X"ED",X"98",X"3A",X"43",X"67",X"3C",X"FE",X"24",X"08",X"02",X"3E",
		X"23",X"1A",X"43",X"67",X"1A",X"44",X"67",X"E5",X"E5",X"3A",X"E1",X"E1",X"45",X"47",X"47",X"67",
		X"52",X"2C",X"43",X"67",X"50",X"71",X"52",X"61",X"47",X"60",X"54",X"08",X"19",X"39",X"38",X"1B",
		X"54",X"45",X"64",X"63",X"67",X"08",X"61",X"66",X"43",X"B7",X"86",X"10",X"97",X"E5",X"52",X"54",
		X"8A",X"09",X"96",X"10",X"C5",X"64",X"54",X"61",X"54",X"0B",X"12",X"A3",X"E5",X"71",X"53",X"91",
		X"32",X"96",X"40",X"C2",X"55",X"53",X"66",X"09",X"F2",X"90",X"C7",X"66",X"61",X"52",X"54",X"53",
		X"3E",X"08",X"95",X"C5",X"64",X"54",X"61",X"54",X"53",X"32",X"37",X"A4",X"E4",X"52",X"53",X"8F",
		X"10",X"F1",X"38",X"C1",X"52",X"53",X"0B",X"15",X"F1",X"28",X"C5",X"43",X"41",X"50",X"53",X"0D",
		X"37",X"A1",X"D0",X"53",X"78",X"00",X"F8",X"18",X"C1",X"64",X"53",X"C2",X"33",X"F1",X"08",X"D2",
		X"60",X"53",X"9C",X"33",X"B7",X"E4",X"60",X"53",X"54",X"36",X"B6",X"D4",X"45",X"53",X"F6",X"33",
		X"F0",X"C0",X"C7",X"45",X"53",X"94",X"00",X"B2",X"E6",X"67",X"61",X"54",X"43",X"45",X"53",X"CA",
		X"14",X"8A",X"00",X"C6",X"43",X"53",X"79",X"37",X"D1",X"1F",X"D2",X"41",X"64",X"41",X"43",X"53",
		X"9E",X"27",X"8F",X"C3",X"42",X"53",X"A0",X"37",X"F4",X"B0",X"42",X"D4",X"53",X"52",X"B2",X"00",
		X"F7",X"C4",X"52",X"52",X"9B",X"36",X"D2",X"4F",X"C1",X"43",X"52",X"52",X"B8",X"00",X"D1",X"27",
		X"C3",X"52",X"52",X"FE",X"35",X"F1",X"20",X"C1",X"52",X"52",X"C2",X"00",X"D1",X"37",X"D2",X"52",
		X"CD",X"00",X"F1",X"30",X"C4",X"64",X"52",X"F6",X"00",X"D2",X"6F",X"C1",X"43",X"64",X"52",X"02",
		X"0B",X"D1",X"07",X"C3",X"64",X"52",X"6B",X"37",X"F1",X"00",X"C1",X"64",X"52",X"6D",X"12",X"D1",
		X"17",X"E4",X"52",X"20",X"01",X"F1",X"10",X"E6",X"54",X"45",X"52",X"13",X"17",X"D2",X"45",X"E1",
		X"54",X"45",X"52",X"22",X"12",X"D2",X"65",X"D4",X"45",X"52",X"6C",X"32",X"D7",X"E1",X"C5",X"65",
		X"55",X"53",X"45",X"52",X"01",X"01",X"8D",X"C5",X"56",X"52",X"45",X"53",X"45",X"52",X"33",X"36",
		X"8C",X"01",X"D3",X"45",X"52",X"7A",X"12",X"F0",X"80",X"D4",X"41",X"45",X"50",X"45",X"52",X"40",
		X"01",X"A7",X"D2",X"27",X"01",X"DB",X"E0",X"53",X"55",X"50",X"EC",X"0A",X"F6",X"C5",X"D0",X"67",
		X"50",X"C4",X"37",X"F6",X"C1",X"E7",X"50",X"17",X"34",X"DA",X"08",X"C5",X"50",X"AB",X"32",X"DA",
		X"28",X"C5",X"47",X"41",X"50",X"70",X"14",X"A0",X"30",X"D0",X"4B",X"01",X"DA",X"18",X"E1",X"54",
		X"55",X"67",X"0F",X"0A",X"D2",X"8B",X"C4",X"54",X"55",X"67",X"26",X"0A",X"D2",X"AB",X"D4",X"55",
		X"67",X"A4",X"01",X"C9",X"41",X"D2",X"61",X"54",X"67",X"74",X"01",X"D2",X"9B",X"D2",X"44",X"54",
		X"67",X"7C",X"01",X"D2",X"BB",X"C7",X"52",X"67",X"85",X"0C",X"81",X"D2",X"67",X"E5",X"0B",X"F2",
		X"98",X"F2",X"66",X"9C",X"10",X"DA",X"00",X"D0",X"67",X"66",X"02",X"0A",X"D1",X"00",X"D4",X"53",
		X"61",X"64",X"67",X"66",X"42",X"0A",X"87",X"C7",X"45",X"66",X"E6",X"31",X"D2",X"44",X"D2",X"60",
		X"43",X"66",X"23",X"32",X"B4",X"C3",X"66",X"2C",X"34",X"DA",X"10",X"C5",X"65",X"41",X"66",X"C0",
		X"36",X"AB",X"C4",X"67",X"65",X"7D",X"33",X"B5",X"C7",X"45",X"65",X"EF",X"35",X"96",X"D8",X"C5",
		X"65",X"A3",X"17",X"96",X"FF",X"E7",X"52",X"43",X"41",X"65",X"1A",X"33",X"91",X"E5",X"DD",X"16",
		X"DA",X"38",X"E7",X"64",X"42",X"16",X"B1",X"D4",X"53",X"61",X"64",X"D9",X"11",X"86",X"D2",X"61",
		X"44",X"64",X"9C",X"15",X"D2",X"98",X"E1",X"44",X"64",X"54",X"12",X"D2",X"88",X"D2",X"44",X"44",
		X"64",X"DF",X"15",X"D2",X"B8",X"C4",X"44",X"64",X"5B",X"15",X"D2",X"A8",X"C4",X"64",X"14",X"02",
		X"D0",X"E4",X"33",X"02",X"DD",X"05",X"D2",X"62",X"4E",X"16",X"D3",X"30",X"D0",X"62",X"1C",X"02",
		X"D5",X"C3",X"F1",X"61",X"18",X"02",X"FC",X"08",X"F0",X"61",X"A1",X"0A",X"FD",X"08",X"C5",X"47");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
