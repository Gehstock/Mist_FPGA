library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity gravitar_vec_rom3 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of gravitar_vec_rom3 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"EC",X"EF",X"40",X"80",X"84",X"64",X"2C",X"00",X"82",X"1D",X"3A",X"46",X"26",X"4D",X"2D",X"46",
		X"26",X"5A",X"26",X"46",X"2D",X"5A",X"26",X"53",X"3A",X"5A",X"26",X"5A",X"3A",X"53",X"33",X"5A",
		X"3A",X"46",X"3A",X"5A",X"33",X"46",X"3A",X"4D",X"26",X"46",X"00",X"C0",X"D4",X"64",X"34",X"40",
		X"26",X"00",X"18",X"00",X"38",X"48",X"F0",X"1F",X"36",X"00",X"20",X"4C",X"E8",X"1F",X"26",X"00",
		X"28",X"48",X"CA",X"1F",X"F0",X"1F",X"2C",X"40",X"DA",X"1F",X"E8",X"1F",X"28",X"58",X"10",X"00",
		X"CA",X"1F",X"20",X"54",X"18",X"00",X"DA",X"1F",X"38",X"58",X"00",X"C0",X"D4",X"64",X"00",X"00",
		X"D0",X"3F",X"26",X"00",X"30",X"00",X"20",X"00",X"E0",X"3F",X"E0",X"1F",X"46",X"00",X"30",X"00",
		X"00",X"20",X"D0",X"1F",X"26",X"00",X"20",X"00",X"20",X"20",X"BA",X"1F",X"E0",X"1F",X"00",X"00",
		X"30",X"20",X"DA",X"1F",X"D0",X"1F",X"E0",X"1F",X"20",X"20",X"1E",X"00",X"BA",X"1F",X"D0",X"1F",
		X"00",X"20",X"30",X"00",X"DA",X"1F",X"31",X"51",X"00",X"C0",X"D4",X"64",X"00",X"00",X"B2",X"DF",
		X"26",X"00",X"4E",X"00",X"34",X"00",X"CC",X"3F",X"CC",X"1F",X"5A",X"00",X"4E",X"00",X"00",X"20",
		X"B2",X"1F",X"26",X"00",X"34",X"00",X"34",X"20",X"A6",X"1F",X"CC",X"1F",X"00",X"00",X"4E",X"20",
		X"DA",X"1F",X"B2",X"1F",X"CC",X"1F",X"34",X"20",X"34",X"00",X"A6",X"1F",X"B2",X"1F",X"00",X"20",
		X"4E",X"00",X"DA",X"1F",X"CC",X"1F",X"CC",X"3F",X"00",X"C0",X"01",X"B0",X"16",X"F0",X"01",X"B0",
		X"2E",X"F0",X"01",X"B0",X"4D",X"F0",X"40",X"80",X"84",X"64",X"C2",X"01",X"38",X"02",X"05",X"F0",
		X"73",X"B0",X"16",X"F0",X"73",X"B0",X"2E",X"F0",X"73",X"B0",X"4D",X"F0",X"40",X"80",X"97",X"64",
		X"9C",X"1F",X"58",X"02",X"88",X"48",X"88",X"44",X"88",X"42",X"88",X"5E",X"88",X"5C",X"88",X"58",
		X"98",X"58",X"98",X"5C",X"98",X"5E",X"98",X"42",X"98",X"44",X"98",X"48",X"00",X"C0",X"77",X"64",
		X"8C",X"56",X"88",X"5E",X"88",X"42",X"8C",X"4A",X"84",X"40",X"00",X"C0",X"84",X"64",X"84",X"40",
		X"8C",X"4A",X"88",X"42",X"88",X"5E",X"8C",X"56",X"84",X"40",X"00",X"00",X"D0",X"1F",X"E0",X"5E",
		X"1A",X"40",X"C0",X"44",X"C4",X"44",X"C0",X"44",X"C4",X"5C",X"C0",X"5C",X"DC",X"5C",X"DC",X"40",
		X"DC",X"44",X"DA",X"42",X"DC",X"5C",X"00",X"44",X"C4",X"44",X"C6",X"5E",X"0C",X"40",X"C6",X"42",
		X"C4",X"5C",X"00",X"5C",X"DC",X"44",X"DA",X"5E",X"00",X"C0",X"7E",X"B0",X"96",X"F0",X"7E",X"B0",
		X"8F",X"F0",X"40",X"80",X"75",X"64",X"38",X"1F",X"88",X"1D",X"20",X"00",X"10",X"80",X"10",X"00",
		X"20",X"80",X"F0",X"1F",X"20",X"80",X"E0",X"1F",X"10",X"80",X"E0",X"1F",X"F0",X"9F",X"F0",X"1F",
		X"E0",X"9F",X"10",X"00",X"E0",X"9F",X"20",X"00",X"F0",X"9F",X"0C",X"40",X"C4",X"48",X"B8",X"48",
		X"08",X"58",X"C8",X"44",X"C8",X"5C",X"A8",X"48",X"18",X"58",X"C4",X"58",X"DC",X"58",X"A8",X"58",
		X"18",X"48",X"D8",X"5C",X"D8",X"44",X"B8",X"58",X"08",X"48",X"DC",X"48",X"74",X"64",X"1C",X"40",
		X"E2",X"40",X"06",X"40",X"E2",X"40",X"06",X"40",X"E0",X"42",X"1E",X"44",X"FE",X"40",X"1C",X"42",
		X"FE",X"40",X"1C",X"5E",X"E0",X"5E",X"00",X"56",X"E2",X"40",X"04",X"5E",X"E2",X"40",X"04",X"42",
		X"E0",X"42",X"1C",X"42",X"E0",X"42",X"00",X"42",X"E2",X"40",X"02",X"40",X"E0",X"5E",X"00",X"5E",
		X"E2",X"40",X"00",X"C0",X"84",X"64",X"20",X"41",X"3F",X"41",X"3F",X"40",X"3F",X"5F",X"20",X"5F",
		X"21",X"5F",X"21",X"40",X"21",X"41",X"00",X"C0",X"40",X"80",X"A2",X"64",X"DA",X"1D",X"14",X"00",
		X"34",X"B2",X"0A",X"F1",X"66",X"64",X"03",X"46",X"35",X"42",X"E0",X"1F",X"50",X"20",X"37",X"46",
		X"23",X"5D",X"16",X"00",X"CA",X"3F",X"24",X"40",X"00",X"C0",X"04",X"B1",X"04",X"48",X"FA",X"F0",
		X"04",X"F1",X"04",X"B1",X"10",X"00",X"28",X"00",X"FA",X"F0",X"04",X"B1",X"0C",X"48",X"FA",X"F0",
		X"3C",X"41",X"22",X"46",X"29",X"5E",X"3D",X"55",X"31",X"44",X"20",X"00",X"0A",X"20",X"F4",X"1F",
		X"2A",X"20",X"D4",X"1F",X"F4",X"3F",X"10",X"00",X"C8",X"3F",X"38",X"00",X"10",X"20",X"EC",X"1F",
		X"44",X"20",X"BC",X"1F",X"EE",X"3F",X"16",X"00",X"AC",X"3F",X"52",X"00",X"18",X"20",X"00",X"C0",
		X"21",X"5C",X"3A",X"5E",X"3D",X"4A",X"2B",X"43",X"E0",X"1F",X"0A",X"20",X"F6",X"1F",X"E0",X"3F",
		X"2C",X"00",X"F2",X"3F",X"0E",X"00",X"2C",X"20",X"C8",X"1F",X"12",X"20",X"EE",X"1F",X"C8",X"3F",
		X"44",X"00",X"EA",X"3F",X"16",X"00",X"46",X"20",X"B0",X"1F",X"1A",X"20",X"E4",X"1F",X"AE",X"3F",
		X"00",X"C0",X"24",X"44",X"24",X"5C",X"38",X"58",X"38",X"48",X"2C",X"4C",X"2C",X"54",X"E0",X"1F",
		X"E0",X"3F",X"20",X"00",X"E0",X"3F",X"28",X"00",X"28",X"20",X"D8",X"1F",X"28",X"20",X"D0",X"1F",
		X"D0",X"3F",X"30",X"00",X"D0",X"3F",X"38",X"00",X"38",X"20",X"C8",X"1F",X"38",X"20",X"00",X"C0",
		X"40",X"80",X"C6",X"64",X"C2",X"01",X"CE",X"1F",X"20",X"F1",X"40",X"80",X"C6",X"64",X"C2",X"01",
		X"CE",X"1F",X"38",X"F1",X"40",X"80",X"C6",X"64",X"C2",X"01",X"CE",X"1F",X"51",X"F1",X"61",X"64",
		X"C2",X"01",X"4C",X"1E",X"24",X"42",X"00",X"00",X"40",X"20",X"24",X"5E",X"3C",X"5E",X"00",X"00",
		X"C0",X"3F",X"3C",X"42",X"00",X"C0",X"C7",X"64",X"28",X"00",X"14",X"00",X"24",X"58",X"20",X"44",
		X"E0",X"1F",X"10",X"20",X"20",X"44",X"E0",X"1F",X"10",X"20",X"20",X"58",X"20",X"00",X"F0",X"3F",
		X"20",X"5C",X"E0",X"1F",X"10",X"20",X"20",X"5C",X"3C",X"48",X"20",X"48",X"D8",X"1F",X"EC",X"1F",
		X"00",X"C0",X"C7",X"64",X"60",X"00",X"20",X"00",X"20",X"58",X"3C",X"58",X"20",X"44",X"E0",X"1F",
		X"F0",X"3F",X"20",X"44",X"E0",X"1F",X"F0",X"3F",X"20",X"48",X"20",X"00",X"10",X"20",X"20",X"5C",
		X"20",X"00",X"10",X"20",X"20",X"5C",X"24",X"48",X"D8",X"1F",X"C4",X"1F",X"00",X"C0",X"61",X"64",
		X"C2",X"01",X"4C",X"1E",X"28",X"00",X"28",X"00",X"22",X"5C",X"C0",X"1F",X"00",X"20",X"3E",X"5C",
		X"3E",X"44",X"40",X"00",X"00",X"20",X"22",X"44",X"00",X"C0",X"C7",X"64",X"EC",X"1F",X"28",X"00",
		X"38",X"5C",X"24",X"40",X"F0",X"1F",X"E0",X"1F",X"24",X"40",X"F0",X"1F",X"E0",X"3F",X"38",X"40",
		X"10",X"00",X"20",X"20",X"3C",X"40",X"10",X"00",X"20",X"20",X"3C",X"40",X"28",X"44",X"28",X"40",
		X"14",X"00",X"D8",X"1F",X"00",X"C0",X"C7",X"64",X"C4",X"1F",X"28",X"00",X"38",X"40",X"38",X"44",
		X"24",X"40",X"10",X"00",X"E0",X"3F",X"3C",X"40",X"10",X"00",X"E0",X"3F",X"28",X"40",X"F0",X"1F",
		X"20",X"20",X"3C",X"40",X"F0",X"1F",X"20",X"20",X"3C",X"40",X"28",X"5C",X"14",X"00",X"B0",X"1F",
		X"00",X"C0",X"40",X"80",X"78",X"F1",X"40",X"80",X"78",X"B1",X"83",X"F1",X"40",X"80",X"78",X"B1",
		X"83",X"B1",X"99",X"F1",X"40",X"80",X"AF",X"F1",X"40",X"80",X"AF",X"B1",X"BD",X"F1",X"40",X"80",
		X"AF",X"B1",X"BD",X"B1",X"D3",X"F1",X"40",X"80",X"A3",X"64",X"70",X"1E",X"40",X"02",X"E4",X"1F",
		X"54",X"20",X"E4",X"1F",X"AC",X"3F",X"48",X"00",X"34",X"20",X"A8",X"1F",X"00",X"20",X"48",X"00",
		X"CC",X"3F",X"07",X"5B",X"EE",X"1F",X"38",X"20",X"EC",X"1F",X"C6",X"3F",X"32",X"00",X"26",X"20",
		X"C4",X"1F",X"00",X"20",X"30",X"00",X"DE",X"3F",X"00",X"C0",X"40",X"80",X"A3",X"64",X"70",X"1E",
		X"40",X"02",X"04",X"45",X"D6",X"1F",X"4A",X"20",X"00",X"00",X"A8",X"3F",X"34",X"00",X"46",X"20",
		X"AA",X"1F",X"E6",X"3F",X"4C",X"00",X"E2",X"3F",X"05",X"5E",X"DE",X"1F",X"32",X"20",X"00",X"00",
		X"C4",X"3F",X"24",X"00",X"30",X"20",X"C6",X"1F",X"EE",X"3F",X"38",X"00",X"EC",X"3F",X"00",X"C0",
		X"40",X"80",X"BC",X"1D",X"8E",X"1D",X"82",X"64",X"24",X"48",X"28",X"44",X"28",X"5C",X"24",X"58",
		X"3C",X"58",X"38",X"5C",X"38",X"44",X"3C",X"48",X"00",X"C0",X"84",X"64",X"0A",X"4B",X"3D",X"44",
		X"39",X"42",X"38",X"41",X"28",X"40",X"2A",X"5D",X"24",X"5C",X"D4",X"1F",X"F8",X"1F",X"24",X"5C",
		X"2A",X"5D",X"28",X"40",X"38",X"41",X"39",X"42",X"3D",X"44",X"12",X"4B",X"00",X"C0",X"87",X"64",
		X"18",X"55",X"28",X"4C",X"2C",X"46",X"20",X"48",X"2C",X"46",X"28",X"41",X"00",X"C0",X"84",X"64",
		X"0A",X"4B",X"24",X"44",X"2A",X"43",X"28",X"40",X"38",X"5F",X"39",X"5E",X"3D",X"5C",X"D4",X"1F",
		X"F8",X"1F",X"3D",X"5C",X"39",X"5E",X"38",X"5F",X"28",X"40",X"2A",X"43",X"24",X"44",X"12",X"4B",
		X"00",X"C0",X"87",X"64",X"18",X"4B",X"28",X"5F",X"2C",X"5A",X"20",X"58",X"2C",X"5A",X"28",X"5F",
		X"00",X"C0",X"30",X"B2",X"3D",X"B2",X"4F",X"F2",X"30",X"B2",X"57",X"B2",X"69",X"F2",X"85",X"64",
		X"20",X"00",X"20",X"20",X"00",X"00",X"20",X"20",X"E0",X"1F",X"20",X"20",X"E0",X"1F",X"00",X"20",
		X"E0",X"1F",X"E0",X"3F",X"00",X"00",X"E0",X"3F",X"20",X"00",X"E0",X"3F",X"20",X"00",X"00",X"20",
		X"00",X"C0",X"A1",X"64",X"08",X"5E",X"2A",X"4A",X"2C",X"40",X"2A",X"56",X"20",X"54",X"36",X"56",
		X"34",X"40",X"36",X"4A",X"20",X"4C",X"18",X"42",X"00",X"C0",X"C4",X"64",X"0E",X"5B",X"25",X"45",
		X"26",X"40",X"25",X"5B",X"20",X"5A",X"3B",X"5B",X"3A",X"40",X"3B",X"45",X"20",X"46",X"00",X"C0",
		X"40",X"80",X"F4",X"01",X"1A",X"02",X"77",X"F2",X"40",X"80",X"F4",X"01",X"1A",X"02",X"77",X"B2",
		X"89",X"F2",X"40",X"80",X"F4",X"01",X"1A",X"02",X"77",X"B2",X"89",X"B2",X"95",X"F2",X"C4",X"64",
		X"C9",X"43",X"C3",X"5D",X"D4",X"5A",X"D4",X"46",X"C3",X"43",X"C9",X"5D",X"A6",X"64",X"C3",X"40",
		X"DD",X"46",X"DD",X"5A",X"C3",X"40",X"00",X"C0",X"C4",X"64",X"14",X"40",X"CC",X"46",X"CC",X"5A",
		X"DA",X"5A",X"D4",X"40",X"DA",X"46",X"A7",X"64",X"02",X"5E",X"00",X"00",X"28",X"20",X"00",X"43",
		X"00",X"00",X"D8",X"3F",X"00",X"C0",X"C4",X"64",X"24",X"42",X"28",X"58",X"3D",X"5D",X"3D",X"40",
		X"23",X"43",X"3D",X"43",X"34",X"40",X"3D",X"5D",X"23",X"5D",X"3D",X"40",X"3D",X"43",X"28",X"48",
		X"24",X"5E",X"00",X"C0",X"00",X"4A",X"FB",X"40",X"FB",X"56",X"E5",X"56",X"EA",X"40",X"E5",X"4A",
		X"FB",X"4A",X"FB",X"40",X"00",X"C0",X"03",X"B3",X"13",X"B3",X"23",X"B3",X"35",X"B3",X"46",X"B3",
		X"56",X"B3",X"65",X"B3",X"77",X"B3",X"87",X"B3",X"97",X"B3",X"A7",X"B3",X"B9",X"B3",X"CA",X"B3",
		X"DA",X"B3",X"E9",X"B3",X"FB",X"B3",X"0B",X"B4",X"1B",X"B4",X"2B",X"B4",X"3D",X"B4",X"4E",X"B4",
		X"5E",X"B4",X"6D",X"B4",X"7F",X"B4",X"8F",X"B4",X"9F",X"B4",X"AF",X"B4",X"C1",X"B4",X"D2",X"B4",
		X"E2",X"B4",X"F1",X"B4",X"03",X"B5",X"00",X"49",X"E9",X"1F",X"0D",X"C0",X"F7",X"1F",X"FB",X"DF",
		X"DE",X"40",X"07",X"00",X"FC",X"DF",X"F9",X"1F",X"FC",X"DF",X"DE",X"40",X"09",X"00",X"FB",X"DF",
		X"17",X"00",X"0D",X"C0",X"00",X"C0",X"02",X"49",X"E7",X"1F",X"08",X"C0",X"F8",X"1F",X"F9",X"DF",
		X"01",X"00",X"FC",X"DF",X"07",X"00",X"FE",X"DF",X"DD",X"5D",X"01",X"00",X"FC",X"DF",X"0A",X"00",
		X"FD",X"DF",X"C9",X"4A",X"00",X"C0",X"11",X"00",X"07",X"00",X"E6",X"1F",X"03",X"C0",X"F9",X"1F",
		X"F8",X"DF",X"DE",X"41",X"08",X"00",X"FF",X"DF",X"FB",X"1F",X"FA",X"DF",X"01",X"00",X"FC",X"DF",
		X"0A",X"00",X"FF",X"DF",X"11",X"00",X"15",X"C0",X"00",X"C0",X"0F",X"00",X"0A",X"00",X"DF",X"53",
		X"FB",X"1F",X"F7",X"DF",X"02",X"00",X"FD",X"DF",X"C0",X"44",X"FD",X"1F",X"F9",X"DF",X"02",X"00",
		X"FD",X"DF",X"0A",X"00",X"01",X"C0",X"0C",X"00",X"17",X"C0",X"00",X"C0",X"0D",X"00",X"0D",X"00",
		X"E6",X"1F",X"F9",X"DF",X"DB",X"5F",X"03",X"00",X"FD",X"DF",X"C1",X"44",X"DC",X"5F",X"03",X"00",
		X"FD",X"DF",X"0A",X"00",X"03",X"C0",X"07",X"00",X"1A",X"C0",X"00",X"C0",X"0A",X"00",X"0F",X"00",
		X"DA",X"54",X"FF",X"1F",X"F6",X"DF",X"DF",X"42",X"07",X"00",X"03",X"C0",X"FF",X"1F",X"F8",X"DF",
		X"DF",X"42",X"09",X"00",X"05",X"C0",X"CD",X"41",X"00",X"C0",X"07",X"00",X"10",X"00",X"EB",X"1F",
		X"F1",X"DF",X"01",X"00",X"F5",X"DF",X"04",X"00",X"FF",X"DF",X"06",X"00",X"05",X"C0",X"01",X"00",
		X"F7",X"DF",X"04",X"00",X"FF",X"DF",X"C3",X"44",X"FD",X"1F",X"1A",X"C0",X"00",X"C0",X"09",X"42",
		X"D6",X"57",X"03",X"00",X"F6",X"DF",X"04",X"00",X"FF",X"DF",X"05",X"00",X"06",X"C0",X"03",X"00",
		X"F9",X"DF",X"04",X"00",X"FF",X"DF",X"07",X"00",X"07",X"C0",X"CD",X"5C",X"00",X"C0",X"09",X"40",
		X"F3",X"1F",X"E9",X"DF",X"05",X"00",X"F7",X"DF",X"C0",X"42",X"04",X"00",X"07",X"C0",X"04",X"00",
		X"F9",X"DF",X"C0",X"42",X"05",X"00",X"09",X"C0",X"F3",X"1F",X"17",X"C0",X"00",X"C0",X"09",X"5E",
		X"F8",X"1F",X"E7",X"DF",X"07",X"00",X"F8",X"DF",X"04",X"00",X"01",X"C0",X"02",X"00",X"07",X"C0",
		X"DD",X"43",X"04",X"00",X"01",X"C0",X"03",X"00",X"0A",X"C0",X"CA",X"57",X"00",X"C0",X"F9",X"1F",
		X"11",X"00",X"FD",X"1F",X"E6",X"DF",X"08",X"00",X"F9",X"DF",X"C1",X"42",X"01",X"00",X"08",X"C0",
		X"06",X"00",X"FB",X"DF",X"04",X"00",X"01",X"C0",X"01",X"00",X"0A",X"C0",X"EB",X"1F",X"11",X"C0",
		X"00",X"C0",X"F6",X"1F",X"0F",X"00",X"D3",X"41",X"09",X"00",X"FB",X"DF",X"03",X"00",X"02",X"C0",
		X"C4",X"40",X"07",X"00",X"FD",X"DF",X"03",X"00",X"02",X"C0",X"FF",X"1F",X"0A",X"C0",X"E9",X"1F",
		X"0C",X"C0",X"00",X"C0",X"F3",X"1F",X"0D",X"00",X"07",X"00",X"E6",X"DF",X"DF",X"45",X"03",X"00",
		X"03",X"C0",X"C4",X"5F",X"DF",X"44",X"03",X"00",X"03",X"C0",X"FD",X"1F",X"0A",X"C0",X"E6",X"1F",
		X"07",X"C0",X"00",X"C0",X"F1",X"1F",X"0A",X"00",X"D4",X"46",X"0A",X"00",X"FF",X"DF",X"C2",X"41",
		X"FD",X"1F",X"07",X"C0",X"08",X"00",X"FF",X"DF",X"C2",X"41",X"FB",X"1F",X"09",X"C0",X"C1",X"53",
		X"00",X"C0",X"F0",X"1F",X"07",X"00",X"0F",X"00",X"EB",X"DF",X"0B",X"00",X"01",X"C0",X"01",X"00",
		X"04",X"C0",X"FB",X"1F",X"06",X"C0",X"09",X"00",X"01",X"C0",X"01",X"00",X"04",X"C0",X"C4",X"5D",
		X"E6",X"1F",X"FD",X"DF",X"00",X"C0",X"02",X"57",X"D7",X"4A",X"0A",X"00",X"03",X"C0",X"01",X"00",
		X"04",X"C0",X"FA",X"1F",X"05",X"C0",X"07",X"00",X"03",X"C0",X"01",X"00",X"04",X"C0",X"F9",X"1F",
		X"07",X"C0",X"DC",X"53",X"00",X"C0",X"00",X"57",X"17",X"00",X"F3",X"DF",X"09",X"00",X"05",X"C0",
		X"C2",X"40",X"F9",X"1F",X"04",X"C0",X"07",X"00",X"04",X"C0",X"C2",X"40",X"F7",X"1F",X"05",X"C0",
		X"E9",X"1F",X"F3",X"DF",X"00",X"C0",X"1E",X"57",X"19",X"00",X"F8",X"DF",X"08",X"00",X"07",X"C0",
		X"FF",X"1F",X"04",X"C0",X"F9",X"1F",X"02",X"C0",X"C3",X"43",X"FF",X"1F",X"04",X"C0",X"F6",X"1F",
		X"03",X"C0",X"D7",X"56",X"00",X"C0",X"EF",X"1F",X"F9",X"1F",X"1A",X"00",X"FD",X"DF",X"07",X"00",
		X"08",X"C0",X"C2",X"5F",X"F8",X"1F",X"01",X"C0",X"05",X"00",X"06",X"C0",X"FF",X"1F",X"04",X"C0",
		X"F6",X"1F",X"01",X"C0",X"EF",X"1F",X"EB",X"DF",X"00",X"C0",X"F1",X"1F",X"F6",X"1F",X"C1",X"4D",
		X"05",X"00",X"09",X"C0",X"FE",X"1F",X"03",X"C0",X"C0",X"5C",X"03",X"00",X"07",X"C0",X"FE",X"1F",
		X"03",X"C0",X"F6",X"1F",X"FF",X"DF",X"F4",X"1F",X"E9",X"DF",X"00",X"C0",X"F3",X"1F",X"F3",X"1F",
		X"1A",X"00",X"07",X"C0",X"C5",X"41",X"FD",X"1F",X"03",X"C0",X"DF",X"5C",X"C4",X"41",X"FD",X"1F",
		X"03",X"C0",X"F6",X"1F",X"FD",X"DF",X"F9",X"1F",X"E6",X"DF",X"00",X"C0",X"F6",X"1F",X"F1",X"1F",
		X"C6",X"4C",X"01",X"00",X"0A",X"C0",X"C1",X"5E",X"F9",X"1F",X"FD",X"DF",X"01",X"00",X"08",X"C0",
		X"C1",X"5E",X"F7",X"1F",X"FB",X"DF",X"D3",X"5F",X"00",X"C0",X"F9",X"1F",X"F0",X"1F",X"15",X"00",
		X"0F",X"C0",X"FF",X"1F",X"0B",X"C0",X"FC",X"1F",X"01",X"C0",X"FA",X"1F",X"FB",X"DF",X"FF",X"1F",
		X"09",X"C0",X"FC",X"1F",X"01",X"C0",X"DD",X"5C",X"03",X"00",X"E6",X"DF",X"00",X"C0",X"17",X"5E",
		X"CA",X"49",X"FD",X"1F",X"0A",X"C0",X"FC",X"1F",X"01",X"C0",X"FB",X"1F",X"FA",X"DF",X"FD",X"1F",
		X"07",X"C0",X"FC",X"1F",X"01",X"C0",X"F9",X"1F",X"F9",X"DF",X"D3",X"44",X"00",X"C0",X"17",X"40",
		X"0D",X"00",X"17",X"C0",X"FB",X"1F",X"09",X"C0",X"C0",X"5E",X"FC",X"1F",X"F9",X"DF",X"FC",X"1F",
		X"07",X"C0",X"C0",X"5E",X"FB",X"1F",X"F7",X"DF",X"0D",X"00",X"E9",X"DF",X"00",X"C0",X"17",X"42",
		X"08",X"00",X"19",X"C0",X"F9",X"1F",X"08",X"C0",X"FC",X"1F",X"FF",X"DF",X"FE",X"1F",X"F9",X"DF",
		X"C3",X"5D",X"FC",X"1F",X"FF",X"DF",X"FD",X"1F",X"F6",X"DF",X"D6",X"49",X"00",X"C0",X"07",X"00",
		X"EF",X"1F",X"03",X"00",X"1A",X"C0",X"F8",X"1F",X"07",X"C0",X"DF",X"5E",X"FF",X"1F",X"F8",X"DF",
		X"FA",X"1F",X"05",X"C0",X"FC",X"1F",X"FF",X"DF",X"01",X"00",X"F6",X"DF",X"15",X"00",X"EF",X"DF",
		X"00",X"C0",X"0A",X"00",X"F1",X"1F",X"CD",X"5F",X"F7",X"1F",X"05",X"C0",X"FD",X"1F",X"FE",X"DF",
		X"DC",X"40",X"F9",X"1F",X"03",X"C0",X"FD",X"1F",X"FE",X"DF",X"01",X"00",X"F6",X"DF",X"17",X"00",
		X"F4",X"DF",X"00",X"C0",X"0D",X"00",X"F3",X"1F",X"F9",X"1F",X"1A",X"C0",X"C1",X"5B",X"FD",X"1F",
		X"FD",X"DF",X"DC",X"41",X"C1",X"5C",X"FD",X"1F",X"FD",X"DF",X"03",X"00",X"F6",X"DF",X"1A",X"00",
		X"F9",X"DF",X"00",X"C0",X"0F",X"00",X"F6",X"1F",X"CC",X"5A",X"F6",X"1F",X"01",X"C0",X"DE",X"5F",
		X"03",X"00",X"F9",X"DF",X"F8",X"1F",X"01",X"C0",X"DE",X"5F",X"05",X"00",X"F7",X"DF",X"DF",X"4D",
		X"00",X"C0",X"10",X"00",X"F9",X"1F",X"F1",X"1F",X"15",X"C0",X"F5",X"1F",X"FF",X"DF",X"FF",X"1F",
		X"FC",X"DF",X"05",X"00",X"FA",X"DF",X"F7",X"1F",X"FF",X"DF",X"FF",X"1F",X"FC",X"DF",X"DC",X"43",
		X"1A",X"00",X"03",X"C0",X"00",X"C0",X"1E",X"49",X"C9",X"56",X"F6",X"1F",X"FD",X"DF",X"FF",X"1F",
		X"FC",X"DF",X"06",X"00",X"FB",X"DF",X"F9",X"1F",X"FD",X"DF",X"FF",X"1F",X"FC",X"DF",X"07",X"00",
		X"F9",X"DF",X"C4",X"4D",X"00",X"C0",X"B0",X"3A",X"C2",X"3A",X"D4",X"3A",X"E2",X"3A",X"F4",X"3A",
		X"04",X"3B",X"14",X"3B",X"26",X"3B",X"38",X"3B",X"4A",X"3B",X"5C",X"3B",X"6A",X"3B",X"7C",X"3B",
		X"8C",X"3B",X"9C",X"3B",X"AE",X"3B",X"C0",X"3B",X"D2",X"3B",X"E4",X"3B",X"F2",X"3B",X"04",X"3C",
		X"14",X"3C",X"24",X"3C",X"36",X"3C",X"48",X"3C",X"5A",X"3C",X"6C",X"3C",X"7A",X"3C",X"8C",X"3C",
		X"9C",X"3C",X"AC",X"3C",X"BE",X"3C",X"D0",X"3C",X"DE",X"3C",X"94",X"4D",X"DA",X"4D",X"3A",X"4E",
		X"92",X"4E",X"D2",X"4E",X"F6",X"4E",X"2A",X"4F",X"82",X"4F",X"5E",X"45",X"78",X"45",X"96",X"45",
		X"96",X"45",X"40",X"80",X"00",X"73",X"00",X"C0",X"40",X"80",X"00",X"71",X"00",X"C0",X"44",X"B5",
		X"81",X"1E",X"60",X"1E",X"00",X"00",X"40",X"23",X"FF",X"02",X"00",X"20",X"00",X"00",X"C0",X"3C",
		X"01",X"1D",X"00",X"20",X"00",X"C0",X"80",X"1E",X"60",X"1E",X"FF",X"02",X"FF",X"82",X"C1",X"1F",
		X"3F",X"80",X"40",X"1D",X"40",X"9D",X"80",X"00",X"80",X"9F",X"80",X"02",X"80",X"82",X"40",X"1F",
		X"C0",X"80",X"C0",X"1D",X"C0",X"9D",X"FF",X"00",X"01",X"9F",X"FF",X"01",X"FF",X"81",X"C2",X"1E",
		X"3E",X"81",X"40",X"1E",X"40",X"9E",X"7F",X"01",X"81",X"9E",X"7F",X"01",X"7F",X"81",X"40",X"1E",
		X"C0",X"81",X"C2",X"1E",X"C2",X"9E",X"FF",X"01",X"01",X"9E",X"FF",X"00",X"FF",X"80",X"C0",X"1D",
		X"40",X"82",X"40",X"1F",X"40",X"9F",X"80",X"02",X"80",X"9D",X"80",X"00",X"80",X"80",X"40",X"1D",
		X"C0",X"82",X"C1",X"1F",X"C1",X"9F",X"FF",X"02",X"01",X"9D",X"01",X"1E",X"00",X"00",X"14",X"71",
		X"A4",X"F6",X"10",X"00",X"00",X"1F",X"00",X"C0",X"00",X"00",X"00",X"E1",X"89",X"B5",X"00",X"00",
		X"00",X"C1",X"89",X"B5",X"00",X"00",X"00",X"A1",X"89",X"B5",X"00",X"00",X"00",X"81",X"89",X"B5",
		X"00",X"00",X"00",X"61",X"89",X"B5",X"00",X"00",X"00",X"41",X"00",X"C0",X"17",X"64",X"00",X"00",
		X"40",X"40",X"10",X"00",X"C0",X"1E",X"00",X"00",X"00",X"21",X"00",X"C0",X"01",X"1D",X"00",X"20",
		X"40",X"80",X"00",X"C0",X"00",X"00",X"40",X"23",X"40",X"80",X"00",X"C0",X"C7",X"64",X"40",X"80",
		X"53",X"F5",X"C8",X"B5",X"00",X"70",X"C0",X"00",X"00",X"00",X"C8",X"B5",X"25",X"40",X"C8",X"B5",
		X"40",X"1F",X"00",X"00",X"C8",X"B5",X"25",X"40",X"C8",X"B5",X"00",X"00",X"00",X"01",X"C8",X"B5",
		X"20",X"45",X"C8",X"B5",X"00",X"00",X"00",X"1F",X"C8",X"B5",X"20",X"45",X"40",X"80",X"00",X"C0",
		X"87",X"64",X"40",X"80",X"40",X"80",X"00",X"C0",X"44",X"B5",X"D4",X"1E",X"D4",X"1E",X"00",X"60",
		X"58",X"02",X"58",X"02",X"00",X"C0",X"40",X"80",X"00",X"70",X"01",X"1F",X"01",X"1F",X"00",X"00",
		X"FF",X"01",X"00",X"00",X"01",X"1E",X"00",X"00",X"FF",X"01",X"00",X"00",X"01",X"1E",X"40",X"80",
		X"00",X"C0",X"00",X"00",X"40",X"23",X"00",X"5F",X"00",X"00",X"C0",X"3C",X"00",X"C0",X"40",X"80",
		X"00",X"71",X"87",X"64",X"20",X"00",X"60",X"1E",X"00",X"C0",X"80",X"48",X"84",X"44",X"84",X"5C",
		X"80",X"58",X"18",X"44",X"88",X"40",X"04",X"5C",X"00",X"C0",X"80",X"4C",X"86",X"40",X"82",X"5E",
		X"80",X"5E",X"9E",X"5E",X"9A",X"40",X"06",X"40",X"82",X"5E",X"80",X"5E",X"9E",X"5E",X"9A",X"40",
		X"3F",X"F6",X"80",X"4C",X"88",X"40",X"18",X"54",X"82",X"F6",X"80",X"4C",X"84",X"40",X"84",X"5C",
		X"80",X"5C",X"9C",X"5C",X"9C",X"40",X"3F",X"F6",X"88",X"40",X"18",X"40",X"80",X"4C",X"88",X"40",
		X"1E",X"5A",X"9A",X"40",X"0C",X"5A",X"00",X"C0",X"80",X"4C",X"88",X"40",X"80",X"5C",X"1C",X"5C",
		X"84",X"40",X"80",X"5C",X"3E",X"F6",X"80",X"4C",X"00",X"5A",X"88",X"40",X"00",X"46",X"9B",X"F6",
		X"88",X"40",X"18",X"4C",X"88",X"40",X"1C",X"40",X"80",X"54",X"08",X"40",X"00",X"C0",X"00",X"44",
		X"84",X"5C",X"84",X"40",X"60",X"F6",X"80",X"4C",X"06",X"40",X"9A",X"5A",X"86",X"5A",X"06",X"40",
		X"00",X"C0",X"00",X"4C",X"80",X"54",X"82",X"F6",X"80",X"4C",X"84",X"5C",X"84",X"44",X"9B",X"F6",
		X"80",X"4C",X"88",X"54",X"60",X"F6",X"80",X"4C",X"88",X"40",X"80",X"54",X"98",X"40",X"0C",X"40",
		X"00",X"C0",X"80",X"4C",X"88",X"40",X"80",X"5A",X"98",X"40",X"12",X"F6",X"80",X"4C",X"88",X"40",
		X"80",X"58",X"9C",X"5C",X"9C",X"40",X"04",X"44",X"84",X"5C",X"83",X"F6",X"80",X"4C",X"88",X"40",
		X"80",X"5A",X"98",X"40",X"02",X"40",X"86",X"5A",X"83",X"F6",X"88",X"40",X"80",X"46",X"98",X"40",
		X"80",X"46",X"88",X"40",X"61",X"F6",X"00",X"4C",X"22",X"F6",X"00",X"4C",X"80",X"54",X"88",X"40",
		X"80",X"4C",X"04",X"54",X"00",X"C0",X"00",X"4C",X"84",X"54",X"84",X"4C",X"61",X"F6",X"00",X"4C",
		X"80",X"54",X"84",X"44",X"84",X"5C",X"60",X"F6",X"88",X"4C",X"18",X"40",X"88",X"54",X"9C",X"F6",
		X"04",X"40",X"80",X"48",X"9C",X"44",X"08",X"40",X"9C",X"5C",X"08",X"58",X"00",X"C0",X"00",X"4C",
		X"88",X"40",X"98",X"54",X"82",X"F6",X"04",X"4C",X"24",X"F6",X"00",X"4C",X"88",X"40",X"80",X"5A",
		X"98",X"40",X"80",X"5A",X"88",X"40",X"04",X"40",X"00",X"C0",X"00",X"4C",X"88",X"40",X"80",X"54",
		X"98",X"40",X"00",X"46",X"88",X"40",X"04",X"5A",X"00",X"C0",X"00",X"4C",X"80",X"5A",X"88",X"40",
		X"00",X"46",X"9B",X"F6",X"00",X"46",X"88",X"40",X"80",X"5A",X"98",X"40",X"80",X"4C",X"0C",X"54",
		X"00",X"C0",X"00",X"4C",X"88",X"40",X"80",X"54",X"04",X"40",X"00",X"C0",X"80",X"4C",X"86",X"F6",
		X"08",X"46",X"98",X"40",X"80",X"46",X"9A",X"F6",X"3F",X"B6",X"3B",X"B6",X"7B",X"B6",X"7D",X"B6",
		X"85",X"B6",X"8D",X"B6",X"55",X"B6",X"92",X"B6",X"99",X"B6",X"9E",X"B6",X"A0",X"B6",X"ED",X"B5",
		X"F5",X"B5",X"01",X"B6",X"05",X"B6",X"0C",X"B6",X"0E",X"B6",X"14",X"B6",X"1B",X"B6",X"20",X"B6",
		X"27",X"B6",X"2B",X"B6",X"31",X"B6",X"34",X"B6",X"38",X"B6",X"3B",X"B6",X"41",X"B6",X"46",X"B6",
		X"4E",X"B6",X"55",X"B6",X"5B",X"B6",X"5D",X"B6",X"63",X"B6",X"67",X"B6",X"6C",X"B6",X"70",X"B6",
		X"77",X"B6",X"00",X"C0",X"44",X"64",X"FC",X"00",X"2F",X"9D",X"11",X"64",X"4B",X"01",X"9A",X"80",
		X"1D",X"00",X"96",X"80",X"BF",X"1F",X"E0",X"9F",X"F1",X"1F",X"AA",X"9F",X"63",X"1F",X"B0",X"9F",
		X"13",X"00",X"4E",X"80",X"2F",X"00",X"13",X"80",X"ED",X"1F",X"CE",X"9F",X"4C",X"00",X"34",X"80",
		X"0E",X"00",X"42",X"80",X"2D",X"1F",X"B9",X"9F",X"40",X"80",X"44",X"64",X"2E",X"01",X"F6",X"9D",
		X"11",X"64",X"D0",X"1F",X"36",X"9F",X"81",X"40",X"00",X"C0",X"44",X"64",X"2B",X"01",X"09",X"9E",
		X"11",X"64",X"38",X"01",X"5C",X"80",X"0F",X"00",X"3D",X"80",X"B5",X"1F",X"51",X"80",X"C2",X"1F",
		X"F2",X"9F",X"97",X"59",X"EF",X"1F",X"11",X"80",X"96",X"1F",X"E0",X"9F",X"40",X"80",X"44",X"64",
		X"3F",X"01",X"49",X"9E",X"11",X"64",X"F1",X"1F",X"C6",X"9F",X"40",X"80",X"44",X"64",X"4F",X"01",
		X"8A",X"9E",X"11",X"64",X"7D",X"00",X"18",X"80",X"93",X"40",X"36",X"00",X"09",X"80",X"01",X"00",
		X"21",X"80",X"23",X"00",X"D6",X"9F",X"1A",X"1F",X"BF",X"9F",X"40",X"80",X"44",X"64",X"5F",X"01",
		X"C5",X"9E",X"11",X"64",X"F1",X"1F",X"C6",X"9F",X"00",X"C0",X"44",X"64",X"5D",X"01",X"D5",X"9E",
		X"11",X"64",X"C9",X"00",X"30",X"80",X"4C",X"00",X"4C",X"80",X"10",X"00",X"4B",X"80",X"DE",X"1E",
		X"E6",X"9F",X"40",X"80",X"44",X"64",X"5E",X"01",X"0E",X"9F",X"11",X"64",X"FF",X"1F",X"C7",X"9F",
		X"40",X"80",X"44",X"64",X"5F",X"01",X"43",X"9F",X"11",X"64",X"D8",X"00",X"1E",X"80",X"DF",X"1F",
		X"DF",X"9F",X"00",X"00",X"11",X"80",X"C6",X"1F",X"F3",X"9F",X"00",X"00",X"DC",X"9F",X"82",X"1F",
		X"EF",X"9F",X"40",X"80",X"44",X"64",X"61",X"01",X"82",X"9F",X"11",X"64",X"FC",X"1F",X"C1",X"9F",
		X"00",X"C0",X"44",X"64",X"5E",X"01",X"C1",X"9F",X"11",X"64",X"6D",X"00",X"CE",X"9F",X"B6",X"00",
		X"0D",X"80",X"00",X"00",X"33",X"80",X"83",X"1F",X"F1",X"9F",X"C8",X"1F",X"20",X"80",X"38",X"00",
		X"20",X"80",X"7D",X"00",X"F2",X"9F",X"FF",X"1F",X"28",X"80",X"4A",X"1F",X"11",X"80",X"95",X"1F",
		X"D6",X"9F",X"40",X"80",X"44",X"64",X"5E",X"01",X"FF",X"9F",X"11",X"64",X"00",X"00",X"C0",X"9F",
		X"00",X"C0",X"44",X"64",X"60",X"01",X"3B",X"80",X"11",X"64",X"21",X"01",X"EF",X"9F",X"FF",X"1F",
		X"42",X"80",X"DF",X"1E",X"10",X"80",X"40",X"80",X"44",X"64",X"5E",X"01",X"7B",X"80",X"11",X"64",
		X"01",X"00",X"BF",X"9F",X"00",X"C0",X"44",X"64",X"5E",X"01",X"B8",X"80",X"11",X"64",X"EA",X"00",
		X"DE",X"9F",X"FF",X"1F",X"E6",X"9F",X"3A",X"00",X"F0",X"9F",X"F1",X"1F",X"8D",X"80",X"C6",X"1F",
		X"09",X"80",X"0F",X"00",X"D5",X"9F",X"18",X"1F",X"22",X"80",X"40",X"80",X"44",X"64",X"5C",X"01",
		X"F7",X"80",X"11",X"64",X"01",X"00",X"C0",X"9F",X"00",X"C0",X"44",X"64",X"5E",X"01",X"35",X"81",
		X"11",X"64",X"B7",X"00",X"DC",X"9F",X"5C",X"00",X"54",X"80",X"F5",X"1F",X"29",X"80",X"C6",X"1E",
		X"65",X"80",X"40",X"80",X"44",X"64",X"4C",X"01",X"75",X"81",X"11",X"64",X"10",X"00",X"C0",X"9F",
		X"40",X"80",X"44",X"64",X"3B",X"01",X"B1",X"81",X"11",X"64",X"EC",X"00",X"C5",X"9F",X"DE",X"1F",
		X"E0",X"9F",X"FF",X"1F",X"1F",X"80",X"C7",X"1F",X"08",X"80",X"FF",X"1F",X"D6",X"9F",X"84",X"1F",
		X"21",X"80",X"40",X"80",X"44",X"64",X"30",X"01",X"F2",X"81",X"11",X"64",X"0D",X"00",X"BE",X"9F",
		X"00",X"C0",X"44",X"64",X"2B",X"01",X"FF",X"81",X"11",X"64",X"3A",X"01",X"92",X"9F",X"F3",X"1F",
		X"62",X"80",X"AB",X"1F",X"5D",X"80",X"C7",X"1F",X"21",X"80",X"98",X"40",X"31",X"1F",X"6B",X"80",
		X"40",X"80",X"44",X"64",X"1C",X"01",X"3E",X"82",X"11",X"64",X"10",X"00",X"C0",X"9F",X"40",X"80",
		X"44",X"64",X"0E",X"01",X"89",X"82",X"11",X"64",X"9D",X"00",X"B6",X"9F",X"10",X"00",X"CF",X"9F",
		X"2C",X"00",X"ED",X"9F",X"03",X"00",X"10",X"80",X"2C",X"00",X"D7",X"9F",X"08",X"1F",X"5B",X"80",
		X"40",X"80",X"44",X"64",X"FB",X"00",X"CC",X"82",X"11",X"64",X"11",X"00",X"BC",X"9F",X"00",X"C0",
		X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
