library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity dderby_sp_bits_2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of dderby_sp_bits_2 is
	type rom is array(0 to  32767) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"97",X"00",X"00",X"99",X"92",X"00",X"03",X"26",X"79",
		X"00",X"0E",X"22",X"97",X"00",X"0E",X"99",X"92",X"00",X"0E",X"22",X"76",X"00",X"00",X"22",X"76",
		X"00",X"00",X"77",X"76",X"00",X"00",X"22",X"76",X"00",X"03",X"22",X"76",X"00",X"37",X"99",X"76",
		X"00",X"37",X"99",X"76",X"00",X"03",X"22",X"76",X"00",X"00",X"22",X"76",X"00",X"00",X"77",X"76",
		X"00",X"00",X"22",X"76",X"00",X"0E",X"22",X"76",X"00",X"0E",X"99",X"92",X"00",X"0E",X"22",X"97",
		X"00",X"03",X"26",X"79",X"00",X"00",X"99",X"92",X"00",X"00",X"99",X"97",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"99",X"99",X"70",X"00",X"22",X"77",X"90",X"00",X"66",X"66",X"66",X"00",
		X"99",X"99",X"00",X"00",X"22",X"92",X"00",X"00",X"66",X"92",X"99",X"00",X"66",X"79",X"99",X"00",
		X"66",X"29",X"00",X"00",X"66",X"29",X"00",X"00",X"66",X"29",X"00",X"00",X"66",X"29",X"00",X"00",
		X"66",X"29",X"00",X"00",X"66",X"29",X"00",X"00",X"66",X"29",X"00",X"00",X"66",X"29",X"00",X"00",
		X"66",X"79",X"99",X"00",X"66",X"92",X"99",X"00",X"22",X"92",X"00",X"00",X"99",X"99",X"00",X"00",
		X"66",X"66",X"66",X"00",X"22",X"77",X"90",X"00",X"99",X"99",X"70",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E3",X"90",X"00",X"00",X"92",X"99",
		X"00",X"00",X"00",X"99",X"00",X"00",X"02",X"62",X"00",X"00",X"22",X"22",X"00",X"00",X"29",X"22",
		X"00",X"00",X"27",X"22",X"00",X"00",X"22",X"29",X"00",X"00",X"62",X"96",X"00",X"00",X"66",X"29",
		X"00",X"00",X"26",X"69",X"00",X"00",X"22",X"99",X"00",X"00",X"72",X"99",X"00",X"0E",X"77",X"99",
		X"00",X"0E",X"22",X"99",X"00",X"0E",X"22",X"92",X"00",X"09",X"92",X"92",X"00",X"00",X"29",X"96",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"97",X"00",X"00",X"00",X"27",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"92",X"00",X"00",X"00",
		X"99",X"70",X"00",X"00",X"29",X"79",X"00",X"00",X"62",X"22",X"00",X"00",X"66",X"22",X"00",X"00",
		X"66",X"72",X"90",X"00",X"66",X"22",X"90",X"00",X"66",X"22",X"99",X"00",X"66",X"22",X"66",X"00",
		X"00",X"00",X"66",X"76",X"00",X"00",X"77",X"22",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"22",
		X"00",X"00",X"00",X"96",X"00",X"00",X"00",X"26",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"97",
		X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"22",X"20",X"00",X"66",X"22",X"70",X"00",X"66",X"29",X"70",X"00",X"66",X"29",X"70",X"00",
		X"62",X"29",X"99",X"00",X"62",X"92",X"09",X"00",X"29",X"92",X"09",X"00",X"69",X"22",X"09",X"00",
		X"26",X"22",X"09",X"00",X"72",X"22",X"99",X"00",X"22",X"22",X"90",X"00",X"72",X"22",X"90",X"00",
		X"09",X"92",X"90",X"00",X"00",X"29",X"00",X"00",X"00",X"62",X"00",X"00",X"00",X"76",X"00",X"00",
		X"00",X"97",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"27",X"00",X"00",X"00",X"22",
		X"00",X"00",X"00",X"62",X"00",X"00",X"99",X"26",X"00",X"00",X"77",X"26",X"00",X"00",X"76",X"92",
		X"00",X"00",X"72",X"29",X"00",X"00",X"72",X"22",X"00",X"00",X"72",X"22",X"00",X"00",X"27",X"29",
		X"00",X"00",X"77",X"92",X"00",X"00",X"27",X"22",X"00",X"00",X"22",X"29",X"00",X"00",X"92",X"96",
		X"00",X"00",X"29",X"69",X"00",X"00",X"67",X"99",X"00",X"00",X"62",X"99",X"00",X"00",X"26",X"99",
		X"00",X"00",X"92",X"96",X"00",X"00",X"97",X"66",X"00",X"00",X"99",X"66",X"00",X"00",X"99",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"79",X"00",X"00",X"00",X"27",X"00",X"00",X"00",X"72",X"00",X"00",X"00",
		X"62",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"27",X"00",X"00",X"00",
		X"62",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"90",X"00",X"00",X"66",X"29",X"00",X"00",
		X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"26",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"97",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"22",
		X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"27",X"00",X"00",X"66",X"22",X"00",X"00",X"66",X"27",X"00",X"00",X"62",X"22",X"00",X"00",
		X"67",X"22",X"00",X"00",X"29",X"29",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"92",X"90",X"00",
		X"99",X"22",X"90",X"00",X"99",X"22",X"70",X"00",X"99",X"22",X"70",X"00",X"92",X"22",X"67",X"00",
		X"22",X"62",X"67",X"00",X"22",X"26",X"79",X"00",X"22",X"62",X"90",X"00",X"22",X"26",X"00",X"00",
		X"76",X"29",X"00",X"00",X"72",X"97",X"00",X"00",X"97",X"70",X"00",X"00",X"97",X"90",X"00",X"00",
		X"99",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"79",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"62",X"00",X"00",X"03",X"62",
		X"00",X"00",X"EE",X"26",X"00",X"00",X"EE",X"66",X"00",X"00",X"33",X"22",X"00",X"00",X"72",X"26",
		X"00",X"00",X"72",X"22",X"00",X"00",X"72",X"29",X"00",X"00",X"79",X"29",X"00",X"00",X"09",X"29",
		X"00",X"00",X"09",X"97",X"00",X"00",X"09",X"22",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"62",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"22",
		X"00",X"00",X"00",X"26",X"00",X"00",X"00",X"26",X"00",X"00",X"00",X"26",X"00",X"00",X"00",X"92",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"79",X"00",X"00",X"00",
		X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"69",X"00",X"00",X"00",
		X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"22",X"00",X"00",X"00",
		X"79",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"29",X"00",X"00",X"00",
		X"22",X"00",X"00",X"00",X"62",X"00",X"00",X"00",X"62",X"00",X"00",X"00",X"62",X"00",X"00",X"00",
		X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",
		X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"69",
		X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"72",X"00",X"00",X"00",X"72",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"70",X"00",X"00",X"66",X"70",X"00",X"00",
		X"22",X"70",X"00",X"00",X"99",X"27",X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"29",X"00",X"00",
		X"99",X"29",X"00",X"00",X"99",X"27",X"00",X"00",X"72",X"22",X"00",X"00",X"22",X"26",X"00",X"00",
		X"22",X"26",X"00",X"00",X"99",X"96",X"00",X"00",X"22",X"92",X"00",X"00",X"22",X"92",X"00",X"00",
		X"22",X"29",X"00",X"00",X"22",X"77",X"00",X"00",X"22",X"90",X"00",X"00",X"22",X"99",X"00",X"00",
		X"22",X"99",X"00",X"00",X"77",X"99",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"09",X"00",
		X"00",X"99",X"99",X"00",X"00",X"90",X"70",X"00",X"00",X"29",X"79",X"00",X"00",X"29",X"22",X"00",
		X"00",X"29",X"72",X"00",X"00",X"29",X"72",X"00",X"00",X"29",X"72",X"00",X"00",X"29",X"72",X"00",
		X"00",X"29",X"72",X"00",X"00",X"29",X"22",X"00",X"00",X"29",X"99",X"00",X"00",X"99",X"22",X"00",
		X"00",X"22",X"77",X"00",X"00",X"29",X"62",X"00",X"00",X"92",X"99",X"00",X"00",X"69",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"97",X"77",X"00",X"00",X"72",X"66",X"00",X"00",X"22",X"66",X"00",
		X"00",X"92",X"66",X"00",X"00",X"92",X"66",X"00",X"00",X"92",X"66",X"00",X"00",X"92",X"66",X"00",
		X"00",X"92",X"66",X"00",X"00",X"92",X"66",X"00",X"00",X"92",X"66",X"00",X"00",X"92",X"66",X"00",
		X"00",X"92",X"66",X"00",X"00",X"26",X"22",X"00",X"00",X"69",X"99",X"00",X"00",X"79",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"29",X"99",X"00",X"00",X"27",X"77",X"00",
		X"00",X"22",X"22",X"00",X"00",X"99",X"29",X"00",X"00",X"92",X"72",X"00",X"00",X"92",X"22",X"00",
		X"00",X"92",X"22",X"00",X"00",X"92",X"22",X"00",X"00",X"92",X"22",X"00",X"00",X"92",X"22",X"00",
		X"00",X"92",X"22",X"00",X"00",X"99",X"99",X"00",X"00",X"77",X"77",X"00",X"00",X"09",X"09",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"9A",X"00",X"00",X"00",X"CA",X"00",X"00",X"00",X"AA",
		X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",
		X"00",X"00",X"09",X"00",X"00",X"00",X"9A",X"00",X"00",X"00",X"AB",X"00",X"00",X"00",X"BA",X"00",
		X"00",X"00",X"AD",X"00",X"00",X"00",X"DD",X"00",X"00",X"09",X"D9",X"00",X"00",X"99",X"99",X"00",
		X"00",X"11",X"90",X"00",X"00",X"11",X"00",X"00",X"00",X"14",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"41",X"00",X"00",X"09",X"11",X"00",X"00",X"91",X"10",X"00",X"00",X"91",X"19",X"00",X"00",
		X"91",X"19",X"00",X"00",X"91",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"09",X"90",X"00",X"00",
		X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"9A",
		X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"D9",X"00",X"00",X"09",X"99",
		X"00",X"00",X"9A",X"99",X"00",X"00",X"AD",X"90",X"00",X"00",X"D9",X"00",X"00",X"00",X"9D",X"00",
		X"00",X"00",X"DA",X"00",X"00",X"99",X"AD",X"00",X"00",X"DD",X"D9",X"00",X"00",X"AA",X"99",X"00",
		X"00",X"AA",X"99",X"00",X"00",X"AA",X"90",X"00",X"00",X"AD",X"00",X"00",X"00",X"DA",X"00",X"00",
		X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"FD",X"00",X"00",X"00",X"DD",X"00",X"00",
		X"00",X"FD",X"00",X"00",X"09",X"DD",X"00",X"00",X"0F",X"99",X"00",X"00",X"0F",X"99",X"00",X"00",
		X"09",X"90",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"99",X"99",X"22",X"00",X"22",X"77",X"22",X"00",X"66",X"66",X"26",X"00",
		X"99",X"99",X"20",X"00",X"22",X"92",X"00",X"00",X"66",X"92",X"99",X"00",X"66",X"79",X"99",X"00",
		X"66",X"29",X"00",X"00",X"66",X"29",X"00",X"00",X"66",X"29",X"00",X"00",X"66",X"29",X"00",X"00",
		X"66",X"29",X"00",X"00",X"66",X"29",X"00",X"00",X"66",X"29",X"00",X"00",X"66",X"29",X"00",X"00",
		X"66",X"79",X"99",X"00",X"66",X"92",X"99",X"00",X"22",X"92",X"00",X"00",X"99",X"99",X"00",X"00",
		X"66",X"66",X"66",X"00",X"22",X"77",X"90",X"00",X"99",X"99",X"70",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"97",X"00",X"00",X"00",X"27",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"92",X"00",X"00",X"00",
		X"99",X"70",X"00",X"00",X"29",X"79",X"00",X"00",X"62",X"22",X"00",X"00",X"66",X"22",X"00",X"00",
		X"66",X"72",X"90",X"00",X"66",X"22",X"90",X"00",X"66",X"22",X"22",X"00",X"66",X"22",X"22",X"00",
		X"66",X"22",X"20",X"00",X"66",X"22",X"70",X"00",X"66",X"29",X"70",X"00",X"66",X"29",X"70",X"00",
		X"62",X"29",X"99",X"00",X"62",X"92",X"09",X"00",X"29",X"92",X"09",X"00",X"69",X"22",X"09",X"00",
		X"26",X"22",X"09",X"00",X"72",X"29",X"99",X"00",X"22",X"99",X"90",X"00",X"72",X"99",X"90",X"00",
		X"09",X"99",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"66",X"00",X"00",
		X"00",X"67",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"27",X"00",X"00",X"66",X"22",X"00",X"00",X"66",X"27",X"00",X"00",X"62",X"22",X"00",X"00",
		X"67",X"22",X"00",X"00",X"29",X"29",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"92",X"90",X"00",
		X"99",X"22",X"90",X"00",X"99",X"22",X"20",X"00",X"99",X"22",X"70",X"00",X"92",X"22",X"97",X"00",
		X"22",X"99",X"97",X"00",X"22",X"99",X"79",X"00",X"22",X"99",X"90",X"00",X"22",X"99",X"00",X"00",
		X"76",X"99",X"00",X"00",X"72",X"97",X"00",X"00",X"97",X"70",X"00",X"00",X"97",X"90",X"00",X"00",
		X"09",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"70",X"00",X"00",X"66",X"70",X"00",X"00",
		X"22",X"70",X"00",X"00",X"99",X"27",X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"29",X"00",X"00",
		X"99",X"29",X"00",X"00",X"99",X"27",X"00",X"00",X"92",X"22",X"00",X"00",X"22",X"26",X"00",X"00",
		X"22",X"96",X"00",X"00",X"99",X"26",X"00",X"00",X"22",X"22",X"00",X"00",X"99",X"22",X"00",X"00",
		X"99",X"22",X"00",X"00",X"99",X"77",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"77",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"69",
		X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"72",X"00",X"00",X"00",X"72",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"92",X"66",X"00",X"00",X"92",X"66",X"00",X"00",X"92",X"66",X"00",X"00",X"92",X"66",X"00",
		X"00",X"92",X"66",X"00",X"00",X"26",X"22",X"00",X"00",X"69",X"99",X"00",X"00",X"79",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"29",X"99",X"00",X"00",X"27",X"77",X"00",
		X"00",X"22",X"22",X"00",X"00",X"99",X"29",X"00",X"00",X"92",X"72",X"00",X"00",X"92",X"22",X"00",
		X"00",X"99",X"22",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"92",X"00",X"00",X"99",X"92",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"97",X"77",X"00",X"00",X"99",X"09",X"00",
		X"00",X"66",X"99",X"00",X"00",X"69",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"97",X"00",X"00",X"99",X"92",X"00",X"00",X"99",X"79",
		X"00",X"00",X"99",X"97",X"00",X"00",X"22",X"92",X"00",X"00",X"29",X"76",X"00",X"00",X"22",X"76",
		X"00",X"00",X"99",X"76",X"00",X"00",X"D9",X"76",X"00",X"00",X"DD",X"76",X"00",X"00",X"9D",X"76",
		X"00",X"00",X"9D",X"76",X"00",X"00",X"9D",X"76",X"00",X"00",X"DD",X"76",X"00",X"00",X"D9",X"76",
		X"00",X"00",X"99",X"76",X"00",X"00",X"99",X"76",X"00",X"0E",X"22",X"92",X"00",X"0E",X"22",X"97",
		X"00",X"0E",X"26",X"79",X"00",X"00",X"99",X"92",X"00",X"00",X"99",X"97",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"9E",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"93",X"00",
		X"00",X"00",X"00",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"92",
		X"00",X"00",X"DD",X"22",X"00",X"00",X"DD",X"99",X"00",X"00",X"9D",X"26",X"00",X"00",X"DD",X"29",
		X"00",X"00",X"D9",X"69",X"00",X"00",X"D9",X"99",X"00",X"00",X"DD",X"99",X"00",X"0E",X"99",X"99",
		X"00",X"00",X"99",X"99",X"00",X"07",X"99",X"92",X"00",X"09",X"29",X"92",X"00",X"00",X"22",X"96",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"90",
		X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"07",X"29",X"00",X"00",X"79",X"22",
		X"00",X"00",X"79",X"92",X"00",X"00",X"79",X"92",X"00",X"00",X"9D",X"22",X"00",X"00",X"DD",X"22",
		X"00",X"00",X"99",X"92",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"96",
		X"00",X"00",X"29",X"69",X"00",X"00",X"62",X"99",X"00",X"00",X"62",X"99",X"00",X"00",X"26",X"99",
		X"00",X"00",X"92",X"96",X"00",X"00",X"97",X"66",X"00",X"00",X"99",X"66",X"00",X"00",X"99",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"29",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"22",X"00",X"00",X"00",
		X"79",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"29",X"00",X"00",X"00",
		X"22",X"00",X"00",X"00",X"62",X"00",X"00",X"00",X"62",X"00",X"00",X"00",X"62",X"00",X"00",X"00",
		X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"79",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"7E",X"DD",X"00",X"00",X"EE",X"D9",X"00",X"00",X"EE",X"9D",X"00",X"00",X"33",X"DD",
		X"00",X"00",X"72",X"D9",X"00",X"00",X"72",X"DD",X"00",X"00",X"79",X"D2",X"00",X"00",X"09",X"22",
		X"00",X"00",X"09",X"22",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"62",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"22",
		X"00",X"00",X"00",X"26",X"00",X"00",X"00",X"26",X"00",X"00",X"00",X"26",X"00",X"00",X"00",X"92",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"EE",X"99",X"00",
		X"00",X"EE",X"99",X"00",X"00",X"90",X"70",X"E0",X"00",X"29",X"79",X"E0",X"00",X"29",X"DD",X"00",
		X"00",X"29",X"D9",X"00",X"00",X"29",X"D9",X"00",X"00",X"29",X"D9",X"00",X"00",X"29",X"D9",X"00",
		X"00",X"29",X"D9",X"00",X"00",X"29",X"22",X"00",X"00",X"29",X"29",X"00",X"00",X"99",X"99",X"00",
		X"00",X"22",X"77",X"00",X"00",X"29",X"62",X"00",X"00",X"92",X"99",X"00",X"00",X"69",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"97",X"77",X"00",X"00",X"72",X"66",X"00",X"00",X"22",X"66",X"00",
		X"00",X"92",X"66",X"00",X"00",X"92",X"66",X"00",X"00",X"92",X"66",X"00",X"00",X"92",X"66",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"97",X"00",X"00",X"99",X"92",X"00",X"00",X"99",X"79",
		X"00",X"00",X"99",X"97",X"00",X"00",X"22",X"92",X"00",X"00",X"29",X"76",X"00",X"00",X"22",X"76",
		X"00",X"00",X"99",X"76",X"00",X"00",X"D9",X"76",X"00",X"00",X"DD",X"76",X"00",X"00",X"9D",X"76",
		X"00",X"00",X"9D",X"76",X"00",X"00",X"9D",X"76",X"00",X"00",X"DD",X"76",X"00",X"00",X"D9",X"76",
		X"00",X"00",X"99",X"76",X"00",X"00",X"99",X"76",X"00",X"00",X"22",X"92",X"00",X"00",X"22",X"97",
		X"00",X"00",X"26",X"79",X"00",X"00",X"99",X"92",X"00",X"00",X"99",X"97",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"97",X"00",X"00",X"00",X"27",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"92",X"00",X"00",X"00",
		X"99",X"70",X"00",X"00",X"29",X"79",X"00",X"00",X"62",X"22",X"00",X"00",X"66",X"22",X"90",X"00",
		X"66",X"72",X"90",X"00",X"66",X"22",X"90",X"00",X"66",X"22",X"22",X"00",X"66",X"22",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"97",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"93",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"92",
		X"00",X"00",X"DD",X"22",X"00",X"00",X"DD",X"99",X"00",X"00",X"9D",X"26",X"00",X"00",X"DD",X"29",
		X"00",X"00",X"D9",X"69",X"00",X"00",X"D9",X"99",X"00",X"00",X"DD",X"99",X"00",X"00",X"99",X"99",
		X"00",X"00",X"99",X"99",X"00",X"07",X"99",X"92",X"00",X"09",X"29",X"92",X"00",X"00",X"22",X"96",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",
		X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"07",X"29",X"00",X"00",X"79",X"22",
		X"00",X"00",X"79",X"92",X"00",X"00",X"79",X"92",X"00",X"00",X"9D",X"22",X"00",X"00",X"DD",X"22",
		X"00",X"00",X"99",X"92",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"96",
		X"00",X"00",X"29",X"69",X"00",X"00",X"62",X"99",X"00",X"00",X"62",X"99",X"00",X"00",X"26",X"99",
		X"00",X"00",X"92",X"96",X"00",X"00",X"97",X"66",X"00",X"00",X"99",X"66",X"00",X"00",X"99",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"29",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"22",X"00",X"00",X"00",
		X"79",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"29",X"00",X"00",X"00",
		X"22",X"00",X"00",X"00",X"62",X"00",X"00",X"00",X"62",X"00",X"00",X"00",X"62",X"00",X"00",X"00",
		X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"79",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"99",X"00",X"00",X"EE",X"99",
		X"00",X"00",X"EE",X"DD",X"00",X"00",X"EE",X"D9",X"00",X"00",X"33",X"9D",X"00",X"00",X"32",X"DD",
		X"00",X"00",X"72",X"D9",X"00",X"00",X"72",X"DD",X"00",X"00",X"79",X"D2",X"00",X"00",X"99",X"22",
		X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"62",
		X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"22",
		X"00",X"00",X"00",X"26",X"00",X"00",X"00",X"26",X"00",X"00",X"00",X"26",X"00",X"00",X"00",X"92",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"90",X"00",X"00",X"E9",X"99",X"E0",
		X"00",X"99",X"99",X"E0",X"00",X"90",X"70",X"E0",X"00",X"29",X"79",X"00",X"00",X"29",X"DD",X"00",
		X"00",X"29",X"D9",X"00",X"00",X"29",X"D9",X"00",X"00",X"29",X"D9",X"00",X"00",X"29",X"D9",X"00",
		X"00",X"29",X"D9",X"00",X"00",X"29",X"22",X"00",X"00",X"29",X"29",X"00",X"00",X"99",X"99",X"00",
		X"00",X"22",X"77",X"00",X"00",X"29",X"62",X"00",X"00",X"92",X"99",X"00",X"00",X"69",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"97",X"77",X"00",X"00",X"72",X"66",X"00",X"00",X"22",X"66",X"00",
		X"00",X"92",X"66",X"00",X"00",X"92",X"66",X"00",X"00",X"92",X"66",X"00",X"00",X"92",X"66",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"99",X"99",X"70",X"00",X"22",X"77",X"70",X"00",X"66",X"66",X"20",X"00",
		X"99",X"99",X"60",X"00",X"22",X"99",X"60",X"00",X"66",X"92",X"29",X"00",X"66",X"79",X"99",X"00",
		X"66",X"29",X"00",X"00",X"66",X"29",X"00",X"00",X"66",X"29",X"00",X"00",X"66",X"29",X"00",X"00",
		X"66",X"29",X"00",X"00",X"66",X"29",X"00",X"00",X"66",X"29",X"00",X"00",X"66",X"29",X"00",X"00",
		X"66",X"79",X"99",X"00",X"66",X"92",X"99",X"00",X"22",X"92",X"00",X"00",X"99",X"99",X"00",X"00",
		X"66",X"66",X"66",X"00",X"22",X"77",X"90",X"00",X"99",X"00",X"70",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"22",X"00",X"00",X"66",X"22",X"70",X"00",X"66",X"29",X"70",X"00",X"66",X"29",X"70",X"00",
		X"62",X"29",X"99",X"00",X"62",X"92",X"09",X"00",X"29",X"92",X"09",X"00",X"69",X"22",X"09",X"00",
		X"26",X"22",X"09",X"00",X"72",X"22",X"99",X"00",X"22",X"29",X"90",X"00",X"72",X"29",X"90",X"00",
		X"09",X"99",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"66",X"00",X"00",
		X"00",X"67",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"66",X"76",X"00",X"00",X"77",X"22",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"22",
		X"00",X"00",X"99",X"96",X"00",X"00",X"00",X"26",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"97",
		X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"22",X"00",X"00",X"66",X"27",X"00",X"00",X"62",X"22",X"00",X"00",X"67",X"22",X"00",X"00",
		X"29",X"29",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"92",X"00",X"00",X"99",X"22",X"00",X"00",
		X"99",X"22",X"00",X"00",X"99",X"22",X"70",X"00",X"92",X"22",X"97",X"00",X"22",X"22",X"97",X"00",
		X"22",X"99",X"79",X"00",X"22",X"99",X"90",X"00",X"22",X"99",X"00",X"00",X"76",X"99",X"00",X"00",
		X"72",X"97",X"00",X"00",X"97",X"70",X"00",X"00",X"07",X"90",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"70",X"00",X"00",X"66",X"70",X"00",X"00",
		X"22",X"70",X"00",X"00",X"99",X"27",X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"29",X"00",X"00",
		X"99",X"29",X"00",X"00",X"99",X"27",X"00",X"00",X"92",X"22",X"00",X"00",X"22",X"26",X"00",X"00",
		X"22",X"96",X"00",X"00",X"99",X"26",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",
		X"92",X"22",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"92",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"77",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"69",
		X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"72",X"00",X"00",X"00",X"72",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"92",X"66",X"00",X"00",X"92",X"66",X"00",X"00",X"92",X"66",X"00",X"00",X"92",X"66",X"00",
		X"00",X"92",X"66",X"00",X"00",X"26",X"22",X"00",X"00",X"69",X"99",X"00",X"00",X"79",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"29",X"99",X"00",X"00",X"27",X"77",X"90",
		X"00",X"22",X"22",X"90",X"00",X"99",X"29",X"90",X"00",X"92",X"72",X"90",X"00",X"92",X"22",X"90",
		X"00",X"99",X"22",X"90",X"00",X"99",X"22",X"90",X"00",X"99",X"22",X"90",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"97",X"77",X"00",X"00",X"99",X"09",X"00",
		X"00",X"66",X"99",X"00",X"00",X"69",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"10",
		X"00",X"09",X"00",X"11",X"00",X"00",X"09",X"01",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"10",X"00",X"10",X"00",X"01",X"01",X"00",X"00",X"01",X"12",X"00",X"00",X"01",X"91",X"10",
		X"00",X"00",X"00",X"10",X"00",X"99",X"F0",X"11",X"00",X"99",X"00",X"11",X"00",X"09",X"00",X"10",
		X"00",X"00",X"22",X"11",X"00",X"11",X"11",X"11",X"00",X"00",X"10",X"90",X"00",X"00",X"00",X"10",
		X"00",X"99",X"99",X"10",X"00",X"99",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"10",X"00",X"10",X"00",X"00",X"00",X"11",X"00",X"00",
		X"00",X"90",X"00",X"00",X"00",X"91",X"11",X"00",X"00",X"01",X"11",X"00",X"00",X"02",X"10",X"00",
		X"09",X"12",X"21",X"00",X"09",X"01",X"22",X"01",X"00",X"00",X"02",X"11",X"00",X"00",X"01",X"10",
		X"00",X"19",X"01",X"00",X"00",X"90",X"01",X"00",X"10",X"90",X"20",X"00",X"11",X"90",X"92",X"09",
		X"00",X"09",X"02",X"99",X"90",X"F9",X"11",X"90",X"09",X"0F",X"01",X"00",X"09",X"1F",X"11",X"00",
		X"00",X"11",X"21",X"00",X"01",X"11",X"11",X"10",X"00",X"00",X"01",X"10",X"00",X"00",X"10",X"00",
		X"00",X"99",X"00",X"99",X"00",X"99",X"99",X"99",X"00",X"09",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"01",X"00",X"10",X"00",X"11",X"00",X"10",X"00",X"10",X"00",X"10",X"00",X"19",
		X"00",X"11",X"00",X"10",X"00",X"01",X"00",X"10",X"00",X"12",X"00",X"02",X"00",X"01",X"00",X"11",
		X"00",X"11",X"00",X"02",X"00",X"11",X"10",X"02",X"00",X"11",X"11",X"01",X"00",X"00",X"99",X"11",
		X"00",X"00",X"01",X"10",X"00",X"00",X"91",X"01",X"00",X"00",X"91",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"F9",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"10",X"99",X"00",X"91",X"09",X"99",X"00",X"09",X"90",X"99",X"01",X"11",X"90",X"90",
		X"00",X"10",X"99",X"00",X"90",X"00",X"99",X"00",X"09",X"01",X"99",X"00",X"00",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"10",X"11",X"00",X"11",X"00",
		X"11",X"00",X"01",X"00",X"11",X"10",X"01",X"00",X"01",X"11",X"01",X"09",X"90",X"01",X"01",X"09",
		X"90",X"11",X"11",X"90",X"00",X"00",X"11",X"00",X"00",X"00",X"10",X"00",X"00",X"09",X"01",X"00",
		X"09",X"09",X"11",X"00",X"90",X"99",X"11",X"00",X"99",X"09",X"10",X"00",X"99",X"99",X"01",X"01",
		X"90",X"99",X"22",X"11",X"99",X"99",X"10",X"00",X"90",X"99",X"00",X"99",X"99",X"99",X"01",X"19",
		X"90",X"90",X"11",X"99",X"99",X"00",X"11",X"09",X"00",X"99",X"10",X"99",X"00",X"99",X"00",X"99",
		X"10",X"10",X"00",X"00",X"11",X"00",X"00",X"00",X"01",X"10",X"00",X"00",X"90",X"10",X"00",X"00",
		X"09",X"11",X"00",X"00",X"00",X"01",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"99",X"00",
		X"01",X"00",X"00",X"00",X"00",X"11",X"10",X"00",X"11",X"10",X"99",X"00",X"00",X"00",X"00",X"00",
		X"99",X"00",X"01",X"00",X"99",X"99",X"10",X"11",X"09",X"99",X"11",X"11",X"09",X"91",X"09",X"01",
		X"00",X"91",X"19",X"01",X"00",X"11",X"11",X"00",X"00",X"01",X"99",X"00",X"00",X"01",X"11",X"00",
		X"00",X"01",X"11",X"11",X"00",X"10",X"00",X"01",X"00",X"01",X"10",X"11",X"00",X"11",X"00",X"10",
		X"00",X"11",X"99",X"01",X"01",X"19",X"99",X"00",X"00",X"19",X"99",X"00",X"00",X"00",X"99",X"99",
		X"00",X"99",X"00",X"99",X"00",X"90",X"00",X"99",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"90",
		X"00",X"00",X"09",X"00",X"00",X"90",X"99",X"00",X"00",X"90",X"90",X"00",X"00",X"01",X"01",X"00",
		X"00",X"F0",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"10",X"00",X"00",
		X"00",X"10",X"10",X"00",X"00",X"99",X"10",X"10",X"00",X"90",X"10",X"00",X"99",X"09",X"10",X"00",
		X"99",X"00",X"10",X"00",X"99",X"00",X"10",X"11",X"11",X"00",X"11",X"01",X"01",X"00",X"01",X"99",
		X"F0",X"11",X"00",X"99",X"00",X"11",X"01",X"99",X"09",X"10",X"00",X"90",X"99",X"01",X"11",X"00",
		X"01",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"10",X"00",X"00",
		X"00",X"10",X"90",X"00",X"00",X"10",X"99",X"00",X"00",X"99",X"90",X"00",X"99",X"00",X"90",X"00",
		X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",
		X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",
		X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",
		X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",
		X"11",X"11",X"00",X"00",X"11",X"99",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",
		X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"10",X"00",X"00",X"10",X"00",
		X"00",X"00",X"11",X"09",X"00",X"01",X"11",X"99",X"00",X"14",X"11",X"90",X"00",X"41",X"41",X"00",
		X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"19",X"00",X"00",X"91",X"90",X"00",
		X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"99",
		X"00",X"01",X"11",X"99",X"00",X"11",X"11",X"00",X"00",X"11",X"00",X"00",X"00",X"99",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"11",X"00",
		X"00",X"00",X"21",X"00",X"00",X"11",X"10",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"11",X"00",
		X"00",X"00",X"21",X"00",X"00",X"00",X"20",X"00",X"00",X"11",X"21",X"00",X"00",X"10",X"01",X"00",
		X"00",X"11",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"11",X"10",X"00",X"00",X"00",X"20",X"00",
		X"00",X"00",X"10",X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"10",X"00",
		X"00",X"11",X"20",X"00",X"00",X"00",X"10",X"00",X"00",X"11",X"11",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"90",X"9F",X"00",X"00",X"9F",X"F0",X"00",
		X"00",X"9F",X"00",X"90",X"00",X"90",X"FF",X"99",X"00",X"99",X"9F",X"F9",X"00",X"99",X"99",X"FF",
		X"00",X"99",X"99",X"F0",X"00",X"FF",X"99",X"FF",X"00",X"F0",X"FF",X"9F",X"00",X"FF",X"0F",X"FF",
		X"00",X"9F",X"0F",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"00",
		X"00",X"99",X"9F",X"F9",X"00",X"9F",X"9F",X"90",X"00",X"9F",X"99",X"F0",X"00",X"FF",X"FF",X"90",
		X"00",X"F9",X"0F",X"00",X"00",X"99",X"90",X"09",X"00",X"99",X"99",X"90",X"00",X"09",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"9F",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"F0",X"90",X"00",X"00",X"F0",X"99",X"00",X"00",X"FF",X"F9",X"00",X"00",X"09",X"FF",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"F0",X"9F",X"00",X"00",X"FF",X"99",X"00",X"00",X"FF",X"99",X"00",
		X"00",X"9F",X"00",X"00",X"0F",X"90",X"F9",X"00",X"09",X"99",X"90",X"00",X"00",X"0F",X"90",X"00",
		X"00",X"F9",X"00",X"00",X"00",X"99",X"09",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"F9",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"0F",X"09",X"9F",X"00",X"09",X"00",X"F9",
		X"00",X"00",X"00",X"0F",X"00",X"0F",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"09",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"F9",X"00",X"00",X"90",X"00",X"90",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",
		X"00",X"00",X"0D",X"A9",X"00",X"00",X"0D",X"A9",X"00",X"00",X"9A",X"A9",X"00",X"00",X"AA",X"90",
		X"00",X"00",X"BD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",X"D9",X"00",
		X"00",X"00",X"90",X"00",X"00",X"09",X"90",X"00",X"00",X"9A",X"00",X"00",X"00",X"AA",X"00",X"00",
		X"00",X"AD",X"00",X"00",X"00",X"DD",X"00",X"00",X"0A",X"DD",X"00",X"00",X"0A",X"99",X"00",X"00",
		X"0A",X"99",X"00",X"00",X"0D",X"90",X"00",X"00",X"09",X"90",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"99",X"00",X"09",X"99",X"22",X"00",X"09",X"22",X"29",
		X"00",X"99",X"66",X"99",X"00",X"99",X"22",X"22",X"00",X"99",X"22",X"99",X"00",X"99",X"22",X"99",
		X"00",X"99",X"22",X"99",X"00",X"99",X"77",X"99",X"00",X"99",X"66",X"99",X"00",X"99",X"22",X"99",
		X"00",X"99",X"22",X"99",X"00",X"99",X"66",X"99",X"00",X"99",X"77",X"99",X"00",X"99",X"22",X"99",
		X"00",X"99",X"22",X"99",X"00",X"99",X"22",X"99",X"00",X"99",X"22",X"22",X"00",X"99",X"66",X"99",
		X"00",X"09",X"22",X"29",X"00",X"09",X"99",X"22",X"00",X"09",X"99",X"99",X"00",X"09",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"99",X"99",X"09",X"00",X"22",X"99",X"09",X"00",X"99",X"77",X"09",X"00",
		X"99",X"22",X"00",X"00",X"99",X"22",X"00",X"00",X"66",X"22",X"70",X"00",X"66",X"22",X"70",X"00",
		X"66",X"92",X"99",X"00",X"66",X"92",X"70",X"00",X"66",X"92",X"70",X"00",X"66",X"92",X"70",X"00",
		X"66",X"92",X"70",X"00",X"66",X"92",X"70",X"00",X"66",X"92",X"70",X"00",X"66",X"92",X"99",X"00",
		X"66",X"22",X"70",X"00",X"66",X"22",X"70",X"00",X"99",X"22",X"00",X"00",X"99",X"22",X"00",X"00",
		X"99",X"77",X"09",X"00",X"22",X"99",X"09",X"00",X"99",X"99",X"09",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"E9",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"92",X"90",
		X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"99",X"00",X"00",X"72",X"22",X"00",X"09",X"27",X"22",
		X"00",X"09",X"29",X"22",X"00",X"09",X"66",X"99",X"00",X"99",X"22",X"22",X"00",X"99",X"22",X"99",
		X"00",X"99",X"22",X"99",X"00",X"99",X"22",X"99",X"00",X"99",X"62",X"99",X"00",X"99",X"99",X"99",
		X"00",X"9E",X"27",X"99",X"00",X"9E",X"22",X"99",X"00",X"9E",X"22",X"99",X"00",X"99",X"62",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"22",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"79",X"99",X"00",X"00",X"67",X"99",X"00",X"00",
		X"66",X"29",X"00",X"00",X"66",X"22",X"00",X"00",X"66",X"22",X"00",X"00",X"66",X"79",X"00",X"00",
		X"00",X"09",X"26",X"99",X"00",X"00",X"22",X"96",X"00",X"00",X"92",X"26",X"00",X"00",X"99",X"99",
		X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"92",X"90",X"00",X"66",X"99",X"90",X"00",X"66",X"92",X"90",X"00",X"66",X"92",X"90",X"00",
		X"66",X"92",X"00",X"00",X"66",X"22",X"00",X"00",X"29",X"29",X"00",X"00",X"92",X"29",X"90",X"00",
		X"99",X"92",X"99",X"00",X"99",X"22",X"09",X"00",X"22",X"22",X"99",X"00",X"99",X"66",X"99",X"00",
		X"99",X"99",X"99",X"00",X"09",X"29",X"90",X"00",X"00",X"22",X"90",X"00",X"00",X"92",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"29",
		X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"22",X"00",X"00",X"22",X"62",X"00",X"00",X"22",X"62",
		X"00",X"00",X"22",X"26",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"72",
		X"00",X"00",X"76",X"22",X"00",X"09",X"27",X"99",X"00",X"09",X"22",X"96",X"00",X"09",X"22",X"69",
		X"00",X"09",X"22",X"99",X"00",X"00",X"62",X"99",X"00",X"00",X"26",X"99",X"00",X"00",X"22",X"99",
		X"00",X"00",X"22",X"99",X"00",X"00",X"92",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"76",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"92",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"69",X"00",X"00",X"00",
		X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"90",X"00",X"00",X"66",X"29",X"00",X"00",
		X"00",X"00",X"09",X"66",X"00",X"00",X"00",X"76",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"92",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"20",X"00",X"00",X"66",X"92",X"00",X"00",X"66",X"22",X"00",X"00",X"66",X"92",X"00",X"00",
		X"66",X"22",X"00",X"00",X"69",X"22",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"29",X"00",X"00",
		X"99",X"29",X"90",X"00",X"99",X"92",X"90",X"00",X"99",X"22",X"00",X"00",X"99",X"22",X"09",X"00",
		X"29",X"22",X"09",X"00",X"22",X"29",X"99",X"00",X"22",X"29",X"99",X"00",X"22",X"92",X"90",X"00",
		X"92",X"66",X"90",X"00",X"99",X"69",X"00",X"00",X"99",X"99",X"00",X"00",X"09",X"09",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"9E",X"00",X"00",X"09",X"9E",X"00",X"00",X"99",X"72",X"00",X"00",X"99",X"27",
		X"00",X"00",X"99",X"27",X"00",X"00",X"9E",X"67",X"00",X"00",X"EE",X"62",X"00",X"00",X"E9",X"62",
		X"00",X"00",X"99",X"22",X"00",X"00",X"92",X"26",X"00",X"00",X"22",X"26",X"00",X"00",X"66",X"22",
		X"00",X"00",X"92",X"29",X"00",X"00",X"92",X"96",X"00",X"00",X"92",X"66",X"00",X"00",X"99",X"69",
		X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"09",X"99",
		X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"96",X"00",X"00",X"00",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"92",X"00",X"00",X"00",
		X"92",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"69",X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"66",X"00",X"00",X"00",
		X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"96",X"00",X"00",X"00",X"96",
		X"00",X"00",X"00",X"96",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"92",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",
		X"66",X"00",X"00",X"00",X"66",X"90",X"00",X"00",X"79",X"90",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"79",X"00",X"00",X"99",X"79",X"00",X"00",
		X"99",X"27",X"00",X"00",X"22",X"27",X"00",X"00",X"29",X"92",X"00",X"00",X"92",X"92",X"00",X"00",
		X"22",X"97",X"00",X"00",X"22",X"77",X"00",X"00",X"22",X"67",X"00",X"00",X"62",X"70",X"00",X"00",
		X"22",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"66",X"99",X"00",X"00",X"77",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"EE",X"79",X"00",X"00",X"E3",X"22",X"00",X"00",X"33",X"67",X"00",X"00",X"22",X"67",X"00",
		X"00",X"22",X"67",X"00",X"00",X"22",X"62",X"00",X"00",X"22",X"72",X"00",X"00",X"22",X"72",X"00",
		X"00",X"22",X"72",X"00",X"00",X"22",X"72",X"00",X"00",X"22",X"72",X"00",X"00",X"22",X"22",X"00",
		X"00",X"22",X"22",X"00",X"00",X"22",X"99",X"00",X"00",X"29",X"29",X"00",X"00",X"99",X"92",X"00",
		X"00",X"92",X"99",X"00",X"00",X"92",X"99",X"00",X"00",X"92",X"99",X"00",X"00",X"99",X"66",X"00",
		X"00",X"96",X"66",X"00",X"00",X"96",X"66",X"00",X"00",X"96",X"66",X"00",X"00",X"96",X"66",X"00",
		X"00",X"96",X"66",X"00",X"00",X"96",X"66",X"00",X"00",X"96",X"66",X"00",X"00",X"96",X"66",X"00",
		X"00",X"96",X"62",X"00",X"00",X"96",X"62",X"00",X"00",X"92",X"99",X"00",X"00",X"92",X"99",X"00",
		X"00",X"27",X"99",X"00",X"00",X"29",X"99",X"00",X"00",X"29",X"99",X"00",X"00",X"72",X"99",X"00",
		X"00",X"27",X"92",X"00",X"00",X"22",X"22",X"00",X"00",X"29",X"99",X"00",X"00",X"96",X"22",X"00",
		X"00",X"96",X"22",X"00",X"00",X"96",X"22",X"00",X"00",X"96",X"22",X"00",X"00",X"96",X"22",X"00",
		X"00",X"99",X"99",X"00",X"00",X"69",X"66",X"00",X"00",X"77",X"77",X"00",X"00",X"97",X"77",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"95",X"00",X"00",X"05",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"59",X"39",X"00",
		X"00",X"99",X"93",X"00",X"00",X"9D",X"93",X"00",X"00",X"93",X"99",X"00",X"00",X"93",X"99",X"00",
		X"00",X"9D",X"93",X"00",X"00",X"93",X"99",X"00",X"00",X"99",X"93",X"00",X"00",X"99",X"33",X"00",
		X"00",X"09",X"39",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"05",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"0B",X"00",X"00",X"BB",X"00",
		X"00",X"B0",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"09",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"9D",X"00",X"00",X"0B",X"99",X"00",X"00",X"00",X"39",X"00",X"00",X"00",X"99",X"0B",X"00",
		X"00",X"39",X"B0",X"00",X"00",X"99",X"B0",X"0B",X"00",X"99",X"B5",X"00",X"00",X"99",X"BB",X"00",
		X"00",X"00",X"BB",X"00",X"0B",X"B0",X"0B",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"50",X"00",
		X"00",X"00",X"05",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"99",X"99",X"09",X"00",X"22",X"99",X"09",X"00",X"99",X"99",X"09",X"00",
		X"99",X"29",X"90",X"00",X"99",X"22",X"90",X"00",X"66",X"22",X"70",X"00",X"66",X"22",X"70",X"00",
		X"66",X"92",X"99",X"00",X"66",X"92",X"99",X"00",X"66",X"92",X"99",X"00",X"66",X"92",X"99",X"00",
		X"66",X"92",X"99",X"00",X"66",X"92",X"90",X"00",X"66",X"92",X"99",X"00",X"66",X"92",X"99",X"00",
		X"66",X"22",X"99",X"00",X"66",X"22",X"79",X"00",X"99",X"22",X"00",X"00",X"99",X"22",X"00",X"00",
		X"22",X"99",X"09",X"00",X"99",X"99",X"09",X"00",X"99",X"99",X"09",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"22",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"79",X"99",X"00",X"00",X"67",X"99",X"00",X"00",
		X"66",X"29",X"00",X"00",X"66",X"22",X"00",X"00",X"66",X"22",X"00",X"00",X"66",X"79",X"00",X"00",
		X"66",X"92",X"90",X"00",X"66",X"99",X"20",X"00",X"66",X"92",X"20",X"00",X"66",X"92",X"22",X"00",
		X"66",X"92",X"00",X"00",X"66",X"22",X"09",X"00",X"29",X"29",X"99",X"00",X"92",X"29",X"99",X"00",
		X"99",X"92",X"99",X"00",X"22",X"22",X"99",X"00",X"99",X"22",X"00",X"00",X"99",X"22",X"00",X"00",
		X"99",X"22",X"00",X"00",X"09",X"92",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"22",X"00",X"00",
		X"00",X"92",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"20",X"00",X"00",X"66",X"92",X"00",X"00",X"66",X"22",X"00",X"00",X"66",X"92",X"00",X"00",
		X"66",X"22",X"00",X"00",X"69",X"22",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"22",X"00",X"00",
		X"99",X"22",X"90",X"00",X"99",X"92",X"90",X"00",X"99",X"22",X"00",X"00",X"99",X"22",X"09",X"00",
		X"29",X"77",X"99",X"00",X"22",X"79",X"99",X"00",X"92",X"99",X"90",X"00",X"99",X"99",X"90",X"00",
		X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"09",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",
		X"66",X"00",X"00",X"00",X"66",X"90",X"00",X"00",X"79",X"90",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"22",X"27",X"00",X"00",X"29",X"92",X"00",X"00",X"92",X"92",X"00",X"00",
		X"22",X"97",X"00",X"00",X"22",X"22",X"00",X"00",X"29",X"22",X"00",X"00",X"99",X"79",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"79",X"90",X"00",X"00",
		X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"96",X"00",X"00",X"00",X"96",X"00",X"00",X"00",X"96",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",
		X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"96",X"66",X"00",X"00",X"96",X"66",X"00",X"00",X"96",X"66",X"00",X"00",X"96",X"66",X"00",
		X"00",X"96",X"62",X"00",X"00",X"96",X"62",X"00",X"00",X"92",X"99",X"00",X"00",X"92",X"99",X"00",
		X"00",X"27",X"99",X"00",X"00",X"29",X"99",X"00",X"00",X"29",X"99",X"00",X"00",X"72",X"99",X"00",
		X"00",X"27",X"92",X"00",X"00",X"22",X"22",X"00",X"00",X"29",X"99",X"00",X"00",X"96",X"22",X"00",
		X"00",X"96",X"22",X"00",X"00",X"96",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"27",X"22",X"00",
		X"00",X"97",X"77",X"00",X"00",X"69",X"77",X"00",X"00",X"79",X"97",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"90",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"99",X"00",X"09",X"99",X"22",X"00",X"09",X"99",X"29",
		X"00",X"99",X"99",X"99",X"00",X"99",X"92",X"22",X"00",X"99",X"22",X"99",X"00",X"99",X"22",X"99",
		X"00",X"99",X"22",X"99",X"00",X"99",X"77",X"99",X"00",X"99",X"66",X"99",X"00",X"99",X"22",X"99",
		X"00",X"99",X"22",X"99",X"00",X"99",X"66",X"99",X"00",X"99",X"77",X"99",X"00",X"99",X"22",X"99",
		X"00",X"09",X"22",X"99",X"00",X"09",X"22",X"99",X"00",X"00",X"22",X"22",X"00",X"00",X"96",X"99",
		X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"E9",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"92",X"90",
		X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"99",X"00",X"00",X"72",X"29",X"00",X"09",X"27",X"99",
		X"00",X"09",X"29",X"99",X"00",X"09",X"66",X"99",X"00",X"09",X"22",X"22",X"00",X"09",X"22",X"99",
		X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"99",X"00",X"09",X"62",X"99",X"00",X"09",X"99",X"99",
		X"00",X"09",X"27",X"99",X"00",X"03",X"22",X"99",X"00",X"03",X"22",X"99",X"00",X"09",X"62",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"29",
		X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"99",X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"99",
		X"00",X"00",X"22",X"29",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"72",
		X"00",X"00",X"76",X"22",X"00",X"00",X"27",X"99",X"00",X"00",X"22",X"96",X"00",X"00",X"22",X"69",
		X"00",X"00",X"22",X"99",X"00",X"00",X"92",X"99",X"00",X"00",X"96",X"99",X"00",X"00",X"92",X"99",
		X"00",X"00",X"92",X"99",X"00",X"00",X"92",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"76",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"92",X"00",X"00",X"00",
		X"92",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"69",X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"66",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"9E",X"00",X"00",X"09",X"9E",X"00",X"00",X"99",X"72",X"00",X"00",X"99",X"27",
		X"00",X"00",X"99",X"27",X"00",X"00",X"9E",X"67",X"00",X"00",X"EE",X"62",X"00",X"00",X"E9",X"62",
		X"00",X"00",X"E9",X"22",X"00",X"00",X"39",X"26",X"00",X"00",X"99",X"26",X"00",X"00",X"99",X"22",
		X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"96",X"00",X"00",X"99",X"66",X"00",X"00",X"99",X"69",
		X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",
		X"00",X"00",X"99",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"96",X"00",X"00",X"00",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"09",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"9E",X"79",X"00",X"00",X"EE",X"29",X"00",X"00",X"E3",X"67",X"00",X"00",X"99",X"67",X"00",
		X"00",X"92",X"67",X"00",X"00",X"32",X"62",X"00",X"00",X"92",X"72",X"00",X"00",X"92",X"72",X"00",
		X"00",X"22",X"72",X"00",X"00",X"22",X"72",X"00",X"00",X"22",X"72",X"00",X"00",X"22",X"22",X"00",
		X"00",X"22",X"22",X"00",X"00",X"22",X"99",X"00",X"00",X"29",X"29",X"00",X"00",X"99",X"92",X"00",
		X"00",X"92",X"99",X"00",X"00",X"92",X"99",X"00",X"00",X"92",X"99",X"00",X"00",X"99",X"66",X"00",
		X"00",X"96",X"66",X"00",X"00",X"96",X"66",X"00",X"00",X"96",X"66",X"00",X"00",X"96",X"66",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"09",X"99",X"99",X"00",X"09",X"99",X"22",X"00",X"09",X"99",X"29",
		X"00",X"99",X"99",X"99",X"00",X"99",X"92",X"22",X"00",X"99",X"22",X"99",X"00",X"99",X"22",X"99",
		X"00",X"99",X"22",X"99",X"00",X"99",X"77",X"99",X"00",X"99",X"66",X"99",X"00",X"99",X"22",X"99",
		X"00",X"99",X"22",X"99",X"00",X"99",X"66",X"99",X"00",X"99",X"77",X"99",X"00",X"99",X"22",X"99",
		X"00",X"09",X"22",X"99",X"00",X"09",X"22",X"99",X"00",X"03",X"22",X"22",X"00",X"03",X"96",X"99",
		X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"22",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"79",X"99",X"00",X"00",X"67",X"99",X"00",X"00",
		X"66",X"29",X"00",X"00",X"66",X"22",X"00",X"00",X"66",X"22",X"90",X"00",X"66",X"79",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"E9",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"92",X"00",
		X"00",X"00",X"22",X"90",X"00",X"00",X"22",X"99",X"00",X"00",X"72",X"29",X"00",X"09",X"27",X"99",
		X"00",X"09",X"29",X"99",X"00",X"09",X"66",X"99",X"00",X"09",X"22",X"22",X"00",X"09",X"22",X"99",
		X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"99",X"00",X"09",X"62",X"99",X"00",X"09",X"99",X"99",
		X"00",X"09",X"27",X"99",X"00",X"09",X"22",X"99",X"00",X"09",X"22",X"99",X"00",X"09",X"62",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"29",
		X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"99",X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"99",
		X"00",X"00",X"22",X"29",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"72",
		X"00",X"00",X"76",X"22",X"00",X"00",X"27",X"99",X"00",X"00",X"22",X"96",X"00",X"00",X"22",X"69",
		X"00",X"00",X"22",X"99",X"00",X"00",X"92",X"99",X"00",X"00",X"96",X"99",X"00",X"00",X"92",X"99",
		X"00",X"00",X"92",X"99",X"00",X"00",X"92",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"76",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"92",X"00",X"00",X"00",
		X"92",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"69",X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"66",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9E",
		X"00",X"00",X"00",X"9E",X"00",X"00",X"09",X"9E",X"00",X"00",X"99",X"72",X"00",X"00",X"99",X"27",
		X"00",X"00",X"99",X"27",X"00",X"00",X"9E",X"67",X"00",X"00",X"EE",X"62",X"00",X"00",X"E9",X"62",
		X"00",X"00",X"E9",X"22",X"00",X"00",X"E9",X"26",X"00",X"00",X"99",X"26",X"00",X"00",X"99",X"22",
		X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"96",X"00",X"00",X"99",X"66",X"00",X"00",X"99",X"69",
		X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",
		X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"96",X"00",X"00",X"00",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"79",X"00",X"00",X"EE",X"29",X"00",X"00",X"E2",X"67",X"00",X"00",X"99",X"67",X"00",
		X"00",X"92",X"67",X"00",X"00",X"22",X"62",X"00",X"00",X"92",X"72",X"00",X"00",X"92",X"72",X"00",
		X"00",X"22",X"72",X"00",X"00",X"22",X"72",X"00",X"00",X"22",X"72",X"00",X"00",X"22",X"22",X"00",
		X"00",X"22",X"22",X"00",X"00",X"22",X"99",X"00",X"00",X"29",X"29",X"00",X"00",X"99",X"92",X"00",
		X"00",X"92",X"99",X"00",X"00",X"92",X"99",X"00",X"00",X"92",X"99",X"00",X"00",X"99",X"66",X"00",
		X"00",X"96",X"66",X"00",X"00",X"96",X"66",X"00",X"00",X"96",X"66",X"00",X"00",X"96",X"66",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"99",X"99",X"09",X"00",X"22",X"99",X"09",X"00",X"99",X"99",X"09",X"00",
		X"99",X"29",X"90",X"00",X"99",X"22",X"90",X"00",X"66",X"22",X"70",X"00",X"66",X"22",X"70",X"00",
		X"66",X"92",X"99",X"00",X"66",X"92",X"99",X"00",X"66",X"92",X"99",X"00",X"66",X"92",X"99",X"00",
		X"66",X"92",X"99",X"00",X"66",X"92",X"90",X"00",X"66",X"92",X"99",X"00",X"66",X"92",X"99",X"00",
		X"66",X"22",X"99",X"00",X"66",X"22",X"79",X"00",X"99",X"22",X"00",X"00",X"99",X"22",X"00",X"00",
		X"22",X"99",X"09",X"00",X"99",X"99",X"09",X"00",X"99",X"99",X"09",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"92",X"90",X"00",X"66",X"99",X"20",X"00",X"66",X"92",X"20",X"00",X"66",X"92",X"22",X"00",
		X"66",X"92",X"00",X"00",X"66",X"22",X"09",X"00",X"29",X"29",X"99",X"00",X"92",X"29",X"99",X"00",
		X"99",X"92",X"99",X"00",X"22",X"22",X"99",X"00",X"99",X"22",X"00",X"00",X"99",X"22",X"00",X"00",
		X"09",X"22",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"22",X"00",X"00",
		X"00",X"92",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"26",X"99",X"00",X"00",X"92",X"96",X"00",X"00",X"92",X"26",X"00",X"00",X"99",X"99",
		X"00",X"00",X"99",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"20",X"00",X"00",X"66",X"92",X"00",X"00",X"66",X"22",X"00",X"00",X"66",X"92",X"00",X"00",
		X"66",X"22",X"00",X"00",X"69",X"22",X"00",X"00",X"99",X"22",X"90",X"00",X"99",X"22",X"90",X"00",
		X"99",X"22",X"90",X"00",X"99",X"92",X"90",X"00",X"99",X"22",X"00",X"00",X"99",X"22",X"09",X"00",
		X"29",X"77",X"99",X"00",X"22",X"79",X"99",X"00",X"92",X"99",X"90",X"00",X"99",X"99",X"90",X"00",
		X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",
		X"66",X"00",X"00",X"00",X"66",X"99",X"00",X"00",X"79",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"22",X"27",X"00",X"00",X"29",X"92",X"00",X"00",X"92",X"92",X"00",X"00",
		X"22",X"97",X"00",X"00",X"22",X"22",X"00",X"00",X"29",X"22",X"00",X"00",X"99",X"79",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"79",X"90",X"00",X"00",
		X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"96",X"00",X"00",X"00",X"96",
		X"00",X"00",X"00",X"96",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",
		X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"96",X"66",X"00",X"00",X"96",X"66",X"00",X"00",X"96",X"66",X"00",X"00",X"96",X"66",X"00",
		X"00",X"96",X"62",X"00",X"00",X"96",X"62",X"00",X"00",X"92",X"99",X"00",X"00",X"92",X"99",X"00",
		X"00",X"27",X"99",X"00",X"00",X"29",X"99",X"00",X"00",X"29",X"99",X"00",X"00",X"72",X"99",X"90",
		X"00",X"27",X"92",X"90",X"00",X"22",X"22",X"90",X"00",X"29",X"99",X"90",X"00",X"96",X"22",X"90",
		X"00",X"96",X"22",X"90",X"00",X"96",X"22",X"90",X"00",X"22",X"22",X"90",X"00",X"27",X"22",X"90",
		X"00",X"97",X"77",X"00",X"00",X"69",X"77",X"00",X"00",X"79",X"97",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"90",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"00",X"00",
		X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",
		X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",
		X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",
		X"22",X"22",X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",
		X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"20",X"00",X"00",X"20",X"00",
		X"00",X"00",X"22",X"09",X"00",X"02",X"22",X"99",X"00",X"26",X"22",X"90",X"00",X"62",X"62",X"00",
		X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"29",X"00",X"00",X"92",X"90",X"00",
		X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"99",
		X"00",X"02",X"22",X"99",X"00",X"22",X"22",X"00",X"00",X"22",X"00",X"00",X"00",X"99",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"11",X"15",X"00",X"00",X"11",X"41",
		X"00",X"00",X"44",X"45",X"00",X"00",X"45",X"95",X"00",X"00",X"55",X"19",X"00",X"00",X"11",X"59",
		X"00",X"00",X"14",X"59",X"00",X"00",X"14",X"99",X"00",X"00",X"14",X"99",X"00",X"00",X"51",X"99",
		X"00",X"00",X"99",X"99",X"00",X"00",X"54",X"99",X"00",X"00",X"14",X"99",X"00",X"00",X"11",X"99",
		X"00",X"00",X"14",X"99",X"00",X"00",X"11",X"59",X"00",X"00",X"99",X"59",X"00",X"00",X"45",X"99",
		X"00",X"00",X"11",X"45",X"00",X"00",X"51",X"11",X"00",X"00",X"99",X"99",X"00",X"00",X"09",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"99",X"00",X"99",X"99",X"91",X"00",X"55",X"15",X"11",X"00",X"55",X"55",X"59",X"00",
		X"99",X"99",X"55",X"00",X"99",X"99",X"55",X"00",X"99",X"59",X"95",X"00",X"11",X"14",X"95",X"00",
		X"44",X"44",X"95",X"00",X"44",X"44",X"95",X"00",X"44",X"44",X"95",X"00",X"44",X"44",X"95",X"00",
		X"44",X"44",X"95",X"00",X"44",X"44",X"95",X"00",X"44",X"44",X"95",X"00",X"44",X"44",X"95",X"00",
		X"44",X"44",X"95",X"00",X"44",X"44",X"95",X"00",X"99",X"99",X"95",X"00",X"99",X"99",X"55",X"00",
		X"99",X"99",X"55",X"00",X"55",X"95",X"49",X"00",X"99",X"99",X"11",X"00",X"00",X"99",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"95",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"9E",X"90",X"00",X"00",X"5E",X"99",
		X"00",X"00",X"13",X"15",X"00",X"00",X"59",X"41",X"00",X"00",X"55",X"44",X"00",X"00",X"51",X"95",
		X"00",X"00",X"51",X"15",X"00",X"00",X"11",X"44",X"00",X"00",X"59",X"41",X"00",X"00",X"59",X"45",
		X"00",X"00",X"55",X"59",X"00",X"00",X"94",X"99",X"00",X"00",X"94",X"59",X"00",X"00",X"44",X"99",
		X"00",X"00",X"51",X"99",X"00",X"00",X"51",X"99",X"00",X"00",X"55",X"99",X"00",X"00",X"45",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"59",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"99",X"90",X"00",X"00",
		X"99",X"59",X"00",X"00",X"45",X"51",X"00",X"00",X"41",X"91",X"00",X"00",X"44",X"99",X"99",X"00",
		X"44",X"99",X"55",X"00",X"44",X"15",X"14",X"00",X"44",X"44",X"14",X"00",X"44",X"44",X"99",X"00",
		X"00",X"00",X"14",X"99",X"00",X"00",X"55",X"95",X"00",X"00",X"95",X"19",X"00",X"00",X"99",X"55",
		X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"44",X"91",X"00",X"44",X"44",X"91",X"00",X"44",X"44",X"55",X"00",X"44",X"44",X"15",X"00",
		X"44",X"44",X"15",X"00",X"54",X"44",X"19",X"00",X"91",X"44",X"59",X"00",X"94",X"44",X"90",X"00",
		X"54",X"44",X"90",X"00",X"91",X"54",X"90",X"00",X"91",X"99",X"00",X"00",X"09",X"99",X"00",X"00",
		X"00",X"49",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"55",
		X"00",X"00",X"09",X"15",X"00",X"00",X"09",X"41",X"00",X"00",X"95",X"44",X"00",X"00",X"54",X"14",
		X"00",X"00",X"45",X"91",X"00",X"00",X"95",X"19",X"00",X"00",X"91",X"45",X"00",X"00",X"54",X"44",
		X"00",X"00",X"59",X"44",X"00",X"00",X"45",X"44",X"00",X"00",X"14",X"44",X"00",X"00",X"54",X"45",
		X"00",X"00",X"51",X"99",X"00",X"00",X"95",X"99",X"00",X"00",X"55",X"99",X"00",X"00",X"45",X"99",
		X"00",X"00",X"14",X"99",X"00",X"00",X"54",X"95",X"00",X"00",X"51",X"95",X"00",X"00",X"95",X"51",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"51",X"00",X"00",X"00",
		X"95",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"59",X"00",X"00",X"00",
		X"49",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"59",X"00",X"00",
		X"00",X"00",X"09",X"11",X"00",X"00",X"00",X"14",X"00",X"00",X"00",X"94",X"00",X"00",X"00",X"95",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"15",
		X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"55",X"00",X"00",X"44",X"91",X"00",X"00",X"44",X"95",X"00",X"00",X"44",X"99",X"00",X"00",
		X"44",X"99",X"00",X"00",X"44",X"59",X"00",X"00",X"44",X"49",X"90",X"00",X"44",X"44",X"59",X"00",
		X"44",X"44",X"59",X"00",X"44",X"44",X"59",X"00",X"44",X"44",X"99",X"00",X"54",X"45",X"00",X"00",
		X"91",X"59",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"59",X"99",X"00",X"00",
		X"55",X"94",X"00",X"00",X"15",X"55",X"00",X"00",X"51",X"19",X"00",X"00",X"95",X"59",X"00",X"00",
		X"99",X"90",X"00",X"00",X"09",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"55",
		X"00",X"00",X"09",X"55",X"00",X"00",X"99",X"55",X"00",X"00",X"9E",X"99",X"00",X"00",X"5E",X"59",
		X"00",X"00",X"53",X"45",X"00",X"00",X"95",X"44",X"00",X"00",X"09",X"44",X"00",X"00",X"09",X"44",
		X"00",X"00",X"09",X"44",X"00",X"00",X"09",X"44",X"00",X"00",X"00",X"41",X"00",X"00",X"00",X"44",
		X"00",X"00",X"00",X"49",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"49",X"00",X"00",X"00",
		X"59",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"15",X"00",X"00",X"00",
		X"15",X"00",X"00",X"00",X"41",X"00",X"00",X"00",X"41",X"00",X"00",X"00",X"41",X"00",X"00",X"00",
		X"54",X"00",X"00",X"00",X"94",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"55",X"00",X"00",X"00",
		X"49",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"91",X"00",X"00",X"00",
		X"91",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"44",X"00",X"00",X"00",
		X"41",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"90",X"00",X"00",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"19",
		X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"91",
		X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"90",X"00",X"00",X"44",X"90",X"00",X"00",X"44",X"90",X"00",X"00",X"44",X"19",X"00",X"00",
		X"44",X"55",X"00",X"00",X"44",X"91",X"00",X"00",X"44",X"91",X"00",X"00",X"44",X"95",X"00",X"00",
		X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",
		X"44",X"44",X"00",X"00",X"14",X"95",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",
		X"44",X"05",X"00",X"00",X"49",X"55",X"00",X"00",X"99",X"54",X"00",X"00",X"99",X"55",X"00",X"00",
		X"09",X"59",X"00",X"00",X"00",X"90",X"00",X"00",X"05",X"00",X"00",X"00",X"55",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"95",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"E9",X"49",X"00",X"00",X"E9",X"99",X"00",
		X"00",X"35",X"55",X"00",X"00",X"95",X"15",X"00",X"00",X"95",X"51",X"00",X"00",X"95",X"11",X"00",
		X"00",X"55",X"11",X"00",X"00",X"55",X"11",X"00",X"00",X"51",X"44",X"00",X"00",X"51",X"14",X"00",
		X"00",X"51",X"14",X"00",X"00",X"51",X"11",X"00",X"00",X"55",X"41",X"00",X"00",X"55",X"95",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"59",X"99",X"00",X"00",X"59",X"95",X"00",
		X"00",X"91",X"41",X"00",X"00",X"51",X"44",X"00",X"00",X"91",X"44",X"00",X"00",X"91",X"44",X"00",
		X"00",X"41",X"44",X"00",X"00",X"91",X"44",X"00",X"00",X"91",X"44",X"00",X"00",X"91",X"44",X"00",
		X"00",X"94",X"44",X"00",X"00",X"91",X"44",X"00",X"00",X"14",X"44",X"00",X"00",X"91",X"44",X"00",
		X"00",X"94",X"41",X"00",X"00",X"91",X"44",X"00",X"00",X"91",X"44",X"00",X"00",X"91",X"44",X"00",
		X"00",X"94",X"44",X"00",X"00",X"91",X"44",X"00",X"00",X"91",X"44",X"00",X"00",X"94",X"44",X"00",
		X"00",X"94",X"44",X"00",X"00",X"51",X"11",X"00",X"00",X"49",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"55",X"55",X"00",X"00",X"15",X"15",X"00",X"00",X"99",X"99",X"00",X"00",X"55",X"55",X"00",
		X"00",X"99",X"59",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"A9",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"93",X"90",X"00",X"99",X"99",X"90",X"00",X"99",X"99",X"90",X"00",
		X"99",X"00",X"99",X"00",X"9A",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"99",X"00",
		X"9A",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"99",X"00",
		X"99",X"00",X"99",X"00",X"99",X"99",X"90",X"00",X"99",X"99",X"95",X"00",X"99",X"93",X"90",X"00",
		X"99",X"33",X"05",X"00",X"99",X"99",X"50",X"00",X"09",X"99",X"05",X"00",X"00",X"99",X"50",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",
		X"00",X"00",X"05",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"50",X"00",
		X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9D",X"00",X"00",X"09",X"9D",X"00",X"00",
		X"09",X"A5",X"00",X"00",X"09",X"55",X"00",X"00",X"99",X"55",X"00",X"00",X"99",X"55",X"00",X"00",
		X"99",X"59",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"99",X"05",X"00",X"09",X"99",X"50",X"00",X"09",X"90",X"05",X"00",X"00",X"00",X"50",X"00",
		X"00",X"00",X"05",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"50",X"00",
		X"00",X"00",X"05",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"50",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"99",X"00",X"99",X"99",X"95",X"00",X"55",X"15",X"15",X"00",X"15",X"55",X"49",X"00",
		X"99",X"99",X"59",X"00",X"99",X"99",X"99",X"00",X"99",X"59",X"95",X"00",X"11",X"14",X"55",X"00",
		X"44",X"44",X"55",X"00",X"44",X"44",X"55",X"00",X"44",X"44",X"59",X"00",X"44",X"44",X"99",X"00",
		X"44",X"44",X"99",X"00",X"44",X"45",X"90",X"00",X"44",X"45",X"90",X"00",X"44",X"44",X"99",X"00",
		X"44",X"44",X"99",X"00",X"44",X"44",X"59",X"00",X"99",X"99",X"59",X"00",X"99",X"99",X"95",X"00",
		X"99",X"99",X"55",X"00",X"51",X"91",X"95",X"00",X"99",X"99",X"55",X"00",X"00",X"99",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"59",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"51",X"09",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"59",X"00",X"00",X"45",X"51",X"90",X"00",X"41",X"91",X"90",X"00",X"44",X"99",X"99",X"00",
		X"44",X"99",X"55",X"00",X"44",X"15",X"14",X"00",X"44",X"44",X"14",X"00",X"44",X"44",X"99",X"00",
		X"44",X"55",X"51",X"00",X"44",X"59",X"99",X"00",X"44",X"99",X"59",X"00",X"44",X"95",X"99",X"00",
		X"44",X"99",X"15",X"00",X"54",X"59",X"19",X"00",X"91",X"59",X"59",X"00",X"94",X"59",X"90",X"00",
		X"54",X"99",X"90",X"00",X"91",X"55",X"90",X"00",X"91",X"49",X"00",X"00",X"09",X"41",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"55",X"00",X"00",X"44",X"91",X"00",X"00",X"44",X"95",X"00",X"00",X"44",X"99",X"00",X"00",
		X"44",X"99",X"00",X"00",X"44",X"59",X"00",X"00",X"44",X"44",X"90",X"00",X"44",X"55",X"59",X"00",
		X"44",X"99",X"59",X"00",X"44",X"99",X"59",X"00",X"44",X"99",X"99",X"00",X"54",X"99",X"00",X"00",
		X"91",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"59",X"59",X"00",X"00",
		X"55",X"95",X"00",X"00",X"15",X"55",X"00",X"00",X"51",X"19",X"00",X"00",X"95",X"59",X"00",X"00",
		X"99",X"90",X"00",X"00",X"09",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"90",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"19",X"00",X"00",
		X"44",X"55",X"00",X"00",X"44",X"91",X"00",X"00",X"44",X"91",X"00",X"00",X"44",X"95",X"00",X"00",
		X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"45",X"51",X"00",X"00",X"54",X"44",X"00",X"00",
		X"45",X"54",X"00",X"00",X"59",X"95",X"00",X"00",X"99",X"95",X"00",X"00",X"99",X"55",X"00",X"00",
		X"99",X"55",X"00",X"00",X"59",X"55",X"00",X"00",X"99",X"54",X"00",X"00",X"55",X"55",X"00",X"00",
		X"55",X"59",X"00",X"00",X"95",X"90",X"00",X"00",X"95",X"00",X"00",X"00",X"55",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"19",
		X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"91",
		X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"41",X"44",X"00",X"00",X"91",X"44",X"00",X"00",X"91",X"44",X"00",X"00",X"91",X"44",X"00",
		X"00",X"94",X"44",X"00",X"00",X"91",X"44",X"00",X"00",X"14",X"44",X"00",X"00",X"91",X"44",X"00",
		X"00",X"94",X"41",X"00",X"00",X"91",X"44",X"00",X"00",X"91",X"44",X"90",X"00",X"91",X"44",X"00",
		X"00",X"94",X"45",X"90",X"00",X"91",X"54",X"00",X"00",X"91",X"54",X"00",X"00",X"19",X"95",X"00",
		X"00",X"19",X"99",X"90",X"00",X"99",X"95",X"00",X"00",X"55",X"99",X"90",X"00",X"55",X"55",X"00",
		X"00",X"95",X"55",X"00",X"00",X"99",X"55",X"00",X"00",X"99",X"99",X"00",X"00",X"55",X"55",X"00",
		X"00",X"99",X"59",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"11",X"15",X"00",X"00",X"11",X"41",
		X"00",X"00",X"44",X"45",X"00",X"00",X"45",X"55",X"00",X"00",X"55",X"19",X"00",X"00",X"99",X"59",
		X"00",X"00",X"D9",X"59",X"00",X"00",X"DD",X"99",X"00",X"00",X"9D",X"99",X"00",X"00",X"D9",X"99",
		X"00",X"00",X"D9",X"99",X"00",X"00",X"9D",X"99",X"00",X"00",X"DD",X"99",X"00",X"00",X"D9",X"99",
		X"00",X"00",X"99",X"99",X"00",X"00",X"59",X"59",X"00",X"00",X"55",X"59",X"00",X"00",X"45",X"99",
		X"00",X"00",X"11",X"45",X"00",X"00",X"51",X"11",X"00",X"00",X"99",X"99",X"00",X"00",X"09",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"95",X"90",X"00",X"00",X"9E",X"99",X"00",X"00",X"EE",X"99",X"00",X"00",X"EE",X"99",
		X"00",X"00",X"EE",X"15",X"00",X"00",X"59",X"41",X"00",X"00",X"55",X"44",X"00",X"00",X"D9",X"55",
		X"00",X"00",X"D9",X"55",X"00",X"00",X"99",X"91",X"00",X"00",X"99",X"11",X"00",X"00",X"99",X"15",
		X"00",X"00",X"D9",X"59",X"00",X"00",X"DD",X"99",X"00",X"00",X"9D",X"59",X"00",X"00",X"99",X"99",
		X"00",X"00",X"59",X"99",X"00",X"00",X"55",X"99",X"00",X"00",X"55",X"99",X"00",X"00",X"45",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"55",
		X"00",X"00",X"09",X"15",X"00",X"00",X"09",X"41",X"00",X"00",X"95",X"44",X"00",X"00",X"54",X"14",
		X"00",X"00",X"4D",X"51",X"00",X"00",X"DD",X"55",X"00",X"00",X"D9",X"95",X"00",X"00",X"99",X"99",
		X"00",X"00",X"99",X"99",X"00",X"00",X"DD",X"55",X"00",X"00",X"9D",X"51",X"00",X"00",X"99",X"15",
		X"00",X"00",X"59",X"99",X"00",X"00",X"55",X"99",X"00",X"00",X"55",X"99",X"00",X"00",X"45",X"99",
		X"00",X"00",X"14",X"99",X"00",X"00",X"54",X"95",X"00",X"00",X"51",X"95",X"00",X"00",X"95",X"51",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"49",X"00",X"00",X"00",
		X"59",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"15",X"00",X"00",X"00",
		X"15",X"00",X"00",X"00",X"41",X"00",X"00",X"00",X"41",X"00",X"00",X"00",X"41",X"00",X"00",X"00",
		X"54",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"55",X"00",X"00",X"00",
		X"49",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"91",X"00",X"00",X"00",
		X"91",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"44",X"00",X"00",X"00",
		X"41",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"90",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"DD",
		X"00",X"00",X"09",X"DD",X"00",X"00",X"99",X"99",X"00",X"00",X"9E",X"9D",X"00",X"00",X"5E",X"9D",
		X"00",X"00",X"53",X"9D",X"00",X"00",X"95",X"D9",X"00",X"00",X"09",X"D9",X"00",X"00",X"09",X"DD",
		X"00",X"00",X"09",X"9D",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"44",
		X"00",X"00",X"00",X"49",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"95",X"90",X"00",X"00",X"90",X"90",X"00",X"00",X"ED",X"99",X"00",X"00",X"E9",X"95",X"00",
		X"00",X"35",X"55",X"00",X"00",X"95",X"D9",X"00",X"00",X"95",X"D5",X"00",X"00",X"95",X"D5",X"90",
		X"00",X"59",X"D9",X"00",X"00",X"59",X"D9",X"00",X"00",X"59",X"D9",X"00",X"00",X"59",X"D9",X"90",
		X"00",X"59",X"99",X"00",X"00",X"55",X"99",X"00",X"00",X"51",X"41",X"90",X"00",X"15",X"95",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"59",X"99",X"00",X"00",X"59",X"95",X"00",
		X"00",X"91",X"41",X"00",X"00",X"51",X"44",X"00",X"00",X"91",X"44",X"00",X"00",X"91",X"44",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"11",X"15",X"00",X"00",X"11",X"41",
		X"00",X"00",X"44",X"45",X"00",X"00",X"45",X"55",X"00",X"00",X"55",X"19",X"00",X"00",X"99",X"59",
		X"00",X"00",X"D9",X"59",X"00",X"00",X"DD",X"99",X"00",X"00",X"9D",X"99",X"00",X"00",X"D9",X"99",
		X"00",X"00",X"D9",X"99",X"00",X"00",X"9D",X"99",X"00",X"00",X"DD",X"99",X"00",X"00",X"D9",X"99",
		X"00",X"00",X"99",X"99",X"00",X"00",X"59",X"59",X"00",X"00",X"55",X"59",X"00",X"00",X"45",X"99",
		X"00",X"00",X"11",X"45",X"00",X"00",X"51",X"11",X"00",X"00",X"99",X"99",X"00",X"00",X"09",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"59",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"59",X"00",X"00",X"45",X"51",X"00",X"00",X"41",X"91",X"90",X"00",X"44",X"99",X"99",X"00",
		X"44",X"99",X"55",X"00",X"44",X"15",X"14",X"00",X"44",X"44",X"14",X"00",X"44",X"44",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"95",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"EE",X"90",X"00",X"00",X"EE",X"99",
		X"00",X"00",X"E3",X"15",X"00",X"00",X"59",X"41",X"00",X"00",X"55",X"44",X"00",X"00",X"D9",X"55",
		X"00",X"00",X"D9",X"55",X"00",X"00",X"99",X"91",X"00",X"00",X"99",X"11",X"00",X"00",X"99",X"15",
		X"00",X"00",X"D9",X"59",X"00",X"00",X"DD",X"99",X"00",X"00",X"9D",X"59",X"00",X"00",X"99",X"99",
		X"00",X"00",X"59",X"99",X"00",X"00",X"55",X"99",X"00",X"00",X"55",X"99",X"00",X"00",X"45",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"55",
		X"00",X"00",X"09",X"15",X"00",X"00",X"09",X"41",X"00",X"00",X"95",X"44",X"00",X"00",X"54",X"14",
		X"00",X"00",X"4D",X"51",X"00",X"00",X"DD",X"55",X"00",X"00",X"D9",X"95",X"00",X"00",X"99",X"99",
		X"00",X"00",X"99",X"99",X"00",X"00",X"DD",X"55",X"00",X"00",X"9D",X"51",X"00",X"00",X"99",X"15",
		X"00",X"00",X"59",X"99",X"00",X"00",X"55",X"99",X"00",X"00",X"55",X"99",X"00",X"00",X"45",X"99",
		X"00",X"00",X"14",X"99",X"00",X"00",X"54",X"95",X"00",X"00",X"51",X"95",X"00",X"00",X"95",X"51",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"49",X"00",X"00",X"00",
		X"59",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"15",X"00",X"00",X"00",
		X"15",X"00",X"00",X"00",X"41",X"00",X"00",X"00",X"41",X"00",X"00",X"00",X"41",X"00",X"00",X"00",
		X"54",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"55",X"00",X"00",X"00",
		X"49",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"91",X"00",X"00",X"00",
		X"91",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"44",X"00",X"00",X"00",
		X"41",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"90",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"DD",
		X"00",X"00",X"09",X"DD",X"00",X"00",X"99",X"99",X"00",X"00",X"95",X"9D",X"00",X"00",X"5E",X"9D",
		X"00",X"00",X"5E",X"9D",X"00",X"00",X"95",X"D9",X"00",X"00",X"09",X"D9",X"00",X"00",X"09",X"DD",
		X"00",X"00",X"09",X"9D",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"91",X"00",X"00",X"09",X"44",
		X"00",X"00",X"09",X"49",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"95",X"90",X"00",X"00",X"90",X"90",X"00",X"00",X"9D",X"99",X"00",X"00",X"E9",X"95",X"00",
		X"00",X"35",X"55",X"00",X"00",X"95",X"D9",X"00",X"00",X"95",X"D5",X"00",X"00",X"95",X"D5",X"00",
		X"00",X"59",X"D9",X"00",X"00",X"59",X"D9",X"00",X"00",X"59",X"D9",X"00",X"00",X"59",X"D9",X"00",
		X"00",X"59",X"99",X"00",X"00",X"55",X"99",X"00",X"00",X"51",X"41",X"00",X"00",X"15",X"95",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"59",X"99",X"00",X"00",X"59",X"95",X"00",
		X"00",X"91",X"41",X"00",X"00",X"51",X"44",X"00",X"00",X"91",X"44",X"00",X"00",X"91",X"44",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"99",X"00",X"99",X"99",X"95",X"00",X"55",X"15",X"15",X"00",X"15",X"55",X"49",X"00",
		X"99",X"99",X"59",X"00",X"99",X"99",X"99",X"00",X"99",X"59",X"95",X"00",X"11",X"14",X"55",X"00",
		X"44",X"44",X"55",X"00",X"44",X"44",X"55",X"00",X"44",X"44",X"59",X"00",X"44",X"44",X"99",X"00",
		X"44",X"44",X"99",X"00",X"44",X"45",X"90",X"00",X"44",X"45",X"90",X"00",X"44",X"44",X"99",X"00",
		X"44",X"44",X"99",X"00",X"44",X"44",X"59",X"00",X"99",X"99",X"59",X"00",X"99",X"99",X"95",X"00",
		X"99",X"99",X"55",X"00",X"51",X"91",X"95",X"00",X"99",X"99",X"55",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"55",X"51",X"00",X"44",X"59",X"99",X"00",X"44",X"99",X"59",X"00",X"44",X"95",X"99",X"00",
		X"44",X"99",X"15",X"00",X"54",X"59",X"19",X"00",X"91",X"59",X"59",X"00",X"94",X"59",X"90",X"00",
		X"54",X"99",X"90",X"00",X"91",X"55",X"90",X"00",X"91",X"49",X"00",X"00",X"99",X"41",X"00",X"00",
		X"99",X"44",X"00",X"00",X"09",X"55",X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"14",X"99",X"00",X"00",X"55",X"95",X"00",X"00",X"95",X"19",X"00",X"00",X"99",X"55",
		X"00",X"00",X"99",X"11",X"00",X"00",X"99",X"55",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"55",X"00",X"00",X"44",X"91",X"00",X"00",X"44",X"95",X"00",X"00",X"44",X"99",X"00",X"00",
		X"44",X"99",X"00",X"00",X"44",X"59",X"00",X"00",X"44",X"44",X"90",X"00",X"44",X"55",X"59",X"00",
		X"44",X"99",X"59",X"00",X"44",X"99",X"59",X"00",X"44",X"99",X"99",X"00",X"54",X"99",X"00",X"00",
		X"91",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"59",X"59",X"00",X"00",
		X"55",X"95",X"00",X"00",X"15",X"55",X"00",X"00",X"51",X"19",X"00",X"00",X"95",X"59",X"00",X"00",
		X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"90",X"00",X"00",X"44",X"90",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"19",X"00",X"00",
		X"44",X"55",X"00",X"00",X"44",X"91",X"00",X"00",X"44",X"91",X"00",X"00",X"44",X"95",X"00",X"00",
		X"44",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"45",X"51",X"00",X"00",X"54",X"44",X"00",X"00",
		X"45",X"54",X"00",X"00",X"59",X"95",X"00",X"00",X"99",X"95",X"00",X"00",X"99",X"55",X"00",X"00",
		X"99",X"55",X"00",X"00",X"59",X"55",X"00",X"00",X"99",X"54",X"00",X"00",X"55",X"55",X"00",X"00",
		X"55",X"59",X"00",X"00",X"95",X"90",X"00",X"00",X"95",X"00",X"00",X"00",X"55",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"19",
		X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"91",
		X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"41",X"44",X"00",X"00",X"91",X"44",X"00",X"00",X"91",X"44",X"00",X"00",X"91",X"44",X"00",
		X"00",X"94",X"44",X"00",X"00",X"91",X"44",X"00",X"00",X"14",X"44",X"00",X"00",X"91",X"44",X"00",
		X"00",X"94",X"41",X"00",X"00",X"91",X"44",X"00",X"00",X"91",X"44",X"00",X"00",X"91",X"44",X"00",
		X"00",X"94",X"45",X"00",X"00",X"91",X"54",X"00",X"00",X"91",X"54",X"00",X"00",X"19",X"95",X"00",
		X"00",X"19",X"99",X"00",X"00",X"99",X"95",X"00",X"00",X"55",X"99",X"00",X"00",X"55",X"55",X"00",
		X"00",X"95",X"55",X"00",X"00",X"99",X"55",X"00",X"00",X"99",X"99",X"00",X"00",X"55",X"55",X"00",
		X"00",X"99",X"59",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"90",X"90",X"00",X"29",X"99",X"99",X"00",X"99",X"29",X"29",X"00",X"00",X"22",X"22",
		X"00",X"00",X"22",X"22",X"00",X"99",X"22",X"22",X"00",X"99",X"22",X"22",X"00",X"29",X"22",X"22",
		X"00",X"29",X"22",X"22",X"00",X"29",X"22",X"22",X"00",X"29",X"22",X"22",X"00",X"29",X"22",X"22",
		X"00",X"29",X"22",X"22",X"00",X"29",X"22",X"22",X"00",X"29",X"29",X"29",X"00",X"99",X"99",X"99",
		X"00",X"90",X"90",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"93",X"99",X"99",X"99",X"92",X"22",X"22",X"22",X"22",X"99",X"99",X"99",X"22",X"99",X"99",X"99",
		X"22",X"09",X"09",X"09",X"22",X"09",X"09",X"09",X"22",X"09",X"09",X"09",X"22",X"09",X"09",X"09",
		X"22",X"09",X"09",X"09",X"22",X"09",X"09",X"09",X"22",X"09",X"09",X"09",X"22",X"09",X"09",X"09",
		X"22",X"09",X"09",X"09",X"22",X"99",X"99",X"99",X"22",X"99",X"99",X"99",X"22",X"22",X"22",X"22",
		X"99",X"99",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"99",X"99",X"99",X"22",X"22",X"22",X"22",X"29",X"99",X"99",X"99",X"29",X"99",X"99",X"99",
		X"29",X"90",X"90",X"90",X"99",X"90",X"90",X"90",X"22",X"90",X"90",X"90",X"22",X"90",X"90",X"90",
		X"99",X"90",X"90",X"90",X"00",X"90",X"90",X"90",X"00",X"90",X"90",X"90",X"99",X"90",X"90",X"90",
		X"29",X"90",X"90",X"90",X"29",X"99",X"99",X"99",X"29",X"99",X"99",X"99",X"92",X"22",X"22",X"22",
		X"99",X"99",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"93",X"99",X"99",X"99",X"22",X"22",X"22",X"22",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"99",X"00",X"09",X"09",X"99",X"99",X"09",X"09",X"92",X"22",X"09",X"09",X"92",X"22",X"09",X"09",
		X"22",X"92",X"09",X"09",X"29",X"92",X"09",X"09",X"29",X"92",X"09",X"09",X"29",X"92",X"09",X"09",
		X"29",X"92",X"09",X"09",X"29",X"92",X"99",X"99",X"29",X"92",X"99",X"99",X"22",X"22",X"22",X"22",
		X"99",X"99",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"99",X"99",X"09",X"00",X"09",X"99",X"99",
		X"00",X"09",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"09",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"9A",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"09",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"A9",X"99",X"00",X"99",X"99",X"99",X"00",X"A9",X"99",X"99",X"00",X"9A",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"09",X"99",X"00",X"09",X"09",X"99",X"00",X"00",X"09",X"99",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"99",
		X"00",X"90",X"00",X"9A",X"00",X"90",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"99",X"99",X"99",X"90",X"99",X"99",X"99",X"90",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"09",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"93",X"00",X"00",X"00",X"93",X"00",X"00",X"00",X"93",X"00",X"00",X"00",X"39",X"00",X"00",
		X"00",X"39",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"99",X"00",X"00",
		X"09",X"90",X"05",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"50",X"00",
		X"00",X"00",X"05",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"50",X"00",
		X"00",X"00",X"05",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"50",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"55",X"11",X"00",X"00",X"44",X"49",
		X"00",X"00",X"11",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"41",X"99",X"00",X"00",X"99",X"99",
		X"00",X"00",X"55",X"99",X"00",X"00",X"11",X"99",X"00",X"00",X"11",X"99",X"00",X"00",X"44",X"99",
		X"00",X"00",X"55",X"99",X"00",X"00",X"11",X"99",X"00",X"00",X"14",X"99",X"00",X"00",X"51",X"99",
		X"00",X"00",X"95",X"99",X"00",X"00",X"59",X"99",X"00",X"00",X"11",X"99",X"00",X"00",X"11",X"99",
		X"00",X"00",X"41",X"99",X"00",X"00",X"14",X"49",X"00",X"00",X"99",X"55",X"00",X"00",X"99",X"99",
		X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"09",X"00",X"00",X"99",X"95",X"00",X"99",X"14",X"99",X"00",X"15",X"11",X"99",X"00",
		X"99",X"55",X"95",X"00",X"99",X"44",X"94",X"00",X"99",X"44",X"91",X"00",X"44",X"91",X"91",X"00",
		X"44",X"91",X"95",X"00",X"44",X"91",X"55",X"00",X"44",X"91",X"55",X"00",X"44",X"94",X"55",X"00",
		X"44",X"91",X"59",X"00",X"44",X"94",X"59",X"00",X"44",X"94",X"59",X"00",X"44",X"94",X"55",X"00",
		X"44",X"91",X"94",X"00",X"44",X"51",X"94",X"00",X"99",X"44",X"94",X"00",X"99",X"11",X"54",X"00",
		X"99",X"55",X"95",X"00",X"51",X"44",X"99",X"00",X"99",X"11",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"9E",X"90",X"00",X"00",X"5E",X"99",
		X"00",X"00",X"EE",X"99",X"00",X"00",X"5E",X"44",X"00",X"00",X"99",X"44",X"00",X"00",X"95",X"14",
		X"00",X"00",X"99",X"99",X"00",X"00",X"55",X"51",X"00",X"00",X"11",X"11",X"00",X"00",X"59",X"44",
		X"00",X"00",X"45",X"14",X"00",X"00",X"15",X"49",X"00",X"00",X"51",X"49",X"00",X"00",X"95",X"59",
		X"00",X"00",X"59",X"99",X"00",X"00",X"45",X"99",X"00",X"00",X"14",X"99",X"00",X"00",X"41",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"95",X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"55",X"00",X"00",X"99",X"99",X"00",X"00",X"44",X"51",X"00",X"00",X"44",X"95",X"90",X"00",
		X"44",X"94",X"59",X"00",X"44",X"14",X"41",X"00",X"44",X"44",X"44",X"00",X"44",X"15",X"44",X"00",
		X"00",X"00",X"11",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"95",X"99",X"00",X"00",X"99",X"91",
		X"00",X"00",X"09",X"55",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"99",X"91",X"00",X"44",X"99",X"59",X"00",X"44",X"99",X"59",X"00",X"44",X"95",X"19",X"00",
		X"44",X"91",X"59",X"00",X"44",X"94",X"59",X"00",X"94",X"54",X"55",X"00",X"94",X"14",X"55",X"00",
		X"94",X"44",X"95",X"00",X"14",X"44",X"95",X"00",X"54",X"44",X"55",X"00",X"09",X"99",X"15",X"00",
		X"00",X"55",X"59",X"00",X"00",X"44",X"55",X"00",X"00",X"44",X"50",X"00",X"00",X"51",X"90",X"00",
		X"00",X"95",X"50",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",
		X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"39",X"00",X"00",X"05",X"49",
		X"00",X"00",X"59",X"44",X"00",X"00",X"95",X"14",X"00",X"00",X"95",X"44",X"00",X"00",X"59",X"44",
		X"00",X"00",X"99",X"94",X"00",X"00",X"91",X"99",X"00",X"00",X"91",X"11",X"00",X"00",X"91",X"41",
		X"00",X"00",X"95",X"44",X"00",X"00",X"59",X"41",X"00",X"00",X"49",X"44",X"00",X"00",X"49",X"45",
		X"00",X"00",X"15",X"59",X"00",X"00",X"14",X"99",X"00",X"00",X"14",X"99",X"00",X"00",X"14",X"99",
		X"00",X"00",X"14",X"99",X"00",X"00",X"94",X"95",X"00",X"00",X"95",X"94",X"00",X"00",X"99",X"54",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"59",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"11",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"49",X"00",X"00",X"00",
		X"45",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"19",X"00",X"00",
		X"00",X"00",X"05",X"14",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"95",
		X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"54",X"00",X"00",X"44",X"94",X"00",X"00",X"44",X"49",X"00",X"00",X"44",X"45",X"00",X"00",
		X"44",X"44",X"00",X"00",X"44",X"14",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"44",X"50",X"00",
		X"44",X"44",X"99",X"00",X"41",X"44",X"95",X"00",X"45",X"45",X"95",X"00",X"45",X"49",X"59",X"00",
		X"44",X"55",X"50",X"00",X"54",X"91",X"90",X"00",X"51",X"55",X"00",X"00",X"15",X"15",X"00",X"00",
		X"45",X"55",X"00",X"00",X"14",X"59",X"00",X"00",X"91",X"95",X"00",X"00",X"95",X"11",X"00",X"00",
		X"59",X"45",X"00",X"00",X"09",X"59",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"50",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"55",
		X"00",X"00",X"00",X"59",X"00",X"00",X"05",X"99",X"00",X"00",X"99",X"15",X"00",X"00",X"99",X"94",
		X"00",X"00",X"5E",X"99",X"00",X"00",X"5E",X"11",X"00",X"00",X"93",X"41",X"00",X"00",X"91",X"45",
		X"00",X"00",X"91",X"41",X"00",X"00",X"95",X"44",X"00",X"00",X"99",X"14",X"00",X"00",X"59",X"44",
		X"00",X"00",X"09",X"44",X"00",X"00",X"09",X"44",X"00",X"00",X"09",X"45",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"95",
		X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"14",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"50",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"19",X"00",X"00",X"00",
		X"49",X"00",X"00",X"00",X"45",X"00",X"00",X"00",X"14",X"00",X"00",X"00",X"44",X"00",X"00",X"00",
		X"44",X"00",X"00",X"00",X"94",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"19",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"91",X"00",X"00",X"00",
		X"45",X"00",X"00",X"00",X"41",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",
		X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"19",
		X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"94",
		X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"05",
		X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"90",X"00",X"00",X"44",X"59",X"00",X"00",
		X"44",X"45",X"00",X"00",X"44",X"45",X"00",X"00",X"44",X"14",X"00",X"00",X"59",X"54",X"00",X"00",
		X"99",X"54",X"00",X"00",X"99",X"54",X"00",X"00",X"99",X"94",X"00",X"00",X"54",X"94",X"00",X"00",
		X"44",X"94",X"00",X"00",X"44",X"55",X"00",X"00",X"44",X"59",X"00",X"00",X"44",X"59",X"00",X"00",
		X"99",X"59",X"00",X"00",X"55",X"99",X"00",X"00",X"15",X"14",X"00",X"00",X"55",X"55",X"00",X"00",
		X"55",X"55",X"00",X"00",X"99",X"50",X"00",X"00",X"44",X"00",X"00",X"00",X"55",X"00",X"00",X"00",
		X"59",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"95",X"99",X"00",X"00",X"E5",X"59",X"00",
		X"00",X"EE",X"99",X"00",X"00",X"E9",X"99",X"00",X"00",X"33",X"95",X"00",X"00",X"44",X"95",X"00",
		X"00",X"44",X"59",X"00",X"00",X"41",X"19",X"00",X"00",X"49",X"49",X"00",X"00",X"49",X"45",X"00",
		X"00",X"19",X"41",X"00",X"00",X"59",X"41",X"00",X"00",X"95",X"44",X"00",X"00",X"95",X"41",X"00",
		X"00",X"91",X"44",X"00",X"00",X"94",X"54",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"55",X"41",X"00",X"00",X"55",X"14",X"00",
		X"00",X"91",X"44",X"00",X"00",X"91",X"44",X"00",X"00",X"91",X"44",X"00",X"00",X"91",X"44",X"00",
		X"00",X"95",X"44",X"00",X"00",X"91",X"44",X"00",X"00",X"91",X"44",X"00",X"00",X"91",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"95",X"44",X"00",X"00",X"95",X"41",X"00",X"00",X"91",X"44",X"00",
		X"00",X"11",X"44",X"00",X"00",X"44",X"54",X"00",X"00",X"11",X"95",X"00",X"00",X"45",X"99",X"00",
		X"00",X"41",X"51",X"00",X"00",X"14",X"44",X"00",X"00",X"54",X"44",X"00",X"00",X"94",X"44",X"00",
		X"00",X"95",X"41",X"00",X"00",X"59",X"99",X"00",X"00",X"55",X"55",X"00",X"00",X"55",X"15",X"00",
		X"00",X"95",X"55",X"00",X"00",X"99",X"55",X"00",X"00",X"45",X"11",X"00",X"00",X"95",X"55",X"00",
		X"00",X"55",X"55",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"93",X"00",X"00",
		X"00",X"39",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"93",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"93",X"00",X"00",X"09",X"39",X"00",X"00",X"09",X"39",X"00",X"00",X"09",X"39",X"00",X"00",
		X"99",X"99",X"00",X"00",X"9A",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"93",X"99",X"00",X"00",
		X"93",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"99",X"05",X"00",X"09",X"90",X"50",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"50",X"00",
		X"00",X"00",X"05",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"50",X"00",
		X"00",X"00",X"05",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"50",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"90",X"00",X"00",X"9D",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"D9",X"90",X"00",
		X"00",X"99",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",X"93",X"05",X"00",X"00",X"39",X"50",X"00",
		X"00",X"99",X"05",X"00",X"00",X"99",X"50",X"00",X"00",X"99",X"05",X"00",X"00",X"99",X"50",X"00",
		X"00",X"00",X"05",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"09",X"00",X"00",X"99",X"95",X"00",X"99",X"14",X"99",X"00",X"15",X"11",X"99",X"00",
		X"99",X"55",X"99",X"00",X"99",X"44",X"99",X"00",X"99",X"44",X"95",X"00",X"44",X"91",X"95",X"00",
		X"44",X"91",X"95",X"00",X"44",X"91",X"99",X"00",X"44",X"91",X"99",X"00",X"44",X"94",X"99",X"00",
		X"44",X"91",X"99",X"00",X"44",X"94",X"99",X"00",X"44",X"94",X"99",X"00",X"44",X"94",X"99",X"00",
		X"44",X"91",X"99",X"00",X"44",X"51",X"99",X"00",X"99",X"44",X"95",X"00",X"99",X"11",X"59",X"00",
		X"99",X"55",X"99",X"00",X"51",X"44",X"99",X"00",X"99",X"11",X"99",X"00",X"00",X"99",X"90",X"00",
		X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"95",X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"55",X"00",X"00",X"99",X"99",X"00",X"00",X"44",X"51",X"99",X"00",X"44",X"95",X"99",X"00",
		X"44",X"94",X"59",X"00",X"44",X"14",X"51",X"00",X"44",X"44",X"45",X"00",X"44",X"15",X"54",X"00",
		X"44",X"99",X"99",X"00",X"44",X"99",X"99",X"00",X"44",X"99",X"99",X"00",X"44",X"95",X"99",X"00",
		X"44",X"91",X"99",X"00",X"44",X"94",X"99",X"00",X"94",X"54",X"99",X"00",X"94",X"14",X"59",X"00",
		X"94",X"44",X"95",X"00",X"14",X"44",X"95",X"00",X"54",X"44",X"00",X"00",X"09",X"99",X"90",X"00",
		X"00",X"55",X"90",X"00",X"00",X"44",X"95",X"00",X"00",X"44",X"50",X"00",X"00",X"55",X"90",X"00",
		X"00",X"95",X"50",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"54",X"00",X"00",X"44",X"94",X"00",X"00",X"44",X"49",X"00",X"00",X"44",X"45",X"90",X"00",
		X"44",X"44",X"90",X"00",X"44",X"14",X"90",X"00",X"44",X"44",X"90",X"00",X"44",X"44",X"50",X"00",
		X"44",X"45",X"99",X"00",X"41",X"55",X"95",X"00",X"45",X"45",X"95",X"00",X"45",X"59",X"99",X"00",
		X"44",X"59",X"50",X"00",X"54",X"99",X"90",X"00",X"51",X"99",X"00",X"00",X"15",X"99",X"00",X"00",
		X"45",X"99",X"00",X"00",X"14",X"99",X"00",X"00",X"91",X"99",X"00",X"00",X"95",X"99",X"00",X"00",
		X"59",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"50",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"99",X"00",X"00",X"44",X"59",X"00",X"00",
		X"44",X"45",X"00",X"00",X"44",X"45",X"00",X"00",X"44",X"14",X"00",X"00",X"59",X"54",X"00",X"00",
		X"99",X"54",X"00",X"00",X"99",X"54",X"00",X"00",X"99",X"94",X"00",X"00",X"54",X"94",X"00",X"00",
		X"44",X"95",X"00",X"00",X"44",X"95",X"00",X"00",X"45",X"99",X"00",X"00",X"54",X"99",X"00",X"00",
		X"49",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"59",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"19",
		X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"94",
		X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"05",
		X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"95",X"44",X"00",X"00",X"91",X"44",X"00",X"00",X"91",X"44",X"00",X"00",X"91",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"95",X"44",X"00",X"00",X"95",X"41",X"00",X"00",X"91",X"44",X"00",
		X"00",X"11",X"44",X"00",X"00",X"44",X"54",X"00",X"00",X"11",X"95",X"90",X"00",X"45",X"99",X"99",
		X"00",X"41",X"51",X"90",X"00",X"14",X"44",X"99",X"00",X"11",X"44",X"90",X"00",X"91",X"54",X"99",
		X"00",X"95",X"55",X"90",X"00",X"99",X"99",X"90",X"00",X"99",X"99",X"90",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"95",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"59",X"00",
		X"00",X"55",X"55",X"00",X"00",X"95",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"55",X"11",X"00",X"00",X"54",X"49",
		X"00",X"00",X"11",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"41",X"99",X"00",X"00",X"99",X"99",
		X"00",X"00",X"99",X"99",X"00",X"00",X"DD",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"9D",X"99",
		X"00",X"00",X"D9",X"99",X"00",X"00",X"9D",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"DD",X"99",
		X"00",X"00",X"99",X"99",X"00",X"00",X"59",X"99",X"00",X"00",X"11",X"99",X"00",X"00",X"11",X"99",
		X"00",X"00",X"41",X"99",X"00",X"00",X"14",X"49",X"00",X"00",X"99",X"55",X"00",X"00",X"99",X"99",
		X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"95",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"5E",X"99",
		X"00",X"00",X"3E",X"99",X"00",X"00",X"EE",X"44",X"00",X"00",X"99",X"44",X"00",X"00",X"95",X"14",
		X"00",X"00",X"99",X"99",X"00",X"00",X"5D",X"99",X"00",X"00",X"D9",X"91",X"00",X"00",X"D9",X"94",
		X"00",X"00",X"99",X"14",X"00",X"00",X"99",X"49",X"00",X"00",X"9D",X"49",X"00",X"00",X"99",X"59",
		X"00",X"00",X"59",X"99",X"00",X"00",X"45",X"99",X"00",X"00",X"14",X"99",X"00",X"00",X"41",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",
		X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"19",X"00",X"00",X"05",X"59",
		X"00",X"00",X"59",X"45",X"00",X"00",X"95",X"54",X"00",X"00",X"95",X"44",X"00",X"00",X"59",X"44",
		X"00",X"00",X"99",X"94",X"00",X"00",X"9D",X"99",X"00",X"00",X"D9",X"99",X"00",X"00",X"99",X"D9",
		X"00",X"00",X"9D",X"D9",X"00",X"00",X"59",X"91",X"00",X"00",X"49",X"44",X"00",X"00",X"49",X"45",
		X"00",X"00",X"15",X"59",X"00",X"00",X"14",X"99",X"00",X"00",X"14",X"99",X"00",X"00",X"14",X"99",
		X"00",X"00",X"14",X"99",X"00",X"00",X"94",X"95",X"00",X"00",X"95",X"94",X"00",X"00",X"99",X"54",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"50",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"59",X"00",X"00",X"00",
		X"49",X"00",X"00",X"00",X"45",X"00",X"00",X"00",X"14",X"00",X"00",X"00",X"44",X"00",X"00",X"00",
		X"44",X"00",X"00",X"00",X"94",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"19",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"91",X"00",X"00",X"00",
		X"45",X"00",X"00",X"00",X"41",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",
		X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"55",
		X"00",X"00",X"00",X"59",X"00",X"00",X"05",X"DD",X"00",X"00",X"99",X"99",X"00",X"00",X"9E",X"99",
		X"00",X"00",X"5E",X"99",X"00",X"00",X"55",X"DD",X"00",X"00",X"91",X"9D",X"00",X"00",X"95",X"9D",
		X"00",X"00",X"91",X"9D",X"00",X"00",X"95",X"D9",X"00",X"00",X"99",X"D9",X"00",X"00",X"59",X"99",
		X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"14",X"00",X"00",X"09",X"45",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"95",
		X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"14",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"95",X"99",X"00",X"00",X"55",X"59",X"00",
		X"00",X"EE",X"99",X"00",X"00",X"EE",X"D9",X"00",X"00",X"35",X"33",X"00",X"00",X"44",X"D5",X"90",
		X"00",X"44",X"D9",X"90",X"00",X"41",X"D9",X"90",X"00",X"49",X"D9",X"90",X"00",X"49",X"D5",X"99",
		X"00",X"19",X"D9",X"90",X"00",X"59",X"D9",X"99",X"00",X"95",X"99",X"90",X"00",X"95",X"99",X"99",
		X"00",X"99",X"11",X"00",X"00",X"94",X"54",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"55",X"41",X"00",X"00",X"55",X"14",X"00",
		X"00",X"91",X"44",X"00",X"00",X"91",X"44",X"00",X"00",X"91",X"44",X"00",X"00",X"91",X"44",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"55",X"11",X"00",X"00",X"54",X"49",
		X"00",X"00",X"11",X"99",X"00",X"00",X"44",X"99",X"00",X"00",X"41",X"99",X"00",X"00",X"99",X"99",
		X"00",X"00",X"99",X"99",X"00",X"00",X"DD",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"9D",X"99",
		X"00",X"00",X"D9",X"99",X"00",X"00",X"9D",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"DD",X"99",
		X"00",X"00",X"99",X"99",X"00",X"00",X"59",X"99",X"00",X"00",X"11",X"99",X"00",X"00",X"11",X"99",
		X"00",X"00",X"41",X"99",X"00",X"00",X"14",X"49",X"00",X"00",X"99",X"55",X"00",X"00",X"99",X"99",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"95",X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"55",X"00",X"00",X"99",X"99",X"00",X"00",X"44",X"51",X"00",X"00",X"44",X"95",X"99",X"00",
		X"44",X"94",X"59",X"00",X"44",X"14",X"51",X"00",X"44",X"44",X"45",X"00",X"44",X"15",X"54",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"5E",X"99",
		X"00",X"00",X"1E",X"99",X"00",X"00",X"5E",X"44",X"00",X"00",X"99",X"44",X"00",X"00",X"95",X"14",
		X"00",X"00",X"99",X"99",X"00",X"00",X"5D",X"99",X"00",X"00",X"D9",X"91",X"00",X"00",X"D9",X"94",
		X"00",X"00",X"99",X"14",X"00",X"00",X"99",X"49",X"00",X"00",X"9D",X"49",X"00",X"00",X"99",X"59",
		X"00",X"00",X"59",X"99",X"00",X"00",X"35",X"99",X"00",X"00",X"14",X"99",X"00",X"00",X"41",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"39",X"00",X"00",X"05",X"59",
		X"00",X"00",X"59",X"45",X"00",X"00",X"95",X"54",X"00",X"00",X"95",X"44",X"00",X"00",X"59",X"44",
		X"00",X"00",X"99",X"94",X"00",X"00",X"9D",X"99",X"00",X"00",X"D9",X"99",X"00",X"00",X"99",X"D9",
		X"00",X"00",X"9D",X"D9",X"00",X"00",X"59",X"91",X"00",X"00",X"49",X"44",X"00",X"00",X"49",X"45",
		X"00",X"00",X"15",X"59",X"00",X"00",X"14",X"99",X"00",X"00",X"14",X"99",X"00",X"00",X"14",X"99",
		X"00",X"00",X"14",X"99",X"00",X"00",X"94",X"95",X"00",X"00",X"95",X"94",X"00",X"00",X"99",X"54",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"50",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"59",X"00",X"00",X"00",
		X"49",X"00",X"00",X"00",X"45",X"00",X"00",X"00",X"14",X"00",X"00",X"00",X"44",X"00",X"00",X"00",
		X"44",X"00",X"00",X"00",X"94",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"19",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"91",X"00",X"00",X"00",
		X"45",X"00",X"00",X"00",X"41",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",
		X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"55",
		X"00",X"00",X"00",X"59",X"00",X"00",X"05",X"DD",X"00",X"00",X"99",X"99",X"00",X"00",X"93",X"99",
		X"00",X"00",X"55",X"99",X"00",X"00",X"55",X"DD",X"00",X"00",X"91",X"9D",X"00",X"00",X"95",X"9D",
		X"00",X"00",X"91",X"9D",X"00",X"00",X"95",X"D9",X"00",X"00",X"99",X"D9",X"00",X"00",X"99",X"99",
		X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"14",X"00",X"00",X"99",X"45",X"00",X"00",X"99",X"99",
		X"00",X"00",X"99",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"95",
		X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"14",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"95",X"99",X"00",X"00",X"55",X"59",X"00",
		X"00",X"E5",X"99",X"00",X"00",X"EE",X"D9",X"00",X"00",X"EE",X"95",X"00",X"00",X"33",X"D5",X"00",
		X"00",X"44",X"D9",X"00",X"00",X"41",X"D9",X"00",X"00",X"49",X"D9",X"00",X"00",X"49",X"D5",X"00",
		X"00",X"19",X"D9",X"00",X"00",X"59",X"D9",X"00",X"00",X"95",X"99",X"00",X"00",X"95",X"99",X"00",
		X"00",X"99",X"11",X"00",X"00",X"94",X"54",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"55",X"41",X"00",X"00",X"55",X"14",X"00",
		X"00",X"91",X"44",X"00",X"00",X"91",X"44",X"00",X"00",X"91",X"44",X"00",X"00",X"91",X"44",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"90",X"09",X"00",X"00",X"99",X"95",X"00",X"99",X"14",X"99",X"00",X"15",X"11",X"99",X"00",
		X"99",X"55",X"99",X"00",X"99",X"44",X"99",X"00",X"99",X"44",X"95",X"00",X"44",X"91",X"95",X"00",
		X"44",X"91",X"95",X"00",X"44",X"91",X"99",X"00",X"44",X"91",X"99",X"00",X"44",X"94",X"99",X"00",
		X"44",X"91",X"99",X"00",X"44",X"94",X"99",X"00",X"44",X"94",X"99",X"00",X"44",X"94",X"99",X"00",
		X"44",X"91",X"99",X"00",X"44",X"51",X"99",X"00",X"99",X"44",X"95",X"00",X"99",X"11",X"59",X"00",
		X"99",X"55",X"99",X"00",X"51",X"44",X"99",X"00",X"99",X"11",X"99",X"00",X"00",X"99",X"90",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"99",X"99",X"00",X"44",X"99",X"99",X"00",X"44",X"99",X"99",X"00",X"44",X"95",X"99",X"00",
		X"44",X"91",X"99",X"00",X"44",X"94",X"99",X"00",X"94",X"54",X"99",X"00",X"94",X"14",X"59",X"00",
		X"94",X"44",X"95",X"00",X"14",X"44",X"95",X"00",X"54",X"44",X"00",X"00",X"09",X"99",X"90",X"00",
		X"09",X"55",X"90",X"00",X"00",X"44",X"95",X"00",X"00",X"44",X"50",X"00",X"00",X"55",X"90",X"00",
		X"00",X"95",X"50",X"00",X"00",X"95",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"51",X"99",X"00",X"00",X"54",X"99",X"00",X"00",X"55",X"99",X"00",X"00",X"99",X"91",
		X"00",X"00",X"99",X"55",X"00",X"00",X"99",X"91",X"00",X"00",X"09",X"59",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"54",X"00",X"00",X"44",X"94",X"00",X"00",X"44",X"49",X"00",X"00",X"44",X"45",X"00",X"00",
		X"44",X"44",X"00",X"00",X"44",X"14",X"90",X"00",X"44",X"44",X"90",X"00",X"44",X"44",X"50",X"00",
		X"44",X"45",X"99",X"00",X"41",X"55",X"95",X"00",X"45",X"45",X"95",X"00",X"45",X"59",X"99",X"00",
		X"44",X"59",X"50",X"00",X"54",X"99",X"90",X"00",X"51",X"99",X"00",X"00",X"15",X"99",X"00",X"00",
		X"45",X"99",X"00",X"00",X"14",X"99",X"00",X"00",X"91",X"99",X"00",X"00",X"95",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"55",X"00",X"00",X"00",X"50",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"90",X"00",X"00",X"44",X"59",X"00",X"00",
		X"44",X"49",X"00",X"00",X"44",X"45",X"00",X"00",X"44",X"14",X"00",X"00",X"59",X"54",X"00",X"00",
		X"99",X"54",X"00",X"00",X"99",X"54",X"00",X"00",X"99",X"94",X"00",X"00",X"54",X"94",X"00",X"00",
		X"44",X"95",X"00",X"00",X"44",X"95",X"00",X"00",X"45",X"99",X"00",X"00",X"54",X"99",X"00",X"00",
		X"49",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"59",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"19",
		X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"94",
		X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"95",X"44",X"00",X"00",X"91",X"44",X"00",X"00",X"91",X"44",X"00",X"00",X"91",X"44",X"00",
		X"00",X"44",X"44",X"00",X"00",X"95",X"44",X"00",X"00",X"95",X"41",X"00",X"00",X"91",X"44",X"00",
		X"00",X"11",X"44",X"00",X"00",X"44",X"54",X"00",X"00",X"11",X"95",X"00",X"00",X"45",X"99",X"00",
		X"00",X"41",X"51",X"00",X"00",X"14",X"44",X"00",X"00",X"11",X"44",X"00",X"00",X"91",X"54",X"00",
		X"00",X"95",X"55",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"95",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"59",X"00",
		X"00",X"55",X"55",X"00",X"00",X"95",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"CC",X"00",X"00",X"C0",X"0C",X"00",X"00",X"C0",X"00",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"0C",X"00",X"09",X"99",X"CC",X"00",X"09",X"99",X"00",
		X"00",X"99",X"99",X"00",X"0C",X"9D",X"99",X"00",X"00",X"99",X"99",X"CC",X"00",X"99",X"99",X"00",
		X"00",X"9D",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"59",X"99",X"00",
		X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"99",X"C0",X"00",X"C0",X"50",X"0C",
		X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"57",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",
		X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",
		X"00",X"00",X"77",X"74",X"00",X"00",X"77",X"12",X"00",X"00",X"77",X"22",X"00",X"00",X"77",X"22",
		X"00",X"00",X"77",X"22",X"00",X"00",X"77",X"23",X"00",X"00",X"77",X"22",X"00",X"00",X"77",X"22",
		X"00",X"00",X"07",X"23",X"00",X"00",X"07",X"22",X"00",X"00",X"07",X"22",X"00",X"00",X"07",X"12",
		X"00",X"00",X"07",X"71",X"00",X"00",X"04",X"74",X"00",X"00",X"00",X"74",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"32",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"07",X"21",X"00",X"00",X"07",X"11",
		X"75",X"77",X"00",X"00",X"77",X"77",X"70",X"00",X"77",X"77",X"77",X"00",X"77",X"77",X"77",X"00",
		X"77",X"77",X"77",X"00",X"77",X"77",X"70",X"00",X"77",X"77",X"70",X"00",X"77",X"77",X"77",X"00",
		X"77",X"77",X"77",X"00",X"44",X"77",X"77",X"00",X"14",X"77",X"77",X"00",X"11",X"77",X"77",X"00",
		X"11",X"77",X"77",X"00",X"11",X"77",X"77",X"70",X"21",X"77",X"77",X"77",X"22",X"77",X"77",X"77",
		X"21",X"77",X"77",X"77",X"21",X"77",X"77",X"70",X"21",X"77",X"77",X"70",X"47",X"77",X"77",X"77",
		X"77",X"77",X"77",X"77",X"41",X"77",X"77",X"77",X"16",X"47",X"77",X"77",X"12",X"47",X"77",X"77",
		X"21",X"47",X"77",X"77",X"22",X"47",X"77",X"77",X"12",X"47",X"77",X"77",X"12",X"77",X"77",X"77",
		X"12",X"77",X"77",X"77",X"12",X"77",X"77",X"77",X"42",X"77",X"77",X"77",X"71",X"77",X"77",X"77",
		X"00",X"00",X"07",X"11",X"00",X"00",X"07",X"41",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"41",
		X"00",X"00",X"00",X"71",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",
		X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"07",
		X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"97",
		X"00",X"00",X"00",X"97",X"00",X"09",X"00",X"74",X"00",X"9B",X"99",X"74",X"00",X"BA",X"99",X"71",
		X"00",X"9A",X"B9",X"74",X"00",X"BB",X"99",X"41",X"00",X"AA",X"A9",X"74",X"00",X"BB",X"9A",X"41",
		X"09",X"BA",X"99",X"74",X"09",X"BA",X"A9",X"41",X"0A",X"BB",X"AA",X"74",X"9A",X"BB",X"AA",X"94",
		X"44",X"77",X"77",X"77",X"11",X"77",X"77",X"77",X"21",X"77",X"77",X"77",X"21",X"77",X"77",X"77",
		X"47",X"77",X"77",X"77",X"41",X"77",X"77",X"77",X"14",X"77",X"77",X"77",X"44",X"47",X"77",X"77",
		X"11",X"77",X"77",X"77",X"12",X"47",X"77",X"77",X"22",X"74",X"77",X"77",X"21",X"47",X"77",X"77",
		X"11",X"44",X"77",X"77",X"47",X"44",X"77",X"77",X"44",X"44",X"A7",X"77",X"11",X"44",X"B7",X"77",
		X"11",X"44",X"AA",X"77",X"11",X"24",X"BA",X"77",X"22",X"14",X"9A",X"77",X"22",X"24",X"BB",X"77",
		X"23",X"14",X"CC",X"44",X"32",X"22",X"BC",X"77",X"32",X"22",X"9C",X"99",X"22",X"21",X"BB",X"99",
		X"22",X"11",X"CC",X"99",X"22",X"22",X"CC",X"99",X"22",X"22",X"CB",X"A9",X"22",X"22",X"BB",X"9A",
		X"22",X"22",X"B9",X"9A",X"22",X"21",X"97",X"9A",X"22",X"12",X"77",X"99",X"22",X"24",X"99",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"9B",X"00",X"00",X"00",X"BB",
		X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"9B",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"31",X"00",X"00",X"00",X"33",
		X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"32",X"00",X"00",X"00",X"32",X"00",X"00",X"00",X"22",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"07",X"22",
		X"9A",X"BB",X"99",X"44",X"BB",X"AA",X"99",X"44",X"BB",X"AB",X"99",X"A4",X"AB",X"AA",X"99",X"A4",
		X"BB",X"BB",X"99",X"A4",X"BB",X"BA",X"99",X"A4",X"B9",X"BB",X"9A",X"A4",X"B9",X"AA",X"A9",X"A4",
		X"BB",X"AB",X"AA",X"A4",X"BB",X"BA",X"AA",X"9A",X"BA",X"AA",X"AA",X"9A",X"BB",X"AB",X"AA",X"9A",
		X"AB",X"AA",X"99",X"6A",X"9B",X"AA",X"9A",X"DA",X"9A",X"9B",X"99",X"9A",X"AA",X"AA",X"99",X"9A",
		X"A9",X"AA",X"99",X"9A",X"A9",X"BA",X"99",X"99",X"A9",X"AB",X"99",X"99",X"99",X"BA",X"99",X"79",
		X"79",X"AA",X"99",X"97",X"77",X"AA",X"99",X"79",X"77",X"99",X"A9",X"77",X"77",X"B7",X"A9",X"77",
		X"77",X"97",X"AA",X"77",X"7A",X"97",X"A9",X"77",X"7A",X"99",X"AA",X"77",X"7A",X"AA",X"AA",X"77",
		X"79",X"BC",X"AA",X"77",X"79",X"CB",X"9A",X"77",X"0A",X"CB",X"AA",X"77",X"09",X"BB",X"AA",X"77",
		X"22",X"24",X"99",X"AA",X"22",X"4A",X"9A",X"AB",X"22",X"AB",X"9A",X"AC",X"22",X"AB",X"9A",X"AB",
		X"22",X"BB",X"99",X"BC",X"21",X"BB",X"B9",X"BB",X"22",X"BA",X"B9",X"CC",X"22",X"A9",X"BB",X"CB",
		X"22",X"A9",X"BA",X"BB",X"22",X"BA",X"BA",X"BB",X"23",X"AA",X"BB",X"BB",X"23",X"AA",X"BB",X"BB",
		X"32",X"AA",X"BB",X"AA",X"32",X"AA",X"BB",X"AA",X"22",X"AA",X"BB",X"A7",X"2A",X"AA",X"BB",X"79",
		X"2A",X"AA",X"BB",X"97",X"49",X"AA",X"BA",X"77",X"4A",X"AA",X"AA",X"77",X"9A",X"AA",X"AA",X"77",
		X"AA",X"AA",X"AA",X"77",X"AB",X"AA",X"AA",X"77",X"AA",X"AA",X"A9",X"79",X"BA",X"BA",X"99",X"79",
		X"BB",X"BB",X"99",X"7A",X"AB",X"BB",X"99",X"7A",X"BA",X"AB",X"97",X"9B",X"AB",X"BB",X"99",X"77",
		X"BB",X"BB",X"99",X"77",X"AB",X"BB",X"97",X"41",X"BB",X"BB",X"99",X"42",X"BB",X"BB",X"97",X"44",
		X"00",X"00",X"00",X"22",X"00",X"00",X"02",X"22",X"00",X"00",X"02",X"21",X"00",X"00",X"22",X"21",
		X"00",X"00",X"22",X"11",X"00",X"00",X"22",X"11",X"00",X"00",X"22",X"14",X"00",X"00",X"22",X"11",
		X"00",X"00",X"22",X"10",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",
		X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"22",X"00",
		X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"32",X"00",X"00",X"00",X"32",X"00",
		X"00",X"00",X"33",X"00",X"00",X"00",X"23",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",
		X"00",X"00",X"23",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"23",X"20",X"00",X"00",X"22",X"20",
		X"00",X"00",X"22",X"20",X"00",X"00",X"22",X"20",X"00",X"00",X"22",X"12",X"00",X"00",X"12",X"12",
		X"09",X"BB",X"A9",X"77",X"00",X"BB",X"99",X"97",X"00",X"BB",X"A9",X"79",X"00",X"AA",X"99",X"9A",
		X"00",X"AA",X"A9",X"99",X"00",X"AA",X"99",X"A9",X"00",X"AA",X"99",X"A9",X"00",X"9A",X"99",X"AA",
		X"00",X"99",X"99",X"AA",X"00",X"99",X"9A",X"AA",X"00",X"99",X"AA",X"99",X"0B",X"99",X"AA",X"99",
		X"0B",X"AA",X"9A",X"99",X"0B",X"9A",X"9A",X"7B",X"00",X"9A",X"99",X"7B",X"00",X"44",X"99",X"7B",
		X"00",X"47",X"A9",X"97",X"00",X"11",X"9A",X"97",X"00",X"11",X"9B",X"A7",X"00",X"21",X"BB",X"AA",
		X"00",X"12",X"49",X"97",X"00",X"12",X"77",X"A9",X"00",X"12",X"47",X"99",X"00",X"12",X"14",X"99",
		X"00",X"22",X"12",X"AB",X"00",X"12",X"24",X"AA",X"00",X"22",X"1B",X"77",X"00",X"12",X"97",X"A7",
		X"00",X"11",X"B9",X"A2",X"00",X"11",X"99",X"AA",X"00",X"12",X"44",X"BA",X"00",X"11",X"47",X"BA",
		X"BB",X"BB",X"99",X"44",X"BB",X"BB",X"99",X"44",X"BB",X"BB",X"99",X"74",X"BB",X"CB",X"79",X"44",
		X"BB",X"CB",X"99",X"74",X"BB",X"CB",X"99",X"47",X"AB",X"BB",X"99",X"74",X"BB",X"CB",X"97",X"47",
		X"9A",X"BB",X"97",X"74",X"AA",X"BA",X"97",X"47",X"AA",X"BA",X"97",X"74",X"AA",X"AB",X"77",X"44",
		X"AA",X"AA",X"77",X"74",X"AA",X"BA",X"77",X"44",X"AA",X"AA",X"77",X"44",X"99",X"99",X"79",X"41",
		X"9A",X"97",X"77",X"41",X"9B",X"79",X"79",X"11",X"BB",X"97",X"97",X"C1",X"B9",X"77",X"79",X"11",
		X"AA",X"77",X"90",X"11",X"AA",X"B7",X"70",X"11",X"BB",X"79",X"70",X"11",X"B9",X"77",X"00",X"11",
		X"99",X"77",X"00",X"11",X"77",X"77",X"00",X"12",X"77",X"77",X"00",X"22",X"44",X"77",X"00",X"22",
		X"21",X"44",X"00",X"22",X"22",X"44",X"00",X"22",X"21",X"44",X"00",X"22",X"22",X"44",X"00",X"22",
		X"00",X"00",X"12",X"12",X"00",X"00",X"11",X"21",X"00",X"00",X"01",X"12",X"00",X"00",X"01",X"21",
		X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"21",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",
		X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"22",X"9B",X"00",X"14",X"21",X"77",X"00",X"21",X"22",X"22",X"00",X"24",X"22",X"12",
		X"00",X"21",X"22",X"22",X"00",X"21",X"22",X"21",X"00",X"24",X"32",X"22",X"00",X"41",X"22",X"22",
		X"00",X"24",X"32",X"22",X"00",X"41",X"22",X"22",X"00",X"24",X"23",X"22",X"00",X"41",X"32",X"22",
		X"00",X"21",X"23",X"22",X"00",X"24",X"22",X"22",X"00",X"41",X"22",X"22",X"00",X"24",X"22",X"22",
		X"40",X"44",X"22",X"22",X"21",X"44",X"22",X"12",X"11",X"22",X"22",X"22",X"22",X"11",X"42",X"12",
		X"22",X"21",X"44",X"22",X"22",X"21",X"44",X"21",X"22",X"22",X"14",X"11",X"22",X"11",X"17",X"11",
		X"22",X"11",X"24",X"15",X"22",X"11",X"12",X"5E",X"22",X"21",X"41",X"EE",X"22",X"22",X"75",X"E5",
		X"11",X"12",X"75",X"55",X"44",X"41",X"45",X"55",X"00",X"14",X"45",X"66",X"00",X"47",X"45",X"65",
		X"22",X"14",X"00",X"22",X"22",X"11",X"00",X"12",X"22",X"21",X"00",X"12",X"22",X"11",X"00",X"22",
		X"22",X"21",X"00",X"12",X"22",X"21",X"E0",X"12",X"22",X"21",X"E0",X"12",X"22",X"21",X"EE",X"11",
		X"22",X"14",X"7E",X"41",X"33",X"11",X"57",X"01",X"32",X"11",X"75",X"04",X"32",X"17",X"75",X"00",
		X"23",X"77",X"77",X"00",X"33",X"E5",X"75",X"00",X"32",X"55",X"77",X"00",X"22",X"EE",X"57",X"00",
		X"22",X"7E",X"77",X"00",X"22",X"77",X"55",X"00",X"22",X"E7",X"57",X"00",X"22",X"5E",X"55",X"00",
		X"55",X"55",X"55",X"50",X"EE",X"5E",X"55",X"50",X"E5",X"55",X"55",X"50",X"7E",X"55",X"55",X"50",
		X"57",X"5E",X"55",X"50",X"57",X"EE",X"55",X"E5",X"77",X"E5",X"55",X"55",X"55",X"EE",X"55",X"E5",
		X"55",X"E5",X"55",X"55",X"55",X"5E",X"55",X"E5",X"55",X"EE",X"55",X"55",X"57",X"E5",X"55",X"5E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",
		X"00",X"00",X"00",X"42",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"23",
		X"00",X"00",X"00",X"32",X"00",X"00",X"00",X"32",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"01",X"22",X"00",X"00",X"12",X"21",
		X"00",X"17",X"47",X"66",X"00",X"77",X"47",X"77",X"00",X"17",X"44",X"75",X"00",X"77",X"47",X"55",
		X"00",X"77",X"77",X"55",X"00",X"77",X"77",X"55",X"E0",X"77",X"57",X"55",X"5E",X"54",X"75",X"55",
		X"05",X"55",X"57",X"75",X"07",X"55",X"55",X"57",X"07",X"55",X"5E",X"75",X"47",X"55",X"77",X"57",
		X"12",X"55",X"55",X"75",X"22",X"55",X"55",X"77",X"23",X"55",X"EE",X"75",X"33",X"55",X"EE",X"77",
		X"33",X"75",X"EE",X"57",X"22",X"27",X"EE",X"77",X"22",X"21",X"E5",X"75",X"22",X"21",X"E5",X"57",
		X"22",X"11",X"EE",X"77",X"22",X"21",X"5E",X"57",X"22",X"12",X"7E",X"77",X"22",X"22",X"77",X"77",
		X"22",X"22",X"11",X"75",X"22",X"22",X"11",X"77",X"22",X"22",X"11",X"77",X"22",X"22",X"17",X"77",
		X"22",X"22",X"71",X"44",X"22",X"22",X"17",X"42",X"12",X"21",X"71",X"42",X"21",X"11",X"77",X"20",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"5E",X"55",X"55",X"55",X"55",X"77",X"55",X"55",X"5E",
		X"75",X"55",X"55",X"55",X"75",X"5E",X"55",X"5E",X"55",X"5E",X"55",X"75",X"5E",X"5E",X"55",X"5E",
		X"5E",X"5E",X"55",X"75",X"EE",X"55",X"55",X"5E",X"E5",X"55",X"55",X"75",X"E5",X"5E",X"55",X"5E",
		X"E5",X"EE",X"55",X"55",X"55",X"5E",X"55",X"5E",X"55",X"55",X"55",X"75",X"E5",X"77",X"77",X"5E",
		X"55",X"51",X"C7",X"55",X"E5",X"51",X"11",X"5E",X"55",X"55",X"22",X"55",X"E7",X"72",X"22",X"55",
		X"71",X"12",X"22",X"77",X"71",X"22",X"22",X"45",X"21",X"22",X"22",X"47",X"11",X"22",X"22",X"12",
		X"21",X"22",X"22",X"41",X"11",X"22",X"22",X"12",X"21",X"22",X"22",X"41",X"12",X"22",X"22",X"12",
		X"11",X"22",X"22",X"40",X"12",X"22",X"22",X"20",X"11",X"22",X"22",X"40",X"12",X"22",X"21",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"C4",X"44",X"44",X"40",
		X"CC",X"CD",X"4D",X"00",X"CC",X"FF",X"CC",X"00",X"7C",X"BB",X"CC",X"00",X"7C",X"CC",X"DD",X"00",
		X"7C",X"CF",X"DD",X"00",X"7D",X"DC",X"DC",X"00",X"4D",X"CF",X"DC",X"00",X"4D",X"BF",X"DC",X"00",
		X"4D",X"BC",X"DC",X"00",X"7D",X"B6",X"DC",X"00",X"4D",X"CC",X"DC",X"00",X"47",X"CC",X"CC",X"00",
		X"07",X"CC",X"C7",X"00",X"07",X"CC",X"C7",X"00",X"07",X"DC",X"C7",X"00",X"00",X"DC",X"C7",X"00",
		X"00",X"DD",X"77",X"00",X"00",X"DD",X"7D",X"00",X"00",X"CD",X"DC",X"00",X"00",X"CD",X"C4",X"00",
		X"00",X"CC",X"C7",X"00",X"00",X"4C",X"97",X"00",X"00",X"44",X"77",X"00",X"00",X"C4",X"70",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"7C",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"CB",X"00",X"00",X"00",X"CD",X"00",X"00",
		X"00",X"DD",X"70",X"00",X"00",X"DC",X"77",X"00",X"00",X"DF",X"CC",X"00",X"00",X"DF",X"CC",X"00",
		X"00",X"DD",X"CC",X"00",X"00",X"DC",X"CC",X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",
		X"00",X"76",X"77",X"00",X"00",X"67",X"77",X"00",X"00",X"76",X"77",X"00",X"00",X"67",X"77",X"00",
		X"00",X"76",X"77",X"00",X"00",X"67",X"77",X"00",X"00",X"76",X"77",X"00",X"00",X"67",X"77",X"00",
		X"00",X"76",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"57",X"77",X"00",
		X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"70",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"9A",X"BB",X"99",X"44",X"BB",X"AA",X"99",X"44",X"BB",X"AB",X"99",X"A4",X"AB",X"AA",X"99",X"A4",
		X"BB",X"BB",X"99",X"A4",X"BB",X"BA",X"99",X"A4",X"B9",X"BB",X"9A",X"A4",X"B9",X"AA",X"A9",X"A4",
		X"BB",X"AB",X"AA",X"A4",X"BB",X"BA",X"AA",X"9A",X"BA",X"AA",X"AA",X"9A",X"BB",X"AB",X"AA",X"9A",
		X"AB",X"AA",X"99",X"6A",X"9B",X"AA",X"9A",X"DA",X"9A",X"9B",X"99",X"9A",X"AA",X"AA",X"99",X"9A",
		X"A9",X"AA",X"99",X"9A",X"A9",X"BA",X"99",X"99",X"A9",X"AB",X"99",X"99",X"99",X"BA",X"99",X"79",
		X"79",X"AA",X"99",X"97",X"77",X"BA",X"99",X"79",X"77",X"B9",X"A9",X"77",X"77",X"BA",X"A9",X"77",
		X"77",X"AB",X"AA",X"77",X"7A",X"9B",X"A9",X"77",X"7A",X"BB",X"AA",X"77",X"7A",X"BB",X"AA",X"77",
		X"79",X"BC",X"AA",X"77",X"79",X"CB",X"9A",X"77",X"0A",X"CB",X"AA",X"77",X"09",X"BB",X"AA",X"77",
		X"BB",X"BB",X"99",X"44",X"BB",X"BB",X"99",X"44",X"BB",X"BB",X"99",X"74",X"BB",X"CB",X"99",X"44",
		X"BB",X"CB",X"99",X"74",X"BB",X"CB",X"99",X"47",X"AB",X"BB",X"99",X"74",X"BB",X"CB",X"97",X"47",
		X"9A",X"BB",X"97",X"74",X"AA",X"BA",X"97",X"47",X"AA",X"BA",X"97",X"74",X"AA",X"AB",X"77",X"44",
		X"AA",X"AA",X"77",X"74",X"AA",X"BA",X"77",X"44",X"AA",X"AA",X"77",X"44",X"99",X"99",X"79",X"41",
		X"9A",X"97",X"77",X"41",X"9B",X"79",X"79",X"11",X"BB",X"97",X"97",X"C1",X"B9",X"77",X"79",X"11",
		X"AA",X"77",X"90",X"11",X"AA",X"B7",X"70",X"11",X"BB",X"79",X"70",X"11",X"B9",X"77",X"00",X"11",
		X"99",X"77",X"00",X"11",X"77",X"77",X"00",X"12",X"77",X"77",X"00",X"22",X"44",X"77",X"00",X"22",
		X"21",X"44",X"00",X"22",X"22",X"44",X"00",X"22",X"21",X"44",X"00",X"22",X"22",X"44",X"00",X"22",
		X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"07",X"77",X"00",X"00",X"77",X"77",X"00",
		X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"70",X"00",X"74",X"77",X"77",X"00",X"71",X"77",X"70",
		X"00",X"42",X"77",X"77",X"00",X"12",X"17",X"77",X"00",X"42",X"17",X"77",X"00",X"42",X"77",X"77",
		X"00",X"74",X"77",X"77",X"00",X"76",X"77",X"77",X"00",X"41",X"41",X"77",X"00",X"12",X"21",X"77",
		X"00",X"42",X"21",X"77",X"00",X"72",X"21",X"77",X"00",X"72",X"24",X"77",X"00",X"71",X"11",X"77",
		X"00",X"77",X"24",X"77",X"00",X"77",X"27",X"77",X"00",X"07",X"17",X"77",X"00",X"07",X"77",X"77",
		X"00",X"00",X"74",X"77",X"00",X"00",X"44",X"77",X"00",X"00",X"11",X"77",X"00",X"0B",X"11",X"47",
		X"00",X"C9",X"11",X"99",X"00",X"B9",X"22",X"A9",X"99",X"99",X"21",X"A9",X"9B",X"79",X"22",X"A9",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"22",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"21",
		X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"32",
		X"00",X"00",X"00",X"32",X"00",X"00",X"00",X"32",X"00",X"00",X"00",X"32",X"00",X"00",X"00",X"23",
		X"BB",X"B7",X"22",X"77",X"BB",X"79",X"22",X"A9",X"BA",X"9A",X"22",X"99",X"BA",X"99",X"22",X"BB",
		X"9A",X"A9",X"24",X"BB",X"99",X"99",X"2B",X"BA",X"A4",X"99",X"4B",X"AA",X"A4",X"99",X"AA",X"AB",
		X"A9",X"99",X"AB",X"BB",X"99",X"99",X"BA",X"AA",X"79",X"9A",X"BA",X"AA",X"79",X"99",X"AA",X"99",
		X"0A",X"99",X"BA",X"77",X"0A",X"99",X"AA",X"77",X"0A",X"AA",X"BB",X"77",X"0A",X"AA",X"BB",X"97",
		X"09",X"AA",X"AA",X"77",X"09",X"AA",X"AA",X"97",X"09",X"99",X"AC",X"97",X"07",X"99",X"AA",X"77",
		X"00",X"9A",X"9A",X"97",X"00",X"AA",X"A9",X"77",X"00",X"AB",X"99",X"77",X"00",X"AB",X"9A",X"77",
		X"00",X"9B",X"99",X"70",X"00",X"9A",X"99",X"70",X"00",X"B9",X"AA",X"00",X"00",X"9A",X"BB",X"00",
		X"00",X"7B",X"97",X"00",X"00",X"7B",X"77",X"00",X"00",X"77",X"22",X"00",X"00",X"42",X"21",X"00",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"02",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"22",
		X"00",X"12",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"12",X"22",X"00",
		X"00",X"22",X"21",X"50",X"00",X"22",X"31",X"E0",X"00",X"22",X"21",X"50",X"00",X"22",X"17",X"75",
		X"00",X"22",X"75",X"75",X"22",X"12",X"55",X"57",X"22",X"77",X"57",X"57",X"21",X"55",X"55",X"55",
		X"22",X"44",X"E5",X"55",X"22",X"47",X"55",X"55",X"12",X"55",X"57",X"55",X"02",X"E7",X"55",X"55",
		X"00",X"57",X"55",X"55",X"00",X"55",X"75",X"55",X"04",X"55",X"55",X"55",X"05",X"55",X"55",X"55",
		X"E5",X"55",X"55",X"55",X"75",X"E5",X"55",X"55",X"24",X"57",X"55",X"55",X"3E",X"EE",X"55",X"55",
		X"22",X"EE",X"55",X"77",X"22",X"55",X"77",X"11",X"22",X"55",X"22",X"21",X"21",X"E5",X"22",X"22",
		X"22",X"77",X"22",X"22",X"21",X"44",X"12",X"21",X"22",X"74",X"12",X"21",X"22",X"41",X"12",X"11",
		X"00",X"FF",X"00",X"DD",X"00",X"00",X"00",X"D0",X"06",X"00",X"00",X"D0",X"6F",X"00",X"00",X"D0",
		X"F0",X"00",X"00",X"DD",X"F0",X"F0",X"00",X"DD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"0D",X"00",X"FF",X"00",X"DD",X"00",X"F0",X"00",X"00",
		X"F0",X"00",X"00",X"00",X"F0",X"00",X"DD",X"0D",X"FF",X"00",X"0D",X"DD",X"6F",X"00",X"0D",X"D0",
		X"06",X"00",X"0D",X"D0",X"00",X"FF",X"0D",X"DD",X"00",X"00",X"0D",X"D0",X"00",X"00",X"0D",X"D0",
		X"00",X"00",X"DD",X"D0",X"00",X"00",X"DD",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0D",X"00",X"00",X"00",X"0D",X"00",X"D0",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0D",
		X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"D0",X"00",X"0D",X"00",X"00",
		X"DD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",
		X"DD",X"00",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"0D",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"D0",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"0D",X"00",X"00",
		X"D0",X"DD",X"00",X"00",X"D0",X"DD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0D",X"00",X"00",X"00",X"D0",X"00",X"00",X"D0",X"D0",X"00",X"00",X"0D",X"00",X"0D",X"00",
		X"0D",X"00",X"D0",X"00",X"00",X"DD",X"D0",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"D0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"00",
		X"00",X"33",X"33",X"00",X"00",X"31",X"31",X"00",X"00",X"31",X"31",X"00",X"00",X"31",X"31",X"00",
		X"00",X"31",X"31",X"00",X"00",X"31",X"31",X"00",X"00",X"31",X"31",X"00",X"00",X"31",X"31",X"00",
		X"00",X"33",X"33",X"00",X"00",X"33",X"03",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"33",X"00",X"00",X"33",X"33",X"30",
		X"00",X"13",X"33",X"33",X"00",X"13",X"00",X"13",X"00",X"13",X"30",X"13",X"00",X"13",X"33",X"13",
		X"00",X"33",X"13",X"13",X"00",X"33",X"13",X"13",X"00",X"30",X"13",X"13",X"00",X"33",X"13",X"13",
		X"00",X"33",X"33",X"33",X"00",X"13",X"30",X"30",X"00",X"33",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"30",X"30",X"30",
		X"00",X"30",X"33",X"33",X"00",X"00",X"13",X"13",X"00",X"30",X"13",X"13",X"00",X"33",X"13",X"13",
		X"00",X"13",X"13",X"13",X"00",X"13",X"13",X"13",X"00",X"13",X"13",X"13",X"00",X"13",X"13",X"13",
		X"00",X"33",X"33",X"33",X"00",X"30",X"30",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"33",X"00",X"00",X"13",X"33",X"30",
		X"00",X"13",X"33",X"33",X"00",X"13",X"00",X"13",X"00",X"13",X"30",X"13",X"00",X"13",X"33",X"13",
		X"00",X"30",X"13",X"13",X"00",X"00",X"13",X"13",X"00",X"00",X"13",X"13",X"00",X"00",X"13",X"13",
		X"00",X"00",X"33",X"33",X"00",X"00",X"30",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"33",X"33",X"33",X"03",X"13",X"13",X"13",
		X"03",X"11",X"11",X"11",X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"11",X"31",X"31",X"31",
		X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"31",
		X"31",X"11",X"11",X"11",X"11",X"13",X"13",X"13",X"33",X"33",X"33",X"33",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"33",X"33",X"33",X"03",X"11",X"11",X"11",
		X"33",X"33",X"33",X"11",X"31",X"33",X"33",X"33",X"11",X"03",X"33",X"33",X"31",X"33",X"11",X"33",
		X"31",X"31",X"33",X"33",X"31",X"11",X"03",X"33",X"31",X"13",X"03",X"33",X"31",X"13",X"33",X"33",
		X"31",X"33",X"31",X"11",X"11",X"11",X"11",X"11",X"33",X"33",X"33",X"33",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"33",X"33",X"33",X"03",X"11",X"11",X"11",
		X"03",X"33",X"11",X"11",X"31",X"33",X"33",X"33",X"31",X"33",X"33",X"33",X"11",X"11",X"33",X"33",
		X"31",X"33",X"33",X"33",X"31",X"03",X"33",X"33",X"31",X"03",X"33",X"33",X"31",X"33",X"33",X"33",
		X"31",X"31",X"11",X"11",X"11",X"11",X"11",X"11",X"33",X"33",X"33",X"33",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"00",
		X"00",X"33",X"33",X"00",X"00",X"32",X"32",X"00",X"00",X"32",X"32",X"00",X"00",X"32",X"32",X"00",
		X"00",X"32",X"32",X"00",X"00",X"32",X"32",X"00",X"00",X"32",X"32",X"00",X"00",X"32",X"32",X"00",
		X"00",X"33",X"33",X"00",X"00",X"33",X"03",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"33",X"00",X"00",X"33",X"33",X"30",
		X"00",X"23",X"33",X"33",X"00",X"23",X"00",X"23",X"00",X"23",X"30",X"23",X"00",X"23",X"33",X"23",
		X"00",X"33",X"23",X"23",X"00",X"33",X"23",X"23",X"00",X"30",X"23",X"23",X"00",X"33",X"23",X"23",
		X"00",X"33",X"33",X"33",X"00",X"23",X"30",X"30",X"00",X"33",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"30",X"30",X"30",
		X"00",X"30",X"33",X"33",X"00",X"00",X"23",X"23",X"00",X"30",X"23",X"23",X"00",X"33",X"23",X"23",
		X"00",X"23",X"23",X"23",X"00",X"23",X"23",X"23",X"00",X"23",X"23",X"23",X"00",X"23",X"23",X"23",
		X"00",X"33",X"33",X"33",X"00",X"30",X"30",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"33",X"00",X"00",X"23",X"33",X"30",
		X"00",X"23",X"33",X"33",X"00",X"23",X"00",X"23",X"00",X"23",X"30",X"23",X"00",X"23",X"33",X"23",
		X"00",X"30",X"23",X"23",X"00",X"00",X"23",X"23",X"00",X"00",X"23",X"23",X"00",X"00",X"23",X"23",
		X"00",X"00",X"33",X"33",X"00",X"00",X"30",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"33",X"33",X"33",X"03",X"23",X"23",X"23",
		X"03",X"22",X"22",X"22",X"32",X"32",X"32",X"32",X"32",X"32",X"32",X"32",X"22",X"32",X"32",X"32",
		X"32",X"32",X"32",X"32",X"32",X"32",X"32",X"32",X"32",X"32",X"32",X"32",X"32",X"32",X"32",X"32",
		X"32",X"22",X"22",X"22",X"22",X"23",X"23",X"23",X"33",X"33",X"33",X"33",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"33",X"33",X"33",X"03",X"22",X"22",X"22",
		X"33",X"33",X"33",X"22",X"32",X"33",X"33",X"33",X"22",X"03",X"33",X"33",X"32",X"33",X"22",X"33",
		X"32",X"32",X"33",X"33",X"32",X"22",X"03",X"33",X"32",X"23",X"03",X"33",X"32",X"23",X"33",X"33",
		X"32",X"33",X"32",X"22",X"22",X"22",X"22",X"22",X"33",X"33",X"33",X"33",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"33",X"33",X"33",X"03",X"22",X"22",X"22",
		X"03",X"33",X"22",X"22",X"32",X"33",X"33",X"33",X"32",X"33",X"33",X"33",X"22",X"22",X"33",X"33",
		X"32",X"33",X"33",X"33",X"32",X"03",X"33",X"33",X"32",X"03",X"33",X"33",X"32",X"33",X"33",X"33",
		X"32",X"32",X"22",X"22",X"22",X"22",X"22",X"22",X"33",X"33",X"33",X"33",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
