library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_SND_0 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_SND_0 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"C3",X"72",X"02",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"08",X"D9",X"3E",X"0E",X"D3",X"40",X"DB",X"80",
		X"B7",X"28",X"13",X"FE",X"30",X"FA",X"64",X"00",X"FE",X"40",X"F2",X"6B",X"00",X"D6",X"10",X"CD",
		X"6F",X"00",X"D9",X"08",X"FB",X"C9",X"06",X"0C",X"21",X"00",X"80",X"77",X"23",X"05",X"20",X"FB",
		X"D9",X"08",X"FB",X"C9",X"CD",X"E7",X"00",X"D9",X"08",X"FB",X"C9",X"D9",X"08",X"FB",X"C9",X"CD",
		X"A6",X"00",X"B7",X"C8",X"FE",X"01",X"28",X"15",X"FE",X"02",X"28",X"16",X"FE",X"03",X"28",X"17",
		X"FE",X"04",X"28",X"18",X"FE",X"05",X"28",X"19",X"AF",X"32",X"0A",X"80",X"C9",X"AF",X"32",X"00",
		X"80",X"C9",X"AF",X"32",X"02",X"80",X"C9",X"AF",X"32",X"04",X"80",X"C9",X"AF",X"32",X"06",X"80",
		X"C9",X"AF",X"32",X"08",X"80",X"C9",X"06",X"00",X"21",X"00",X"80",X"BE",X"28",X"1B",X"23",X"23",
		X"BE",X"28",X"1B",X"23",X"23",X"BE",X"28",X"1B",X"23",X"23",X"BE",X"28",X"1B",X"23",X"23",X"BE",
		X"28",X"1B",X"23",X"23",X"BE",X"28",X"1B",X"AF",X"C9",X"23",X"70",X"3E",X"01",X"C9",X"23",X"70",
		X"3E",X"02",X"C9",X"23",X"70",X"3E",X"03",X"C9",X"23",X"70",X"3E",X"04",X"C9",X"23",X"70",X"3E",
		X"05",X"C9",X"23",X"70",X"3E",X"06",X"C9",X"32",X"1A",X"80",X"CD",X"A6",X"00",X"B7",X"C0",X"AF",
		X"CD",X"A6",X"00",X"B7",X"20",X"73",X"3A",X"00",X"80",X"CD",X"F1",X"01",X"32",X"12",X"80",X"3A",
		X"02",X"80",X"CD",X"F1",X"01",X"32",X"13",X"80",X"3A",X"04",X"80",X"CD",X"F1",X"01",X"32",X"14",
		X"80",X"3A",X"1A",X"80",X"CD",X"F1",X"01",X"32",X"15",X"80",X"CD",X"FA",X"01",X"32",X"17",X"80",
		X"3A",X"06",X"80",X"CD",X"F1",X"01",X"32",X"12",X"80",X"3A",X"08",X"80",X"CD",X"F1",X"01",X"32",
		X"13",X"80",X"3A",X"0A",X"80",X"CD",X"F1",X"01",X"32",X"14",X"80",X"CD",X"FA",X"01",X"32",X"18",
		X"80",X"B7",X"28",X"63",X"3A",X"17",X"80",X"B7",X"28",X"79",X"3A",X"18",X"80",X"21",X"06",X"80",
		X"CD",X"E3",X"01",X"CD",X"F1",X"01",X"47",X"3A",X"17",X"80",X"21",X"00",X"80",X"CD",X"E3",X"01",
		X"CD",X"F1",X"01",X"B8",X"F2",X"C3",X"01",X"18",X"3E",X"FE",X"01",X"28",X"17",X"FE",X"02",X"28",
		X"1A",X"FE",X"03",X"28",X"1D",X"FE",X"04",X"28",X"20",X"FE",X"05",X"28",X"23",X"3A",X"1A",X"80",
		X"32",X"0A",X"80",X"C9",X"3A",X"1A",X"80",X"32",X"00",X"80",X"C9",X"3A",X"1A",X"80",X"32",X"02",
		X"80",X"C9",X"3A",X"1A",X"80",X"32",X"04",X"80",X"C9",X"3A",X"1A",X"80",X"32",X"06",X"80",X"C9",
		X"3A",X"1A",X"80",X"32",X"08",X"80",X"C9",X"3A",X"17",X"80",X"B7",X"C8",X"FE",X"01",X"28",X"09",
		X"FE",X"02",X"28",X"0A",X"21",X"04",X"80",X"18",X"18",X"21",X"00",X"80",X"18",X"13",X"21",X"02",
		X"80",X"18",X"0E",X"3A",X"18",X"80",X"FE",X"01",X"28",X"0F",X"FE",X"02",X"28",X"10",X"21",X"0A",
		X"80",X"3A",X"1A",X"80",X"77",X"23",X"36",X"00",X"C9",X"21",X"06",X"80",X"18",X"F3",X"21",X"08",
		X"80",X"18",X"EE",X"FE",X"01",X"28",X"08",X"23",X"23",X"FE",X"02",X"28",X"02",X"23",X"23",X"7E",
		X"C9",X"21",X"42",X"02",X"5F",X"16",X"00",X"19",X"7E",X"C9",X"3A",X"12",X"80",X"21",X"13",X"80",
		X"BE",X"FA",X"15",X"02",X"3A",X"14",X"80",X"BE",X"FA",X"34",X"02",X"3A",X"15",X"80",X"BE",X"FA",
		X"40",X"02",X"3E",X"02",X"C9",X"21",X"14",X"80",X"BE",X"FA",X"26",X"02",X"3A",X"15",X"80",X"BE",
		X"FA",X"32",X"02",X"3E",X"03",X"C9",X"21",X"15",X"80",X"BE",X"FA",X"2F",X"02",X"AF",X"C9",X"3E",
		X"01",X"C9",X"AF",X"C9",X"21",X"15",X"80",X"BE",X"FA",X"3D",X"02",X"AF",X"C9",X"3E",X"03",X"C9",
		X"AF",X"C9",X"00",X"01",X"02",X"03",X"04",X"05",X"06",X"07",X"08",X"09",X"0A",X"0B",X"0C",X"0D",
		X"0E",X"0F",X"10",X"11",X"12",X"13",X"14",X"15",X"16",X"17",X"18",X"19",X"1A",X"1B",X"1C",X"1D",
		X"1E",X"1F",X"20",X"21",X"22",X"23",X"24",X"25",X"26",X"27",X"28",X"29",X"2A",X"2B",X"2C",X"2D",
		X"2E",X"2F",X"06",X"00",X"21",X"00",X"80",X"70",X"23",X"7C",X"FE",X"84",X"20",X"F9",X"31",X"00",
		X"84",X"ED",X"56",X"21",X"00",X"90",X"22",X"0C",X"80",X"77",X"3E",X"07",X"D3",X"40",X"3E",X"3F",
		X"32",X"0E",X"80",X"D3",X"80",X"3E",X"07",X"D3",X"10",X"3E",X"3F",X"32",X"0F",X"80",X"D3",X"20",
		X"CD",X"2D",X"04",X"CD",X"35",X"04",X"CD",X"3D",X"04",X"CD",X"45",X"04",X"CD",X"4D",X"04",X"CD",
		X"55",X"04",X"FB",X"3E",X"0F",X"D3",X"40",X"DB",X"80",X"E6",X"80",X"20",X"F6",X"3E",X"0F",X"D3",
		X"40",X"DB",X"80",X"E6",X"80",X"28",X"F6",X"F3",X"3E",X"01",X"32",X"10",X"80",X"3A",X"01",X"80",
		X"B7",X"CA",X"4B",X"03",X"3A",X"00",X"80",X"CD",X"04",X"08",X"FB",X"00",X"00",X"F3",X"3E",X"02",
		X"32",X"10",X"80",X"3A",X"03",X"80",X"B7",X"CA",X"54",X"03",X"3A",X"02",X"80",X"CD",X"04",X"08",
		X"FB",X"00",X"00",X"F3",X"3E",X"03",X"32",X"10",X"80",X"3A",X"05",X"80",X"B7",X"CA",X"5D",X"03",
		X"3A",X"04",X"80",X"CD",X"04",X"08",X"FB",X"00",X"00",X"F3",X"3E",X"04",X"32",X"10",X"80",X"3A",
		X"07",X"80",X"B7",X"CA",X"66",X"03",X"3A",X"06",X"80",X"CD",X"04",X"08",X"FB",X"00",X"00",X"F3",
		X"3E",X"05",X"32",X"10",X"80",X"3A",X"09",X"80",X"B7",X"CA",X"6F",X"03",X"3A",X"08",X"80",X"CD",
		X"04",X"08",X"FB",X"00",X"00",X"F3",X"3E",X"06",X"32",X"10",X"80",X"3A",X"0B",X"80",X"B7",X"CA",
		X"78",X"03",X"3A",X"0A",X"80",X"CD",X"04",X"08",X"C3",X"B2",X"02",X"3A",X"00",X"80",X"CD",X"81",
		X"03",X"C3",X"DA",X"02",X"3A",X"02",X"80",X"CD",X"81",X"03",X"C3",X"F0",X"02",X"3A",X"04",X"80",
		X"CD",X"81",X"03",X"C3",X"06",X"03",X"3A",X"06",X"80",X"CD",X"81",X"03",X"C3",X"1C",X"03",X"3A",
		X"08",X"80",X"CD",X"81",X"03",X"C3",X"32",X"03",X"3A",X"0A",X"80",X"CD",X"81",X"03",X"C3",X"B2",
		X"02",X"21",X"92",X"03",X"E5",X"87",X"5F",X"16",X"00",X"21",X"CD",X"03",X"19",X"5E",X"23",X"56",
		X"EB",X"E9",X"3A",X"10",X"80",X"FE",X"01",X"28",X"16",X"FE",X"02",X"28",X"18",X"FE",X"03",X"28",
		X"1A",X"FE",X"04",X"28",X"1C",X"FE",X"05",X"28",X"1E",X"3E",X"01",X"32",X"0B",X"80",X"C9",X"3E",
		X"01",X"32",X"01",X"80",X"C9",X"3E",X"01",X"32",X"03",X"80",X"C9",X"3E",X"01",X"32",X"05",X"80",
		X"C9",X"3E",X"01",X"32",X"07",X"80",X"C9",X"3E",X"01",X"32",X"09",X"80",X"C9",X"5D",X"04",X"C0",
		X"08",X"3C",X"09",X"B8",X"09",X"34",X"0A",X"B0",X"0A",X"F9",X"0C",X"1D",X"12",X"A9",X"13",X"B9",
		X"0D",X"C7",X"0D",X"2E",X"10",X"3C",X"10",X"43",X"10",X"B2",X"10",X"C0",X"10",X"00",X"00",X"00",
		X"00",X"00",X"11",X"3C",X"0B",X"E3",X"0B",X"6D",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7A",X"0D",X"80",
		X"11",X"19",X"12",X"B6",X"12",X"34",X"13",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"08",X"D3",
		X"40",X"AF",X"D3",X"80",X"C9",X"3E",X"09",X"D3",X"40",X"AF",X"D3",X"80",X"C9",X"3E",X"0A",X"D3",
		X"40",X"AF",X"D3",X"80",X"C9",X"3E",X"08",X"D3",X"10",X"AF",X"D3",X"20",X"C9",X"3E",X"09",X"D3",
		X"10",X"AF",X"D3",X"20",X"C9",X"3E",X"0A",X"D3",X"10",X"AF",X"D3",X"20",X"C9",X"3A",X"10",X"80",
		X"FE",X"01",X"28",X"19",X"FE",X"02",X"28",X"1E",X"FE",X"03",X"28",X"23",X"FE",X"04",X"28",X"28",
		X"FE",X"05",X"28",X"2D",X"06",X"24",X"CD",X"B8",X"04",X"CD",X"55",X"04",X"C9",X"06",X"09",X"CD",
		X"AA",X"04",X"CD",X"2D",X"04",X"C9",X"06",X"12",X"CD",X"AA",X"04",X"CD",X"35",X"04",X"C9",X"06",
		X"24",X"CD",X"AA",X"04",X"CD",X"3D",X"04",X"C9",X"06",X"09",X"CD",X"B8",X"04",X"CD",X"45",X"04",
		X"C9",X"06",X"12",X"CD",X"B8",X"04",X"CD",X"4D",X"04",X"C9",X"3E",X"07",X"D3",X"40",X"3A",X"0E",
		X"80",X"B0",X"32",X"0E",X"80",X"D3",X"80",X"C9",X"3E",X"07",X"D3",X"10",X"3A",X"0F",X"80",X"B0",
		X"32",X"0F",X"80",X"D3",X"20",X"C9",X"3A",X"10",X"80",X"FE",X"01",X"28",X"20",X"FE",X"02",X"28",
		X"2C",X"FE",X"03",X"28",X"2C",X"FE",X"04",X"28",X"2C",X"FE",X"05",X"28",X"2C",X"06",X"04",X"78",
		X"D3",X"10",X"7D",X"D3",X"20",X"04",X"78",X"D3",X"10",X"7C",X"D3",X"20",X"C9",X"06",X"00",X"78",
		X"D3",X"40",X"7D",X"D3",X"80",X"04",X"78",X"D3",X"40",X"7C",X"D3",X"80",X"C9",X"06",X"02",X"18",
		X"EE",X"06",X"04",X"18",X"EA",X"06",X"00",X"18",X"D6",X"06",X"02",X"18",X"D2",X"3A",X"10",X"80",
		X"FE",X"01",X"28",X"18",X"FE",X"02",X"28",X"1C",X"FE",X"03",X"28",X"1E",X"FE",X"04",X"28",X"20",
		X"FE",X"05",X"28",X"22",X"16",X"FB",X"1E",X"20",X"CD",X"71",X"05",X"C9",X"16",X"FE",X"1E",X"08",
		X"CD",X"62",X"05",X"C9",X"16",X"FD",X"1E",X"10",X"18",X"F6",X"16",X"FB",X"1E",X"20",X"18",X"F0",
		X"16",X"FE",X"1E",X"08",X"18",X"E2",X"16",X"FD",X"1E",X"10",X"18",X"DC",X"3A",X"10",X"80",X"FE",
		X"04",X"FA",X"5B",X"05",X"7A",X"D3",X"10",X"7B",X"D3",X"20",X"C9",X"7A",X"D3",X"40",X"7B",X"D3",
		X"80",X"C9",X"3E",X"07",X"D3",X"40",X"3A",X"0E",X"80",X"A2",X"B3",X"32",X"0E",X"80",X"D3",X"80",
		X"C9",X"3E",X"07",X"D3",X"10",X"3A",X"0F",X"80",X"A2",X"B3",X"32",X"0F",X"80",X"D3",X"20",X"C9",
		X"3A",X"10",X"80",X"FE",X"01",X"28",X"18",X"FE",X"02",X"28",X"1C",X"FE",X"03",X"28",X"1E",X"FE",
		X"04",X"28",X"20",X"FE",X"05",X"28",X"22",X"16",X"DF",X"1E",X"04",X"CD",X"71",X"05",X"C9",X"16",
		X"F7",X"1E",X"01",X"CD",X"62",X"05",X"C9",X"16",X"EF",X"1E",X"02",X"18",X"F6",X"16",X"DF",X"1E",
		X"04",X"18",X"F0",X"16",X"F7",X"1E",X"01",X"18",X"E2",X"16",X"EF",X"1E",X"02",X"18",X"DC",X"3A",
		X"10",X"80",X"FE",X"01",X"28",X"18",X"FE",X"02",X"28",X"1C",X"FE",X"03",X"28",X"1E",X"FE",X"04",
		X"28",X"20",X"FE",X"05",X"28",X"22",X"16",X"DB",X"1E",X"00",X"CD",X"71",X"05",X"C9",X"16",X"F6",
		X"1E",X"00",X"CD",X"62",X"05",X"C9",X"16",X"ED",X"1E",X"00",X"18",X"F6",X"16",X"DB",X"1E",X"00",
		X"18",X"F0",X"16",X"F6",X"1E",X"00",X"18",X"E2",X"16",X"ED",X"1E",X"00",X"18",X"DC",X"3A",X"10",
		X"80",X"FE",X"01",X"28",X"18",X"FE",X"02",X"28",X"1C",X"FE",X"03",X"28",X"1C",X"FE",X"04",X"28",
		X"1C",X"FE",X"05",X"28",X"1C",X"3E",X"0A",X"D3",X"10",X"78",X"D3",X"20",X"C9",X"3E",X"08",X"D3",
		X"40",X"78",X"D3",X"80",X"C9",X"3E",X"09",X"18",X"F6",X"3E",X"0A",X"18",X"F2",X"3E",X"08",X"18",
		X"E6",X"3E",X"09",X"18",X"E2",X"3A",X"10",X"80",X"FE",X"04",X"FA",X"44",X"06",X"7A",X"D3",X"10",
		X"DB",X"20",X"5F",X"C9",X"7A",X"D3",X"40",X"DB",X"80",X"5F",X"C9",X"3A",X"10",X"80",X"FE",X"01",
		X"28",X"17",X"FE",X"02",X"28",X"1A",X"FE",X"03",X"28",X"1A",X"FE",X"04",X"28",X"1A",X"FE",X"05",
		X"28",X"1A",X"3E",X"0A",X"D3",X"10",X"DB",X"20",X"C9",X"3E",X"08",X"D3",X"40",X"DB",X"80",X"C9",
		X"3E",X"09",X"18",X"F7",X"3E",X"0A",X"18",X"F3",X"3E",X"08",X"18",X"E8",X"3E",X"09",X"18",X"E4",
		X"3A",X"10",X"80",X"FE",X"01",X"28",X"20",X"FE",X"02",X"28",X"2C",X"FE",X"03",X"28",X"2C",X"FE",
		X"04",X"28",X"2C",X"FE",X"05",X"28",X"2C",X"06",X"04",X"78",X"D3",X"10",X"DB",X"20",X"6F",X"04",
		X"78",X"D3",X"10",X"DB",X"20",X"67",X"C9",X"06",X"00",X"78",X"D3",X"40",X"DB",X"80",X"6F",X"04",
		X"78",X"D3",X"40",X"DB",X"80",X"67",X"C9",X"06",X"02",X"18",X"EE",X"06",X"04",X"18",X"EA",X"06",
		X"00",X"18",X"D6",X"06",X"02",X"18",X"D2",X"3A",X"10",X"80",X"FE",X"04",X"28",X"21",X"FE",X"05",
		X"28",X"22",X"FE",X"06",X"28",X"23",X"FE",X"01",X"28",X"24",X"FE",X"02",X"28",X"25",X"11",X"FF",
		X"F3",X"2A",X"0C",X"80",X"7A",X"A4",X"67",X"7B",X"A5",X"6F",X"22",X"0C",X"80",X"77",X"C9",X"11",
		X"FC",X"FF",X"18",X"ED",X"11",X"F3",X"FF",X"18",X"E8",X"11",X"CF",X"FF",X"18",X"E3",X"11",X"3F",
		X"FF",X"18",X"DE",X"11",X"FF",X"FC",X"18",X"D9",X"3A",X"10",X"80",X"FE",X"04",X"28",X"20",X"FE",
		X"05",X"28",X"21",X"FE",X"06",X"28",X"22",X"FE",X"01",X"28",X"23",X"FE",X"02",X"28",X"24",X"11",
		X"FF",X"F3",X"2A",X"0C",X"80",X"7A",X"A4",X"67",X"7B",X"A5",X"6F",X"22",X"0C",X"80",X"C9",X"11",
		X"FC",X"FF",X"18",X"EE",X"11",X"F3",X"FF",X"18",X"E9",X"11",X"CF",X"FF",X"18",X"E4",X"11",X"3F",
		X"FF",X"18",X"DF",X"11",X"FF",X"FC",X"18",X"DA",X"CD",X"08",X"07",X"3A",X"10",X"80",X"FE",X"04",
		X"28",X"17",X"FE",X"05",X"28",X"18",X"FE",X"06",X"28",X"19",X"FE",X"01",X"28",X"1A",X"FE",X"02",
		X"28",X"1B",X"11",X"00",X"08",X"CD",X"F6",X"07",X"C9",X"11",X"02",X"00",X"18",X"F7",X"11",X"08",
		X"00",X"18",X"F2",X"11",X"20",X"00",X"18",X"ED",X"11",X"80",X"00",X"18",X"E8",X"11",X"00",X"02",
		X"18",X"E3",X"CD",X"08",X"07",X"3A",X"10",X"80",X"FE",X"04",X"28",X"17",X"FE",X"05",X"28",X"18",
		X"FE",X"06",X"28",X"19",X"FE",X"01",X"28",X"1A",X"FE",X"02",X"28",X"1B",X"11",X"00",X"04",X"CD",
		X"F6",X"07",X"C9",X"11",X"01",X"00",X"18",X"F7",X"11",X"04",X"00",X"18",X"F2",X"11",X"10",X"00",
		X"18",X"ED",X"11",X"40",X"00",X"18",X"E8",X"11",X"00",X"01",X"18",X"E3",X"CD",X"08",X"07",X"3A",
		X"10",X"80",X"FE",X"04",X"28",X"17",X"FE",X"05",X"28",X"18",X"FE",X"06",X"28",X"19",X"FE",X"01",
		X"28",X"1A",X"FE",X"02",X"28",X"1B",X"11",X"00",X"0C",X"CD",X"F6",X"07",X"C9",X"11",X"03",X"00",
		X"18",X"F7",X"11",X"0C",X"00",X"18",X"F2",X"11",X"30",X"00",X"18",X"ED",X"11",X"C0",X"00",X"18",
		X"E8",X"11",X"00",X"03",X"18",X"E3",X"2A",X"0C",X"80",X"7A",X"B4",X"67",X"7B",X"B5",X"6F",X"22");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
