library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity swimmer_tile_bit2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of swimmer_tile_bit2 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"1C",X"1E",X"1F",X"00",X"00",X"00",X"00",X"40",X"C0",X"80",X"00",
		X"3E",X"7F",X"FF",X"FF",X"7F",X"F7",X"C7",X"88",X"00",X"C0",X"F0",X"F0",X"F0",X"80",X"00",X"00",
		X"00",X"01",X"01",X"03",X"3F",X"FF",X"FF",X"FF",X"00",X"00",X"80",X"A0",X"FC",X"F8",X"F0",X"FC",
		X"E7",X"F3",X"71",X"00",X"06",X"07",X"07",X"00",X"FE",X"F8",X"F0",X"F0",X"F0",X"F0",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"78",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"E0",X"40",X"01",X"03",X"07",X"03",X"00",X"00",X"00",X"80",X"C0",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",
		X"60",X"71",X"33",X"34",X"1E",X"0F",X"03",X"00",X"C0",X"80",X"00",X"00",X"80",X"C0",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"18",X"3C",X"39",X"3D",X"00",X"00",X"00",X"00",X"60",X"C0",X"80",X"00",
		X"1E",X"3C",X"3F",X"3F",X"3F",X"1E",X"00",X"00",X"00",X"00",X"A0",X"F0",X"F0",X"E0",X"00",X"00",
		X"02",X"02",X"00",X"07",X"03",X"01",X"01",X"00",X"00",X"00",X"50",X"90",X"38",X"FA",X"F2",X"E7",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"6F",X"3C",X"18",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"38",X"38",X"3C",X"38",X"3C",X"3C",X"00",X"00",X"00",X"00",X"10",X"30",X"60",X"C0",
		X"7D",X"FF",X"FF",X"7F",X"7F",X"FF",X"EE",X"CC",X"00",X"A0",X"F8",X"F8",X"F8",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"7B",X"44",X"78",X"40",X"40",X"00",X"00",X"00",X"EF",X"90",X"8E",X"81",X"9E",X"00",
		X"07",X"0F",X"1F",X"3E",X"3F",X"3D",X"78",X"78",X"80",X"80",X"80",X"00",X"80",X"80",X"C8",X"79",
		X"30",X"00",X"01",X"03",X"03",X"01",X"00",X"00",X"19",X"3A",X"FE",X"FC",X"F8",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"1E",X"1E",X"0E",X"00",X"40",X"40",X"C0",X"B0",X"78",X"78",X"70",
		X"00",X"00",X"00",X"19",X"0C",X"08",X"08",X"01",X"00",X"00",X"00",X"98",X"D8",X"B8",X"90",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"3C",X"66",X"66",X"66",X"66",X"66",X"3C",X"00",X"18",X"38",X"18",X"18",X"18",X"18",X"3C",
		X"00",X"3C",X"66",X"0E",X"1C",X"38",X"70",X"7E",X"00",X"3C",X"66",X"06",X"1C",X"06",X"66",X"3C",
		X"00",X"0C",X"1C",X"2C",X"6C",X"6C",X"7E",X"0C",X"00",X"7C",X"60",X"60",X"7C",X"06",X"66",X"3C",
		X"00",X"3C",X"66",X"60",X"7C",X"66",X"66",X"3C",X"00",X"7E",X"66",X"06",X"0C",X"18",X"18",X"18",
		X"00",X"3C",X"66",X"66",X"3C",X"66",X"66",X"3C",X"00",X"3C",X"66",X"66",X"3E",X"06",X"66",X"3C",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",
		X"00",X"00",X"00",X"00",X"01",X"01",X"41",X"21",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"08",
		X"11",X"08",X"00",X"00",X"00",X"F0",X"00",X"00",X"10",X"20",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"1C",X"22",X"5D",X"51",X"5D",X"22",X"1C",X"00",X"1C",X"36",X"63",X"63",X"7F",X"63",X"63",
		X"00",X"7E",X"63",X"63",X"7E",X"63",X"63",X"7E",X"00",X"3E",X"63",X"60",X"60",X"63",X"63",X"3E",
		X"00",X"7C",X"62",X"63",X"63",X"63",X"63",X"7E",X"00",X"7F",X"60",X"60",X"7E",X"60",X"60",X"7F",
		X"00",X"7F",X"60",X"60",X"7E",X"60",X"60",X"60",X"00",X"3E",X"63",X"60",X"67",X"63",X"63",X"3E",
		X"00",X"63",X"63",X"63",X"7F",X"63",X"63",X"63",X"00",X"7E",X"18",X"18",X"18",X"18",X"18",X"7E",
		X"00",X"0F",X"03",X"03",X"03",X"63",X"63",X"3E",X"00",X"63",X"66",X"6C",X"7C",X"6E",X"67",X"63",
		X"00",X"78",X"30",X"30",X"30",X"30",X"31",X"7F",X"00",X"63",X"63",X"77",X"7F",X"6B",X"63",X"63",
		X"00",X"63",X"63",X"73",X"6B",X"67",X"63",X"63",X"00",X"3E",X"63",X"63",X"63",X"63",X"63",X"3E",
		X"00",X"7E",X"63",X"63",X"7E",X"60",X"60",X"60",X"00",X"3E",X"63",X"63",X"6B",X"67",X"62",X"3D",
		X"00",X"7E",X"63",X"63",X"7E",X"7C",X"6E",X"67",X"00",X"3E",X"63",X"78",X"3E",X"0F",X"63",X"3E",
		X"00",X"7E",X"18",X"18",X"18",X"18",X"18",X"18",X"00",X"63",X"63",X"63",X"63",X"63",X"63",X"3E",
		X"00",X"63",X"63",X"63",X"63",X"36",X"1C",X"08",X"00",X"63",X"63",X"6B",X"7F",X"7F",X"77",X"63",
		X"00",X"63",X"77",X"3E",X"1C",X"3E",X"77",X"63",X"00",X"63",X"63",X"36",X"1C",X"1C",X"1C",X"1C",
		X"00",X"7E",X"46",X"0E",X"1C",X"38",X"72",X"7E",X"00",X"18",X"1C",X"1C",X"18",X"10",X"00",X"20",
		X"00",X"F0",X"60",X"60",X"60",X"60",X"62",X"FE",X"00",X"FD",X"C0",X"C0",X"F8",X"C0",X"C0",X"FC",
		X"03",X"FB",X"61",X"62",X"60",X"60",X"60",X"60",X"FF",X"81",X"81",X"81",X"81",X"81",X"81",X"FF",
		X"00",X"00",X"03",X"07",X"1C",X"3C",X"78",X"70",X"00",X"00",X"E0",X"E0",X"00",X"0C",X"1C",X"1C",
		X"78",X"F9",X"FF",X"FF",X"FF",X"7F",X"7F",X"FE",X"6C",X"CC",X"38",X"78",X"F0",X"E0",X"C0",X"00",
		X"1C",X"1E",X"0E",X"0F",X"0E",X"0F",X"1F",X"1F",X"00",X"00",X"00",X"06",X"0C",X"18",X"30",X"40",
		X"3F",X"3F",X"4F",X"9F",X"1F",X"3B",X"F6",X"00",X"E8",X"FE",X"FF",X"FF",X"C3",X"80",X"00",X"00",
		X"00",X"00",X"0F",X"3F",X"7F",X"FF",X"FF",X"1F",X"00",X"00",X"02",X"06",X"8C",X"98",X"A0",X"F0",
		X"1F",X"27",X"CF",X"8F",X"9F",X"F9",X"F3",X"F7",X"FC",X"FC",X"FC",X"F8",X"F8",X"F0",X"E0",X"C0",
		X"00",X"00",X"00",X"00",X"3C",X"3E",X"3E",X"0F",X"00",X"00",X"00",X"00",X"00",X"04",X"0C",X"18",
		X"1F",X"3F",X"3F",X"3F",X"4F",X"9F",X"1F",X"3F",X"30",X"40",X"E0",X"F8",X"FC",X"FC",X"9C",X"1C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"1E",X"00",X"00",X"00",X"40",X"40",X"C0",X"B0",X"78",
		X"3F",X"1F",X"0F",X"0C",X"04",X"00",X"05",X"0F",X"FC",X"F8",X"F0",X"F0",X"C8",X"88",X"D8",X"D8",
		X"00",X"00",X"00",X"01",X"01",X"1D",X"0F",X"0F",X"00",X"00",X"00",X"00",X"C0",X"DC",X"F8",X"F8",
		X"0F",X"3F",X"7F",X"FF",X"F8",X"F0",X"F8",X"78",X"F8",X"FC",X"FE",X"FF",X"1F",X"0F",X"1F",X"1E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"20",
		X"00",X"00",X"00",X"00",X"1D",X"3F",X"0F",X"00",X"70",X"60",X"60",X"C0",X"F8",X"FC",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"20",
		X"00",X"00",X"00",X"30",X"7D",X"7F",X"3F",X"1F",X"70",X"60",X"60",X"CC",X"FE",X"FE",X"FC",X"F8",
		X"00",X"18",X"31",X"7E",X"7E",X"3C",X"1F",X"39",X"40",X"40",X"80",X"00",X"00",X"7E",X"CC",X"DC",
		X"31",X"03",X"07",X"06",X"00",X"00",X"00",X"00",X"9C",X"FC",X"FC",X"F8",X"70",X"00",X"00",X"00",
		X"03",X"06",X"1F",X"3F",X"7F",X"FF",X"E0",X"00",X"00",X"00",X"C0",X"C0",X"C0",X"C0",X"00",X"1B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"1F",X"1F",X"1E",X"1E",X"3C",X"38",X"30",
		X"03",X"06",X"00",X"00",X"0F",X"0F",X"1F",X"1F",X"80",X"00",X"00",X"40",X"90",X"18",X"38",X"F3",
		X"3F",X"3F",X"3F",X"7F",X"7F",X"7F",X"38",X"00",X"E7",X"EF",X"FF",X"F8",X"E0",X"00",X"00",X"00",
		X"00",X"01",X"06",X"0C",X"1F",X"1F",X"1E",X"1C",X"00",X"80",X"00",X"00",X"80",X"80",X"80",X"FB",
		X"3C",X"3C",X"18",X"00",X"00",X"01",X"01",X"00",X"77",X"37",X"1F",X"3F",X"FE",X"FC",X"F8",X"C0",
		X"5F",X"7F",X"78",X"78",X"7C",X"3C",X"1C",X"1C",X"FE",X"FE",X"1E",X"1E",X"3E",X"3C",X"38",X"38",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"1C",X"1C",X"1C",X"1C",X"00",X"00",X"00",X"30",X"38",X"38",X"38",X"38",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"20",X"70",X"60",X"60",
		X"00",X"3D",X"3F",X"1F",X"07",X"07",X"03",X"00",X"C0",X"FC",X"F8",X"F8",X"E0",X"E0",X"C0",X"00",
		X"0F",X"0F",X"0F",X"1D",X"0C",X"08",X"0C",X"0D",X"F0",X"F0",X"F0",X"F8",X"D8",X"B8",X"D8",X"D8",
		X"0D",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"60",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"03",X"02",X"01",X"00",X"00",X"00",X"08",X"FF",X"DF",X"07",X"8F",
		X"01",X"03",X"02",X"01",X"00",X"00",X"00",X"00",X"FF",X"DF",X"2F",X"FF",X"F8",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"00",X"18",X"18",X"00",X"00",X"18",X"18",X"00",
		X"00",X"00",X"00",X"00",X"30",X"30",X"10",X"20",X"F8",X"20",X"20",X"20",X"11",X"1B",X"15",X"11",
		X"00",X"00",X"06",X"0E",X"0E",X"3E",X"FC",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"3E",X"0E",X"0E",X"02",X"00",X"00",X"00",X"E8",X"F0",X"20",X"00",X"00",X"00",X"00",
		X"00",X"00",X"20",X"30",X"70",X"70",X"60",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"7F",X"77",X"71",X"30",X"20",X"00",X"00",X"00",X"40",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"3E",X"FF",X"FF",X"F3",X"03",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"F3",X"FF",X"FF",X"3F",X"1F",X"00",
		X"00",X"00",X"01",X"03",X"8F",X"DF",X"87",X"C7",X"00",X"00",X"00",X"80",X"C0",X"C0",X"80",X"00",
		X"FF",X"DF",X"0F",X"CF",X"F3",X"C1",X"00",X"00",X"60",X"B8",X"C0",X"C0",X"80",X"00",X"00",X"00",
		X"78",X"FC",X"FE",X"FE",X"DF",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"20",X"E0",X"E0",X"C0",X"F8",
		X"0F",X"0F",X"0F",X"DF",X"FF",X"FE",X"FC",X"78",X"F0",X"F0",X"C0",X"E0",X"E0",X"20",X"00",X"00",
		X"00",X"00",X"00",X"1E",X"1F",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"1F",X"1F",X"1E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"06",X"0E",X"1C",X"18",X"10",X"38",X"00",X"00",X"60",X"70",X"78",X"38",X"28",X"7C",
		X"30",X"30",X"3C",X"3F",X"1F",X"1F",X"0F",X"0F",X"2C",X"6C",X"FC",X"FC",X"F8",X"F8",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"20",X"70",X"60",X"60",
		X"E0",X"FD",X"7F",X"3F",X"1F",X"0F",X"0F",X"0F",X"C7",X"FF",X"FE",X"FC",X"F8",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"00",X"40",X"20",X"70",X"20",X"20",X"40",X"B8",
		X"3F",X"7F",X"7F",X"FF",X"FF",X"EF",X"FD",X"FC",X"7C",X"FE",X"FE",X"FF",X"FF",X"F7",X"FF",X"DF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"20",X"70",X"60",X"60",
		X"00",X"7D",X"FF",X"FF",X"EF",X"0F",X"0F",X"0F",X"C0",X"FE",X"FF",X"FF",X"F7",X"F0",X"F0",X"F0",
		X"3E",X"3F",X"3F",X"07",X"01",X"00",X"00",X"00",X"00",X"F0",X"C0",X"F9",X"FF",X"7B",X"40",X"31",
		X"00",X"00",X"00",X"01",X"07",X"3F",X"3F",X"3E",X"3F",X"3B",X"45",X"FF",X"FF",X"FC",X"F0",X"00",
		X"03",X"07",X"0F",X"1E",X"FE",X"FE",X"FC",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FE",X"FE",X"1E",X"0F",X"07",X"03",X"00",X"E8",X"F0",X"20",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"07",X"1F",X"1F",X"03",X"01",X"08",X"3E",X"FF",X"FE",X"F8",X"FC",
		X"1F",X"1F",X"07",X"00",X"00",X"00",X"00",X"00",X"FF",X"FE",X"F9",X"FF",X"3F",X"01",X"01",X"03",
		X"F8",X"FE",X"7F",X"DF",X"FF",X"FF",X"3F",X"7F",X"00",X"00",X"00",X"80",X"80",X"80",X"00",X"00",
		X"FF",X"FF",X"7F",X"FF",X"DF",X"FF",X"FE",X"F8",X"80",X"4A",X"BC",X"88",X"80",X"00",X"00",X"00",
		X"0F",X"1D",X"0C",X"08",X"4C",X"5D",X"7F",X"7E",X"F0",X"F8",X"D8",X"BC",X"DE",X"DE",X"FE",X"7E",
		X"3E",X"06",X"06",X"00",X"00",X"00",X"00",X"00",X"7C",X"60",X"60",X"00",X"00",X"00",X"00",X"00",
		X"1D",X"0C",X"08",X"1C",X"5D",X"5D",X"7E",X"78",X"F8",X"D8",X"BC",X"DC",X"DE",X"DE",X"3E",X"1E",
		X"78",X"F0",X"F0",X"E0",X"E0",X"E0",X"00",X"00",X"1E",X"0F",X"0F",X"07",X"07",X"07",X"00",X"00",
		X"C8",X"9C",X"1D",X"3F",X"1F",X"1F",X"0F",X"0F",X"BF",X"D9",X"D8",X"F8",X"F8",X"F8",X"F0",X"F0",
		X"07",X"07",X"07",X"03",X"03",X"00",X"00",X"00",X"E0",X"E0",X"E0",X"C0",X"C0",X"00",X"00",X"00",
		X"1D",X"0C",X"08",X"0C",X"5D",X"5D",X"7A",X"78",X"F8",X"D8",X"BC",X"DC",X"DE",X"DE",X"3E",X"1E",
		X"7C",X"3C",X"1C",X"1C",X"00",X"00",X"00",X"00",X"3E",X"3C",X"38",X"38",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"01",X"01",X"07",X"07",X"00",X"00",X"F0",X"C0",X"E2",X"FF",X"F7",X"C1",X"63",
		X"00",X"07",X"07",X"01",X"01",X"01",X"00",X"00",X"7F",X"F7",X"CB",X"FF",X"FE",X"F8",X"F0",X"00",
		X"00",X"00",X"0F",X"3F",X"FC",X"FC",X"F8",X"F8",X"00",X"00",X"80",X"F0",X"B8",X"1C",X"0C",X"00",
		X"FC",X"FE",X"FF",X"FC",X"3F",X"0F",X"00",X"00",X"00",X"9C",X"FC",X"B8",X"F0",X"80",X"00",X"00",
		X"00",X"01",X"03",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"F0",X"C0",X"F1",X"FF",X"3B",X"40",X"31",
		X"00",X"00",X"0F",X"0F",X"0F",X"03",X"01",X"00",X"3F",X"3B",X"45",X"FF",X"FF",X"FC",X"F0",X"00",
		X"1C",X"1E",X"1E",X"0E",X"FE",X"FE",X"FC",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FE",X"FE",X"0E",X"1E",X"1E",X"1C",X"00",X"E8",X"F0",X"20",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"7E",X"18",X"18",X"18",X"18",X"18",X"18",X"00",X"7F",X"60",X"60",X"7E",X"60",X"60",X"7F",
		X"00",X"63",X"63",X"63",X"7F",X"63",X"63",X"63",X"00",X"63",X"66",X"6C",X"7C",X"6E",X"67",X"63",
		X"00",X"1C",X"36",X"63",X"63",X"7F",X"63",X"63",X"00",X"63",X"63",X"73",X"6B",X"67",X"63",X"63",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"78",X"30",X"30",X"30",X"30",X"31",X"7F",
		X"00",X"00",X"00",X"00",X"01",X"06",X"04",X"08",X"00",X"00",X"00",X"00",X"C0",X"30",X"10",X"88",
		X"09",X"08",X"04",X"06",X"01",X"00",X"00",X"00",X"C8",X"88",X"10",X"30",X"C0",X"00",X"00",X"00",
		X"00",X"7E",X"18",X"18",X"18",X"18",X"18",X"18",X"00",X"7C",X"62",X"63",X"63",X"63",X"63",X"7E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"03",X"03",X"03",X"07",X"0F",X"1F",X"E0",X"F0",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"1F",X"1F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"07",X"07",X"07",X"1F",X"1F",X"3F",X"3F",X"7F",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"01",X"01",X"03",X"03",X"03",X"07",X"07",X"C0",X"E0",X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"44",X"C6",X"C6",X"82",X"C6",X"7C",X"7C",X"7C",X"7C",X"FE",X"FE",X"EE",X"6C",X"6C",X"00",
		X"00",X"10",X"1C",X"1E",X"00",X"00",X"00",X"14",X"00",X"00",X"00",X"00",X"30",X"7C",X"78",X"38",
		X"3E",X"14",X"00",X"00",X"00",X"1E",X"1C",X"10",X"00",X"38",X"78",X"7C",X"30",X"00",X"00",X"00",
		X"06",X"0E",X"0E",X"04",X"01",X"01",X"04",X"3E",X"00",X"00",X"18",X"FC",X"FE",X"FF",X"CF",X"07",
		X"04",X"01",X"01",X"04",X"0E",X"0E",X"06",X"00",X"CF",X"FF",X"FE",X"FC",X"18",X"00",X"00",X"00",
		X"00",X"00",X"08",X"0E",X"1E",X"1E",X"0C",X"00",X"00",X"00",X"20",X"E0",X"F0",X"F0",X"60",X"00",
		X"00",X"21",X"63",X"61",X"E3",X"01",X"00",X"00",X"00",X"08",X"8C",X"0C",X"8E",X"00",X"00",X"00",
		X"07",X"0F",X"1F",X"3E",X"3C",X"1C",X"1E",X"1E",X"C0",X"E0",X"F0",X"F8",X"78",X"70",X"F0",X"F0",
		X"0C",X"E1",X"F3",X"61",X"01",X"01",X"00",X"00",X"60",X"0E",X"9E",X"0C",X"00",X"00",X"00",X"00",
		X"01",X"07",X"0D",X"09",X"19",X"1F",X"01",X"1D",X"80",X"E0",X"B0",X"90",X"98",X"F8",X"80",X"B8",
		X"01",X"1D",X"01",X"0D",X"01",X"01",X"07",X"1F",X"80",X"B8",X"80",X"B0",X"80",X"80",X"E0",X"F8",
		X"00",X"00",X"00",X"82",X"8A",X"CA",X"C0",X"FF",X"00",X"00",X"00",X"B0",X"BC",X"A6",X"22",X"FF",
		X"FF",X"C0",X"CA",X"8A",X"82",X"00",X"00",X"00",X"FF",X"22",X"A6",X"BC",X"B0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"0E",X"0E",X"0C",X"00",X"00",X"00",X"00",X"10",X"38",X"38",X"18",
		X"00",X"10",X"31",X"30",X"20",X"00",X"00",X"00",X"00",X"84",X"C6",X"86",X"82",X"80",X"00",X"00",
		X"00",X"00",X"1C",X"0E",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"E0",X"F0",X"60",X"00",
		X"3E",X"04",X"00",X"00",X"00",X"0E",X"1C",X"00",X"00",X"00",X"60",X"F0",X"E0",X"00",X"00",X"00",
		X"70",X"F9",X"C3",X"FB",X"73",X"07",X"0F",X"19",X"1C",X"3E",X"06",X"3E",X"1C",X"00",X"60",X"30",
		X"19",X"0C",X"60",X"EC",X"CC",X"DC",X"FC",X"78",X"30",X"60",X"0C",X"6E",X"66",X"76",X"7E",X"3C",
		X"70",X"F8",X"C1",X"F9",X"73",X"03",X"07",X"03",X"0E",X"9F",X"83",X"9F",X"8E",X"00",X"60",X"30",
		X"03",X"06",X"60",X"EC",X"CC",X"DC",X"FC",X"78",X"30",X"60",X"06",X"37",X"33",X"3B",X"3F",X"1E",
		X"00",X"F8",X"F8",X"F0",X"F1",X"00",X"00",X"00",X"00",X"3C",X"7E",X"FF",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"E3",X"F3",X"F3",X"FB",X"FB",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"C3",X"C3",X"00",
		X"00",X"00",X"00",X"02",X"07",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"06",X"1C",X"3E",X"3E",X"3E",X"1C",X"00",X"00",X"00",X"70",X"F8",X"F8",X"F8",X"70",X"00",
		X"00",X"1F",X"1F",X"1F",X"9F",X"00",X"00",X"00",X"00",X"3E",X"3E",X"BE",X"BE",X"00",X"00",X"00",
		X"00",X"00",X"DF",X"DF",X"DF",X"DF",X"DF",X"00",X"00",X"00",X"FE",X"7E",X"7E",X"3E",X"3E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"00",X"00",X"00",X"00",X"3F",X"FF",X"FF",X"FF",
		X"07",X"07",X"0F",X"0F",X"0F",X"0F",X"07",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"FE",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",X"F0",X"F0",
		X"01",X"07",X"0F",X"0F",X"0F",X"07",X"03",X"01",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"7F",X"3F",X"7F",X"7F",X"FF",X"FF",X"FF",X"C0",X"F0",X"F8",X"F8",X"F8",X"F0",X"E0",X"C0",
		X"0E",X"1E",X"1C",X"1F",X"1F",X"1F",X"1F",X"06",X"00",X"00",X"00",X"00",X"B0",X"78",X"78",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"1E",X"1C",X"1F",X"1F",X"1E",X"1E",X"0C",X"00",X"00",X"00",X"00",X"60",X"F0",X"F0",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"78",X"F0",X"E0",X"FB",X"FF",X"F7",X"F3",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"1F",X"1F",X"0F",X"06",X"0A",X"15",X"0A",X"30",X"78",X"F8",X"78",X"30",X"A8",X"54",X"A8",
		X"00",X"01",X"03",X"0B",X"23",X"03",X"02",X"83",X"7F",X"FB",X"FF",X"DF",X"FE",X"FF",X"FB",X"BF",
		X"2B",X"52",X"03",X"A3",X"07",X"07",X"2E",X"0C",X"FF",X"F8",X"C2",X"80",X"0A",X"50",X"82",X"00",
		X"FF",X"FF",X"7F",X"FF",X"FD",X"FF",X"FF",X"AF",X"00",X"C8",X"E4",X"E0",X"61",X"E8",X"E0",X"E9",
		X"FD",X"47",X"01",X"20",X"88",X"00",X"25",X"00",X"64",X"E0",X"E0",X"E1",X"74",X"70",X"38",X"18",
		X"03",X"1C",X"24",X"48",X"58",X"59",X"3A",X"44",X"80",X"5C",X"E6",X"EE",X"FE",X"F6",X"63",X"EF",
		X"9C",X"9D",X"8E",X"4C",X"3C",X"7C",X"3A",X"01",X"FE",X"FC",X"FC",X"FE",X"FE",X"6E",X"44",X"B8",
		X"00",X"00",X"00",X"00",X"03",X"0F",X"1F",X"3E",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",
		X"3F",X"0F",X"7F",X"7F",X"3B",X"00",X"00",X"00",X"C0",X"FE",X"FE",X"FE",X"DC",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"0F",X"1F",X"3C",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",
		X"3E",X"0F",X"7F",X"7E",X"38",X"00",X"00",X"00",X"60",X"FE",X"FE",X"7E",X"1C",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"0F",X"1F",X"3C",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",
		X"3E",X"0F",X"0F",X"0E",X"08",X"00",X"00",X"00",X"60",X"FE",X"F0",X"70",X"10",X"00",X"00",X"00",
		X"00",X"00",X"00",X"02",X"02",X"02",X"02",X"00",X"40",X"50",X"58",X"DC",X"DC",X"DC",X"4C",X"4C",
		X"05",X"04",X"01",X"01",X"01",X"01",X"01",X"05",X"4C",X"4C",X"5C",X"5C",X"5C",X"1C",X"5C",X"4C",
		X"20",X"63",X"70",X"F0",X"F0",X"F0",X"F8",X"78",X"00",X"F6",X"00",X"00",X"1F",X"00",X"00",X"20",
		X"3D",X"1F",X"0F",X"00",X"00",X"00",X"00",X"00",X"F8",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"00",X"00",X"ED",X"00",X"00",X"00",X"00",X"C0",X"00",X"38",X"00",X"00",X"00",X"00",
		X"18",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"E6",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"CF",X"86",X"06",X"02",X"00",X"00",X"00",X"00",X"F8",X"D8",X"08",X"08",X"0C",X"0C",X"0C",X"1C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"18",X"18",X"18",X"38",X"38",X"18",X"30",
		X"00",X"00",X"00",X"05",X"0D",X"0F",X"0F",X"1F",X"7F",X"FE",X"FC",X"F8",X"F8",X"FC",X"FE",X"FF",
		X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",X"F8",X"E0",X"C0",X"E0",X"F0",X"F0",X"F0",X"F0",
		X"50",X"3A",X"C8",X"4D",X"10",X"26",X"08",X"A2",X"00",X"00",X"00",X"00",X"5D",X"28",X"E2",X"10",
		X"00",X"00",X"00",X"00",X"01",X"16",X"22",X"74",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"08",X"2A",X"E3",X"5A",X"04",X"20",X"52",X"00",X"00",X"00",X"00",X"01",X"05",X"0A",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"06",X"0A",X"00",X"03",X"10",X"04",X"0A",X"02",X"10",X"00",
		X"1F",X"10",X"10",X"1E",X"01",X"01",X"1E",X"00",X"00",X"38",X"44",X"44",X"44",X"44",X"38",X"00",
		X"00",X"FE",X"28",X"FE",X"AA",X"AA",X"AA",X"FE",X"00",X"DF",X"11",X"D1",X"1F",X"12",X"51",X"D1",
		X"00",X"04",X"04",X"05",X"05",X"01",X"09",X"09",X"5C",X"5C",X"5C",X"4C",X"4C",X"DC",X"DC",X"CC",
		X"08",X"00",X"00",X"01",X"07",X"0F",X"1F",X"1F",X"4C",X"5C",X"4C",X"CC",X"FC",X"FC",X"FC",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"00",X"1C",X"06",X"02",X"02",X"02",X"00",X"00",
		X"78",X"79",X"73",X"23",X"03",X"01",X"00",X"00",X"E0",X"E0",X"E0",X"F0",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"03",X"0F",X"1F",X"3F",X"3F",X"00",X"00",X"00",X"C0",X"F0",X"F8",X"F8",X"F8",
		X"7F",X"7F",X"7F",X"7F",X"3F",X"2A",X"10",X"00",X"F8",X"F0",X"C0",X"40",X"00",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"18",X"78",X"20",X"30",X"78",X"58",X"D8",X"BC",
		X"3E",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"3C",X"F8",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"06",X"0F",X"1F",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",
		X"1F",X"1F",X"1F",X"0F",X"0F",X"0E",X"04",X"00",X"C0",X"E0",X"80",X"20",X"00",X"00",X"00",X"00",
		X"28",X"8A",X"84",X"80",X"96",X"96",X"96",X"96",X"04",X"11",X"D2",X"D0",X"D1",X"D9",X"D8",X"D2",
		X"B6",X"96",X"96",X"96",X"16",X"16",X"06",X"06",X"F6",X"EC",X"ED",X"ED",X"DB",X"DB",X"DB",X"DB",
		X"17",X"17",X"17",X"07",X"03",X"00",X"00",X"00",X"68",X"20",X"02",X"F2",X"F2",X"FA",X"FA",X"FA",
		X"FA",X"FA",X"FA",X"FA",X"FA",X"F8",X"00",X"00",X"00",X"46",X"53",X"52",X"50",X"56",X"57",X"37",
		X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"49",X"54",X"88",X"40",X"92",X"00",X"78",X"78",
		X"7A",X"FA",X"7A",X"7A",X"78",X"78",X"7A",X"7A",X"18",X"8A",X"A6",X"A1",X"88",X"8B",X"8B",X"AB",
		X"AB",X"AB",X"AB",X"8B",X"8B",X"AB",X"AB",X"AB",X"44",X"D6",X"4D",X"24",X"48",X"00",X"BF",X"BF",
		X"BF",X"BF",X"FF",X"BF",X"BF",X"BF",X"BF",X"BF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"08",X"1B",X"17",X"07",X"0A",X"18",X"00",X"00",X"00",X"00",X"18",X"38",X"30",X"50",
		X"12",X"06",X"06",X"08",X"1D",X"1D",X"08",X"00",X"E0",X"40",X"40",X"80",X"80",X"00",X"00",X"00",
		X"00",X"20",X"67",X"28",X"28",X"28",X"28",X"27",X"00",X"00",X"70",X"88",X"88",X"88",X"88",X"70",
		X"00",X"2F",X"68",X"28",X"2F",X"20",X"28",X"27",X"00",X"80",X"38",X"44",X"44",X"C4",X"C4",X"38",
		X"00",X"38",X"44",X"05",X"19",X"21",X"41",X"7C",X"00",X"00",X"EE",X"11",X"11",X"11",X"11",X"EE",
		X"00",X"38",X"44",X"05",X"19",X"05",X"45",X"38",X"00",X"00",X"EE",X"11",X"11",X"11",X"11",X"EE",
		X"00",X"08",X"18",X"29",X"49",X"49",X"7D",X"08",X"00",X"00",X"EE",X"11",X"11",X"11",X"11",X"EE",
		X"00",X"38",X"44",X"41",X"79",X"45",X"45",X"38",X"00",X"00",X"EE",X"11",X"11",X"11",X"11",X"EE",
		X"00",X"00",X"00",X"00",X"0E",X"1C",X"1F",X"1F",X"00",X"00",X"00",X"F0",X"38",X"44",X"E0",X"C0",
		X"1F",X"1F",X"0F",X"0E",X"07",X"03",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"0E",X"1F",X"1F",X"00",X"00",X"00",X"00",X"80",X"70",X"F0",X"E0",
		X"3F",X"3F",X"3F",X"1F",X"1E",X"08",X"00",X"00",X"E0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"0E",X"1E",X"1F",X"3F",X"3F",X"00",X"00",X"C0",X"70",X"78",X"F0",X"F0",X"F0",
		X"3F",X"3F",X"1F",X"07",X"00",X"00",X"00",X"00",X"E0",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"07",X"0F",X"1F",X"1F",X"00",X"00",X"80",X"E0",X"F0",X"F8",X"FC",X"FC",
		X"3F",X"3F",X"1F",X"0E",X"00",X"00",X"00",X"00",X"FC",X"FC",X"FC",X"F8",X"00",X"00",X"00",X"00",
		X"00",X"38",X"44",X"45",X"39",X"45",X"45",X"38",X"00",X"00",X"EE",X"11",X"11",X"11",X"11",X"EE",
		X"00",X"38",X"44",X"45",X"3D",X"05",X"45",X"38",X"00",X"00",X"EE",X"11",X"11",X"11",X"11",X"EE",
		X"00",X"4E",X"D1",X"41",X"46",X"48",X"50",X"5F",X"00",X"00",X"36",X"49",X"49",X"49",X"49",X"36",
		X"00",X"4E",X"D1",X"50",X"5E",X"51",X"51",X"4E",X"00",X"00",X"36",X"49",X"49",X"49",X"49",X"36",
		X"00",X"00",X"78",X"9D",X"9D",X"1D",X"1D",X"39",X"00",X"00",X"EE",X"33",X"33",X"33",X"33",X"33",
		X"71",X"E1",X"E1",X"E1",X"FC",X"00",X"00",X"00",X"33",X"33",X"33",X"FF",X"EE",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0E",X"7F",X"3F",X"3F",X"3F",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"E0",
		X"1F",X"1F",X"07",X"01",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F8",X"38",X"08",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
