library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity BASIC11 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of BASIC11 is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"4C",X"CC",X"EC",X"4C",X"71",X"C4",X"72",X"C9",X"91",X"C6",X"86",X"E9",X"D0",X"E9",X"15",X"CD",
		X"18",X"CD",X"11",X"CA",X"50",X"DA",X"A0",X"DA",X"DD",X"D9",X"66",X"D9",X"84",X"DA",X"A0",X"DA",
		X"54",X"C8",X"FC",X"C7",X"08",X"C8",X"97",X"CE",X"3B",X"CA",X"54",X"CD",X"7D",X"D1",X"CD",X"CC",
		X"88",X"CD",X"1B",X"CB",X"E4",X"C9",X"BC",X"C9",X"6F",X"CA",X"51",X"C9",X"C7",X"C9",X"11",X"CA",
		X"98",X"CA",X"CD",X"EB",X"E6",X"EB",X"0B",X"EC",X"20",X"EC",X"32",X"EC",X"B4",X"FA",X"CA",X"FA",
		X"E0",X"FA",X"9E",X"FA",X"FB",X"EA",X"FB",X"EA",X"FB",X"EA",X"EF",X"EA",X"EF",X"EA",X"EF",X"EA",
		X"EF",X"EA",X"EF",X"EA",X"EF",X"EA",X"EF",X"EA",X"FB",X"EA",X"FB",X"EA",X"70",X"C9",X"C1",X"CA",
		X"57",X"D9",X"5A",X"E8",X"08",X"E9",X"B9",X"D4",X"4E",X"D9",X"AA",X"CB",X"9F",X"C9",X"47",X"C7",
		X"0C",X"C7",X"45",X"CD",X"45",X"E9",X"12",X"CD",X"ED",X"C6",X"21",X"DF",X"BD",X"DF",X"49",X"DF",
		X"21",X"00",X"7E",X"D4",X"A6",X"D4",X"B5",X"D9",X"FB",X"02",X"2E",X"E2",X"4F",X"E3",X"AF",X"DC",
		X"AA",X"E2",X"8B",X"E3",X"92",X"E3",X"DB",X"E3",X"3F",X"E4",X"38",X"D9",X"83",X"D9",X"D4",X"DD",
		X"A6",X"D8",X"93",X"D5",X"D7",X"D8",X"B5",X"D8",X"16",X"D8",X"77",X"DE",X"0F",X"DF",X"0B",X"DF",
		X"DA",X"DA",X"3F",X"DA",X"45",X"EC",X"2A",X"D8",X"56",X"D8",X"61",X"D8",X"79",X"24",X"DB",X"79",
		X"0D",X"DB",X"7B",X"EF",X"DC",X"7B",X"E6",X"DD",X"7F",X"37",X"E2",X"50",X"E5",X"D0",X"46",X"E2",
		X"D0",X"7D",X"70",X"E2",X"5A",X"3B",X"D0",X"64",X"12",X"D1",X"45",X"4E",X"C4",X"45",X"44",X"49",
		X"D4",X"53",X"54",X"4F",X"52",X"C5",X"52",X"45",X"43",X"41",X"4C",X"CC",X"54",X"52",X"4F",X"CE",
		X"54",X"52",X"4F",X"46",X"C6",X"50",X"4F",X"D0",X"50",X"4C",X"4F",X"D4",X"50",X"55",X"4C",X"CC",
		X"4C",X"4F",X"52",X"45",X"D3",X"44",X"4F",X"4B",X"C5",X"52",X"45",X"50",X"45",X"41",X"D4",X"55",
		X"4E",X"54",X"49",X"CC",X"46",X"4F",X"D2",X"4C",X"4C",X"49",X"53",X"D4",X"4C",X"50",X"52",X"49",
		X"4E",X"D4",X"4E",X"45",X"58",X"D4",X"44",X"41",X"54",X"C1",X"49",X"4E",X"50",X"55",X"D4",X"44",
		X"49",X"CD",X"43",X"4C",X"D3",X"52",X"45",X"41",X"C4",X"4C",X"45",X"D4",X"47",X"4F",X"54",X"CF",
		X"52",X"55",X"CE",X"49",X"C6",X"52",X"45",X"53",X"54",X"4F",X"52",X"C5",X"47",X"4F",X"53",X"55",
		X"C2",X"52",X"45",X"54",X"55",X"52",X"CE",X"52",X"45",X"CD",X"48",X"49",X"4D",X"45",X"CD",X"47",
		X"52",X"41",X"C2",X"52",X"45",X"4C",X"45",X"41",X"53",X"C5",X"54",X"45",X"58",X"D4",X"48",X"49",
		X"52",X"45",X"D3",X"53",X"48",X"4F",X"4F",X"D4",X"45",X"58",X"50",X"4C",X"4F",X"44",X"C5",X"5A",
		X"41",X"D0",X"50",X"49",X"4E",X"C7",X"53",X"4F",X"55",X"4E",X"C4",X"4D",X"55",X"53",X"49",X"C3",
		X"50",X"4C",X"41",X"D9",X"43",X"55",X"52",X"53",X"45",X"D4",X"43",X"55",X"52",X"4D",X"4F",X"D6",
		X"44",X"52",X"41",X"D7",X"43",X"49",X"52",X"43",X"4C",X"C5",X"50",X"41",X"54",X"54",X"45",X"52",
		X"CE",X"46",X"49",X"4C",X"CC",X"43",X"48",X"41",X"D2",X"50",X"41",X"50",X"45",X"D2",X"49",X"4E",
		X"CB",X"53",X"54",X"4F",X"D0",X"4F",X"CE",X"57",X"41",X"49",X"D4",X"43",X"4C",X"4F",X"41",X"C4",
		X"43",X"53",X"41",X"56",X"C5",X"44",X"45",X"C6",X"50",X"4F",X"4B",X"C5",X"50",X"52",X"49",X"4E",
		X"D4",X"43",X"4F",X"4E",X"D4",X"4C",X"49",X"53",X"D4",X"43",X"4C",X"45",X"41",X"D2",X"47",X"45",
		X"D4",X"43",X"41",X"4C",X"CC",X"A1",X"4E",X"45",X"D7",X"54",X"41",X"42",X"A8",X"54",X"CF",X"46",
		X"CE",X"53",X"50",X"43",X"A8",X"C0",X"41",X"55",X"54",X"CF",X"45",X"4C",X"53",X"C5",X"54",X"48",
		X"45",X"CE",X"4E",X"4F",X"D4",X"53",X"54",X"45",X"D0",X"AB",X"AD",X"AA",X"AF",X"DE",X"41",X"4E",
		X"C4",X"4F",X"D2",X"BE",X"BD",X"BC",X"53",X"47",X"CE",X"49",X"4E",X"D4",X"41",X"42",X"D3",X"55",
		X"53",X"D2",X"46",X"52",X"C5",X"50",X"4F",X"D3",X"48",X"45",X"58",X"A4",X"A6",X"53",X"51",X"D2",
		X"52",X"4E",X"C4",X"4C",X"CE",X"45",X"58",X"D0",X"43",X"4F",X"D3",X"53",X"49",X"CE",X"54",X"41",
		X"CE",X"41",X"54",X"CE",X"50",X"45",X"45",X"CB",X"44",X"45",X"45",X"CB",X"4C",X"4F",X"C7",X"4C",
		X"45",X"CE",X"53",X"54",X"52",X"A4",X"56",X"41",X"CC",X"41",X"53",X"C3",X"43",X"48",X"52",X"A4",
		X"50",X"C9",X"54",X"52",X"55",X"C5",X"46",X"41",X"4C",X"53",X"C5",X"4B",X"45",X"59",X"A4",X"53",
		X"43",X"52",X"CE",X"50",X"4F",X"49",X"4E",X"D4",X"4C",X"45",X"46",X"54",X"A4",X"52",X"49",X"47",
		X"48",X"54",X"A4",X"4D",X"49",X"44",X"A4",X"00",X"4E",X"45",X"58",X"54",X"20",X"57",X"49",X"54",
		X"48",X"4F",X"55",X"54",X"20",X"46",X"4F",X"D2",X"53",X"59",X"4E",X"54",X"41",X"D8",X"52",X"45",
		X"54",X"55",X"52",X"4E",X"20",X"57",X"49",X"54",X"48",X"4F",X"55",X"54",X"20",X"47",X"4F",X"53",
		X"55",X"C2",X"4F",X"55",X"54",X"20",X"4F",X"46",X"20",X"44",X"41",X"54",X"C1",X"49",X"4C",X"4C",
		X"45",X"47",X"41",X"4C",X"20",X"51",X"55",X"41",X"4E",X"54",X"49",X"54",X"D9",X"4F",X"56",X"45",
		X"52",X"46",X"4C",X"4F",X"D7",X"4F",X"55",X"54",X"20",X"4F",X"46",X"20",X"4D",X"45",X"4D",X"4F",
		X"52",X"D9",X"55",X"4E",X"44",X"45",X"46",X"27",X"44",X"20",X"53",X"54",X"41",X"54",X"45",X"4D",
		X"45",X"4E",X"D4",X"42",X"41",X"44",X"20",X"53",X"55",X"42",X"53",X"43",X"52",X"49",X"50",X"D4",
		X"52",X"45",X"44",X"49",X"4D",X"27",X"44",X"20",X"41",X"52",X"52",X"41",X"D9",X"44",X"49",X"56",
		X"49",X"53",X"49",X"4F",X"4E",X"20",X"42",X"59",X"20",X"5A",X"45",X"52",X"CF",X"49",X"4C",X"4C",
		X"45",X"47",X"41",X"4C",X"20",X"44",X"49",X"52",X"45",X"43",X"D4",X"44",X"49",X"53",X"50",X"20",
		X"54",X"59",X"50",X"45",X"20",X"4D",X"49",X"53",X"4D",X"41",X"54",X"43",X"C8",X"53",X"54",X"52",
		X"49",X"4E",X"47",X"20",X"54",X"4F",X"4F",X"20",X"4C",X"4F",X"4E",X"C7",X"46",X"4F",X"52",X"4D",
		X"55",X"4C",X"41",X"20",X"54",X"4F",X"4F",X"20",X"43",X"4F",X"4D",X"50",X"4C",X"45",X"D8",X"43",
		X"41",X"4E",X"27",X"54",X"20",X"43",X"4F",X"4E",X"54",X"49",X"4E",X"55",X"C5",X"55",X"4E",X"44",
		X"45",X"46",X"27",X"44",X"20",X"46",X"55",X"4E",X"43",X"54",X"49",X"4F",X"CE",X"42",X"41",X"44",
		X"20",X"55",X"4E",X"54",X"49",X"CC",X"20",X"45",X"52",X"52",X"4F",X"52",X"00",X"20",X"49",X"4E",
		X"20",X"00",X"0D",X"0A",X"52",X"65",X"61",X"64",X"79",X"20",X"0D",X"0A",X"00",X"0D",X"0A",X"20",
		X"42",X"52",X"45",X"41",X"4B",X"00",X"BA",X"E8",X"E8",X"E8",X"E8",X"BD",X"01",X"01",X"C9",X"8D",
		X"D0",X"21",X"A5",X"B9",X"D0",X"0A",X"BD",X"02",X"01",X"85",X"B8",X"BD",X"03",X"01",X"85",X"B9",
		X"DD",X"03",X"01",X"D0",X"07",X"A5",X"B8",X"DD",X"02",X"01",X"F0",X"07",X"8A",X"18",X"69",X"12",
		X"AA",X"D0",X"D8",X"60",X"20",X"44",X"C4",X"85",X"A0",X"84",X"A1",X"38",X"A5",X"C9",X"E5",X"CE",
		X"85",X"91",X"A8",X"A5",X"CA",X"E5",X"CF",X"AA",X"E8",X"98",X"F0",X"23",X"A5",X"C9",X"38",X"E5",
		X"91",X"85",X"C9",X"B0",X"03",X"C6",X"CA",X"38",X"A5",X"C7",X"E5",X"91",X"85",X"C7",X"B0",X"08",
		X"C6",X"C8",X"90",X"04",X"B1",X"C9",X"91",X"C7",X"88",X"D0",X"F9",X"B1",X"C9",X"91",X"C7",X"C6",
		X"CA",X"C6",X"C8",X"CA",X"D0",X"F2",X"60",X"0A",X"69",X"3E",X"B0",X"40",X"85",X"91",X"BA",X"E4",
		X"91",X"90",X"39",X"60",X"C4",X"A3",X"90",X"28",X"D0",X"04",X"C5",X"A2",X"90",X"22",X"48",X"A2",
		X"09",X"98",X"48",X"B5",X"C6",X"CA",X"10",X"FA",X"20",X"50",X"D6",X"A2",X"F7",X"68",X"95",X"D0",
		X"E8",X"30",X"FA",X"68",X"A8",X"68",X"C4",X"A3",X"90",X"06",X"D0",X"10",X"C5",X"A2",X"B0",X"0C",
		X"60",X"AD",X"C0",X"02",X"29",X"FE",X"8D",X"C0",X"02",X"4C",X"A8",X"C4",X"A2",X"4D",X"20",X"2F",
		X"C8",X"46",X"2E",X"20",X"F0",X"CB",X"20",X"D7",X"CC",X"BD",X"A8",X"C2",X"48",X"29",X"7F",X"20",
		X"D9",X"CC",X"E8",X"68",X"10",X"F3",X"20",X"26",X"C7",X"A9",X"A6",X"A0",X"C3",X"20",X"B0",X"CC",
		X"A4",X"A9",X"C8",X"F0",X"03",X"20",X"BA",X"E0",X"4E",X"52",X"02",X"46",X"2E",X"4E",X"F2",X"02",
		X"A9",X"B2",X"A0",X"C3",X"20",X"1A",X"00",X"20",X"2F",X"C8",X"20",X"92",X"C5",X"86",X"E9",X"84",
		X"EA",X"20",X"E2",X"00",X"AA",X"F0",X"F0",X"A2",X"FF",X"86",X"A9",X"90",X"06",X"20",X"FA",X"C5",
		X"4C",X"0C",X"C9",X"20",X"E2",X"CA",X"20",X"FA",X"C5",X"84",X"26",X"20",X"B3",X"C6",X"90",X"44",
		X"A0",X"01",X"B1",X"CE",X"85",X"92",X"A5",X"9C",X"85",X"91",X"A5",X"CF",X"85",X"94",X"A5",X"CE",
		X"88",X"F1",X"CE",X"18",X"65",X"9C",X"85",X"9C",X"85",X"93",X"A5",X"9D",X"69",X"FF",X"85",X"9D",
		X"E5",X"CF",X"AA",X"38",X"A5",X"CE",X"E5",X"9C",X"A8",X"B0",X"03",X"E8",X"C6",X"94",X"18",X"65",
		X"91",X"90",X"03",X"C6",X"92",X"18",X"B1",X"91",X"91",X"93",X"C8",X"D0",X"F9",X"E6",X"92",X"E6",
		X"94",X"CA",X"D0",X"F2",X"20",X"08",X"C7",X"20",X"5F",X"C5",X"A5",X"35",X"F0",X"89",X"18",X"A5",
		X"9C",X"85",X"C9",X"65",X"26",X"85",X"C7",X"A4",X"9D",X"84",X"CA",X"90",X"01",X"C8",X"84",X"C8",
		X"20",X"F4",X"C3",X"A5",X"A0",X"A4",X"A1",X"85",X"9C",X"84",X"9D",X"A4",X"26",X"88",X"B9",X"31",
		X"00",X"91",X"CE",X"88",X"10",X"F8",X"20",X"08",X"C7",X"20",X"5F",X"C5",X"4C",X"B7",X"C4",X"A5",
		X"9A",X"A4",X"9B",X"85",X"91",X"84",X"92",X"18",X"A0",X"01",X"B1",X"91",X"F0",X"1D",X"A0",X"04",
		X"C8",X"B1",X"91",X"D0",X"FB",X"C8",X"98",X"65",X"91",X"AA",X"A0",X"00",X"91",X"91",X"A5",X"92",
		X"69",X"00",X"C8",X"91",X"91",X"86",X"91",X"85",X"92",X"90",X"DD",X"60",X"CA",X"10",X"05",X"20",
		X"F0",X"CB",X"A2",X"00",X"20",X"E8",X"C5",X"C9",X"01",X"D0",X"0D",X"AC",X"69",X"02",X"B1",X"12",
		X"29",X"7F",X"C9",X"20",X"B0",X"02",X"A9",X"09",X"48",X"20",X"D9",X"CC",X"68",X"C9",X"7F",X"F0",
		X"DB",X"C9",X"0D",X"F0",X"30",X"C9",X"03",X"F0",X"28",X"C9",X"18",X"F0",X"0B",X"C9",X"20",X"90",
		X"D3",X"95",X"35",X"E8",X"E0",X"4F",X"90",X"07",X"A9",X"5C",X"20",X"D9",X"CC",X"D0",X"C0",X"E0",
		X"4C",X"90",X"C1",X"8A",X"48",X"98",X"48",X"20",X"9F",X"FA",X"68",X"A8",X"68",X"AA",X"4C",X"94",
		X"C5",X"E6",X"17",X"A2",X"00",X"4C",X"EA",X"CB",X"20",X"3B",X"02",X"10",X"FB",X"C9",X"0F",X"D0",
		X"08",X"48",X"A5",X"2E",X"49",X"FF",X"85",X"2E",X"68",X"60",X"A6",X"E9",X"A0",X"04",X"84",X"2A",
		X"B5",X"00",X"C9",X"20",X"F0",X"41",X"85",X"25",X"C9",X"22",X"F0",X"5F",X"24",X"2A",X"70",X"37",
		X"C9",X"3F",X"D0",X"04",X"A9",X"BA",X"D0",X"2F",X"C9",X"30",X"90",X"04",X"C9",X"3C",X"90",X"27",
		X"84",X"E0",X"A0",X"00",X"84",X"26",X"A9",X"E9",X"85",X"18",X"A9",X"C0",X"85",X"19",X"86",X"E9",
		X"CA",X"E8",X"E6",X"18",X"D0",X"02",X"E6",X"19",X"B5",X"00",X"38",X"F1",X"18",X"F0",X"F2",X"C9",
		X"80",X"D0",X"2F",X"05",X"26",X"A4",X"E0",X"E8",X"C8",X"99",X"30",X"00",X"B9",X"30",X"00",X"F0",
		X"39",X"38",X"E9",X"3A",X"F0",X"04",X"C9",X"57",X"D0",X"02",X"85",X"2A",X"38",X"E9",X"63",X"D0",
		X"9F",X"85",X"25",X"B5",X"00",X"F0",X"E0",X"C5",X"25",X"F0",X"DC",X"C8",X"99",X"30",X"00",X"E8",
		X"D0",X"F1",X"A6",X"E9",X"E6",X"26",X"B1",X"18",X"08",X"E6",X"18",X"D0",X"02",X"E6",X"19",X"28",
		X"10",X"F4",X"B1",X"18",X"D0",X"B2",X"B5",X"00",X"10",X"BB",X"99",X"32",X"00",X"A9",X"34",X"85",
		X"E9",X"60",X"20",X"E2",X"CA",X"20",X"B3",X"C6",X"90",X"16",X"6E",X"F2",X"02",X"20",X"6C",X"C7",
		X"4E",X"F2",X"02",X"20",X"F0",X"CB",X"A9",X"0B",X"20",X"D9",X"CC",X"68",X"68",X"4C",X"B7",X"C4",
		X"4C",X"23",X"CA",X"A9",X"00",X"85",X"1D",X"85",X"1E",X"A5",X"9A",X"A6",X"9B",X"A0",X"01",X"85",
		X"CE",X"86",X"CF",X"B1",X"CE",X"F0",X"25",X"C8",X"C8",X"E6",X"1D",X"D0",X"02",X"E6",X"1E",X"A5",
		X"34",X"D1",X"CE",X"90",X"18",X"F0",X"03",X"88",X"D0",X"09",X"A5",X"33",X"88",X"D1",X"CE",X"90",
		X"0C",X"F0",X"0A",X"88",X"B1",X"CE",X"AA",X"88",X"B1",X"CE",X"B0",X"D1",X"18",X"60",X"D0",X"FD",
		X"A9",X"00",X"4E",X"F4",X"02",X"A8",X"91",X"9A",X"C8",X"91",X"9A",X"A5",X"9A",X"18",X"69",X"02",
		X"85",X"9C",X"A5",X"9B",X"69",X"00",X"85",X"9D",X"20",X"3A",X"C7",X"A9",X"00",X"D0",X"2A",X"A5",
		X"A6",X"A4",X"A7",X"85",X"A2",X"84",X"A3",X"A5",X"9C",X"A4",X"9D",X"85",X"9E",X"84",X"9F",X"85",
		X"A0",X"84",X"A1",X"20",X"52",X"C9",X"A2",X"88",X"86",X"85",X"68",X"A8",X"68",X"A2",X"FE",X"9A",
		X"48",X"98",X"48",X"A9",X"00",X"85",X"AD",X"85",X"2B",X"60",X"18",X"A5",X"9A",X"69",X"FF",X"85",
		X"E9",X"A5",X"9B",X"69",X"FF",X"85",X"EA",X"60",X"08",X"20",X"E2",X"CA",X"20",X"B3",X"C6",X"28",
		X"F0",X"14",X"20",X"E8",X"00",X"F0",X"15",X"C9",X"CD",X"D0",X"92",X"20",X"E2",X"00",X"F0",X"06",
		X"20",X"E2",X"CA",X"F0",X"07",X"60",X"A9",X"FF",X"85",X"33",X"85",X"34",X"A0",X"01",X"B1",X"CE",
		X"F0",X"4D",X"20",X"62",X"C9",X"C9",X"20",X"D0",X"0E",X"4E",X"DF",X"02",X"AD",X"DF",X"02",X"10",
		X"FB",X"20",X"62",X"C9",X"4E",X"DF",X"02",X"C8",X"B1",X"CE",X"AA",X"C8",X"B1",X"CE",X"C5",X"34",
		X"D0",X"04",X"E4",X"33",X"F0",X"02",X"B0",X"27",X"84",X"B8",X"48",X"20",X"F0",X"CB",X"68",X"20",
		X"C5",X"E0",X"A9",X"20",X"A4",X"B8",X"29",X"7F",X"20",X"D9",X"CC",X"C8",X"F0",X"11",X"B1",X"CE",
		X"D0",X"1E",X"A8",X"B1",X"CE",X"AA",X"C8",X"B1",X"CE",X"86",X"CE",X"85",X"CF",X"D0",X"AD",X"2C",
		X"F2",X"02",X"10",X"01",X"60",X"20",X"F0",X"CB",X"20",X"2F",X"C8",X"68",X"68",X"4C",X"A8",X"C4",
		X"10",X"D6",X"38",X"E9",X"7F",X"AA",X"84",X"B8",X"A0",X"00",X"A9",X"E9",X"85",X"18",X"A9",X"C0",
		X"85",X"19",X"CA",X"F0",X"0D",X"E6",X"18",X"D0",X"02",X"E6",X"19",X"B1",X"18",X"10",X"F6",X"4C",
		X"E2",X"C7",X"C8",X"B1",X"18",X"30",X"AD",X"20",X"D9",X"CC",X"4C",X"F2",X"C7",X"20",X"16",X"C8",
		X"4E",X"F2",X"02",X"20",X"E8",X"00",X"4C",X"48",X"C7",X"20",X"16",X"C8",X"20",X"E8",X"00",X"20",
		X"AB",X"CB",X"20",X"2F",X"C8",X"60",X"2C",X"F1",X"02",X"30",X"39",X"A5",X"30",X"8D",X"59",X"02",
		X"AD",X"58",X"02",X"85",X"30",X"38",X"6E",X"F1",X"02",X"AD",X"56",X"02",X"4C",X"44",X"C8",X"2C",
		X"F1",X"02",X"10",X"20",X"A5",X"30",X"8D",X"58",X"02",X"AD",X"59",X"02",X"85",X"30",X"4E",X"F1",
		X"02",X"AD",X"57",X"02",X"85",X"31",X"38",X"E9",X"08",X"B0",X"FB",X"49",X"FF",X"E9",X"06",X"18",
		X"65",X"31",X"85",X"32",X"60",X"A9",X"80",X"85",X"2B",X"20",X"1C",X"CB",X"20",X"C6",X"C3",X"D0",
		X"05",X"8A",X"69",X"0F",X"AA",X"9A",X"68",X"68",X"A9",X"09",X"20",X"37",X"C4",X"20",X"4E",X"CA",
		X"18",X"98",X"65",X"E9",X"48",X"A5",X"EA",X"69",X"00",X"48",X"A5",X"A9",X"48",X"A5",X"A8",X"48",
		X"A9",X"C3",X"20",X"67",X"D0",X"20",X"06",X"CF",X"20",X"03",X"CF",X"A5",X"D5",X"09",X"7F",X"25",
		X"D1",X"85",X"D1",X"A9",X"9E",X"A0",X"C8",X"85",X"91",X"84",X"92",X"4C",X"C0",X"CF",X"A9",X"81",
		X"A0",X"DC",X"20",X"7B",X"DE",X"20",X"E8",X"00",X"C9",X"CB",X"D0",X"06",X"20",X"E2",X"00",X"20",
		X"03",X"CF",X"20",X"13",X"DF",X"20",X"B1",X"CF",X"A5",X"B9",X"48",X"A5",X"B8",X"48",X"A9",X"8D",
		X"48",X"20",X"62",X"C9",X"A5",X"E9",X"A4",X"EA",X"F0",X"06",X"85",X"AC",X"84",X"AD",X"A0",X"00",
		X"B1",X"E9",X"D0",X"5B",X"4E",X"52",X"02",X"A0",X"02",X"B1",X"E9",X"18",X"D0",X"03",X"4C",X"8A",
		X"C9",X"C8",X"B1",X"E9",X"85",X"A8",X"C8",X"B1",X"E9",X"85",X"A9",X"98",X"65",X"E9",X"85",X"E9",
		X"90",X"02",X"E6",X"EA",X"2C",X"F4",X"02",X"10",X"13",X"48",X"A9",X"5B",X"20",X"FB",X"CC",X"A5",
		X"A9",X"A6",X"A8",X"20",X"C5",X"E0",X"A9",X"5D",X"20",X"FB",X"CC",X"68",X"20",X"E2",X"00",X"20",
		X"15",X"C9",X"4C",X"C1",X"C8",X"F0",X"49",X"E9",X"80",X"90",X"11",X"C9",X"42",X"B0",X"30",X"0A",
		X"A8",X"B9",X"07",X"C0",X"48",X"B9",X"06",X"C0",X"48",X"4C",X"E2",X"00",X"4C",X"1C",X"CB",X"C9",
		X"3A",X"F0",X"C1",X"C9",X"C8",X"D0",X"0E",X"2C",X"52",X"02",X"10",X"13",X"20",X"B1",X"CA",X"4E",
		X"52",X"02",X"4C",X"C1",X"C8",X"C9",X"27",X"D0",X"06",X"20",X"99",X"CA",X"4C",X"C1",X"C8",X"4C",
		X"70",X"D0",X"38",X"A5",X"9A",X"E9",X"01",X"A4",X"9B",X"B0",X"01",X"88",X"85",X"B0",X"84",X"B1",
		X"60",X"60",X"AD",X"DF",X"02",X"10",X"F9",X"29",X"7F",X"A2",X"08",X"C9",X"03",X"D0",X"F2",X"C9",
		X"03",X"B0",X"01",X"18",X"D0",X"43",X"A5",X"E9",X"A4",X"EA",X"F0",X"0C",X"85",X"AC",X"84",X"AD",
		X"A5",X"A8",X"A4",X"A9",X"85",X"AA",X"84",X"AB",X"68",X"68",X"A9",X"BD",X"A0",X"C3",X"A2",X"00",
		X"8E",X"F1",X"02",X"8E",X"DF",X"02",X"86",X"2E",X"90",X"03",X"4C",X"9D",X"C4",X"4C",X"A8",X"C4",
		X"D0",X"17",X"A2",X"D7",X"A4",X"AD",X"D0",X"03",X"4C",X"7E",X"C4",X"A5",X"AC",X"85",X"E9",X"84",
		X"EA",X"A5",X"AA",X"A4",X"AB",X"85",X"A8",X"84",X"A9",X"60",X"4C",X"36",X"D3",X"D0",X"03",X"4C",
		X"08",X"C7",X"20",X"0F",X"C7",X"4C",X"DC",X"C9",X"A9",X"03",X"20",X"37",X"C4",X"A5",X"EA",X"48",
		X"A5",X"E9",X"48",X"A5",X"A9",X"48",X"A5",X"A8",X"48",X"A9",X"9B",X"48",X"20",X"E8",X"00",X"20",
		X"E5",X"C9",X"4C",X"C1",X"C8",X"20",X"53",X"E8",X"20",X"51",X"CA",X"A5",X"A9",X"C5",X"34",X"B0",
		X"0B",X"98",X"38",X"65",X"E9",X"A6",X"EA",X"90",X"07",X"E8",X"B0",X"04",X"A5",X"9A",X"A6",X"9B",
		X"20",X"BD",X"C6",X"90",X"1E",X"A5",X"CE",X"E9",X"01",X"85",X"E9",X"A5",X"CF",X"E9",X"00",X"85",
		X"EA",X"60",X"D0",X"FD",X"A9",X"FF",X"85",X"B9",X"20",X"C6",X"C3",X"9A",X"C9",X"9B",X"F0",X"0B",
		X"A2",X"16",X"2C",X"A2",X"5A",X"4C",X"7E",X"C4",X"4C",X"70",X"D0",X"68",X"68",X"C0",X"0C",X"F0",
		X"19",X"85",X"A8",X"68",X"85",X"A9",X"68",X"85",X"E9",X"68",X"85",X"EA",X"20",X"4E",X"CA",X"98",
		X"18",X"65",X"E9",X"85",X"E9",X"90",X"02",X"E6",X"EA",X"60",X"68",X"68",X"68",X"60",X"A2",X"3A",
		X"2C",X"A2",X"00",X"86",X"24",X"A0",X"00",X"84",X"25",X"A5",X"25",X"A6",X"24",X"85",X"24",X"86",
		X"25",X"B1",X"E9",X"F0",X"E4",X"C5",X"25",X"F0",X"E0",X"C8",X"C9",X"22",X"D0",X"F3",X"F0",X"E9",
		X"20",X"17",X"CF",X"20",X"E8",X"00",X"C9",X"97",X"F0",X"05",X"A9",X"C9",X"20",X"67",X"D0",X"A5",
		X"D0",X"D0",X"05",X"20",X"9E",X"CA",X"F0",X"B7",X"20",X"E8",X"00",X"B0",X"03",X"4C",X"E5",X"C9",
		X"08",X"38",X"6E",X"52",X"02",X"28",X"4C",X"15",X"C9",X"20",X"51",X"CA",X"F0",X"A1",X"A0",X"00",
		X"B1",X"E9",X"F0",X"0C",X"C8",X"C9",X"C9",X"F0",X"F0",X"C9",X"C8",X"D0",X"F3",X"4C",X"3F",X"CA",
		X"60",X"A0",X"FF",X"C8",X"B1",X"E9",X"F0",X"04",X"C9",X"3A",X"D0",X"F7",X"4C",X"3F",X"CA",X"4C",
		X"70",X"D0",X"20",X"C8",X"D8",X"48",X"C9",X"9B",X"F0",X"04",X"C9",X"97",X"D0",X"F1",X"C6",X"D4",
		X"D0",X"04",X"68",X"4C",X"17",X"C9",X"20",X"E2",X"00",X"20",X"E2",X"CA",X"C9",X"2C",X"F0",X"EE",
		X"68",X"60",X"A2",X"00",X"86",X"33",X"86",X"34",X"B0",X"F7",X"E9",X"2F",X"85",X"24",X"A5",X"34",
		X"85",X"91",X"C9",X"19",X"B0",X"D4",X"A5",X"33",X"0A",X"26",X"91",X"0A",X"26",X"91",X"65",X"33",
		X"85",X"33",X"A5",X"91",X"65",X"34",X"85",X"34",X"06",X"33",X"26",X"34",X"A5",X"33",X"65",X"24",
		X"85",X"33",X"90",X"02",X"E6",X"34",X"20",X"E2",X"00",X"4C",X"E8",X"CA",X"20",X"88",X"D1",X"85",
		X"B8",X"84",X"B9",X"A9",X"D4",X"20",X"67",X"D0",X"A5",X"29",X"48",X"A5",X"28",X"48",X"20",X"17",
		X"CF",X"68",X"2A",X"20",X"09",X"CF",X"D0",X"18",X"68",X"10",X"12",X"20",X"F4",X"DE",X"20",X"A9",
		X"D2",X"A0",X"00",X"A5",X"D3",X"91",X"B8",X"C8",X"A5",X"D4",X"91",X"B8",X"60",X"4C",X"A9",X"DE",
		X"68",X"A0",X"02",X"B1",X"D3",X"C5",X"A3",X"90",X"17",X"D0",X"07",X"88",X"B1",X"D3",X"C5",X"A2",
		X"90",X"0E",X"A4",X"D4",X"C4",X"9D",X"90",X"08",X"D0",X"0D",X"A5",X"D3",X"C5",X"9C",X"B0",X"07",
		X"A5",X"D3",X"A4",X"D4",X"4C",X"8D",X"CB",X"A0",X"00",X"B1",X"D3",X"20",X"A3",X"D5",X"A5",X"BF",
		X"A4",X"C0",X"85",X"DE",X"84",X"DF",X"20",X"A4",X"D7",X"A9",X"D0",X"A0",X"00",X"85",X"BF",X"84",
		X"C0",X"20",X"05",X"D8",X"A0",X"00",X"B1",X"BF",X"91",X"B8",X"C8",X"B1",X"BF",X"91",X"B8",X"C8",
		X"B1",X"BF",X"91",X"B8",X"60",X"20",X"B3",X"CC",X"20",X"E8",X"00",X"F0",X"43",X"F0",X"5C",X"C9",
		X"C2",X"F0",X"7B",X"C9",X"C5",X"18",X"F0",X"76",X"C9",X"2C",X"F0",X"50",X"C9",X"3B",X"F0",X"6B",
		X"C9",X"C6",X"D0",X"03",X"4C",X"59",X"CC",X"20",X"17",X"CF",X"24",X"28",X"30",X"D7",X"20",X"D5",
		X"E0",X"20",X"B5",X"D5",X"A0",X"00",X"B1",X"D3",X"18",X"65",X"30",X"C5",X"31",X"90",X"03",X"20",
		X"F0",X"CB",X"20",X"B3",X"CC",X"20",X"D4",X"CC",X"D0",X"BE",X"A0",X"00",X"94",X"35",X"A2",X"34",
		X"A5",X"30",X"48",X"A9",X"0D",X"20",X"D9",X"CC",X"68",X"2C",X"F1",X"02",X"30",X"04",X"C5",X"31",
		X"F0",X"09",X"A9",X"00",X"85",X"30",X"A9",X"0A",X"20",X"D9",X"CC",X"60",X"A5",X"30",X"2C",X"F1",
		X"02",X"30",X"04",X"38",X"ED",X"53",X"02",X"38",X"E9",X"08",X"B0",X"FC",X"49",X"FF",X"69",X"01",
		X"AA",X"18",X"65",X"30",X"C5",X"31",X"90",X"1F",X"20",X"F0",X"CB",X"4C",X"4B",X"CC",X"08",X"20",
		X"C5",X"D8",X"C9",X"29",X"D0",X"20",X"28",X"90",X"0E",X"8A",X"C5",X"31",X"90",X"03",X"4C",X"36",
		X"D3",X"38",X"E5",X"30",X"90",X"05",X"AA",X"E8",X"CA",X"D0",X"06",X"20",X"E2",X"00",X"4C",X"AD",
		X"CB",X"20",X"D4",X"CC",X"D0",X"F2",X"4C",X"70",X"D0",X"2C",X"F1",X"02",X"30",X"F8",X"AE",X"1F",
		X"02",X"F0",X"03",X"4C",X"F7",X"EA",X"20",X"C5",X"D8",X"E0",X"28",X"B0",X"40",X"86",X"0C",X"20",
		X"65",X"D0",X"20",X"C8",X"D8",X"E8",X"E0",X"1C",X"B0",X"33",X"AD",X"6A",X"02",X"48",X"29",X"FE",
		X"8D",X"6A",X"02",X"A9",X"00",X"20",X"01",X"F8",X"A5",X"0C",X"8D",X"69",X"02",X"8A",X"8D",X"68",
		X"02",X"20",X"0C",X"DA",X"A5",X"1F",X"A4",X"20",X"85",X"12",X"84",X"13",X"68",X"8D",X"6A",X"02",
		X"A9",X"01",X"20",X"01",X"F8",X"A9",X"3B",X"20",X"67",X"D0",X"4C",X"AD",X"CB",X"4C",X"C2",X"D8",
		X"20",X"B5",X"D5",X"20",X"D0",X"D7",X"AA",X"A0",X"00",X"E8",X"CA",X"F0",X"10",X"B1",X"91",X"20",
		X"D9",X"CC",X"C8",X"C9",X"0D",X"D0",X"F3",X"20",X"0B",X"CC",X"4C",X"BA",X"CC",X"60",X"A9",X"0C",
		X"2C",X"A9",X"11",X"2C",X"A9",X"20",X"2C",X"A9",X"3F",X"24",X"2E",X"30",X"33",X"48",X"C9",X"20",
		X"90",X"0B",X"A5",X"30",X"C5",X"31",X"D0",X"03",X"20",X"F0",X"CB",X"E6",X"30",X"68",X"2C",X"F1",
		X"02",X"10",X"08",X"48",X"20",X"3E",X"02",X"68",X"29",X"FF",X"60",X"86",X"27",X"AA",X"20",X"38",
		X"02",X"C9",X"20",X"90",X"04",X"C9",X"7F",X"D0",X"05",X"AE",X"69",X"02",X"86",X"30",X"A6",X"27",
		X"29",X"FF",X"60",X"6C",X"F5",X"02",X"A9",X"80",X"2C",X"A9",X"00",X"8D",X"F4",X"02",X"60",X"A5",
		X"2C",X"F0",X"13",X"30",X"04",X"A0",X"FF",X"D0",X"04",X"A5",X"AE",X"A4",X"AF",X"85",X"A8",X"84",
		X"A9",X"A2",X"A8",X"4C",X"7E",X"C4",X"A9",X"85",X"A0",X"CE",X"20",X"B0",X"CC",X"A5",X"AC",X"A4",
		X"AD",X"85",X"E9",X"84",X"EA",X"60",X"20",X"D2",X"D4",X"A2",X"36",X"A0",X"00",X"84",X"36",X"A9",
		X"40",X"20",X"8F",X"CD",X"60",X"46",X"2E",X"C9",X"22",X"D0",X"0B",X"20",X"25",X"D0",X"A9",X"3B",
		X"20",X"67",X"D0",X"20",X"B3",X"CC",X"20",X"D2",X"D4",X"A9",X"2C",X"85",X"34",X"A9",X"00",X"85",
		X"17",X"20",X"80",X"CD",X"A5",X"35",X"D0",X"16",X"A5",X"17",X"F0",X"F1",X"18",X"4C",X"80",X"C9",
		X"20",X"D7",X"CC",X"20",X"D4",X"CC",X"4C",X"92",X"C5",X"A6",X"B0",X"A4",X"B1",X"A9",X"98",X"85",
		X"2C",X"86",X"B2",X"84",X"B3",X"20",X"88",X"D1",X"85",X"B8",X"84",X"B9",X"A5",X"E9",X"A4",X"EA",
		X"85",X"BA",X"84",X"BB",X"A6",X"B2",X"A4",X"B3",X"86",X"E9",X"84",X"EA",X"20",X"E8",X"00",X"D0",
		X"1D",X"24",X"2C",X"50",X"0D",X"20",X"78",X"EB",X"10",X"FB",X"85",X"35",X"A2",X"34",X"A0",X"00",
		X"F0",X"08",X"30",X"71",X"20",X"D7",X"CC",X"20",X"80",X"CD",X"86",X"E9",X"84",X"EA",X"20",X"E2",
		X"00",X"24",X"28",X"10",X"31",X"24",X"2C",X"50",X"09",X"E8",X"86",X"E9",X"A9",X"00",X"85",X"24",
		X"F0",X"0C",X"85",X"24",X"C9",X"22",X"F0",X"07",X"A9",X"3A",X"85",X"24",X"A9",X"2C",X"18",X"85",
		X"25",X"A5",X"E9",X"A4",X"EA",X"69",X"00",X"90",X"01",X"C8",X"20",X"BB",X"D5",X"20",X"0D",X"D9",
		X"20",X"51",X"CB",X"4C",X"0E",X"CE",X"20",X"E7",X"DF",X"A5",X"29",X"20",X"39",X"CB",X"20",X"E8",
		X"00",X"F0",X"07",X"C9",X"2C",X"F0",X"03",X"4C",X"1F",X"CD",X"A5",X"E9",X"A4",X"EA",X"85",X"B2",
		X"84",X"B3",X"A5",X"BA",X"A4",X"BB",X"85",X"E9",X"84",X"EA",X"20",X"E8",X"00",X"F0",X"2C",X"20",
		X"65",X"D0",X"4C",X"95",X"CD",X"20",X"4E",X"CA",X"C8",X"AA",X"D0",X"12",X"A2",X"2A",X"C8",X"B1",
		X"E9",X"F0",X"69",X"C8",X"B1",X"E9",X"85",X"AE",X"C8",X"B1",X"E9",X"C8",X"85",X"AF",X"B1",X"E9",
		X"AA",X"20",X"3F",X"CA",X"E0",X"91",X"D0",X"DD",X"4C",X"CE",X"CD",X"A5",X"B2",X"A4",X"B3",X"A6",
		X"2C",X"10",X"03",X"4C",X"5C",X"C9",X"A0",X"00",X"B1",X"B2",X"F0",X"07",X"A9",X"74",X"A0",X"CE",
		X"4C",X"B0",X"CC",X"60",X"3F",X"45",X"58",X"54",X"52",X"41",X"20",X"49",X"47",X"4E",X"4F",X"52",
		X"45",X"44",X"0D",X"0A",X"00",X"3F",X"52",X"45",X"44",X"4F",X"20",X"46",X"52",X"4F",X"4D",X"20",
		X"53",X"54",X"41",X"52",X"54",X"0D",X"0A",X"00",X"D0",X"04",X"A0",X"00",X"F0",X"03",X"20",X"88",
		X"D1",X"85",X"B8",X"84",X"B9",X"20",X"C6",X"C3",X"F0",X"04",X"A2",X"00",X"F0",X"66",X"9A",X"8A",
		X"18",X"69",X"04",X"48",X"69",X"06",X"85",X"93",X"68",X"A0",X"01",X"20",X"7B",X"DE",X"BA",X"BD",
		X"09",X"01",X"85",X"D5",X"A5",X"B8",X"A4",X"B9",X"20",X"22",X"DB",X"20",X"A9",X"DE",X"A0",X"01",
		X"20",X"4E",X"DF",X"BA",X"38",X"FD",X"09",X"01",X"F0",X"17",X"BD",X"0F",X"01",X"85",X"A8",X"BD",
		X"10",X"01",X"85",X"A9",X"BD",X"12",X"01",X"85",X"E9",X"BD",X"11",X"01",X"85",X"EA",X"4C",X"C1",
		X"C8",X"8A",X"69",X"11",X"AA",X"9A",X"20",X"E8",X"00",X"C9",X"2C",X"D0",X"F1",X"20",X"E2",X"00",
		X"20",X"9E",X"CE",X"20",X"17",X"CF",X"18",X"24",X"38",X"24",X"28",X"30",X"03",X"B0",X"03",X"60",
		X"B0",X"FD",X"A2",X"A8",X"4C",X"7E",X"C4",X"A6",X"E9",X"D0",X"02",X"C6",X"EA",X"C6",X"E9",X"A2",
		X"00",X"24",X"48",X"8A",X"48",X"A9",X"01",X"20",X"37",X"C4",X"20",X"00",X"D0",X"A9",X"00",X"85",
		X"BC",X"20",X"E8",X"00",X"38",X"E9",X"D3",X"90",X"17",X"C9",X"03",X"B0",X"13",X"C9",X"01",X"2A",
		X"49",X"01",X"45",X"BC",X"C5",X"BC",X"90",X"61",X"85",X"BC",X"20",X"E2",X"00",X"4C",X"34",X"CF",
		X"A6",X"BC",X"D0",X"2C",X"B0",X"7F",X"69",X"07",X"90",X"7B",X"65",X"28",X"D0",X"03",X"4C",X"67",
		X"D7",X"69",X"FF",X"85",X"91",X"0A",X"65",X"91",X"A8",X"68",X"D9",X"CC",X"C0",X"B0",X"6B",X"20",
		X"06",X"CF",X"48",X"20",X"99",X"CF",X"68",X"A4",X"BA",X"10",X"17",X"AA",X"F0",X"5A",X"D0",X"63",
		X"46",X"28",X"8A",X"2A",X"A6",X"E9",X"D0",X"02",X"C6",X"EA",X"C6",X"E9",X"A0",X"1B",X"85",X"BC",
		X"D0",X"D7",X"D9",X"CC",X"C0",X"B0",X"4C",X"90",X"D9",X"B9",X"CE",X"C0",X"48",X"B9",X"CD",X"C0",
		X"48",X"20",X"AC",X"CF",X"A5",X"BC",X"4C",X"22",X"CF",X"4C",X"70",X"D0",X"A5",X"D5",X"BE",X"CC",
		X"C0",X"A8",X"68",X"85",X"91",X"68",X"85",X"92",X"E6",X"91",X"D0",X"02",X"E6",X"92",X"98",X"48",
		X"20",X"F4",X"DE",X"A5",X"D4",X"48",X"A5",X"D3",X"48",X"A5",X"D2",X"48",X"A5",X"D1",X"48",X"A5",
		X"D0",X"48",X"6C",X"91",X"00",X"A0",X"FF",X"68",X"F0",X"23",X"C9",X"64",X"F0",X"03",X"20",X"06",
		X"CF",X"84",X"BA",X"68",X"4A",X"85",X"2D",X"68",X"85",X"D8",X"68",X"85",X"D9",X"68",X"85",X"DA",
		X"68",X"85",X"DB",X"68",X"85",X"DC",X"68",X"85",X"DD",X"45",X"D5",X"85",X"DE",X"A5",X"D0",X"60",
		X"A9",X"00",X"85",X"28",X"20",X"E2",X"00",X"B0",X"03",X"4C",X"E7",X"DF",X"20",X"16",X"D2",X"B0",
		X"6B",X"C9",X"2E",X"F0",X"F4",X"C9",X"23",X"F0",X"F0",X"C9",X"CD",X"F0",X"58",X"C9",X"CC",X"F0",
		X"E3",X"C9",X"22",X"D0",X"0F",X"A5",X"E9",X"A4",X"EA",X"69",X"00",X"90",X"01",X"C8",X"20",X"B5",
		X"D5",X"4C",X"0D",X"D9",X"C9",X"CA",X"D0",X"13",X"A0",X"18",X"D0",X"3B",X"20",X"A9",X"D2",X"A5",
		X"D4",X"49",X"FF",X"A8",X"A5",X"D3",X"49",X"FF",X"4C",X"99",X"D4",X"C9",X"C4",X"D0",X"03",X"4C",
		X"22",X"D5",X"C9",X"D6",X"90",X"03",X"4C",X"A0",X"D0",X"20",X"62",X"D0",X"20",X"17",X"CF",X"A9",
		X"29",X"2C",X"A9",X"28",X"2C",X"A9",X"2C",X"A0",X"00",X"D1",X"E9",X"D0",X"03",X"4C",X"E2",X"00",
		X"A2",X"10",X"4C",X"7E",X"C4",X"A0",X"15",X"68",X"68",X"4C",X"73",X"CF",X"20",X"88",X"D1",X"85",
		X"D3",X"84",X"D4",X"A6",X"28",X"F0",X"05",X"A2",X"00",X"86",X"DF",X"60",X"A6",X"29",X"10",X"0D",
		X"A0",X"00",X"B1",X"D3",X"AA",X"C8",X"B1",X"D3",X"A8",X"8A",X"4C",X"99",X"D4",X"4C",X"7B",X"DE",
		X"0A",X"48",X"AA",X"20",X"E2",X"00",X"E0",X"DB",X"90",X"24",X"E0",X"E7",X"90",X"23",X"20",X"62",
		X"D0",X"20",X"17",X"CF",X"20",X"65",X"D0",X"20",X"08",X"CF",X"68",X"AA",X"A5",X"D4",X"48",X"A5",
		X"D3",X"48",X"8A",X"48",X"20",X"C8",X"D8",X"68",X"A8",X"8A",X"48",X"4C",X"D3",X"D0",X"20",X"59",
		X"D0",X"68",X"A8",X"B9",X"DE",X"BF",X"85",X"C4",X"B9",X"DF",X"BF",X"85",X"C5",X"20",X"C3",X"00",
		X"4C",X"06",X"CF",X"A0",X"FF",X"2C",X"A0",X"00",X"84",X"26",X"20",X"A9",X"D2",X"A5",X"D3",X"45",
		X"26",X"85",X"24",X"A5",X"D4",X"45",X"26",X"85",X"25",X"20",X"D5",X"DE",X"20",X"A9",X"D2",X"A5",
		X"D4",X"45",X"26",X"25",X"25",X"45",X"26",X"A8",X"A5",X"D3",X"45",X"26",X"25",X"24",X"45",X"26",
		X"4C",X"99",X"D4",X"20",X"09",X"CF",X"B0",X"13",X"A5",X"DD",X"09",X"7F",X"25",X"D9",X"85",X"D9",
		X"A9",X"D8",X"A0",X"00",X"20",X"4C",X"DF",X"AA",X"4C",X"5E",X"D1",X"A9",X"00",X"85",X"28",X"C6",
		X"BC",X"20",X"D0",X"D7",X"85",X"D0",X"86",X"D1",X"84",X"D2",X"A5",X"DB",X"A4",X"DC",X"20",X"D4",
		X"D7",X"86",X"DB",X"84",X"DC",X"AA",X"38",X"E5",X"D0",X"F0",X"08",X"A9",X"01",X"90",X"04",X"A6",
		X"D0",X"A9",X"FF",X"85",X"D5",X"A0",X"FF",X"E8",X"C8",X"CA",X"D0",X"07",X"A6",X"D5",X"30",X"0F",
		X"18",X"90",X"0C",X"B1",X"DB",X"D1",X"D1",X"F0",X"EF",X"A2",X"FF",X"B0",X"02",X"A2",X"01",X"E8",
		X"8A",X"2A",X"25",X"2D",X"F0",X"02",X"A9",X"FF",X"4C",X"24",X"DF",X"20",X"65",X"D0",X"AA",X"20",
		X"8D",X"D1",X"20",X"E8",X"00",X"D0",X"F4",X"60",X"A2",X"00",X"20",X"E8",X"00",X"86",X"27",X"85",
		X"B4",X"20",X"E8",X"00",X"20",X"16",X"D2",X"B0",X"03",X"4C",X"70",X"D0",X"A2",X"00",X"86",X"28",
		X"86",X"29",X"20",X"E2",X"00",X"90",X"05",X"20",X"16",X"D2",X"90",X"0B",X"AA",X"20",X"E2",X"00",
		X"90",X"FB",X"20",X"16",X"D2",X"B0",X"F6",X"C9",X"24",X"D0",X"06",X"A9",X"FF",X"85",X"28",X"D0",
		X"10",X"C9",X"25",X"D0",X"13",X"A5",X"2B",X"30",X"D0",X"A9",X"80",X"85",X"29",X"05",X"B4",X"85",
		X"B4",X"8A",X"09",X"80",X"AA",X"20",X"E2",X"00",X"86",X"B5",X"38",X"05",X"2B",X"E9",X"28",X"D0",
		X"03",X"4C",X"BB",X"D2",X"24",X"2B",X"70",X"F9",X"A9",X"00",X"85",X"2B",X"A5",X"9C",X"A6",X"9D",
		X"A0",X"00",X"86",X"CF",X"85",X"CE",X"E4",X"9F",X"D0",X"04",X"C5",X"9E",X"F0",X"24",X"A5",X"B4",
		X"D1",X"CE",X"D0",X"08",X"A5",X"B5",X"C8",X"D1",X"CE",X"F0",X"6C",X"88",X"18",X"A5",X"CE",X"69",
		X"07",X"90",X"E1",X"E8",X"D0",X"DC",X"C9",X"41",X"90",X"07",X"E9",X"5B",X"38",X"E9",X"A5",X"B0",
		X"00",X"60",X"68",X"48",X"C9",X"7E",X"D0",X"0D",X"BA",X"BD",X"02",X"01",X"C9",X"D0",X"D0",X"05",
		X"A9",X"07",X"A0",X"E2",X"60",X"A5",X"9E",X"A4",X"9F",X"85",X"CE",X"84",X"CF",X"A5",X"A0",X"A4",
		X"A1",X"85",X"C9",X"84",X"CA",X"18",X"69",X"07",X"90",X"01",X"C8",X"85",X"C7",X"84",X"C8",X"20",
		X"F4",X"C3",X"A5",X"C7",X"A4",X"C8",X"C8",X"85",X"9E",X"84",X"9F",X"A0",X"00",X"A5",X"B4",X"91",
		X"CE",X"C8",X"A5",X"B5",X"91",X"CE",X"A9",X"00",X"C8",X"91",X"CE",X"C8",X"91",X"CE",X"C8",X"91",
		X"CE",X"C8",X"91",X"CE",X"C8",X"91",X"CE",X"A5",X"CE",X"18",X"69",X"02",X"A4",X"CF",X"90",X"01",
		X"C8",X"85",X"B6",X"84",X"B7",X"60",X"A5",X"26",X"0A",X"69",X"05",X"65",X"CE",X"A4",X"CF",X"90",
		X"01",X"C8",X"85",X"C7",X"84",X"C8",X"60",X"90",X"80",X"00",X"00",X"00",X"20",X"E2",X"00",X"20",
		X"17",X"CF",X"20",X"06",X"CF",X"A5",X"D5",X"30",X"0D",X"A5",X"D0",X"C9",X"90",X"90",X"09",X"A9",
		X"97",X"A0",X"D2",X"20",X"4C",X"DF",X"D0",X"7E",X"4C",X"8C",X"DF",X"A5",X"2B",X"D0",X"47",X"A5",
		X"27",X"05",X"29",X"48",X"A5",X"28",X"48",X"A0",X"00",X"98",X"48",X"A5",X"B5",X"48",X"A5",X"B4",
		X"48",X"20",X"9C",X"D2",X"68",X"85",X"B4",X"68",X"85",X"B5",X"68",X"A8",X"BA",X"BD",X"02",X"01",
		X"48",X"BD",X"01",X"01",X"48",X"A5",X"D3",X"9D",X"02",X"01",X"A5",X"D4",X"9D",X"01",X"01",X"C8",
		X"20",X"E8",X"00",X"C9",X"2C",X"F0",X"D2",X"84",X"26",X"20",X"5F",X"D0",X"68",X"85",X"28",X"68",
		X"85",X"29",X"29",X"7F",X"85",X"27",X"A6",X"9E",X"A5",X"9F",X"86",X"CE",X"85",X"CF",X"C5",X"A1",
		X"D0",X"04",X"E4",X"A0",X"F0",X"3F",X"A0",X"00",X"B1",X"CE",X"C8",X"C5",X"B4",X"D0",X"06",X"A5",
		X"B5",X"D1",X"CE",X"F0",X"16",X"C8",X"B1",X"CE",X"18",X"65",X"CE",X"AA",X"C8",X"B1",X"CE",X"65",
		X"CF",X"90",X"D7",X"A2",X"6B",X"2C",X"A2",X"35",X"4C",X"7E",X"C4",X"A2",X"78",X"A5",X"27",X"D0",
		X"F7",X"A5",X"2B",X"F0",X"02",X"38",X"60",X"20",X"86",X"D2",X"A5",X"26",X"A0",X"04",X"D1",X"CE",
		X"D0",X"E1",X"4C",X"EB",X"D3",X"A5",X"2B",X"F0",X"08",X"20",X"3D",X"E9",X"A2",X"2A",X"4C",X"7E",
		X"C4",X"20",X"86",X"D2",X"20",X"44",X"C4",X"A9",X"00",X"A8",X"85",X"E1",X"A2",X"05",X"A5",X"B4",
		X"91",X"CE",X"10",X"01",X"CA",X"C8",X"A5",X"B5",X"91",X"CE",X"10",X"02",X"CA",X"CA",X"86",X"E0",
		X"A5",X"26",X"C8",X"C8",X"C8",X"91",X"CE",X"A2",X"0B",X"A9",X"00",X"24",X"27",X"50",X"08",X"68",
		X"18",X"69",X"01",X"AA",X"68",X"69",X"00",X"C8",X"91",X"CE",X"C8",X"8A",X"91",X"CE",X"20",X"4D",
		X"D4",X"86",X"E0",X"85",X"E1",X"A4",X"91",X"C6",X"26",X"D0",X"DC",X"65",X"C8",X"B0",X"5D",X"85",
		X"C8",X"A8",X"8A",X"65",X"C7",X"90",X"03",X"C8",X"F0",X"52",X"20",X"44",X"C4",X"85",X"A0",X"84",
		X"A1",X"A9",X"00",X"E6",X"E1",X"A4",X"E0",X"F0",X"05",X"88",X"91",X"C7",X"D0",X"FB",X"C6",X"C8",
		X"C6",X"E1",X"D0",X"F5",X"E6",X"C8",X"38",X"A5",X"A0",X"E5",X"CE",X"A0",X"02",X"91",X"CE",X"A5",
		X"A1",X"C8",X"E5",X"CF",X"91",X"CE",X"A5",X"27",X"D0",X"62",X"C8",X"B1",X"CE",X"85",X"26",X"A9",
		X"00",X"85",X"E0",X"85",X"E1",X"C8",X"68",X"AA",X"85",X"D3",X"68",X"85",X"D4",X"D1",X"CE",X"90",
		X"0E",X"D0",X"06",X"C8",X"8A",X"D1",X"CE",X"90",X"07",X"4C",X"33",X"D3",X"4C",X"7C",X"C4",X"C8",
		X"A5",X"E1",X"05",X"E0",X"18",X"F0",X"0A",X"20",X"4D",X"D4",X"8A",X"65",X"D3",X"AA",X"98",X"A4",
		X"91",X"65",X"D4",X"86",X"E0",X"C6",X"26",X"D0",X"CA",X"85",X"E1",X"A2",X"05",X"A5",X"B4",X"10",
		X"01",X"CA",X"A5",X"B5",X"10",X"02",X"CA",X"CA",X"86",X"97",X"A9",X"00",X"20",X"56",X"D4",X"8A",
		X"65",X"C7",X"85",X"B6",X"98",X"65",X"C8",X"85",X"B7",X"A8",X"A5",X"B6",X"60",X"84",X"91",X"B1",
		X"CE",X"85",X"97",X"88",X"B1",X"CE",X"85",X"98",X"A9",X"10",X"85",X"CC",X"A2",X"00",X"A0",X"00",
		X"8A",X"0A",X"AA",X"98",X"2A",X"A8",X"B0",X"A4",X"06",X"E0",X"26",X"E1",X"90",X"0B",X"18",X"8A",
		X"65",X"97",X"AA",X"98",X"65",X"98",X"A8",X"B0",X"93",X"C6",X"CC",X"D0",X"E3",X"60",X"A5",X"28",
		X"F0",X"03",X"20",X"D0",X"D7",X"20",X"50",X"D6",X"38",X"A5",X"A2",X"E5",X"A0",X"A8",X"A5",X"A3",
		X"E5",X"A1",X"A2",X"00",X"86",X"28",X"4C",X"40",X"DF",X"A2",X"00",X"86",X"28",X"85",X"D1",X"84",
		X"D2",X"A2",X"90",X"4C",X"2C",X"DF",X"20",X"CB",X"D8",X"8A",X"F0",X"08",X"AC",X"58",X"02",X"2C",
		X"F1",X"02",X"10",X"02",X"A4",X"30",X"A9",X"00",X"F0",X"DF",X"C9",X"D9",X"D0",X"21",X"20",X"E2",
		X"00",X"A9",X"D4",X"20",X"67",X"D0",X"20",X"53",X"E8",X"A5",X"33",X"A4",X"34",X"85",X"22",X"84",
		X"23",X"60",X"A6",X"A9",X"E8",X"D0",X"FA",X"A2",X"95",X"2C",X"A2",X"E5",X"4C",X"7E",X"C4",X"20",
		X"0D",X"D5",X"20",X"D2",X"D4",X"20",X"62",X"D0",X"A9",X"80",X"85",X"2B",X"20",X"88",X"D1",X"20",
		X"06",X"CF",X"20",X"5F",X"D0",X"A9",X"D4",X"20",X"67",X"D0",X"48",X"A5",X"B7",X"48",X"A5",X"B6",
		X"48",X"A5",X"EA",X"48",X"A5",X"E9",X"48",X"20",X"3C",X"CA",X"4C",X"7D",X"D5",X"A9",X"C4",X"20",
		X"67",X"D0",X"09",X"80",X"A2",X"80",X"86",X"2B",X"20",X"8F",X"D1",X"85",X"BD",X"84",X"BE",X"4C",
		X"06",X"CF",X"20",X"0D",X"D5",X"A5",X"BE",X"48",X"A5",X"BD",X"48",X"20",X"59",X"D0",X"20",X"06",
		X"CF",X"68",X"85",X"BD",X"68",X"85",X"BE",X"A0",X"02",X"B1",X"BD",X"85",X"B6",X"AA",X"C8",X"B1",
		X"BD",X"F0",X"97",X"85",X"B7",X"C8",X"B1",X"B6",X"48",X"88",X"10",X"FA",X"A4",X"B7",X"20",X"AD",
		X"DE",X"A5",X"EA",X"48",X"A5",X"E9",X"48",X"B1",X"BD",X"85",X"E9",X"C8",X"B1",X"BD",X"85",X"EA",
		X"A5",X"B7",X"48",X"A5",X"B6",X"48",X"20",X"03",X"CF",X"68",X"85",X"BD",X"68",X"85",X"BE",X"20",
		X"E8",X"00",X"F0",X"03",X"4C",X"70",X"D0",X"68",X"85",X"E9",X"68",X"85",X"EA",X"A0",X"00",X"68",
		X"91",X"BD",X"68",X"C8",X"91",X"BD",X"68",X"C8",X"91",X"BD",X"68",X"C8",X"91",X"BD",X"68",X"C8",
		X"91",X"BD",X"60",X"20",X"06",X"CF",X"A0",X"00",X"20",X"D7",X"E0",X"68",X"68",X"A9",X"FF",X"A0",
		X"00",X"F0",X"12",X"A6",X"D3",X"A4",X"D4",X"86",X"BF",X"84",X"C0",X"20",X"1E",X"D6",X"86",X"D1",
		X"84",X"D2",X"85",X"D0",X"60",X"A2",X"22",X"86",X"24",X"86",X"25",X"85",X"DE",X"84",X"DF",X"85",
		X"D1",X"84",X"D2",X"A0",X"FF",X"C8",X"B1",X"DE",X"F0",X"0C",X"C5",X"24",X"F0",X"04",X"C5",X"25",
		X"D0",X"F3",X"C9",X"22",X"F0",X"01",X"18",X"84",X"D0",X"98",X"65",X"DE",X"85",X"E0",X"A6",X"DF",
		X"90",X"01",X"E8",X"86",X"E1",X"A5",X"DF",X"D0",X"0B",X"98",X"20",X"A3",X"D5",X"A6",X"DE",X"A4",
		X"DF",X"20",X"B2",X"D7",X"A6",X"85",X"E0",X"91",X"D0",X"05",X"A2",X"C4",X"4C",X"7E",X"C4",X"A5",
		X"D0",X"95",X"00",X"A5",X"D1",X"95",X"01",X"A5",X"D2",X"95",X"02",X"A0",X"00",X"86",X"D3",X"84",
		X"D4",X"84",X"DF",X"88",X"84",X"28",X"86",X"86",X"E8",X"E8",X"E8",X"86",X"85",X"60",X"46",X"2A",
		X"48",X"49",X"FF",X"38",X"65",X"A2",X"A4",X"A3",X"B0",X"01",X"88",X"C4",X"A1",X"90",X"11",X"D0",
		X"04",X"C5",X"A0",X"90",X"0B",X"85",X"A2",X"84",X"A3",X"85",X"A4",X"84",X"A5",X"AA",X"68",X"60",
		X"A2",X"4D",X"A5",X"2A",X"30",X"B6",X"20",X"50",X"D6",X"A9",X"80",X"85",X"2A",X"68",X"D0",X"D0",
		X"A6",X"A6",X"A5",X"A7",X"86",X"A2",X"85",X"A3",X"A0",X"00",X"84",X"BE",X"84",X"BD",X"A5",X"A0",
		X"A6",X"A1",X"85",X"CE",X"86",X"CF",X"A9",X"88",X"A2",X"00",X"85",X"91",X"86",X"92",X"C5",X"85",
		X"F0",X"05",X"20",X"F1",X"D6",X"F0",X"F7",X"A9",X"07",X"85",X"C2",X"A5",X"9C",X"A6",X"9D",X"85",
		X"91",X"86",X"92",X"E4",X"9F",X"D0",X"04",X"C5",X"9E",X"F0",X"05",X"20",X"E7",X"D6",X"F0",X"F3",
		X"85",X"C7",X"86",X"C8",X"A9",X"03",X"85",X"C2",X"A5",X"C7",X"A6",X"C8",X"E4",X"A1",X"D0",X"07",
		X"C5",X"A0",X"D0",X"03",X"4C",X"30",X"D7",X"85",X"91",X"86",X"92",X"A0",X"00",X"B1",X"91",X"AA",
		X"C8",X"B1",X"91",X"08",X"C8",X"B1",X"91",X"65",X"C7",X"85",X"C7",X"C8",X"B1",X"91",X"65",X"C8",
		X"85",X"C8",X"28",X"10",X"D3",X"8A",X"30",X"D0",X"C8",X"B1",X"91",X"A0",X"00",X"0A",X"69",X"05",
		X"65",X"91",X"85",X"91",X"90",X"02",X"E6",X"92",X"A6",X"92",X"E4",X"C8",X"D0",X"04",X"C5",X"C7",
		X"F0",X"BA",X"20",X"F1",X"D6",X"F0",X"F3",X"B1",X"91",X"30",X"35",X"C8",X"B1",X"91",X"10",X"30",
		X"C8",X"B1",X"91",X"F0",X"2B",X"C8",X"B1",X"91",X"AA",X"C8",X"B1",X"91",X"C5",X"A3",X"90",X"06",
		X"D0",X"1E",X"E4",X"A2",X"B0",X"1A",X"C5",X"CF",X"90",X"16",X"D0",X"04",X"E4",X"CE",X"90",X"10",
		X"86",X"CE",X"85",X"CF",X"A5",X"91",X"A6",X"92",X"85",X"BD",X"86",X"BE",X"A5",X"C2",X"85",X"C4",
		X"A5",X"C2",X"18",X"65",X"91",X"85",X"91",X"90",X"02",X"E6",X"92",X"A6",X"92",X"A0",X"00",X"60",
		X"A5",X"BE",X"05",X"BD",X"F0",X"F5",X"A5",X"C4",X"29",X"04",X"4A",X"A8",X"85",X"C4",X"B1",X"BD",
		X"65",X"CE",X"85",X"C9",X"A5",X"CF",X"69",X"00",X"85",X"CA",X"A5",X"A2",X"A6",X"A3",X"85",X"C7",
		X"86",X"C8",X"20",X"FB",X"C3",X"A4",X"C4",X"C8",X"A5",X"C7",X"91",X"BD",X"AA",X"E6",X"C8",X"A5",
		X"C8",X"C8",X"91",X"BD",X"4C",X"54",X"D6",X"A5",X"D4",X"48",X"A5",X"D3",X"48",X"20",X"00",X"D0",
		X"20",X"08",X"CF",X"68",X"85",X"DE",X"68",X"85",X"DF",X"A0",X"00",X"B1",X"DE",X"18",X"71",X"D3",
		X"90",X"05",X"A2",X"B5",X"4C",X"7E",X"C4",X"20",X"A3",X"D5",X"20",X"A4",X"D7",X"A5",X"BF",X"A4",
		X"C0",X"20",X"D4",X"D7",X"20",X"B6",X"D7",X"A5",X"DE",X"A4",X"DF",X"20",X"D4",X"D7",X"20",X"F4",
		X"D5",X"4C",X"31",X"CF",X"A0",X"00",X"B1",X"DE",X"48",X"C8",X"B1",X"DE",X"AA",X"C8",X"B1",X"DE",
		X"A8",X"68",X"86",X"91",X"84",X"92",X"A8",X"F0",X"0A",X"48",X"88",X"B1",X"91",X"91",X"A4",X"98",
		X"D0",X"F8",X"68",X"18",X"65",X"A4",X"85",X"A4",X"90",X"02",X"E6",X"A5",X"60",X"20",X"08",X"CF",
		X"A5",X"D3",X"A4",X"D4",X"85",X"91",X"84",X"92",X"20",X"05",X"D8",X"08",X"A0",X"00",X"B1",X"91",
		X"48",X"C8",X"B1",X"91",X"AA",X"C8",X"B1",X"91",X"A8",X"68",X"28",X"D0",X"13",X"C4",X"A3",X"D0",
		X"0F",X"E4",X"A2",X"D0",X"0B",X"48",X"18",X"65",X"A2",X"85",X"A2",X"90",X"02",X"E6",X"A3",X"68",
		X"86",X"91",X"84",X"92",X"60",X"C4",X"87",X"D0",X"0C",X"C5",X"86",X"D0",X"08",X"85",X"85",X"E9",
		X"03",X"85",X"86",X"A0",X"00",X"60",X"20",X"CB",X"D8",X"8A",X"48",X"A9",X"01",X"20",X"AB",X"D5",
		X"68",X"A0",X"00",X"91",X"D1",X"68",X"68",X"4C",X"F4",X"D5",X"20",X"8B",X"D8",X"D1",X"BF",X"98",
		X"90",X"04",X"B1",X"BF",X"AA",X"98",X"48",X"8A",X"48",X"20",X"AB",X"D5",X"A5",X"BF",X"A4",X"C0",
		X"20",X"D4",X"D7",X"68",X"A8",X"68",X"18",X"65",X"91",X"85",X"91",X"90",X"02",X"E6",X"92",X"98",
		X"20",X"B6",X"D7",X"4C",X"F4",X"D5",X"20",X"8B",X"D8",X"18",X"F1",X"BF",X"49",X"FF",X"4C",X"30",
		X"D8",X"A9",X"FF",X"85",X"D4",X"20",X"E8",X"00",X"C9",X"29",X"F0",X"06",X"20",X"65",X"D0",X"20",
		X"C8",X"D8",X"20",X"8B",X"D8",X"F0",X"4B",X"CA",X"8A",X"48",X"18",X"A2",X"00",X"F1",X"BF",X"B0",
		X"B6",X"49",X"FF",X"C5",X"D4",X"90",X"B1",X"A5",X"D4",X"B0",X"AD",X"20",X"5F",X"D0",X"68",X"A8",
		X"68",X"85",X"C4",X"68",X"68",X"68",X"AA",X"68",X"85",X"BF",X"68",X"85",X"C0",X"A5",X"C4",X"48",
		X"98",X"48",X"A0",X"00",X"8A",X"60",X"20",X"AC",X"D8",X"4C",X"B6",X"D4",X"20",X"CD",X"D7",X"A2",
		X"00",X"86",X"28",X"A8",X"60",X"20",X"AC",X"D8",X"F0",X"08",X"A0",X"00",X"B1",X"91",X"A8",X"4C",
		X"B6",X"D4",X"4C",X"36",X"D3",X"20",X"E2",X"00",X"20",X"03",X"CF",X"20",X"A2",X"D2",X"A6",X"D3",
		X"D0",X"F0",X"A6",X"D4",X"4C",X"E8",X"00",X"20",X"AC",X"D8",X"D0",X"03",X"4C",X"B2",X"DB",X"A6",
		X"E9",X"A4",X"EA",X"86",X"E0",X"84",X"E1",X"A6",X"91",X"86",X"E9",X"18",X"65",X"91",X"85",X"93",
		X"A6",X"92",X"86",X"EA",X"90",X"01",X"E8",X"86",X"94",X"A0",X"00",X"B1",X"93",X"48",X"A9",X"00",
		X"91",X"93",X"20",X"E8",X"00",X"20",X"E7",X"DF",X"68",X"A0",X"00",X"91",X"93",X"A6",X"E0",X"A4",
		X"E1",X"86",X"E9",X"84",X"EA",X"60",X"20",X"03",X"CF",X"20",X"22",X"D9",X"20",X"65",X"D0",X"4C",
		X"C8",X"D8",X"A5",X"D5",X"30",X"9C",X"A5",X"D0",X"C9",X"91",X"B0",X"96",X"20",X"8C",X"DF",X"A5",
		X"D3",X"A4",X"D4",X"84",X"33",X"85",X"34",X"60",X"A5",X"34",X"48",X"A5",X"33",X"48",X"20",X"22",
		X"D9",X"A0",X"00",X"B1",X"33",X"A8",X"68",X"85",X"33",X"68",X"85",X"34",X"4C",X"B6",X"D4",X"20",
		X"16",X"D9",X"8A",X"A0",X"00",X"91",X"33",X"60",X"20",X"03",X"CF",X"20",X"22",X"D9",X"A4",X"33",
		X"A6",X"34",X"A9",X"02",X"4C",X"C9",X"EE",X"20",X"53",X"E8",X"A5",X"33",X"A4",X"34",X"85",X"1D",
		X"84",X"1E",X"20",X"65",X"D0",X"20",X"53",X"E8",X"A0",X"01",X"B9",X"33",X"00",X"91",X"1D",X"88",
		X"10",X"F8",X"60",X"20",X"22",X"D9",X"A0",X"01",X"B1",X"33",X"48",X"88",X"B1",X"33",X"A8",X"68",
		X"4C",X"40",X"DF",X"48",X"4A",X"4A",X"4A",X"4A",X"20",X"9C",X"D9",X"68",X"29",X"0F",X"09",X"30",
		X"C9",X"3A",X"90",X"02",X"69",X"06",X"C9",X"30",X"D0",X"04",X"A4",X"2F",X"F0",X"06",X"85",X"2F",
		X"9D",X"00",X"01",X"E8",X"60",X"20",X"22",X"D9",X"A2",X"00",X"86",X"2F",X"A9",X"23",X"85",X"FF",
		X"A5",X"34",X"20",X"93",X"D9",X"A5",X"33",X"20",X"93",X"D9",X"8A",X"D0",X"06",X"A9",X"30",X"9D",
		X"00",X"01",X"E8",X"A9",X"00",X"9D",X"00",X"01",X"4C",X"9B",X"D5",X"4C",X"70",X"D0",X"20",X"21",
		X"EC",X"20",X"C8",X"D8",X"8A",X"F0",X"06",X"CA",X"D0",X"F1",X"A9",X"09",X"2C",X"A9",X"08",X"A2",
		X"10",X"8E",X"F8",X"02",X"A2",X"1B",X"48",X"8A",X"20",X"0C",X"DA",X"AD",X"F8",X"02",X"A0",X"27",
		X"91",X"1F",X"88",X"D0",X"FB",X"68",X"91",X"1F",X"CA",X"D0",X"EB",X"60",X"20",X"31",X"F7",X"84",
		X"20",X"18",X"69",X"80",X"48",X"85",X"1F",X"A9",X"BB",X"65",X"20",X"85",X"20",X"68",X"60",X"4C",
		X"C2",X"D8",X"20",X"F6",X"DA",X"20",X"C8",X"D8",X"E0",X"28",X"B0",X"F3",X"8E",X"F8",X"02",X"20",
		X"65",X"D0",X"20",X"C8",X"D8",X"E0",X"1B",X"B0",X"E6",X"E8",X"8A",X"20",X"0C",X"DA",X"60",X"20",
		X"62",X"D0",X"20",X"22",X"DA",X"20",X"5F",X"D0",X"AC",X"F8",X"02",X"B1",X"1F",X"A8",X"4C",X"B6",
		X"D4",X"20",X"22",X"DA",X"20",X"65",X"D0",X"20",X"17",X"CF",X"24",X"28",X"10",X"1D",X"20",X"D0",
		X"D7",X"AA",X"18",X"AD",X"F8",X"02",X"65",X"1F",X"90",X"02",X"E6",X"20",X"85",X"1F",X"A0",X"00",
		X"E8",X"CA",X"F0",X"10",X"B1",X"91",X"91",X"1F",X"C8",X"D0",X"F6",X"20",X"CB",X"D8",X"8A",X"AC",
		X"F8",X"02",X"91",X"1F",X"60",X"D0",X"17",X"A9",X"03",X"20",X"37",X"C4",X"A5",X"EA",X"48",X"A5",
		X"E9",X"48",X"A5",X"A9",X"48",X"A5",X"A8",X"48",X"A9",X"8B",X"48",X"4C",X"C1",X"C8",X"4C",X"70",
		X"D0",X"A9",X"FF",X"85",X"B9",X"20",X"C6",X"C3",X"9A",X"C9",X"8B",X"F0",X"05",X"A2",X"F5",X"4C",
		X"7E",X"C4",X"C0",X"10",X"D0",X"05",X"84",X"D0",X"98",X"D0",X"06",X"20",X"E8",X"00",X"20",X"17",
		X"CF",X"68",X"A5",X"D0",X"F0",X"05",X"68",X"68",X"68",X"68",X"60",X"68",X"85",X"A8",X"68",X"85",
		X"A9",X"68",X"85",X"E9",X"68",X"85",X"EA",X"4C",X"8C",X"DA",X"20",X"78",X"EB",X"08",X"48",X"10",
		X"03",X"A9",X"01",X"2C",X"A9",X"00",X"20",X"AB",X"D5",X"68",X"28",X"10",X"04",X"A0",X"00",X"91",
		X"D1",X"68",X"68",X"4C",X"F4",X"D5",X"AD",X"C0",X"02",X"29",X"01",X"F0",X"05",X"A2",X"A3",X"4C",
		X"7E",X"C4",X"60",X"60",X"A9",X"05",X"A0",X"E2",X"4C",X"22",X"DB",X"20",X"51",X"DD",X"A5",X"D5",
		X"49",X"FF",X"85",X"D5",X"45",X"DD",X"85",X"DE",X"A5",X"D0",X"4C",X"25",X"DB",X"20",X"54",X"DC",
		X"90",X"3C",X"20",X"51",X"DD",X"D0",X"03",X"4C",X"D5",X"DE",X"A6",X"DF",X"86",X"C5",X"A2",X"D8",
		X"A5",X"D8",X"A8",X"F0",X"CE",X"38",X"E5",X"D0",X"F0",X"24",X"90",X"12",X"84",X"D0",X"A4",X"DD",
		X"84",X"D5",X"49",X"FF",X"69",X"00",X"A0",X"00",X"84",X"C5",X"A2",X"D0",X"D0",X"04",X"A0",X"00",
		X"84",X"DF",X"C9",X"F9",X"30",X"C7",X"A8",X"A5",X"DF",X"56",X"01",X"20",X"6B",X"DC",X"24",X"DE",
		X"10",X"57",X"A0",X"D0",X"E0",X"D8",X"F0",X"02",X"A0",X"D8",X"38",X"49",X"FF",X"65",X"C5",X"85",
		X"DF",X"B9",X"04",X"00",X"F5",X"04",X"85",X"D4",X"B9",X"03",X"00",X"F5",X"03",X"85",X"D3",X"B9",
		X"02",X"00",X"F5",X"02",X"85",X"D2",X"B9",X"01",X"00",X"F5",X"01",X"85",X"D1",X"B0",X"03",X"20",
		X"02",X"DC",X"A0",X"00",X"98",X"18",X"A6",X"D1",X"D0",X"4A",X"A6",X"D2",X"86",X"D1",X"A6",X"D3",
		X"86",X"D2",X"A6",X"D4",X"86",X"D3",X"A6",X"DF",X"86",X"D4",X"84",X"DF",X"69",X"08",X"C9",X"28",
		X"D0",X"E4",X"A9",X"00",X"85",X"D0",X"85",X"D5",X"60",X"65",X"C5",X"85",X"DF",X"A5",X"D4",X"65",
		X"DC",X"85",X"D4",X"A5",X"D3",X"65",X"DB",X"85",X"D3",X"A5",X"D2",X"65",X"DA",X"85",X"D2",X"A5",
		X"D1",X"65",X"D9",X"85",X"D1",X"4C",X"F1",X"DB",X"69",X"01",X"06",X"DF",X"26",X"D4",X"26",X"D3",
		X"26",X"D2",X"26",X"D1",X"10",X"F2",X"38",X"E5",X"D0",X"B0",X"C7",X"49",X"FF",X"69",X"01",X"85",
		X"D0",X"90",X"0E",X"E6",X"D0",X"F0",X"42",X"66",X"D1",X"66",X"D2",X"66",X"D3",X"66",X"D4",X"66",
		X"DF",X"60",X"A5",X"D5",X"49",X"FF",X"85",X"D5",X"A5",X"D1",X"49",X"FF",X"85",X"D1",X"A5",X"D2",
		X"49",X"FF",X"85",X"D2",X"A5",X"D3",X"49",X"FF",X"85",X"D3",X"A5",X"D4",X"49",X"FF",X"85",X"D4",
		X"A5",X"DF",X"49",X"FF",X"85",X"DF",X"E6",X"DF",X"D0",X"0E",X"E6",X"D4",X"D0",X"0A",X"E6",X"D3",
		X"D0",X"06",X"E6",X"D2",X"D0",X"02",X"E6",X"D1",X"60",X"A2",X"45",X"4C",X"7E",X"C4",X"A2",X"94",
		X"B4",X"04",X"84",X"DF",X"B4",X"03",X"94",X"04",X"B4",X"02",X"94",X"03",X"B4",X"01",X"94",X"02",
		X"A4",X"D7",X"94",X"01",X"69",X"08",X"30",X"E8",X"F0",X"E6",X"E9",X"08",X"A8",X"A5",X"DF",X"B0",
		X"14",X"16",X"01",X"90",X"02",X"F6",X"01",X"76",X"01",X"76",X"01",X"76",X"02",X"76",X"03",X"76",
		X"04",X"6A",X"C8",X"D0",X"EC",X"18",X"60",X"82",X"13",X"5D",X"8D",X"DE",X"82",X"49",X"0F",X"DA",
		X"9E",X"81",X"00",X"00",X"00",X"00",X"03",X"7F",X"5E",X"56",X"CB",X"79",X"80",X"13",X"9B",X"0B",
		X"64",X"80",X"76",X"38",X"93",X"16",X"82",X"38",X"AA",X"3B",X"20",X"80",X"35",X"04",X"F3",X"34",
		X"81",X"35",X"04",X"F3",X"34",X"80",X"80",X"00",X"00",X"00",X"80",X"31",X"72",X"17",X"F8",X"20",
		X"13",X"DF",X"F0",X"02",X"10",X"03",X"4C",X"36",X"D3",X"A5",X"D0",X"E9",X"7F",X"48",X"A9",X"80",
		X"85",X"D0",X"A9",X"9B",X"A0",X"DC",X"20",X"22",X"DB",X"A9",X"A0",X"A0",X"DC",X"20",X"E4",X"DD",
		X"A9",X"81",X"A0",X"DC",X"20",X"0B",X"DB",X"A9",X"86",X"A0",X"DC",X"20",X"FD",X"E2",X"A9",X"A5",
		X"A0",X"DC",X"20",X"22",X"DB",X"68",X"20",X"76",X"E0",X"A9",X"AA",X"A0",X"DC",X"20",X"51",X"DD",
		X"D0",X"03",X"4C",X"50",X"DD",X"20",X"7C",X"DD",X"A9",X"00",X"85",X"95",X"85",X"96",X"85",X"97",
		X"85",X"98",X"A5",X"DF",X"20",X"1E",X"DD",X"A5",X"D4",X"20",X"1E",X"DD",X"A5",X"D3",X"20",X"1E",
		X"DD",X"A5",X"D2",X"20",X"1E",X"DD",X"A5",X"D1",X"20",X"23",X"DD",X"4C",X"64",X"DE",X"D0",X"03",
		X"4C",X"3E",X"DC",X"4A",X"09",X"80",X"A8",X"90",X"19",X"18",X"A5",X"98",X"65",X"DC",X"85",X"98",
		X"A5",X"97",X"65",X"DB",X"85",X"97",X"A5",X"96",X"65",X"DA",X"85",X"96",X"A5",X"95",X"65",X"D9",
		X"85",X"95",X"66",X"95",X"66",X"96",X"66",X"97",X"66",X"98",X"66",X"DF",X"98",X"4A",X"D0",X"D6",
		X"60",X"85",X"91",X"84",X"92",X"A0",X"04",X"B1",X"91",X"85",X"DC",X"88",X"B1",X"91",X"85",X"DB",
		X"88",X"B1",X"91",X"85",X"DA",X"88",X"B1",X"91",X"85",X"DD",X"45",X"D5",X"85",X"DE",X"A5",X"DD",
		X"09",X"80",X"85",X"D9",X"88",X"B1",X"91",X"85",X"D8",X"A5",X"D0",X"60",X"A5",X"D8",X"F0",X"1F",
		X"18",X"65",X"D0",X"90",X"04",X"30",X"1D",X"18",X"2C",X"10",X"14",X"69",X"80",X"85",X"D0",X"D0",
		X"03",X"4C",X"B6",X"DB",X"A5",X"DE",X"85",X"D5",X"60",X"A5",X"D5",X"49",X"FF",X"30",X"05",X"68",
		X"68",X"4C",X"B2",X"DB",X"4C",X"39",X"DC",X"20",X"E5",X"DE",X"AA",X"F0",X"10",X"18",X"69",X"02",
		X"B0",X"F2",X"A2",X"00",X"86",X"DE",X"20",X"32",X"DB",X"E6",X"D0",X"F0",X"E7",X"60",X"84",X"20",
		X"00",X"00",X"00",X"20",X"E5",X"DE",X"A9",X"BE",X"A0",X"DD",X"A2",X"00",X"86",X"DE",X"20",X"7B",
		X"DE",X"4C",X"E7",X"DD",X"20",X"AF",X"DC",X"20",X"E5",X"DE",X"A9",X"77",X"A0",X"DC",X"20",X"7B",
		X"DE",X"4C",X"E7",X"DD",X"20",X"51",X"DD",X"F0",X"76",X"20",X"F4",X"DE",X"A9",X"00",X"38",X"E5",
		X"D0",X"85",X"D0",X"20",X"7C",X"DD",X"E6",X"D0",X"F0",X"AA",X"A2",X"FC",X"A9",X"01",X"A4",X"D9",
		X"C4",X"D1",X"D0",X"10",X"A4",X"DA",X"C4",X"D2",X"D0",X"0A",X"A4",X"DB",X"C4",X"D3",X"D0",X"04",
		X"A4",X"DC",X"C4",X"D4",X"08",X"2A",X"90",X"09",X"E8",X"95",X"98",X"F0",X"32",X"10",X"34",X"A9",
		X"01",X"28",X"B0",X"0E",X"06",X"DC",X"26",X"DB",X"26",X"DA",X"26",X"D9",X"B0",X"E6",X"30",X"CE",
		X"10",X"E2",X"A8",X"A5",X"DC",X"E5",X"D4",X"85",X"DC",X"A5",X"DB",X"E5",X"D3",X"85",X"DB",X"A5",
		X"DA",X"E5",X"D2",X"85",X"DA",X"A5",X"D9",X"E5",X"D1",X"85",X"D9",X"98",X"4C",X"24",X"DE",X"A9",
		X"40",X"D0",X"CE",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"85",X"DF",X"28",X"4C",X"64",X"DE",X"A2",
		X"85",X"4C",X"7E",X"C4",X"A5",X"95",X"85",X"D1",X"A5",X"96",X"85",X"D2",X"A5",X"97",X"85",X"D3",
		X"A5",X"98",X"85",X"D4",X"4C",X"92",X"DB",X"A9",X"7C",X"A0",X"DC",X"85",X"91",X"84",X"92",X"A0",
		X"04",X"B1",X"91",X"85",X"D4",X"88",X"B1",X"91",X"85",X"D3",X"88",X"B1",X"91",X"85",X"D2",X"88",
		X"B1",X"91",X"85",X"D5",X"09",X"80",X"85",X"D1",X"88",X"B1",X"91",X"85",X"D0",X"84",X"DF",X"60",
		X"A2",X"CB",X"2C",X"A2",X"C6",X"A0",X"00",X"F0",X"04",X"A6",X"B8",X"A4",X"B9",X"20",X"F4",X"DE",
		X"86",X"91",X"84",X"92",X"A0",X"04",X"A5",X"D4",X"91",X"91",X"88",X"A5",X"D3",X"91",X"91",X"88",
		X"A5",X"D2",X"91",X"91",X"88",X"A5",X"D5",X"09",X"7F",X"25",X"D1",X"91",X"91",X"88",X"A5",X"D0",
		X"91",X"91",X"84",X"DF",X"60",X"A5",X"DD",X"85",X"D5",X"A2",X"05",X"B5",X"D7",X"95",X"CF",X"CA",
		X"D0",X"F9",X"86",X"DF",X"60",X"20",X"F4",X"DE",X"A2",X"06",X"B5",X"CF",X"95",X"D7",X"CA",X"D0",
		X"F9",X"86",X"DF",X"60",X"A5",X"D0",X"F0",X"FB",X"06",X"DF",X"90",X"F7",X"20",X"2A",X"DC",X"D0",
		X"F2",X"4C",X"F3",X"DB",X"20",X"A9",X"D2",X"46",X"D4",X"B0",X"04",X"A9",X"00",X"F0",X"15",X"A9",
		X"FF",X"30",X"11",X"A5",X"D0",X"F0",X"09",X"A5",X"D5",X"2A",X"A9",X"FF",X"B0",X"02",X"A9",X"01",
		X"60",X"20",X"13",X"DF",X"85",X"D1",X"A9",X"00",X"85",X"D2",X"A2",X"88",X"A5",X"D1",X"49",X"FF",
		X"2A",X"A9",X"00",X"85",X"D4",X"85",X"D3",X"86",X"D0",X"85",X"DF",X"85",X"D5",X"4C",X"8D",X"DB",
		X"85",X"D1",X"84",X"D2",X"A2",X"90",X"38",X"B0",X"E8",X"46",X"D5",X"60",X"85",X"93",X"84",X"94",
		X"A0",X"00",X"B1",X"93",X"C8",X"AA",X"F0",X"BB",X"B1",X"93",X"45",X"D5",X"30",X"B9",X"E4",X"D0",
		X"D0",X"21",X"B1",X"93",X"09",X"80",X"C5",X"D1",X"D0",X"19",X"C8",X"B1",X"93",X"C5",X"D2",X"D0",
		X"12",X"C8",X"B1",X"93",X"C5",X"D3",X"D0",X"0B",X"C8",X"A9",X"7F",X"C5",X"DF",X"B1",X"93",X"E5",
		X"D4",X"F0",X"28",X"A5",X"D5",X"90",X"02",X"49",X"FF",X"4C",X"19",X"DF",X"A5",X"D0",X"F0",X"4A",
		X"38",X"E9",X"A0",X"24",X"D5",X"10",X"09",X"AA",X"A9",X"FF",X"85",X"D7",X"20",X"08",X"DC",X"8A",
		X"A2",X"D0",X"C9",X"F9",X"10",X"06",X"20",X"54",X"DC",X"84",X"D7",X"60",X"A8",X"A5",X"D5",X"29",
		X"80",X"46",X"D1",X"05",X"D1",X"85",X"D1",X"20",X"6B",X"DC",X"84",X"D7",X"60",X"A5",X"D0",X"C9",
		X"A0",X"B0",X"20",X"20",X"8C",X"DF",X"84",X"DF",X"A5",X"D5",X"84",X"D5",X"49",X"80",X"2A",X"A9",
		X"A0",X"85",X"D0",X"A5",X"D4",X"85",X"24",X"4C",X"8D",X"DB",X"85",X"D1",X"85",X"D2",X"85",X"D3",
		X"85",X"D4",X"A8",X"60",X"4C",X"81",X"E9",X"A0",X"00",X"A2",X"0A",X"94",X"CC",X"CA",X"10",X"FB",
		X"90",X"13",X"C9",X"23",X"F0",X"EE",X"C9",X"2D",X"D0",X"04",X"86",X"D6",X"F0",X"04",X"C9",X"2B",
		X"D0",X"05",X"20",X"E2",X"00",X"90",X"5B",X"C9",X"2E",X"F0",X"2E",X"C9",X"45",X"D0",X"30",X"20",
		X"E2",X"00",X"90",X"17",X"C9",X"CD",X"F0",X"0E",X"C9",X"2D",X"F0",X"0A",X"C9",X"CC",X"F0",X"08",
		X"C9",X"2B",X"F0",X"04",X"D0",X"07",X"66",X"CF",X"20",X"E2",X"00",X"90",X"5C",X"24",X"CF",X"10",
		X"0E",X"A9",X"00",X"38",X"E5",X"CD",X"4C",X"41",X"E0",X"66",X"CE",X"24",X"CE",X"50",X"C3",X"A5",
		X"CD",X"38",X"E5",X"CC",X"85",X"CD",X"F0",X"12",X"10",X"09",X"20",X"C3",X"DD",X"E6",X"CD",X"D0",
		X"F9",X"F0",X"07",X"20",X"A7",X"DD",X"C6",X"CD",X"D0",X"F9",X"A5",X"D6",X"30",X"01",X"60",X"4C",
		X"71",X"E2",X"48",X"24",X"CE",X"10",X"02",X"E6",X"CC",X"20",X"A7",X"DD",X"68",X"38",X"E9",X"30",
		X"20",X"76",X"E0",X"4C",X"02",X"E0",X"48",X"20",X"E5",X"DE",X"68",X"20",X"24",X"DF",X"A5",X"DD",
		X"45",X"D5",X"85",X"DE",X"A6",X"D0",X"4C",X"25",X"DB",X"A5",X"CD",X"C9",X"0A",X"90",X"09",X"A9",
		X"64",X"24",X"CF",X"30",X"11",X"4C",X"39",X"DC",X"0A",X"0A",X"18",X"65",X"CD",X"0A",X"18",X"A0",
		X"00",X"71",X"E9",X"38",X"E9",X"30",X"85",X"CD",X"4C",X"28",X"E0",X"9B",X"3E",X"BC",X"1F",X"FD",
		X"9E",X"6E",X"6B",X"27",X"FD",X"9E",X"6E",X"6B",X"28",X"00",X"A9",X"AD",X"A0",X"C3",X"20",X"D2",
		X"E0",X"A5",X"A9",X"A6",X"A8",X"85",X"D1",X"86",X"D2",X"A2",X"90",X"38",X"20",X"31",X"DF",X"20",
		X"D5",X"E0",X"4C",X"B0",X"CC",X"A0",X"01",X"A9",X"20",X"24",X"D5",X"10",X"02",X"A9",X"2D",X"99",
		X"FF",X"00",X"85",X"D5",X"84",X"E0",X"C8",X"A9",X"30",X"A6",X"D0",X"D0",X"03",X"4C",X"F8",X"E1",
		X"A9",X"00",X"E0",X"80",X"F0",X"02",X"B0",X"09",X"A9",X"B5",X"A0",X"E0",X"20",X"ED",X"DC",X"A9",
		X"F7",X"85",X"CC",X"A9",X"B0",X"A0",X"E0",X"20",X"4C",X"DF",X"F0",X"1E",X"10",X"12",X"A9",X"AB",
		X"A0",X"E0",X"20",X"4C",X"DF",X"F0",X"02",X"10",X"0E",X"20",X"A7",X"DD",X"C6",X"CC",X"D0",X"EE",
		X"20",X"C3",X"DD",X"E6",X"CC",X"D0",X"DC",X"20",X"04",X"DB",X"20",X"8C",X"DF",X"A2",X"01",X"A5",
		X"CC",X"18",X"69",X"0A",X"30",X"09",X"C9",X"0B",X"B0",X"06",X"69",X"FF",X"AA",X"A9",X"02",X"38",
		X"E9",X"02",X"85",X"CD",X"86",X"CC",X"8A",X"F0",X"02",X"10",X"13",X"A4",X"E0",X"A9",X"2E",X"C8",
		X"99",X"FF",X"00",X"8A",X"F0",X"06",X"A9",X"30",X"C8",X"99",X"FF",X"00",X"84",X"E0",X"A0",X"00",
		X"A2",X"80",X"A5",X"D4",X"18",X"79",X"0D",X"E2",X"85",X"D4",X"A5",X"D3",X"79",X"0C",X"E2",X"85",
		X"D3",X"A5",X"D2",X"79",X"0B",X"E2",X"85",X"D2",X"A5",X"D1",X"79",X"0A",X"E2",X"85",X"D1",X"E8",
		X"B0",X"04",X"10",X"DE",X"30",X"02",X"30",X"DA",X"8A",X"90",X"04",X"49",X"FF",X"69",X"0A",X"69",
		X"2F",X"C8",X"C8",X"C8",X"C8",X"84",X"B6",X"A4",X"E0",X"C8",X"AA",X"29",X"7F",X"99",X"FF",X"00",
		X"C6",X"CC",X"D0",X"06",X"A9",X"2E",X"C8",X"99",X"FF",X"00",X"84",X"E0",X"A4",X"B6",X"8A",X"49",
		X"FF",X"29",X"80",X"AA",X"C0",X"24",X"D0",X"AA",X"A4",X"E0",X"B9",X"FF",X"00",X"88",X"C9",X"30",
		X"F0",X"F8",X"C9",X"2E",X"F0",X"01",X"C8",X"A9",X"2B",X"A6",X"CD",X"F0",X"2E",X"10",X"08",X"A9",
		X"00",X"38",X"E5",X"CD",X"AA",X"A9",X"2D",X"99",X"01",X"01",X"A9",X"45",X"99",X"00",X"01",X"8A",
		X"A2",X"2F",X"38",X"E8",X"E9",X"0A",X"B0",X"FB",X"69",X"3A",X"99",X"03",X"01",X"8A",X"99",X"02",
		X"01",X"A9",X"00",X"99",X"04",X"01",X"F0",X"08",X"99",X"FF",X"00",X"A9",X"00",X"99",X"00",X"01",
		X"A9",X"00",X"A0",X"01",X"60",X"80",X"00",X"00",X"00",X"00",X"FA",X"0A",X"1F",X"00",X"00",X"98",
		X"96",X"80",X"FF",X"F0",X"BD",X"C0",X"00",X"01",X"86",X"A0",X"FF",X"FF",X"D8",X"F0",X"00",X"00",
		X"03",X"E8",X"FF",X"FF",X"FF",X"9C",X"00",X"00",X"00",X"0A",X"FF",X"FF",X"FF",X"FF",X"20",X"E5",
		X"DE",X"A9",X"05",X"A0",X"E2",X"20",X"7B",X"DE",X"F0",X"70",X"A5",X"D8",X"D0",X"03",X"4C",X"B4",
		X"DB",X"A2",X"BD",X"A0",X"00",X"20",X"AD",X"DE",X"A5",X"DD",X"10",X"0F",X"20",X"BD",X"DF",X"A9",
		X"BD",X"A0",X"00",X"20",X"4C",X"DF",X"D0",X"03",X"98",X"A4",X"24",X"20",X"D7",X"DE",X"98",X"48",
		X"20",X"AF",X"DC",X"A9",X"BD",X"A0",X"00",X"20",X"ED",X"DC",X"20",X"AA",X"E2",X"68",X"4A",X"90",
		X"0A",X"A5",X"D0",X"F0",X"06",X"A5",X"D5",X"49",X"FF",X"85",X"D5",X"60",X"81",X"38",X"AA",X"3B",
		X"29",X"07",X"71",X"34",X"58",X"3E",X"56",X"74",X"16",X"7E",X"B3",X"1B",X"77",X"2F",X"EE",X"E3",
		X"85",X"7A",X"1D",X"84",X"1C",X"2A",X"7C",X"63",X"59",X"58",X"0A",X"7E",X"75",X"FD",X"E7",X"C6",
		X"80",X"31",X"72",X"18",X"10",X"81",X"00",X"00",X"00",X"00",X"A9",X"7C",X"A0",X"E2",X"20",X"ED",
		X"DC",X"A5",X"DF",X"69",X"50",X"90",X"03",X"20",X"FC",X"DE",X"85",X"C5",X"20",X"E8",X"DE",X"A5",
		X"D0",X"C9",X"88",X"90",X"03",X"20",X"99",X"DD",X"20",X"BD",X"DF",X"A5",X"24",X"18",X"69",X"81",
		X"F0",X"F3",X"38",X"E9",X"01",X"48",X"A2",X"05",X"B5",X"D8",X"B4",X"D0",X"95",X"D0",X"94",X"D8",
		X"CA",X"10",X"F5",X"A5",X"C5",X"85",X"DF",X"20",X"0E",X"DB",X"20",X"71",X"E2",X"A9",X"81",X"A0",
		X"E2",X"20",X"13",X"E3",X"A9",X"00",X"85",X"DE",X"68",X"20",X"7E",X"DD",X"60",X"85",X"E0",X"84",
		X"E1",X"20",X"A3",X"DE",X"A9",X"C6",X"20",X"ED",X"DC",X"20",X"17",X"E3",X"A9",X"C6",X"A0",X"00",
		X"4C",X"ED",X"DC",X"85",X"E0",X"84",X"E1",X"20",X"A0",X"DE",X"B1",X"E0",X"85",X"D6",X"A4",X"E0",
		X"C8",X"98",X"D0",X"02",X"E6",X"E1",X"85",X"E0",X"A4",X"E1",X"20",X"ED",X"DC",X"A5",X"E0",X"A4",
		X"E1",X"18",X"69",X"05",X"90",X"01",X"C8",X"85",X"E0",X"84",X"E1",X"20",X"22",X"DB",X"A9",X"CB",
		X"A0",X"00",X"C6",X"D6",X"D0",X"E4",X"60",X"98",X"35",X"44",X"7A",X"68",X"28",X"B1",X"46",X"20",
		X"13",X"DF",X"AA",X"30",X"18",X"A9",X"FA",X"A0",X"00",X"20",X"7B",X"DE",X"8A",X"F0",X"E7",X"A9",
		X"47",X"A0",X"E3",X"20",X"ED",X"DC",X"A9",X"4B",X"A0",X"E3",X"20",X"22",X"DB",X"A6",X"D4",X"A5",
		X"D1",X"85",X"D4",X"86",X"D1",X"A9",X"00",X"85",X"D5",X"A5",X"D0",X"85",X"DF",X"A9",X"80",X"85",
		X"D0",X"20",X"92",X"DB",X"A2",X"FA",X"A0",X"00",X"4C",X"AD",X"DE",X"A9",X"07",X"A0",X"E4",X"20",
		X"22",X"DB",X"20",X"E5",X"DE",X"A9",X"0C",X"A0",X"E4",X"A6",X"DD",X"20",X"CC",X"DD",X"20",X"E5",
		X"DE",X"20",X"BD",X"DF",X"A9",X"00",X"85",X"DE",X"20",X"0E",X"DB",X"A9",X"11",X"A0",X"E4",X"20",
		X"0B",X"DB",X"A5",X"D5",X"48",X"10",X"0D",X"20",X"04",X"DB",X"A5",X"D5",X"30",X"09",X"A5",X"2D",
		X"49",X"FF",X"85",X"2D",X"20",X"71",X"E2",X"A9",X"11",X"A0",X"E4",X"20",X"22",X"DB",X"68",X"10",
		X"03",X"20",X"71",X"E2",X"A9",X"16",X"A0",X"E4",X"4C",X"FD",X"E2",X"20",X"A3",X"DE",X"A9",X"00",
		X"85",X"2D",X"20",X"92",X"E3",X"A2",X"BD",X"A0",X"00",X"20",X"88",X"E3",X"A9",X"C6",X"A0",X"00",
		X"20",X"7B",X"DE",X"A9",X"00",X"85",X"D5",X"A5",X"2D",X"20",X"03",X"E4",X"A9",X"BD",X"A0",X"00",
		X"4C",X"E4",X"DD",X"48",X"4C",X"C4",X"E3",X"81",X"49",X"0F",X"DA",X"A2",X"83",X"49",X"0F",X"DA",
		X"A2",X"7F",X"00",X"00",X"00",X"00",X"05",X"84",X"E6",X"1A",X"2D",X"1B",X"86",X"28",X"07",X"FB",
		X"F8",X"87",X"99",X"68",X"89",X"01",X"87",X"23",X"35",X"DF",X"E1",X"86",X"A5",X"5D",X"E7",X"28",
		X"83",X"49",X"0F",X"DA",X"A2",X"A1",X"54",X"46",X"8F",X"13",X"8F",X"52",X"43",X"89",X"CD",X"A5",
		X"D5",X"48",X"10",X"03",X"20",X"71",X"E2",X"A5",X"D0",X"48",X"C9",X"81",X"90",X"07",X"A9",X"81",
		X"A0",X"DC",X"20",X"E4",X"DD",X"A9",X"6F",X"A0",X"E4",X"20",X"FD",X"E2",X"68",X"C9",X"81",X"90",
		X"07",X"A9",X"07",X"A0",X"E4",X"20",X"0B",X"DB",X"68",X"10",X"03",X"4C",X"71",X"E2",X"60",X"0B",
		X"76",X"B3",X"83",X"BD",X"D3",X"79",X"1E",X"F4",X"A6",X"F5",X"7B",X"83",X"FC",X"B0",X"10",X"7C",
		X"0C",X"1F",X"67",X"CA",X"7C",X"DE",X"53",X"CB",X"C1",X"7D",X"14",X"64",X"70",X"4C",X"7D",X"B7",
		X"EA",X"51",X"7A",X"7D",X"63",X"30",X"88",X"7E",X"7E",X"92",X"44",X"99",X"3A",X"7E",X"4C",X"CC",
		X"91",X"C7",X"7F",X"AA",X"AA",X"AA",X"13",X"81",X"00",X"00",X"00",X"00",X"20",X"35",X"E7",X"20",
		X"C9",X"E6",X"C9",X"24",X"D0",X"F9",X"8E",X"B1",X"02",X"A2",X"09",X"20",X"C9",X"E6",X"9D",X"A7",
		X"02",X"CA",X"D0",X"F7",X"20",X"C9",X"E6",X"F0",X"0A",X"E0",X"10",X"B0",X"F7",X"9D",X"93",X"02",
		X"E8",X"D0",X"F1",X"9D",X"93",X"02",X"20",X"94",X"E5",X"20",X"90",X"E7",X"8A",X"D0",X"CD",X"60",
		X"AD",X"A9",X"02",X"AC",X"AA",X"02",X"85",X"33",X"84",X"34",X"A0",X"00",X"20",X"C9",X"E6",X"AE",
		X"5B",X"02",X"D0",X"05",X"91",X"33",X"4C",X"05",X"E5",X"D1",X"33",X"F0",X"08",X"EE",X"5C",X"02",
		X"D0",X"03",X"EE",X"5D",X"02",X"20",X"6C",X"E5",X"90",X"E2",X"60",X"10",X"07",X"53",X"65",X"61",
		X"72",X"63",X"68",X"69",X"6E",X"67",X"20",X"2E",X"2E",X"00",X"10",X"07",X"4C",X"6F",X"61",X"64",
		X"69",X"6E",X"67",X"20",X"2E",X"2E",X"00",X"0A",X"0D",X"45",X"72",X"72",X"6F",X"72",X"73",X"20",
		X"66",X"6F",X"75",X"6E",X"64",X"0D",X"0A",X"00",X"10",X"07",X"46",X"6F",X"75",X"6E",X"64",X"20",
		X"2E",X"2E",X"00",X"10",X"07",X"56",X"65",X"72",X"69",X"66",X"79",X"69",X"6E",X"67",X"20",X"2E",
		X"2E",X"00",X"20",X"56",X"65",X"72",X"69",X"66",X"79",X"20",X"65",X"72",X"72",X"6F",X"72",X"73",
		X"20",X"64",X"65",X"74",X"65",X"63",X"74",X"65",X"64",X"0D",X"0A",X"00",X"A5",X"33",X"CD",X"AB",
		X"02",X"A5",X"34",X"ED",X"AC",X"02",X"E6",X"33",X"D0",X"02",X"E6",X"34",X"60",X"A9",X"0B",X"A0",
		X"E5",X"20",X"EA",X"E5",X"60",X"A9",X"45",X"A0",X"E6",X"20",X"EA",X"E5",X"A9",X"7F",X"A0",X"02",
		X"20",X"B6",X"E5",X"60",X"A9",X"38",X"A0",X"E5",X"4C",X"AB",X"E5",X"AD",X"5B",X"02",X"D0",X"07",
		X"A9",X"1A",X"A0",X"E5",X"4C",X"AB",X"E5",X"A9",X"43",X"A0",X"E5",X"20",X"EA",X"E5",X"A9",X"93",
		X"A0",X"02",X"20",X"B6",X"E5",X"60",X"20",X"65",X"F8",X"E8",X"A0",X"00",X"8C",X"5F",X"02",X"AD",
		X"AE",X"02",X"F0",X"13",X"C8",X"2C",X"AE",X"02",X"30",X"0D",X"C8",X"2C",X"AF",X"02",X"30",X"07",
		X"C8",X"2C",X"B0",X"02",X"30",X"01",X"C8",X"B9",X"E5",X"E5",X"8D",X"5E",X"02",X"A9",X"5E",X"A0",
		X"02",X"20",X"65",X"F8",X"60",X"42",X"43",X"53",X"49",X"52",X"20",X"F5",X"E5",X"A2",X"00",X"20",
		X"65",X"F8",X"E8",X"E8",X"60",X"48",X"AD",X"1F",X"02",X"D0",X"0A",X"A2",X"22",X"A9",X"10",X"9D",
		X"80",X"BB",X"CA",X"10",X"FA",X"68",X"60",X"20",X"5A",X"E7",X"A9",X"24",X"20",X"5E",X"E6",X"A2",
		X"09",X"BD",X"A7",X"02",X"20",X"5E",X"E6",X"CA",X"D0",X"F7",X"BD",X"7F",X"02",X"F0",X"06",X"20",
		X"5E",X"E6",X"E8",X"D0",X"F5",X"20",X"5E",X"E6",X"A2",X"00",X"CA",X"D0",X"FD",X"60",X"AD",X"A9",
		X"02",X"AC",X"AA",X"02",X"85",X"33",X"84",X"34",X"A0",X"00",X"B1",X"33",X"20",X"5E",X"E6",X"20",
		X"6C",X"E5",X"90",X"F6",X"60",X"10",X"07",X"53",X"61",X"76",X"69",X"6E",X"67",X"20",X"2E",X"2E",
		X"00",X"AD",X"B1",X"02",X"F0",X"07",X"A9",X"27",X"A0",X"E5",X"20",X"B0",X"CC",X"60",X"85",X"2F",
		X"8A",X"48",X"98",X"48",X"20",X"C0",X"E6",X"18",X"A0",X"09",X"A9",X"00",X"F0",X"06",X"46",X"2F",
		X"08",X"69",X"00",X"28",X"20",X"8B",X"E6",X"88",X"D0",X"F4",X"49",X"01",X"4A",X"A0",X"04",X"20",
		X"8B",X"E6",X"38",X"88",X"D0",X"F9",X"68",X"A8",X"68",X"AA",X"60",X"48",X"08",X"AD",X"4D",X"02",
		X"D0",X"0A",X"38",X"20",X"B2",X"E6",X"28",X"20",X"B2",X"E6",X"68",X"60",X"20",X"B2",X"E6",X"A2",
		X"0F",X"28",X"B0",X"02",X"A2",X"07",X"20",X"AB",X"E6",X"68",X"60",X"20",X"C0",X"E6",X"CA",X"D0",
		X"FA",X"60",X"A9",X"D0",X"A2",X"00",X"B0",X"02",X"0A",X"E8",X"8D",X"06",X"03",X"8E",X"07",X"03",
		X"AD",X"04",X"03",X"2C",X"0D",X"03",X"50",X"FB",X"60",X"98",X"48",X"8A",X"48",X"20",X"1C",X"E7",
		X"20",X"1C",X"E7",X"B0",X"FB",X"20",X"FF",X"E6",X"B0",X"16",X"A9",X"00",X"A0",X"08",X"20",X"FC",
		X"E6",X"08",X"66",X"2F",X"28",X"69",X"00",X"88",X"D0",X"F4",X"20",X"FC",X"E6",X"E9",X"00",X"4A",
		X"90",X"03",X"2E",X"B1",X"02",X"68",X"AA",X"68",X"A8",X"A5",X"2F",X"60",X"20",X"1C",X"E7",X"48",
		X"AD",X"4D",X"02",X"F0",X"15",X"20",X"1C",X"E7",X"A2",X"02",X"90",X"02",X"A2",X"06",X"A9",X"00",
		X"20",X"1C",X"E7",X"69",X"00",X"CA",X"D0",X"F8",X"C9",X"04",X"68",X"60",X"48",X"AD",X"00",X"03",
		X"AD",X"0D",X"03",X"29",X"10",X"F0",X"F9",X"AD",X"09",X"03",X"48",X"A9",X"FF",X"8D",X"09",X"03",
		X"68",X"C9",X"FE",X"68",X"60",X"20",X"FC",X"E6",X"66",X"2F",X"A9",X"16",X"C5",X"2F",X"D0",X"F5",
		X"AD",X"4D",X"02",X"F0",X"08",X"20",X"1C",X"E7",X"20",X"1C",X"E7",X"B0",X"FB",X"A2",X"03",X"20",
		X"C9",X"E6",X"C9",X"16",X"D0",X"DF",X"CA",X"D0",X"F6",X"60",X"A2",X"02",X"A0",X"03",X"A9",X"16",
		X"20",X"5E",X"E6",X"88",X"D0",X"F8",X"CA",X"D0",X"F5",X"60",X"20",X"1A",X"EE",X"A0",X"06",X"78",
		X"BE",X"82",X"E7",X"B9",X"89",X"E7",X"9D",X"00",X"03",X"88",X"10",X"F4",X"A9",X"40",X"8D",X"00",
		X"03",X"60",X"05",X"04",X"0B",X"02",X"0C",X"08",X"0E",X"00",X"D0",X"C0",X"FF",X"10",X"F4",X"7F",
		X"A0",X"00",X"A2",X"00",X"AD",X"7F",X"02",X"F0",X"15",X"B9",X"7F",X"02",X"D9",X"93",X"02",X"F0",
		X"01",X"E8",X"99",X"93",X"02",X"C8",X"C0",X"11",X"B0",X"04",X"48",X"68",X"D0",X"EB",X"60",X"4C",
		X"70",X"D0",X"A9",X"00",X"8D",X"4D",X"02",X"8D",X"AD",X"02",X"8D",X"AE",X"02",X"8D",X"5B",X"02",
		X"8D",X"5A",X"02",X"8D",X"5C",X"02",X"8D",X"5D",X"02",X"8D",X"B1",X"02",X"20",X"17",X"CF",X"24",
		X"28",X"10",X"DC",X"20",X"D0",X"D7",X"AA",X"A0",X"00",X"E8",X"CA",X"F0",X"0A",X"B1",X"91",X"99",
		X"7F",X"02",X"C8",X"C0",X"10",X"D0",X"F3",X"A9",X"00",X"99",X"7F",X"02",X"20",X"E8",X"00",X"F0",
		X"61",X"C9",X"2C",X"D0",X"BA",X"20",X"E2",X"00",X"F0",X"58",X"C9",X"2C",X"F0",X"F7",X"C9",X"C7",
		X"D0",X"05",X"8D",X"AD",X"02",X"B0",X"EE",X"C9",X"53",X"D0",X"05",X"8D",X"4D",X"02",X"B0",X"E5",
		X"C9",X"56",X"D0",X"05",X"8D",X"5B",X"02",X"B0",X"DC",X"C9",X"4A",X"D0",X"05",X"8D",X"5A",X"02",
		X"B0",X"D3",X"C9",X"41",X"F0",X"04",X"C9",X"45",X"D0",X"47",X"85",X"0E",X"20",X"E2",X"00",X"A2",
		X"80",X"8E",X"AE",X"02",X"20",X"53",X"E8",X"A5",X"33",X"A4",X"34",X"A6",X"0E",X"E0",X"41",X"D0",
		X"08",X"8D",X"A9",X"02",X"8C",X"AA",X"02",X"B0",X"A3",X"8D",X"AB",X"02",X"8C",X"AC",X"02",X"4C",
		X"EC",X"E7",X"60",X"20",X"03",X"CF",X"20",X"22",X"D9",X"18",X"60",X"08",X"20",X"B2",X"E7",X"AD",
		X"AD",X"02",X"0D",X"AE",X"02",X"D0",X"0A",X"AD",X"5A",X"02",X"F0",X"08",X"AD",X"5B",X"02",X"F0",
		X"03",X"4C",X"70",X"D0",X"20",X"6A",X"E7",X"20",X"7D",X"E5",X"20",X"AC",X"E4",X"2C",X"AE",X"02",
		X"70",X"F8",X"AD",X"5A",X"02",X"F0",X"2C",X"AD",X"AE",X"02",X"D0",X"EE",X"A5",X"9C",X"A4",X"9D",
		X"38",X"E9",X"02",X"B0",X"01",X"88",X"8D",X"A9",X"02",X"8C",X"AA",X"02",X"38",X"E5",X"9A",X"AA",
		X"98",X"E5",X"9B",X"A8",X"18",X"8A",X"6D",X"AB",X"02",X"8D",X"AB",X"02",X"98",X"6D",X"AC",X"02",
		X"8D",X"AC",X"02",X"20",X"9B",X"E5",X"20",X"E0",X"E4",X"20",X"3D",X"E9",X"28",X"AD",X"5B",X"02",
		X"F0",X"11",X"AE",X"5C",X"02",X"AD",X"5D",X"02",X"20",X"C5",X"E0",X"A9",X"52",X"A0",X"E5",X"20",
		X"B0",X"CC",X"60",X"20",X"51",X"E6",X"AD",X"AE",X"02",X"F0",X"0E",X"AD",X"AD",X"02",X"F0",X"08",
		X"AD",X"B1",X"02",X"EA",X"EA",X"6C",X"A9",X"02",X"60",X"AE",X"AB",X"02",X"AD",X"AC",X"02",X"86",
		X"9C",X"85",X"9D",X"20",X"5F",X"C5",X"AD",X"AD",X"02",X"F0",X"08",X"AD",X"B1",X"02",X"EA",X"EA",
		X"4C",X"08",X"C7",X"20",X"08",X"C7",X"4C",X"A8",X"C4",X"A5",X"9A",X"A4",X"9B",X"8D",X"A9",X"02",
		X"8C",X"AA",X"02",X"A5",X"9C",X"A4",X"9D",X"8D",X"AB",X"02",X"8C",X"AC",X"02",X"08",X"20",X"B2",
		X"E7",X"AD",X"5A",X"02",X"0D",X"5B",X"02",X"F0",X"03",X"4C",X"70",X"D0",X"20",X"6A",X"E7",X"20",
		X"85",X"E5",X"20",X"07",X"E6",X"20",X"2E",X"E6",X"20",X"3D",X"E9",X"28",X"60",X"20",X"F5",X"E5",
		X"20",X"AA",X"F9",X"4C",X"E0",X"ED",X"20",X"53",X"E8",X"6C",X"33",X"00",X"A2",X"00",X"86",X"0C",
		X"86",X"0D",X"F0",X"13",X"A2",X"03",X"0A",X"0A",X"0A",X"0A",X"0A",X"26",X"0C",X"26",X"0D",X"90",
		X"03",X"4C",X"39",X"DC",X"CA",X"10",X"F3",X"20",X"E2",X"00",X"C9",X"80",X"B0",X"0E",X"09",X"80",
		X"49",X"B0",X"C9",X"0A",X"90",X"DE",X"69",X"88",X"C9",X"FA",X"B0",X"D8",X"A5",X"0D",X"A4",X"0C",
		X"60",X"20",X"4C",X"E9",X"4C",X"40",X"DF",X"08",X"20",X"57",X"EA",X"A9",X"40",X"8D",X"AE",X"02",
		X"A5",X"28",X"8D",X"AF",X"02",X"A5",X"29",X"8D",X"B0",X"02",X"20",X"85",X"E5",X"20",X"07",X"E6",
		X"20",X"9E",X"EA",X"20",X"2E",X"E6",X"24",X"28",X"10",X"22",X"A0",X"00",X"B1",X"0C",X"F0",X"17",
		X"AA",X"A0",X"02",X"B1",X"0C",X"99",X"D0",X"00",X"88",X"D0",X"F8",X"E8",X"CA",X"F0",X"08",X"B1",
		X"D1",X"20",X"5E",X"E6",X"C8",X"D0",X"F5",X"20",X"42",X"EA",X"90",X"DE",X"20",X"3D",X"E9",X"28",
		X"60",X"20",X"50",X"D6",X"08",X"20",X"57",X"EA",X"20",X"7D",X"E5",X"20",X"AC",X"E4",X"2C",X"AE",
		X"02",X"50",X"F8",X"AD",X"AF",X"02",X"45",X"28",X"D0",X"F1",X"AD",X"B0",X"02",X"45",X"29",X"D0",
		X"EA",X"20",X"9B",X"E5",X"A0",X"02",X"B1",X"CE",X"CD",X"A9",X"02",X"C8",X"B1",X"CE",X"ED",X"AA",
		X"02",X"B0",X"06",X"20",X"3D",X"E9",X"4C",X"7C",X"C4",X"20",X"9E",X"EA",X"20",X"E0",X"E4",X"24",
		X"28",X"10",X"27",X"A0",X"00",X"B1",X"0C",X"F0",X"1C",X"20",X"AB",X"D5",X"A0",X"00",X"AA",X"E8",
		X"CA",X"F0",X"08",X"20",X"C9",X"E6",X"91",X"D1",X"C8",X"D0",X"F5",X"A0",X"02",X"B9",X"D0",X"00",
		X"91",X"0C",X"88",X"D0",X"F8",X"20",X"42",X"EA",X"90",X"D9",X"20",X"3D",X"E9",X"20",X"51",X"E6",
		X"28",X"60",X"18",X"A9",X"03",X"65",X"0C",X"85",X"0C",X"90",X"02",X"E6",X"0D",X"A8",X"A5",X"0D",
		X"CC",X"AB",X"02",X"ED",X"AC",X"02",X"60",X"A9",X"40",X"85",X"2B",X"20",X"88",X"D1",X"A9",X"00",
		X"85",X"2B",X"A0",X"03",X"B1",X"CE",X"8D",X"AA",X"02",X"88",X"B1",X"CE",X"8D",X"A9",X"02",X"D0",
		X"03",X"CE",X"AA",X"02",X"CE",X"A9",X"02",X"20",X"65",X"D0",X"A5",X"29",X"48",X"A5",X"28",X"48",
		X"20",X"B2",X"E7",X"68",X"85",X"28",X"68",X"85",X"29",X"AD",X"5B",X"02",X"0D",X"AD",X"02",X"0D",
		X"AE",X"02",X"0D",X"5A",X"02",X"F0",X"03",X"4C",X"70",X"D0",X"20",X"6A",X"E7",X"60",X"18",X"A5",
		X"CE",X"6D",X"A9",X"02",X"8D",X"AB",X"02",X"A5",X"CF",X"6D",X"AA",X"02",X"8D",X"AC",X"02",X"A0",
		X"04",X"B1",X"CE",X"20",X"88",X"D2",X"8D",X"A9",X"02",X"8C",X"AA",X"02",X"85",X"0C",X"84",X"0D",
		X"60",X"3F",X"FB",X"17",X"FC",X"CF",X"FB",X"C7",X"F0",X"FC",X"F0",X"0F",X"F1",X"7E",X"F3",X"1C",
		X"F1",X"67",X"F2",X"2C",X"F1",X"03",X"F2",X"0F",X"F2",X"03",X"04",X"04",X"03",X"03",X"03",X"02",
		X"01",X"03",X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",
		X"AD",X"C0",X"02",X"29",X"01",X"D0",X"05",X"A2",X"A3",X"4C",X"7E",X"C4",X"C0",X"4E",X"B0",X"03",
		X"4C",X"70",X"D0",X"C0",X"66",X"B0",X"F9",X"98",X"38",X"E9",X"4E",X"A8",X"B9",X"C2",X"EA",X"48",
		X"B9",X"C1",X"EA",X"48",X"98",X"4A",X"A8",X"B9",X"D9",X"EA",X"48",X"B9",X"E5",X"EA",X"8D",X"C3",
		X"02",X"A9",X"00",X"8D",X"F0",X"02",X"20",X"03",X"CF",X"AD",X"C3",X"02",X"D0",X"06",X"20",X"22",
		X"D9",X"4C",X"3B",X"EB",X"A5",X"D0",X"C9",X"90",X"20",X"2A",X"D9",X"AC",X"F0",X"02",X"A5",X"33",
		X"99",X"E1",X"02",X"A5",X"34",X"99",X"E2",X"02",X"C8",X"C8",X"8C",X"F0",X"02",X"68",X"A8",X"88",
		X"F0",X"08",X"98",X"48",X"20",X"65",X"D0",X"4C",X"26",X"EB",X"A9",X"00",X"8D",X"E0",X"02",X"68",
		X"AA",X"68",X"A8",X"A9",X"EB",X"48",X"A9",X"6D",X"48",X"98",X"48",X"8A",X"48",X"60",X"A9",X"01",
		X"2C",X"E0",X"02",X"F0",X"F8",X"4C",X"36",X"D3",X"AD",X"DF",X"02",X"10",X"0B",X"08",X"29",X"7F",
		X"48",X"A9",X"00",X"8D",X"DF",X"02",X"68",X"28",X"60",X"C4",X"9D",X"B0",X"02",X"38",X"60",X"D0",
		X"06",X"C5",X"9C",X"90",X"F9",X"F0",X"F7",X"20",X"B5",X"EB",X"90",X"F2",X"AA",X"AD",X"C0",X"02",
		X"29",X"02",X"08",X"8A",X"28",X"D0",X"E6",X"98",X"48",X"38",X"E9",X"1C",X"A8",X"8A",X"20",X"B5",
		X"EB",X"68",X"A8",X"8A",X"60",X"CC",X"C2",X"02",X"90",X"02",X"F0",X"01",X"60",X"CD",X"C1",X"02",
		X"60",X"AC",X"C2",X"02",X"AD",X"C1",X"02",X"D0",X"01",X"88",X"38",X"E9",X"01",X"60",X"20",X"03",
		X"CF",X"20",X"22",X"D9",X"A5",X"33",X"A4",X"34",X"20",X"89",X"EB",X"90",X"03",X"4C",X"7C",X"C4",
		X"85",X"A6",X"84",X"A7",X"4C",X"0F",X"C7",X"AD",X"60",X"02",X"D0",X"F1",X"AD",X"C0",X"02",X"48",
		X"29",X"01",X"F0",X"05",X"A2",X"A3",X"4C",X"7E",X"C4",X"68",X"29",X"FD",X"8D",X"C0",X"02",X"20",
		X"C1",X"EB",X"48",X"98",X"18",X"69",X"1C",X"A8",X"68",X"4C",X"E0",X"EB",X"20",X"C1",X"EB",X"20",
		X"89",X"EB",X"B0",X"C9",X"48",X"AD",X"C0",X"02",X"09",X"02",X"8D",X"C0",X"02",X"68",X"4C",X"E0",
		X"EB",X"AD",X"C0",X"02",X"A8",X"29",X"01",X"F0",X"09",X"98",X"29",X"FE",X"8D",X"C0",X"02",X"20",
		X"67",X"F9",X"60",X"AD",X"C0",X"02",X"48",X"29",X"02",X"F0",X"B9",X"68",X"09",X"01",X"8D",X"C0",
		X"02",X"20",X"20",X"F9",X"60",X"20",X"62",X"D0",X"20",X"17",X"CF",X"A5",X"34",X"48",X"A5",X"33",
		X"48",X"20",X"22",X"D9",X"A5",X"33",X"8D",X"E1",X"02",X"A5",X"34",X"8D",X"E2",X"02",X"68",X"85",
		X"33",X"68",X"85",X"34",X"20",X"65",X"D0",X"20",X"17",X"CF",X"A5",X"34",X"48",X"A5",X"33",X"48",
		X"20",X"22",X"D9",X"A5",X"34",X"8D",X"E4",X"02",X"A5",X"33",X"8D",X"E3",X"02",X"68",X"85",X"33",
		X"68",X"85",X"34",X"20",X"C8",X"F1",X"AC",X"E1",X"02",X"AD",X"E0",X"02",X"29",X"01",X"D0",X"09",
		X"AD",X"E2",X"02",X"20",X"99",X"D4",X"4C",X"5F",X"D0",X"4C",X"C2",X"D8",X"E6",X"E9",X"D0",X"02",
		X"E6",X"EA",X"AD",X"60",X"EA",X"C9",X"20",X"F0",X"F3",X"20",X"B9",X"EC",X"60",X"2C",X"60",X"EA",
		X"2C",X"60",X"EA",X"60",X"80",X"4F",X"C7",X"52",X"58",X"C9",X"C8",X"F0",X"0E",X"C9",X"27",X"F0",
		X"0A",X"C9",X"3A",X"B0",X"06",X"38",X"E9",X"30",X"38",X"E9",X"D0",X"60",X"D8",X"A2",X"FF",X"86",
		X"A9",X"9A",X"A9",X"CC",X"A0",X"EC",X"85",X"1B",X"84",X"1C",X"A9",X"4C",X"85",X"1A",X"85",X"C3",
		X"85",X"21",X"8D",X"FB",X"02",X"A9",X"36",X"A0",X"D3",X"85",X"22",X"84",X"23",X"8D",X"FC",X"02",
		X"8C",X"FD",X"02",X"8D",X"F5",X"02",X"8C",X"F6",X"02",X"A2",X"1C",X"BD",X"9B",X"EC",X"95",X"E1",
		X"CA",X"D0",X"F8",X"A9",X"03",X"85",X"C2",X"8A",X"85",X"D7",X"85",X"87",X"85",X"2F",X"48",X"85",
		X"2E",X"8D",X"F2",X"02",X"A2",X"88",X"86",X"85",X"A8",X"A9",X"02",X"8D",X"C0",X"02",X"A9",X"28",
		X"8D",X"57",X"02",X"A9",X"50",X"8D",X"56",X"02",X"A9",X"00",X"85",X"30",X"8D",X"58",X"02",X"8D",
		X"59",X"02",X"20",X"3E",X"C8",X"20",X"CE",X"CC",X"A9",X"96",X"A0",X"ED",X"20",X"B0",X"CC",X"20",
		X"F0",X"CB",X"A2",X"00",X"A0",X"05",X"86",X"9A",X"84",X"9B",X"A0",X"00",X"98",X"91",X"9A",X"E6",
		X"9A",X"D0",X"02",X"E6",X"9B",X"20",X"F0",X"C6",X"A5",X"9A",X"A4",X"9B",X"20",X"44",X"C4",X"20",
		X"F0",X"CB",X"A5",X"A6",X"38",X"E5",X"9A",X"AA",X"A5",X"A7",X"E5",X"9B",X"20",X"C5",X"E0",X"A9",
		X"88",X"A0",X"ED",X"20",X"B0",X"CC",X"A9",X"B0",X"A0",X"CC",X"85",X"1B",X"84",X"1C",X"A9",X"10",
		X"8D",X"F8",X"02",X"4C",X"A8",X"C4",X"00",X"00",X"20",X"42",X"59",X"54",X"45",X"53",X"20",X"46",
		X"52",X"45",X"45",X"0A",X"0D",X"00",X"4F",X"52",X"49",X"43",X"20",X"45",X"58",X"54",X"45",X"4E",
		X"44",X"45",X"44",X"20",X"42",X"41",X"53",X"49",X"43",X"20",X"56",X"31",X"2E",X"31",X"75",X"6B",
		X"0D",X"0A",X"31",X"39",X"38",X"33",X"20",X"54",X"41",X"4E",X"47",X"45",X"52",X"49",X"4E",X"45",
		X"0D",X"0A",X"00",X"00",X"A2",X"00",X"A0",X"00",X"C4",X"10",X"D0",X"04",X"E4",X"11",X"F0",X"0F",
		X"B1",X"0C",X"91",X"0E",X"C8",X"D0",X"F1",X"E6",X"0D",X"E6",X"0F",X"E8",X"4C",X"C8",X"ED",X"60",
		X"48",X"20",X"8C",X"EE",X"A9",X"00",X"A2",X"00",X"A0",X"03",X"20",X"AB",X"EE",X"A9",X"01",X"A0",
		X"19",X"20",X"AB",X"EE",X"A9",X"00",X"8D",X"71",X"02",X"AD",X"0B",X"03",X"29",X"7F",X"09",X"40",
		X"8D",X"0B",X"03",X"A9",X"C0",X"8D",X"0E",X"03",X"A9",X"10",X"8D",X"06",X"03",X"8D",X"04",X"03",
		X"A9",X"27",X"8D",X"07",X"03",X"8D",X"05",X"03",X"68",X"60",X"48",X"A9",X"40",X"8D",X"0E",X"03",
		X"68",X"60",X"48",X"AD",X"0D",X"03",X"29",X"40",X"F0",X"06",X"8D",X"0D",X"03",X"20",X"34",X"EE",
		X"68",X"4C",X"4A",X"02",X"48",X"8A",X"48",X"98",X"48",X"A0",X"00",X"B9",X"72",X"02",X"38",X"E9",
		X"01",X"99",X"72",X"02",X"C8",X"B9",X"72",X"02",X"E9",X"00",X"99",X"72",X"02",X"C8",X"C0",X"06",
		X"D0",X"E9",X"A9",X"00",X"20",X"9D",X"EE",X"C0",X"00",X"D0",X"10",X"A2",X"00",X"A0",X"03",X"20",
		X"AB",X"EE",X"20",X"95",X"F4",X"8A",X"10",X"03",X"8E",X"DF",X"02",X"A9",X"01",X"20",X"9D",X"EE",
		X"C0",X"00",X"D0",X"12",X"A2",X"00",X"A0",X"19",X"20",X"AB",X"EE",X"AD",X"71",X"02",X"49",X"01",
		X"8D",X"71",X"02",X"20",X"01",X"F8",X"68",X"A8",X"68",X"AA",X"68",X"60",X"48",X"98",X"48",X"A0",
		X"05",X"A9",X"00",X"99",X"72",X"02",X"88",X"10",X"FA",X"68",X"A8",X"68",X"60",X"48",X"0A",X"A8",
		X"78",X"B9",X"72",X"02",X"BE",X"73",X"02",X"58",X"A8",X"68",X"60",X"48",X"8A",X"48",X"98",X"48",
		X"BA",X"BD",X"03",X"01",X"0A",X"A8",X"68",X"48",X"78",X"99",X"72",X"02",X"BD",X"02",X"01",X"99",
		X"73",X"02",X"58",X"68",X"A8",X"68",X"AA",X"68",X"60",X"20",X"AB",X"EE",X"20",X"9D",X"EE",X"C0",
		X"00",X"D0",X"F9",X"E0",X"00",X"D0",X"F5",X"60",X"AD",X"13",X"02",X"8D",X"14",X"02",X"4E",X"12",
		X"02",X"6E",X"12",X"02",X"6E",X"12",X"02",X"60",X"48",X"98",X"48",X"20",X"DE",X"EE",X"20",X"49",
		X"F0",X"20",X"24",X"F0",X"68",X"A8",X"68",X"60",X"D8",X"20",X"D8",X"EE",X"2C",X"E2",X"02",X"10",
		X"0A",X"A9",X"FF",X"4D",X"E1",X"02",X"AA",X"E8",X"8E",X"E1",X"02",X"2C",X"E4",X"02",X"10",X"0A",
		X"A9",X"FF",X"4D",X"E3",X"02",X"AA",X"E8",X"8E",X"E3",X"02",X"AD",X"E1",X"02",X"CD",X"E3",X"02",
		X"90",X"0F",X"AE",X"E1",X"02",X"F0",X"09",X"AD",X"E3",X"02",X"20",X"40",X"EF",X"20",X"84",X"EF",
		X"60",X"AE",X"E3",X"02",X"F0",X"09",X"AD",X"E1",X"02",X"20",X"40",X"EF",X"20",X"5C",X"EF",X"60",
		X"85",X"0D",X"8E",X"00",X"02",X"A9",X"00",X"85",X"0C",X"8D",X"01",X"02",X"20",X"C8",X"EF",X"20",
		X"FA",X"EF",X"A9",X"00",X"85",X"0E",X"85",X"0F",X"8D",X"00",X"02",X"60",X"2C",X"E4",X"02",X"10",
		X"06",X"20",X"95",X"F0",X"4C",X"6A",X"EF",X"20",X"89",X"F0",X"20",X"AC",X"EF",X"F0",X"0E",X"2C",
		X"E2",X"02",X"10",X"06",X"20",X"B2",X"F0",X"4C",X"7D",X"EF",X"20",X"A1",X"F0",X"20",X"16",X"F0",
		X"CA",X"D0",X"D9",X"60",X"2C",X"E2",X"02",X"10",X"06",X"20",X"B2",X"F0",X"4C",X"92",X"EF",X"20",
		X"A1",X"F0",X"20",X"AC",X"EF",X"F0",X"0E",X"2C",X"E4",X"02",X"10",X"06",X"20",X"95",X"F0",X"4C",
		X"A5",X"EF",X"20",X"89",X"F0",X"20",X"16",X"F0",X"CA",X"D0",X"D9",X"60",X"D8",X"18",X"A5",X"0E",
		X"65",X"0C",X"85",X"0E",X"A5",X"0F",X"65",X"0D",X"85",X"0F",X"24",X"0E",X"10",X"03",X"18",X"69",
		X"01",X"CD",X"00",X"02",X"8D",X"00",X"02",X"60",X"48",X"8A",X"48",X"98",X"48",X"A9",X"00",X"85",
		X"0E",X"85",X"0F",X"A2",X"10",X"06",X"0C",X"26",X"0D",X"26",X"0E",X"26",X"0F",X"A5",X"0E",X"38",
		X"ED",X"00",X"02",X"A8",X"A5",X"0F",X"ED",X"01",X"02",X"90",X"06",X"E6",X"0C",X"84",X"0E",X"85",
		X"0F",X"CA",X"D0",X"E1",X"68",X"A8",X"68",X"AA",X"68",X"60",X"48",X"0E",X"00",X"02",X"2E",X"01",
		X"02",X"AD",X"00",X"02",X"38",X"E5",X"0E",X"AD",X"01",X"02",X"E5",X"0F",X"B0",X"06",X"E6",X"0C",
		X"D0",X"02",X"E6",X"0D",X"68",X"60",X"2C",X"14",X"02",X"18",X"10",X"04",X"20",X"24",X"F0",X"38",
		X"2E",X"14",X"02",X"60",X"A0",X"00",X"B1",X"10",X"29",X"40",X"F0",X"1C",X"AD",X"15",X"02",X"2C",
		X"12",X"02",X"30",X"0E",X"70",X"07",X"49",X"FF",X"31",X"10",X"91",X"10",X"60",X"11",X"10",X"91",
		X"10",X"60",X"70",X"04",X"51",X"10",X"91",X"10",X"60",X"D8",X"48",X"98",X"48",X"20",X"31",X"F7",
		X"18",X"69",X"00",X"85",X"10",X"98",X"69",X"A0",X"85",X"11",X"A9",X"00",X"85",X"0D",X"8D",X"01",
		X"02",X"86",X"0C",X"A9",X"06",X"8D",X"00",X"02",X"20",X"C8",X"EF",X"18",X"A5",X"0C",X"65",X"10",
		X"85",X"10",X"A9",X"00",X"65",X"11",X"85",X"11",X"A9",X"20",X"A4",X"0E",X"F0",X"04",X"4A",X"88",
		X"90",X"FA",X"8D",X"15",X"02",X"68",X"A8",X"68",X"60",X"18",X"A5",X"10",X"69",X"28",X"85",X"10",
		X"90",X"02",X"E6",X"11",X"60",X"38",X"A5",X"10",X"E9",X"28",X"85",X"10",X"B0",X"02",X"C6",X"11",
		X"60",X"4E",X"15",X"02",X"90",X"0B",X"A9",X"20",X"8D",X"15",X"02",X"E6",X"10",X"D0",X"02",X"E6",
		X"11",X"60",X"0E",X"15",X"02",X"2C",X"15",X"02",X"50",X"0D",X"A9",X"01",X"8D",X"15",X"02",X"A5",
		X"10",X"D0",X"02",X"C6",X"11",X"C6",X"10",X"60",X"A9",X"04",X"A2",X"E5",X"20",X"F8",X"F2",X"B0",
		X"28",X"AD",X"E5",X"02",X"8D",X"12",X"02",X"A9",X"F0",X"A2",X"E1",X"20",X"F8",X"F2",X"B0",X"19",
		X"A9",X"C8",X"A2",X"E3",X"20",X"F8",X"F2",X"B0",X"10",X"AE",X"E1",X"02",X"8E",X"19",X"02",X"AC",
		X"E3",X"02",X"8C",X"1A",X"02",X"20",X"E8",X"EE",X"60",X"EE",X"E0",X"02",X"60",X"20",X"0A",X"F3",
		X"B0",X"0A",X"AE",X"19",X"02",X"AC",X"1A",X"02",X"20",X"E8",X"EE",X"60",X"EE",X"E0",X"02",X"60",
		X"20",X"0A",X"F3",X"B0",X"04",X"20",X"F8",X"EE",X"60",X"EE",X"E0",X"02",X"60",X"AE",X"E2",X"02",
		X"D0",X"07",X"AE",X"E1",X"02",X"8E",X"13",X"02",X"60",X"EE",X"E0",X"02",X"60",X"AE",X"E2",X"02",
		X"D0",X"3B",X"AE",X"E1",X"02",X"E0",X"20",X"90",X"34",X"E0",X"80",X"B0",X"30",X"A9",X"02",X"A2",
		X"E3",X"20",X"F8",X"F2",X"B0",X"27",X"A9",X"04",X"A2",X"E5",X"20",X"F8",X"F2",X"B0",X"1E",X"AD",
		X"19",X"02",X"C9",X"EB",X"B0",X"17",X"AD",X"1A",X"02",X"C9",X"C1",X"B0",X"10",X"20",X"71",X"F1",
		X"20",X"9B",X"F1",X"AE",X"19",X"02",X"AC",X"1A",X"02",X"20",X"49",X"F0",X"60",X"EE",X"E0",X"02",
		X"60",X"D8",X"AD",X"E5",X"02",X"8D",X"12",X"02",X"20",X"DE",X"EE",X"AD",X"E1",X"02",X"85",X"0C",
		X"A9",X"00",X"85",X"0D",X"A2",X"03",X"06",X"0C",X"26",X"0D",X"CA",X"D0",X"F9",X"AD",X"E3",X"02",
		X"0A",X"0A",X"18",X"69",X"98",X"18",X"65",X"0D",X"85",X"0D",X"60",X"D8",X"A0",X"00",X"84",X"0F",
		X"B1",X"0C",X"85",X"0E",X"20",X"5D",X"F3",X"26",X"0E",X"26",X"0E",X"A2",X"06",X"26",X"0E",X"90",
		X"03",X"20",X"24",X"F0",X"20",X"A1",X"F0",X"CA",X"D0",X"F3",X"20",X"6E",X"F3",X"20",X"89",X"F0",
		X"A4",X"0F",X"C8",X"C0",X"08",X"D0",X"D7",X"60",X"A9",X"F0",X"A2",X"E1",X"20",X"F8",X"F2",X"B0",
		X"2F",X"A9",X"C8",X"A2",X"E3",X"20",X"F8",X"F2",X"B0",X"26",X"AE",X"E1",X"02",X"8E",X"19",X"02",
		X"AC",X"E3",X"02",X"8C",X"1A",X"02",X"20",X"49",X"F0",X"A0",X"00",X"B1",X"10",X"2D",X"15",X"02",
		X"F0",X"05",X"A9",X"FF",X"4C",X"F9",X"F1",X"A9",X"00",X"8D",X"E1",X"02",X"8D",X"E2",X"02",X"60",
		X"EE",X"E0",X"02",X"60",X"A9",X"10",X"85",X"0C",X"A9",X"00",X"85",X"0D",X"20",X"1C",X"F2",X"60",
		X"A9",X"00",X"85",X"0C",X"A9",X"01",X"85",X"0D",X"20",X"1C",X"F2",X"60",X"A9",X"08",X"A2",X"E1",
		X"20",X"F8",X"F2",X"B0",X"3F",X"20",X"5D",X"F3",X"AD",X"E1",X"02",X"05",X"0C",X"8D",X"02",X"02",
		X"AE",X"1F",X"02",X"D0",X"12",X"A6",X"0D",X"9D",X"6B",X"02",X"A9",X"A8",X"18",X"65",X"0D",X"AA",
		X"A0",X"BB",X"A9",X"1B",X"4C",X"51",X"F2",X"A9",X"00",X"18",X"65",X"0D",X"AA",X"A0",X"A0",X"A9",
		X"C8",X"8D",X"00",X"02",X"86",X"10",X"84",X"11",X"A9",X"01",X"8D",X"01",X"02",X"20",X"CD",X"F2",
		X"20",X"6E",X"F3",X"60",X"EE",X"E0",X"02",X"60",X"D8",X"AD",X"E3",X"02",X"8D",X"01",X"02",X"F0",
		X"58",X"A0",X"00",X"AD",X"19",X"02",X"38",X"E9",X"06",X"90",X"04",X"C8",X"4C",X"76",X"F2",X"98",
		X"18",X"6D",X"E3",X"02",X"A8",X"AD",X"E4",X"02",X"69",X"00",X"D0",X"3D",X"C0",X"29",X"B0",X"39",
		X"AD",X"E6",X"02",X"D0",X"34",X"AD",X"E1",X"02",X"8D",X"00",X"02",X"F0",X"2C",X"18",X"6D",X"1A",
		X"02",X"A8",X"AD",X"E2",X"02",X"69",X"00",X"D0",X"20",X"C0",X"C9",X"B0",X"1C",X"C0",X"C8",X"D0",
		X"02",X"A0",X"00",X"8C",X"1A",X"02",X"AD",X"E5",X"02",X"8D",X"02",X"02",X"20",X"CD",X"F2",X"AC",
		X"1A",X"02",X"AE",X"19",X"02",X"20",X"49",X"F0",X"60",X"EE",X"E0",X"02",X"60",X"D8",X"AD",X"02",
		X"02",X"A0",X"00",X"91",X"10",X"C8",X"CC",X"01",X"02",X"D0",X"F8",X"20",X"89",X"F0",X"CE",X"00",
		X"02",X"D0",X"EB",X"60",X"8D",X"04",X"02",X"BD",X"01",X"02",X"D0",X"0A",X"BD",X"00",X"02",X"F0",
		X"05",X"CD",X"04",X"02",X"90",X"01",X"38",X"60",X"8D",X"04",X"02",X"BD",X"01",X"02",X"D0",X"08",
		X"BD",X"00",X"02",X"CD",X"04",X"02",X"90",X"01",X"38",X"60",X"A9",X"04",X"A2",X"E5",X"20",X"F8",
		X"F2",X"B0",X"49",X"18",X"AD",X"E1",X"02",X"6D",X"19",X"02",X"8D",X"00",X"02",X"AD",X"E2",X"02",
		X"69",X"00",X"8D",X"01",X"02",X"A2",X"00",X"A9",X"F0",X"20",X"F8",X"F2",X"B0",X"2E",X"18",X"AD",
		X"E3",X"02",X"6D",X"1A",X"02",X"8D",X"02",X"02",X"AD",X"E4",X"02",X"69",X"00",X"8D",X"03",X"02",
		X"A2",X"02",X"A9",X"C8",X"20",X"F8",X"F2",X"B0",X"13",X"AD",X"E5",X"02",X"8D",X"12",X"02",X"AD",
		X"00",X"02",X"8D",X"19",X"02",X"AD",X"02",X"02",X"8D",X"1A",X"02",X"18",X"60",X"A5",X"10",X"8D",
		X"16",X"02",X"A5",X"11",X"8D",X"17",X"02",X"AD",X"15",X"02",X"8D",X"18",X"02",X"60",X"AD",X"16",
		X"02",X"85",X"10",X"AD",X"17",X"02",X"85",X"11",X"AD",X"18",X"02",X"8D",X"15",X"02",X"60",X"D8",
		X"AD",X"E2",X"02",X"D0",X"3D",X"AD",X"E1",X"02",X"F0",X"38",X"AD",X"19",X"02",X"CD",X"E1",X"02",
		X"90",X"30",X"18",X"6D",X"E1",X"02",X"C9",X"F0",X"B0",X"28",X"AD",X"1A",X"02",X"CD",X"E1",X"02",
		X"90",X"20",X"18",X"6D",X"E1",X"02",X"C9",X"C8",X"B0",X"18",X"A2",X"E3",X"A9",X"04",X"20",X"F8",
		X"F2",X"B0",X"0F",X"AD",X"E3",X"02",X"8D",X"12",X"02",X"20",X"D8",X"EE",X"20",X"C6",X"F3",X"4C",
		X"C5",X"F3",X"EE",X"E0",X"02",X"60",X"20",X"5D",X"F3",X"AD",X"1A",X"02",X"38",X"ED",X"E1",X"02",
		X"A8",X"AE",X"19",X"02",X"20",X"49",X"F0",X"AD",X"E1",X"02",X"85",X"0F",X"20",X"85",X"F4",X"A9",
		X"80",X"8D",X"1B",X"02",X"8D",X"1D",X"02",X"A9",X"00",X"8D",X"1C",X"02",X"AD",X"E1",X"02",X"8D",
		X"1E",X"02",X"A9",X"00",X"85",X"0F",X"20",X"14",X"F4",X"20",X"44",X"F4",X"A5",X"0F",X"F0",X"03",
		X"20",X"16",X"F0",X"AD",X"1C",X"02",X"D0",X"EA",X"AD",X"1E",X"02",X"CD",X"E1",X"02",X"D0",X"E2",
		X"20",X"6E",X"F3",X"60",X"AD",X"1D",X"02",X"AE",X"1E",X"02",X"20",X"74",X"F4",X"A5",X"0C",X"18",
		X"6D",X"1B",X"02",X"8D",X"1B",X"02",X"AD",X"1C",X"02",X"85",X"0C",X"65",X"0D",X"8D",X"1C",X"02",
		X"C5",X"0C",X"F0",X"0F",X"B0",X"06",X"20",X"A1",X"F0",X"4C",X"3F",X"F4",X"20",X"B2",X"F0",X"A9",
		X"01",X"85",X"0F",X"60",X"AD",X"1B",X"02",X"AE",X"1C",X"02",X"20",X"74",X"F4",X"38",X"AD",X"1D",
		X"02",X"E5",X"0C",X"8D",X"1D",X"02",X"AD",X"1E",X"02",X"85",X"0C",X"E5",X"0D",X"8D",X"1E",X"02",
		X"C5",X"0C",X"F0",X"0F",X"B0",X"06",X"20",X"89",X"F0",X"4C",X"6F",X"F4",X"20",X"95",X"F0",X"A9",
		X"01",X"85",X"0F",X"60",X"85",X"0C",X"86",X"0D",X"A6",X"0E",X"A5",X"0D",X"2A",X"66",X"0D",X"66",
		X"0C",X"CA",X"D0",X"F6",X"60",X"E6",X"0F",X"A9",X"00",X"85",X"0E",X"A9",X"01",X"0A",X"E6",X"0E",
		X"C5",X"0F",X"90",X"F9",X"60",X"48",X"08",X"98",X"48",X"D8",X"AD",X"08",X"02",X"10",X"1E",X"29",
		X"87",X"8D",X"10",X"02",X"AE",X"0A",X"02",X"20",X"61",X"F5",X"CD",X"10",X"02",X"D0",X"0E",X"CE",
		X"0E",X"02",X"D0",X"33",X"AD",X"4F",X"02",X"8D",X"0E",X"02",X"4C",X"C6",X"F4",X"AD",X"4E",X"02",
		X"8D",X"0E",X"02",X"20",X"23",X"F5",X"20",X"EF",X"F4",X"AA",X"10",X"1D",X"48",X"AD",X"6A",X"02",
		X"29",X"08",X"D0",X"0F",X"68",X"48",X"C9",X"A0",X"90",X"06",X"20",X"14",X"FB",X"4C",X"E3",X"F4",
		X"20",X"2A",X"FB",X"68",X"4C",X"E9",X"F4",X"A9",X"00",X"AA",X"68",X"A8",X"28",X"68",X"60",X"AD",
		X"09",X"02",X"A8",X"A9",X"00",X"C0",X"A4",X"F0",X"04",X"C0",X"A7",X"D0",X"03",X"18",X"69",X"40",
		X"18",X"6D",X"08",X"02",X"10",X"1C",X"29",X"7F",X"AA",X"BD",X"78",X"FF",X"2D",X"0C",X"02",X"10",
		X"03",X"38",X"E9",X"20",X"29",X"7F",X"C0",X"A2",X"D0",X"06",X"C9",X"40",X"30",X"02",X"29",X"1F",
		X"09",X"80",X"60",X"A9",X"38",X"8D",X"0D",X"02",X"8D",X"08",X"02",X"8D",X"09",X"02",X"A9",X"7F",
		X"48",X"68",X"48",X"AA",X"A9",X"07",X"20",X"61",X"F5",X"0D",X"0D",X"02",X"10",X"12",X"A2",X"00",
		X"A0",X"20",X"CC",X"0D",X"02",X"D0",X"01",X"E8",X"9D",X"08",X"02",X"68",X"48",X"9D",X"0A",X"02",
		X"38",X"68",X"6A",X"48",X"38",X"AD",X"0D",X"02",X"E9",X"08",X"8D",X"0D",X"02",X"10",X"D2",X"68",
		X"60",X"48",X"A9",X"0E",X"20",X"90",X"F5",X"68",X"29",X"07",X"AA",X"8D",X"11",X"02",X"09",X"B8",
		X"8D",X"00",X"03",X"A0",X"04",X"88",X"D0",X"FD",X"AD",X"00",X"03",X"29",X"08",X"D0",X"0D",X"CA",
		X"8A",X"29",X"07",X"AA",X"CD",X"11",X"02",X"D0",X"E5",X"A9",X"00",X"60",X"8A",X"09",X"80",X"60",
		X"08",X"78",X"8D",X"0F",X"03",X"A8",X"8A",X"C0",X"07",X"D0",X"02",X"09",X"40",X"48",X"AD",X"0C",
		X"03",X"09",X"EE",X"8D",X"0C",X"03",X"29",X"11",X"09",X"CC",X"8D",X"0C",X"03",X"AA",X"68",X"8D",
		X"0F",X"03",X"8A",X"09",X"EC",X"8D",X"0C",X"03",X"29",X"11",X"09",X"CC",X"8D",X"0C",X"03",X"28",
		X"60",X"08",X"78",X"8D",X"01",X"03",X"AD",X"00",X"03",X"29",X"EF",X"8D",X"00",X"03",X"AD",X"00",
		X"03",X"09",X"10",X"8D",X"00",X"03",X"28",X"AD",X"0D",X"03",X"29",X"02",X"F0",X"F9",X"AD",X"0D",
		X"03",X"60",X"CF",X"CF",X"CF",X"CF",X"A3",X"CF",X"A6",X"CC",X"00",X"27",X"34",X"0F",X"66",X"99",
		X"60",X"CF",X"A7",X"B3",X"CF",X"A8",X"BE",X"CF",X"CF",X"CF",X"CF",X"CF",X"A5",X"A5",X"CF",X"A4",
		X"84",X"CF",X"29",X"1F",X"AA",X"BD",X"E2",X"F5",X"18",X"69",X"2F",X"8D",X"61",X"02",X"A9",X"00",
		X"69",X"F6",X"8D",X"62",X"02",X"AD",X"6A",X"02",X"48",X"29",X"FE",X"8D",X"6A",X"02",X"68",X"29",
		X"01",X"8D",X"51",X"02",X"A9",X"00",X"20",X"01",X"F8",X"38",X"A9",X"00",X"6C",X"61",X"02",X"CE",
		X"69",X"02",X"30",X"05",X"20",X"D7",X"F7",X"D0",X"40",X"A9",X"27",X"8D",X"69",X"02",X"AD",X"68",
		X"02",X"C9",X"01",X"F0",X"34",X"CE",X"68",X"02",X"38",X"A5",X"12",X"E9",X"28",X"85",X"12",X"B0",
		X"02",X"C6",X"13",X"4C",X"FE",X"F6",X"EE",X"69",X"02",X"A2",X"27",X"EC",X"69",X"02",X"10",X"19",
		X"20",X"0D",X"F7",X"AD",X"68",X"02",X"CD",X"7E",X"02",X"F0",X"11",X"EE",X"68",X"02",X"18",X"A5",
		X"12",X"69",X"28",X"85",X"12",X"90",X"02",X"E6",X"13",X"4C",X"FE",X"F6",X"20",X"5D",X"F3",X"A2",
		X"06",X"BD",X"77",X"02",X"95",X"0B",X"CA",X"D0",X"F8",X"20",X"C4",X"ED",X"20",X"6E",X"F3",X"20",
		X"1A",X"F7",X"4C",X"FE",X"F6",X"AE",X"7E",X"02",X"AD",X"7A",X"02",X"85",X"12",X"AD",X"7B",X"02",
		X"85",X"13",X"20",X"1A",X"F7",X"18",X"A5",X"12",X"69",X"28",X"85",X"12",X"90",X"02",X"E6",X"13",
		X"CA",X"D0",X"EF",X"20",X"0D",X"F7",X"A9",X"01",X"8D",X"68",X"02",X"AD",X"7A",X"02",X"85",X"12",
		X"AD",X"7B",X"02",X"85",X"13",X"4C",X"FE",X"F6",X"20",X"0D",X"F7",X"8E",X"53",X"02",X"4C",X"FE",
		X"F6",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"4D",X"6A",X"02",X"8D",X"6A",X"02",X"4C",
		X"FE",X"F6",X"AD",X"51",X"02",X"49",X"01",X"8D",X"51",X"02",X"4C",X"FE",X"F6",X"AD",X"0C",X"02",
		X"49",X"80",X"8D",X"0C",X"02",X"20",X"5A",X"F7",X"4C",X"FE",X"F6",X"20",X"9F",X"FA",X"AD",X"6A",
		X"02",X"0D",X"51",X"02",X"8D",X"6A",X"02",X"A9",X"01",X"20",X"01",X"F8",X"60",X"A2",X"00",X"20",
		X"DE",X"F7",X"D0",X"02",X"E8",X"E8",X"8E",X"69",X"02",X"60",X"A0",X"27",X"A9",X"20",X"91",X"12",
		X"88",X"10",X"FB",X"A0",X"00",X"AD",X"6B",X"02",X"91",X"12",X"AD",X"6C",X"02",X"C8",X"91",X"12",
		X"60",X"A0",X"00",X"8C",X"63",X"02",X"8D",X"64",X"02",X"0A",X"2E",X"63",X"02",X"0A",X"2E",X"63",
		X"02",X"18",X"6D",X"64",X"02",X"90",X"03",X"EE",X"63",X"02",X"0A",X"2E",X"63",X"02",X"0A",X"2E",
		X"63",X"02",X"0A",X"2E",X"63",X"02",X"AC",X"63",X"02",X"60",X"AD",X"0C",X"02",X"10",X"07",X"A9",
		X"70",X"A0",X"F7",X"4C",X"6A",X"F7",X"A9",X"76",X"A0",X"F7",X"A2",X"23",X"20",X"65",X"F8",X"60",
		X"07",X"43",X"41",X"50",X"53",X"00",X"07",X"20",X"20",X"20",X"20",X"00",X"48",X"08",X"98",X"48",
		X"8A",X"48",X"D8",X"E0",X"13",X"F0",X"46",X"E0",X"14",X"F0",X"42",X"E0",X"06",X"F0",X"3E",X"AD",
		X"6A",X"02",X"29",X"02",X"F0",X"3A",X"8A",X"C9",X"20",X"90",X"32",X"AD",X"6A",X"02",X"29",X"10",
		X"F0",X"13",X"8A",X"38",X"E9",X"40",X"30",X"09",X"29",X"1F",X"20",X"E4",X"F7",X"A9",X"1B",X"D0",
		X"1C",X"A9",X"20",X"10",X"F5",X"E0",X"7F",X"F0",X"08",X"68",X"48",X"20",X"E4",X"F7",X"4C",X"D0",
		X"F7",X"A9",X"08",X"20",X"02",X"F6",X"A9",X"20",X"20",X"E4",X"F7",X"A9",X"08",X"20",X"02",X"F6",
		X"68",X"AA",X"68",X"A8",X"28",X"68",X"60",X"AD",X"69",X"02",X"29",X"FE",X"D0",X"05",X"AD",X"6A",
		X"02",X"29",X"20",X"60",X"48",X"AC",X"69",X"02",X"91",X"12",X"2C",X"6A",X"02",X"50",X"0B",X"AD",
		X"69",X"02",X"18",X"69",X"28",X"A8",X"68",X"48",X"91",X"12",X"A9",X"09",X"20",X"02",X"F6",X"68",
		X"60",X"2D",X"6A",X"02",X"4A",X"6A",X"8D",X"65",X"02",X"AC",X"69",X"02",X"B1",X"12",X"29",X"7F",
		X"0D",X"65",X"02",X"91",X"12",X"60",X"A9",X"00",X"85",X"0C",X"A9",X"B9",X"85",X"0D",X"A9",X"00",
		X"20",X"2D",X"F8",X"A0",X"BA",X"84",X"0D",X"A9",X"20",X"20",X"2D",X"F8",X"60",X"A0",X"00",X"48",
		X"20",X"54",X"F8",X"91",X"0C",X"C8",X"68",X"48",X"20",X"52",X"F8",X"68",X"48",X"20",X"50",X"F8",
		X"91",X"0C",X"C8",X"C0",X"00",X"F0",X"07",X"68",X"18",X"69",X"01",X"4C",X"2F",X"F8",X"68",X"60",
		X"4A",X"4A",X"4A",X"4A",X"29",X"03",X"AA",X"BD",X"61",X"F8",X"91",X"0C",X"C8",X"91",X"0C",X"C8",
		X"60",X"00",X"38",X"07",X"3F",X"85",X"0C",X"84",X"0D",X"AD",X"1F",X"02",X"D0",X"0D",X"A0",X"00",
		X"B1",X"0C",X"F0",X"07",X"9D",X"80",X"BB",X"E8",X"C8",X"D0",X"F5",X"60",X"4C",X"7C",X"F7",X"4C",
		X"78",X"EB",X"4C",X"C1",X"F5",X"4C",X"65",X"F8",X"4C",X"22",X"EE",X"4C",X"B2",X"F8",X"40",X"A2",
		X"FF",X"9A",X"58",X"D8",X"A2",X"12",X"BD",X"7C",X"F8",X"9D",X"38",X"02",X"CA",X"10",X"F7",X"A9",
		X"20",X"8D",X"4E",X"02",X"A9",X"04",X"8D",X"4F",X"02",X"20",X"14",X"FA",X"20",X"B8",X"F8",X"4C",
		X"CC",X"EC",X"20",X"B8",X"F8",X"4C",X"71",X"C4",X"20",X"AA",X"F9",X"A9",X"07",X"A2",X"40",X"20",
		X"90",X"F5",X"20",X"E0",X"ED",X"20",X"0E",X"F9",X"A9",X"FF",X"8D",X"0C",X"02",X"20",X"C9",X"F9",
		X"A2",X"05",X"20",X"82",X"F9",X"20",X"16",X"F8",X"20",X"5A",X"F7",X"60",X"48",X"8A",X"48",X"A9",
		X"01",X"8D",X"1F",X"02",X"A9",X"BF",X"8D",X"7B",X"02",X"8D",X"79",X"02",X"A9",X"68",X"8D",X"7A",
		X"02",X"A9",X"90",X"8D",X"78",X"02",X"A9",X"03",X"8D",X"7E",X"02",X"A9",X"00",X"8D",X"7D",X"02",
		X"A9",X"50",X"8D",X"7C",X"02",X"A2",X"0C",X"20",X"38",X"02",X"68",X"AA",X"68",X"60",X"48",X"A9",
		X"03",X"8D",X"6A",X"02",X"A9",X"00",X"8D",X"6C",X"02",X"A9",X"17",X"8D",X"6B",X"02",X"68",X"60",
		X"48",X"AD",X"1F",X"02",X"D0",X"05",X"A2",X"0B",X"20",X"82",X"F9",X"A9",X"FE",X"2D",X"6A",X"02",
		X"8D",X"6A",X"02",X"A9",X"1E",X"8D",X"DF",X"BF",X"A9",X"40",X"8D",X"00",X"A0",X"A2",X"17",X"20",
		X"82",X"F9",X"A9",X"00",X"8D",X"19",X"02",X"8D",X"1A",X"02",X"85",X"10",X"A9",X"A0",X"85",X"11",
		X"A9",X"20",X"8D",X"15",X"02",X"A9",X"FF",X"8D",X"13",X"02",X"20",X"DC",X"F8",X"A9",X"01",X"0D",
		X"6A",X"02",X"8D",X"6A",X"02",X"68",X"60",X"48",X"A9",X"FE",X"2D",X"6A",X"02",X"8D",X"6A",X"02",
		X"A2",X"11",X"20",X"82",X"F9",X"20",X"C9",X"F9",X"A9",X"01",X"0D",X"6A",X"02",X"8D",X"6A",X"02",
		X"68",X"60",X"A0",X"06",X"BD",X"92",X"F9",X"99",X"0B",X"00",X"CA",X"88",X"D0",X"F6",X"20",X"C4",
		X"ED",X"60",X"78",X"FC",X"00",X"B5",X"00",X"03",X"00",X"B4",X"00",X"98",X"80",X"07",X"00",X"98",
		X"00",X"B4",X"80",X"07",X"00",X"A0",X"01",X"A0",X"3F",X"1F",X"A9",X"FF",X"8D",X"03",X"03",X"A9",
		X"F7",X"8D",X"02",X"03",X"A9",X"B7",X"8D",X"00",X"03",X"A9",X"DD",X"8D",X"0C",X"03",X"A9",X"7F",
		X"8D",X"0E",X"03",X"A9",X"00",X"8D",X"0B",X"03",X"60",X"A9",X"1A",X"20",X"07",X"FA",X"A9",X"20",
		X"A0",X"28",X"99",X"7F",X"BB",X"88",X"D0",X"FA",X"A9",X"00",X"8D",X"1F",X"02",X"A9",X"BB",X"8D",
		X"7B",X"02",X"8D",X"79",X"02",X"A9",X"A8",X"8D",X"7A",X"02",X"A9",X"D0",X"8D",X"78",X"02",X"A9",
		X"1B",X"8D",X"7E",X"02",X"A9",X"04",X"8D",X"7D",X"02",X"A9",X"10",X"8D",X"7C",X"02",X"A2",X"0C",
		X"20",X"38",X"02",X"20",X"5A",X"F7",X"60",X"8D",X"DF",X"BF",X"A9",X"02",X"A2",X"00",X"A0",X"03",
		X"20",X"C9",X"EE",X"60",X"A0",X"00",X"8C",X"60",X"02",X"8C",X"20",X"02",X"8C",X"00",X"05",X"84",
		X"0E",X"88",X"84",X"0C",X"8C",X"00",X"45",X"AD",X"00",X"05",X"D0",X"04",X"A9",X"C0",X"D0",X"05",
		X"EE",X"20",X"02",X"A9",X"40",X"85",X"0F",X"C8",X"A9",X"03",X"85",X"0D",X"E6",X"0C",X"D0",X"02",
		X"E6",X"0D",X"A5",X"0C",X"C5",X"0E",X"D0",X"06",X"A5",X"0D",X"C5",X"0F",X"F0",X"0F",X"A9",X"AA",
		X"91",X"0C",X"D1",X"0C",X"D0",X"07",X"4A",X"91",X"0C",X"D1",X"0C",X"F0",X"DF",X"38",X"A5",X"0F",
		X"E9",X"28",X"85",X"0F",X"A5",X"0E",X"C5",X"0C",X"A5",X"0F",X"E5",X"0D",X"90",X"09",X"A5",X"0C",
		X"A4",X"0D",X"EE",X"60",X"02",X"D0",X"04",X"A5",X"0E",X"A4",X"0F",X"85",X"A6",X"84",X"A7",X"8D",
		X"C1",X"02",X"8C",X"C2",X"02",X"60",X"08",X"78",X"86",X"14",X"84",X"15",X"A0",X"00",X"B1",X"14",
		X"AA",X"98",X"48",X"20",X"90",X"F5",X"68",X"A8",X"C8",X"C0",X"0E",X"D0",X"F1",X"28",X"60",X"A2",
		X"A7",X"A0",X"FA",X"20",X"86",X"FA",X"60",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"10",
		X"00",X"00",X"00",X"0F",X"00",X"A2",X"BD",X"A0",X"FA",X"20",X"86",X"FA",X"60",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"07",X"10",X"10",X"10",X"00",X"08",X"00",X"A2",X"D3",X"A0",X"FA",X"20",
		X"86",X"FA",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"07",X"10",X"10",X"10",X"00",X"18",
		X"00",X"A2",X"06",X"A0",X"FB",X"20",X"86",X"FA",X"A9",X"00",X"AA",X"8A",X"48",X"A9",X"00",X"20",
		X"90",X"F5",X"A2",X"00",X"CA",X"D0",X"FD",X"68",X"AA",X"E8",X"E0",X"70",X"D0",X"ED",X"A9",X"08",
		X"A2",X"00",X"20",X"90",X"F5",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"0F",X"00",
		X"00",X"00",X"00",X"00",X"A2",X"1C",X"A0",X"FB",X"20",X"86",X"FA",X"60",X"1F",X"00",X"00",X"00",
		X"00",X"00",X"00",X"3E",X"10",X"00",X"00",X"1F",X"00",X"00",X"A2",X"32",X"A0",X"FB",X"20",X"86",
		X"FA",X"60",X"2F",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"10",X"00",X"00",X"1F",X"00",X"00",
		X"AD",X"E1",X"02",X"C9",X"01",X"D0",X"22",X"A9",X"00",X"AE",X"E3",X"02",X"20",X"90",X"F5",X"A9",
		X"01",X"AE",X"E4",X"02",X"20",X"90",X"F5",X"AD",X"E5",X"02",X"29",X"0F",X"D0",X"04",X"A2",X"10",
		X"D0",X"01",X"AA",X"A9",X"08",X"20",X"90",X"F5",X"60",X"C9",X"02",X"D0",X"22",X"A9",X"02",X"AE",
		X"E3",X"02",X"20",X"90",X"F5",X"A9",X"03",X"AE",X"E4",X"02",X"20",X"90",X"F5",X"AD",X"E5",X"02",
		X"29",X"0F",X"D0",X"04",X"A2",X"10",X"D0",X"01",X"AA",X"A9",X"09",X"20",X"90",X"F5",X"60",X"C9",
		X"03",X"D0",X"22",X"A9",X"04",X"AE",X"E3",X"02",X"20",X"90",X"F5",X"A9",X"05",X"AE",X"E4",X"02",
		X"20",X"90",X"F5",X"AD",X"E5",X"02",X"29",X"0F",X"D0",X"04",X"A2",X"10",X"D0",X"01",X"AA",X"A9",
		X"0A",X"20",X"90",X"F5",X"60",X"A9",X"06",X"AE",X"E3",X"02",X"20",X"90",X"F5",X"AD",X"E1",X"02",
		X"C9",X"04",X"F0",X"93",X"C9",X"05",X"F0",X"B5",X"C9",X"06",X"F0",X"D7",X"EE",X"E0",X"02",X"60",
		X"AD",X"E3",X"02",X"0A",X"0A",X"0A",X"0D",X"E1",X"02",X"49",X"3F",X"AA",X"A9",X"07",X"20",X"90",
		X"F5",X"18",X"AD",X"E7",X"02",X"0A",X"8D",X"E7",X"02",X"AD",X"E8",X"02",X"2A",X"8D",X"E8",X"02",
		X"A9",X"0B",X"AE",X"E7",X"02",X"20",X"90",X"F5",X"A9",X"0C",X"AE",X"E8",X"02",X"20",X"90",X"F5",
		X"AD",X"E5",X"02",X"29",X"07",X"A8",X"B9",X"10",X"FC",X"AA",X"A9",X"0D",X"20",X"90",X"F5",X"60",
		X"00",X"00",X"04",X"08",X"0A",X"0B",X"0C",X"0D",X"A2",X"E1",X"A9",X"04",X"20",X"E4",X"F2",X"B0",
		X"39",X"A2",X"E3",X"A9",X"08",X"20",X"F8",X"F2",X"B0",X"30",X"A2",X"E5",X"A9",X"0D",X"20",X"E4",
		X"F2",X"B0",X"27",X"AC",X"E3",X"02",X"AE",X"E5",X"02",X"BD",X"5E",X"FC",X"8D",X"E4",X"02",X"BD",
		X"6B",X"FC",X"8D",X"E3",X"02",X"AD",X"E7",X"02",X"8D",X"E5",X"02",X"88",X"30",X"09",X"4E",X"E4",
		X"02",X"6E",X"E3",X"02",X"4C",X"4B",X"FC",X"4C",X"40",X"FB",X"EE",X"E0",X"02",X"60",X"00",X"07",
		X"07",X"06",X"06",X"05",X"05",X"05",X"04",X"04",X"04",X"04",X"03",X"00",X"77",X"0B",X"A6",X"47",
		X"EC",X"97",X"47",X"FB",X"B3",X"70",X"30",X"F4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"08",X"08",X"08",X"08",X"00",X"08",X"00",X"14",X"14",X"14",X"00",X"00",X"00",X"00",X"00",
		X"14",X"14",X"3E",X"14",X"3E",X"14",X"14",X"00",X"08",X"1E",X"28",X"1C",X"0A",X"3C",X"08",X"00",
		X"30",X"32",X"04",X"08",X"10",X"26",X"06",X"00",X"10",X"28",X"28",X"10",X"2A",X"24",X"1A",X"00",
		X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"08",X"10",X"20",X"20",X"20",X"10",X"08",X"00",
		X"08",X"04",X"02",X"02",X"02",X"04",X"08",X"00",X"08",X"2A",X"1C",X"08",X"1C",X"2A",X"08",X"00",
		X"00",X"08",X"08",X"3E",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"10",
		X"00",X"00",X"00",X"3E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",
		X"00",X"02",X"04",X"08",X"10",X"20",X"00",X"00",X"1C",X"22",X"26",X"2A",X"32",X"22",X"1C",X"00",
		X"08",X"18",X"08",X"08",X"08",X"08",X"1C",X"00",X"1C",X"22",X"02",X"04",X"08",X"10",X"3E",X"00",
		X"3E",X"02",X"04",X"0C",X"02",X"22",X"1C",X"00",X"04",X"0C",X"14",X"24",X"3E",X"04",X"04",X"00",
		X"3E",X"20",X"3C",X"02",X"02",X"22",X"1C",X"00",X"0C",X"10",X"20",X"3C",X"22",X"22",X"1C",X"00",
		X"3E",X"02",X"04",X"08",X"10",X"10",X"10",X"00",X"1C",X"22",X"22",X"1C",X"22",X"22",X"1C",X"00",
		X"1C",X"22",X"22",X"1E",X"02",X"04",X"18",X"00",X"00",X"00",X"08",X"00",X"00",X"08",X"00",X"00",
		X"00",X"00",X"08",X"00",X"00",X"08",X"08",X"10",X"04",X"08",X"10",X"20",X"10",X"08",X"04",X"00",
		X"00",X"00",X"3E",X"00",X"3E",X"00",X"00",X"00",X"10",X"08",X"04",X"02",X"04",X"08",X"10",X"00",
		X"1C",X"22",X"04",X"08",X"08",X"00",X"08",X"00",X"1C",X"22",X"2A",X"2E",X"2C",X"20",X"1E",X"00",
		X"08",X"14",X"22",X"22",X"3E",X"22",X"22",X"00",X"3C",X"22",X"22",X"3C",X"22",X"22",X"3C",X"00",
		X"1C",X"22",X"20",X"20",X"20",X"22",X"1C",X"00",X"3C",X"22",X"22",X"22",X"22",X"22",X"3C",X"00",
		X"3E",X"20",X"20",X"3C",X"20",X"20",X"3E",X"00",X"3E",X"20",X"20",X"3C",X"20",X"20",X"20",X"00",
		X"1E",X"20",X"20",X"20",X"26",X"22",X"1E",X"00",X"22",X"22",X"22",X"3E",X"22",X"22",X"22",X"00",
		X"1C",X"08",X"08",X"08",X"08",X"08",X"1C",X"00",X"02",X"02",X"02",X"02",X"02",X"22",X"1C",X"00",
		X"22",X"24",X"28",X"30",X"28",X"24",X"22",X"00",X"20",X"20",X"20",X"20",X"20",X"20",X"3E",X"00",
		X"22",X"36",X"2A",X"2A",X"22",X"22",X"22",X"00",X"22",X"22",X"32",X"2A",X"26",X"22",X"22",X"00",
		X"1C",X"22",X"22",X"22",X"22",X"22",X"1C",X"00",X"3C",X"22",X"22",X"3C",X"20",X"20",X"20",X"00",
		X"1C",X"22",X"22",X"22",X"2A",X"24",X"1A",X"00",X"3C",X"22",X"22",X"3C",X"28",X"24",X"22",X"00",
		X"1C",X"22",X"20",X"1C",X"02",X"22",X"1C",X"00",X"3E",X"08",X"08",X"08",X"08",X"08",X"08",X"00",
		X"22",X"22",X"22",X"22",X"22",X"22",X"1C",X"00",X"22",X"22",X"22",X"22",X"22",X"14",X"08",X"00",
		X"22",X"22",X"22",X"2A",X"2A",X"36",X"22",X"00",X"22",X"22",X"14",X"08",X"14",X"22",X"22",X"00",
		X"22",X"22",X"14",X"08",X"08",X"08",X"08",X"00",X"3E",X"02",X"04",X"08",X"10",X"20",X"3E",X"00",
		X"1E",X"10",X"10",X"10",X"10",X"10",X"1E",X"00",X"00",X"20",X"10",X"08",X"04",X"02",X"00",X"00",
		X"3C",X"04",X"04",X"04",X"04",X"04",X"3C",X"00",X"08",X"14",X"2A",X"08",X"08",X"08",X"08",X"00",
		X"0E",X"10",X"10",X"10",X"3C",X"10",X"3E",X"00",X"0C",X"12",X"2D",X"29",X"29",X"2D",X"12",X"0C",
		X"00",X"00",X"1C",X"02",X"1E",X"22",X"1E",X"00",X"20",X"20",X"3C",X"22",X"22",X"22",X"3C",X"00",
		X"00",X"00",X"1E",X"20",X"20",X"20",X"1E",X"00",X"02",X"02",X"1E",X"22",X"22",X"22",X"1E",X"00",
		X"00",X"00",X"1C",X"22",X"3E",X"20",X"1E",X"00",X"0C",X"12",X"10",X"3C",X"10",X"10",X"10",X"00",
		X"00",X"00",X"1C",X"22",X"22",X"1E",X"02",X"1C",X"20",X"20",X"3C",X"22",X"22",X"22",X"22",X"00",
		X"08",X"00",X"18",X"08",X"08",X"08",X"1C",X"00",X"04",X"00",X"0C",X"04",X"04",X"04",X"24",X"18",
		X"20",X"20",X"22",X"24",X"38",X"24",X"22",X"00",X"18",X"08",X"08",X"08",X"08",X"08",X"1C",X"00",
		X"00",X"00",X"36",X"2A",X"2A",X"2A",X"22",X"00",X"00",X"00",X"3C",X"22",X"22",X"22",X"22",X"00",
		X"00",X"00",X"1C",X"22",X"22",X"22",X"1C",X"00",X"00",X"00",X"3C",X"22",X"22",X"3C",X"20",X"20",
		X"00",X"00",X"1E",X"22",X"22",X"1E",X"02",X"02",X"00",X"00",X"2E",X"30",X"20",X"20",X"20",X"00",
		X"00",X"00",X"1E",X"20",X"1C",X"02",X"3C",X"00",X"10",X"10",X"3C",X"10",X"10",X"12",X"0C",X"00",
		X"00",X"00",X"22",X"22",X"22",X"26",X"1A",X"00",X"00",X"00",X"22",X"22",X"22",X"14",X"08",X"00",
		X"00",X"00",X"22",X"22",X"2A",X"2A",X"36",X"00",X"00",X"00",X"22",X"14",X"08",X"14",X"22",X"00",
		X"00",X"00",X"22",X"22",X"22",X"1E",X"02",X"1C",X"00",X"00",X"3E",X"04",X"08",X"10",X"3E",X"00",
		X"0E",X"18",X"18",X"30",X"18",X"18",X"0E",X"00",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"38",X"0C",X"0C",X"06",X"0C",X"0C",X"38",X"00",X"2A",X"15",X"2A",X"15",X"2A",X"15",X"2A",X"15",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"37",X"EA",X"ED",X"EB",X"20",X"F5",X"F9",X"38",
		X"EE",X"F4",X"36",X"39",X"2C",X"E9",X"E8",X"EC",X"35",X"F2",X"E2",X"3B",X"2E",X"EF",X"E7",X"30",
		X"F6",X"E6",X"34",X"2D",X"0B",X"F0",X"E5",X"2F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"31",X"1B",X"FA",X"5C",X"08",X"7F",X"E1",X"0D",X"F8",X"F1",X"32",X"23",X"0A",X"5D",X"F3",X"00",
		X"33",X"E4",X"E3",X"27",X"09",X"5B",X"F7",X"3D",X"26",X"4A",X"4D",X"4B",X"20",X"55",X"59",X"2A",
		X"4E",X"54",X"5E",X"28",X"3C",X"49",X"48",X"4C",X"25",X"52",X"42",X"3A",X"3E",X"4F",X"47",X"29",
		X"56",X"46",X"24",X"5F",X"0B",X"50",X"45",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"21",X"1B",X"5A",X"7C",X"08",X"7F",X"41",X"0D",X"58",X"51",X"22",X"7E",X"0A",X"7D",X"53",X"00",
		X"5F",X"44",X"43",X"40",X"09",X"7B",X"57",X"2B",X"D0",X"01",X"47",X"02",X"8F",X"F8",X"44",X"02");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
