library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity bg_graphx is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of bg_graphx is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"88",X"CC",X"22",X"22",X"66",X"CC",X"88",X"00",X"33",X"77",X"CC",X"88",X"88",X"77",X"33",X"00",
		X"22",X"22",X"EE",X"EE",X"22",X"22",X"00",X"00",X"00",X"00",X"FF",X"FF",X"44",X"00",X"00",X"00",
		X"22",X"22",X"AA",X"AA",X"EE",X"EE",X"66",X"00",X"66",X"FF",X"BB",X"99",X"99",X"CC",X"44",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"66",X"44",X"00",X"88",X"DD",X"FF",X"BB",X"99",X"88",X"00",X"00",
		X"88",X"EE",X"EE",X"88",X"88",X"88",X"88",X"00",X"00",X"FF",X"FF",X"CC",X"66",X"33",X"11",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"66",X"44",X"00",X"11",X"BB",X"AA",X"AA",X"AA",X"EE",X"EE",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"EE",X"CC",X"00",X"00",X"99",X"99",X"99",X"DD",X"77",X"33",X"00",
		X"00",X"00",X"00",X"EE",X"EE",X"00",X"00",X"00",X"CC",X"EE",X"BB",X"99",X"88",X"CC",X"CC",X"00",
		X"CC",X"EE",X"AA",X"AA",X"22",X"22",X"CC",X"00",X"00",X"66",X"99",X"99",X"BB",X"FF",X"66",X"00",
		X"88",X"CC",X"66",X"22",X"22",X"22",X"00",X"00",X"77",X"FF",X"99",X"99",X"99",X"FF",X"66",X"00",
		X"EE",X"EE",X"88",X"88",X"88",X"EE",X"EE",X"00",X"33",X"77",X"CC",X"88",X"CC",X"77",X"33",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"EE",X"EE",X"00",X"66",X"FF",X"99",X"99",X"99",X"FF",X"FF",X"00",
		X"44",X"66",X"22",X"22",X"66",X"CC",X"88",X"00",X"44",X"CC",X"88",X"88",X"CC",X"77",X"33",X"00",
		X"88",X"CC",X"66",X"22",X"22",X"EE",X"EE",X"00",X"33",X"77",X"CC",X"88",X"88",X"FF",X"FF",X"00",
		X"22",X"22",X"22",X"22",X"EE",X"EE",X"00",X"00",X"88",X"99",X"99",X"99",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"00",X"88",X"99",X"99",X"99",X"99",X"FF",X"FF",X"00",
		X"EE",X"EE",X"22",X"22",X"66",X"CC",X"88",X"00",X"99",X"99",X"99",X"88",X"CC",X"77",X"33",X"00",
		X"EE",X"EE",X"00",X"00",X"00",X"EE",X"EE",X"00",X"FF",X"FF",X"11",X"11",X"11",X"FF",X"FF",X"00",
		X"22",X"22",X"EE",X"EE",X"22",X"22",X"00",X"00",X"88",X"88",X"FF",X"FF",X"88",X"88",X"00",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"66",X"44",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"22",X"66",X"EE",X"CC",X"88",X"EE",X"EE",X"00",X"88",X"CC",X"66",X"33",X"11",X"FF",X"FF",X"00",
		X"22",X"22",X"22",X"22",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"EE",X"EE",X"00",X"88",X"00",X"EE",X"EE",X"00",X"FF",X"FF",X"77",X"33",X"77",X"FF",X"FF",X"00",
		X"EE",X"EE",X"CC",X"88",X"00",X"EE",X"EE",X"00",X"FF",X"FF",X"11",X"33",X"77",X"FF",X"FF",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"EE",X"CC",X"00",X"77",X"FF",X"88",X"88",X"88",X"FF",X"77",X"00",
		X"00",X"88",X"88",X"88",X"88",X"EE",X"EE",X"00",X"77",X"FF",X"88",X"88",X"88",X"FF",X"FF",X"00",
		X"AA",X"CC",X"EE",X"AA",X"22",X"EE",X"CC",X"00",X"77",X"FF",X"88",X"88",X"88",X"FF",X"77",X"00",
		X"22",X"66",X"EE",X"CC",X"88",X"EE",X"EE",X"00",X"77",X"FF",X"99",X"88",X"88",X"FF",X"FF",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"66",X"44",X"00",X"00",X"55",X"DD",X"99",X"99",X"FF",X"66",X"00",
		X"00",X"00",X"EE",X"EE",X"00",X"00",X"00",X"00",X"88",X"88",X"FF",X"FF",X"88",X"88",X"00",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"EE",X"CC",X"00",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"00",
		X"00",X"88",X"CC",X"EE",X"CC",X"88",X"00",X"00",X"FF",X"FF",X"11",X"00",X"11",X"FF",X"FF",X"00",
		X"EE",X"EE",X"CC",X"88",X"CC",X"EE",X"EE",X"00",X"FF",X"FF",X"11",X"33",X"11",X"FF",X"FF",X"00",
		X"66",X"EE",X"CC",X"88",X"CC",X"EE",X"66",X"00",X"CC",X"EE",X"77",X"33",X"77",X"EE",X"CC",X"00",
		X"00",X"00",X"EE",X"EE",X"00",X"00",X"00",X"00",X"EE",X"FF",X"11",X"11",X"FF",X"EE",X"00",X"00",
		X"22",X"22",X"22",X"AA",X"EE",X"EE",X"66",X"00",X"CC",X"EE",X"FF",X"BB",X"99",X"88",X"88",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"FF",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"44",X"AA",X"44",X"00",X"88",X"44",X"22",X"00",X"88",X"44",X"22",X"11",X"44",X"AA",X"44",X"00",
		X"00",X"00",X"00",X"00",X"66",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"00",X"CC",X"EE",X"FF",X"33",X"00",X"00",
		X"FF",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"22",X"11",X"55",X"55",X"99",X"22",X"CC",X"33",X"44",X"88",X"AA",X"AA",X"99",X"44",X"33",
		X"00",X"00",X"00",X"00",X"0F",X"0F",X"00",X"00",X"0C",X"0C",X"0C",X"0C",X"0F",X"0F",X"00",X"00",
		X"0B",X"0B",X"0F",X"0F",X"00",X"00",X"0F",X"0F",X"0D",X"0D",X"0D",X"01",X"00",X"00",X"07",X"0F",
		X"0F",X"00",X"00",X"0F",X"0F",X"0F",X"0B",X"0B",X"0F",X"00",X"00",X"07",X"0F",X"0F",X"0D",X"0D",
		X"0F",X"00",X"00",X"0F",X"0F",X"00",X"00",X"0F",X"0F",X"0C",X"0C",X"0F",X"0F",X"0C",X"0C",X"0F",
		X"03",X"03",X"03",X"0F",X"0E",X"00",X"00",X"0F",X"0C",X"0C",X"0C",X"0F",X"07",X"00",X"00",X"07",
		X"03",X"0F",X"0E",X"00",X"00",X"03",X"03",X"03",X"0C",X"0F",X"07",X"00",X"00",X"0C",X"0C",X"0C",
		X"00",X"00",X"0E",X"0F",X"03",X"03",X"03",X"03",X"00",X"00",X"07",X"0F",X"0C",X"0C",X"0C",X"0C",
		X"00",X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"88",X"CC",X"6E",X"BF",X"6E",X"CC",X"88",X"00",X"F3",X"E3",X"F3",X"F3",X"F3",X"E3",X"F3",
		X"00",X"F0",X"FB",X"FB",X"FA",X"FE",X"FE",X"F0",X"00",X"32",X"32",X"32",X"32",X"32",X"32",X"32",
		X"00",X"88",X"4C",X"AE",X"DF",X"AE",X"4C",X"88",X"00",X"F3",X"FB",X"FB",X"FB",X"FB",X"FB",X"F3",
		X"0F",X"6F",X"CF",X"8F",X"AF",X"BF",X"FF",X"00",X"23",X"33",X"33",X"33",X"33",X"33",X"33",X"00",
		X"7F",X"EE",X"CC",X"88",X"00",X"00",X"00",X"00",X"0F",X"7F",X"0F",X"BF",X"FF",X"EE",X"CC",X"00",
		X"00",X"00",X"FF",X"BF",X"AF",X"8F",X"CF",X"6F",X"00",X"00",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"88",X"CC",X"EE",X"00",X"00",X"CC",X"EE",X"FF",X"BF",X"0F",X"7F",
		X"0F",X"96",X"3C",X"78",X"78",X"2D",X"87",X"F0",X"87",X"D2",X"F0",X"E1",X"E1",X"F0",X"F0",X"F0",
		X"78",X"68",X"48",X"80",X"00",X"00",X"00",X"00",X"5A",X"D2",X"C3",X"96",X"3C",X"68",X"C0",X"80",
		X"00",X"F0",X"87",X"2D",X"78",X"78",X"3C",X"96",X"00",X"F0",X"F0",X"F0",X"E1",X"E1",X"F0",X"D2",
		X"00",X"00",X"00",X"00",X"00",X"80",X"48",X"68",X"00",X"80",X"C0",X"68",X"3C",X"96",X"C3",X"D2",
		X"FF",X"FF",X"DD",X"FF",X"BB",X"FF",X"FF",X"0F",X"7F",X"7F",X"0F",X"0F",X"1F",X"3F",X"1F",X"0F",
		X"0F",X"0E",X"8C",X"08",X"00",X"00",X"00",X"00",X"FF",X"77",X"9F",X"0F",X"8F",X"0E",X"CC",X"08",
		X"00",X"0F",X"FF",X"FF",X"BB",X"FF",X"DD",X"FF",X"00",X"0F",X"1F",X"3F",X"1F",X"2F",X"2F",X"5D",
		X"00",X"00",X"00",X"00",X"00",X"08",X"8C",X"0E",X"00",X"08",X"CC",X"0E",X"8F",X"0F",X"9F",X"77",
		X"DF",X"DF",X"F0",X"F0",X"F0",X"F0",X"DF",X"DF",X"EF",X"EF",X"FC",X"FC",X"FC",X"FC",X"EF",X"EF",
		X"F7",X"EE",X"CC",X"88",X"00",X"00",X"00",X"00",X"F8",X"F0",X"F1",X"F3",X"F7",X"EE",X"CC",X"88",
		X"00",X"DF",X"DF",X"F0",X"F0",X"F0",X"F0",X"DF",X"00",X"EF",X"EF",X"FC",X"FC",X"FC",X"FC",X"EF",
		X"00",X"00",X"00",X"00",X"00",X"88",X"CC",X"EE",X"00",X"88",X"CC",X"EE",X"F7",X"F3",X"F1",X"F0",
		X"FE",X"FF",X"11",X"00",X"71",X"00",X"10",X"00",X"77",X"11",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"00",X"71",X"00",X"11",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",
		X"EE",X"88",X"C0",X"C0",X"88",X"CC",X"EE",X"00",X"F7",X"F3",X"FE",X"7F",X"BF",X"11",X"F7",X"00",
		X"00",X"00",X"EE",X"CC",X"88",X"C0",X"C0",X"88",X"00",X"00",X"F7",X"11",X"BF",X"7F",X"FE",X"F3",
		X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"18",X"18",X"10",X"20",X"40",X"51",X"91",X"22",X"00",X"00",X"01",X"01",X"0E",X"00",X"10",X"E0",
		X"22",X"91",X"51",X"40",X"20",X"10",X"18",X"18",X"E0",X"10",X"00",X"0E",X"01",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"51",X"91",X"22",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"18",X"18",X"18",X"10",X"10",X"20",X"20",X"40",X"44",X"44",X"44",X"89",X"89",X"01",X"02",X"02",
		X"40",X"20",X"20",X"10",X"10",X"18",X"18",X"18",X"02",X"02",X"01",X"89",X"89",X"44",X"44",X"44",
		X"00",X"00",X"00",X"00",X"00",X"22",X"91",X"51",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",
		X"51",X"51",X"51",X"A2",X"00",X"00",X"00",X"00",X"02",X"02",X"04",X"00",X"00",X"00",X"00",X"00",
		X"18",X"18",X"18",X"18",X"18",X"20",X"20",X"20",X"44",X"44",X"44",X"44",X"44",X"45",X"89",X"89",
		X"20",X"20",X"20",X"18",X"18",X"18",X"18",X"18",X"89",X"89",X"45",X"44",X"44",X"44",X"44",X"44",
		X"00",X"00",X"00",X"00",X"A2",X"51",X"51",X"51",X"00",X"00",X"00",X"00",X"00",X"04",X"02",X"02",
		X"20",X"20",X"51",X"51",X"91",X"22",X"00",X"00",X"01",X"02",X"02",X"02",X"04",X"00",X"00",X"00",
		X"18",X"18",X"18",X"18",X"18",X"18",X"20",X"20",X"44",X"44",X"44",X"44",X"44",X"44",X"89",X"89",
		X"20",X"20",X"18",X"18",X"18",X"18",X"18",X"18",X"89",X"89",X"44",X"44",X"44",X"44",X"44",X"44",
		X"00",X"00",X"22",X"91",X"51",X"51",X"20",X"20",X"00",X"00",X"00",X"04",X"02",X"02",X"02",X"01",
		X"20",X"20",X"20",X"40",X"40",X"40",X"80",X"00",X"89",X"89",X"01",X"02",X"02",X"04",X"00",X"00",
		X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"20",X"44",X"44",X"44",X"44",X"44",X"44",X"88",X"89",
		X"20",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"89",X"88",X"44",X"44",X"44",X"44",X"44",X"44",
		X"00",X"80",X"40",X"40",X"40",X"20",X"20",X"20",X"00",X"00",X"04",X"02",X"02",X"01",X"89",X"89",
		X"91",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"20",X"20",X"20",X"40",X"40",X"40",X"40",X"89",X"89",X"89",X"89",X"8A",X"8A",X"8A",X"8C",
		X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"28",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"28",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"40",X"40",X"40",X"40",X"20",X"20",X"20",X"20",X"8C",X"8A",X"8A",X"8A",X"89",X"89",X"89",X"89",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"91",X"91",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"04",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"20",X"20",X"40",X"40",X"40",X"40",X"80",X"89",X"89",X"89",X"8A",X"8A",X"8A",X"8A",X"8C",
		X"18",X"18",X"18",X"18",X"18",X"28",X"28",X"28",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"28",X"28",X"28",X"18",X"18",X"18",X"18",X"18",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"80",X"40",X"40",X"40",X"40",X"20",X"20",X"20",X"8C",X"8A",X"8A",X"8A",X"8A",X"89",X"89",X"89",
		X"00",X"00",X"00",X"00",X"00",X"00",X"91",X"91",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"04",
		X"51",X"91",X"A2",X"A2",X"00",X"00",X"00",X"00",X"04",X"04",X"04",X"00",X"00",X"00",X"00",X"00",
		X"20",X"20",X"20",X"20",X"20",X"40",X"40",X"40",X"89",X"89",X"89",X"89",X"8A",X"8A",X"8A",X"8A",
		X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"88",
		X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"88",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"40",X"40",X"40",X"20",X"20",X"20",X"20",X"20",X"8A",X"8A",X"8A",X"8A",X"89",X"89",X"89",X"89",
		X"00",X"00",X"00",X"00",X"A2",X"A2",X"91",X"51",X"00",X"00",X"00",X"00",X"00",X"04",X"04",X"04",
		X"51",X"51",X"91",X"A2",X"A2",X"22",X"00",X"00",X"02",X"02",X"02",X"04",X"04",X"00",X"00",X"00",
		X"20",X"20",X"20",X"20",X"20",X"40",X"40",X"40",X"89",X"89",X"89",X"89",X"89",X"89",X"8A",X"8A",
		X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"40",X"40",X"40",X"20",X"20",X"20",X"20",X"20",X"8A",X"8A",X"89",X"89",X"89",X"89",X"89",X"89",
		X"00",X"00",X"22",X"A2",X"A2",X"91",X"51",X"51",X"00",X"00",X"00",X"04",X"04",X"02",X"02",X"02",
		X"40",X"40",X"40",X"40",X"80",X"80",X"80",X"00",X"02",X"02",X"04",X"04",X"04",X"04",X"00",X"00",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"89",X"89",X"89",X"89",X"89",X"8A",X"8A",X"8A",
		X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"8A",X"8A",X"8A",X"89",X"89",X"89",X"89",X"89",
		X"00",X"80",X"80",X"80",X"40",X"40",X"40",X"40",X"00",X"00",X"04",X"04",X"04",X"04",X"02",X"02",
		X"11",X"33",X"44",X"44",X"66",X"33",X"11",X"00",X"CC",X"EE",X"33",X"11",X"11",X"EE",X"CC",X"00",
		X"44",X"44",X"77",X"77",X"44",X"44",X"00",X"00",X"00",X"00",X"FF",X"FF",X"22",X"00",X"00",X"00",
		X"44",X"44",X"55",X"55",X"77",X"77",X"66",X"00",X"66",X"FF",X"DD",X"99",X"99",X"33",X"22",X"00",
		X"33",X"77",X"44",X"44",X"44",X"66",X"22",X"00",X"11",X"BB",X"FF",X"DD",X"99",X"11",X"00",X"00",
		X"11",X"77",X"77",X"11",X"11",X"11",X"11",X"00",X"00",X"FF",X"FF",X"33",X"66",X"CC",X"88",X"00",
		X"33",X"77",X"44",X"44",X"44",X"66",X"22",X"00",X"88",X"DD",X"55",X"55",X"55",X"77",X"77",X"00",
		X"33",X"77",X"44",X"44",X"44",X"77",X"33",X"00",X"00",X"99",X"99",X"99",X"BB",X"EE",X"CC",X"00",
		X"00",X"00",X"00",X"77",X"77",X"00",X"00",X"00",X"33",X"77",X"DD",X"99",X"11",X"33",X"33",X"00",
		X"33",X"77",X"55",X"55",X"44",X"44",X"33",X"00",X"00",X"66",X"99",X"99",X"DD",X"FF",X"66",X"00",
		X"11",X"33",X"66",X"44",X"44",X"44",X"00",X"00",X"EE",X"FF",X"99",X"99",X"99",X"FF",X"66",X"00",
		X"77",X"77",X"11",X"11",X"11",X"77",X"77",X"00",X"CC",X"EE",X"33",X"11",X"33",X"EE",X"CC",X"00",
		X"33",X"77",X"44",X"44",X"44",X"77",X"77",X"00",X"66",X"FF",X"99",X"99",X"99",X"FF",X"FF",X"00",
		X"22",X"66",X"44",X"44",X"66",X"33",X"11",X"00",X"22",X"33",X"11",X"11",X"33",X"EE",X"CC",X"00",
		X"11",X"33",X"66",X"44",X"44",X"77",X"77",X"00",X"CC",X"EE",X"33",X"11",X"11",X"FF",X"FF",X"00",
		X"44",X"44",X"44",X"44",X"77",X"77",X"00",X"00",X"11",X"99",X"99",X"99",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"77",X"77",X"00",X"11",X"99",X"99",X"99",X"99",X"FF",X"FF",X"00",
		X"77",X"77",X"44",X"44",X"66",X"33",X"11",X"00",X"99",X"99",X"99",X"11",X"33",X"EE",X"CC",X"00",
		X"77",X"77",X"00",X"00",X"00",X"77",X"77",X"00",X"FF",X"FF",X"88",X"88",X"88",X"FF",X"FF",X"00",
		X"44",X"44",X"77",X"77",X"44",X"44",X"00",X"00",X"11",X"11",X"FF",X"FF",X"11",X"11",X"00",X"00",
		X"33",X"77",X"44",X"44",X"44",X"66",X"22",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"66",X"77",X"33",X"11",X"77",X"77",X"00",X"11",X"33",X"66",X"CC",X"88",X"FF",X"FF",X"00",
		X"44",X"44",X"44",X"44",X"77",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"77",X"77",X"00",X"11",X"00",X"77",X"77",X"00",X"FF",X"FF",X"EE",X"CC",X"EE",X"FF",X"FF",X"00",
		X"77",X"77",X"33",X"11",X"00",X"77",X"77",X"00",X"FF",X"FF",X"88",X"CC",X"EE",X"FF",X"FF",X"00",
		X"33",X"77",X"44",X"44",X"44",X"77",X"33",X"00",X"EE",X"FF",X"11",X"11",X"11",X"FF",X"EE",X"00",
		X"00",X"11",X"11",X"11",X"11",X"77",X"77",X"00",X"EE",X"FF",X"11",X"11",X"11",X"FF",X"FF",X"00",
		X"55",X"33",X"77",X"55",X"44",X"77",X"33",X"00",X"EE",X"FF",X"11",X"11",X"11",X"FF",X"EE",X"00",
		X"44",X"66",X"77",X"33",X"11",X"77",X"77",X"00",X"EE",X"FF",X"99",X"11",X"11",X"FF",X"FF",X"00",
		X"33",X"77",X"44",X"44",X"44",X"66",X"22",X"00",X"00",X"AA",X"BB",X"99",X"99",X"FF",X"66",X"00",
		X"00",X"00",X"77",X"77",X"00",X"00",X"00",X"00",X"11",X"11",X"FF",X"FF",X"11",X"11",X"00",X"00",
		X"33",X"77",X"44",X"44",X"44",X"77",X"33",X"00",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"00",
		X"00",X"11",X"33",X"77",X"33",X"11",X"00",X"00",X"FF",X"FF",X"88",X"00",X"88",X"FF",X"FF",X"00",
		X"77",X"77",X"33",X"11",X"33",X"77",X"77",X"00",X"FF",X"FF",X"88",X"CC",X"88",X"FF",X"FF",X"00",
		X"66",X"77",X"33",X"11",X"33",X"77",X"66",X"00",X"33",X"77",X"EE",X"CC",X"EE",X"77",X"33",X"00",
		X"00",X"00",X"77",X"77",X"00",X"00",X"00",X"00",X"77",X"FF",X"88",X"88",X"FF",X"77",X"00",X"00",
		X"44",X"44",X"44",X"55",X"77",X"77",X"66",X"00",X"33",X"77",X"FF",X"DD",X"99",X"11",X"11",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"FF",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"22",X"55",X"22",X"00",X"11",X"22",X"44",X"00",X"11",X"22",X"44",X"88",X"22",X"55",X"22",X"00",
		X"00",X"00",X"00",X"00",X"66",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"00",X"33",X"77",X"FF",X"CC",X"00",X"00",
		X"FF",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"44",X"88",X"AA",X"AA",X"99",X"44",X"33",X"CC",X"22",X"11",X"55",X"55",X"99",X"22",X"CC",
		X"00",X"00",X"00",X"00",X"0F",X"0F",X"00",X"00",X"03",X"03",X"03",X"03",X"0F",X"0F",X"00",X"00",
		X"0D",X"0D",X"0F",X"0F",X"00",X"00",X"0F",X"0F",X"0B",X"0B",X"0B",X"08",X"00",X"00",X"0E",X"0F",
		X"0F",X"00",X"00",X"0F",X"0F",X"0F",X"0D",X"0D",X"0F",X"00",X"00",X"0E",X"0F",X"0F",X"0B",X"0B",
		X"0F",X"00",X"00",X"0F",X"0F",X"00",X"00",X"0F",X"0F",X"03",X"03",X"0F",X"0F",X"03",X"03",X"0F",
		X"0C",X"0C",X"0C",X"0F",X"07",X"00",X"00",X"0F",X"03",X"03",X"03",X"0F",X"0E",X"00",X"00",X"0E",
		X"0C",X"0F",X"07",X"00",X"00",X"0C",X"0C",X"0C",X"03",X"0F",X"0E",X"00",X"00",X"03",X"03",X"03",
		X"00",X"00",X"07",X"0F",X"0C",X"0C",X"0C",X"0C",X"00",X"00",X"0E",X"0F",X"03",X"03",X"03",X"03",
		X"00",X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"33",X"67",X"DF",X"67",X"33",X"11",X"00",X"FC",X"7C",X"FC",X"FC",X"FC",X"7C",X"FC",
		X"00",X"F0",X"FD",X"FD",X"F5",X"F7",X"F7",X"F0",X"00",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",
		X"00",X"11",X"23",X"57",X"BF",X"57",X"23",X"11",X"00",X"FC",X"FD",X"FD",X"FD",X"FD",X"FD",X"FC",
		X"0F",X"6F",X"3F",X"1F",X"5F",X"DF",X"FF",X"00",X"4C",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"00",
		X"EF",X"77",X"33",X"11",X"00",X"00",X"00",X"00",X"0F",X"EF",X"0F",X"DF",X"FF",X"77",X"33",X"00",
		X"00",X"00",X"FF",X"DF",X"5F",X"1F",X"3F",X"6F",X"00",X"00",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"77",X"00",X"00",X"33",X"77",X"FF",X"DF",X"0F",X"EF",
		X"0F",X"96",X"C3",X"E1",X"E1",X"4B",X"1E",X"F0",X"1E",X"B4",X"F0",X"78",X"78",X"F0",X"F0",X"F0",
		X"E1",X"61",X"21",X"10",X"00",X"00",X"00",X"00",X"A5",X"B4",X"3C",X"96",X"C3",X"61",X"30",X"10",
		X"00",X"F0",X"1E",X"4B",X"E1",X"E1",X"C3",X"96",X"00",X"F0",X"F0",X"F0",X"78",X"78",X"F0",X"B4",
		X"00",X"00",X"00",X"00",X"00",X"10",X"21",X"61",X"00",X"10",X"30",X"61",X"C3",X"96",X"3C",X"B4",
		X"FF",X"FF",X"BB",X"FF",X"DD",X"FF",X"FF",X"0F",X"EF",X"EF",X"0F",X"0F",X"8F",X"CF",X"8F",X"0F",
		X"0F",X"07",X"13",X"01",X"00",X"00",X"00",X"00",X"FF",X"EE",X"9F",X"0F",X"1F",X"07",X"33",X"01",
		X"00",X"0F",X"FF",X"FF",X"DD",X"FF",X"BB",X"FF",X"00",X"0F",X"8F",X"CF",X"8F",X"4F",X"4F",X"AB",
		X"00",X"00",X"00",X"00",X"00",X"01",X"13",X"07",X"00",X"01",X"33",X"07",X"1F",X"0F",X"9F",X"EE",
		X"BF",X"BF",X"F0",X"F0",X"F0",X"F0",X"BF",X"BF",X"7F",X"7F",X"F3",X"F3",X"F3",X"F3",X"7F",X"7F",
		X"FE",X"77",X"33",X"11",X"00",X"00",X"00",X"00",X"F1",X"F0",X"F8",X"FC",X"FE",X"77",X"33",X"11",
		X"00",X"BF",X"BF",X"F0",X"F0",X"F0",X"F0",X"BF",X"00",X"7F",X"7F",X"F3",X"F3",X"F3",X"F3",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"77",X"00",X"11",X"33",X"77",X"FE",X"FC",X"F8",X"F0",
		X"F7",X"FF",X"88",X"00",X"E8",X"00",X"80",X"00",X"EE",X"88",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"00",X"E8",X"00",X"88",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",
		X"77",X"11",X"30",X"30",X"11",X"33",X"77",X"00",X"FE",X"FC",X"F7",X"EF",X"DF",X"88",X"FE",X"00",
		X"00",X"00",X"77",X"33",X"11",X"30",X"30",X"11",X"00",X"00",X"FE",X"88",X"DF",X"EF",X"F7",X"FC",
		X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"81",X"81",X"80",X"40",X"20",X"A8",X"98",X"44",X"00",X"00",X"08",X"08",X"07",X"00",X"80",X"70",
		X"44",X"98",X"A8",X"20",X"40",X"80",X"81",X"81",X"70",X"80",X"00",X"07",X"08",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A8",X"98",X"44",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"81",X"81",X"81",X"80",X"80",X"40",X"40",X"20",X"22",X"22",X"22",X"19",X"19",X"08",X"04",X"04",
		X"20",X"40",X"40",X"80",X"80",X"81",X"81",X"81",X"04",X"04",X"08",X"19",X"19",X"22",X"22",X"22",
		X"00",X"00",X"00",X"00",X"00",X"44",X"98",X"A8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",
		X"A8",X"A8",X"A8",X"54",X"00",X"00",X"00",X"00",X"04",X"04",X"02",X"00",X"00",X"00",X"00",X"00",
		X"81",X"81",X"81",X"81",X"81",X"40",X"40",X"40",X"22",X"22",X"22",X"22",X"22",X"2A",X"19",X"19",
		X"40",X"40",X"40",X"81",X"81",X"81",X"81",X"81",X"19",X"19",X"2A",X"22",X"22",X"22",X"22",X"22",
		X"00",X"00",X"00",X"00",X"54",X"A8",X"A8",X"A8",X"00",X"00",X"00",X"00",X"00",X"02",X"04",X"04",
		X"40",X"40",X"A8",X"A8",X"98",X"44",X"00",X"00",X"08",X"04",X"04",X"04",X"02",X"00",X"00",X"00",
		X"81",X"81",X"81",X"81",X"81",X"81",X"40",X"40",X"22",X"22",X"22",X"22",X"22",X"22",X"19",X"19",
		X"40",X"40",X"81",X"81",X"81",X"81",X"81",X"81",X"19",X"19",X"22",X"22",X"22",X"22",X"22",X"22",
		X"00",X"00",X"44",X"98",X"A8",X"A8",X"40",X"40",X"00",X"00",X"00",X"02",X"04",X"04",X"04",X"08",
		X"40",X"40",X"40",X"20",X"20",X"20",X"10",X"00",X"19",X"19",X"08",X"04",X"04",X"02",X"00",X"00",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"40",X"22",X"22",X"22",X"22",X"22",X"22",X"11",X"19",
		X"40",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"19",X"11",X"22",X"22",X"22",X"22",X"22",X"22",
		X"00",X"10",X"20",X"20",X"20",X"40",X"40",X"40",X"00",X"00",X"02",X"04",X"04",X"08",X"19",X"19",
		X"98",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"40",X"40",X"40",X"20",X"20",X"20",X"20",X"19",X"19",X"19",X"19",X"15",X"15",X"15",X"13",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"41",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"41",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"20",X"20",X"20",X"20",X"40",X"40",X"40",X"40",X"13",X"15",X"15",X"15",X"19",X"19",X"19",X"19",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"98",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"98",X"98",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"40",X"40",X"20",X"20",X"20",X"20",X"10",X"19",X"19",X"19",X"15",X"15",X"15",X"15",X"13",
		X"81",X"81",X"81",X"81",X"81",X"41",X"41",X"41",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"41",X"41",X"41",X"81",X"81",X"81",X"81",X"81",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"10",X"20",X"20",X"20",X"20",X"40",X"40",X"40",X"13",X"15",X"15",X"15",X"15",X"19",X"19",X"19",
		X"00",X"00",X"00",X"00",X"00",X"00",X"98",X"98",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"02",
		X"A8",X"98",X"54",X"54",X"00",X"00",X"00",X"00",X"02",X"02",X"02",X"00",X"00",X"00",X"00",X"00",
		X"40",X"40",X"40",X"40",X"40",X"20",X"20",X"20",X"19",X"19",X"19",X"19",X"15",X"15",X"15",X"15",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"11",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"11",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"20",X"20",X"20",X"40",X"40",X"40",X"40",X"40",X"15",X"15",X"15",X"15",X"19",X"19",X"19",X"19",
		X"00",X"00",X"00",X"00",X"54",X"54",X"98",X"A8",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"02",
		X"A8",X"A8",X"98",X"54",X"54",X"44",X"00",X"00",X"04",X"04",X"04",X"02",X"02",X"00",X"00",X"00",
		X"40",X"40",X"40",X"40",X"40",X"20",X"20",X"20",X"19",X"19",X"19",X"19",X"19",X"19",X"15",X"15",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"20",X"20",X"20",X"40",X"40",X"40",X"40",X"40",X"15",X"15",X"19",X"19",X"19",X"19",X"19",X"19",
		X"00",X"00",X"44",X"54",X"54",X"98",X"A8",X"A8",X"00",X"00",X"00",X"02",X"02",X"04",X"04",X"04",
		X"20",X"20",X"20",X"20",X"10",X"10",X"10",X"00",X"04",X"04",X"02",X"02",X"02",X"02",X"00",X"00",
		X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"19",X"19",X"19",X"19",X"19",X"15",X"15",X"15",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"15",X"15",X"15",X"19",X"19",X"19",X"19",X"19",
		X"00",X"10",X"10",X"10",X"20",X"20",X"20",X"20",X"00",X"00",X"02",X"02",X"02",X"02",X"04",X"04");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
