`define BUILD_DATE "190901"
`define BUILD_TIME "150452"
