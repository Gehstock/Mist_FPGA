library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity cmd_chr_rom is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of cmd_chr_rom is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"CC",X"EE",X"22",X"22",X"22",X"EE",X"CC",X"00",X"77",X"FF",X"88",X"88",X"88",X"FF",X"77",
		X"00",X"00",X"00",X"44",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"44",X"66",X"22",X"22",X"AA",X"EE",X"CC",X"00",X"CC",X"EE",X"FF",X"FF",X"BB",X"99",X"88",
		X"00",X"22",X"22",X"22",X"AA",X"EE",X"66",X"22",X"00",X"44",X"CC",X"99",X"99",X"99",X"FF",X"66",
		X"00",X"00",X"88",X"CC",X"66",X"EE",X"EE",X"00",X"00",X"33",X"33",X"22",X"22",X"FF",X"FF",X"22",
		X"00",X"EE",X"EE",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"44",X"CC",X"88",X"88",X"88",X"FF",X"77",
		X"00",X"88",X"CC",X"66",X"22",X"22",X"22",X"00",X"00",X"77",X"FF",X"99",X"99",X"99",X"FF",X"66",
		X"00",X"66",X"66",X"22",X"22",X"AA",X"EE",X"66",X"00",X"00",X"00",X"EE",X"FF",X"11",X"00",X"00",
		X"00",X"CC",X"EE",X"22",X"22",X"22",X"EE",X"CC",X"00",X"66",X"FF",X"99",X"99",X"99",X"FF",X"66",
		X"00",X"CC",X"EE",X"22",X"22",X"22",X"EE",X"CC",X"00",X"00",X"99",X"99",X"99",X"DD",X"77",X"33",
		X"00",X"88",X"CC",X"66",X"22",X"66",X"CC",X"88",X"00",X"FF",X"FF",X"22",X"22",X"22",X"FF",X"FF",
		X"00",X"EE",X"EE",X"22",X"22",X"22",X"EE",X"CC",X"00",X"FF",X"FF",X"99",X"99",X"99",X"FF",X"66",
		X"00",X"88",X"CC",X"66",X"22",X"22",X"66",X"44",X"00",X"33",X"77",X"CC",X"88",X"88",X"CC",X"44",
		X"00",X"EE",X"EE",X"22",X"22",X"66",X"CC",X"88",X"00",X"FF",X"FF",X"88",X"88",X"CC",X"77",X"33",
		X"00",X"EE",X"EE",X"22",X"22",X"22",X"22",X"22",X"00",X"FF",X"FF",X"99",X"99",X"99",X"99",X"88",
		X"00",X"EE",X"EE",X"22",X"22",X"22",X"22",X"22",X"00",X"FF",X"FF",X"11",X"11",X"11",X"11",X"00",
		X"00",X"88",X"CC",X"66",X"22",X"22",X"22",X"22",X"00",X"33",X"77",X"CC",X"88",X"99",X"FF",X"FF",
		X"00",X"EE",X"EE",X"00",X"00",X"00",X"EE",X"EE",X"00",X"FF",X"FF",X"11",X"11",X"11",X"FF",X"FF",
		X"00",X"00",X"00",X"22",X"EE",X"EE",X"22",X"00",X"00",X"00",X"00",X"88",X"FF",X"FF",X"88",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"00",X"44",X"CC",X"88",X"88",X"88",X"FF",X"77",
		X"00",X"EE",X"EE",X"00",X"88",X"CC",X"66",X"22",X"00",X"FF",X"FF",X"33",X"77",X"EE",X"CC",X"88",
		X"00",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"88",X"88",X"88",X"88",X"88",
		X"00",X"EE",X"EE",X"CC",X"88",X"CC",X"EE",X"EE",X"00",X"FF",X"FF",X"11",X"33",X"11",X"FF",X"FF",
		X"00",X"EE",X"EE",X"CC",X"88",X"00",X"EE",X"EE",X"00",X"FF",X"FF",X"11",X"33",X"77",X"FF",X"FF",
		X"00",X"CC",X"EE",X"22",X"22",X"22",X"EE",X"CC",X"00",X"77",X"FF",X"88",X"88",X"88",X"FF",X"77",
		X"00",X"EE",X"EE",X"22",X"22",X"22",X"EE",X"CC",X"00",X"FF",X"FF",X"22",X"22",X"22",X"33",X"11",
		X"00",X"CC",X"EE",X"22",X"22",X"22",X"EE",X"CC",X"00",X"77",X"FF",X"88",X"AA",X"EE",X"77",X"BB",
		X"00",X"EE",X"EE",X"22",X"22",X"22",X"EE",X"CC",X"00",X"FF",X"FF",X"22",X"66",X"FF",X"DD",X"99",
		X"00",X"CC",X"EE",X"22",X"22",X"22",X"66",X"44",X"00",X"44",X"DD",X"99",X"99",X"99",X"FF",X"66",
		X"00",X"22",X"22",X"EE",X"EE",X"22",X"22",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",
		X"00",X"EE",X"EE",X"00",X"00",X"00",X"EE",X"EE",X"00",X"77",X"FF",X"88",X"88",X"88",X"FF",X"77",
		X"00",X"EE",X"EE",X"00",X"00",X"00",X"EE",X"EE",X"00",X"11",X"33",X"77",X"EE",X"77",X"33",X"11",
		X"00",X"EE",X"EE",X"00",X"88",X"00",X"EE",X"EE",X"00",X"33",X"FF",X"77",X"33",X"77",X"FF",X"33",
		X"00",X"66",X"EE",X"CC",X"88",X"CC",X"EE",X"66",X"00",X"CC",X"EE",X"77",X"33",X"77",X"EE",X"CC",
		X"00",X"66",X"EE",X"00",X"00",X"EE",X"66",X"00",X"00",X"00",X"11",X"FF",X"FF",X"11",X"00",X"00",
		X"00",X"22",X"22",X"22",X"AA",X"EE",X"EE",X"66",X"00",X"CC",X"EE",X"FF",X"BB",X"99",X"88",X"88",
		X"CC",X"22",X"99",X"55",X"55",X"11",X"22",X"CC",X"33",X"44",X"99",X"AA",X"AA",X"88",X"44",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"33",X"FF",X"CC",X"00",X"00",X"00",X"00",X"CC",X"CC",X"FF",X"FF",X"EE",X"00",X"00",X"00",
		X"BB",X"BB",X"BB",X"00",X"00",X"00",X"CC",X"FF",X"00",X"FF",X"FF",X"00",X"CC",X"FF",X"FF",X"33",
		X"BB",X"33",X"00",X"00",X"EE",X"FF",X"33",X"33",X"DD",X"CC",X"00",X"00",X"77",X"FF",X"CC",X"CC",
		X"33",X"00",X"00",X"EE",X"FF",X"FF",X"BB",X"BB",X"77",X"00",X"00",X"77",X"FF",X"FF",X"DD",X"DD",
		X"00",X"00",X"EE",X"FF",X"FF",X"BB",X"BB",X"BB",X"00",X"00",X"CC",X"DD",X"DD",X"DD",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"D0",X"A0",X"50",X"A0",X"40",X"C0",X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"B0",X"70",X"B0",X"10",X"80",X"10",X"80",X"10",X"80",X"50",X"A0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"A0",X"C0",X"A0",X"40",X"80",
		X"70",X"B0",X"F0",X"70",X"F0",X"F0",X"D0",X"E0",X"F0",X"F0",X"E0",X"F0",X"D0",X"F0",X"F0",X"F0",
		X"00",X"00",X"80",X"80",X"40",X"80",X"40",X"A0",X"C0",X"F0",X"F0",X"E0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"40",X"80",X"60",X"E0",X"D0",X"E0",X"D0",X"A0",X"50",X"A0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"30",X"10",X"20",X"10",X"30",X"10",X"30",X"10",X"00",X"10",X"00",X"10",X"10",X"10",X"10",
		X"10",X"20",X"10",X"30",X"10",X"30",X"10",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"00",X"10",X"00",X"30",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"D0",X"E0",X"50",X"A0",X"40",X"80",X"80",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",
		X"70",X"F0",X"50",X"A0",X"00",X"00",X"00",X"00",X"10",X"00",X"10",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"D0",X"A0",X"D0",X"A0",X"40",X"80",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"A0",X"C0",
		X"48",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"4B",X"4B",X"5A",X"78",X"84",X"0C",X"00",X"00",
		X"78",X"78",X"D2",X"D2",X"96",X"96",X"E1",X"E1",X"C3",X"78",X"78",X"5A",X"4B",X"4B",X"D2",X"E1",
		X"B4",X"B4",X"96",X"96",X"D2",X"F0",X"5A",X"5A",X"96",X"96",X"C3",X"78",X"3C",X"69",X"69",X"4B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"48",X"00",X"00",X"C0",X"C0",X"B4",X"96",X"78",X"B4",
		X"0F",X"FF",X"FF",X"EE",X"EE",X"EE",X"CC",X"44",X"0F",X"77",X"33",X"33",X"11",X"11",X"00",X"00",
		X"7B",X"F3",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"4B",X"4B",X"5A",X"78",X"B7",X"3F",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F3",X"7B",X"FF",X"FF",X"F3",X"F3",X"B4",X"96",X"78",X"B4",
		X"0F",X"FF",X"FF",X"FE",X"FE",X"FE",X"FC",X"F4",X"0F",X"F7",X"F3",X"F3",X"F1",X"F0",X"F0",X"F0",
		X"00",X"22",X"44",X"88",X"00",X"88",X"44",X"22",X"00",X"88",X"44",X"22",X"11",X"22",X"44",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"00",
		X"0C",X"0E",X"0F",X"87",X"87",X"0F",X"0E",X"0C",X"61",X"41",X"C2",X"87",X"87",X"C2",X"41",X"A1",
		X"0F",X"0F",X"0F",X"0E",X"0E",X"0C",X"08",X"00",X"1E",X"0D",X"0B",X"07",X"0F",X"0F",X"0F",X"0E",
		X"0F",X"0F",X"0F",X"0F",X"0E",X"87",X"C3",X"61",X"C3",X"C3",X"C3",X"61",X"70",X"70",X"D0",X"80",
		X"00",X"08",X"0C",X"0E",X"0E",X"0F",X"0F",X"87",X"0E",X"0F",X"0F",X"07",X"0B",X"0D",X"1E",X"10",
		X"43",X"C3",X"86",X"0F",X"0F",X"0F",X"0F",X"00",X"80",X"D0",X"70",X"70",X"61",X"C3",X"C3",X"C2",
		X"0C",X"0E",X"0F",X"87",X"87",X"0F",X"0E",X"0C",X"A1",X"41",X"C2",X"87",X"87",X"C2",X"41",X"61",
		X"86",X"86",X"0C",X"0A",X"84",X"C0",X"84",X"80",X"42",X"86",X"94",X"96",X"1E",X"3C",X"48",X"18",
		X"08",X"0C",X"00",X"E0",X"80",X"48",X"2C",X"00",X"E0",X"30",X"12",X"21",X"21",X"21",X"52",X"52",
		X"08",X"2C",X"78",X"A4",X"0C",X"48",X"A4",X"B4",X"52",X"43",X"21",X"29",X"A5",X"90",X"30",X"E0",
		X"00",X"08",X"08",X"00",X"08",X"86",X"E0",X"87",X"09",X"1C",X"3C",X"29",X"A5",X"94",X"86",X"42",
		X"3F",X"1F",X"0F",X"87",X"87",X"0F",X"1F",X"3F",X"E9",X"EB",X"D3",X"87",X"87",X"D3",X"EB",X"E5",
		X"0F",X"0F",X"0F",X"1F",X"1F",X"3F",X"7F",X"FF",X"1E",X"2F",X"4F",X"8F",X"0F",X"0F",X"0F",X"1F",
		X"0F",X"0F",X"0F",X"0F",X"1F",X"87",X"C3",X"E9",X"C3",X"C3",X"C3",X"E9",X"F8",X"F8",X"F2",X"F7",
		X"FF",X"7F",X"3F",X"1F",X"1F",X"0F",X"0F",X"87",X"1F",X"0F",X"0F",X"8F",X"4F",X"2F",X"1E",X"FE",
		X"CB",X"C3",X"97",X"0F",X"0F",X"0F",X"0F",X"FF",X"F7",X"F2",X"F8",X"F8",X"E9",X"C3",X"C3",X"D3",
		X"3F",X"1F",X"0F",X"87",X"87",X"0F",X"1F",X"3F",X"E5",X"EB",X"D3",X"87",X"87",X"D3",X"EB",X"E9",
		X"97",X"97",X"3F",X"5F",X"B7",X"F3",X"B7",X"F7",X"DB",X"97",X"B6",X"96",X"1E",X"3C",X"7B",X"79",
		X"7F",X"3F",X"FF",X"F1",X"F7",X"7B",X"3D",X"FF",X"F1",X"FC",X"DE",X"ED",X"ED",X"ED",X"DA",X"DA",
		X"7F",X"3D",X"78",X"B5",X"3F",X"7B",X"B5",X"B4",X"DA",X"CB",X"ED",X"6D",X"A5",X"F6",X"FC",X"F1",
		X"FF",X"7F",X"7F",X"FF",X"7F",X"97",X"F1",X"87",X"6F",X"3E",X"3C",X"6D",X"A5",X"B6",X"97",X"DB",
		X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"FF",X"CC",X"88",X"00",X"00",X"00",X"00",
		X"8F",X"8F",X"0F",X"8E",X"0E",X"0C",X"08",X"00",X"FF",X"8F",X"0F",X"FF",X"8F",X"8F",X"0F",X"0E",
		X"6F",X"CF",X"6F",X"EF",X"6F",X"CF",X"6F",X"67",X"0F",X"0F",X"0F",X"07",X"07",X"03",X"01",X"00",
		X"00",X"08",X"0C",X"8E",X"8E",X"0F",X"0F",X"8F",X"0E",X"0F",X"7F",X"FF",X"8F",X"7F",X"0F",X"8F",
		X"67",X"CF",X"6F",X"EF",X"6F",X"CF",X"6F",X"EF",X"00",X"01",X"03",X"07",X"07",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"00",X"88",X"CC",X"FF",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"2E",X"26",X"00",X"00",X"00",X"00",X"00",
		X"CE",X"6F",X"7F",X"7F",X"7F",X"2E",X"2E",X"0F",X"1F",X"2F",X"2F",X"0F",X"07",X"07",X"4F",X"0C",
		X"0E",X"0C",X"88",X"CC",X"6E",X"2E",X"4C",X"8C",X"0D",X"4D",X"07",X"27",X"1F",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"08",X"0C",X"8F",X"AE",X"8E",
		X"FC",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F9",X"FF",X"FC",X"F8",X"F0",X"F0",X"F0",X"F0",
		X"8F",X"8F",X"0F",X"9E",X"1E",X"3C",X"78",X"F0",X"FF",X"8F",X"0F",X"FF",X"8F",X"8F",X"0F",X"1E",
		X"6F",X"CF",X"6F",X"EF",X"6F",X"CF",X"6F",X"E7",X"0F",X"0F",X"0F",X"87",X"87",X"C3",X"E1",X"F0",
		X"F0",X"78",X"3C",X"9E",X"9E",X"0F",X"0F",X"8F",X"1E",X"0F",X"7F",X"FF",X"8F",X"7F",X"0F",X"8F",
		X"E7",X"CF",X"6F",X"EF",X"6F",X"CF",X"6F",X"EF",X"F0",X"E1",X"C3",X"87",X"87",X"0F",X"0F",X"0F",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"FC",X"F0",X"F0",X"F0",X"F0",X"F8",X"FC",X"FF",X"F9",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"1E",X"3E",X"B6",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"DE",X"6F",X"7F",X"7F",X"7F",X"3E",X"3E",X"0F",X"1F",X"2F",X"2F",X"0F",X"87",X"87",X"4F",X"3C",
		X"1E",X"3C",X"F8",X"FC",X"7E",X"3E",X"7C",X"BC",X"2D",X"6D",X"87",X"A7",X"1F",X"0F",X"0F",X"0F",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"B4",X"F0",X"F0",X"F0",X"78",X"3C",X"8F",X"BE",X"9E",
		X"F0",X"B4",X"1E",X"1E",X"5A",X"5A",X"F0",X"F0",X"F0",X"D2",X"96",X"B4",X"A5",X"87",X"C3",X"F0",
		X"F0",X"1E",X"F0",X"1E",X"1E",X"F0",X"1E",X"1E",X"87",X"87",X"F0",X"C3",X"87",X"B4",X"87",X"C3",
		X"1E",X"D2",X"1E",X"3C",X"F0",X"1E",X"1E",X"3C",X"87",X"B4",X"87",X"C3",X"F0",X"87",X"87",X"E1",
		X"F0",X"1E",X"1E",X"5A",X"1E",X"96",X"F0",X"3C",X"F0",X"87",X"87",X"B4",X"87",X"87",X"F0",X"C3",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"FF",X"33",X"3D",X"A5",X"42",X"86",X"16",X"92",X"FF",X"FC",X"8B",X"9A",X"A4",X"96",X"06",X"14",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",X"F3",X"FF",X"FF",X"FF",X"3F",X"1F",X"69",X"2D",X"0F",
		X"82",X"06",X"96",X"52",X"85",X"1D",X"F3",X"FF",X"94",X"86",X"16",X"24",X"DA",X"CB",X"CC",X"FF",
		X"F3",X"FB",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"0F",X"0F",X"1F",X"3F",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"50",X"0F",X"20",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"0C",X"0C",X"0E",X"0E",X"0E",X"00",X"0C",X"0F",X"0F",X"0F",X"03",X"01",X"01",
		X"1E",X"0F",X"0F",X"87",X"E0",X"C0",X"C0",X"C0",X"0F",X"0F",X"0F",X"1E",X"1E",X"1E",X"1E",X"1E",
		X"0F",X"0F",X"F0",X"50",X"F0",X"F0",X"F0",X"F0",X"0F",X"00",X"00",X"10",X"20",X"10",X"20",X"50",
		X"00",X"0C",X"0E",X"0E",X"0E",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"80",X"00",X"80",
		X"87",X"0F",X"0F",X"0F",X"0F",X"E0",X"D0",X"E0",X"F0",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"F0",X"70",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"18",X"0F",X"0F",X"0F",
		X"0E",X"0E",X"0E",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"00",X"80",X"80",X"80",X"0C",
		X"0F",X"0F",X"0F",X"F0",X"F0",X"3C",X"0F",X"0F",X"0F",X"0F",X"0F",X"3C",X"0F",X"0F",X"87",X"E1",
		X"E1",X"0F",X"0F",X"0F",X"87",X"61",X"F0",X"F0",X"10",X"01",X"01",X"01",X"00",X"00",X"10",X"18",
		X"0E",X"00",X"00",X"00",X"00",X"00",X"08",X"0E",X"0F",X"00",X"00",X"00",X"00",X"0E",X"0F",X"0F",
		X"0F",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"F0",
		X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"70",X"F0",X"08",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"0E",X"0E",X"80",X"00",X"00",X"0C",X"0F",X"0F",X"0F",X"0F",
		X"F0",X"2C",X"0F",X"0F",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"01",X"00",X"0F",X"0F",X"0F",
		X"07",X"01",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"08",X"0F",X"0F",X"0F",X"0F",
		X"00",X"00",X"08",X"0E",X"0E",X"0E",X"0E",X"00",X"C0",X"0E",X"0F",X"0F",X"0F",X"0F",X"0F",X"C0",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"0F",X"0F",X"0F",X"F0",X"0F",X"0F",X"0F",X"3C",
		X"0F",X"0F",X"10",X"00",X"01",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"01",X"01",X"01",
		X"0E",X"0C",X"0C",X"08",X"80",X"00",X"00",X"00",X"C3",X"0F",X"0F",X"0F",X"0F",X"78",X"00",X"80",
		X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"E0",X"F0",X"70",X"3C",X"0F",X"0F",X"0F",X"87",X"F0",X"0F",
		X"1E",X"0F",X"0F",X"0F",X"03",X"10",X"0F",X"0F",X"07",X"03",X"03",X"00",X"08",X"0F",X"0F",X"0F",
		X"0C",X"0C",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0F",X"C3",X"C3",X"E1",X"E1",X"E1",X"E1",X"E1",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"70",X"F0",X"30",X"B0",X"50",X"B0",X"70",X"B0",
		X"18",X"08",X"00",X"00",X"10",X"00",X"18",X"28",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",
		X"0C",X"00",X"00",X"00",X"80",X"80",X"80",X"08",X"0F",X"0F",X"0C",X"F0",X"78",X"1E",X"0F",X"0F",
		X"C3",X"C3",X"C3",X"3C",X"0F",X"0F",X"0F",X"87",X"B0",X"50",X"F0",X"0F",X"0F",X"0F",X"0F",X"F0",
		X"0F",X"03",X"00",X"03",X"0F",X"0F",X"0F",X"1E",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"07",
		X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0C",X"03",X"01",X"01",X"C1",X"C1",X"C3",X"0F",X"0F",
		X"00",X"00",X"70",X"F0",X"F0",X"70",X"F0",X"43",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",
		X"00",X"00",X"08",X"08",X"0C",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"07",X"07",X"03",X"01",
		X"00",X"00",X"00",X"00",X"08",X"0C",X"0C",X"0E",X"00",X"08",X"0E",X"0F",X"0F",X"0F",X"07",X"03",
		X"0E",X"0F",X"0F",X"0F",X"07",X"01",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",
		X"07",X"0F",X"0F",X"0F",X"0E",X"08",X"08",X"00",X"00",X"01",X"03",X"07",X"07",X"0F",X"0F",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"13",X"13",X"1F",X"1F",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",
		X"00",X"80",X"84",X"0C",X"0C",X"0C",X"0C",X"C0",X"30",X"BC",X"9E",X"8F",X"BC",X"BC",X"AD",X"8F",
		X"1F",X"0F",X"0F",X"07",X"07",X"01",X"00",X"00",X"07",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"80",X"00",X"00",X"CC",X"EE",X"EE",X"00",X"8F",X"AD",X"2D",X"0C",X"0F",X"0F",X"07",X"00",
		X"00",X"00",X"00",X"13",X"13",X"1F",X"1F",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",
		X"00",X"80",X"84",X"0C",X"0C",X"0C",X"0C",X"C0",X"30",X"BC",X"9E",X"8F",X"BC",X"BC",X"AD",X"8F",
		X"1F",X"0F",X"4F",X"EF",X"EF",X"6F",X"0F",X"06",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"8F",X"AD",X"2D",X"08",X"08",X"00",X"00",X"00",
		X"00",X"00",X"01",X"07",X"07",X"0F",X"0F",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",
		X"00",X"EE",X"EE",X"CC",X"00",X"00",X"80",X"84",X"00",X"07",X"0F",X"0F",X"0C",X"3C",X"BC",X"9E",
		X"1F",X"1F",X"1F",X"13",X"13",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"0C",X"0C",X"0C",X"C0",X"C0",X"80",X"00",X"8F",X"BC",X"BC",X"AD",X"8F",X"8F",X"AD",X"21",
		X"06",X"0F",X"6F",X"EF",X"EF",X"4F",X"0F",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"84",X"00",X"00",X"00",X"08",X"08",X"3C",X"BC",X"9E",
		X"1F",X"1F",X"1F",X"13",X"13",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"0C",X"0C",X"0C",X"C0",X"C0",X"80",X"00",X"8F",X"BC",X"BC",X"AD",X"8F",X"8F",X"AD",X"21",
		X"00",X"00",X"0F",X"8F",X"8F",X"87",X"87",X"0F",X"00",X"00",X"00",X"11",X"10",X"30",X"30",X"10",
		X"00",X"00",X"00",X"C0",X"E0",X"69",X"0F",X"C3",X"00",X"00",X"00",X"0B",X"2F",X"6F",X"6F",X"6F",
		X"0F",X"0F",X"0F",X"97",X"B7",X"37",X"03",X"00",X"01",X"34",X"34",X"34",X"34",X"00",X"00",X"00",
		X"C3",X"87",X"3C",X"3C",X"A4",X"84",X"00",X"00",X"6F",X"6F",X"6F",X"6F",X"2F",X"0F",X"08",X"00",
		X"CF",X"CF",X"4F",X"87",X"87",X"87",X"87",X"87",X"00",X"07",X"03",X"21",X"30",X"30",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"84",X"A4",X"3C",X"00",X"08",X"0C",X"0E",X"0E",X"0F",X"0F",X"2F",
		X"87",X"C3",X"C3",X"83",X"67",X"66",X"00",X"00",X"07",X"34",X"34",X"10",X"00",X"00",X"00",X"00",
		X"3C",X"87",X"C3",X"C3",X"0F",X"69",X"E0",X"C0",X"6F",X"0F",X"EF",X"EF",X"EF",X"EF",X"67",X"01",
		X"E1",X"69",X"C3",X"87",X"87",X"0F",X"EF",X"CF",X"03",X"01",X"07",X"34",X"30",X"30",X"30",X"31",
		X"00",X"00",X"00",X"00",X"00",X"84",X"A4",X"3C",X"00",X"00",X"08",X"0C",X"0E",X"0F",X"0F",X"2F",
		X"87",X"07",X"07",X"03",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3C",X"87",X"C3",X"C3",X"07",X"69",X"E0",X"C0",X"6F",X"0F",X"EF",X"EF",X"EF",X"EF",X"67",X"01",
		X"0C",X"86",X"F0",X"E1",X"E1",X"C3",X"C3",X"87",X"01",X"10",X"10",X"00",X"00",X"07",X"34",X"30",
		X"00",X"00",X"00",X"00",X"00",X"84",X"A4",X"3C",X"00",X"00",X"08",X"0C",X"0E",X"0F",X"0F",X"2F",
		X"87",X"C3",X"87",X"0E",X"0C",X"CC",X"88",X"00",X"30",X"10",X"10",X"00",X"11",X"11",X"00",X"00",
		X"3C",X"87",X"C3",X"C3",X"0F",X"69",X"E0",X"C0",X"6F",X"0F",X"EF",X"EF",X"EF",X"EF",X"67",X"01",
		X"00",X"88",X"CC",X"0C",X"0E",X"87",X"C3",X"87",X"00",X"00",X"11",X"11",X"00",X"10",X"10",X"30",
		X"C0",X"E0",X"69",X"0F",X"C3",X"C3",X"87",X"3C",X"01",X"67",X"EF",X"EF",X"EF",X"EF",X"0F",X"6F",
		X"87",X"C3",X"C3",X"E1",X"E1",X"F0",X"86",X"0C",X"30",X"34",X"07",X"00",X"00",X"10",X"10",X"01",
		X"3C",X"A4",X"84",X"00",X"00",X"00",X"00",X"00",X"2F",X"0F",X"0F",X"0E",X"0C",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"0F",X"0F",X"87",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",
		X"C0",X"E0",X"69",X"0F",X"C3",X"C3",X"87",X"3C",X"01",X"67",X"EF",X"EF",X"EF",X"EF",X"0F",X"6F",
		X"CF",X"EF",X"0F",X"87",X"87",X"C3",X"69",X"E0",X"31",X"30",X"30",X"30",X"34",X"07",X"01",X"03",
		X"3C",X"A4",X"84",X"00",X"00",X"00",X"00",X"00",X"2F",X"0F",X"0F",X"0E",X"0C",X"08",X"00",X"00",
		X"00",X"00",X"66",X"67",X"83",X"C3",X"C3",X"87",X"00",X"00",X"00",X"00",X"10",X"30",X"34",X"07",
		X"C0",X"E0",X"69",X"0F",X"C3",X"C3",X"87",X"3C",X"01",X"67",X"EF",X"EF",X"EF",X"EF",X"0F",X"6F",
		X"87",X"87",X"87",X"87",X"C3",X"4F",X"CF",X"CF",X"00",X"10",X"30",X"30",X"21",X"03",X"07",X"00",
		X"3C",X"A4",X"84",X"00",X"00",X"00",X"00",X"00",X"2F",X"0F",X"0F",X"0E",X"0E",X"0C",X"08",X"00",
		X"66",X"EF",X"47",X"83",X"87",X"0F",X"0F",X"0F",X"00",X"07",X"07",X"03",X"43",X"70",X"70",X"61",
		X"00",X"00",X"84",X"A4",X"3C",X"3C",X"87",X"C3",X"00",X"00",X"01",X"2B",X"6F",X"6F",X"0F",X"EF",
		X"0F",X"0F",X"0F",X"0F",X"86",X"C0",X"0C",X"0E",X"21",X"21",X"21",X"10",X"10",X"10",X"01",X"01",
		X"C3",X"0F",X"69",X"E0",X"C0",X"00",X"00",X"00",X"EF",X"EF",X"EF",X"67",X"01",X"00",X"00",X"00",
		X"0E",X"0C",X"C0",X"86",X"0F",X"0F",X"0F",X"0F",X"01",X"01",X"10",X"10",X"10",X"21",X"21",X"21",
		X"00",X"00",X"00",X"C0",X"E0",X"69",X"0F",X"C3",X"00",X"00",X"00",X"01",X"67",X"EF",X"EF",X"EF",
		X"0F",X"0F",X"0F",X"87",X"87",X"47",X"EF",X"66",X"61",X"70",X"70",X"43",X"03",X"07",X"07",X"00",
		X"C3",X"87",X"3C",X"3C",X"A4",X"84",X"00",X"00",X"EF",X"0F",X"6F",X"6F",X"2B",X"01",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"01",X"33",X"33",X"F7",X"A7",X"87",X"0F",X"0F",X"00",X"00",X"04",X"34",X"16",X"34",X"30",X"10",
		X"00",X"00",X"00",X"C0",X"E0",X"69",X"0F",X"C3",X"08",X"0C",X"0C",X"0F",X"2F",X"6F",X"6F",X"6F",
		X"0F",X"0F",X"87",X"87",X"87",X"83",X"00",X"00",X"10",X"10",X"10",X"30",X"34",X"16",X"34",X"04",
		X"C3",X"87",X"3C",X"3C",X"A4",X"B7",X"FF",X"44",X"6F",X"6F",X"6F",X"6F",X"2F",X"0F",X"0F",X"00",
		X"08",X"0E",X"E0",X"78",X"F0",X"C3",X"87",X"0F",X"03",X"34",X"07",X"43",X"70",X"70",X"70",X"30",
		X"00",X"00",X"00",X"00",X"84",X"A4",X"3C",X"3C",X"00",X"00",X"00",X"00",X"01",X"2B",X"6F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"03",X"01",X"00",X"00",X"30",X"01",X"01",X"00",X"00",X"00",X"00",X"00",
		X"87",X"C3",X"C3",X"0F",X"69",X"E0",X"C0",X"00",X"6F",X"6F",X"6F",X"6F",X"2F",X"2F",X"0D",X"EE",
		X"00",X"08",X"C0",X"C2",X"4B",X"0F",X"2F",X"6F",X"07",X"21",X"70",X"70",X"61",X"43",X"07",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"84",X"A4",X"3C",X"3C",
		X"0F",X"6F",X"6F",X"6F",X"EF",X"67",X"01",X"00",X"07",X"07",X"07",X"07",X"47",X"67",X"22",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"87",X"C3",X"C3",X"0F",X"69",X"E0",X"C0",X"00",
		X"00",X"08",X"C0",X"C2",X"4B",X"0F",X"2F",X"6F",X"07",X"21",X"70",X"70",X"61",X"43",X"07",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"84",X"A4",X"3C",X"3C",
		X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"4B",X"61",X"61",X"01",X"01",X"00",X"00",X"00",
		X"00",X"00",X"01",X"03",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"30",
		X"00",X"C0",X"E0",X"69",X"0F",X"C3",X"C3",X"87",X"EE",X"0D",X"2F",X"2F",X"6F",X"6F",X"6F",X"6F",
		X"0F",X"87",X"C3",X"F0",X"78",X"E0",X"0E",X"08",X"30",X"70",X"70",X"70",X"43",X"07",X"34",X"03",
		X"3C",X"3C",X"A4",X"84",X"00",X"00",X"00",X"00",X"0F",X"6F",X"2B",X"01",X"00",X"00",X"00",X"00",
		X"00",X"01",X"67",X"EF",X"6F",X"6F",X"6F",X"0F",X"66",X"22",X"67",X"47",X"07",X"07",X"07",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",X"69",X"0F",X"C3",X"C3",X"87",
		X"6F",X"2F",X"0F",X"4B",X"C3",X"C0",X"08",X"00",X"07",X"07",X"43",X"61",X"70",X"70",X"21",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"3C",X"A4",X"84",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"43",X"43",X"0F",
		X"6F",X"2F",X"0F",X"4B",X"C2",X"C0",X"08",X"00",X"07",X"07",X"43",X"61",X"70",X"70",X"21",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"3C",X"A4",X"84",X"00",X"00",X"00",X"00",
		X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"88",X"7F",X"7F",X"3F",X"0E",X"68",X"C0",X"00",X"BB",
		X"69",X"69",X"4B",X"0F",X"B4",X"F0",X"30",X"22",X"01",X"01",X"01",X"01",X"10",X"00",X"00",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"0E",X"0C",X"08",X"08",X"6E",X"7F",
		X"10",X"10",X"12",X"1E",X"0F",X"2D",X"69",X"69",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",
		X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"88",X"88",X"00",X"00",X"00",X"00",X"6E",X"7F",X"7F",X"7F",X"3F",X"0E",X"68",X"C0",
		X"69",X"69",X"69",X"69",X"4B",X"0F",X"B4",X"F0",X"01",X"01",X"01",X"01",X"01",X"01",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"0E",X"0C",X"08",X"08",
		X"00",X"00",X"10",X"10",X"12",X"1E",X"0F",X"2D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"68",X"C0",X"00",X"CC",X"00",X"00",X"00",X"00",
		X"B4",X"F0",X"30",X"DD",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"88",X"88",X"00",X"00",X"80",X"80",X"6E",X"7F",X"7F",X"7F",X"3F",X"0E",
		X"0F",X"2D",X"69",X"69",X"69",X"69",X"4B",X"0F",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"0E",X"0C",
		X"00",X"00",X"00",X"00",X"10",X"10",X"12",X"1E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"88",X"00",X"00",X"3F",X"0E",X"68",X"C0",X"00",X"DD",X"00",X"00",
		X"4B",X"0F",X"B4",X"F0",X"30",X"AA",X"00",X"00",X"01",X"01",X"10",X"00",X"00",X"11",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"0E",X"0C",X"08",X"08",X"6E",X"7F",X"7F",X"7F",
		X"12",X"1E",X"0F",X"2D",X"69",X"69",X"69",X"69",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"8C",X"A8",X"88",X"20",X"20",X"20",X"00",X"00",X"1F",X"FF",X"F0",X"D0",X"D0",X"A0",X"C0",X"80",
		X"CF",X"CF",X"DF",X"FE",X"FE",X"FC",X"FC",X"FC",X"3B",X"3B",X"3F",X"3B",X"3B",X"1D",X"11",X"00",
		X"00",X"80",X"80",X"20",X"20",X"20",X"88",X"A8",X"EE",X"EF",X"88",X"88",X"EE",X"FF",X"FF",X"3F",
		X"11",X"77",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",X"00",X"00",X"00",X"11",X"11",X"3B",X"3F",X"3B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A8",X"A8",X"8C",X"A8",X"A8",X"00",X"20",X"20",X"FF",X"3F",X"1F",X"FF",X"F0",X"D0",X"D0",X"A0",
		X"FF",X"EF",X"CF",X"CF",X"DF",X"FE",X"FE",X"FC",X"3F",X"3B",X"3B",X"3B",X"3F",X"3B",X"3B",X"1D",
		X"00",X"00",X"80",X"80",X"00",X"20",X"20",X"00",X"00",X"00",X"EE",X"EF",X"88",X"88",X"EE",X"FF",
		X"00",X"00",X"11",X"77",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"3B",
		X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"A0",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"FE",X"FC",X"FC",X"FC",X"00",X"00",X"00",X"00",X"3B",X"1D",X"11",X"00",X"00",X"00",X"00",X"00",
		X"00",X"20",X"A8",X"A8",X"8C",X"A8",X"A8",X"20",X"EE",X"FF",X"FF",X"3F",X"1F",X"FF",X"F0",X"D0",
		X"FF",X"FF",X"FF",X"EF",X"CF",X"CF",X"DF",X"FE",X"11",X"3B",X"3F",X"3B",X"3B",X"3B",X"3F",X"3B",
		X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"20",X"00",X"00",X"00",X"00",X"EE",X"EF",X"88",X"88",
		X"00",X"00",X"00",X"00",X"11",X"77",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",
		X"A8",X"00",X"20",X"20",X"00",X"00",X"00",X"00",X"F0",X"D0",X"D0",X"A0",X"C0",X"80",X"00",X"00",
		X"DF",X"FE",X"FE",X"FC",X"FC",X"FC",X"00",X"00",X"3F",X"3B",X"3B",X"1D",X"11",X"00",X"00",X"00",
		X"00",X"20",X"20",X"00",X"A8",X"A8",X"8C",X"A8",X"88",X"88",X"EE",X"FF",X"FF",X"3F",X"1F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",X"CF",X"CF",X"00",X"11",X"11",X"3B",X"3F",X"3B",X"3B",X"3B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"EF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"44",X"CC",X"88",X"00",X"00",X"00",X"00",X"F7",X"E6",X"4C",X"7F",X"E6",X"08",X"08",X"00",
		X"5A",X"1E",X"C3",X"C3",X"96",X"0F",X"0F",X"07",X"61",X"43",X"03",X"30",X"10",X"01",X"00",X"00",
		X"08",X"C0",X"C0",X"CA",X"CE",X"EE",X"AA",X"AA",X"E1",X"4B",X"3C",X"3F",X"7F",X"7F",X"F7",X"FF",
		X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",X"4F",X"FB",X"16",X"34",X"34",X"34",X"16",X"07",X"34",X"75",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"08",X"08",X"0C",X"A4",X"F0",
		X"B4",X"A5",X"0F",X"6F",X"6F",X"6F",X"EF",X"EF",X"12",X"30",X"30",X"21",X"61",X"61",X"61",X"07",
		X"00",X"00",X"08",X"0C",X"C0",X"80",X"00",X"00",X"00",X"E1",X"C3",X"1E",X"1E",X"3C",X"3C",X"84",
		X"22",X"27",X"2F",X"2F",X"A7",X"A7",X"87",X"1E",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"66",X"44",X"CC",X"88",X"00",X"00",X"F7",X"F7",X"F7",X"E6",X"4C",X"7F",X"E6",X"08",
		X"4F",X"F7",X"5A",X"1E",X"C3",X"C3",X"96",X"0F",X"34",X"73",X"61",X"43",X"03",X"30",X"10",X"01",
		X"00",X"00",X"08",X"C0",X"C0",X"CA",X"CE",X"EE",X"A4",X"F0",X"E1",X"4B",X"3C",X"3F",X"7F",X"7F",
		X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",X"61",X"07",X"16",X"34",X"34",X"34",X"16",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"84",X"80",X"80",X"80",X"08",X"08",X"0C",
		X"87",X"1E",X"B4",X"A5",X"0F",X"6F",X"6F",X"6F",X"10",X"03",X"12",X"30",X"30",X"21",X"61",X"61",
		X"00",X"00",X"00",X"00",X"08",X"0C",X"C0",X"80",X"00",X"00",X"00",X"E1",X"C3",X"1E",X"1E",X"3C",
		X"00",X"00",X"22",X"27",X"2F",X"2F",X"A7",X"A7",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E6",X"08",X"08",X"00",X"00",X"00",X"00",X"00",
		X"96",X"0F",X"0F",X"07",X"00",X"00",X"00",X"00",X"10",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CE",X"EE",X"AA",X"AA",X"66",X"44",X"CC",X"88",X"7F",X"7F",X"F7",X"FF",X"F7",X"E6",X"4C",X"7F",
		X"EF",X"EF",X"4F",X"FE",X"5A",X"1E",X"C3",X"C3",X"16",X"07",X"34",X"76",X"61",X"43",X"03",X"30",
		X"00",X"00",X"00",X"00",X"08",X"C0",X"C0",X"CA",X"08",X"0C",X"A4",X"F0",X"E1",X"4B",X"3C",X"3F",
		X"6F",X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",X"61",X"61",X"61",X"07",X"16",X"34",X"34",X"34",
		X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"1E",X"3C",X"3C",X"84",X"80",X"80",X"80",X"08",
		X"A7",X"A7",X"87",X"1E",X"B4",X"A5",X"0F",X"6F",X"10",X"10",X"10",X"03",X"12",X"30",X"30",X"21",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"0C",X"00",X"00",X"00",X"00",X"00",X"E1",X"C3",X"1E",
		X"00",X"00",X"00",X"00",X"22",X"27",X"2F",X"2F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"4C",X"7F",X"E6",X"08",X"08",X"00",X"00",X"00",
		X"C3",X"C3",X"96",X"0F",X"0F",X"07",X"00",X"00",X"03",X"30",X"10",X"01",X"00",X"00",X"00",X"00",
		X"C0",X"CA",X"CE",X"EE",X"AA",X"AA",X"66",X"44",X"3C",X"3F",X"7F",X"7F",X"F7",X"F7",X"F7",X"E6",
		X"EF",X"EF",X"EF",X"EF",X"4F",X"FB",X"5A",X"1E",X"34",X"34",X"16",X"07",X"34",X"73",X"61",X"43",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"C0",X"80",X"08",X"08",X"0C",X"A4",X"F0",X"E1",X"4B",
		X"0F",X"6F",X"6F",X"EF",X"EF",X"EF",X"EF",X"EF",X"30",X"21",X"61",X"61",X"61",X"07",X"16",X"34",
		X"08",X"0C",X"C0",X"80",X"00",X"00",X"00",X"00",X"C3",X"1E",X"1E",X"3C",X"3C",X"84",X"80",X"80",
		X"2F",X"2F",X"A7",X"A7",X"87",X"1E",X"B4",X"A5",X"00",X"00",X"10",X"10",X"10",X"03",X"12",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E1",
		X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"27",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"02",X"08",X"6E",X"7B",X"F3",X"EE",X"88",X"97",X"F1",X"F3",X"E7",X"CF",X"16",X"32",X"11",
		X"CF",X"7E",X"3D",X"F1",X"E4",X"CD",X"00",X"04",X"03",X"23",X"74",X"FC",X"FE",X"FF",X"77",X"00",
		X"00",X"CC",X"EE",X"F8",X"7B",X"6A",X"4C",X"E6",X"02",X"00",X"DD",X"FC",X"E1",X"79",X"2F",X"4B",
		X"00",X"9B",X"8F",X"2F",X"7C",X"EF",X"4B",X"F7",X"33",X"77",X"FE",X"ED",X"65",X"23",X"09",X"03",
		X"8C",X"C0",X"C0",X"60",X"60",X"30",X"30",X"10",X"7E",X"F3",X"E6",X"C0",X"C1",X"80",X"80",X"80",
		X"CB",X"FD",X"FE",X"FE",X"FF",X"66",X"00",X"00",X"FC",X"30",X"31",X"60",X"40",X"C0",X"81",X"80",
		X"78",X"E6",X"EC",X"80",X"C4",X"EE",X"F7",X"E6",X"1E",X"A5",X"4B",X"0F",X"3D",X"E3",X"C3",X"9F",
		X"6D",X"C3",X"69",X"BC",X"4B",X"CB",X"6D",X"9E",X"E1",X"63",X"31",X"32",X"77",X"FE",X"77",X"FE",
		X"C4",X"EA",X"7F",X"7F",X"EA",X"C4",X"C8",X"68",X"4F",X"A5",X"F5",X"5A",X"69",X"C3",X"F9",X"B4",
		X"D6",X"BD",X"E5",X"0F",X"5A",X"0F",X"DA",X"4B",X"77",X"FE",X"77",X"77",X"36",X"31",X"71",X"F0",
		X"10",X"10",X"30",X"60",X"60",X"C0",X"C9",X"C0",X"00",X"00",X"80",X"A2",X"F7",X"FF",X"FA",X"FD",
		X"10",X"10",X"54",X"FE",X"FC",X"FC",X"F5",X"CB",X"80",X"40",X"60",X"20",X"30",X"14",X"19",X"77",
		X"60",X"30",X"30",X"10",X"00",X"00",X"00",X"00",X"C1",X"80",X"80",X"80",X"00",X"00",X"00",X"00",
		X"FF",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"C0",X"81",X"80",X"00",X"00",X"00",X"00",
		X"C4",X"EE",X"F7",X"E6",X"8C",X"C0",X"C0",X"60",X"3D",X"E3",X"C3",X"9F",X"7E",X"F3",X"E6",X"C0",
		X"4F",X"CB",X"6D",X"9E",X"CB",X"FD",X"FE",X"FE",X"77",X"FE",X"77",X"FE",X"FC",X"30",X"31",X"60",
		X"EA",X"C4",X"C8",X"68",X"78",X"E8",X"E2",X"80",X"69",X"C3",X"F9",X"B4",X"1E",X"A5",X"4B",X"0F",
		X"5A",X"0F",X"DA",X"4B",X"6D",X"C3",X"69",X"BC",X"36",X"31",X"71",X"F0",X"E1",X"63",X"31",X"32",
		X"60",X"C0",X"C9",X"C0",X"C4",X"EA",X"7F",X"7F",X"F7",X"FF",X"FA",X"FD",X"4F",X"A5",X"F5",X"5A",
		X"FC",X"FC",X"F5",X"CB",X"D6",X"BD",X"E5",X"0F",X"30",X"14",X"19",X"77",X"77",X"FE",X"77",X"77",
		X"00",X"00",X"00",X"00",X"10",X"10",X"30",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"A2",
		X"00",X"00",X"00",X"00",X"10",X"10",X"54",X"FE",X"00",X"00",X"00",X"00",X"80",X"40",X"60",X"20",
		X"0E",X"0E",X"0E",X"0C",X"0C",X"08",X"00",X"00",X"81",X"81",X"03",X"0F",X"0F",X"0F",X"0F",X"08",
		X"F0",X"F0",X"E0",X"00",X"0F",X"0F",X"0F",X"0F",X"F0",X"70",X"30",X"0C",X"0F",X"0F",X"0F",X"07",
		X"08",X"08",X"0E",X"0F",X"0F",X"0F",X"03",X"00",X"0F",X"07",X"07",X"03",X"03",X"00",X"00",X"00",
		X"80",X"08",X"0C",X"0E",X"0E",X"0E",X"0E",X"0E",X"0F",X"0F",X"0F",X"C3",X"C3",X"C1",X"C1",X"C1",
		X"0F",X"C3",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"70",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"0F",X"0E",X"08",X"18",X"10",X"10",X"10",X"00",X"07",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0C",X"08",X"00",X"80",X"80",X"80",X"C0",X"80",X"0F",X"0F",X"0F",X"0E",X"78",X"F0",X"78",X"1E",
		X"F0",X"0F",X"0F",X"0F",X"0F",X"3C",X"0F",X"0F",X"78",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"87",X"E1",X"C3",X"0F",X"0F",X"03",X"01",X"10",X"30",X"30",X"10",X"01",X"03",
		X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0C",X"0F",X"01",X"81",X"01",X"01",X"01",X"83",X"43",
		X"E0",X"D0",X"E0",X"D0",X"A0",X"D0",X"A0",X"D0",X"F0",X"F0",X"F0",X"F0",X"E0",X"F0",X"F0",X"F0",
		X"30",X"10",X"30",X"70",X"78",X"78",X"3C",X"1E",X"0F",X"0F",X"0F",X"0F",X"07",X"07",X"07",X"03",
		X"0E",X"0E",X"0E",X"0E",X"00",X"08",X"0E",X"0E",X"0F",X"0F",X"0F",X"01",X"08",X"0F",X"0F",X"0F",
		X"0F",X"07",X"80",X"08",X"0F",X"0F",X"0F",X"0F",X"43",X"D0",X"68",X"0F",X"0F",X"0F",X"0F",X"F0",
		X"10",X"70",X"0F",X"0F",X"0F",X"0F",X"07",X"07",X"08",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"08",X"0F",
		X"0F",X"0F",X"00",X"00",X"00",X"0C",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"0E",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"01",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"01",X"00",
		X"00",X"00",X"08",X"0E",X"0E",X"0E",X"0E",X"0E",X"00",X"08",X"0F",X"0F",X"0F",X"07",X"0F",X"0F",
		X"08",X"0F",X"0F",X"0F",X"07",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"80",X"00",X"00",X"0F",
		X"0F",X"0F",X"0F",X"50",X"20",X"00",X"00",X"00",X"0F",X"0F",X"20",X"10",X"00",X"00",X"00",X"00",
		X"0E",X"0E",X"0E",X"0E",X"0C",X"00",X"00",X"00",X"81",X"81",X"0F",X"0F",X"0F",X"0E",X"80",X"80",
		X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"1E",X"1E",X"0F",X"0F",X"0F",X"0F",X"F0",X"78",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"66",X"EF",X"C7",X"C3",X"87",X"87",X"0F",X"00",X"00",X"00",X"14",X"34",X"16",X"34",X"10",
		X"00",X"00",X"00",X"C0",X"E0",X"69",X"0F",X"C3",X"00",X"00",X"00",X"DB",X"2F",X"6F",X"6F",X"6F",
		X"0F",X"0F",X"87",X"87",X"C3",X"C7",X"EF",X"66",X"10",X"10",X"34",X"16",X"34",X"14",X"00",X"00",
		X"C3",X"87",X"3C",X"3C",X"A4",X"84",X"00",X"00",X"6F",X"6F",X"6F",X"6F",X"2F",X"0B",X"00",X"00",
		X"00",X"00",X"80",X"C3",X"C3",X"C3",X"87",X"87",X"00",X"04",X"16",X"16",X"34",X"30",X"10",X"10",
		X"00",X"44",X"FF",X"F3",X"E0",X"69",X"0F",X"C3",X"00",X"00",X"0F",X"0F",X"2B",X"6F",X"6F",X"6F",
		X"87",X"87",X"87",X"C3",X"C3",X"C1",X"80",X"00",X"10",X"10",X"10",X"30",X"34",X"16",X"16",X"04",
		X"C3",X"87",X"3C",X"3C",X"A4",X"B7",X"FF",X"44",X"6F",X"6F",X"6F",X"6F",X"2B",X"0F",X"0F",X"00",
		X"61",X"E1",X"E1",X"E1",X"0F",X"0F",X"87",X"87",X"00",X"00",X"00",X"00",X"00",X"01",X"10",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"0E",X"0E",X"0E",X"08",X"0C",X"0C",X"1E",X"DE",
		X"87",X"87",X"87",X"0F",X"D2",X"F0",X"30",X"CC",X"70",X"70",X"70",X"01",X"10",X"00",X"00",X"44",
		X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"88",X"EF",X"EF",X"EF",X"0E",X"E0",X"C0",X"00",X"44",
		X"30",X"30",X"30",X"B4",X"B4",X"0F",X"B7",X"B7",X"00",X"00",X"00",X"44",X"10",X"10",X"74",X"30",
		X"00",X"00",X"00",X"C0",X"E0",X"E0",X"2C",X"E0",X"00",X"00",X"80",X"80",X"C0",X"0F",X"8F",X"CF",
		X"B7",X"B7",X"0F",X"B4",X"B4",X"30",X"30",X"30",X"74",X"30",X"10",X"54",X"00",X"00",X"00",X"00",
		X"E0",X"2C",X"E0",X"E0",X"C0",X"00",X"00",X"00",X"CF",X"8F",X"0F",X"C0",X"80",X"80",X"00",X"00",
		X"88",X"30",X"F0",X"D2",X"0F",X"87",X"87",X"87",X"22",X"00",X"00",X"10",X"01",X"70",X"70",X"70",
		X"88",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"99",X"00",X"C0",X"E0",X"0E",X"EF",X"EF",X"EF",
		X"87",X"87",X"0F",X"0F",X"E1",X"E1",X"E1",X"61",X"30",X"10",X"01",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DE",X"1E",X"0C",X"0C",X"08",X"0C",X"0E",X"0E",
		X"40",X"68",X"2C",X"0F",X"0F",X"1F",X"1F",X"0F",X"00",X"01",X"03",X"43",X"43",X"61",X"61",X"01",
		X"00",X"00",X"80",X"C0",X"C0",X"08",X"0C",X"48",X"00",X"00",X"10",X"3C",X"CF",X"EF",X"EF",X"CF",
		X"87",X"C3",X"E1",X"E1",X"C0",X"00",X"00",X"00",X"00",X"10",X"30",X"70",X"30",X"10",X"00",X"00",
		X"C0",X"91",X"80",X"44",X"00",X"00",X"00",X"00",X"0F",X"1E",X"3C",X"78",X"C0",X"11",X"22",X"00",
		X"00",X"00",X"00",X"C0",X"E1",X"E1",X"C3",X"87",X"00",X"00",X"10",X"30",X"70",X"30",X"10",X"00",
		X"00",X"00",X"00",X"88",X"44",X"80",X"91",X"C0",X"44",X"00",X"00",X"C0",X"78",X"3C",X"1E",X"0F",
		X"0F",X"1F",X"1F",X"0F",X"0F",X"2C",X"68",X"40",X"01",X"61",X"61",X"43",X"43",X"03",X"01",X"00",
		X"48",X"0C",X"08",X"C0",X"C0",X"80",X"00",X"00",X"CF",X"EF",X"EF",X"CF",X"3C",X"10",X"00",X"00",
		X"C0",X"E0",X"F0",X"F0",X"E1",X"0F",X"0F",X"0F",X"00",X"00",X"10",X"10",X"00",X"00",X"01",X"01",
		X"80",X"C0",X"86",X"0F",X"0F",X"0F",X"3C",X"28",X"10",X"30",X"30",X"83",X"0F",X"0F",X"0F",X"6F",
		X"1F",X"97",X"C3",X"E1",X"30",X"00",X"44",X"22",X"10",X"10",X"44",X"00",X"11",X"00",X"00",X"00",
		X"08",X"C0",X"E0",X"E0",X"C0",X"80",X"00",X"00",X"EF",X"EF",X"CF",X"1E",X"1C",X"00",X"00",X"00",
		X"22",X"00",X"88",X"30",X"E1",X"C3",X"97",X"1F",X"00",X"00",X"00",X"11",X"00",X"44",X"10",X"10",
		X"00",X"00",X"80",X"C0",X"E0",X"E0",X"C0",X"08",X"00",X"00",X"00",X"1C",X"1E",X"CF",X"EF",X"EF",
		X"0F",X"0F",X"0F",X"E1",X"F0",X"F0",X"E0",X"C0",X"01",X"01",X"00",X"00",X"10",X"10",X"00",X"00",
		X"28",X"3C",X"0F",X"0F",X"0F",X"86",X"C0",X"80",X"6F",X"0F",X"0F",X"0F",X"83",X"30",X"30",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"0E",
		X"01",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"08",X"08",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F1",X"F7",X"FF",X"FF",X"FF",X"FF",X"80",X"00",X"10",X"30",X"22",X"22",X"22",X"22",X"22",
		X"00",X"00",X"C0",X"C0",X"E2",X"E2",X"E2",X"F3",X"80",X"FF",X"FF",X"FE",X"FC",X"FC",X"F8",X"70",
		X"80",X"0C",X"0E",X"1F",X"08",X"34",X"00",X"00",X"22",X"22",X"02",X"01",X"07",X"01",X"01",X"00",
		X"F3",X"F7",X"F7",X"77",X"66",X"C4",X"00",X"00",X"70",X"70",X"70",X"88",X"00",X"F0",X"00",X"00",
		X"00",X"11",X"22",X"44",X"88",X"10",X"60",X"0C",X"00",X"00",X"00",X"00",X"00",X"01",X"05",X"03",
		X"00",X"80",X"C0",X"E0",X"E8",X"FE",X"FF",X"FF",X"E0",X"70",X"30",X"30",X"77",X"FF",X"77",X"33",
		X"0C",X"66",X"11",X"80",X"40",X"20",X"10",X"00",X"03",X"05",X"01",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F1",X"E6",X"EE",X"CC",X"88",X"00",X"30",X"70",X"F0",X"70",X"33",X"33",X"77",X"EE",
		X"00",X"00",X"37",X"08",X"1E",X"0E",X"0C",X"88",X"00",X"01",X"01",X"07",X"01",X"02",X"20",X"20",
		X"00",X"00",X"C8",X"60",X"70",X"F8",X"F8",X"FC",X"00",X"00",X"FF",X"00",X"80",X"77",X"77",X"77",
		X"88",X"F0",X"F0",X"F0",X"F0",X"F8",X"FE",X"FF",X"20",X"20",X"20",X"20",X"20",X"33",X"11",X"00",
		X"FC",X"EC",X"EC",X"EC",X"CC",X"CC",X"00",X"00",X"77",X"F7",X"F3",X"F3",X"F1",X"F0",X"F0",X"88",
		X"00",X"33",X"77",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"15",X"17",X"15",
		X"00",X"48",X"40",X"10",X"10",X"88",X"DC",X"DC",X"FF",X"FF",X"CC",X"CC",X"FF",X"FF",X"FF",X"1F",
		X"EF",X"EF",X"EF",X"FF",X"FF",X"FE",X"FE",X"76",X"15",X"15",X"17",X"15",X"15",X"06",X"00",X"00",
		X"DE",X"DC",X"D4",X"80",X"90",X"10",X"00",X"00",X"0F",X"7F",X"F8",X"E0",X"E0",X"D0",X"E0",X"C0",
		X"00",X"33",X"77",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"15",X"17",X"15",
		X"40",X"48",X"00",X"10",X"00",X"98",X"DC",X"CC",X"FF",X"FF",X"CC",X"CC",X"FF",X"FF",X"FF",X"1F",
		X"EF",X"EF",X"EF",X"FF",X"FF",X"FE",X"FE",X"76",X"15",X"15",X"17",X"15",X"15",X"06",X"00",X"00",
		X"DE",X"CC",X"D4",X"90",X"80",X"10",X"00",X"00",X"0F",X"7F",X"F8",X"E0",X"E0",X"D0",X"E0",X"C0",
		X"00",X"23",X"47",X"7F",X"FF",X"FE",X"FE",X"FE",X"00",X"00",X"00",X"01",X"07",X"00",X"11",X"11",
		X"00",X"00",X"00",X"98",X"98",X"C4",X"D0",X"D2",X"00",X"2E",X"FF",X"F3",X"F0",X"F0",X"F0",X"F0",
		X"FE",X"FE",X"FE",X"FF",X"7F",X"47",X"23",X"00",X"11",X"11",X"00",X"07",X"01",X"00",X"00",X"00",
		X"52",X"50",X"C4",X"98",X"98",X"00",X"00",X"00",X"F0",X"F0",X"E0",X"F0",X"F3",X"FF",X"2E",X"00",
		X"76",X"FE",X"FE",X"FF",X"FF",X"EF",X"EF",X"EF",X"00",X"00",X"06",X"15",X"15",X"17",X"15",X"15",
		X"00",X"00",X"10",X"80",X"90",X"D4",X"CC",X"DE",X"C0",X"E0",X"D0",X"E0",X"E0",X"F8",X"7F",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"77",X"33",X"00",X"15",X"17",X"15",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"DC",X"98",X"00",X"10",X"40",X"48",X"00",X"1F",X"FF",X"FF",X"FF",X"CC",X"CC",X"FF",X"FF",
		X"76",X"FE",X"FE",X"FF",X"FF",X"EF",X"EF",X"EF",X"00",X"00",X"06",X"15",X"15",X"17",X"15",X"15",
		X"00",X"00",X"10",X"90",X"80",X"D4",X"DC",X"CE",X"C0",X"E0",X"D0",X"E0",X"E0",X"F8",X"7F",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"77",X"33",X"00",X"15",X"17",X"15",X"00",X"00",X"00",X"00",X"00",
		X"DC",X"DC",X"88",X"10",X"10",X"00",X"48",X"40",X"1F",X"FF",X"FF",X"FF",X"CC",X"CC",X"FF",X"FF",
		X"00",X"00",X"11",X"77",X"7F",X"FF",X"EF",X"CF",X"00",X"00",X"00",X"01",X"03",X"02",X"06",X"15",
		X"10",X"CE",X"DC",X"88",X"00",X"10",X"98",X"DC",X"00",X"77",X"FF",X"FF",X"FF",X"7F",X"3F",X"1F",
		X"BF",X"FE",X"FC",X"F8",X"F0",X"F0",X"F0",X"30",X"17",X"33",X"37",X"33",X"33",X"11",X"00",X"00",
		X"CC",X"DC",X"CE",X"DC",X"98",X"98",X"00",X"10",X"CF",X"F7",X"F3",X"F1",X"F1",X"B1",X"73",X"C4",
		X"30",X"F0",X"F0",X"F0",X"F8",X"FC",X"FE",X"BF",X"00",X"00",X"11",X"33",X"33",X"37",X"33",X"17",
		X"10",X"10",X"88",X"98",X"DC",X"CE",X"DC",X"DC",X"C4",X"73",X"B1",X"F1",X"F1",X"F3",X"F7",X"CF",
		X"CF",X"EF",X"FF",X"7F",X"77",X"11",X"00",X"00",X"15",X"06",X"02",X"03",X"01",X"00",X"00",X"00",
		X"DC",X"88",X"10",X"00",X"88",X"DC",X"CE",X"10",X"1F",X"3F",X"7F",X"FF",X"FF",X"FF",X"77",X"00",
		X"E8",X"1F",X"DF",X"E3",X"E3",X"CF",X"C3",X"ED",X"11",X"21",X"21",X"57",X"57",X"43",X"43",X"12",
		X"00",X"00",X"00",X"08",X"08",X"8C",X"8D",X"3F",X"00",X"00",X"0E",X"87",X"B7",X"9F",X"8F",X"87",
		X"ED",X"C3",X"CF",X"E3",X"E3",X"DF",X"1F",X"E8",X"56",X"43",X"43",X"57",X"57",X"21",X"21",X"11",
		X"3F",X"1D",X"0C",X"08",X"08",X"00",X"00",X"00",X"87",X"8F",X"8F",X"87",X"87",X"0E",X"00",X"00",
		X"E6",X"1E",X"DE",X"E3",X"E3",X"CF",X"C3",X"ED",X"10",X"23",X"23",X"53",X"53",X"47",X"47",X"52",
		X"00",X"00",X"00",X"08",X"08",X"8C",X"9D",X"3F",X"00",X"00",X"0E",X"8F",X"BF",X"97",X"87",X"8F",
		X"ED",X"C3",X"CF",X"E3",X"E3",X"DE",X"1E",X"E6",X"52",X"47",X"47",X"53",X"53",X"23",X"23",X"10",
		X"3F",X"1D",X"0C",X"08",X"08",X"00",X"00",X"00",X"8F",X"87",X"87",X"8F",X"8F",X"0E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"CC",X"EE",X"FF",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"86",X"00",X"00",X"00",X"00",X"00",X"00",X"25",X"1E",
		X"FF",X"FF",X"EE",X"CC",X"00",X"00",X"00",X"00",X"77",X"77",X"33",X"11",X"00",X"00",X"00",X"00",
		X"78",X"80",X"20",X"00",X"00",X"00",X"00",X"00",X"0F",X"34",X"52",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"CC",X"EE",X"FF",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"68",X"00",X"00",X"00",X"00",X"00",X"00",X"52",X"E1",
		X"FF",X"FF",X"EE",X"CC",X"00",X"00",X"00",X"00",X"77",X"77",X"33",X"11",X"00",X"00",X"00",X"00",
		X"87",X"08",X"02",X"00",X"00",X"00",X"00",X"00",X"F0",X"43",X"25",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"00",X"14",X"5B",X"3E",X"78",X"00",X"00",X"00",X"02",X"01",X"00",X"00",X"50",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"18",X"84",X"CA",
		X"16",X"29",X"10",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B4",X"84",X"02",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"13",X"36",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"0C",X"84",
		X"12",X"01",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"64",X"70",X"F5",X"E1",X"DA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"84",X"C0",X"58",X"F4",X"3D",
		X"C3",X"A5",X"72",X"21",X"22",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B4",X"E8",X"20",X"80",X"00",X"00",X"00",X"00",
		X"80",X"C0",X"42",X"60",X"B4",X"DA",X"87",X"D3",X"00",X"44",X"00",X"01",X"64",X"41",X"30",X"10",
		X"80",X"22",X"00",X"08",X"74",X"C0",X"80",X"00",X"00",X"18",X"30",X"F0",X"7C",X"5A",X"78",X"2C",
		X"0F",X"1E",X"A7",X"C3",X"5A",X"65",X"61",X"90",X"31",X"61",X"10",X"30",X"60",X"50",X"44",X"00",
		X"A4",X"01",X"80",X"E0",X"30",X"08",X"22",X"80",X"87",X"9E",X"3C",X"5A",X"78",X"E0",X"30",X"11",
		X"EE",X"FF",X"99",X"88",X"00",X"77",X"FF",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"11",X"FF",X"EE",X"00",X"EE",X"FF",X"11",
		X"FF",X"77",X"00",X"77",X"FF",X"88",X"FF",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"EE",X"00",X"EE",X"FF",X"11",X"FF",X"EE",
		X"44",X"88",X"FF",X"77",X"00",X"77",X"FF",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"99",X"FF",X"66",X"00",X"EE",X"FF",X"11",
		X"FF",X"77",X"00",X"77",X"FF",X"88",X"FF",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"EE",X"00",X"EE",X"FF",X"11",X"FF",X"EE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
