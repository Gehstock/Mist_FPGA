library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity tcs_rom5 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of tcs_rom5 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"7F",X"82",X"85",X"88",X"8B",X"8F",X"92",X"95",X"98",X"9B",X"9E",X"A1",X"A4",X"A7",X"AA",X"AD",
		X"B0",X"B3",X"B5",X"B8",X"BB",X"BE",X"C0",X"C3",X"C6",X"C8",X"CB",X"CD",X"D0",X"D2",X"D4",X"D7",
		X"D9",X"DB",X"DD",X"DF",X"E1",X"E3",X"E5",X"E7",X"E9",X"EA",X"EC",X"EE",X"EF",X"F0",X"F2",X"F3",
		X"F4",X"F6",X"F7",X"F8",X"F9",X"F9",X"FA",X"FB",X"FC",X"FC",X"FD",X"FD",X"FD",X"FE",X"FE",X"FE",
		X"FE",X"FE",X"FE",X"FE",X"FD",X"FD",X"FD",X"FC",X"FC",X"FB",X"FA",X"F9",X"F9",X"F8",X"F7",X"F5",
		X"F4",X"F3",X"F2",X"F0",X"EF",X"ED",X"EC",X"EA",X"E9",X"E7",X"E5",X"E3",X"E1",X"DF",X"DD",X"DB",
		X"D9",X"D7",X"D4",X"D2",X"D0",X"CD",X"CB",X"C8",X"C6",X"C3",X"C0",X"BE",X"BB",X"B8",X"B5",X"B2",
		X"B0",X"AD",X"AA",X"A7",X"A4",X"A1",X"9E",X"9B",X"98",X"95",X"92",X"8F",X"8B",X"88",X"85",X"82",
		X"7F",X"7C",X"79",X"76",X"73",X"6F",X"6C",X"69",X"66",X"63",X"60",X"5D",X"5A",X"57",X"54",X"51",
		X"4E",X"4C",X"49",X"46",X"43",X"40",X"3E",X"3B",X"38",X"36",X"33",X"31",X"2E",X"2C",X"2A",X"27",
		X"25",X"23",X"21",X"1F",X"1D",X"1B",X"19",X"17",X"15",X"14",X"12",X"10",X"0F",X"0E",X"0C",X"0B",
		X"0A",X"09",X"07",X"06",X"05",X"05",X"04",X"03",X"02",X"02",X"01",X"01",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"02",X"02",X"03",X"04",X"05",X"05",X"06",X"07",X"09",
		X"0A",X"0B",X"0C",X"0E",X"0F",X"11",X"12",X"14",X"15",X"17",X"19",X"1B",X"1D",X"1F",X"21",X"23",
		X"25",X"27",X"2A",X"2C",X"2E",X"31",X"33",X"36",X"38",X"3B",X"3E",X"40",X"43",X"46",X"49",X"4C",
		X"4E",X"51",X"54",X"57",X"5A",X"5D",X"60",X"63",X"66",X"69",X"6C",X"6F",X"73",X"76",X"79",X"7C",
		X"00",X"01",X"02",X"03",X"04",X"05",X"06",X"07",X"08",X"09",X"0A",X"0B",X"0C",X"0D",X"0E",X"0F",
		X"10",X"11",X"12",X"13",X"14",X"15",X"16",X"17",X"18",X"19",X"1A",X"1B",X"1C",X"1D",X"1E",X"1F",
		X"20",X"21",X"22",X"23",X"24",X"25",X"26",X"27",X"28",X"29",X"2A",X"2B",X"2C",X"2D",X"2E",X"2F",
		X"30",X"31",X"32",X"33",X"34",X"35",X"36",X"37",X"38",X"39",X"3A",X"3B",X"3C",X"3D",X"3E",X"3F",
		X"40",X"41",X"42",X"43",X"44",X"45",X"46",X"47",X"48",X"49",X"4A",X"4B",X"4C",X"4D",X"4E",X"4F",
		X"50",X"51",X"52",X"53",X"54",X"55",X"56",X"57",X"58",X"59",X"5A",X"5B",X"5C",X"5D",X"5E",X"5F",
		X"60",X"61",X"62",X"63",X"64",X"65",X"66",X"67",X"68",X"69",X"6A",X"6B",X"6C",X"6D",X"6E",X"6F",
		X"70",X"71",X"72",X"73",X"74",X"75",X"76",X"77",X"78",X"79",X"7A",X"7B",X"7C",X"7D",X"7E",X"7F",
		X"80",X"81",X"82",X"83",X"84",X"85",X"86",X"87",X"88",X"89",X"8A",X"8B",X"8C",X"8D",X"8E",X"8F",
		X"90",X"91",X"92",X"93",X"94",X"95",X"96",X"97",X"98",X"99",X"9A",X"9B",X"9C",X"9D",X"9E",X"9F",
		X"A0",X"A1",X"A2",X"A3",X"A4",X"A5",X"A6",X"A7",X"A8",X"A9",X"AA",X"AB",X"AC",X"AD",X"AE",X"AF",
		X"B0",X"B1",X"B2",X"B3",X"B4",X"B5",X"B6",X"B7",X"B8",X"B9",X"BA",X"BB",X"BC",X"BD",X"BE",X"BF",
		X"C0",X"C1",X"C2",X"C3",X"C4",X"C5",X"C6",X"C7",X"C8",X"C9",X"CA",X"CB",X"CC",X"CD",X"CE",X"CF",
		X"D0",X"D1",X"D2",X"D3",X"D4",X"D5",X"D6",X"D7",X"D8",X"D9",X"DA",X"DB",X"DC",X"DD",X"DE",X"DF",
		X"E0",X"E1",X"E2",X"E3",X"E4",X"E5",X"E6",X"E7",X"E8",X"E9",X"EA",X"EB",X"EC",X"ED",X"EE",X"EF",
		X"F0",X"F1",X"F2",X"F3",X"F4",X"F5",X"F6",X"F7",X"F8",X"F9",X"FA",X"FB",X"FC",X"FD",X"FE",X"FF",
		X"FF",X"FE",X"FD",X"FC",X"FB",X"FA",X"F9",X"F8",X"F7",X"F6",X"F5",X"F4",X"F3",X"F2",X"F1",X"F0",
		X"EF",X"EE",X"ED",X"EC",X"EB",X"EA",X"E9",X"E8",X"E7",X"E6",X"E5",X"E4",X"E3",X"E2",X"E1",X"E0",
		X"DF",X"DE",X"DD",X"DC",X"DB",X"DA",X"D9",X"D8",X"D7",X"D6",X"D5",X"D4",X"D3",X"D2",X"D1",X"D0",
		X"CF",X"CE",X"CD",X"CC",X"CB",X"CA",X"C9",X"C8",X"C7",X"C6",X"C5",X"C4",X"C3",X"C2",X"C1",X"C0",
		X"BF",X"BE",X"BD",X"BC",X"BB",X"BA",X"B9",X"B8",X"B7",X"B6",X"B5",X"B4",X"B3",X"B2",X"B1",X"B0",
		X"AF",X"AE",X"AD",X"AC",X"AB",X"AA",X"A9",X"A8",X"A7",X"A6",X"A5",X"A4",X"A3",X"A2",X"A1",X"A0",
		X"9F",X"9E",X"9D",X"9C",X"9B",X"9A",X"99",X"98",X"97",X"96",X"95",X"94",X"93",X"92",X"91",X"90",
		X"8F",X"8E",X"8D",X"8C",X"8B",X"8A",X"89",X"88",X"87",X"86",X"85",X"84",X"83",X"82",X"81",X"80",
		X"7F",X"7E",X"7D",X"7C",X"7B",X"7A",X"79",X"78",X"77",X"76",X"75",X"74",X"73",X"72",X"71",X"70",
		X"6F",X"6E",X"6D",X"6C",X"6B",X"6A",X"69",X"68",X"67",X"66",X"65",X"64",X"63",X"62",X"61",X"60",
		X"5F",X"5E",X"5D",X"5C",X"5B",X"5A",X"59",X"58",X"57",X"56",X"55",X"54",X"53",X"52",X"51",X"50",
		X"4F",X"4E",X"4D",X"4C",X"4B",X"4A",X"49",X"48",X"47",X"46",X"45",X"44",X"43",X"42",X"41",X"40",
		X"3F",X"3E",X"3D",X"3C",X"3B",X"3A",X"39",X"38",X"37",X"36",X"35",X"34",X"33",X"32",X"31",X"30",
		X"2F",X"2E",X"2D",X"2C",X"2B",X"2A",X"29",X"28",X"27",X"26",X"25",X"24",X"23",X"22",X"21",X"20",
		X"1F",X"1E",X"1D",X"1C",X"1B",X"1A",X"19",X"18",X"17",X"16",X"15",X"14",X"13",X"12",X"11",X"10",
		X"0F",X"0E",X"0D",X"0C",X"0B",X"0A",X"09",X"08",X"07",X"06",X"05",X"04",X"03",X"02",X"01",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",
		X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",X"E7",X"E7",X"E7",X"E7",X"E7",X"E7",X"E7",X"E7",
		X"DF",X"DF",X"DF",X"DF",X"DF",X"DF",X"DF",X"DF",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",
		X"CF",X"CF",X"CF",X"CF",X"CF",X"CF",X"CF",X"CF",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"B7",X"B7",X"B7",X"B7",X"B7",X"B7",X"B7",X"B7",
		X"AF",X"AF",X"AF",X"AF",X"AF",X"AF",X"AF",X"AF",X"A7",X"A7",X"A7",X"A7",X"A7",X"A7",X"A7",X"A7",
		X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"97",X"97",X"97",X"97",X"97",X"97",X"97",X"97",
		X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",
		X"6F",X"6F",X"6F",X"6F",X"6F",X"6F",X"6F",X"6F",X"67",X"67",X"67",X"67",X"67",X"67",X"67",X"67",
		X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"57",X"57",X"57",X"57",X"57",X"57",X"57",X"57",
		X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"4F",X"47",X"47",X"47",X"47",X"47",X"47",X"47",X"47",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"37",
		X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"17",X"17",X"17",X"17",X"17",X"17",X"17",X"17",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",
		X"FF",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",
		X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",
		X"7F",X"85",X"8B",X"92",X"98",X"9E",X"A3",X"A9",X"AF",X"B4",X"BA",X"BF",X"C4",X"C8",X"CC",X"D0",
		X"D4",X"D8",X"DB",X"DE",X"E0",X"E2",X"E4",X"E6",X"E7",X"E8",X"E9",X"E9",X"E9",X"E8",X"E8",X"E7",
		X"E5",X"E4",X"E2",X"E0",X"DD",X"DB",X"D8",X"D5",X"D2",X"CE",X"CB",X"C7",X"C3",X"C0",X"BC",X"B8",
		X"B4",X"B0",X"AC",X"A8",X"A4",X"A0",X"9D",X"99",X"96",X"92",X"8F",X"8C",X"89",X"86",X"84",X"81",
		X"7F",X"7D",X"7B",X"7A",X"78",X"77",X"76",X"76",X"75",X"75",X"75",X"75",X"75",X"76",X"76",X"77",
		X"78",X"79",X"7A",X"7C",X"7D",X"7E",X"80",X"82",X"83",X"85",X"87",X"88",X"8A",X"8C",X"8D",X"8F",
		X"91",X"92",X"93",X"95",X"96",X"97",X"98",X"98",X"99",X"99",X"9A",X"9A",X"9A",X"9A",X"99",X"99",
		X"98",X"98",X"97",X"96",X"94",X"93",X"92",X"90",X"8F",X"8D",X"8B",X"89",X"87",X"85",X"83",X"81",
		X"7F",X"7D",X"7B",X"79",X"77",X"75",X"73",X"71",X"6F",X"6E",X"6C",X"6B",X"6A",X"68",X"67",X"66",
		X"66",X"65",X"65",X"64",X"64",X"64",X"64",X"65",X"65",X"66",X"66",X"67",X"68",X"69",X"6B",X"6C",
		X"6D",X"6F",X"71",X"72",X"74",X"76",X"77",X"79",X"7B",X"7C",X"7E",X"80",X"81",X"82",X"84",X"85",
		X"86",X"87",X"88",X"88",X"89",X"89",X"89",X"89",X"89",X"88",X"88",X"87",X"86",X"85",X"83",X"81",
		X"7F",X"7D",X"7A",X"78",X"75",X"72",X"6F",X"6C",X"68",X"65",X"61",X"5E",X"5A",X"56",X"52",X"4E",
		X"4A",X"46",X"42",X"3E",X"3B",X"37",X"33",X"30",X"2C",X"29",X"26",X"23",X"21",X"1E",X"1C",X"1A",
		X"19",X"17",X"16",X"16",X"15",X"15",X"15",X"16",X"17",X"18",X"1A",X"1C",X"1E",X"20",X"23",X"26",
		X"2A",X"2E",X"32",X"36",X"3A",X"3F",X"44",X"4A",X"4F",X"55",X"5A",X"60",X"66",X"6C",X"73",X"79",
		X"FF",X"00",X"FE",X"01",X"FD",X"02",X"FC",X"03",X"FB",X"04",X"FA",X"05",X"F9",X"06",X"F8",X"07",
		X"F7",X"08",X"F6",X"09",X"F5",X"0A",X"F4",X"0B",X"F3",X"0C",X"F2",X"0D",X"F1",X"0E",X"F0",X"0F",
		X"EF",X"10",X"EE",X"11",X"ED",X"12",X"EC",X"13",X"EB",X"14",X"EA",X"15",X"E9",X"16",X"E8",X"17",
		X"E7",X"18",X"E6",X"19",X"E5",X"1A",X"E4",X"1B",X"E3",X"1C",X"E2",X"1D",X"E1",X"1E",X"E0",X"1F",
		X"DF",X"20",X"DE",X"21",X"DD",X"22",X"DC",X"23",X"DB",X"24",X"DA",X"25",X"D9",X"26",X"D8",X"27",
		X"D7",X"28",X"D6",X"29",X"D5",X"2A",X"D4",X"2B",X"D3",X"2C",X"D2",X"2D",X"D1",X"2E",X"D0",X"2F",
		X"CF",X"30",X"CE",X"31",X"CD",X"32",X"CC",X"33",X"CB",X"34",X"CA",X"35",X"C9",X"36",X"C8",X"37",
		X"C7",X"38",X"C6",X"39",X"C5",X"3A",X"C4",X"3B",X"C3",X"3C",X"C2",X"3D",X"C1",X"3E",X"C0",X"3F",
		X"BF",X"40",X"BE",X"41",X"BD",X"42",X"BC",X"43",X"BB",X"44",X"BA",X"45",X"B9",X"46",X"B8",X"47",
		X"B7",X"48",X"B6",X"49",X"B5",X"4A",X"B4",X"4B",X"B3",X"4C",X"B2",X"4D",X"B1",X"4E",X"B0",X"4F",
		X"AF",X"50",X"AE",X"51",X"AD",X"52",X"AC",X"53",X"AB",X"54",X"AA",X"55",X"A9",X"56",X"A8",X"57",
		X"A7",X"58",X"A6",X"59",X"A5",X"5A",X"A4",X"5B",X"A3",X"5C",X"A2",X"5D",X"A1",X"5E",X"A0",X"5F",
		X"9F",X"60",X"9E",X"61",X"9D",X"62",X"9C",X"63",X"9B",X"64",X"9A",X"65",X"99",X"66",X"98",X"67",
		X"97",X"68",X"96",X"69",X"95",X"6A",X"94",X"6B",X"93",X"6C",X"92",X"6D",X"91",X"6E",X"90",X"6F",
		X"8F",X"70",X"8E",X"71",X"8D",X"72",X"8C",X"73",X"8B",X"74",X"8A",X"75",X"89",X"76",X"88",X"77",
		X"87",X"78",X"86",X"79",X"85",X"7A",X"84",X"7B",X"83",X"7C",X"82",X"7D",X"81",X"7E",X"80",X"7F",
		X"7F",X"80",X"7E",X"81",X"7D",X"82",X"7C",X"83",X"7B",X"84",X"7A",X"85",X"79",X"86",X"78",X"87",
		X"77",X"88",X"76",X"89",X"75",X"8A",X"74",X"8B",X"73",X"8C",X"72",X"8D",X"71",X"8E",X"70",X"8F",
		X"6F",X"90",X"6E",X"91",X"6D",X"92",X"6C",X"93",X"6B",X"94",X"6A",X"95",X"69",X"96",X"68",X"97",
		X"67",X"98",X"66",X"99",X"65",X"9A",X"64",X"9B",X"63",X"9C",X"62",X"9D",X"61",X"9E",X"60",X"9F",
		X"5F",X"A0",X"5E",X"A1",X"5D",X"A2",X"5C",X"A3",X"5B",X"A4",X"5A",X"A5",X"59",X"A6",X"58",X"A7",
		X"57",X"A8",X"56",X"A9",X"55",X"AA",X"54",X"AB",X"53",X"AC",X"52",X"AD",X"51",X"AE",X"50",X"AF",
		X"4F",X"B0",X"4E",X"B1",X"4D",X"B2",X"4C",X"B3",X"4B",X"B4",X"4A",X"B5",X"49",X"B6",X"48",X"B7",
		X"47",X"B8",X"46",X"B9",X"45",X"BA",X"44",X"BB",X"43",X"BC",X"42",X"BD",X"41",X"BE",X"40",X"BF",
		X"3F",X"C0",X"3E",X"C1",X"3D",X"C2",X"3C",X"C3",X"3B",X"C4",X"3A",X"C5",X"39",X"C6",X"38",X"C7",
		X"37",X"C8",X"36",X"C9",X"35",X"CA",X"34",X"CB",X"33",X"CC",X"32",X"CD",X"31",X"CE",X"30",X"CF",
		X"2F",X"D0",X"2E",X"D1",X"2D",X"D2",X"2C",X"D3",X"2B",X"D4",X"2A",X"D5",X"29",X"D6",X"28",X"D7",
		X"27",X"D8",X"26",X"D9",X"25",X"DA",X"24",X"DB",X"23",X"DC",X"22",X"DD",X"21",X"DE",X"20",X"DF",
		X"1F",X"E0",X"1E",X"E1",X"1D",X"E2",X"1C",X"E3",X"1B",X"E4",X"1A",X"E5",X"19",X"E6",X"18",X"E7",
		X"17",X"E8",X"16",X"E9",X"15",X"EA",X"14",X"EB",X"13",X"EC",X"12",X"ED",X"11",X"EE",X"10",X"EF",
		X"0F",X"F0",X"0E",X"F1",X"0D",X"F2",X"0C",X"F3",X"0B",X"F4",X"0A",X"F5",X"09",X"F6",X"08",X"F7",
		X"07",X"F8",X"06",X"F9",X"05",X"FA",X"04",X"FB",X"03",X"FC",X"02",X"FD",X"01",X"FE",X"00",X"FF",
		X"FF",X"FE",X"FD",X"FC",X"00",X"00",X"00",X"00",X"F7",X"F6",X"F5",X"F4",X"00",X"00",X"00",X"00",
		X"EF",X"EE",X"ED",X"EC",X"00",X"00",X"00",X"00",X"E7",X"E6",X"E5",X"E4",X"00",X"00",X"00",X"00",
		X"DF",X"DE",X"DD",X"DC",X"00",X"00",X"00",X"00",X"D7",X"D6",X"D5",X"D4",X"00",X"00",X"00",X"00",
		X"CF",X"CE",X"CD",X"CC",X"00",X"00",X"00",X"00",X"C7",X"C6",X"C5",X"C4",X"00",X"00",X"00",X"00",
		X"BF",X"BE",X"BD",X"BC",X"00",X"00",X"00",X"00",X"B7",X"B6",X"B5",X"B4",X"00",X"00",X"00",X"00",
		X"AF",X"AE",X"AD",X"AC",X"00",X"00",X"00",X"00",X"A7",X"A6",X"A5",X"A4",X"00",X"00",X"00",X"00",
		X"9F",X"9E",X"9D",X"9C",X"00",X"00",X"00",X"00",X"97",X"96",X"95",X"94",X"00",X"00",X"00",X"00",
		X"8F",X"8E",X"8D",X"8C",X"00",X"00",X"00",X"00",X"87",X"86",X"85",X"84",X"00",X"00",X"00",X"00",
		X"7F",X"7E",X"7D",X"7C",X"00",X"00",X"00",X"00",X"77",X"76",X"75",X"74",X"00",X"00",X"00",X"00",
		X"6F",X"6E",X"6D",X"6C",X"00",X"00",X"00",X"00",X"67",X"66",X"65",X"64",X"00",X"00",X"00",X"00",
		X"5F",X"5E",X"5D",X"5C",X"00",X"00",X"00",X"00",X"57",X"56",X"55",X"54",X"00",X"00",X"00",X"00",
		X"4F",X"4E",X"4D",X"4C",X"00",X"00",X"00",X"00",X"47",X"46",X"45",X"44",X"00",X"00",X"00",X"00",
		X"3F",X"3E",X"3D",X"3C",X"00",X"00",X"00",X"00",X"37",X"36",X"35",X"34",X"00",X"00",X"00",X"00",
		X"2F",X"2E",X"2D",X"2C",X"00",X"00",X"00",X"00",X"27",X"26",X"25",X"24",X"00",X"00",X"00",X"00",
		X"1F",X"1E",X"1D",X"1C",X"00",X"00",X"00",X"00",X"17",X"16",X"15",X"14",X"00",X"00",X"00",X"00",
		X"0F",X"0E",X"0D",X"0C",X"00",X"00",X"00",X"00",X"07",X"06",X"05",X"04",X"00",X"00",X"00",X"00",
		X"7E",X"81",X"7C",X"83",X"7A",X"85",X"78",X"87",X"76",X"89",X"74",X"8B",X"72",X"8D",X"70",X"8F",
		X"6E",X"91",X"6C",X"93",X"6A",X"95",X"68",X"97",X"66",X"99",X"64",X"9B",X"62",X"9D",X"60",X"9F",
		X"5E",X"A1",X"5C",X"A3",X"5A",X"A5",X"58",X"A7",X"56",X"A9",X"54",X"AB",X"52",X"AD",X"50",X"AF",
		X"4E",X"B1",X"4C",X"B3",X"4A",X"B5",X"48",X"B7",X"46",X"B9",X"44",X"BB",X"42",X"BD",X"40",X"BF",
		X"3E",X"C1",X"3C",X"C3",X"3A",X"C5",X"38",X"C7",X"36",X"C9",X"34",X"CB",X"32",X"CD",X"30",X"CF",
		X"2E",X"D1",X"2C",X"D3",X"2A",X"D5",X"28",X"D7",X"26",X"D9",X"24",X"DB",X"22",X"DD",X"20",X"DF",
		X"1E",X"E1",X"1C",X"E3",X"1A",X"E5",X"18",X"E7",X"16",X"E9",X"14",X"EB",X"12",X"ED",X"10",X"EF",
		X"0E",X"F1",X"0C",X"F3",X"0A",X"F5",X"08",X"F7",X"06",X"F9",X"04",X"FB",X"02",X"FD",X"00",X"FF",
		X"01",X"FE",X"03",X"FC",X"05",X"FA",X"07",X"F8",X"09",X"F6",X"0B",X"F4",X"0D",X"F2",X"0F",X"F0",
		X"11",X"EE",X"13",X"EC",X"15",X"EA",X"17",X"E8",X"19",X"E6",X"1B",X"E4",X"1D",X"E2",X"1F",X"E0",
		X"21",X"DE",X"23",X"DC",X"25",X"DA",X"27",X"D8",X"29",X"D6",X"2B",X"D4",X"2D",X"D2",X"2F",X"D0",
		X"31",X"CE",X"33",X"CC",X"35",X"CA",X"37",X"C8",X"39",X"C6",X"3B",X"C4",X"3D",X"C2",X"3F",X"C0",
		X"41",X"BE",X"43",X"BC",X"45",X"BA",X"47",X"B8",X"49",X"B6",X"4B",X"B4",X"4D",X"B2",X"4F",X"B0",
		X"51",X"AE",X"53",X"AC",X"55",X"AA",X"57",X"A8",X"59",X"A6",X"5B",X"A4",X"5D",X"A2",X"5F",X"A0",
		X"61",X"9E",X"63",X"9C",X"65",X"9A",X"67",X"98",X"69",X"96",X"6B",X"94",X"6D",X"92",X"6F",X"90",
		X"71",X"8E",X"73",X"8C",X"75",X"8A",X"77",X"88",X"79",X"86",X"7B",X"84",X"7D",X"82",X"7F",X"80",
		X"00",X"FF",X"02",X"FD",X"04",X"FB",X"06",X"F9",X"08",X"F7",X"0A",X"F5",X"0C",X"F3",X"0E",X"F1",
		X"10",X"EF",X"12",X"ED",X"14",X"EB",X"16",X"E9",X"18",X"E7",X"1A",X"E5",X"1C",X"E3",X"1E",X"E1",
		X"20",X"DF",X"22",X"DD",X"24",X"DB",X"26",X"D9",X"28",X"D7",X"2A",X"D5",X"2C",X"D3",X"2E",X"D1",
		X"30",X"CF",X"32",X"CD",X"34",X"CB",X"36",X"C9",X"38",X"C7",X"3A",X"C5",X"3C",X"C3",X"3E",X"C1",
		X"40",X"BF",X"42",X"BD",X"44",X"BB",X"46",X"B9",X"48",X"B7",X"4A",X"B5",X"4C",X"B3",X"4E",X"B1",
		X"50",X"AF",X"52",X"AD",X"54",X"AB",X"56",X"A9",X"58",X"A7",X"5A",X"A5",X"5C",X"A3",X"5E",X"A1",
		X"60",X"9F",X"62",X"9D",X"64",X"9B",X"66",X"99",X"68",X"97",X"6A",X"95",X"6C",X"93",X"6E",X"91",
		X"70",X"8F",X"72",X"8D",X"74",X"8B",X"76",X"89",X"78",X"87",X"7A",X"85",X"7C",X"83",X"7E",X"81",
		X"80",X"7F",X"82",X"7D",X"84",X"7B",X"86",X"79",X"88",X"77",X"8A",X"75",X"8C",X"73",X"8E",X"71",
		X"90",X"6F",X"92",X"6D",X"94",X"6B",X"96",X"69",X"98",X"67",X"9A",X"65",X"9C",X"63",X"9E",X"61",
		X"A0",X"5F",X"A2",X"5D",X"A4",X"5B",X"A6",X"59",X"A8",X"57",X"AA",X"55",X"AC",X"53",X"AE",X"51",
		X"B0",X"4F",X"B2",X"4D",X"B4",X"4B",X"B6",X"49",X"B8",X"47",X"BA",X"45",X"BC",X"43",X"BE",X"41",
		X"C0",X"3F",X"C2",X"3D",X"C4",X"3B",X"C6",X"39",X"C8",X"37",X"CA",X"35",X"CC",X"33",X"CE",X"31",
		X"D0",X"2F",X"D2",X"2D",X"D4",X"2B",X"D6",X"29",X"D8",X"27",X"DA",X"25",X"DC",X"23",X"DE",X"21",
		X"E0",X"1F",X"E2",X"1D",X"E4",X"1B",X"E6",X"19",X"E8",X"17",X"EA",X"15",X"EC",X"13",X"EE",X"11",
		X"F0",X"0F",X"F2",X"0D",X"F4",X"0B",X"F6",X"09",X"F8",X"07",X"FA",X"05",X"FC",X"03",X"FE",X"01",
		X"FF",X"F5",X"EB",X"E2",X"D9",X"D0",X"C8",X"C0",X"B8",X"B1",X"AA",X"A3",X"9C",X"96",X"90",X"8A",
		X"85",X"7F",X"7A",X"75",X"71",X"6C",X"68",X"64",X"60",X"5C",X"58",X"55",X"51",X"68",X"85",X"90",
		X"B8",X"B1",X"AA",X"A3",X"9C",X"96",X"90",X"8A",X"85",X"7F",X"7A",X"75",X"71",X"6C",X"68",X"64",
		X"60",X"5C",X"58",X"55",X"51",X"4E",X"4B",X"48",X"45",X"42",X"40",X"3D",X"3B",X"4B",X"60",X"68",
		X"85",X"7F",X"7A",X"75",X"71",X"6C",X"68",X"64",X"60",X"5C",X"58",X"55",X"51",X"4E",X"4B",X"48",
		X"45",X"42",X"40",X"3D",X"3B",X"38",X"36",X"34",X"32",X"30",X"2E",X"2C",X"2A",X"36",X"45",X"4B",
		X"60",X"5C",X"58",X"55",X"51",X"4E",X"4B",X"48",X"45",X"42",X"40",X"3D",X"3B",X"38",X"36",X"34",
		X"32",X"30",X"2E",X"2C",X"2A",X"29",X"27",X"25",X"24",X"23",X"21",X"20",X"1F",X"27",X"32",X"36",
		X"45",X"42",X"40",X"3D",X"3B",X"38",X"36",X"34",X"32",X"30",X"2E",X"2C",X"2A",X"29",X"27",X"25",
		X"24",X"23",X"21",X"20",X"1F",X"1D",X"1C",X"1B",X"1A",X"19",X"18",X"17",X"16",X"1C",X"24",X"27",
		X"32",X"30",X"2E",X"2C",X"2A",X"29",X"27",X"25",X"24",X"23",X"21",X"20",X"1F",X"1D",X"1C",X"1B",
		X"1A",X"19",X"18",X"17",X"16",X"15",X"14",X"14",X"13",X"12",X"11",X"11",X"10",X"14",X"1A",X"1C",
		X"24",X"23",X"21",X"20",X"1F",X"1D",X"1C",X"1B",X"1A",X"19",X"18",X"17",X"16",X"15",X"14",X"14",
		X"13",X"12",X"11",X"11",X"10",X"0F",X"0F",X"0E",X"0E",X"0D",X"0C",X"0C",X"0B",X"0F",X"13",X"14",
		X"1A",X"19",X"18",X"17",X"16",X"15",X"14",X"14",X"13",X"12",X"11",X"11",X"10",X"0F",X"0F",X"0E",
		X"0E",X"0D",X"0C",X"0C",X"0B",X"0B",X"0B",X"0A",X"09",X"09",X"09",X"08",X"07",X"06",X"05",X"04",
		X"7F",X"DB",X"FE",X"D7",X"7F",X"2A",X"0A",X"2E",X"7F",X"CD",X"EC",X"CA",X"7F",X"37",X"1B",X"39",
		X"7F",X"C2",X"DC",X"BF",X"7F",X"41",X"29",X"43",X"7F",X"B8",X"CE",X"B6",X"7F",X"4A",X"35",X"4C",
		X"7F",X"B0",X"C3",X"AE",X"7F",X"52",X"40",X"53",X"7F",X"A9",X"B9",X"A7",X"7F",X"58",X"49",X"5A",
		X"7F",X"A3",X"B1",X"A1",X"7F",X"5E",X"51",X"5F",X"7F",X"9E",X"AA",X"9C",X"7F",X"63",X"58",X"64",
		X"7F",X"99",X"A3",X"98",X"7F",X"67",X"5D",X"68",X"7F",X"95",X"9E",X"95",X"7F",X"6A",X"62",X"6B",
		X"7F",X"92",X"9A",X"91",X"7F",X"6D",X"66",X"6E",X"7F",X"8F",X"96",X"8F",X"7F",X"70",X"6A",X"70",
		X"7F",X"8D",X"92",X"8D",X"7F",X"72",X"6D",X"73",X"7F",X"8B",X"90",X"8B",X"7F",X"74",X"70",X"74",
		X"7F",X"89",X"8D",X"89",X"7F",X"75",X"72",X"76",X"7F",X"88",X"8B",X"87",X"7F",X"77",X"74",X"77",
		X"7F",X"87",X"89",X"86",X"7F",X"78",X"75",X"78",X"7F",X"85",X"88",X"85",X"7F",X"79",X"77",X"79",
		X"7F",X"84",X"87",X"84",X"7F",X"7A",X"78",X"7A",X"7F",X"84",X"86",X"84",X"7F",X"7B",X"79",X"7B",
		X"7F",X"83",X"85",X"83",X"7F",X"7B",X"7A",X"7B",X"7F",X"82",X"84",X"82",X"7F",X"7C",X"7B",X"7C",
		X"7F",X"82",X"83",X"82",X"7F",X"7C",X"7B",X"7C",X"7F",X"82",X"82",X"81",X"7F",X"7D",X"7C",X"7D",
		X"7F",X"81",X"82",X"81",X"7F",X"7D",X"7C",X"7D",X"7F",X"81",X"82",X"81",X"7F",X"7D",X"7D",X"7D",
		X"7F",X"81",X"81",X"81",X"7F",X"7E",X"7D",X"7E",X"7F",X"80",X"81",X"80",X"7F",X"7E",X"7D",X"7E",
		X"7F",X"80",X"81",X"80",X"7F",X"7E",X"7E",X"7E",X"7F",X"80",X"80",X"80",X"7F",X"7E",X"7E",X"7E",
		X"7F",X"80",X"80",X"80",X"7F",X"7E",X"7E",X"7E",X"7F",X"80",X"80",X"80",X"7F",X"7E",X"7E",X"7E",
		X"FF",X"FA",X"F5",X"F0",X"EC",X"E7",X"E3",X"DE",X"DA",X"D6",X"D2",X"CE",X"CA",X"C6",X"C2",X"BE",
		X"BB",X"B7",X"B3",X"B0",X"AD",X"A9",X"A6",X"A3",X"A0",X"9C",X"99",X"96",X"94",X"91",X"8E",X"8B",
		X"88",X"86",X"83",X"81",X"7E",X"7C",X"79",X"77",X"75",X"72",X"70",X"6E",X"6C",X"6A",X"68",X"66",
		X"64",X"62",X"60",X"5E",X"5C",X"5B",X"59",X"57",X"55",X"54",X"52",X"51",X"4F",X"4D",X"4C",X"4A",
		X"49",X"48",X"46",X"45",X"44",X"42",X"41",X"40",X"3E",X"3D",X"3C",X"3B",X"3A",X"39",X"38",X"37",
		X"35",X"34",X"33",X"32",X"31",X"30",X"30",X"2F",X"2E",X"2D",X"2C",X"2B",X"2A",X"29",X"29",X"28",
		X"27",X"26",X"26",X"25",X"24",X"23",X"23",X"22",X"21",X"21",X"20",X"20",X"1F",X"1E",X"1E",X"1D",
		X"1D",X"1C",X"1C",X"1B",X"1A",X"1A",X"19",X"19",X"18",X"18",X"18",X"17",X"17",X"16",X"16",X"15",
		X"15",X"15",X"14",X"14",X"14",X"13",X"13",X"12",X"12",X"12",X"11",X"11",X"11",X"10",X"10",X"10",
		X"0F",X"0F",X"0F",X"0E",X"0E",X"0E",X"0E",X"0D",X"0D",X"0D",X"0D",X"0C",X"0C",X"0C",X"0C",X"0B",
		X"0B",X"0B",X"0B",X"0B",X"0A",X"0A",X"0A",X"0A",X"0A",X"09",X"09",X"09",X"09",X"09",X"08",X"08",
		X"08",X"08",X"08",X"08",X"08",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"06",X"06",X"06",X"06",
		X"06",X"06",X"06",X"06",X"06",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"04",
		X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"03",X"03",X"03",X"03",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"FE",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",
		X"FD",X"FD",X"FD",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"FC",X"FC",X"FC",X"FC",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",
		X"FB",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"F9",X"F9",X"F9",X"F9",X"F9",
		X"F9",X"F9",X"F9",X"F9",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F7",X"F7",X"F7",X"F7",X"F7",
		X"F7",X"F7",X"F6",X"F6",X"F6",X"F6",X"F6",X"F5",X"F5",X"F5",X"F5",X"F5",X"F4",X"F4",X"F4",X"F4",
		X"F4",X"F3",X"F3",X"F3",X"F3",X"F2",X"F2",X"F2",X"F2",X"F1",X"F1",X"F1",X"F1",X"F0",X"F0",X"F0",
		X"EF",X"EF",X"EF",X"EE",X"EE",X"EE",X"ED",X"ED",X"ED",X"EC",X"EC",X"EB",X"EB",X"EB",X"EA",X"EA",
		X"EA",X"E9",X"E9",X"E8",X"E8",X"E7",X"E7",X"E7",X"E6",X"E6",X"E5",X"E5",X"E4",X"E3",X"E3",X"E2",
		X"E2",X"E1",X"E1",X"E0",X"DF",X"DF",X"DE",X"DE",X"DD",X"DC",X"DC",X"DB",X"DA",X"D9",X"D9",X"D8",
		X"D7",X"D6",X"D6",X"D5",X"D4",X"D3",X"D2",X"D1",X"D0",X"CF",X"CF",X"CE",X"CD",X"CC",X"CB",X"CA",
		X"C8",X"C7",X"C6",X"C5",X"C4",X"C3",X"C2",X"C1",X"BF",X"BE",X"BD",X"BB",X"BA",X"B9",X"B7",X"B6",
		X"B5",X"B3",X"B2",X"B0",X"AE",X"AD",X"AB",X"AA",X"A8",X"A6",X"A4",X"A3",X"A1",X"9F",X"9D",X"9B",
		X"99",X"97",X"95",X"93",X"91",X"8F",X"8D",X"8A",X"88",X"86",X"83",X"81",X"7E",X"7C",X"79",X"77",
		X"74",X"71",X"6E",X"6B",X"69",X"66",X"63",X"5F",X"5C",X"59",X"56",X"52",X"4F",X"4C",X"48",X"44",
		X"41",X"3D",X"39",X"35",X"31",X"2D",X"29",X"25",X"21",X"1C",X"18",X"13",X"0F",X"0A",X"05",X"00",
		X"7F",X"9C",X"B3",X"C6",X"D2",X"D6",X"D2",X"C7",X"BA",X"A8",X"98",X"8C",X"83",X"7F",X"7F",X"82",
		X"86",X"8A",X"8D",X"8C",X"88",X"82",X"79",X"71",X"6B",X"68",X"69",X"6F",X"79",X"87",X"95",X"A2",
		X"AC",X"B1",X"B0",X"AA",X"A0",X"92",X"84",X"78",X"72",X"71",X"77",X"84",X"96",X"AC",X"C1",X"D5",
		X"E3",X"EB",X"EB",X"E3",X"D5",X"C3",X"AF",X"9B",X"8A",X"7D",X"76",X"73",X"74",X"77",X"7B",X"7E",
		X"7F",X"7E",X"7B",X"77",X"74",X"73",X"76",X"7E",X"8A",X"9B",X"AF",X"C3",X"D5",X"E3",X"EB",X"EB",
		X"E3",X"D5",X"C1",X"AC",X"96",X"84",X"77",X"71",X"72",X"78",X"84",X"92",X"9F",X"AA",X"B0",X"B1",
		X"AC",X"A2",X"95",X"87",X"79",X"6F",X"69",X"68",X"6B",X"71",X"79",X"82",X"88",X"8C",X"8D",X"8A",
		X"86",X"82",X"7F",X"7F",X"83",X"8C",X"98",X"A8",X"B9",X"C7",X"D2",X"D6",X"D2",X"C6",X"B3",X"9B",
		X"7F",X"63",X"4B",X"38",X"2C",X"28",X"2C",X"37",X"45",X"56",X"66",X"72",X"7B",X"7F",X"7F",X"7C",
		X"78",X"74",X"71",X"72",X"76",X"7C",X"85",X"8D",X"93",X"96",X"95",X"8F",X"85",X"77",X"69",X"5C",
		X"52",X"4D",X"4E",X"54",X"5F",X"6C",X"7A",X"86",X"8D",X"8D",X"86",X"7A",X"68",X"52",X"3D",X"29",
		X"1B",X"13",X"13",X"1B",X"29",X"3B",X"4F",X"63",X"74",X"80",X"88",X"8B",X"8A",X"87",X"83",X"80",
		X"7F",X"80",X"83",X"87",X"8A",X"8B",X"88",X"80",X"74",X"63",X"4F",X"3B",X"29",X"1B",X"13",X"13",
		X"1B",X"29",X"3D",X"52",X"68",X"7A",X"87",X"8D",X"8C",X"85",X"7A",X"6C",X"5F",X"54",X"4E",X"4D",
		X"52",X"5C",X"69",X"77",X"85",X"8F",X"95",X"96",X"93",X"8D",X"85",X"7C",X"76",X"72",X"71",X"74",
		X"78",X"7C",X"7F",X"7F",X"7B",X"72",X"65",X"56",X"45",X"37",X"2C",X"28",X"2C",X"38",X"4B",X"64",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"FE",X"01",X"FD",X"02",X"FC",X"03",X"FB",X"04",X"FA",X"05",X"F9",X"06",X"F8",X"07",
		X"F7",X"08",X"F6",X"09",X"F5",X"0A",X"F4",X"0B",X"F3",X"0C",X"F2",X"0D",X"F1",X"0E",X"F0",X"0F",
		X"EF",X"10",X"EE",X"11",X"ED",X"12",X"EC",X"13",X"EB",X"14",X"EA",X"15",X"E9",X"16",X"E8",X"17",
		X"E7",X"18",X"E6",X"19",X"E5",X"1A",X"E4",X"1B",X"E3",X"1C",X"E2",X"1D",X"E1",X"1E",X"E0",X"1F",
		X"DF",X"20",X"DE",X"21",X"DD",X"22",X"DC",X"23",X"DB",X"24",X"DA",X"25",X"D9",X"26",X"D8",X"27",
		X"D7",X"28",X"D6",X"29",X"D5",X"2A",X"D4",X"2B",X"D3",X"2C",X"D2",X"2D",X"D1",X"2E",X"D0",X"2F",
		X"CF",X"30",X"CE",X"31",X"CD",X"32",X"CC",X"33",X"CB",X"34",X"CA",X"35",X"C9",X"36",X"C8",X"37",
		X"C0",X"38",X"C6",X"39",X"C5",X"3A",X"C4",X"3B",X"C3",X"3C",X"C2",X"3D",X"C1",X"3E",X"C0",X"3F",
		X"BF",X"40",X"BE",X"41",X"BD",X"42",X"BC",X"43",X"BB",X"44",X"BA",X"45",X"B9",X"46",X"B8",X"47",
		X"B7",X"48",X"B6",X"49",X"B5",X"4A",X"B4",X"4B",X"B3",X"4C",X"B2",X"4D",X"B1",X"4E",X"B0",X"4F",
		X"AF",X"50",X"AE",X"51",X"AD",X"52",X"AC",X"53",X"AB",X"54",X"AA",X"55",X"A9",X"56",X"A8",X"57",
		X"A7",X"58",X"A6",X"59",X"A5",X"5A",X"A4",X"5B",X"A3",X"5C",X"A2",X"5D",X"A1",X"5E",X"A0",X"5F",
		X"9F",X"60",X"9E",X"61",X"9D",X"62",X"9C",X"63",X"9B",X"64",X"9A",X"65",X"99",X"66",X"98",X"67",
		X"97",X"68",X"96",X"69",X"95",X"6A",X"94",X"6B",X"93",X"6C",X"92",X"6D",X"91",X"6E",X"90",X"6F",
		X"8F",X"70",X"8E",X"71",X"8D",X"72",X"8C",X"73",X"8B",X"74",X"8A",X"75",X"89",X"76",X"88",X"77",
		X"87",X"78",X"86",X"79",X"85",X"7A",X"84",X"7B",X"83",X"7C",X"82",X"7D",X"81",X"7E",X"80",X"7F",
		X"FF",X"7F",X"FE",X"7E",X"FD",X"7D",X"FC",X"7C",X"FB",X"7B",X"FA",X"7A",X"F9",X"79",X"F8",X"78",
		X"F7",X"77",X"F6",X"76",X"F5",X"75",X"F4",X"74",X"F3",X"73",X"F2",X"72",X"F1",X"71",X"F0",X"70",
		X"EF",X"6F",X"EE",X"6E",X"ED",X"6D",X"EC",X"6C",X"EB",X"6B",X"EA",X"6A",X"E9",X"69",X"E8",X"68",
		X"E7",X"67",X"E6",X"66",X"E5",X"65",X"E4",X"64",X"E3",X"63",X"E2",X"62",X"E1",X"61",X"E0",X"60",
		X"DF",X"5F",X"DE",X"5E",X"DD",X"5D",X"DC",X"5C",X"DB",X"5B",X"DA",X"5A",X"D9",X"59",X"D8",X"58",
		X"D7",X"57",X"D6",X"56",X"D5",X"55",X"D4",X"54",X"D3",X"53",X"D2",X"52",X"D1",X"51",X"D0",X"50",
		X"CF",X"4F",X"CE",X"4E",X"CD",X"4D",X"CC",X"4C",X"CB",X"4B",X"CA",X"4A",X"C9",X"49",X"C8",X"48",
		X"C7",X"47",X"C6",X"46",X"C5",X"45",X"C4",X"44",X"C3",X"43",X"C2",X"42",X"C1",X"41",X"C0",X"40",
		X"BF",X"3F",X"BE",X"3E",X"BD",X"3D",X"BC",X"3C",X"BB",X"3B",X"BA",X"3A",X"B9",X"39",X"B8",X"38",
		X"B7",X"37",X"B6",X"36",X"B5",X"35",X"B4",X"34",X"B3",X"33",X"B2",X"32",X"B1",X"31",X"B0",X"30",
		X"AF",X"2F",X"AE",X"2E",X"AD",X"2D",X"AC",X"2C",X"AB",X"2B",X"AA",X"2A",X"A9",X"29",X"A8",X"28",
		X"A7",X"27",X"A6",X"26",X"A5",X"25",X"A4",X"24",X"A3",X"23",X"A2",X"22",X"A1",X"21",X"A0",X"20",
		X"9F",X"1F",X"9E",X"1E",X"9D",X"1D",X"9C",X"1C",X"9B",X"1B",X"9A",X"1A",X"99",X"19",X"98",X"18",
		X"97",X"17",X"96",X"16",X"95",X"15",X"94",X"14",X"93",X"13",X"92",X"12",X"91",X"11",X"90",X"10",
		X"8F",X"0F",X"8E",X"0E",X"8D",X"0D",X"8C",X"0C",X"8B",X"0B",X"8A",X"0A",X"89",X"09",X"88",X"08",
		X"87",X"07",X"86",X"06",X"85",X"05",X"84",X"04",X"83",X"03",X"82",X"02",X"81",X"01",X"80",X"00",
		X"7F",X"8D",X"9B",X"A9",X"B6",X"C1",X"CD",X"D7",X"E0",X"E8",X"EF",X"F4",X"F8",X"FC",X"FD",X"FE",
		X"FD",X"FB",X"F8",X"F4",X"EF",X"E9",X"E2",X"DA",X"D1",X"C8",X"BF",X"B4",X"AA",X"9F",X"94",X"8A",
		X"7F",X"75",X"6A",X"61",X"57",X"4F",X"47",X"3F",X"39",X"33",X"2E",X"2A",X"27",X"25",X"23",X"23",
		X"23",X"25",X"27",X"2A",X"2E",X"32",X"37",X"3D",X"43",X"4A",X"51",X"58",X"60",X"68",X"6F",X"77",
		X"7F",X"87",X"8E",X"95",X"9C",X"A2",X"A8",X"AD",X"B2",X"B6",X"BA",X"BD",X"BF",X"C1",X"C2",X"C2",
		X"C2",X"C1",X"BF",X"BD",X"BA",X"B7",X"B3",X"AF",X"AA",X"A6",X"A0",X"9B",X"96",X"90",X"8A",X"85",
		X"7F",X"79",X"74",X"6F",X"6A",X"66",X"61",X"5D",X"5A",X"57",X"54",X"52",X"50",X"4F",X"4F",X"4E",
		X"4F",X"4F",X"50",X"52",X"54",X"56",X"59",X"5C",X"5F",X"63",X"67",X"6B",X"6F",X"73",X"77",X"7B",
		X"7F",X"83",X"87",X"8B",X"8E",X"91",X"95",X"97",X"9A",X"9C",X"9E",X"A0",X"A1",X"A2",X"A2",X"A2",
		X"A2",X"A2",X"A1",X"A0",X"9E",X"9C",X"9B",X"98",X"96",X"93",X"91",X"8E",X"8B",X"88",X"85",X"82",
		X"7F",X"7C",X"79",X"77",X"74",X"72",X"6F",X"6D",X"6B",X"6A",X"68",X"67",X"66",X"66",X"65",X"65",
		X"65",X"66",X"66",X"67",X"68",X"6A",X"6B",X"6D",X"6E",X"70",X"72",X"74",X"76",X"78",X"7B",X"7D",
		X"7F",X"81",X"83",X"85",X"87",X"89",X"8A",X"8C",X"8D",X"8E",X"8F",X"90",X"91",X"91",X"92",X"92",
		X"92",X"91",X"91",X"90",X"8F",X"8F",X"8E",X"8C",X"8B",X"8A",X"88",X"87",X"85",X"84",X"82",X"81",
		X"7F",X"7D",X"7C",X"7B",X"79",X"78",X"77",X"76",X"75",X"74",X"73",X"73",X"72",X"72",X"72",X"71",
		X"72",X"72",X"72",X"73",X"73",X"74",X"74",X"75",X"76",X"77",X"78",X"79",X"7A",X"7C",X"7D",X"7E",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7E",X"7E",X"7E",X"7E",X"7D",X"7D",X"7D",X"7D",X"7D",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7D",X"7D",X"7D",X"7D",X"7E",X"7E",X"7E",X"7F",
		X"7F",X"7F",X"80",X"80",X"81",X"81",X"82",X"82",X"82",X"83",X"83",X"83",X"84",X"84",X"84",X"84",
		X"84",X"85",X"85",X"85",X"84",X"84",X"84",X"84",X"84",X"83",X"83",X"82",X"82",X"81",X"80",X"80",
		X"7F",X"7E",X"7D",X"7D",X"7C",X"7B",X"7A",X"7A",X"79",X"78",X"77",X"77",X"76",X"76",X"75",X"75",
		X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"76",X"77",X"77",X"78",X"79",X"7A",X"7B",X"7C",X"7E",
		X"7F",X"80",X"82",X"83",X"85",X"86",X"88",X"89",X"8B",X"8C",X"8D",X"8E",X"8F",X"90",X"91",X"92",
		X"92",X"92",X"92",X"92",X"92",X"92",X"91",X"90",X"8F",X"8D",X"8C",X"8A",X"88",X"86",X"84",X"82",
		X"7F",X"7C",X"7A",X"77",X"74",X"71",X"6F",X"6C",X"69",X"67",X"65",X"62",X"61",X"5F",X"5D",X"5C",
		X"5B",X"5B",X"5B",X"5B",X"5B",X"5C",X"5E",X"5F",X"62",X"64",X"67",X"6A",X"6E",X"72",X"76",X"7A",
		X"7F",X"84",X"89",X"8E",X"93",X"98",X"9D",X"A2",X"A7",X"AC",X"B0",X"B4",X"B8",X"BB",X"BE",X"C0",
		X"C2",X"C3",X"C3",X"C3",X"C2",X"C0",X"BD",X"BA",X"B6",X"B1",X"AC",X"A6",X"9F",X"98",X"90",X"88",
		X"7F",X"76",X"6D",X"63",X"59",X"50",X"46",X"3D",X"34",X"2B",X"23",X"1B",X"15",X"0F",X"0A",X"05",
		X"02",X"01",X"00",X"01",X"03",X"06",X"0B",X"11",X"18",X"21",X"2B",X"36",X"43",X"50",X"5F",X"6F",
		X"7F",X"8E",X"9C",X"A9",X"B6",X"C0",X"CA",X"D2",X"D8",X"DE",X"E2",X"E6",X"E9",X"EB",X"ED",X"EE",
		X"EF",X"F0",X"F0",X"F0",X"F1",X"F1",X"F0",X"F0",X"F0",X"EF",X"EF",X"EE",X"EE",X"ED",X"EC",X"EB",
		X"EA",X"E9",X"E8",X"E7",X"E6",X"E5",X"E4",X"E3",X"E2",X"E1",X"E0",X"DF",X"DE",X"DD",X"DC",X"DB",
		X"DA",X"D9",X"D7",X"D6",X"D5",X"D4",X"D3",X"D2",X"D1",X"D0",X"CE",X"CD",X"CC",X"CB",X"CA",X"C9",
		X"C8",X"C7",X"C5",X"C4",X"C3",X"C2",X"C1",X"C0",X"BF",X"BD",X"BC",X"BB",X"BA",X"B9",X"B8",X"B7",
		X"B6",X"B4",X"B3",X"B2",X"B1",X"B0",X"AF",X"AE",X"AC",X"AB",X"AA",X"A9",X"A8",X"A7",X"A6",X"A4",
		X"A3",X"A2",X"A1",X"A0",X"9F",X"9E",X"9D",X"9B",X"9A",X"99",X"98",X"97",X"96",X"95",X"93",X"92",
		X"91",X"90",X"8F",X"8E",X"8D",X"8B",X"8A",X"89",X"88",X"87",X"86",X"85",X"84",X"82",X"81",X"80",
		X"7F",X"7E",X"7D",X"7C",X"7A",X"79",X"78",X"77",X"76",X"75",X"74",X"73",X"71",X"70",X"6F",X"6E",
		X"6D",X"6C",X"6B",X"69",X"68",X"67",X"66",X"65",X"64",X"63",X"61",X"60",X"5F",X"5E",X"5D",X"5C",
		X"5B",X"5A",X"58",X"57",X"56",X"55",X"54",X"53",X"52",X"50",X"4F",X"4E",X"4D",X"4C",X"4B",X"4A",
		X"48",X"47",X"46",X"45",X"44",X"43",X"42",X"41",X"3F",X"3E",X"3D",X"3C",X"3B",X"3A",X"39",X"37",
		X"36",X"35",X"34",X"33",X"32",X"31",X"30",X"2E",X"2D",X"2C",X"2B",X"2A",X"29",X"28",X"27",X"25",
		X"24",X"23",X"22",X"21",X"20",X"1F",X"1E",X"1D",X"1C",X"1B",X"1A",X"19",X"18",X"17",X"16",X"15",
		X"14",X"13",X"12",X"11",X"10",X"10",X"0F",X"0F",X"0E",X"0E",X"0E",X"0D",X"0D",X"0E",X"0E",X"0E",
		X"0F",X"10",X"11",X"13",X"15",X"18",X"1C",X"20",X"26",X"2C",X"34",X"3E",X"48",X"55",X"62",X"70",
		X"7F",X"8A",X"94",X"9F",X"A8",X"B1",X"B9",X"C1",X"C8",X"CD",X"D2",X"D7",X"DA",X"DE",X"E0",X"E2",
		X"E4",X"E5",X"E7",X"E7",X"E8",X"E9",X"E9",X"E9",X"E9",X"E9",X"E9",X"E9",X"E9",X"E8",X"E8",X"E7",
		X"E7",X"E6",X"E5",X"E5",X"E4",X"E3",X"E2",X"E2",X"E1",X"E0",X"DF",X"DE",X"DD",X"DC",X"DB",X"DA",
		X"D9",X"D8",X"D7",X"D6",X"D5",X"D4",X"D2",X"D1",X"D0",X"CF",X"CE",X"CD",X"CC",X"CB",X"CA",X"C9",
		X"C7",X"C6",X"C5",X"C4",X"C3",X"C2",X"C1",X"C0",X"BF",X"BD",X"BC",X"BB",X"BA",X"B9",X"B8",X"B7",
		X"B5",X"B4",X"B3",X"B2",X"B1",X"B0",X"AF",X"AE",X"AC",X"AB",X"AA",X"A9",X"A8",X"A7",X"A6",X"A4",
		X"A3",X"A2",X"A1",X"A0",X"9F",X"9E",X"9D",X"9B",X"9A",X"99",X"98",X"97",X"96",X"95",X"93",X"92",
		X"91",X"90",X"8F",X"8E",X"8D",X"8B",X"8A",X"89",X"88",X"87",X"86",X"85",X"84",X"82",X"81",X"80",
		X"7F",X"7E",X"7D",X"7C",X"7A",X"79",X"78",X"77",X"76",X"75",X"74",X"73",X"71",X"70",X"6F",X"6E",
		X"6D",X"6C",X"6B",X"69",X"68",X"67",X"66",X"65",X"64",X"63",X"61",X"60",X"5F",X"5E",X"5D",X"5C",
		X"5B",X"5A",X"58",X"57",X"56",X"55",X"54",X"53",X"52",X"50",X"4F",X"4E",X"4D",X"4C",X"4B",X"4A",
		X"49",X"47",X"46",X"45",X"44",X"43",X"42",X"41",X"3F",X"3E",X"3D",X"3C",X"3B",X"3A",X"39",X"38",
		X"37",X"35",X"34",X"33",X"32",X"31",X"30",X"2F",X"2E",X"2D",X"2C",X"2A",X"29",X"28",X"27",X"26",
		X"25",X"24",X"23",X"22",X"21",X"20",X"1F",X"1E",X"1D",X"1C",X"1C",X"1B",X"1A",X"19",X"19",X"18",
		X"17",X"17",X"16",X"16",X"15",X"15",X"15",X"15",X"15",X"15",X"15",X"15",X"16",X"17",X"17",X"19",
		X"1A",X"1C",X"1E",X"20",X"24",X"27",X"2C",X"31",X"36",X"3D",X"45",X"4D",X"56",X"5F",X"6A",X"74",
		X"7F",X"86",X"8D",X"93",X"9A",X"A0",X"A6",X"AC",X"B1",X"B6",X"BB",X"BF",X"C3",X"C7",X"CA",X"CD",
		X"CF",X"D2",X"D4",X"D5",X"D7",X"D8",X"D9",X"DA",X"DB",X"DC",X"DC",X"DC",X"DD",X"DD",X"DD",X"DD",
		X"DD",X"DC",X"DC",X"DC",X"DC",X"DB",X"DB",X"DA",X"DA",X"D9",X"D9",X"D8",X"D7",X"D7",X"D6",X"D5",
		X"D5",X"D4",X"D3",X"D2",X"D1",X"D0",X"D0",X"CF",X"CE",X"CD",X"CC",X"CB",X"CA",X"C9",X"C8",X"C7",
		X"C6",X"C5",X"C4",X"C3",X"C2",X"C1",X"C0",X"BF",X"BE",X"BD",X"BB",X"BA",X"B9",X"B8",X"B7",X"B6",
		X"B5",X"B4",X"B3",X"B2",X"B1",X"AF",X"AE",X"AD",X"AC",X"AB",X"AA",X"A9",X"A8",X"A7",X"A5",X"A4",
		X"A3",X"A2",X"A1",X"A0",X"9F",X"9E",X"9C",X"9B",X"9A",X"99",X"98",X"97",X"96",X"95",X"93",X"92",
		X"91",X"90",X"8F",X"8E",X"8D",X"8B",X"8A",X"89",X"88",X"87",X"86",X"85",X"84",X"82",X"81",X"80",
		X"7F",X"7E",X"7D",X"7C",X"7A",X"79",X"78",X"77",X"76",X"75",X"74",X"73",X"71",X"70",X"6F",X"6E",
		X"6D",X"6C",X"6B",X"69",X"68",X"67",X"66",X"65",X"64",X"63",X"62",X"60",X"5F",X"5E",X"5D",X"5C",
		X"5B",X"5A",X"59",X"57",X"56",X"55",X"54",X"53",X"52",X"51",X"50",X"4F",X"4D",X"4C",X"4B",X"4A",
		X"49",X"48",X"47",X"46",X"45",X"44",X"43",X"41",X"40",X"3F",X"3E",X"3D",X"3C",X"3B",X"3A",X"39",
		X"38",X"37",X"36",X"35",X"34",X"33",X"32",X"31",X"30",X"2F",X"2E",X"2E",X"2D",X"2C",X"2B",X"2A",
		X"29",X"29",X"28",X"27",X"27",X"26",X"25",X"25",X"24",X"24",X"23",X"23",X"22",X"22",X"22",X"22",
		X"21",X"21",X"21",X"21",X"21",X"22",X"22",X"22",X"23",X"24",X"25",X"26",X"27",X"29",X"2A",X"2C",
		X"2F",X"31",X"34",X"37",X"3B",X"3F",X"43",X"48",X"4D",X"52",X"58",X"5E",X"64",X"6B",X"71",X"78",
		X"7F",X"84",X"89",X"8D",X"92",X"97",X"9B",X"A0",X"A4",X"A8",X"AC",X"AF",X"B3",X"B6",X"B9",X"BC",
		X"BE",X"C1",X"C3",X"C5",X"C7",X"C9",X"CA",X"CC",X"CD",X"CE",X"CF",X"D0",X"D0",X"D1",X"D1",X"D2",
		X"D2",X"D2",X"D2",X"D2",X"D2",X"D2",X"D2",X"D2",X"D1",X"D1",X"D1",X"D0",X"D0",X"D0",X"CF",X"CF",
		X"CE",X"CD",X"CD",X"CC",X"CC",X"CB",X"CA",X"CA",X"C9",X"C8",X"C7",X"C7",X"C6",X"C5",X"C4",X"C3",
		X"C2",X"C2",X"C1",X"C0",X"BF",X"BE",X"BD",X"BC",X"BB",X"BA",X"B9",X"B8",X"B7",X"B6",X"B5",X"B4",
		X"B3",X"B2",X"B1",X"B0",X"AF",X"AE",X"AD",X"AC",X"AB",X"AA",X"A9",X"A8",X"A7",X"A6",X"A5",X"A3",
		X"A2",X"A1",X"A0",X"9F",X"9E",X"9D",X"9C",X"9B",X"9A",X"99",X"97",X"96",X"95",X"94",X"93",X"92",
		X"91",X"90",X"8F",X"8D",X"8C",X"8B",X"8A",X"89",X"88",X"87",X"86",X"85",X"83",X"82",X"81",X"80",
		X"7F",X"7E",X"7D",X"7C",X"7B",X"79",X"78",X"77",X"76",X"75",X"74",X"73",X"72",X"71",X"6F",X"6E",
		X"6D",X"6C",X"6B",X"6A",X"69",X"68",X"67",X"65",X"64",X"63",X"62",X"61",X"60",X"5F",X"5E",X"5D",
		X"5C",X"5B",X"59",X"58",X"57",X"56",X"55",X"54",X"53",X"52",X"51",X"50",X"4F",X"4E",X"4D",X"4C",
		X"4B",X"4A",X"49",X"48",X"47",X"46",X"45",X"44",X"43",X"42",X"41",X"40",X"3F",X"3E",X"3D",X"3C",
		X"3C",X"3B",X"3A",X"39",X"38",X"37",X"37",X"36",X"35",X"34",X"34",X"33",X"32",X"32",X"31",X"31",
		X"30",X"2F",X"2F",X"2E",X"2E",X"2E",X"2D",X"2D",X"2D",X"2C",X"2C",X"2C",X"2C",X"2C",X"2C",X"2C",
		X"2C",X"2C",X"2D",X"2D",X"2E",X"2E",X"2F",X"30",X"31",X"32",X"34",X"35",X"37",X"39",X"3B",X"3D",
		X"40",X"42",X"45",X"48",X"4B",X"4F",X"52",X"56",X"5A",X"5E",X"63",X"67",X"6C",X"71",X"75",X"7A",
		X"7F",X"82",X"85",X"88",X"8A",X"8D",X"90",X"93",X"95",X"98",X"9A",X"9D",X"9F",X"A2",X"A4",X"A6",
		X"A8",X"AA",X"AC",X"AE",X"AF",X"B1",X"B3",X"B4",X"B5",X"B7",X"B8",X"B9",X"BA",X"BB",X"BC",X"BD",
		X"BD",X"BE",X"BE",X"BF",X"BF",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"C0",X"C0",X"BF",X"BF",X"BF",X"BE",X"BE",X"BD",X"BD",X"BC",X"BC",X"BB",X"BB",X"BA",X"BA",X"B9",
		X"B8",X"B8",X"B7",X"B7",X"B6",X"B5",X"B4",X"B4",X"B3",X"B2",X"B1",X"B1",X"B0",X"AF",X"AE",X"AE",
		X"AD",X"AC",X"AB",X"AA",X"A9",X"A9",X"A8",X"A7",X"A6",X"A5",X"A4",X"A3",X"A2",X"A1",X"A0",X"A0",
		X"9F",X"9E",X"9D",X"9C",X"9B",X"9A",X"99",X"98",X"97",X"96",X"95",X"94",X"93",X"92",X"91",X"90",
		X"8F",X"8E",X"8D",X"8C",X"8B",X"8A",X"89",X"88",X"87",X"86",X"85",X"84",X"83",X"82",X"81",X"80",
		X"7F",X"7E",X"7D",X"7C",X"7B",X"7A",X"79",X"78",X"77",X"76",X"75",X"74",X"73",X"72",X"71",X"70",
		X"6F",X"6E",X"6D",X"6C",X"6B",X"6A",X"69",X"68",X"67",X"66",X"65",X"64",X"63",X"62",X"61",X"60",
		X"5F",X"5E",X"5E",X"5D",X"5C",X"5B",X"5A",X"59",X"58",X"57",X"56",X"55",X"55",X"54",X"53",X"52",
		X"51",X"50",X"50",X"4F",X"4E",X"4D",X"4D",X"4C",X"4B",X"4A",X"4A",X"49",X"48",X"47",X"47",X"46",
		X"46",X"45",X"44",X"44",X"43",X"43",X"42",X"42",X"41",X"41",X"40",X"40",X"3F",X"3F",X"3F",X"3E",
		X"3E",X"3E",X"3E",X"3E",X"3E",X"3E",X"3E",X"3E",X"3E",X"3E",X"3E",X"3E",X"3F",X"3F",X"40",X"40",
		X"41",X"41",X"42",X"43",X"44",X"45",X"46",X"47",X"49",X"4A",X"4B",X"4D",X"4F",X"50",X"52",X"54",
		X"56",X"58",X"5A",X"5C",X"5F",X"61",X"64",X"66",X"69",X"6B",X"6E",X"71",X"74",X"76",X"79",X"7C",
		X"7F",X"81",X"83",X"85",X"86",X"88",X"8A",X"8C",X"8E",X"8F",X"91",X"93",X"95",X"96",X"98",X"99",
		X"9B",X"9C",X"9E",X"9F",X"A0",X"A2",X"A3",X"A4",X"A5",X"A6",X"A7",X"A8",X"A9",X"AA",X"AB",X"AC",
		X"AD",X"AD",X"AE",X"AF",X"AF",X"B0",X"B0",X"B0",X"B1",X"B1",X"B1",X"B2",X"B2",X"B2",X"B2",X"B2",
		X"B2",X"B2",X"B2",X"B2",X"B2",X"B2",X"B2",X"B1",X"B1",X"B1",X"B1",X"B0",X"B0",X"B0",X"AF",X"AF",
		X"AF",X"AE",X"AE",X"AD",X"AD",X"AC",X"AC",X"AB",X"AA",X"AA",X"A9",X"A9",X"A8",X"A7",X"A7",X"A6",
		X"A6",X"A5",X"A4",X"A3",X"A3",X"A2",X"A1",X"A1",X"A0",X"9F",X"9E",X"9E",X"9D",X"9C",X"9B",X"9B",
		X"9A",X"99",X"98",X"97",X"97",X"96",X"95",X"94",X"93",X"93",X"92",X"91",X"90",X"8F",X"8E",X"8E",
		X"8D",X"8C",X"8B",X"8A",X"89",X"88",X"88",X"87",X"86",X"85",X"84",X"83",X"82",X"82",X"81",X"80",
		X"7F",X"7E",X"7D",X"7C",X"7C",X"7B",X"7A",X"79",X"78",X"77",X"76",X"76",X"75",X"74",X"73",X"72",
		X"71",X"70",X"70",X"6F",X"6E",X"6D",X"6C",X"6B",X"6B",X"6A",X"69",X"68",X"67",X"67",X"66",X"65",
		X"64",X"63",X"63",X"62",X"61",X"60",X"60",X"5F",X"5E",X"5D",X"5D",X"5C",X"5B",X"5B",X"5A",X"59",
		X"58",X"58",X"57",X"57",X"56",X"55",X"55",X"54",X"54",X"53",X"52",X"52",X"51",X"51",X"50",X"50",
		X"4F",X"4F",X"4F",X"4E",X"4E",X"4E",X"4D",X"4D",X"4D",X"4D",X"4C",X"4C",X"4C",X"4C",X"4C",X"4C",
		X"4C",X"4C",X"4C",X"4C",X"4C",X"4C",X"4D",X"4D",X"4D",X"4E",X"4E",X"4E",X"4F",X"4F",X"50",X"51",
		X"51",X"52",X"53",X"54",X"55",X"56",X"57",X"58",X"59",X"5A",X"5B",X"5C",X"5E",X"5F",X"60",X"62",
		X"63",X"65",X"66",X"68",X"69",X"6B",X"6D",X"6F",X"70",X"72",X"74",X"76",X"78",X"79",X"7B",X"7D",
		X"7F",X"80",X"81",X"82",X"83",X"84",X"84",X"85",X"86",X"87",X"88",X"89",X"8A",X"8B",X"8B",X"8C",
		X"8D",X"8E",X"8F",X"8F",X"90",X"91",X"92",X"92",X"93",X"94",X"94",X"95",X"96",X"96",X"97",X"97",
		X"98",X"98",X"99",X"99",X"9A",X"9A",X"9B",X"9B",X"9B",X"9C",X"9C",X"9C",X"9D",X"9D",X"9D",X"9D",
		X"9D",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",
		X"9E",X"9D",X"9D",X"9D",X"9D",X"9D",X"9C",X"9C",X"9C",X"9C",X"9B",X"9B",X"9B",X"9A",X"9A",X"9A",
		X"99",X"99",X"99",X"98",X"98",X"97",X"97",X"96",X"96",X"96",X"95",X"95",X"94",X"94",X"93",X"93",
		X"92",X"92",X"91",X"90",X"90",X"8F",X"8F",X"8E",X"8E",X"8D",X"8D",X"8C",X"8B",X"8B",X"8A",X"8A",
		X"89",X"88",X"88",X"87",X"87",X"86",X"85",X"85",X"84",X"83",X"83",X"82",X"82",X"81",X"80",X"80",
		X"7F",X"7E",X"7E",X"7D",X"7C",X"7C",X"7B",X"7B",X"7A",X"79",X"79",X"78",X"77",X"77",X"76",X"76",
		X"75",X"74",X"74",X"73",X"73",X"72",X"71",X"71",X"70",X"70",X"6F",X"6F",X"6E",X"6E",X"6D",X"6C",
		X"6C",X"6B",X"6B",X"6A",X"6A",X"69",X"69",X"68",X"68",X"68",X"67",X"67",X"66",X"66",X"65",X"65",
		X"65",X"64",X"64",X"64",X"63",X"63",X"63",X"62",X"62",X"62",X"62",X"61",X"61",X"61",X"61",X"61",
		X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",
		X"61",X"61",X"61",X"61",X"61",X"62",X"62",X"62",X"63",X"63",X"63",X"64",X"64",X"65",X"65",X"66",
		X"66",X"67",X"67",X"68",X"68",X"69",X"6A",X"6A",X"6B",X"6C",X"6C",X"6D",X"6E",X"6F",X"6F",X"70",
		X"71",X"72",X"73",X"73",X"74",X"75",X"76",X"77",X"78",X"79",X"7A",X"7A",X"7B",X"7C",X"7D",X"7E",
		X"7F",X"80",X"80",X"81",X"81",X"82",X"82",X"82",X"83",X"83",X"84",X"84",X"85",X"85",X"86",X"86",
		X"87",X"87",X"88",X"88",X"89",X"89",X"89",X"8A",X"8A",X"8B",X"8B",X"8B",X"8C",X"8C",X"8C",X"8D",
		X"8D",X"8D",X"8E",X"8E",X"8E",X"8F",X"8F",X"8F",X"8F",X"90",X"90",X"90",X"90",X"90",X"91",X"91",
		X"91",X"91",X"91",X"91",X"91",X"92",X"92",X"92",X"92",X"92",X"92",X"92",X"92",X"92",X"92",X"92",
		X"92",X"92",X"92",X"92",X"92",X"92",X"91",X"91",X"91",X"91",X"91",X"91",X"91",X"90",X"90",X"90",
		X"90",X"90",X"90",X"8F",X"8F",X"8F",X"8F",X"8E",X"8E",X"8E",X"8D",X"8D",X"8D",X"8D",X"8C",X"8C",
		X"8C",X"8B",X"8B",X"8B",X"8A",X"8A",X"8A",X"89",X"89",X"88",X"88",X"88",X"87",X"87",X"87",X"86",
		X"86",X"85",X"85",X"85",X"84",X"84",X"83",X"83",X"82",X"82",X"82",X"81",X"81",X"80",X"80",X"7F",
		X"7F",X"7F",X"7E",X"7E",X"7D",X"7D",X"7C",X"7C",X"7C",X"7B",X"7B",X"7A",X"7A",X"79",X"79",X"79",
		X"78",X"78",X"77",X"77",X"77",X"76",X"76",X"76",X"75",X"75",X"74",X"74",X"74",X"73",X"73",X"73",
		X"72",X"72",X"72",X"71",X"71",X"71",X"71",X"70",X"70",X"70",X"6F",X"6F",X"6F",X"6F",X"6E",X"6E",
		X"6E",X"6E",X"6E",X"6E",X"6D",X"6D",X"6D",X"6D",X"6D",X"6D",X"6D",X"6C",X"6C",X"6C",X"6C",X"6C",
		X"6C",X"6C",X"6C",X"6C",X"6C",X"6C",X"6C",X"6C",X"6C",X"6C",X"6C",X"6C",X"6D",X"6D",X"6D",X"6D",
		X"6D",X"6D",X"6D",X"6E",X"6E",X"6E",X"6E",X"6E",X"6F",X"6F",X"6F",X"6F",X"70",X"70",X"70",X"71",
		X"71",X"71",X"72",X"72",X"72",X"73",X"73",X"73",X"74",X"74",X"75",X"75",X"75",X"76",X"76",X"77",
		X"77",X"78",X"78",X"79",X"79",X"7A",X"7A",X"7B",X"7B",X"7C",X"7C",X"7C",X"7D",X"7D",X"7E",X"7E",
		X"43",X"4F",X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"20",X"31",X"39",X"38",X"35",X"2C",X"20",
		X"42",X"41",X"4C",X"4C",X"59",X"20",X"4D",X"49",X"44",X"57",X"41",X"59",X"20",X"4D",X"46",X"47",
		X"2E",X"20",X"43",X"4F",X"2E",X"20",X"20",X"41",X"4C",X"4C",X"20",X"52",X"49",X"47",X"48",X"54",
		X"53",X"20",X"52",X"45",X"53",X"45",X"52",X"56",X"45",X"44",X"4E",X"41",X"35",X"39",X"2D",X"30",
		X"58",X"58",X"2D",X"55",X"35",X"20",X"20",X"00",X"00",X"FF",X"0D",X"01",X"10",X"26",X"01",X"57",
		X"DC",X"2D",X"D3",X"2F",X"DD",X"2D",X"DC",X"25",X"D3",X"27",X"DD",X"25",X"A6",X"9F",X"00",X"2C",
		X"E6",X"9F",X"00",X"24",X"3D",X"D3",X"1D",X"D3",X"1F",X"DD",X"1D",X"A6",X"9F",X"00",X"1C",X"D6",
		X"3A",X"3D",X"97",X"22",X"DC",X"4D",X"D3",X"4F",X"DD",X"4D",X"DC",X"45",X"D3",X"47",X"DD",X"45",
		X"A6",X"9F",X"00",X"4C",X"E6",X"9F",X"00",X"44",X"3D",X"D3",X"3D",X"D3",X"3F",X"DD",X"3D",X"A6",
		X"9F",X"00",X"3C",X"D6",X"5A",X"3D",X"97",X"42",X"DC",X"65",X"D3",X"67",X"DD",X"65",X"DC",X"5D",
		X"D3",X"5F",X"AB",X"9F",X"00",X"64",X"DD",X"5D",X"A6",X"9F",X"00",X"5C",X"D6",X"7A",X"3D",X"97",
		X"62",X"DC",X"85",X"D3",X"87",X"DD",X"85",X"DC",X"7D",X"D3",X"7F",X"AB",X"9F",X"00",X"84",X"DD",
		X"7D",X"A6",X"9F",X"00",X"7C",X"D6",X"9A",X"3D",X"97",X"82",X"DC",X"A5",X"D3",X"A7",X"DD",X"A5",
		X"DC",X"9D",X"D3",X"9F",X"AB",X"9F",X"00",X"A4",X"DD",X"9D",X"A6",X"9F",X"00",X"9C",X"D6",X"BA",
		X"3D",X"9B",X"82",X"46",X"D6",X"22",X"DB",X"42",X"56",X"DB",X"62",X"56",X"34",X"04",X"5F",X"AB",
		X"E0",X"46",X"56",X"FD",X"60",X"00",X"8E",X"E0",X"D8",X"96",X"00",X"48",X"48",X"10",X"AE",X"86",
		X"8B",X"02",X"EE",X"86",X"EC",X"C4",X"E3",X"42",X"ED",X"C4",X"A6",X"D8",X"FF",X"A7",X"45",X"EC",
		X"A4",X"83",X"00",X"01",X"ED",X"A4",X"27",X"15",X"96",X"00",X"80",X"01",X"97",X"00",X"24",X"07",
		X"86",X"04",X"97",X"00",X"7E",X"DE",X"4A",X"12",X"12",X"12",X"7E",X"DE",X"4A",X"8E",X"E0",X"EC",
		X"96",X"00",X"48",X"48",X"30",X"86",X"10",X"AE",X"94",X"EE",X"02",X"10",X"AE",X"A9",X"00",X"0E",
		X"26",X"06",X"6F",X"C4",X"10",X"BE",X"E1",X"00",X"10",X"AF",X"94",X"8E",X"E0",X"D8",X"96",X"00",
		X"48",X"48",X"30",X"86",X"EE",X"84",X"AE",X"02",X"30",X"88",X"E7",X"34",X"10",X"EC",X"A1",X"ED",
		X"C4",X"A6",X"A0",X"A7",X"84",X"30",X"03",X"EC",X"A1",X"ED",X"84",X"30",X"05",X"A6",X"A0",X"A7",
		X"84",X"30",X"03",X"EC",X"A1",X"ED",X"84",X"30",X"05",X"A6",X"A0",X"A7",X"84",X"30",X"03",X"EC",
		X"A1",X"ED",X"84",X"30",X"05",X"A6",X"A0",X"A7",X"84",X"30",X"03",X"EC",X"A4",X"ED",X"84",X"CC",
		X"00",X"00",X"30",X"03",X"ED",X"84",X"35",X"10",X"30",X"01",X"ED",X"84",X"ED",X"08",X"ED",X"88",
		X"10",X"ED",X"88",X"18",X"7E",X"DE",X"4A",X"DC",X"1D",X"D3",X"1F",X"DD",X"1D",X"DC",X"25",X"D3",
		X"27",X"DD",X"25",X"DC",X"2D",X"D3",X"2F",X"DD",X"2D",X"DC",X"35",X"D3",X"37",X"DD",X"35",X"DC",
		X"3D",X"D3",X"3F",X"DD",X"3D",X"DC",X"45",X"D3",X"47",X"DD",X"45",X"DC",X"55",X"D3",X"57",X"DD",
		X"55",X"4F",X"E6",X"9F",X"00",X"1C",X"58",X"49",X"EB",X"9F",X"00",X"24",X"89",X"00",X"EB",X"9F",
		X"00",X"2C",X"89",X"00",X"EB",X"9F",X"00",X"34",X"89",X"00",X"EB",X"9F",X"00",X"3C",X"89",X"00",
		X"EB",X"9F",X"00",X"44",X"89",X"00",X"EB",X"9F",X"00",X"54",X"89",X"00",X"58",X"49",X"58",X"49");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
