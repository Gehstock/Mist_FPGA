library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
--use IEEE.STD_LOGIC_ARITH.All;
--use ieee.std_logic_unsigned.all;

entity CharTable_ROM is
    Port ( ADDR : in  STD_LOGIC_VECTOR (8 downto 0);
           DATA_OUT : out  STD_LOGIC_VECTOR (7 downto 0));
end CharTable_ROM;

architecture Behavioral of CharTable_ROM is

	type ROM_TYPE is array (0 to 511)
        of std_logic_vector(7 downto 0);
		  
	constant ROM : ROM_TYPE :=
            (
-- addr=0x0000
X"00",X"0e",X"11",X"01",X"0d",X"15",X"15",X"0e",
X"00",X"04",X"0a",X"11",X"11",X"1f",X"11",X"11",
X"00",X"1e",X"09",X"09",X"0e",X"09",X"09",X"1e",
X"00",X"0e",X"11",X"10",X"10",X"10",X"11",X"0e",
X"00",X"1e",X"09",X"09",X"09",X"09",X"09",X"1e",
X"00",X"1f",X"10",X"10",X"1c",X"10",X"10",X"1f",
X"00",X"1f",X"10",X"10",X"1c",X"10",X"10",X"10",
X"00",X"0f",X"10",X"10",X"13",X"11",X"11",X"0f",
-- addr=0x0040
X"00",X"11",X"11",X"11",X"1f",X"11",X"11",X"11",
X"00",X"0e",X"04",X"04",X"04",X"04",X"04",X"0e",
X"00",X"01",X"01",X"01",X"01",X"01",X"11",X"0e",
X"00",X"11",X"12",X"14",X"18",X"14",X"12",X"11",
X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"1f",
X"00",X"11",X"1b",X"15",X"15",X"11",X"11",X"11",
X"00",X"11",X"19",X"15",X"13",X"11",X"11",X"11",
X"00",X"1f",X"11",X"11",X"11",X"11",X"11",X"1f",
-- addr=0x0080
X"00",X"1e",X"11",X"11",X"1e",X"10",X"10",X"10",
X"00",X"0e",X"11",X"11",X"11",X"15",X"12",X"0d",
X"00",X"1e",X"11",X"11",X"1e",X"14",X"12",X"11",
X"00",X"0e",X"11",X"08",X"04",X"02",X"11",X"0e",
X"00",X"1f",X"04",X"04",X"04",X"04",X"04",X"04",
X"00",X"11",X"11",X"11",X"11",X"11",X"11",X"0e",
X"00",X"11",X"11",X"11",X"0a",X"0a",X"04",X"04",
X"00",X"11",X"11",X"11",X"11",X"15",X"1b",X"11",
-- addr=0x00c0
X"00",X"11",X"11",X"0a",X"04",X"0a",X"11",X"11",
X"00",X"11",X"11",X"0a",X"04",X"04",X"04",X"04",
X"00",X"1f",X"01",X"02",X"04",X"08",X"10",X"1f",
X"00",X"0e",X"08",X"08",X"08",X"08",X"08",X"0e",
X"00",X"10",X"10",X"08",X"04",X"02",X"01",X"01",
X"00",X"0e",X"02",X"02",X"02",X"02",X"02",X"0e",
X"00",X"04",X"0e",X"15",X"04",X"04",X"04",X"04",
X"00",X"00",X"04",X"08",X"1f",X"08",X"04",X"00",
-- addr=0x0100
X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
X"00",X"04",X"04",X"04",X"04",X"04",X"00",X"04",
X"00",X"0a",X"0a",X"0a",X"00",X"00",X"00",X"00",
X"00",X"0a",X"0a",X"1b",X"00",X"1b",X"0a",X"0a",
X"00",X"04",X"0f",X"10",X"0e",X"01",X"1e",X"04",
X"00",X"19",X"19",X"02",X"04",X"08",X"13",X"13",
X"00",X"08",X"14",X"14",X"08",X"15",X"12",X"0d",
X"00",X"0c",X"0c",X"0c",X"00",X"00",X"00",X"00",
-- addr=0x0140
X"00",X"02",X"04",X"08",X"08",X"08",X"04",X"02",
X"00",X"08",X"04",X"02",X"02",X"02",X"04",X"08",
X"00",X"15",X"0e",X"1f",X"0e",X"15",X"00",X"00",
X"00",X"00",X"04",X"04",X"1f",X"04",X"04",X"00",
X"00",X"00",X"00",X"00",X"0c",X"0c",X"04",X"08",
X"00",X"00",X"00",X"00",X"1f",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"00",X"0c",X"0c",
X"00",X"01",X"01",X"02",X"04",X"08",X"10",X"10",
-- addr=0x0180
X"00",X"0c",X"12",X"12",X"12",X"12",X"12",X"0c",
X"00",X"04",X"0c",X"04",X"04",X"04",X"04",X"0e",
X"00",X"0e",X"11",X"01",X"0e",X"10",X"10",X"1f",
X"00",X"0e",X"11",X"01",X"06",X"01",X"11",X"0e",
X"00",X"02",X"06",X"0a",X"12",X"1f",X"02",X"02",
X"00",X"1f",X"10",X"1e",X"01",X"01",X"11",X"0e",
X"00",X"06",X"08",X"10",X"1e",X"11",X"11",X"0e",
X"00",X"1f",X"01",X"02",X"04",X"08",X"10",X"10",
-- addr=0x01c0
X"00",X"0e",X"11",X"11",X"0e",X"11",X"11",X"0e",
X"00",X"0e",X"11",X"11",X"0f",X"01",X"02",X"0c",
X"00",X"00",X"0c",X"0c",X"00",X"0c",X"0c",X"00",
X"00",X"0c",X"0c",X"00",X"0c",X"0c",X"04",X"08",
X"00",X"02",X"04",X"08",X"10",X"08",X"04",X"02",
X"00",X"00",X"00",X"1f",X"00",X"1f",X"00",X"00",
X"00",X"08",X"04",X"02",X"01",X"02",X"04",X"08",
X"00",X"0c",X"12",X"02",X"04",X"04",X"00",X"04"

-- 512 bytes
-- file: MCY7304NAA.bin
				);
				 
begin

	DATA_OUT <= ROM(to_integer(unsigned(ADDR)));

end Behavioral;

