`define BUILD_DATE "190308"
`define BUILD_TIME "223352"
