library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity rom_sprite_l is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of rom_sprite_l is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"3F",X"03",X"F5",X"0F",X"A5",X"3D",X"69",X"E5",X"59",X"DA",X"57",X"D5",X"AB",X"D5",X"57",
		X"F0",X"00",X"BF",X"00",X"95",X"C0",X"65",X"70",X"65",X"5C",X"FD",X"5C",X"0D",X"5C",X"33",X"5C",
		X"D6",X"81",X"EA",X"80",X"EA",X"80",X"35",X"55",X"0D",X"55",X"03",X"55",X"00",X"FF",X"00",X"00",
		X"C3",X"DC",X"CC",X"3C",X"F0",X"FC",X"4F",X"0C",X"57",X"3C",X"57",X"C0",X"FF",X"C0",X"00",X"00",
		X"0F",X"FF",X"3D",X"5A",X"3A",X"95",X"D5",X"6A",X"E9",X"55",X"D6",X"A9",X"D5",X"55",X"D6",X"05",
		X"FF",X"00",X"95",X"C0",X"65",X"70",X"59",X"5F",X"96",X"57",X"7F",X"FF",X"F0",X"C3",X"C3",X"C3",
		X"DA",X"03",X"EA",X"03",X"EA",X"95",X"35",X"55",X"0D",X"55",X"03",X"55",X"00",X"D5",X"00",X"3F",
		X"03",X"0F",X"C0",X"0C",X"F0",X"00",X"C0",X"00",X"CC",X"00",X"70",X"C0",X"73",X"00",X"FC",X"00",
		X"00",X"3F",X"03",X"D5",X"0D",X"55",X"3A",X"AA",X"35",X"57",X"3A",X"AC",X"F5",X"5C",X"D6",X"AC",
		X"F0",X"00",X"5C",X"00",X"57",X"00",X"95",X"C0",X"FF",X"FC",X"CC",X"FF",X"CC",X"CF",X"CC",X"CC",
		X"EA",X"5F",X"D5",X"60",X"DA",X"A0",X"FA",X"A0",X"3E",X"A9",X"0F",X"55",X"03",X"FF",X"00",X"00",
		X"FF",X"FF",X"15",X"57",X"15",X"5C",X"15",X"70",X"55",X"C0",X"57",X"00",X"FC",X"00",X"00",X"00",
		X"00",X"FF",X"0F",X"55",X"35",X"55",X"EA",X"AA",X"D5",X"55",X"DA",X"AA",X"E9",X"55",X"E5",X"AA",
		X"FF",X"F0",X"55",X"5C",X"55",X"FF",X"AB",X"CF",X"5C",X"C3",X"BC",X"C3",X"70",X"C0",X"B0",X"00",
		X"D6",X"95",X"DA",X"50",X"39",X"60",X"39",X"A8",X"0D",X"AA",X"03",X"A9",X"00",X"D5",X"00",X"3F",
		X"70",X"00",X"3C",X"00",X"0F",X"30",X"17",X"33",X"57",X"F3",X"55",X"FF",X"55",X"5F",X"FF",X"F0",
		X"00",X"3F",X"00",X"D6",X"03",X"A6",X"0E",X"A6",X"36",X"A5",X"36",X"A9",X"36",X"03",X"35",X"03",
		X"F0",X"00",X"7F",X"C0",X"59",X"B0",X"99",X"9C",X"99",X"9C",X"99",X"97",X"FF",X"97",X"03",X"97",
		X"35",X"03",X"35",X"57",X"35",X"57",X"0D",X"57",X"03",X"57",X"00",X"D7",X"00",X"37",X"00",X"0F",
		X"FF",X"97",X"03",X"57",X"FF",X"5C",X"03",X"70",X"FF",X"C0",X"0F",X"00",X"FC",X"00",X"3C",X"00",
		X"00",X"0F",X"00",X"F5",X"03",X"A9",X"0D",X"5A",X"3A",X"96",X"DA",X"A5",X"DA",X"81",X"D6",X"01",
		X"FF",X"C0",X"A5",X"B0",X"69",X"9C",X"59",X"9C",X"99",X"97",X"99",X"97",X"99",X"97",X"99",X"97",
		X"D5",X"01",X"D5",X"4F",X"D5",X"7C",X"D7",X"F0",X"DF",X"00",X"DF",X"F0",X"3C",X"00",X"3F",X"C0",
		X"99",X"97",X"FD",X"97",X"0F",X"97",X"00",X"D7",X"3F",X"F7",X"00",X"37",X"00",X"FC",X"0F",X"F0",
		X"02",X"00",X"0F",X"FF",X"3F",X"FF",X"FF",X"FF",X"00",X"05",X"00",X"54",X"01",X"50",X"01",X"40",
		X"02",X"00",X"FF",X"C0",X"FF",X"F0",X"FF",X"FC",X"40",X"00",X"54",X"00",X"15",X"00",X"05",X"00",
		X"00",X"00",X"2A",X"00",X"2A",X"00",X"55",X"55",X"5A",X"81",X"5A",X"81",X"5A",X"A9",X"15",X"55",
		X"00",X"00",X"02",X"A0",X"02",X"A0",X"55",X"54",X"0A",X"94",X"0A",X"94",X"AA",X"94",X"55",X"50",
		X"00",X"AA",X"0A",X"A0",X"2A",X"00",X"AA",X"FC",X"AA",X"CF",X"55",X"50",X"55",X"EC",X"57",X"EF",
		X"AA",X"A8",X"00",X"00",X"00",X"00",X"3F",X"C0",X"F0",X"FC",X"00",X"00",X"00",X"00",X"55",X"55",
		X"16",X"AA",X"07",X"EF",X"00",X"ED",X"00",X"00",X"00",X"3F",X"03",X"FF",X"0F",X"C0",X"00",X"FF",
		X"55",X"55",X"55",X"50",X"55",X"00",X"00",X"00",X"FF",X"00",X"0F",X"F0",X"00",X"FC",X"FF",X"C0",
		X"02",X"00",X"02",X"00",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"A0",X"54",X"A1",X"45",X"A0",X"00",
		X"02",X"00",X"02",X"00",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"A8",
		X"A0",X"00",X"55",X"55",X"59",X"99",X"59",X"99",X"59",X"99",X"15",X"55",X"00",X"00",X"00",X"00",
		X"00",X"A8",X"55",X"55",X"6A",X"05",X"6A",X"05",X"6A",X"A5",X"55",X"54",X"00",X"00",X"00",X"00",
		X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"A0",X"50",X"A1",X"55",X"A1",X"45",X"A0",X"00",X"A0",X"00",
		X"FF",X"F0",X"FF",X"FC",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"55",X"55",X"59",X"99",X"15",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A8",X"55",X"55",X"6A",X"15",X"55",X"54",
		X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"55",X"55",
		X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"55",X"55",
		X"59",X"99",X"59",X"99",X"59",X"99",X"15",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"42",X"A5",X"42",X"A5",X"6A",X"A5",X"55",X"54",X"30",X"00",X"30",X"14",X"0C",X"14",X"03",X"C0",
		X"0F",X"FF",X"0C",X"F5",X"F0",X"CD",X"DF",X"0F",X"D7",X"30",X"D5",X"C3",X"D5",X"FC",X"D5",X"0F",
		X"FC",X"00",X"57",X"00",X"55",X"C0",X"55",X"70",X"F5",X"70",X"3A",X"7C",X"35",X"AC",X"F5",X"5C",
		X"D5",X"03",X"D5",X"01",X"D5",X"A9",X"35",X"A9",X"0D",X"A5",X"03",X"A5",X"00",X"FF",X"00",X"00",
		X"9A",X"5C",X"96",X"BC",X"95",X"B0",X"65",X"F0",X"67",X"C0",X"5F",X"00",X"FC",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"80",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"80",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",
		X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",
		X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",
		X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",
		X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",
		X"01",X"00",X"05",X"40",X"17",X"50",X"1F",X"D0",X"17",X"50",X"05",X"40",X"01",X"00",X"02",X"00",
		X"05",X"40",X"17",X"50",X"5F",X"D4",X"17",X"50",X"05",X"40",X"02",X"00",X"02",X"00",X"02",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"1A",X"00",X"6B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"90",X"00",X"A4",X"00",
		X"00",X"6F",X"00",X"6B",X"00",X"1A",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"24",X"00",X"A4",X"00",X"90",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"80",X"02",X"05",X"00",X"1F",X"00",X"7E",X"08",X"7A",
		X"00",X"00",X"00",X"00",X"80",X"00",X"02",X"00",X"50",X"80",X"F4",X"00",X"BD",X"00",X"AD",X"20",
		X"08",X"7A",X"00",X"7E",X"00",X"1F",X"02",X"05",X"00",X"80",X"00",X"02",X"00",X"00",X"00",X"00",
		X"AD",X"20",X"BD",X"00",X"F4",X"00",X"50",X"80",X"02",X"00",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"54",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"20",X"00",X"90",X"00",
		X"00",X"01",X"00",X"15",X"00",X"55",X"00",X"54",X"00",X"50",X"00",X"00",X"00",X"04",X"00",X"00",
		X"00",X"10",X"80",X"90",X"00",X"90",X"02",X"40",X"02",X"40",X"05",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"08",X"04",X"02",
		X"00",X"00",X"00",X"00",X"02",X"00",X"0C",X"00",X"02",X"80",X"00",X"20",X"00",X"00",X"00",X"00",
		X"0C",X"02",X"06",X"00",X"06",X"00",X"02",X"00",X"02",X"00",X"00",X"00",X"00",X"20",X"00",X"00",
		X"80",X"20",X"A0",X"00",X"9C",X"00",X"19",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"08",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"02",X"80",X"02",X"B0",X"00",X"7A",X"00",X"05",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"0B",X"00",X"03",X"80",X"C0",X"80",
		X"00",X"02",X"00",X"00",X"03",X"00",X"07",X"C0",X"06",X"0C",X"02",X"02",X"00",X"00",X"00",X"00",
		X"C0",X"40",X"A0",X"20",X"28",X"00",X"02",X"00",X"00",X"00",X"80",X"00",X"20",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"51",X"02",X"50",X"01",X"50",X"01",X"10",X"10",X"40",
		X"00",X"00",X"10",X"00",X"00",X"00",X"01",X"40",X"01",X"40",X"0D",X"00",X"20",X"04",X"40",X"00",
		X"07",X"02",X"04",X"00",X"04",X"00",X"20",X"10",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"C0",X"05",X"C0",X"20",X"00",X"00",X"04",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"26",X"00",X"66",X"01",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"43",X"F0",X"4F",X"FC",X"7F",X"0F",X"7C",X"03",
		X"01",X"66",X"01",X"66",X"00",X"66",X"00",X"26",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"00",X"7C",X"03",X"7F",X"0F",X"4F",X"FC",X"43",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"3C",X"10",X"FF",X"13",X"FF",X"9F",X"C3",X"9F",X"03",X"9C",X"03",
		X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"90",X"00",X"9C",X"03",X"9F",X"03",X"9F",X"03",X"13",X"FF",X"10",X"FF",X"00",X"3C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"69",X"0A",X"69",X"1A",X"69",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"C0",X"FF",X"FF",
		X"5A",X"69",X"1A",X"69",X"0A",X"69",X"00",X"69",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"3C",X"00",X"CF",X"00",X"03",X"00",X"03",X"00",X"0F",X"00",X"0D",X"00",X"05",X"00",X"2A",
		X"0F",X"00",X"3C",X"C0",X"30",X"00",X"30",X"00",X"3C",X"00",X"5C",X"00",X"54",X"00",X"AA",X"00",
		X"00",X"2A",X"00",X"2A",X"00",X"05",X"00",X"05",X"00",X"02",X"00",X"02",X"00",X"00",X"00",X"00",
		X"AA",X"00",X"AA",X"00",X"54",X"00",X"54",X"00",X"A0",X"00",X"A0",X"00",X"40",X"00",X"00",X"00",
		X"00",X"3C",X"00",X"F0",X"03",X"C0",X"03",X"C0",X"03",X"F0",X"00",X"35",X"00",X"15",X"00",X"AA",
		X"0F",X"00",X"03",X"C0",X"00",X"F0",X"00",X"F0",X"03",X"F0",X"57",X"00",X"55",X"00",X"AA",X"80",
		X"00",X"AA",X"00",X"15",X"00",X"15",X"00",X"0A",X"00",X"0A",X"00",X"01",X"00",X"00",X"00",X"00",
		X"AA",X"80",X"55",X"00",X"55",X"00",X"A8",X"00",X"A8",X"00",X"50",X"00",X"00",X"00",X"00",X"00",
		X"03",X"F0",X"0F",X"00",X"3C",X"00",X"3C",X"00",X"0F",X"F0",X"03",X"D5",X"05",X"55",X"0A",X"AA",
		X"03",X"F0",X"00",X"3C",X"00",X"0F",X"00",X"0F",X"03",X"FC",X"55",X"F0",X"55",X"54",X"AA",X"A8",
		X"02",X"AA",X"00",X"55",X"00",X"15",X"00",X"0A",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"A0",X"55",X"40",X"55",X"00",X"A8",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"0F",X"00",X"0F",X"00",X"0F",
		X"05",X"40",X"15",X"50",X"D5",X"54",X"D5",X"05",X"D4",X"01",X"DA",X"03",X"EA",X"03",X"EA",X"0F",
		X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"03",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EA",X"FF",X"FF",X"CF",X"FF",X"CF",X"FC",X"00",X"FF",X"CF",X"FF",X"CC",X"3F",X"F0",X"0F",X"C0",
		X"00",X"55",X"05",X"55",X"15",X"57",X"55",X"15",X"55",X"15",X"50",X"01",X"55",X"15",X"15",X"14",
		X"55",X"40",X"FD",X"50",X"FE",X"94",X"4A",X"94",X"4E",X"A4",X"0E",X"A8",X"0C",X"28",X"0F",X"08",
		X"05",X"50",X"00",X"54",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"28",X"03",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"41",X"00",X"41",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"51",X"50",X"11",X"10",
		X"00",X"41",X"00",X"41",X"01",X"41",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"10",X"11",X"10",X"51",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"41",X"00",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"51",X"50",X"11",X"10",
		X"00",X"41",X"00",X"41",X"01",X"41",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"51",X"10",X"01",X"10",X"51",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"51",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"51",X"50",X"11",X"10",
		X"01",X"51",X"00",X"11",X"01",X"51",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"10",X"11",X"10",X"51",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"51",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"51",X"50",X"11",X"10",
		X"01",X"51",X"00",X"11",X"01",X"51",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"51",X"10",X"01",X"10",X"51",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"51",X"00",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"51",X"50",X"11",X"10",
		X"01",X"51",X"00",X"11",X"01",X"51",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"10",X"11",X"10",X"51",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"51",X"00",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"51",X"50",X"11",X"10",
		X"01",X"51",X"00",X"11",X"01",X"51",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"51",X"10",X"01",X"10",X"51",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"01",X"51",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"51",X"50",X"11",X"10",
		X"01",X"11",X"01",X"11",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"10",X"11",X"10",X"51",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"01",X"50",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"51",X"50",X"11",X"10",
		X"01",X"11",X"01",X"11",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"51",X"10",X"01",X"10",X"51",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"2A",X"00",X"AA",X"00",X"AB",X"03",X"FF",X"03",X"FF",X"3F",X"FF",X"FF",X"FF",X"55",X"55",
		X"55",X"80",X"FE",X"80",X"FE",X"00",X"FF",X"F0",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"55",X"54",
		X"55",X"5A",X"55",X"6A",X"55",X"6A",X"55",X"6A",X"15",X"6A",X"15",X"5A",X"05",X"55",X"00",X"55",
		X"AA",X"95",X"80",X"15",X"00",X"15",X"00",X"54",X"81",X"50",X"A5",X"50",X"55",X"40",X"50",X"00",
		X"00",X"2A",X"00",X"AA",X"00",X"AB",X"03",X"FF",X"0F",X"FF",X"3F",X"FF",X"FF",X"FF",X"55",X"55",
		X"55",X"80",X"FE",X"80",X"FE",X"00",X"FF",X"C0",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"55",X"54",
		X"55",X"5A",X"55",X"6A",X"55",X"6A",X"55",X"6A",X"15",X"6A",X"15",X"5A",X"05",X"55",X"00",X"55",
		X"AA",X"95",X"80",X"15",X"00",X"15",X"00",X"54",X"81",X"50",X"A5",X"50",X"55",X"40",X"50",X"00",
		X"00",X"05",X"00",X"15",X"00",X"15",X"00",X"57",X"00",X"5F",X"00",X"5D",X"00",X"5F",X"00",X"57",
		X"40",X"00",X"50",X"00",X"50",X"00",X"54",X"00",X"D4",X"00",X"D4",X"00",X"D4",X"00",X"54",X"00",
		X"00",X"15",X"00",X"15",X"00",X"05",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",
		X"50",X"00",X"50",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"15",X"01",X"55",X"05",X"5F",X"05",X"7D",X"05",X"5F",X"01",X"55",X"00",X"15",X"00",X"02",
		X"50",X"00",X"55",X"00",X"D5",X"00",X"F5",X"40",X"D5",X"40",X"55",X"00",X"50",X"00",X"00",X"00",
		X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"00",X"2A",X"00",X"A9",X"03",X"E6",X"0B",X"FE",X"2A",X"FF",X"29",X"FF",X"A6",X"BF",
		X"A4",X"00",X"5A",X"80",X"AA",X"90",X"AA",X"68",X"A9",X"A8",X"A6",X"A9",X"DA",X"A6",X"FA",X"A6",
		X"9A",X"AF",X"9A",X"A7",X"6A",X"9A",X"2A",X"6A",X"29",X"AA",X"06",X"AA",X"02",X"A5",X"00",X"1A",
		X"FE",X"9A",X"FF",X"68",X"FF",X"A8",X"BF",X"E0",X"9B",X"C0",X"6A",X"00",X"A8",X"00",X"80",X"00",
		X"00",X"00",X"00",X"AB",X"2A",X"AB",X"AA",X"5F",X"95",X"AF",X"6A",X"AF",X"AA",X"AF",X"5A",X"5F",
		X"00",X"00",X"EA",X"00",X"EA",X"A8",X"F5",X"AA",X"FA",X"56",X"FA",X"A9",X"FA",X"AA",X"FA",X"5A",
		X"A5",X"AF",X"AA",X"AF",X"6A",X"AF",X"95",X"AF",X"AA",X"5F",X"2A",X"AB",X"00",X"AB",X"00",X"00",
		X"F5",X"A5",X"FA",X"AA",X"FA",X"A9",X"FA",X"56",X"F5",X"AA",X"EA",X"A8",X"EA",X"00",X"00",X"00",
		X"3F",X"0F",X"0C",X"3F",X"3F",X"FF",X"3F",X"FF",X"FF",X"FF",X"6A",X"6A",X"6A",X"6A",X"6A",X"6A",
		X"F0",X"FC",X"FC",X"30",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"A9",X"A9",X"A9",X"A9",X"A9",X"A9",
		X"6A",X"6A",X"6A",X"5A",X"5A",X"9A",X"16",X"96",X"05",X"A6",X"01",X"55",X"00",X"0C",X"00",X"3F",
		X"A9",X"A9",X"A5",X"A9",X"A6",X"A5",X"96",X"94",X"9A",X"50",X"55",X"40",X"30",X"00",X"FC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"A0",X"0A",X"14",X"14",X"05",X"50",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"A0",X"0A",X"14",X"14",X"05",X"50",
		X"05",X"50",X"14",X"14",X"A0",X"0A",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"05",X"50",X"14",X"14",X"A0",X"0A",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"9A",X"0A",X"6A",X"0A",X"69",X"2A",X"69",X"29",X"AA",X"29",X"AA",X"2B",X"FF",X"3F",X"FF",
		X"66",X"80",X"69",X"A0",X"A9",X"A0",X"A9",X"A8",X"6A",X"68",X"6A",X"68",X"FF",X"E8",X"FF",X"FC",
		X"3F",X"FF",X"2B",X"FF",X"29",X"A9",X"29",X"A9",X"2A",X"6A",X"0A",X"6A",X"0A",X"69",X"02",X"99",
		X"FF",X"FC",X"FF",X"E8",X"AA",X"68",X"AA",X"68",X"69",X"68",X"69",X"A0",X"A9",X"A0",X"A6",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"01",X"00",X"30",X"00",X"C0",X"C0",X"0C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"84",X"00",X"02",X"00",X"00",X"40",X"48",X"00",
		X"00",X"00",X"C0",X"CC",X"0C",X"01",X"00",X"C1",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"48",X"00",X"24",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"C2",X"0C",X"C0",X"C0",X"CC",X"C0",X"0E",X"00",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"44",X"00",X"66",X"00",X"A4",X"40",X"92",X"40",
		X"C0",X"0E",X"C0",X"CD",X"0C",X"C1",X"0C",X"C1",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"19",X"40",X"89",X"00",X"20",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"00",X"0F",X"00",X"00",X"0C",X"00",X"30",X"03",X"C3",X"00",X"FC",X"30",X"D7",X"FC",
		X"FF",X"C0",X"0D",X"C0",X"0D",X"70",X"FD",X"5C",X"CE",X"57",X"0D",X"97",X"3D",X"67",X"F6",X"5B",
		X"D5",X"5F",X"D5",X"50",X"D5",X"50",X"35",X"60",X"0D",X"6A",X"03",X"6A",X"00",X"E9",X"00",X"3F",
		X"65",X"9B",X"59",X"9B",X"19",X"97",X"19",X"67",X"59",X"67",X"56",X"6F",X"56",X"70",X"FF",X"C0");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
