library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity TRIPLEDRAWPOKER_1K is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of TRIPLEDRAWPOKER_1K is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"0F",X"1F",X"3F",X"7F",X"FF",
		X"FF",X"7F",X"3F",X"1F",X"0F",X"07",X"03",X"01",X"F0",X"F8",X"FC",X"FC",X"FC",X"F8",X"F0",X"E0",
		X"E0",X"F0",X"F8",X"FC",X"FC",X"FC",X"F8",X"F0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"00",X"00",X"60",X"70",X"78",X"7C",X"6E",X"67",
		X"00",X"00",X"60",X"70",X"78",X"7C",X"7E",X"7F",X"00",X"00",X"1C",X"1E",X"1F",X"0F",X"07",X"07",
		X"7F",X"77",X"73",X"71",X"70",X"70",X"70",X"00",X"87",X"C7",X"E7",X"FF",X"FF",X"7E",X"3C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"18",X"38",X"78",X"70",X"70",X"71",X"00",X"00",X"0C",X"0E",X"0F",X"07",X"07",X"C7",
		X"FF",X"E0",X"E0",X"FE",X"FE",X"FE",X"E0",X"E0",X"FF",X"07",X"07",X"7F",X"7F",X"7F",X"07",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"E0",X"E0",X"E6",X"E6",X"E6",X"E7",X"E7",X"FF",X"07",X"07",X"67",X"67",X"67",X"E7",X"E7",
		X"00",X"0E",X"0F",X"0F",X"0F",X"0F",X"0E",X"0E",X"00",X"00",X"00",X"80",X"C0",X"E0",X"F0",X"78",
		X"6E",X"6E",X"7F",X"7F",X"7F",X"6E",X"6E",X"00",X"3C",X"1E",X"FF",X"FF",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"18",X"39",X"79",X"79",X"71",X"71",X"00",X"00",X"FF",X"FF",X"FF",X"C7",X"C7",X"C7",
		X"FF",X"E0",X"E0",X"E7",X"E7",X"E7",X"E7",X"FF",X"C7",X"C7",X"C7",X"C7",X"C7",X"87",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"07",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"1F",X"3F",X"7F",X"7B",X"71",X"71",X"00",X"00",X"FC",X"FE",X"FF",X"EF",X"C7",X"C7",
		X"07",X"07",X"E7",X"E7",X"C7",X"0F",X"1F",X"FF",X"C7",X"C7",X"C7",X"C7",X"CF",X"8E",X"0C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"E0",X"E7",X"E7",X"E3",X"F0",X"F8",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"60",X"78",X"7E",X"00",X"00",X"1F",X"1F",X"1F",X"07",X"07",X"07",
		X"7F",X"1F",X"07",X"01",X"00",X"00",X"00",X"00",X"87",X"E7",X"FF",X"FF",X"7F",X"1F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"1E",X"3F",X"7F",X"7B",X"71",X"71",X"00",X"00",X"3C",X"FE",X"FF",X"EF",X"C7",X"C7",
		X"71",X"71",X"71",X"7B",X"7F",X"3F",X"1E",X"00",X"C7",X"C7",X"C7",X"EF",X"FF",X"FE",X"3C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"18",X"38",X"79",X"71",X"71",X"71",X"00",X"00",X"7C",X"FE",X"FF",X"EF",X"C7",X"C7",
		X"71",X"71",X"71",X"78",X"7F",X"3F",X"1F",X"00",X"C7",X"C7",X"C7",X"EF",X"FF",X"FE",X"FC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"3F",X"3F",X"3F",X"00",X"00",X"1F",X"3F",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"FE",X"FF",
		X"3F",X"38",X"38",X"38",X"3F",X"3F",X"1F",X"00",X"FF",X"07",X"07",X"07",X"FF",X"FF",X"FE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0C",X"1C",X"3C",X"38",X"38",X"38",X"38",X"00",X"00",X"00",X"07",X"07",X"07",X"07",X"07",
		X"3C",X"3F",X"1F",X"0F",X"00",X"00",X"00",X"00",X"07",X"FF",X"FF",X"FF",X"07",X"07",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"3F",X"7F",X"7F",X"78",X"70",X"70",X"00",X"00",X"FE",X"FF",X"FF",X"0F",X"07",X"E7",
		X"71",X"7B",X"7F",X"7F",X"3F",X"1E",X"3C",X"38",X"E7",X"CF",X"FF",X"FF",X"FE",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"60",X"7F",X"7F",X"7F",X"63",X"01",X"03",X"00",X"03",X"FF",X"FF",X"FF",X"C3",X"E0",X"F0",
		X"07",X"6F",X"7E",X"7C",X"78",X"70",X"60",X"00",X"FB",X"3F",X"1F",X"0F",X"07",X"03",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"60",X"7C",X"7F",X"7F",X"67",X"07",X"06",X"06",X"00",X"00",X"00",X"C0",X"F0",X"FC",X"3F",X"1F",
		X"06",X"06",X"07",X"67",X"7F",X"7F",X"7C",X"60",X"1F",X"3F",X"FC",X"F0",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"03",X"07",X"0F",X"1F",X"3F",X"7F",X"FF",X"00",X"80",X"C0",X"E0",X"F0",X"F8",X"FC",X"FE",
		X"FF",X"7F",X"3F",X"1F",X"0F",X"07",X"03",X"01",X"FE",X"FC",X"F8",X"F0",X"E0",X"C0",X"80",X"00",
		X"83",X"43",X"24",X"18",X"18",X"24",X"42",X"81",X"81",X"42",X"24",X"18",X"18",X"24",X"43",X"83",
		X"C1",X"C2",X"24",X"18",X"18",X"24",X"42",X"81",X"81",X"42",X"24",X"18",X"18",X"24",X"C2",X"C1",
		X"81",X"42",X"24",X"18",X"18",X"24",X"42",X"81",X"81",X"42",X"24",X"18",X"18",X"00",X"00",X"81",
		X"81",X"00",X"00",X"00",X"00",X"00",X"00",X"81",X"81",X"00",X"00",X"00",X"00",X"00",X"00",X"81",
		X"80",X"00",X"00",X"18",X"18",X"24",X"42",X"81",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"1F",X"1F",X"03",X"07",X"0F",X"1D",X"18",X"00",
		X"F8",X"F8",X"18",X"18",X"18",X"F8",X"F0",X"00",X"00",X"1F",X"1F",X"19",X"19",X"19",X"18",X"18",
		X"00",X"F8",X"F8",X"98",X"98",X"98",X"18",X"18",X"00",X"1F",X"1F",X"18",X"18",X"1C",X"0F",X"07",
		X"00",X"F8",X"F8",X"18",X"18",X"38",X"F0",X"E0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E7",X"DB",X"DB",X"DB",X"FF",X"FF",
		X"FF",X"E0",X"E0",X"E6",X"E6",X"E6",X"E0",X"F1",X"FF",X"07",X"07",X"67",X"67",X"67",X"07",X"8F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E0",X"E0",X"E6",X"E6",X"E6",X"E7",X"E7",
		X"FF",X"07",X"07",X"67",X"67",X"67",X"E7",X"E7",X"FF",X"FF",X"FF",X"E0",X"E0",X"FF",X"FF",X"FF",
		X"FF",X"E7",X"E7",X"07",X"07",X"E7",X"E7",X"FF",X"FF",X"E0",X"E0",X"E7",X"E7",X"E3",X"F0",X"F8",
		X"FF",X"07",X"07",X"E7",X"E7",X"C7",X"0F",X"1F",X"FF",X"E0",X"E0",X"FE",X"FE",X"FE",X"E0",X"E0",
		X"FF",X"0F",X"07",X"67",X"67",X"67",X"07",X"0F",X"FF",X"E0",X"E0",X"E7",X"E7",X"E7",X"E7",X"FF",
		X"FF",X"07",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
