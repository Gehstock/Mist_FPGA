library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity silverland_program is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of silverland_program is
	type rom is array(0 to  24575) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"08",X"D9",X"ED",X"56",X"C3",X"52",X"00",X"0B",X"F5",X"E5",X"D5",X"C5",X"C3",X"2D",X"04",X"2A",
		X"F5",X"E5",X"D5",X"C5",X"C3",X"8A",X"04",X"32",X"8F",X"0B",X"21",X"9F",X"0B",X"06",X"B1",X"36",
		X"F5",X"E5",X"D5",X"C5",X"C3",X"3A",X"05",X"0B",X"F5",X"E5",X"D5",X"C5",X"C3",X"5F",X"05",X"5E",
		X"22",X"09",X"80",X"C3",X"69",X"05",X"C1",X"0B",X"CD",X"28",X"09",X"CD",X"64",X"09",X"C1",X"CB",
		X"40",X"20",X"0D",X"E5",X"21",X"C1",X"0B",X"11",X"3A",X"00",X"B8",X"C3",X"D1",X"02",X"B0",X"E1",
		X"06",X"01",X"01",X"00",X"00",X"3A",X"00",X"B8",X"3E",X"05",X"3D",X"20",X"FD",X"10",X"F9",X"0D",
		X"20",X"F3",X"C3",X"48",X"00",X"28",X"08",X"D9",X"FD",X"E5",X"DD",X"E5",X"AF",X"32",X"00",X"A0",
		X"3A",X"13",X"80",X"FE",X"FF",X"C2",X"EC",X"00",X"21",X"04",X"80",X"3A",X"00",X"B8",X"CB",X"47",
		X"28",X"04",X"36",X"01",X"18",X"0F",X"7E",X"36",X"00",X"B7",X"28",X"09",X"2B",X"7E",X"3C",X"3C",
		X"FE",X"C8",X"30",X"01",X"77",X"CD",X"25",X"01",X"CD",X"E7",X"47",X"2A",X"09",X"80",X"7C",X"B5",
		X"28",X"04",X"2B",X"22",X"09",X"80",X"21",X"11",X"80",X"35",X"3E",X"18",X"86",X"20",X"3D",X"36",
		X"00",X"11",X"14",X"80",X"EB",X"CB",X"7E",X"20",X"30",X"23",X"3E",X"05",X"BE",X"20",X"2A",X"13",
		X"1A",X"EE",X"01",X"12",X"20",X"15",X"3A",X"16",X"80",X"CB",X"77",X"20",X"07",X"3E",X"12",X"CD",
		X"12",X"0D",X"18",X"15",X"3E",X"13",X"CD",X"12",X"0D",X"18",X"0E",X"3A",X"16",X"80",X"CB",X"77",
		X"3E",X"02",X"20",X"02",X"3E",X"00",X"CD",X"12",X"0D",X"CD",X"07",X"01",X"21",X"11",X"80",X"3E",
		X"01",X"CB",X"46",X"28",X"02",X"3E",X"02",X"32",X"06",X"80",X"3E",X"01",X"32",X"00",X"A0",X"DD",
		X"E1",X"FD",X"E1",X"D9",X"08",X"ED",X"45",X"21",X"24",X"24",X"22",X"BB",X"93",X"22",X"BD",X"93",
		X"21",X"BD",X"93",X"3A",X"03",X"80",X"0F",X"0E",X"00",X"0C",X"D6",X"0A",X"30",X"FB",X"0D",X"C6",
		X"0A",X"77",X"2B",X"71",X"C9",X"06",X"08",X"11",X"80",X"98",X"21",X"47",X"82",X"0E",X"04",X"7E",
		X"CB",X"7F",X"20",X"14",X"23",X"B7",X"28",X"07",X"13",X"23",X"0D",X"20",X"FB",X"18",X"12",X"AF",
		X"12",X"23",X"13",X"0D",X"20",X"FA",X"18",X"09",X"CB",X"BE",X"23",X"ED",X"A0",X"AF",X"B1",X"20",
		X"FA",X"10",X"DA",X"C9",X"E5",X"21",X"47",X"82",X"06",X"08",X"3A",X"00",X"80",X"4F",X"16",X"00",
		X"7E",X"E6",X"7F",X"B9",X"20",X"02",X"16",X"01",X"23",X"23",X"23",X"23",X"23",X"10",X"F1",X"E1",
		X"7A",X"B7",X"C0",X"7D",X"45",X"21",X"05",X"80",X"86",X"FE",X"09",X"3F",X"D8",X"77",X"21",X"47",
		X"82",X"7E",X"B7",X"20",X"07",X"3A",X"00",X"80",X"77",X"10",X"F6",X"C9",X"11",X"05",X"00",X"19",
		X"18",X"EF",X"7C",X"C6",X"20",X"67",X"7D",X"C6",X"10",X"6F",X"D5",X"FD",X"E1",X"50",X"59",X"DD",
		X"21",X"47",X"82",X"06",X"08",X"3A",X"00",X"80",X"4F",X"DD",X"7E",X"00",X"E6",X"7F",X"B9",X"20",
		X"21",X"DD",X"72",X"01",X"14",X"DD",X"73",X"02",X"7C",X"FD",X"86",X"00",X"DD",X"77",X"04",X"FD",
		X"23",X"7D",X"FD",X"86",X"00",X"DD",X"77",X"03",X"FD",X"23",X"78",X"FE",X"06",X"30",X"03",X"DD",
		X"35",X"03",X"D5",X"11",X"05",X"00",X"DD",X"19",X"D1",X"10",X"CE",X"3E",X"00",X"32",X"00",X"A0",
		X"21",X"47",X"82",X"06",X"08",X"11",X"05",X"00",X"3A",X"00",X"80",X"4F",X"7E",X"E6",X"7F",X"B9",
		X"20",X"02",X"CB",X"FE",X"19",X"10",X"F5",X"3E",X"01",X"32",X"00",X"A0",X"C9",X"21",X"47",X"82",
		X"06",X"08",X"3A",X"00",X"80",X"4F",X"7E",X"E6",X"7F",X"B9",X"20",X"08",X"36",X"00",X"11",X"05",
		X"80",X"1A",X"3D",X"12",X"11",X"05",X"00",X"19",X"10",X"EC",X"C9",X"3A",X"23",X"80",X"E6",X"F8",
		X"32",X"23",X"80",X"3A",X"14",X"80",X"CB",X"47",X"20",X"20",X"CB",X"7F",X"20",X"35",X"3A",X"16",
		X"80",X"CB",X"77",X"20",X"05",X"3A",X"00",X"A8",X"18",X"03",X"3A",X"00",X"A0",X"E6",X"C1",X"07",
		X"07",X"47",X"3A",X"23",X"80",X"B0",X"32",X"23",X"80",X"C9",X"2A",X"0B",X"80",X"11",X"0F",X"80",
		X"CD",X"B7",X"02",X"22",X"0B",X"80",X"30",X"E9",X"21",X"7C",X"02",X"22",X"0B",X"80",X"EB",X"36",
		X"00",X"18",X"E7",X"2A",X"0D",X"80",X"11",X"10",X"80",X"CD",X"B7",X"02",X"22",X"0D",X"80",X"30",
		X"D0",X"21",X"85",X"02",X"22",X"0D",X"80",X"EB",X"36",X"00",X"18",X"E7",X"A4",X"F4",X"65",X"F4",
		X"F4",X"84",X"F6",X"F4",X"FF",X"F5",X"55",X"F4",X"64",X"72",X"66",X"F6",X"52",X"80",X"F5",X"45",
		X"F4",X"F4",X"24",X"86",X"A2",X"F6",X"26",X"F4",X"A4",X"F5",X"F4",X"F4",X"F4",X"86",X"F2",X"82",
		X"66",X"F4",X"F5",X"55",X"F4",X"11",X"F4",X"F4",X"F6",X"F4",X"80",X"F4",X"F0",X"F4",X"F0",X"F4",
		X"F0",X"F4",X"F0",X"F4",X"F4",X"F4",X"FF",X"1A",X"47",X"3C",X"12",X"7E",X"FE",X"FF",X"37",X"C8",
		X"E6",X"F0",X"0F",X"0F",X"0F",X"0F",X"4E",X"B8",X"20",X"03",X"23",X"AF",X"12",X"79",X"E6",X"07",
		X"C9",X"AF",X"A7",X"DD",X"21",X"D9",X"02",X"18",X"1C",X"08",X"3C",X"DD",X"21",X"E1",X"02",X"18",
		X"14",X"08",X"AF",X"37",X"DD",X"21",X"EA",X"02",X"18",X"0B",X"08",X"3C",X"DD",X"21",X"F2",X"02",
		X"18",X"03",X"C3",X"D0",X"03",X"11",X"B6",X"03",X"21",X"1F",X"03",X"28",X"03",X"21",X"33",X"03",
		X"38",X"05",X"08",X"1A",X"2F",X"18",X"02",X"08",X"1A",X"FD",X"21",X"14",X"03",X"4F",X"13",X"1A",
		X"47",X"13",X"1A",X"E9",X"13",X"1A",X"FE",X"ED",X"28",X"03",X"08",X"18",X"DB",X"DD",X"E9",X"67",
		X"2E",X"00",X"3A",X"00",X"B8",X"71",X"2C",X"20",X"FC",X"24",X"10",X"F6",X"1A",X"67",X"79",X"2F",
		X"77",X"FD",X"E9",X"67",X"2E",X"00",X"7E",X"2F",X"A9",X"20",X"1F",X"2C",X"3A",X"00",X"B8",X"7E",
		X"A9",X"20",X"17",X"1A",X"FE",X"98",X"20",X"0A",X"2C",X"CB",X"6D",X"28",X"04",X"7D",X"C6",X"20",
		X"6F",X"2D",X"2C",X"20",X"EA",X"24",X"10",X"E4",X"FD",X"E9",X"4F",X"D9",X"AF",X"37",X"DD",X"21",
		X"64",X"03",X"18",X"91",X"21",X"18",X"91",X"D9",X"EB",X"79",X"21",X"6F",X"03",X"18",X"30",X"D9",
		X"2D",X"D9",X"7B",X"21",X"78",X"03",X"18",X"27",X"7A",X"21",X"7E",X"03",X"18",X"21",X"D9",X"21",
		X"B0",X"03",X"11",X"08",X"91",X"01",X"06",X"00",X"ED",X"B0",X"D9",X"3A",X"00",X"B0",X"CB",X"7F",
		X"CA",X"00",X"00",X"3A",X"00",X"B8",X"AF",X"12",X"1A",X"3E",X"FF",X"12",X"1A",X"18",X"EC",X"D9",
		X"4F",X"E6",X"0F",X"77",X"2D",X"79",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"77",X"2B",X"D9",X"E9",
		X"0B",X"0A",X"0D",X"1B",X"0A",X"16",X"00",X"04",X"80",X"FF",X"01",X"88",X"24",X"04",X"90",X"00",
		X"08",X"98",X"ED",X"00",X"0B",X"0A",X"0D",X"1B",X"18",X"16",X"90",X"01",X"0C",X"00",X"ED",X"B0",
		X"21",X"00",X"00",X"01",X"00",X"0A",X"11",X"F4",X"03",X"79",X"86",X"4F",X"3A",X"00",X"B8",X"2C",
		X"20",X"F7",X"24",X"3E",X"07",X"A4",X"20",X"F1",X"1A",X"B9",X"00",X"00",X"0E",X"00",X"13",X"10",
		X"E8",X"C3",X"74",X"05",X"0C",X"6A",X"29",X"F3",X"DC",X"B6",X"FD",X"44",X"63",X"D5",X"F4",X"D9",
		X"21",X"C4",X"03",X"11",X"A6",X"90",X"01",X"06",X"00",X"ED",X"B0",X"D9",X"EB",X"21",X"B0",X"90",
		X"3E",X"F8",X"A2",X"0F",X"0F",X"0F",X"77",X"79",X"D9",X"21",X"BA",X"90",X"D9",X"21",X"23",X"04",
		X"C3",X"9F",X"03",X"00",X"00",X"00",X"00",X"3A",X"00",X"B8",X"1A",X"18",X"FA",X"E6",X"1F",X"5F",
		X"21",X"70",X"04",X"06",X"0D",X"BE",X"28",X"07",X"23",X"23",X"10",X"F9",X"37",X"18",X"25",X"23",
		X"7E",X"06",X"01",X"B7",X"28",X"01",X"47",X"7B",X"CD",X"AB",X"04",X"CB",X"7E",X"28",X"06",X"1C",
		X"10",X"F5",X"37",X"18",X"0F",X"73",X"CB",X"FE",X"23",X"36",X"00",X"01",X"0E",X"00",X"54",X"5D",
		X"13",X"ED",X"B0",X"B7",X"C1",X"D1",X"E1",X"C1",X"C9",X"C1",X"D1",X"E1",X"E3",X"7C",X"E1",X"C9",
		X"00",X"00",X"01",X"00",X"02",X"00",X"03",X"03",X"06",X"03",X"09",X"03",X"0C",X"00",X"0D",X"00",
		X"0E",X"00",X"0F",X"00",X"10",X"03",X"13",X"00",X"14",X"00",X"E6",X"1F",X"5F",X"CD",X"AB",X"04",
		X"CB",X"BE",X"CB",X"F6",X"7B",X"D5",X"CD",X"31",X"06",X"D1",X"CB",X"76",X"28",X"F4",X"36",X"00",
		X"4B",X"21",X"47",X"82",X"06",X"08",X"CD",X"06",X"02",X"18",X"BE",X"21",X"00",X"B8",X"BE",X"21",
		X"00",X"80",X"BE",X"21",X"2F",X"80",X"C8",X"26",X"00",X"D5",X"6F",X"29",X"29",X"29",X"29",X"11",
		X"3F",X"80",X"19",X"D1",X"C9",X"C5",X"D5",X"AF",X"ED",X"A0",X"B1",X"20",X"FA",X"3A",X"00",X"B8",
		X"11",X"20",X"00",X"E3",X"19",X"EB",X"E1",X"C1",X"10",X"EB",X"C9",X"C5",X"D5",X"AF",X"ED",X"A0",
		X"B1",X"20",X"FA",X"3A",X"00",X"B8",X"11",X"10",X"00",X"E3",X"19",X"EB",X"E1",X"C1",X"10",X"EB",
		X"C9",X"C5",X"D5",X"12",X"13",X"0D",X"20",X"FB",X"21",X"00",X"B8",X"BE",X"11",X"20",X"00",X"E1",
		X"19",X"EB",X"C1",X"10",X"EC",X"C9",X"E5",X"62",X"6B",X"13",X"0B",X"77",X"ED",X"B0",X"E1",X"3A",
		X"00",X"B8",X"C9",X"E5",X"EB",X"1E",X"20",X"57",X"7A",X"77",X"16",X"00",X"19",X"57",X"0B",X"78",
		X"B1",X"20",X"F5",X"E1",X"3A",X"00",X"B8",X"C9",X"06",X"05",X"1A",X"BE",X"C0",X"23",X"13",X"10",
		X"F9",X"C9",X"CB",X"D2",X"CB",X"DA",X"CD",X"F1",X"04",X"C9",X"E6",X"1F",X"06",X"00",X"4F",X"EB",
		X"21",X"31",X"82",X"09",X"34",X"06",X"28",X"21",X"B9",X"81",X"7E",X"B7",X"28",X"09",X"23",X"23",
		X"23",X"10",X"F7",X"37",X"C3",X"69",X"04",X"71",X"23",X"73",X"23",X"72",X"C3",X"69",X"04",X"E6",
		X"1F",X"CD",X"AB",X"04",X"CB",X"F6",X"C3",X"69",X"04",X"2A",X"09",X"80",X"7C",X"B5",X"C8",X"3A",
		X"00",X"B8",X"18",X"F5",X"31",X"00",X"84",X"AF",X"32",X"07",X"A0",X"3E",X"07",X"D3",X"08",X"3E",
		X"3F",X"D3",X"09",X"11",X"00",X"90",X"3E",X"24",X"CD",X"76",X"08",X"11",X"00",X"9C",X"3E",X"00",
		X"CD",X"76",X"08",X"21",X"00",X"80",X"3E",X"00",X"01",X"F0",X"04",X"CD",X"79",X"08",X"11",X"00",
		X"98",X"3E",X"00",X"CD",X"76",X"08",X"11",X"00",X"88",X"3E",X"FF",X"CD",X"76",X"08",X"3E",X"3F",
		X"32",X"A0",X"81",X"3E",X"FF",X"32",X"00",X"80",X"21",X"7C",X"02",X"22",X"0B",X"80",X"21",X"85",
		X"02",X"22",X"0D",X"80",X"21",X"2F",X"80",X"22",X"07",X"80",X"3E",X"81",X"32",X"14",X"80",X"3E",
		X"00",X"CF",X"3E",X"01",X"32",X"00",X"A0",X"01",X"10",X"00",X"09",X"EB",X"21",X"00",X"80",X"34",
		X"7E",X"FE",X"15",X"20",X"05",X"36",X"00",X"11",X"3F",X"80",X"3A",X"00",X"B8",X"EB",X"CB",X"7E",
		X"28",X"E5",X"22",X"07",X"80",X"CB",X"76",X"3A",X"00",X"80",X"C4",X"31",X"06",X"CB",X"76",X"20",
		X"D6",X"11",X"2F",X"80",X"01",X"10",X"00",X"ED",X"B0",X"26",X"00",X"3A",X"00",X"80",X"87",X"6F",
		X"01",X"63",X"06",X"09",X"5E",X"23",X"56",X"EB",X"01",X"1D",X"06",X"C5",X"E9",X"3A",X"00",X"B8",
		X"11",X"2F",X"80",X"2A",X"07",X"80",X"01",X"10",X"00",X"EB",X"ED",X"B0",X"2A",X"07",X"80",X"18",
		X"A6",X"E5",X"EB",X"21",X"31",X"82",X"06",X"00",X"4F",X"09",X"7E",X"B7",X"28",X"23",X"35",X"06",
		X"28",X"21",X"B9",X"81",X"79",X"BE",X"20",X"14",X"1A",X"E6",X"9F",X"12",X"36",X"00",X"23",X"13",
		X"7E",X"36",X"00",X"12",X"23",X"13",X"7E",X"36",X"00",X"12",X"18",X"05",X"23",X"23",X"23",X"10",
		X"E4",X"E1",X"C9",X"8D",X"06",X"6D",X"35",X"6F",X"0F",X"3D",X"3D",X"3D",X"3D",X"3D",X"3D",X"6B",
		X"42",X"6B",X"42",X"6B",X"42",X"6B",X"42",X"6B",X"42",X"6B",X"42",X"9F",X"34",X"BC",X"33",X"12",
		X"33",X"68",X"3F",X"CD",X"44",X"CD",X"44",X"CD",X"44",X"6E",X"46",X"7F",X"0A",X"21",X"32",X"80",
		X"CB",X"7E",X"C2",X"26",X"07",X"CB",X"FE",X"21",X"00",X"00",X"22",X"BC",X"93",X"01",X"00",X"12",
		X"C5",X"79",X"CD",X"12",X"0D",X"C1",X"0C",X"10",X"F7",X"3E",X"E4",X"11",X"A1",X"90",X"01",X"18",
		X"00",X"00",X"00",X"00",X"3E",X"08",X"11",X"A1",X"90",X"01",X"01",X"18",X"00",X"00",X"00",X"3E",
		X"E4",X"11",X"A2",X"90",X"01",X"18",X"00",X"C3",X"00",X"52",X"3E",X"09",X"11",X"A2",X"90",X"01",
		X"01",X"18",X"CD",X"32",X"05",X"3A",X"00",X"B0",X"E6",X"0C",X"0F",X"0F",X"C6",X"03",X"32",X"01",
		X"80",X"3A",X"00",X"B0",X"E6",X"03",X"21",X"02",X"80",X"36",X"00",X"FE",X"03",X"28",X"0E",X"36",
		X"04",X"FE",X"02",X"28",X"08",X"36",X"01",X"FE",X"01",X"28",X"02",X"36",X"02",X"3E",X"FF",X"32",
		X"13",X"80",X"3E",X"81",X"32",X"14",X"80",X"3E",X"00",X"CD",X"12",X"0D",X"3A",X"16",X"80",X"CB",
		X"7F",X"28",X"05",X"3E",X"02",X"CD",X"12",X"0D",X"AF",X"32",X"01",X"A0",X"32",X"02",X"A0",X"32",
		X"15",X"80",X"3E",X"14",X"CF",X"C9",X"21",X"14",X"80",X"CB",X"7E",X"28",X"33",X"3A",X"03",X"80",
		X"21",X"02",X"80",X"BE",X"3E",X"03",X"38",X"28",X"32",X"15",X"80",X"21",X"14",X"80",X"CB",X"BE",
		X"21",X"7C",X"02",X"22",X"0B",X"80",X"21",X"85",X"02",X"22",X"0D",X"80",X"21",X"0F",X"80",X"36",
		X"00",X"23",X"36",X"00",X"06",X"14",X"3E",X"01",X"D7",X"3C",X"10",X"FC",X"3E",X"14",X"CF",X"C9",
		X"3A",X"15",X"80",X"FE",X"05",X"20",X"0D",X"3A",X"00",X"B8",X"3A",X"06",X"80",X"B7",X"28",X"F0",
		X"3D",X"32",X"06",X"80",X"21",X"14",X"80",X"7E",X"E6",X"60",X"C8",X"EB",X"21",X"7C",X"02",X"22",
		X"0B",X"80",X"21",X"85",X"02",X"22",X"0D",X"80",X"21",X"0F",X"80",X"36",X"00",X"23",X"36",X"00",
		X"06",X"14",X"3E",X"01",X"D7",X"3C",X"10",X"FC",X"EB",X"CB",X"7E",X"C2",X"FD",X"06",X"CB",X"76",
		X"20",X"16",X"CB",X"AE",X"21",X"17",X"80",X"3A",X"16",X"80",X"CB",X"77",X"28",X"01",X"23",X"7E",
		X"C6",X"01",X"27",X"77",X"3E",X"05",X"18",X"80",X"CB",X"B6",X"3A",X"16",X"80",X"21",X"19",X"80",
		X"01",X"10",X"20",X"CB",X"77",X"28",X"04",X"01",X"20",X"10",X"23",X"7E",X"B7",X"20",X"1B",X"C5",
		X"CD",X"0D",X"08",X"3E",X"21",X"CD",X"12",X"0D",X"21",X"64",X"00",X"F7",X"C1",X"21",X"16",X"80",
		X"7E",X"B0",X"77",X"E6",X"30",X"FE",X"30",X"CA",X"8A",X"08",X"21",X"16",X"80",X"7E",X"EE",X"40",
		X"47",X"A1",X"20",X"14",X"70",X"78",X"07",X"07",X"E6",X"01",X"21",X"00",X"B0",X"CB",X"66",X"28",
		X"01",X"AF",X"32",X"01",X"A0",X"32",X"02",X"A0",X"3E",X"04",X"C3",X"38",X"07",X"3A",X"00",X"B8",
		X"21",X"00",X"88",X"11",X"01",X"88",X"01",X"FF",X"00",X"36",X"FF",X"ED",X"B0",X"3A",X"00",X"B8",
		X"21",X"00",X"98",X"11",X"01",X"98",X"01",X"1F",X"00",X"36",X"00",X"ED",X"B0",X"3A",X"00",X"B8",
		X"3E",X"00",X"11",X"04",X"90",X"01",X"16",X"20",X"CD",X"32",X"05",X"11",X"04",X"90",X"01",X"16",
		X"20",X"3E",X"24",X"CD",X"F1",X"04",X"3A",X"00",X"B8",X"3E",X"E4",X"11",X"A1",X"90",X"01",X"18",
		X"00",X"00",X"00",X"00",X"3E",X"08",X"11",X"A1",X"90",X"01",X"01",X"18",X"00",X"00",X"00",X"3E",
		X"E4",X"11",X"A2",X"90",X"01",X"18",X"00",X"CD",X"13",X"05",X"3E",X"09",X"11",X"A2",X"90",X"01",
		X"01",X"18",X"CD",X"32",X"05",X"C9",X"01",X"FF",X"03",X"62",X"6B",X"77",X"13",X"ED",X"A0",X"AF",
		X"B1",X"20",X"FA",X"B0",X"C8",X"3A",X"00",X"B8",X"18",X"F3",X"CD",X"0D",X"08",X"AF",X"32",X"01",
		X"A0",X"32",X"02",X"A0",X"21",X"2B",X"80",X"7E",X"B7",X"CA",X"2A",X"09",X"32",X"39",X"80",X"11",
		X"00",X"A8",X"21",X"34",X"80",X"CB",X"46",X"28",X"03",X"11",X"00",X"A0",X"ED",X"53",X"37",X"80",
		X"21",X"00",X"F0",X"22",X"3D",X"80",X"01",X"10",X"00",X"11",X"67",X"91",X"21",X"59",X"0A",X"ED",
		X"B0",X"01",X"10",X"00",X"11",X"07",X"92",X"21",X"69",X"0A",X"ED",X"B0",X"3A",X"39",X"80",X"FE",
		X"01",X"20",X"05",X"11",X"9B",X"92",X"18",X"0C",X"FE",X"02",X"20",X"05",X"11",X"1B",X"92",X"18",
		X"03",X"11",X"9B",X"91",X"ED",X"53",X"35",X"80",X"3E",X"25",X"12",X"21",X"6E",X"92",X"3E",X"0A",
		X"77",X"2A",X"3D",X"80",X"23",X"22",X"3D",X"80",X"CD",X"6A",X"09",X"3A",X"34",X"80",X"CB",X"5F",
		X"20",X"28",X"2A",X"3D",X"80",X"7C",X"B5",X"28",X"21",X"21",X"3A",X"80",X"34",X"7E",X"E6",X"0F",
		X"20",X"DF",X"21",X"34",X"80",X"CB",X"4E",X"20",X"06",X"CB",X"CE",X"3E",X"24",X"18",X"04",X"CB",
		X"8E",X"3E",X"25",X"ED",X"5B",X"35",X"80",X"12",X"18",X"C7",X"21",X"34",X"80",X"CB",X"46",X"20",
		X"29",X"CB",X"C6",X"01",X"09",X"00",X"21",X"35",X"80",X"11",X"36",X"80",X"36",X"00",X"ED",X"B0",
		X"21",X"34",X"80",X"CB",X"9E",X"21",X"00",X"B0",X"CB",X"66",X"20",X"08",X"3E",X"01",X"32",X"01",
		X"A0",X"32",X"02",X"A0",X"21",X"2C",X"80",X"C3",X"97",X"08",X"01",X"0A",X"00",X"11",X"35",X"80",
		X"21",X"34",X"80",X"36",X"00",X"ED",X"B0",X"C3",X"FD",X"06",X"3A",X"00",X"B8",X"3A",X"03",X"80",
		X"B7",X"28",X"07",X"3A",X"00",X"B8",X"E6",X"0C",X"20",X"3D",X"21",X"3B",X"80",X"34",X"20",X"EA",
		X"2A",X"37",X"80",X"7E",X"CB",X"47",X"28",X"52",X"21",X"34",X"80",X"CB",X"7E",X"C0",X"CB",X"FE",
		X"3A",X"3C",X"80",X"FE",X"1C",X"28",X"20",X"FE",X"1B",X"28",X"28",X"FE",X"1A",X"28",X"08",X"C6",
		X"0A",X"2A",X"35",X"80",X"77",X"18",X"06",X"3E",X"26",X"2A",X"35",X"80",X"77",X"23",X"7E",X"FE",
		X"28",X"28",X"0A",X"22",X"35",X"80",X"C9",X"3E",X"24",X"2A",X"35",X"80",X"77",X"21",X"34",X"80",
		X"CB",X"DE",X"C9",X"2A",X"35",X"80",X"2B",X"7E",X"FE",X"27",X"20",X"03",X"23",X"18",X"03",X"3E",
		X"24",X"77",X"22",X"35",X"80",X"23",X"3E",X"24",X"77",X"C9",X"21",X"34",X"80",X"CB",X"BE",X"21",
		X"3C",X"80",X"CB",X"77",X"20",X"05",X"CB",X"7F",X"20",X"0B",X"C9",X"34",X"7E",X"FE",X"1D",X"20",
		X"0B",X"AF",X"77",X"18",X"07",X"35",X"CB",X"7E",X"28",X"02",X"36",X"1C",X"E5",X"21",X"3B",X"80",
		X"E5",X"21",X"01",X"00",X"F7",X"E1",X"34",X"3A",X"00",X"B8",X"7E",X"E6",X"0F",X"20",X"F1",X"36",
		X"00",X"3E",X"24",X"11",X"6E",X"92",X"01",X"03",X"00",X"CD",X"06",X"05",X"E1",X"7E",X"FE",X"1B",
		X"28",X"13",X"30",X"16",X"FE",X"1A",X"28",X"24",X"C6",X"0A",X"21",X"6E",X"92",X"77",X"21",X"00",
		X"F0",X"22",X"3D",X"80",X"C9",X"21",X"79",X"0A",X"18",X"03",X"21",X"7C",X"0A",X"11",X"6E",X"92",
		X"01",X"03",X"00",X"ED",X"B0",X"21",X"00",X"F0",X"22",X"3D",X"80",X"C9",X"3E",X"26",X"21",X"6E",
		X"92",X"77",X"21",X"00",X"F0",X"22",X"3D",X"80",X"C9",X"17",X"0A",X"16",X"0E",X"24",X"1B",X"0E",
		X"10",X"12",X"1C",X"1D",X"0A",X"1D",X"12",X"18",X"17",X"1C",X"0E",X"15",X"0E",X"0C",X"1D",X"24",
		X"0C",X"11",X"0A",X"1B",X"0A",X"0C",X"1D",X"0E",X"1B",X"1B",X"1E",X"0B",X"0E",X"17",X"0D",X"21",
		X"15",X"80",X"7E",X"FE",X"00",X"C2",X"B2",X"0A",X"CD",X"0D",X"08",X"01",X"19",X"00",X"21",X"15",
		X"80",X"11",X"16",X"80",X"36",X"00",X"ED",X"B0",X"21",X"01",X"01",X"22",X"17",X"80",X"3A",X"01",
		X"80",X"32",X"19",X"80",X"32",X"1A",X"80",X"CD",X"DC",X"0C",X"21",X"15",X"80",X"34",X"23",X"36",
		X"30",X"C9",X"7E",X"FE",X"01",X"C2",X"3A",X"0B",X"21",X"32",X"80",X"7E",X"34",X"B7",X"20",X"4F",
		X"CD",X"0D",X"08",X"01",X"13",X"06",X"21",X"5A",X"0C",X"11",X"86",X"90",X"CD",X"C5",X"04",X"01",
		X"13",X"06",X"11",X"86",X"90",X"3E",X"12",X"CD",X"32",X"05",X"3E",X"15",X"CD",X"12",X"0D",X"3E",
		X"16",X"CD",X"12",X"0D",X"3E",X"17",X"CD",X"12",X"0D",X"01",X"04",X"04",X"21",X"CC",X"0C",X"11",
		X"4C",X"92",X"CD",X"C5",X"04",X"11",X"4C",X"92",X"3E",X"10",X"01",X"04",X"04",X"CD",X"32",X"05",
		X"3E",X"18",X"CD",X"12",X"0D",X"3E",X"19",X"CD",X"12",X"0D",X"21",X"32",X"00",X"F7",X"C9",X"7E",
		X"FE",X"08",X"28",X"1E",X"CB",X"47",X"20",X"0A",X"3E",X"15",X"CD",X"12",X"0D",X"21",X"32",X"00",
		X"F7",X"C9",X"3E",X"24",X"11",X"49",X"91",X"01",X"0B",X"00",X"CD",X"06",X"05",X"21",X"32",X"00",
		X"F7",X"C9",X"36",X"00",X"21",X"15",X"80",X"36",X"05",X"C9",X"FE",X"03",X"C2",X"BB",X"0B",X"21",
		X"32",X"80",X"7E",X"B7",X"20",X"0F",X"36",X"01",X"CD",X"0D",X"08",X"3E",X"1D",X"CD",X"12",X"0D",
		X"3E",X"20",X"CD",X"12",X"0D",X"3A",X"03",X"80",X"21",X"02",X"80",X"4E",X"B7",X"CB",X"11",X"B9",
		X"30",X"1F",X"3E",X"1E",X"CD",X"12",X"0D",X"3A",X"00",X"B8",X"CB",X"57",X"C8",X"3A",X"03",X"80",
		X"21",X"02",X"80",X"96",X"32",X"03",X"80",X"CD",X"07",X"01",X"21",X"16",X"80",X"36",X"10",X"18",
		X"22",X"3E",X"1F",X"CD",X"12",X"0D",X"3A",X"00",X"B8",X"CB",X"57",X"20",X"E0",X"CB",X"5F",X"C8",
		X"3A",X"03",X"80",X"21",X"02",X"80",X"96",X"96",X"32",X"03",X"80",X"CD",X"07",X"01",X"21",X"16",
		X"80",X"36",X"80",X"21",X"2E",X"80",X"36",X"00",X"3A",X"01",X"80",X"67",X"6F",X"22",X"19",X"80",
		X"21",X"01",X"01",X"22",X"17",X"80",X"21",X"15",X"80",X"34",X"C9",X"FE",X"04",X"20",X"1B",X"CD",
		X"0D",X"08",X"21",X"16",X"80",X"3E",X"1B",X"CB",X"76",X"28",X"02",X"3E",X"1C",X"CD",X"12",X"0D",
		X"3E",X"1A",X"CD",X"12",X"0D",X"21",X"15",X"80",X"34",X"C9",X"FE",X"05",X"C0",X"CD",X"DC",X"0C",
		X"21",X"C8",X"00",X"F7",X"21",X"14",X"80",X"CB",X"C6",X"CB",X"96",X"23",X"23",X"7E",X"E6",X"F0",
		X"77",X"CD",X"0D",X"08",X"21",X"14",X"80",X"CB",X"7E",X"20",X"16",X"3E",X"13",X"CD",X"12",X"0D",
		X"3E",X"00",X"CD",X"12",X"0D",X"3A",X"16",X"80",X"CB",X"7F",X"28",X"05",X"3E",X"02",X"CD",X"12",
		X"0D",X"AF",X"32",X"A1",X"81",X"32",X"A9",X"81",X"32",X"B1",X"81",X"32",X"9F",X"81",X"CD",X"DC",
		X"0C",X"3E",X"07",X"D3",X"08",X"3E",X"3F",X"32",X"A0",X"81",X"D3",X"09",X"3E",X"14",X"D7",X"3E",
		X"01",X"CF",X"3E",X"02",X"CF",X"3E",X"0E",X"CF",X"3E",X"0D",X"CF",X"3E",X"0F",X"CF",X"21",X"14",
		X"80",X"CB",X"7E",X"C0",X"3E",X"13",X"CD",X"12",X"0D",X"3E",X"00",X"CD",X"12",X"0D",X"3A",X"16",
		X"80",X"CB",X"7F",X"C8",X"3E",X"02",X"CD",X"12",X"0D",X"C9",X"91",X"92",X"93",X"94",X"95",X"96",
		X"97",X"98",X"99",X"9A",X"9B",X"9C",X"9D",X"9E",X"9F",X"A0",X"A1",X"A2",X"A3",X"A4",X"A5",X"A6",
		X"A7",X"A8",X"A9",X"AA",X"AB",X"AC",X"AD",X"AE",X"AF",X"B0",X"B1",X"B2",X"B3",X"B4",X"B5",X"B6",
		X"B7",X"B8",X"B9",X"BA",X"BB",X"BC",X"BD",X"BE",X"BF",X"C0",X"C1",X"C2",X"C3",X"C4",X"C5",X"C6",
		X"C7",X"C8",X"C9",X"CA",X"CB",X"CC",X"CD",X"CE",X"CF",X"D0",X"D1",X"D2",X"D3",X"D4",X"D5",X"D6",
		X"D7",X"D8",X"D9",X"DA",X"DB",X"DC",X"DD",X"DE",X"DF",X"E0",X"E1",X"E2",X"E3",X"E4",X"E5",X"E6",
		X"E7",X"E8",X"E9",X"EA",X"EB",X"EC",X"ED",X"EE",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"75",X"76",X"77",X"78",
		X"79",X"7A",X"7B",X"7C",X"7D",X"7E",X"7F",X"80",X"81",X"82",X"83",X"84",X"21",X"5B",X"93",X"36",
		X"85",X"11",X"20",X"00",X"19",X"36",X"FF",X"11",X"00",X"0C",X"19",X"36",X"10",X"21",X"5D",X"93",
		X"11",X"19",X"80",X"01",X"17",X"80",X"3A",X"16",X"80",X"CB",X"77",X"28",X"02",X"13",X"03",X"1A",
		X"77",X"0A",X"21",X"1C",X"93",X"E6",X"F0",X"0F",X"0F",X"0F",X"0F",X"77",X"23",X"0A",X"E6",X"0F",
		X"77",X"C9",X"21",X"4F",X"0D",X"16",X"00",X"87",X"5F",X"87",X"83",X"5F",X"19",X"46",X"23",X"4E",
		X"C5",X"23",X"4E",X"23",X"46",X"23",X"5E",X"23",X"56",X"60",X"69",X"C1",X"7E",X"FE",X"FF",X"C8",
		X"12",X"3A",X"00",X"B8",X"23",X"E5",X"CB",X"D2",X"CB",X"DA",X"EB",X"71",X"EB",X"CB",X"92",X"CB",
		X"9A",X"21",X"20",X"00",X"CB",X"40",X"20",X"02",X"2E",X"01",X"19",X"EB",X"E1",X"18",X"DD",X"00",
		X"00",X"27",X"0E",X"7B",X"90",X"00",X"00",X"2B",X"0E",X"BA",X"90",X"00",X"00",X"32",X"0E",X"FB",
		X"90",X"00",X"00",X"2B",X"0E",X"3A",X"91",X"00",X"00",X"36",X"0E",X"7B",X"91",X"00",X"00",X"3A",
		X"0E",X"9A",X"91",X"00",X"00",X"41",X"0E",X"BA",X"91",X"00",X"00",X"48",X"0E",X"FB",X"91",X"00",
		X"00",X"3A",X"0E",X"1A",X"92",X"00",X"00",X"41",X"0E",X"3A",X"92",X"00",X"00",X"4C",X"0E",X"7B",
		X"92",X"00",X"00",X"3A",X"0E",X"9A",X"92",X"00",X"00",X"41",X"0E",X"BA",X"92",X"00",X"00",X"50",
		X"0E",X"FA",X"92",X"00",X"00",X"57",X"0E",X"1B",X"93",X"00",X"00",X"5C",X"0E",X"9A",X"93",X"01",
		X"00",X"63",X"0E",X"40",X"91",X"01",X"00",X"6E",X"0E",X"42",X"91",X"00",X"00",X"7A",X"0E",X"7B",
		X"90",X"00",X"00",X"7A",X"0E",X"FB",X"90",X"00",X"00",X"7E",X"0E",X"BB",X"93",X"00",X"00",X"83",
		X"0E",X"49",X"91",X"00",X"00",X"8F",X"0E",X"85",X"91",X"00",X"00",X"A4",X"0E",X"C5",X"91",X"00",
		X"00",X"BA",X"0E",X"29",X"93",X"00",X"00",X"CA",X"0E",X"65",X"93",X"00",X"00",X"E0",X"0E",X"0A",
		X"92",X"00",X"00",X"EB",X"0E",X"28",X"91",X"00",X"00",X"FC",X"0E",X"28",X"91",X"00",X"00",X"0D",
		X"0F",X"4D",X"91",X"00",X"00",X"12",X"0F",X"87",X"91",X"00",X"00",X"22",X"0F",X"86",X"91",X"00",
		X"00",X"34",X"0F",X"C8",X"91",X"00",X"00",X"41",X"0F",X"CB",X"91",X"00",X"00",X"4B",X"0F",X"68",
		X"91",X"00",X"00",X"5B",X"0F",X"A6",X"91",X"01",X"1E",X"19",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"02",X"1E",X"19",X"FF",X"1D",X"18",X"19",X"FF",X"27",X"0F",X"0A",X"15",X"26",X"28",
		X"FF",X"00",X"01",X"00",X"00",X"00",X"00",X"FF",X"02",X"17",X"0D",X"FF",X"03",X"1B",X"0D",X"FF",
		X"1B",X"18",X"1E",X"17",X"0D",X"1C",X"FF",X"27",X"00",X"01",X"28",X"FF",X"0C",X"1B",X"0E",X"0D",
		X"12",X"1D",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"24",X"24",X"24",X"FF",X"0F",X"1B",
		X"0E",X"0E",X"FF",X"12",X"17",X"1C",X"0E",X"1B",X"1D",X"24",X"0C",X"18",X"12",X"17",X"FF",X"24",
		X"24",X"01",X"24",X"0C",X"18",X"12",X"17",X"24",X"24",X"24",X"24",X"01",X"24",X"19",X"15",X"0A",
		X"22",X"0E",X"1B",X"FF",X"24",X"24",X"02",X"24",X"0C",X"18",X"12",X"17",X"1C",X"24",X"24",X"24",
		X"02",X"24",X"19",X"15",X"0A",X"22",X"0E",X"1B",X"1C",X"FF",X"24",X"24",X"24",X"24",X"24",X"24",
		X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"FF",X"24",X"24",X"24",X"24",X"24",X"24",
		X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"FF",
		X"10",X"18",X"18",X"0D",X"24",X"24",X"15",X"1E",X"0C",X"14",X"FF",X"19",X"15",X"0A",X"22",X"0E",
		X"1B",X"24",X"18",X"17",X"0E",X"24",X"1C",X"1D",X"0A",X"1B",X"1D",X"FF",X"19",X"15",X"0A",X"22",
		X"0E",X"1B",X"24",X"1D",X"20",X"18",X"24",X"1C",X"1D",X"0A",X"1B",X"1D",X"FF",X"19",X"1E",X"1C",
		X"11",X"FF",X"18",X"17",X"15",X"22",X"24",X"18",X"17",X"0E",X"24",X"19",X"15",X"0A",X"22",X"0E",
		X"1B",X"FF",X"18",X"17",X"0E",X"24",X"18",X"1B",X"24",X"1D",X"20",X"18",X"24",X"19",X"15",X"0A",
		X"22",X"0E",X"1B",X"FF",X"1C",X"1D",X"0A",X"1B",X"1D",X"24",X"0B",X"1E",X"1D",X"1D",X"18",X"17",
		X"FF",X"10",X"0A",X"16",X"0E",X"24",X"18",X"1F",X"0E",X"1B",X"FF",X"24",X"24",X"24",X"24",X"24",
		X"10",X"18",X"0A",X"15",X"24",X"24",X"24",X"24",X"24",X"24",X"FF",X"24",X"24",X"24",X"24",X"24",
		X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"FF",X"21",
		X"32",X"80",X"CB",X"7E",X"C2",X"45",X"10",X"CB",X"FE",X"CB",X"EE",X"21",X"17",X"80",X"3A",X"16",
		X"80",X"CB",X"77",X"28",X"01",X"23",X"3A",X"14",X"80",X"CB",X"7F",X"3E",X"0A",X"20",X"07",X"7E",
		X"FE",X"0A",X"38",X"02",X"3E",X"0A",X"3D",X"0F",X"E6",X"7F",X"32",X"33",X"80",X"32",X"28",X"80",
		X"ED",X"44",X"C6",X"A8",X"32",X"29",X"80",X"3A",X"14",X"80",X"CB",X"7F",X"11",X"BC",X"31",X"20",
		X"2A",X"7E",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"28",X"06",X"47",X"AF",X"C6",X"0A",X"10",X"FC",
		X"47",X"7E",X"E6",X"0F",X"80",X"FE",X"11",X"38",X"04",X"D6",X"07",X"18",X"F8",X"3D",X"E6",X"0F",
		X"6F",X"26",X"00",X"29",X"11",X"0C",X"13",X"19",X"5E",X"23",X"56",X"ED",X"53",X"38",X"80",X"11",
		X"04",X"90",X"01",X"16",X"20",X"3E",X"35",X"CD",X"F1",X"04",X"11",X"04",X"9C",X"01",X"16",X"20",
		X"3E",X"1E",X"CD",X"F1",X"04",X"ED",X"5F",X"E6",X"03",X"28",X"02",X"EE",X"03",X"07",X"07",X"C6",
		X"00",X"32",X"3C",X"80",X"21",X"00",X"00",X"22",X"3D",X"80",X"01",X"00",X"20",X"11",X"04",X"90",
		X"21",X"19",X"90",X"C5",X"06",X"00",X"79",X"E6",X"0F",X"4F",X"DD",X"21",X"85",X"12",X"DD",X"09",
		X"DD",X"7E",X"00",X"12",X"77",X"CB",X"D4",X"CB",X"DC",X"36",X"5E",X"CB",X"94",X"CB",X"9C",X"EB",
		X"CB",X"D4",X"CB",X"DC",X"36",X"1E",X"CB",X"94",X"CB",X"9C",X"01",X"20",X"00",X"09",X"EB",X"09",
		X"C1",X"0C",X"10",X"CF",X"C9",X"3A",X"21",X"80",X"21",X"36",X"80",X"96",X"21",X"32",X"80",X"CA",
		X"E8",X"10",X"FA",X"71",X"10",X"CB",X"EE",X"CD",X"F8",X"12",X"2A",X"21",X"80",X"11",X"E0",X"00",
		X"19",X"22",X"3A",X"80",X"45",X"2A",X"21",X"80",X"B7",X"ED",X"52",X"68",X"38",X"14",X"68",X"18",
		X"11",X"CB",X"AE",X"CD",X"F8",X"12",X"2A",X"21",X"80",X"11",X"08",X"00",X"B7",X"ED",X"52",X"22",
		X"3A",X"80",X"3A",X"3A",X"80",X"E6",X"07",X"20",X"5F",X"26",X"00",X"CD",X"46",X"46",X"ED",X"53",
		X"34",X"80",X"01",X"16",X"00",X"3E",X"35",X"CD",X"06",X"05",X"ED",X"5B",X"34",X"80",X"01",X"16",
		X"01",X"3E",X"1E",X"CD",X"32",X"05",X"16",X"00",X"3A",X"3A",X"80",X"E6",X"78",X"0F",X"0F",X"0F",
		X"5F",X"21",X"85",X"12",X"19",X"4E",X"2A",X"34",X"80",X"3A",X"33",X"80",X"B7",X"47",X"28",X"05",
		X"36",X"34",X"23",X"10",X"FB",X"71",X"C5",X"11",X"15",X"0C",X"2A",X"34",X"80",X"19",X"EB",X"2A",
		X"34",X"80",X"01",X"15",X"00",X"09",X"C1",X"3A",X"33",X"80",X"B7",X"28",X"07",X"47",X"36",X"34",
		X"2B",X"1B",X"10",X"FA",X"71",X"EB",X"36",X"5E",X"21",X"30",X"80",X"34",X"3E",X"03",X"A6",X"20",
		X"32",X"3A",X"1F",X"80",X"6F",X"3A",X"33",X"80",X"07",X"07",X"07",X"D6",X"06",X"67",X"01",X"08",
		X"20",X"C5",X"CD",X"D0",X"3E",X"C1",X"38",X"16",X"3A",X"33",X"80",X"ED",X"44",X"C6",X"15",X"07",
		X"07",X"07",X"C6",X"06",X"67",X"3A",X"1F",X"80",X"6F",X"CD",X"D0",X"3E",X"30",X"05",X"21",X"16",
		X"80",X"CB",X"DE",X"21",X"36",X"80",X"3A",X"21",X"80",X"BE",X"C8",X"77",X"2A",X"3D",X"80",X"ED",
		X"5B",X"3A",X"80",X"B7",X"ED",X"52",X"30",X"04",X"ED",X"53",X"3D",X"80",X"3A",X"3A",X"80",X"E6",
		X"07",X"C0",X"21",X"32",X"80",X"CB",X"66",X"C2",X"DB",X"11",X"CD",X"95",X"12",X"11",X"C0",X"0E",
		X"2A",X"21",X"80",X"B7",X"ED",X"52",X"38",X"0D",X"21",X"32",X"80",X"CB",X"E6",X"21",X"14",X"80",
		X"CB",X"D6",X"C3",X"DB",X"11",X"CD",X"C2",X"12",X"D8",X"DD",X"7E",X"01",X"E6",X"F8",X"0F",X"0F",
		X"0F",X"FE",X"00",X"20",X"2C",X"DD",X"7E",X"02",X"E6",X"1F",X"5F",X"16",X"00",X"2A",X"34",X"80",
		X"19",X"DD",X"7E",X"02",X"E6",X"E0",X"07",X"07",X"07",X"47",X"3A",X"3C",X"80",X"57",X"3A",X"3A",
		X"80",X"CB",X"5F",X"20",X"02",X"14",X"14",X"7A",X"77",X"23",X"3C",X"77",X"23",X"10",X"F8",X"18",
		X"C4",X"2A",X"3D",X"80",X"ED",X"5B",X"3A",X"80",X"B7",X"ED",X"52",X"28",X"02",X"30",X"B6",X"21",
		X"32",X"80",X"CB",X"6E",X"28",X"AF",X"21",X"3A",X"80",X"CB",X"5E",X"20",X"A8",X"FE",X"13",X"20",
		X"07",X"21",X"16",X"80",X"CB",X"56",X"20",X"9D",X"CF",X"38",X"9A",X"2E",X"E0",X"F5",X"DD",X"7E",
		X"02",X"E6",X"1F",X"07",X"07",X"07",X"67",X"F1",X"E7",X"18",X"8A",X"2A",X"21",X"80",X"11",X"C0",
		X"0E",X"B7",X"ED",X"52",X"3E",X"F8",X"A5",X"0F",X"0F",X"FE",X"10",X"D0",X"6F",X"11",X"1D",X"12",
		X"19",X"5E",X"23",X"56",X"2A",X"34",X"80",X"06",X"0B",X"1A",X"77",X"13",X"23",X"10",X"FA",X"06",
		X"0B",X"1B",X"1A",X"77",X"23",X"10",X"FA",X"11",X"00",X"0C",X"2A",X"34",X"80",X"19",X"06",X"0B",
		X"36",X"1E",X"23",X"10",X"FB",X"06",X"0B",X"36",X"5E",X"23",X"10",X"FB",X"C9",X"2D",X"12",X"2D",
		X"12",X"2D",X"12",X"2D",X"12",X"2D",X"12",X"2D",X"12",X"2D",X"12",X"2D",X"12",X"35",X"35",X"35",
		X"35",X"35",X"35",X"35",X"35",X"35",X"35",X"35",X"35",X"35",X"35",X"35",X"35",X"35",X"35",X"35",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"2C",X"2D",X"2E",X"2F",X"2F",X"30",X"31",X"32",X"32",X"2C",X"2D",
		X"31",X"32",X"33",X"30",X"31",X"3A",X"00",X"B8",X"01",X"FD",X"FF",X"ED",X"5B",X"3A",X"80",X"CB",
		X"9B",X"DD",X"2A",X"38",X"80",X"DD",X"7E",X"01",X"E6",X"07",X"67",X"DD",X"6E",X"00",X"29",X"29",
		X"29",X"7C",X"B5",X"C8",X"ED",X"52",X"D8",X"DD",X"09",X"DD",X"22",X"38",X"80",X"3A",X"00",X"B8",
		X"18",X"E3",X"3A",X"00",X"B8",X"01",X"03",X"00",X"ED",X"5B",X"3A",X"80",X"CB",X"9B",X"DD",X"2A",
		X"38",X"80",X"DD",X"7E",X"01",X"E6",X"07",X"67",X"DD",X"6E",X"00",X"29",X"29",X"29",X"B7",X"ED",
		X"52",X"28",X"0D",X"3F",X"D8",X"DD",X"09",X"DD",X"22",X"38",X"80",X"3A",X"00",X"B8",X"18",X"E2",
		X"2A",X"38",X"80",X"09",X"22",X"38",X"80",X"C9",X"ED",X"44",X"4F",X"3A",X"37",X"80",X"81",X"32",
		X"37",X"80",X"06",X"16",X"21",X"04",X"98",X"77",X"23",X"10",X"FC",X"C9",X"2C",X"13",X"E2",X"14",
		X"E9",X"16",X"E1",X"18",X"D0",X"1A",X"07",X"1D",X"FC",X"1E",X"B5",X"20",X"E0",X"22",X"B4",X"24",
		X"2B",X"26",X"5F",X"28",X"87",X"2A",X"2E",X"2C",X"C9",X"2D",X"D3",X"2F",X"00",X"00",X"00",X"20",
		X"00",X"42",X"20",X"00",X"2A",X"20",X"00",X"32",X"22",X"00",X"6C",X"26",X"00",X"26",X"28",X"00",
		X"64",X"36",X"00",X"24",X"3C",X"80",X"0C",X"42",X"80",X"03",X"42",X"00",X"27",X"44",X"00",X"47",
		X"44",X"48",X"10",X"4C",X"00",X"51",X"4E",X"00",X"6F",X"50",X"00",X"31",X"58",X"30",X"03",X"5C",
		X"00",X"48",X"62",X"00",X"22",X"64",X"00",X"41",X"66",X"00",X"41",X"66",X"98",X"0E",X"66",X"80",
		X"12",X"70",X"00",X"23",X"7A",X"48",X"08",X"7A",X"80",X"0B",X"7A",X"00",X"4F",X"7C",X"00",X"4F",
		X"7E",X"00",X"31",X"80",X"00",X"33",X"86",X"00",X"22",X"8A",X"00",X"2D",X"92",X"00",X"51",X"94",
		X"00",X"33",X"98",X"00",X"25",X"98",X"80",X"0A",X"9C",X"48",X"0C",X"A2",X"00",X"45",X"A2",X"00",
		X"2B",X"A8",X"80",X"12",X"AA",X"00",X"21",X"AC",X"00",X"21",X"AC",X"00",X"30",X"AE",X"00",X"4E",
		X"B6",X"30",X"05",X"B8",X"00",X"29",X"BE",X"00",X"23",X"C0",X"00",X"23",X"C2",X"80",X"0E",X"C6",
		X"00",X"6C",X"C8",X"00",X"8A",X"CA",X"00",X"6C",X"CC",X"00",X"2E",X"DA",X"00",X"51",X"DC",X"80",
		X"0A",X"DE",X"00",X"25",X"E0",X"00",X"27",X"E2",X"00",X"29",X"E2",X"60",X"02",X"F2",X"00",X"22",
		X"F2",X"48",X"11",X"F8",X"00",X"2B",X"FA",X"00",X"2D",X"FA",X"00",X"33",X"FC",X"98",X"06",X"FC",
		X"00",X"33",X"06",X"01",X"24",X"0E",X"81",X"11",X"10",X"01",X"24",X"12",X"01",X"44",X"14",X"01",
		X"44",X"1A",X"01",X"27",X"1A",X"01",X"4C",X"1C",X"01",X"2E",X"1E",X"61",X"0C",X"26",X"01",X"27",
		X"2E",X"01",X"22",X"2E",X"01",X"51",X"2E",X"81",X"0A",X"30",X"01",X"33",X"34",X"01",X"25",X"36",
		X"01",X"25",X"38",X"01",X"2D",X"3A",X"01",X"2F",X"48",X"01",X"27",X"48",X"81",X"12",X"4A",X"01",
		X"27",X"4C",X"01",X"29",X"4C",X"01",X"30",X"4E",X"01",X"29",X"4E",X"01",X"30",X"50",X"01",X"27",
		X"50",X"31",X"13",X"56",X"01",X"21",X"5A",X"01",X"2E",X"5C",X"01",X"6C",X"5E",X"01",X"6C",X"60",
		X"99",X"04",X"60",X"01",X"2E",X"68",X"01",X"33",X"6A",X"01",X"45",X"6A",X"01",X"33",X"6C",X"01",
		X"45",X"6E",X"01",X"65",X"70",X"01",X"67",X"72",X"01",X"49",X"74",X"61",X"0F",X"78",X"01",X"21",
		X"7A",X"01",X"41",X"7A",X"01",X"2F",X"7C",X"01",X"4D",X"7E",X"01",X"2D",X"7E",X"81",X"07",X"82",
		X"01",X"23",X"8A",X"01",X"2A",X"8A",X"31",X"0E",X"8A",X"01",X"33",X"92",X"99",X"0B",X"94",X"01",
		X"25",X"9C",X"01",X"21",X"9E",X"49",X"07",X"9E",X"01",X"6F",X"A8",X"01",X"49",X"AC",X"81",X"11",
		X"B0",X"01",X"31",X"B2",X"01",X"23",X"B2",X"01",X"30",X"B4",X"01",X"25",X"B4",X"01",X"2E",X"B6",
		X"01",X"27",X"B6",X"01",X"2C",X"BA",X"81",X"09",X"BC",X"01",X"33",X"C2",X"01",X"21",X"C2",X"01",
		X"26",X"C2",X"01",X"2E",X"C4",X"01",X"28",X"C4",X"01",X"2C",X"C6",X"01",X"2A",X"CC",X"81",X"10",
		X"D0",X"99",X"05",X"D4",X"01",X"2F",X"D6",X"01",X"2F",X"DC",X"81",X"05",X"DE",X"31",X"0A",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"20",X"00",X"42",X"20",X"00",X"4A",X"20",X"00",X"32",X"22",X"00",
		X"6C",X"26",X"00",X"26",X"28",X"00",X"64",X"3C",X"00",X"29",X"3E",X"00",X"4D",X"3E",X"30",X"03",
		X"40",X"00",X"2F",X"44",X"00",X"22",X"44",X"80",X"07",X"46",X"00",X"42",X"48",X"00",X"42",X"4A",
		X"00",X"22",X"52",X"00",X"2E",X"54",X"00",X"2E",X"56",X"00",X"4C",X"56",X"48",X"13",X"58",X"00",
		X"2C",X"5C",X"00",X"41",X"5E",X"00",X"41",X"5E",X"80",X"07",X"66",X"00",X"48",X"68",X"00",X"46",
		X"6A",X"00",X"46",X"70",X"00",X"2F",X"72",X"00",X"4D",X"74",X"98",X"04",X"74",X"00",X"2D",X"80",
		X"80",X"02",X"88",X"00",X"23",X"8A",X"00",X"43",X"8A",X"30",X"0C",X"8C",X"00",X"63",X"8E",X"00",
		X"43",X"90",X"00",X"23",X"96",X"00",X"2A",X"98",X"00",X"68",X"9A",X"00",X"68",X"9C",X"00",X"2A",
		X"9E",X"80",X"13",X"A0",X"98",X"11",X"A8",X"60",X"0D",X"AC",X"00",X"29",X"AE",X"00",X"2F",X"B0",
		X"00",X"23",X"B4",X"80",X"0C",X"B4",X"00",X"51",X"B6",X"00",X"21",X"B6",X"00",X"28",X"BA",X"00",
		X"2D",X"BE",X"00",X"27",X"C0",X"00",X"33",X"C4",X"00",X"23",X"C4",X"00",X"2D",X"CC",X"00",X"24",
		X"CE",X"00",X"44",X"D0",X"00",X"64",X"D0",X"00",X"31",X"D2",X"00",X"64",X"D4",X"00",X"46",X"D4",
		X"00",X"31",X"D6",X"00",X"28",X"DA",X"00",X"21",X"DE",X"00",X"2B",X"E0",X"00",X"4B",X"E2",X"30",
		X"11",X"EA",X"00",X"25",X"EA",X"80",X"10",X"EC",X"00",X"63",X"EE",X"00",X"63",X"F0",X"00",X"63",
		X"F2",X"00",X"26",X"F8",X"00",X"33",X"FA",X"00",X"6F",X"FC",X"80",X"09",X"FC",X"00",X"8D",X"FE",
		X"00",X"8D",X"00",X"01",X"6F",X"02",X"01",X"26",X"0C",X"01",X"26",X"0E",X"01",X"45",X"0E",X"01",
		X"2F",X"10",X"01",X"64",X"10",X"81",X"0B",X"10",X"01",X"4E",X"12",X"61",X"01",X"12",X"01",X"45",
		X"12",X"01",X"2F",X"14",X"01",X"26",X"1A",X"01",X"21",X"1E",X"01",X"2D",X"20",X"01",X"69",X"22",
		X"01",X"49",X"22",X"99",X"02",X"24",X"01",X"2A",X"2A",X"81",X"13",X"2E",X"01",X"2E",X"30",X"01",
		X"4D",X"32",X"01",X"2E",X"36",X"01",X"25",X"38",X"61",X"11",X"3A",X"01",X"63",X"3C",X"01",X"64",
		X"3C",X"81",X"13",X"3E",X"01",X"46",X"42",X"31",X"0D",X"48",X"01",X"29",X"4A",X"01",X"2A",X"4C",
		X"01",X"2B",X"4E",X"01",X"2C",X"4E",X"01",X"33",X"54",X"81",X"03",X"58",X"01",X"64",X"5A",X"01",
		X"65",X"5C",X"01",X"66",X"5C",X"49",X"0F",X"62",X"01",X"21",X"64",X"01",X"22",X"6C",X"01",X"26",
		X"6C",X"01",X"2D",X"6E",X"01",X"25",X"6E",X"01",X"2E",X"70",X"01",X"44",X"70",X"01",X"2F",X"70",
		X"81",X"09",X"72",X"01",X"25",X"7C",X"01",X"29",X"7E",X"01",X"67",X"7E",X"81",X"11",X"80",X"01",
		X"24",X"82",X"01",X"25",X"84",X"01",X"26",X"86",X"01",X"87",X"8C",X"01",X"21",X"90",X"99",X"0F",
		X"94",X"01",X"45",X"9E",X"01",X"41",X"9E",X"61",X"10",X"9E",X"01",X"33",X"A8",X"01",X"2A",X"AA",
		X"01",X"2A",X"AC",X"01",X"2C",X"AE",X"01",X"2E",X"B0",X"01",X"2E",X"B0",X"81",X"12",X"B2",X"61",
		X"09",X"B2",X"01",X"2E",X"B4",X"01",X"2E",X"B6",X"01",X"25",X"B6",X"01",X"2F",X"B8",X"01",X"30",
		X"BA",X"01",X"30",X"BC",X"01",X"21",X"BC",X"61",X"05",X"BC",X"01",X"31",X"BE",X"01",X"31",X"C0",
		X"01",X"31",X"C2",X"61",X"0A",X"C2",X"01",X"31",X"C4",X"01",X"31",X"C6",X"99",X"05",X"C6",X"01",
		X"31",X"CE",X"01",X"21",X"CE",X"01",X"33",X"D0",X"01",X"49",X"D2",X"31",X"05",X"D4",X"01",X"30",
		X"D8",X"01",X"69",X"DA",X"01",X"41",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"20",X"00",X"42",X"20",
		X"00",X"2A",X"20",X"00",X"32",X"22",X"00",X"6C",X"26",X"00",X"26",X"28",X"00",X"64",X"32",X"00",
		X"49",X"34",X"00",X"49",X"3A",X"00",X"31",X"3A",X"60",X"0E",X"3C",X"00",X"50",X"3E",X"00",X"31",
		X"46",X"80",X"0B",X"4E",X"80",X"03",X"4E",X"00",X"2A",X"50",X"00",X"68",X"52",X"00",X"68",X"54",
		X"00",X"2A",X"56",X"30",X"03",X"5C",X"00",X"42",X"5E",X"00",X"62",X"60",X"00",X"42",X"62",X"00",
		X"22",X"64",X"00",X"22",X"64",X"00",X"6D",X"66",X"00",X"6D",X"6E",X"00",X"49",X"70",X"00",X"48",
		X"72",X"00",X"29",X"76",X"30",X"10",X"7A",X"00",X"25",X"7C",X"00",X"24",X"7E",X"00",X"43",X"7E",
		X"80",X"12",X"80",X"00",X"62",X"82",X"00",X"62",X"84",X"00",X"42",X"84",X"80",X"12",X"86",X"00",
		X"22",X"88",X"00",X"29",X"8A",X"00",X"49",X"8C",X"00",X"2B",X"92",X"00",X"50",X"98",X"00",X"49",
		X"9A",X"00",X"2A",X"9C",X"00",X"2A",X"9E",X"00",X"2B",X"A2",X"98",X"02",X"A2",X"80",X"0F",X"AA",
		X"00",X"4B",X"AA",X"48",X"11",X"AC",X"00",X"69",X"AE",X"00",X"4A",X"B2",X"60",X"02",X"B6",X"00",
		X"44",X"B6",X"80",X"08",X"B8",X"00",X"25",X"BE",X"00",X"42",X"C0",X"00",X"62",X"C2",X"00",X"22",
		X"C4",X"00",X"23",X"C4",X"80",X"13",X"C6",X"00",X"23",X"CC",X"00",X"49",X"CE",X"30",X"06",X"D4",
		X"00",X"32",X"D6",X"00",X"50",X"D8",X"00",X"6E",X"D8",X"80",X"04",X"DA",X"00",X"8C",X"DC",X"00",
		X"4F",X"DE",X"00",X"4F",X"E2",X"00",X"22",X"E4",X"00",X"42",X"E6",X"00",X"22",X"EC",X"80",X"10",
		X"F8",X"80",X"12",X"FA",X"00",X"29",X"FC",X"00",X"46",X"FC",X"98",X"0E",X"FE",X"00",X"46",X"00",
		X"61",X"02",X"00",X"01",X"24",X"0A",X"01",X"6B",X"0C",X"49",X"06",X"0C",X"01",X"6B",X"0E",X"01",
		X"6B",X"16",X"81",X"08",X"18",X"01",X"32",X"1A",X"01",X"50",X"1C",X"01",X"46",X"1C",X"01",X"32",
		X"1E",X"01",X"46",X"1E",X"01",X"32",X"20",X"01",X"45",X"20",X"01",X"32",X"22",X"01",X"45",X"22",
		X"01",X"50",X"24",X"01",X"50",X"26",X"01",X"6E",X"28",X"01",X"50",X"28",X"31",X"0B",X"2A",X"01",
		X"32",X"2C",X"01",X"22",X"2E",X"01",X"22",X"2E",X"99",X"0A",X"34",X"81",X"12",X"38",X"01",X"49",
		X"3A",X"01",X"49",X"3C",X"01",X"67",X"40",X"61",X"03",X"40",X"01",X"31",X"46",X"01",X"4B",X"48",
		X"01",X"4B",X"4A",X"01",X"22",X"4C",X"01",X"42",X"4E",X"01",X"42",X"4E",X"81",X"0B",X"50",X"01",
		X"43",X"5C",X"01",X"23",X"5E",X"01",X"42",X"5E",X"01",X"2C",X"60",X"01",X"42",X"60",X"01",X"4B",
		X"62",X"01",X"42",X"62",X"01",X"2C",X"64",X"01",X"42",X"64",X"49",X"08",X"68",X"99",X"0E",X"6C",
		X"81",X"07",X"6E",X"01",X"27",X"70",X"01",X"46",X"72",X"01",X"27",X"72",X"01",X"50",X"74",X"01",
		X"4F",X"74",X"31",X"0B",X"80",X"01",X"82",X"80",X"81",X"0F",X"88",X"81",X"04",X"88",X"01",X"A8",
		X"92",X"01",X"82",X"92",X"81",X"0F",X"9A",X"81",X"04",X"9A",X"01",X"A8",X"A2",X"01",X"28",X"A4",
		X"99",X"04",X"A8",X"01",X"2C",X"A8",X"01",X"31",X"AC",X"01",X"25",X"B0",X"01",X"30",X"B2",X"01",
		X"22",X"B4",X"01",X"29",X"B4",X"01",X"2D",X"BA",X"01",X"2E",X"BC",X"81",X"04",X"BE",X"01",X"2A",
		X"BE",X"01",X"32",X"C0",X"49",X"04",X"C6",X"01",X"44",X"CA",X"01",X"2B",X"CE",X"01",X"22",X"CE",
		X"81",X"0F",X"D2",X"99",X"0B",X"D8",X"01",X"24",X"D8",X"01",X"28",X"D8",X"01",X"4F",X"FF",X"FF",
		X"FF",X"00",X"00",X"00",X"20",X"00",X"42",X"20",X"00",X"2A",X"20",X"00",X"32",X"22",X"00",X"6C",
		X"26",X"00",X"26",X"28",X"00",X"64",X"2E",X"00",X"2E",X"30",X"00",X"2D",X"32",X"00",X"2B",X"3C",
		X"80",X"0B",X"3C",X"00",X"32",X"3E",X"00",X"50",X"40",X"00",X"50",X"42",X"00",X"46",X"42",X"00",
		X"50",X"44",X"00",X"27",X"44",X"00",X"32",X"4A",X"30",X"0E",X"4E",X"80",X"06",X"52",X"00",X"22",
		X"54",X"00",X"42",X"56",X"00",X"42",X"58",X"00",X"22",X"58",X"00",X"2B",X"58",X"80",X"12",X"60",
		X"98",X"0F",X"64",X"00",X"47",X"66",X"00",X"46",X"68",X"48",X"0C",X"6E",X"00",X"4A",X"70",X"00",
		X"4A",X"72",X"00",X"22",X"72",X"00",X"4A",X"74",X"00",X"42",X"76",X"00",X"22",X"76",X"60",X"0F",
		X"7A",X"80",X"08",X"7C",X"00",X"4C",X"7E",X"00",X"6A",X"80",X"00",X"4B",X"84",X"00",X"26",X"86",
		X"00",X"28",X"90",X"00",X"22",X"90",X"80",X"10",X"96",X"00",X"27",X"96",X"00",X"30",X"98",X"00",
		X"27",X"98",X"00",X"31",X"9A",X"00",X"50",X"9C",X"30",X"02",X"9C",X"00",X"4F",X"A0",X"00",X"2B",
		X"A2",X"00",X"24",X"A2",X"00",X"4C",X"A8",X"80",X"07",X"AC",X"00",X"42",X"AC",X"98",X"08",X"AE",
		X"00",X"24",X"AE",X"48",X"11",X"B4",X"00",X"50",X"B6",X"00",X"50",X"B8",X"00",X"6E",X"B8",X"80",
		X"07",X"C0",X"00",X"2B",X"C2",X"00",X"22",X"C4",X"00",X"42",X"C4",X"00",X"32",X"C6",X"00",X"62",
		X"C8",X"00",X"82",X"CE",X"00",X"2E",X"D2",X"48",X"08",X"D4",X"00",X"32",X"DC",X"80",X"0B",X"E0",
		X"00",X"2B",X"E0",X"60",X"10",X"E2",X"00",X"2B",X"E4",X"00",X"2A",X"E4",X"98",X"10",X"E6",X"00",
		X"49",X"E8",X"00",X"48",X"EA",X"00",X"47",X"EC",X"00",X"26",X"FC",X"00",X"22",X"FC",X"00",X"2C",
		X"FC",X"80",X"10",X"FE",X"00",X"2C",X"00",X"01",X"4B",X"02",X"01",X"4B",X"04",X"01",X"4B",X"06",
		X"61",X"06",X"06",X"01",X"6A",X"08",X"01",X"2B",X"0A",X"01",X"2C",X"0C",X"01",X"2D",X"14",X"81",
		X"08",X"18",X"01",X"26",X"1A",X"01",X"64",X"1C",X"01",X"45",X"1C",X"01",X"32",X"1E",X"01",X"32",
		X"30",X"01",X"2F",X"30",X"81",X"13",X"32",X"01",X"2E",X"34",X"01",X"4D",X"36",X"01",X"27",X"36",
		X"01",X"4D",X"3C",X"01",X"22",X"3E",X"49",X"09",X"48",X"99",X"0B",X"4C",X"01",X"22",X"4E",X"01",
		X"42",X"4E",X"81",X"10",X"52",X"01",X"4D",X"54",X"01",X"6D",X"56",X"81",X"07",X"56",X"01",X"8C",
		X"58",X"01",X"8C",X"5A",X"01",X"23",X"5A",X"01",X"6E",X"5C",X"01",X"42",X"5E",X"01",X"22",X"64",
		X"01",X"28",X"64",X"01",X"32",X"66",X"01",X"29",X"66",X"01",X"32",X"66",X"81",X"0E",X"68",X"01",
		X"32",X"6A",X"01",X"32",X"6C",X"01",X"42",X"6C",X"01",X"50",X"6E",X"01",X"42",X"6E",X"01",X"6E",
		X"70",X"31",X"0B",X"70",X"01",X"6E",X"72",X"01",X"6E",X"74",X"81",X"06",X"74",X"01",X"50",X"80",
		X"01",X"24",X"80",X"49",X"09",X"84",X"01",X"2D",X"88",X"31",X"11",X"8A",X"01",X"27",X"92",X"49",
		X"07",X"94",X"01",X"2E",X"9A",X"61",X"02",X"9E",X"01",X"25",X"A0",X"49",X"0D",X"A8",X"01",X"2A",
		X"A8",X"61",X"10",X"AC",X"01",X"22",X"B0",X"01",X"2E",X"B2",X"31",X"03",X"B6",X"81",X"0A",X"BC",
		X"01",X"25",X"BC",X"49",X"09",X"C0",X"01",X"32",X"C6",X"01",X"22",X"C6",X"01",X"2C",X"C8",X"31",
		X"0F",X"D0",X"81",X"07",X"D4",X"01",X"25",X"D6",X"61",X"09",X"D8",X"01",X"2D",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"20",X"00",X"24",X"20",X"00",X"2A",X"20",X"00",X"31",X"22",X"00",X"6C",X"26",
		X"00",X"26",X"28",X"00",X"64",X"34",X"00",X"2C",X"36",X"00",X"4A",X"38",X"00",X"68",X"3A",X"00",
		X"86",X"3C",X"00",X"86",X"3E",X"00",X"68",X"40",X"00",X"4A",X"40",X"30",X"11",X"42",X"80",X"03",
		X"42",X"00",X"2C",X"46",X"00",X"23",X"48",X"00",X"23",X"48",X"98",X"0E",X"54",X"00",X"2D",X"56",
		X"00",X"69",X"58",X"00",X"69",X"5A",X"00",X"4B",X"5C",X"00",X"23",X"5E",X"00",X"23",X"60",X"00",
		X"23",X"64",X"60",X"0E",X"66",X"00",X"48",X"68",X"00",X"66",X"6A",X"00",X"46",X"6C",X"00",X"46",
		X"6C",X"18",X"14",X"6E",X"80",X"10",X"74",X"00",X"31",X"76",X"00",X"4F",X"78",X"00",X"6D",X"7A",
		X"00",X"6D",X"7C",X"00",X"6D",X"80",X"00",X"4F",X"82",X"98",X"03",X"82",X"00",X"31",X"86",X"00",
		X"2C",X"88",X"00",X"2B",X"8A",X"00",X"2A",X"8C",X"80",X"11",X"90",X"80",X"11",X"92",X"00",X"6A",
		X"94",X"00",X"68",X"98",X"30",X"04",X"9C",X"00",X"27",X"9E",X"00",X"28",X"A0",X"00",X"29",X"A2",
		X"00",X"2A",X"A6",X"00",X"23",X"A8",X"00",X"23",X"A8",X"80",X"05",X"AA",X"00",X"23",X"AB",X"30",
		X"11",X"AE",X"00",X"28",X"B0",X"00",X"27",X"B2",X"00",X"26",X"B2",X"98",X"0D",X"B8",X"80",X"11",
		X"C0",X"00",X"23",X"C2",X"00",X"23",X"C4",X"00",X"23",X"C4",X"00",X"29",X"C6",X"00",X"23",X"C6",
		X"00",X"2A",X"C8",X"00",X"49",X"CA",X"00",X"4A",X"CE",X"80",X"10",X"DA",X"00",X"31",X"DA",X"48",
		X"09",X"DC",X"00",X"4F",X"DE",X"00",X"4F",X"E0",X"00",X"4F",X"E2",X"00",X"4F",X"E4",X"00",X"4F",
		X"E6",X"00",X"29",X"E6",X"00",X"4F",X"E8",X"00",X"47",X"E8",X"00",X"4F",X"E9",X"60",X"03",X"EA",
		X"00",X"47",X"EC",X"00",X"47",X"EE",X"00",X"67",X"F0",X"00",X"67",X"F2",X"00",X"49",X"F6",X"80",
		X"11",X"FC",X"00",X"23",X"FC",X"00",X"30",X"FE",X"00",X"23",X"FE",X"00",X"30",X"00",X"01",X"23",
		X"00",X"01",X"31",X"00",X"61",X"0C",X"02",X"01",X"23",X"02",X"01",X"29",X"04",X"01",X"23",X"04",
		X"01",X"29",X"06",X"01",X"23",X"06",X"99",X"0E",X"0A",X"31",X"0F",X"10",X"01",X"2B",X"12",X"81",
		X"04",X"12",X"01",X"2B",X"14",X"01",X"2B",X"16",X"01",X"2B",X"18",X"01",X"4B",X"1A",X"01",X"4B",
		X"1C",X"01",X"4C",X"20",X"49",X"0A",X"22",X"01",X"26",X"24",X"01",X"26",X"26",X"01",X"27",X"28",
		X"01",X"28",X"2A",X"01",X"29",X"2A",X"01",X"2F",X"2A",X"01",X"31",X"2E",X"01",X"23",X"3E",X"81",
		X"04",X"40",X"01",X"2A",X"42",X"01",X"49",X"44",X"01",X"68",X"46",X"01",X"87",X"48",X"01",X"87",
		X"4A",X"01",X"87",X"4C",X"01",X"87",X"4E",X"01",X"87",X"50",X"01",X"87",X"52",X"01",X"68",X"54",
		X"01",X"49",X"56",X"01",X"2A",X"58",X"01",X"31",X"58",X"19",X"00",X"5E",X"81",X"04",X"5E",X"01",
		X"48",X"60",X"01",X"49",X"62",X"01",X"48",X"62",X"31",X"10",X"64",X"01",X"47",X"66",X"01",X"46",
		X"68",X"01",X"27",X"6A",X"01",X"27",X"6A",X"01",X"31",X"6C",X"01",X"27",X"6C",X"01",X"4F",X"6E",
		X"01",X"4E",X"70",X"81",X"0A",X"74",X"01",X"23",X"74",X"01",X"29",X"7A",X"99",X"05",X"7A",X"01",
		X"2E",X"80",X"99",X"05",X"80",X"61",X"0F",X"88",X"01",X"25",X"8A",X"61",X"0A",X"8A",X"01",X"2E",
		X"90",X"01",X"31",X"94",X"01",X"43",X"94",X"31",X"0F",X"9C",X"01",X"2D",X"9E",X"61",X"07",X"A2",
		X"01",X"2A",X"A2",X"81",X"0F",X"A8",X"01",X"24",X"A8",X"99",X"09",X"A8",X"01",X"30",X"B2",X"81",
		X"05",X"B2",X"01",X"2A",X"B2",X"61",X"0F",X"B6",X"01",X"27",X"BA",X"01",X"24",X"BC",X"49",X"0A",
		X"BC",X"01",X"2F",X"C4",X"01",X"2A",X"C6",X"61",X"08",X"CA",X"01",X"24",X"CA",X"81",X"0C",X"CA",
		X"01",X"31",X"CE",X"99",X"0C",X"D0",X"61",X"05",X"D8",X"01",X"25",X"D8",X"01",X"29",X"D8",X"01",
		X"2E",X"DA",X"01",X"2F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"20",X"00",X"24",X"20",X"00",X"8A",
		X"22",X"00",X"6C",X"26",X"00",X"25",X"28",X"00",X"63",X"2A",X"00",X"43",X"2C",X"00",X"23",X"2E",
		X"00",X"31",X"34",X"00",X"25",X"3C",X"00",X"2D",X"3E",X"00",X"2B",X"3E",X"80",X"06",X"42",X"00",
		X"2B",X"44",X"60",X"06",X"44",X"00",X"2D",X"46",X"00",X"4F",X"4C",X"00",X"23",X"4C",X"80",X"08",
		X"4E",X"48",X"0F",X"50",X"00",X"2A",X"54",X"00",X"2A",X"54",X"80",X"0F",X"58",X"00",X"29",X"5C",
		X"80",X"03",X"5C",X"00",X"28",X"60",X"00",X"27",X"60",X"18",X"14",X"62",X"00",X"25",X"64",X"00",
		X"23",X"64",X"80",X"0A",X"6A",X"30",X"11",X"6C",X"00",X"2D",X"70",X"00",X"2A",X"74",X"00",X"27",
		X"76",X"60",X"0F",X"78",X"00",X"26",X"7C",X"00",X"26",X"7E",X"80",X"0D",X"82",X"00",X"6D",X"84",
		X"00",X"6D",X"86",X"60",X"08",X"8C",X"80",X"06",X"8E",X"00",X"2C",X"90",X"30",X"05",X"90",X"00",
		X"2E",X"92",X"00",X"30",X"98",X"98",X"05",X"9A",X"80",X"0F",X"9E",X"80",X"05",X"A2",X"00",X"4A",
		X"A4",X"00",X"4C",X"A6",X"00",X"4E",X"A8",X"00",X"4F",X"AC",X"18",X"00",X"AE",X"00",X"2A",X"B0",
		X"00",X"28",X"B4",X"48",X"05",X"B4",X"00",X"28",X"B6",X"00",X"2A",X"B6",X"80",X"0F",X"B8",X"00",
		X"2C",X"BA",X"00",X"2E",X"BC",X"00",X"30",X"BE",X"00",X"23",X"C0",X"00",X"43",X"C2",X"00",X"63",
		X"C4",X"00",X"83",X"C6",X"00",X"A3",X"C8",X"00",X"A3",X"C8",X"80",X"11",X"CA",X"00",X"83",X"D0",
		X"80",X"0A",X"D0",X"60",X"0F",X"D4",X"00",X"2B",X"D6",X"00",X"2E",X"DA",X"00",X"31",X"DC",X"30",
		X"03",X"DC",X"80",X"0A",X"E2",X"00",X"2A",X"E4",X"00",X"2C",X"EA",X"00",X"30",X"EE",X"00",X"29",
		X"F0",X"80",X"06",X"F2",X"00",X"26",X"F6",X"00",X"2F",X"F8",X"00",X"23",X"F8",X"80",X"0D",X"FA",
		X"00",X"2A",X"FC",X"00",X"2F",X"FE",X"00",X"28",X"00",X"01",X"2A",X"02",X"01",X"2D",X"04",X"01",
		X"23",X"06",X"01",X"43",X"06",X"01",X"30",X"08",X"01",X"63",X"0A",X"01",X"43",X"0C",X"01",X"23",
		X"0E",X"81",X"0D",X"12",X"61",X"07",X"14",X"01",X"6D",X"1C",X"01",X"29",X"1E",X"01",X"2B",X"20",
		X"01",X"83",X"22",X"81",X"0F",X"26",X"49",X"05",X"28",X"01",X"2A",X"2A",X"01",X"28",X"32",X"01",
		X"2B",X"34",X"31",X"05",X"34",X"01",X"2D",X"36",X"01",X"30",X"3C",X"81",X"05",X"40",X"01",X"23",
		X"42",X"01",X"43",X"44",X"01",X"63",X"46",X"01",X"43",X"4A",X"81",X"03",X"4C",X"01",X"49",X"4C",
		X"81",X"11",X"4E",X"01",X"29",X"50",X"01",X"47",X"52",X"01",X"63",X"54",X"01",X"43",X"54",X"19",
		X"14",X"56",X"99",X"0B",X"5C",X"01",X"31",X"5E",X"81",X"07",X"5E",X"01",X"4F",X"60",X"01",X"8B",
		X"62",X"01",X"A9",X"64",X"01",X"31",X"6C",X"49",X"0F",X"6E",X"81",X"03",X"70",X"01",X"2A",X"72",
		X"01",X"28",X"72",X"81",X"10",X"74",X"01",X"26",X"76",X"01",X"25",X"78",X"01",X"23",X"7C",X"01",
		X"A9",X"7E",X"01",X"8B",X"84",X"01",X"2D",X"8C",X"01",X"29",X"8C",X"81",X"0F",X"94",X"01",X"25",
		X"98",X"01",X"2A",X"98",X"81",X"0F",X"9E",X"01",X"23",X"A2",X"01",X"2F",X"A4",X"31",X"05",X"A6",
		X"01",X"2A",X"AC",X"01",X"2D",X"B0",X"81",X"08",X"B2",X"01",X"23",X"B8",X"81",X"07",X"B8",X"01",
		X"2F",X"BE",X"01",X"29",X"C2",X"01",X"27",X"C6",X"01",X"27",X"CA",X"01",X"25",X"D4",X"01",X"2A",
		X"D8",X"81",X"0F",X"DA",X"01",X"2A",X"DC",X"49",X"09",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"20",
		X"00",X"24",X"20",X"00",X"4A",X"22",X"00",X"6C",X"26",X"00",X"26",X"28",X"00",X"64",X"2A",X"00",
		X"44",X"30",X"00",X"4D",X"32",X"00",X"2C",X"3E",X"80",X"07",X"42",X"00",X"2A",X"42",X"60",X"0F",
		X"44",X"00",X"28",X"48",X"00",X"27",X"4A",X"00",X"24",X"4A",X"48",X"10",X"4E",X"00",X"2A",X"50",
		X"80",X"0E",X"52",X"00",X"2A",X"56",X"00",X"2A",X"58",X"00",X"4C",X"5A",X"00",X"30",X"5E",X"00",
		X"28",X"60",X"00",X"2A",X"62",X"00",X"2C",X"64",X"00",X"2C",X"66",X"80",X"07",X"66",X"00",X"2C",
		X"68",X"00",X"2C",X"6A",X"00",X"2A",X"6C",X"00",X"28",X"6C",X"80",X"0F",X"6E",X"00",X"25",X"74",
		X"30",X"05",X"74",X"00",X"2A",X"78",X"00",X"2C",X"7C",X"00",X"2E",X"7E",X"00",X"30",X"80",X"00",
		X"26",X"82",X"80",X"09",X"86",X"00",X"2B",X"8A",X"00",X"2D",X"8C",X"00",X"30",X"90",X"00",X"29",
		X"96",X"80",X"05",X"98",X"60",X"0A",X"9A",X"00",X"30",X"9E",X"00",X"2B",X"A2",X"80",X"0D",X"A6",
		X"00",X"27",X"AA",X"00",X"24",X"AE",X"80",X"07",X"B0",X"00",X"2C",X"B2",X"48",X"08",X"B4",X"00",
		X"2E",X"BA",X"00",X"28",X"BC",X"00",X"25",X"C0",X"80",X"0E",X"C2",X"00",X"2A",X"C6",X"00",X"2C",
		X"CA",X"00",X"2E",X"CE",X"80",X"05",X"CE",X"00",X"30",X"D4",X"98",X"07",X"DA",X"60",X"10",X"DC",
		X"00",X"24",X"DE",X"00",X"84",X"E4",X"00",X"29",X"EA",X"80",X"0F",X"EC",X"00",X"2A",X"F0",X"00",
		X"2C",X"F4",X"00",X"4D",X"F6",X"80",X"07",X"FA",X"00",X"28",X"FE",X"00",X"44",X"FE",X"60",X"0D",
		X"04",X"01",X"2A",X"04",X"81",X"0F",X"06",X"01",X"2C",X"0A",X"01",X"2F",X"0C",X"81",X"07",X"10",
		X"01",X"24",X"10",X"01",X"28",X"12",X"01",X"44",X"14",X"31",X"0F",X"18",X"01",X"2A",X"1A",X"01",
		X"6C",X"20",X"01",X"44",X"22",X"81",X"0F",X"24",X"61",X"08",X"26",X"01",X"4B",X"2A",X"81",X"08",
		X"2A",X"01",X"30",X"2E",X"01",X"28",X"30",X"49",X"0D",X"32",X"01",X"26",X"34",X"01",X"24",X"36",
		X"01",X"2D",X"38",X"01",X"2F",X"3C",X"61",X"0D",X"3E",X"81",X"05",X"3E",X"01",X"2A",X"42",X"01",
		X"2A",X"46",X"81",X"06",X"46",X"01",X"2A",X"4A",X"01",X"2A",X"4E",X"01",X"2A",X"4E",X"81",X"0F",
		X"52",X"01",X"28",X"52",X"31",X"10",X"54",X"01",X"24",X"54",X"31",X"06",X"58",X"81",X"0F",X"5A",
		X"01",X"2B",X"5E",X"01",X"2C",X"60",X"81",X"09",X"62",X"01",X"4E",X"66",X"61",X"05",X"68",X"01",
		X"2A",X"6C",X"01",X"2A",X"6E",X"01",X"26",X"74",X"99",X"0C",X"7C",X"01",X"64",X"7E",X"01",X"84",
		X"86",X"01",X"29",X"8C",X"01",X"28",X"8E",X"81",X"0C",X"90",X"01",X"26",X"94",X"01",X"24",X"98",
		X"01",X"2C",X"9C",X"81",X"0F",X"9E",X"81",X"06",X"A4",X"01",X"24",X"A4",X"49",X"0F",X"AE",X"81",
		X"05",X"B2",X"01",X"4D",X"B8",X"61",X"06",X"BA",X"81",X"0D",X"C2",X"99",X"07",X"CA",X"01",X"2A",
		X"CC",X"01",X"28",X"CE",X"01",X"26",X"D0",X"01",X"24",X"D8",X"01",X"2A",X"DC",X"01",X"2C",X"DE",
		X"01",X"4E",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"20",X"00",X"24",X"20",X"00",X"8A",X"22",X"00",
		X"6C",X"26",X"00",X"26",X"28",X"00",X"64",X"2A",X"00",X"44",X"2C",X"00",X"24",X"30",X"00",X"30",
		X"32",X"00",X"30",X"34",X"00",X"2E",X"3C",X"00",X"26",X"3E",X"00",X"44",X"40",X"00",X"44",X"40",
		X"80",X"0E",X"42",X"00",X"26",X"46",X"00",X"2E",X"48",X"00",X"6C",X"4A",X"00",X"6C",X"4C",X"80",
		X"08",X"4C",X"00",X"4E",X"50",X"00",X"26",X"52",X"00",X"44",X"52",X"18",X"14",X"54",X"00",X"44",
		X"56",X"00",X"64",X"58",X"00",X"84",X"5A",X"00",X"84",X"5A",X"48",X"0E",X"5C",X"00",X"64",X"5E",
		X"00",X"44",X"60",X"00",X"30",X"62",X"00",X"4E",X"64",X"80",X"06",X"64",X"00",X"6C",X"66",X"00",
		X"8A",X"68",X"00",X"4E",X"6C",X"00",X"24",X"6E",X"00",X"44",X"70",X"00",X"44",X"72",X"00",X"64",
		X"72",X"80",X"0E",X"74",X"00",X"64",X"76",X"00",X"44",X"7C",X"00",X"44",X"7E",X"00",X"44",X"80",
		X"00",X"64",X"80",X"48",X"0E",X"82",X"00",X"44",X"86",X"80",X"0E",X"88",X"00",X"2A",X"88",X"18",
		X"14",X"8A",X"00",X"2A",X"8C",X"00",X"4A",X"8E",X"00",X"4A",X"90",X"00",X"6A",X"92",X"00",X"4A",
		X"94",X"00",X"4A",X"96",X"00",X"6A",X"98",X"00",X"4E",X"9A",X"80",X"06",X"9A",X"00",X"30",X"9E",
		X"00",X"24",X"A0",X"00",X"44",X"A2",X"00",X"44",X"A4",X"00",X"64",X"A6",X"00",X"64",X"A6",X"48",
		X"0E",X"A8",X"00",X"84",X"AA",X"00",X"64",X"AC",X"00",X"44",X"AE",X"00",X"24",X"B2",X"00",X"6C",
		X"B4",X"00",X"8A",X"B6",X"00",X"6C",X"BA",X"80",X"0C",X"BC",X"00",X"2C",X"BE",X"00",X"6A",X"C0",
		X"00",X"6A",X"C0",X"18",X"14",X"C2",X"00",X"4C",X"C6",X"80",X"04",X"CC",X"00",X"26",X"CE",X"00",
		X"44",X"D0",X"00",X"64",X"D2",X"00",X"66",X"D2",X"30",X"10",X"D4",X"00",X"2A",X"DA",X"00",X"46",
		X"DC",X"00",X"48",X"DE",X"18",X"14",X"E0",X"60",X"08",X"E4",X"80",X"0A",X"E6",X"00",X"26",X"E8",
		X"00",X"46",X"EA",X"00",X"66",X"EC",X"00",X"84",X"EE",X"00",X"64",X"EE",X"80",X"10",X"F4",X"00",
		X"4E",X"F6",X"00",X"6C",X"F8",X"00",X"6C",X"FA",X"00",X"6A",X"FE",X"80",X"06",X"04",X"01",X"4C",
		X"06",X"01",X"6C",X"08",X"49",X"06",X"08",X"01",X"4C",X"0E",X"19",X"00",X"12",X"01",X"44",X"14",
		X"01",X"A4",X"16",X"01",X"A4",X"18",X"01",X"A4",X"1A",X"01",X"84",X"1C",X"01",X"64",X"1E",X"01",
		X"64",X"20",X"01",X"44",X"20",X"81",X"0E",X"22",X"01",X"24",X"26",X"01",X"30",X"28",X"01",X"4E",
		X"2A",X"81",X"06",X"2A",X"01",X"6C",X"2C",X"01",X"8A",X"2E",X"01",X"8A",X"30",X"01",X"8A",X"32",
		X"01",X"6C",X"36",X"19",X"00",X"3A",X"81",X"08",X"3C",X"01",X"24",X"3E",X"01",X"24",X"40",X"01",
		X"44",X"42",X"01",X"64",X"44",X"01",X"64",X"46",X"01",X"64",X"46",X"49",X"0C",X"46",X"81",X"10",
		X"48",X"01",X"44",X"4E",X"31",X"06",X"50",X"01",X"4C",X"52",X"01",X"6A",X"54",X"01",X"6A",X"56",
		X"01",X"6C",X"5A",X"81",X"08",X"5E",X"01",X"24",X"60",X"01",X"24",X"60",X"61",X"0C",X"62",X"01",
		X"44",X"62",X"19",X"14",X"64",X"01",X"44",X"66",X"01",X"64",X"66",X"81",X"10",X"6C",X"99",X"0A",
		X"72",X"01",X"44",X"74",X"01",X"64",X"76",X"01",X"64",X"78",X"01",X"44",X"7A",X"19",X"00",X"7A",
		X"81",X"0E",X"7E",X"49",X"08",X"82",X"81",X"0F",X"84",X"01",X"2A",X"88",X"01",X"2C",X"8C",X"81",
		X"06",X"90",X"01",X"30",X"92",X"01",X"47",X"9A",X"81",X"08",X"9E",X"01",X"2A",X"A0",X"49",X"05",
		X"A2",X"01",X"4D",X"A6",X"81",X"08",X"A8",X"01",X"24",X"AC",X"61",X"0D",X"AE",X"99",X"06",X"B2",
		X"01",X"4D",X"BA",X"01",X"49",X"BC",X"01",X"44",X"BE",X"81",X"0F",X"C6",X"01",X"2A",X"C8",X"01",
		X"2E",X"CA",X"81",X"06",X"D0",X"01",X"64",X"DA",X"01",X"2C",X"DC",X"01",X"30",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"20",X"00",X"6A",X"22",X"00",X"4C",X"26",X"00",X"25",X"28",X"00",X"45",X"2A",
		X"00",X"25",X"2C",X"00",X"25",X"2E",X"00",X"2F",X"30",X"00",X"4D",X"32",X"00",X"6B",X"34",X"00",
		X"4D",X"36",X"00",X"2F",X"3A",X"00",X"25",X"3C",X"00",X"2B",X"3E",X"80",X"07",X"42",X"00",X"29",
		X"44",X"00",X"2A",X"48",X"48",X"07",X"48",X"00",X"2F",X"4E",X"00",X"27",X"50",X"00",X"25",X"50",
		X"80",X"0B",X"54",X"00",X"2B",X"56",X"00",X"2D",X"58",X"00",X"2F",X"5E",X"00",X"2A",X"5E",X"80",
		X"05",X"64",X"80",X"05",X"66",X"00",X"29",X"6A",X"00",X"27",X"6C",X"60",X"0A",X"6C",X"00",X"2F",
		X"70",X"80",X"0D",X"72",X"00",X"28",X"74",X"00",X"2A",X"78",X"00",X"2C",X"7C",X"80",X"08",X"80",
		X"00",X"2A",X"82",X"80",X"0F",X"84",X"00",X"28",X"86",X"00",X"2F",X"88",X"00",X"29",X"8C",X"00",
		X"2D",X"8E",X"00",X"25",X"90",X"18",X"00",X"94",X"00",X"29",X"94",X"80",X"0D",X"98",X"00",X"28",
		X"98",X"18",X"14",X"9A",X"00",X"25",X"9C",X"48",X"0D",X"A2",X"80",X"08",X"A4",X"00",X"2D",X"A6",
		X"00",X"25",X"A6",X"00",X"2F",X"A8",X"00",X"45",X"AC",X"60",X"0A",X"B4",X"80",X"08",X"B4",X"00",
		X"2B",X"B6",X"00",X"2D",X"B8",X"00",X"2F",X"BA",X"98",X"07",X"C2",X"00",X"2B",X"C4",X"00",X"65",
		X"C6",X"00",X"45",X"C8",X"00",X"25",X"CC",X"80",X"08",X"CE",X"00",X"4D",X"D0",X"00",X"2F",X"D2",
		X"00",X"28",X"DA",X"00",X"47",X"DA",X"48",X"0D",X"DC",X"00",X"45",X"E2",X"00",X"28",X"E4",X"00",
		X"29",X"E6",X"30",X"06",X"E8",X"00",X"4D",X"EC",X"00",X"28",X"F0",X"80",X"0D",X"F2",X"00",X"25",
		X"F4",X"00",X"45",X"F4",X"98",X"0B",X"F6",X"00",X"45",X"F8",X"00",X"25",X"FA",X"60",X"0F",X"FE",
		X"00",X"29",X"02",X"01",X"2B",X"04",X"81",X"0F",X"06",X"01",X"25",X"06",X"01",X"2C",X"0A",X"81",
		X"08",X"0A",X"01",X"2C",X"0E",X"61",X"06",X"10",X"01",X"2F",X"12",X"81",X"0B",X"16",X"01",X"28",
		X"18",X"01",X"2A",X"1C",X"01",X"2F",X"1E",X"81",X"06",X"22",X"01",X"2A",X"26",X"01",X"25",X"26",
		X"81",X"0E",X"2A",X"01",X"2D",X"2C",X"31",X"08",X"30",X"01",X"2B",X"32",X"01",X"29",X"36",X"01",
		X"2F",X"38",X"61",X"09",X"3E",X"01",X"27",X"40",X"01",X"25",X"40",X"81",X"0D",X"44",X"01",X"2C",
		X"48",X"81",X"08",X"4C",X"01",X"27",X"4E",X"01",X"2F",X"50",X"01",X"25",X"56",X"01",X"2A",X"58",
		X"01",X"68",X"5A",X"01",X"2A",X"5C",X"01",X"68",X"5E",X"01",X"2A",X"60",X"31",X"0D",X"66",X"81",
		X"0A",X"66",X"01",X"2D",X"68",X"01",X"2F",X"6C",X"01",X"27",X"6E",X"01",X"25",X"74",X"81",X"07",
		X"74",X"01",X"2F",X"78",X"01",X"29",X"7C",X"99",X"0A",X"82",X"01",X"2A",X"88",X"81",X"08",X"8C",
		X"01",X"2D",X"90",X"81",X"05",X"94",X"01",X"28",X"94",X"81",X"0D",X"9A",X"81",X"0D",X"9C",X"01",
		X"25",X"A0",X"01",X"2D",X"A2",X"81",X"06",X"A6",X"01",X"2A",X"AC",X"01",X"2F",X"AE",X"81",X"07",
		X"B6",X"81",X"08",X"B8",X"81",X"0E",X"BC",X"81",X"06",X"C0",X"01",X"2B",X"C6",X"01",X"2F",X"C8",
		X"01",X"2F",X"CC",X"01",X"25",X"CC",X"81",X"0B",X"D2",X"01",X"2D",X"D6",X"81",X"08",X"DA",X"01",
		X"27",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"20",X"00",X"2A",X"22",X"00",X"4C",X"26",X"00",X"25",
		X"28",X"00",X"45",X"30",X"00",X"2A",X"34",X"00",X"25",X"36",X"00",X"2D",X"38",X"00",X"26",X"3A",
		X"00",X"2B",X"3E",X"00",X"2F",X"46",X"00",X"2A",X"4C",X"00",X"2E",X"4E",X"60",X"08",X"50",X"00",
		X"25",X"52",X"00",X"2F",X"56",X"00",X"28",X"5C",X"00",X"2C",X"60",X"80",X"08",X"62",X"00",X"25",
		X"62",X"00",X"2A",X"66",X"00",X"2F",X"6A",X"00",X"29",X"6C",X"00",X"2D",X"70",X"00",X"25",X"74",
		X"60",X"0D",X"76",X"00",X"2B",X"78",X"00",X"25",X"7E",X"00",X"28",X"7E",X"00",X"4D",X"84",X"00",
		X"25",X"84",X"00",X"2C",X"8E",X"60",X"0D",X"90",X"00",X"2A",X"9A",X"98",X"05",X"A0",X"00",X"2D",
		X"A6",X"80",X"0A",X"AC",X"00",X"2D",X"AE",X"00",X"27",X"B4",X"80",X"0D",X"BA",X"00",X"2E",X"BE",
		X"80",X"06",X"C2",X"00",X"2A",X"C8",X"80",X"0D",X"CC",X"00",X"28",X"D0",X"00",X"25",X"D2",X"80",
		X"07",X"D4",X"00",X"2F",X"D8",X"80",X"0C",X"DC",X"00",X"2B",X"DE",X"80",X"06",X"E4",X"00",X"27",
		X"E8",X"80",X"0B",X"EA",X"00",X"4D",X"F0",X"98",X"09",X"F6",X"00",X"27",X"F8",X"00",X"25",X"FA",
		X"80",X"0A",X"FA",X"00",X"2F",X"FE",X"00",X"2A",X"00",X"01",X"2A",X"02",X"01",X"2A",X"04",X"01",
		X"2A",X"06",X"81",X"06",X"06",X"01",X"2A",X"08",X"01",X"2A",X"0A",X"01",X"2A",X"0C",X"01",X"2A",
		X"0C",X"81",X"0E",X"0E",X"01",X"2A",X"10",X"01",X"2A",X"12",X"01",X"68",X"14",X"01",X"2A",X"18",
		X"49",X"0A",X"24",X"01",X"2B",X"26",X"01",X"2B",X"2A",X"01",X"2B",X"2C",X"01",X"2A",X"2E",X"01",
		X"29",X"30",X"01",X"29",X"30",X"31",X"0E",X"32",X"01",X"27",X"34",X"01",X"25",X"34",X"01",X"2E",
		X"3A",X"01",X"2A",X"3C",X"01",X"2A",X"3E",X"01",X"2A",X"40",X"01",X"2B",X"42",X"01",X"2C",X"44",
		X"99",X"06",X"4E",X"01",X"2F",X"54",X"01",X"28",X"54",X"49",X"0D",X"56",X"01",X"26",X"60",X"31",
		X"09",X"60",X"01",X"2C",X"68",X"01",X"2F",X"6A",X"61",X"05",X"6E",X"31",X"0E",X"70",X"01",X"27",
		X"7A",X"01",X"28",X"7A",X"31",X"0F",X"7C",X"01",X"2A",X"80",X"01",X"2A",X"84",X"61",X"0D",X"8A",
		X"81",X"07",X"8C",X"01",X"2D",X"92",X"81",X"0E",X"96",X"01",X"28",X"9C",X"31",X"08",X"A4",X"49",
		X"0D",X"AA",X"81",X"06",X"AC",X"01",X"2A",X"B0",X"01",X"2C",X"B6",X"01",X"2E",X"BC",X"81",X"0D",
		X"BE",X"61",X"07",X"C6",X"01",X"25",X"C8",X"99",X"0A",X"D0",X"01",X"2A",X"D2",X"01",X"2A",X"D4",
		X"81",X"08",X"DA",X"01",X"25",X"DC",X"01",X"45",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"20",X"00",
		X"6A",X"22",X"00",X"2C",X"26",X"00",X"25",X"28",X"00",X"45",X"2A",X"00",X"45",X"2C",X"00",X"25",
		X"30",X"00",X"2F",X"32",X"00",X"2F",X"34",X"00",X"4D",X"3C",X"00",X"45",X"3E",X"00",X"45",X"3E",
		X"80",X"0C",X"40",X"00",X"45",X"42",X"00",X"65",X"44",X"48",X"0E",X"44",X"00",X"45",X"4A",X"80",
		X"08",X"4C",X"00",X"2F",X"4E",X"00",X"4D",X"50",X"00",X"4D",X"52",X"00",X"6B",X"5A",X"00",X"25",
		X"5C",X"00",X"45",X"5C",X"80",X"0E",X"5E",X"00",X"65",X"60",X"00",X"65",X"62",X"00",X"65",X"62",
		X"18",X"14",X"64",X"00",X"45",X"64",X"48",X"0C",X"66",X"00",X"25",X"6A",X"00",X"2F",X"6C",X"00",
		X"4D",X"6E",X"00",X"6B",X"70",X"00",X"6B",X"74",X"60",X"0C",X"78",X"00",X"29",X"7A",X"00",X"29",
		X"7C",X"00",X"47",X"7C",X"80",X"0E",X"7E",X"00",X"45",X"80",X"00",X"45",X"82",X"00",X"25",X"86",
		X"00",X"25",X"88",X"48",X"06",X"88",X"00",X"4D",X"8A",X"00",X"4D",X"8C",X"18",X"00",X"8C",X"00",
		X"6B",X"8E",X"00",X"6B",X"90",X"00",X"4D",X"92",X"80",X"08",X"92",X"00",X"2F",X"94",X"00",X"2F",
		X"98",X"00",X"29",X"9A",X"00",X"49",X"9A",X"80",X"0E",X"9C",X"00",X"49",X"9E",X"00",X"49",X"A0",
		X"00",X"69",X"A2",X"00",X"4B",X"A4",X"00",X"4B",X"A6",X"00",X"4D",X"A8",X"80",X"06",X"AC",X"00",
		X"25",X"AE",X"00",X"25",X"B0",X"00",X"45",X"B2",X"00",X"45",X"B2",X"30",X"0C",X"B4",X"00",X"25",
		X"B4",X"18",X"14",X"B8",X"00",X"2F",X"BA",X"00",X"4D",X"BC",X"00",X"4D",X"BE",X"00",X"4D",X"C0",
		X"80",X"08",X"C4",X"00",X"25",X"C6",X"00",X"25",X"C8",X"00",X"45",X"CA",X"00",X"45",X"CC",X"00",
		X"45",X"CE",X"00",X"25",X"D2",X"80",X"08",X"D2",X"00",X"2F",X"D6",X"00",X"6B",X"D8",X"00",X"4D",
		X"DA",X"30",X"08",X"E0",X"00",X"29",X"E2",X"00",X"49",X"E2",X"80",X"0E",X"E4",X"00",X"49",X"E6",
		X"00",X"49",X"E8",X"00",X"49",X"EA",X"00",X"4B",X"EC",X"00",X"4B",X"EE",X"00",X"4D",X"F0",X"80",
		X"06",X"F0",X"00",X"2F",X"F4",X"60",X"08",X"F8",X"00",X"25",X"FA",X"00",X"45",X"FC",X"00",X"45",
		X"FE",X"00",X"45",X"00",X"01",X"45",X"02",X"01",X"25",X"04",X"81",X"0E",X"08",X"49",X"0E",X"0A",
		X"01",X"65",X"0C",X"01",X"65",X"0E",X"01",X"45",X"16",X"01",X"2F",X"16",X"19",X"00",X"18",X"01",
		X"6B",X"1A",X"01",X"6B",X"1C",X"01",X"6B",X"1E",X"01",X"4D",X"20",X"01",X"2F",X"22",X"81",X"08",
		X"26",X"01",X"25",X"28",X"01",X"45",X"2A",X"01",X"45",X"2C",X"01",X"45",X"2C",X"31",X"0E",X"2E",
		X"01",X"45",X"30",X"01",X"65",X"32",X"01",X"65",X"34",X"01",X"45",X"36",X"01",X"25",X"3A",X"81",
		X"0E",X"3C",X"99",X"0A",X"40",X"19",X"14",X"44",X"01",X"2F",X"46",X"49",X"06",X"46",X"01",X"4D",
		X"48",X"01",X"6B",X"4A",X"01",X"6B",X"4C",X"01",X"89",X"4E",X"01",X"6B",X"50",X"81",X"06",X"50",
		X"01",X"4D",X"58",X"01",X"69",X"5A",X"01",X"49",X"5C",X"01",X"49",X"5C",X"81",X"0F",X"5E",X"01",
		X"69",X"60",X"01",X"2D",X"64",X"19",X"00",X"64",X"81",X"08",X"66",X"81",X"0E",X"68",X"01",X"25",
		X"6A",X"01",X"45",X"6C",X"01",X"45",X"70",X"01",X"2F",X"72",X"01",X"2F",X"74",X"01",X"4D",X"76",
		X"01",X"4D",X"76",X"31",X"08",X"78",X"01",X"4D",X"7A",X"01",X"2F",X"7C",X"81",X"0A",X"7C",X"01",
		X"25",X"7E",X"01",X"25",X"80",X"19",X"14",X"80",X"01",X"45",X"86",X"61",X"0E",X"88",X"01",X"27",
		X"8E",X"01",X"2A",X"92",X"01",X"2A",X"96",X"81",X"0E",X"9C",X"81",X"06",X"9E",X"01",X"2E",X"A2",
		X"01",X"2A",X"A8",X"81",X"09",X"AE",X"31",X"0F",X"B0",X"01",X"28",X"B4",X"81",X"0C",X"B8",X"99",
		X"0C",X"BC",X"49",X"07",X"C2",X"01",X"2D",X"CA",X"01",X"45",X"CC",X"01",X"25",X"CE",X"81",X"0E",
		X"D4",X"01",X"2B",X"D8",X"61",X"06",X"DA",X"01",X"2E",X"DE",X"01",X"25",X"FF",X"FF",X"FF",X"00",
		X"00",X"00",X"20",X"00",X"6A",X"22",X"00",X"4C",X"26",X"00",X"25",X"28",X"00",X"45",X"2A",X"00",
		X"45",X"2C",X"00",X"25",X"2E",X"00",X"2F",X"30",X"00",X"2F",X"32",X"00",X"4D",X"3A",X"00",X"25",
		X"3C",X"00",X"45",X"3E",X"00",X"45",X"40",X"00",X"25",X"42",X"00",X"2F",X"44",X"00",X"4D",X"46",
		X"00",X"4D",X"48",X"80",X"08",X"48",X"00",X"2F",X"4C",X"00",X"2C",X"4E",X"00",X"4A",X"50",X"00",
		X"6A",X"52",X"00",X"2C",X"54",X"30",X"08",X"58",X"80",X"0E",X"5A",X"00",X"2B",X"5C",X"00",X"49",
		X"5E",X"00",X"49",X"60",X"00",X"49",X"62",X"00",X"2B",X"64",X"00",X"4B",X"66",X"00",X"4B",X"68",
		X"18",X"00",X"68",X"00",X"4D",X"6A",X"80",X"06",X"6A",X"00",X"4D",X"6E",X"00",X"25",X"6E",X"48",
		X"0E",X"70",X"00",X"25",X"72",X"00",X"65",X"74",X"00",X"65",X"76",X"00",X"45",X"78",X"00",X"45",
		X"7E",X"18",X"14",X"80",X"00",X"2F",X"82",X"00",X"4D",X"84",X"00",X"6B",X"86",X"00",X"6B",X"88",
		X"00",X"4D",X"8A",X"80",X"08",X"8A",X"00",X"2F",X"8E",X"80",X"0E",X"92",X"00",X"2B",X"94",X"00",
		X"49",X"96",X"00",X"49",X"98",X"00",X"2B",X"9C",X"30",X"08",X"9E",X"80",X"0E",X"A0",X"00",X"2B",
		X"A2",X"00",X"2B",X"A4",X"00",X"4B",X"A6",X"00",X"4B",X"A8",X"00",X"4B",X"AA",X"00",X"4D",X"AC",
		X"00",X"4D",X"B0",X"48",X"0E",X"B4",X"80",X"08",X"B6",X"18",X"00",X"B6",X"00",X"29",X"B8",X"00",
		X"47",X"BA",X"00",X"47",X"BC",X"00",X"47",X"BE",X"00",X"65",X"C0",X"00",X"45",X"C2",X"60",X"08",
		X"C2",X"80",X"0E",X"C6",X"00",X"2F",X"C8",X"00",X"4D",X"CA",X"00",X"4D",X"CC",X"00",X"6B",X"CE",
		X"00",X"6B",X"D0",X"00",X"4D",X"D2",X"00",X"2F",X"D4",X"48",X"0A",X"D8",X"00",X"2A",X"DA",X"00",
		X"4A",X"DA",X"80",X"0E",X"DC",X"00",X"4A",X"DE",X"00",X"6A",X"E0",X"00",X"6A",X"E4",X"98",X"0C",
		X"EE",X"18",X"14",X"F0",X"00",X"27",X"F2",X"00",X"65",X"F4",X"00",X"65",X"F6",X"00",X"65",X"F8",
		X"00",X"25",X"FC",X"18",X"00",X"00",X"01",X"2F",X"02",X"81",X"08",X"02",X"01",X"4D",X"04",X"01",
		X"4D",X"06",X"01",X"6B",X"08",X"01",X"4D",X"0A",X"01",X"4D",X"0C",X"01",X"2F",X"0E",X"31",X"08",
		X"12",X"01",X"25",X"14",X"01",X"45",X"16",X"01",X"65",X"16",X"81",X"0E",X"18",X"01",X"45",X"1E",
		X"01",X"2F",X"20",X"01",X"4D",X"22",X"01",X"4D",X"24",X"01",X"6B",X"26",X"01",X"4D",X"28",X"01",
		X"4D",X"2A",X"01",X"2F",X"2C",X"49",X"08",X"2C",X"81",X"0A",X"30",X"01",X"29",X"32",X"01",X"49",
		X"34",X"01",X"49",X"36",X"19",X"00",X"36",X"01",X"2B",X"38",X"01",X"4B",X"3A",X"01",X"6B",X"3C",
		X"01",X"4D",X"3E",X"61",X"2F",X"3E",X"01",X"2F",X"42",X"01",X"25",X"44",X"01",X"45",X"46",X"01",
		X"65",X"48",X"01",X"65",X"48",X"81",X"0E",X"4A",X"01",X"45",X"4C",X"01",X"25",X"50",X"49",X"08",
		X"54",X"01",X"2F",X"56",X"01",X"4D",X"58",X"81",X"0A",X"58",X"01",X"4D",X"5A",X"01",X"6B",X"5C",
		X"01",X"6B",X"5E",X"01",X"4D",X"60",X"01",X"2F",X"66",X"01",X"2D",X"68",X"81",X"06",X"68",X"01",
		X"4D",X"6A",X"01",X"4D",X"72",X"01",X"2B",X"74",X"81",X"06",X"74",X"01",X"6B",X"76",X"01",X"4D",
		X"7C",X"01",X"25",X"7E",X"01",X"25",X"80",X"01",X"45",X"80",X"81",X"0C",X"84",X"01",X"2B",X"86",
		X"01",X"47",X"88",X"01",X"27",X"8A",X"01",X"25",X"8E",X"81",X"0E",X"94",X"99",X"08",X"9C",X"61",
		X"0F",X"9E",X"81",X"08",X"A4",X"49",X"0D",X"A8",X"01",X"28",X"AC",X"81",X"0D",X"B0",X"81",X"09",
		X"B6",X"01",X"2A",X"B8",X"61",X"07",X"B8",X"01",X"2C",X"BA",X"01",X"2E",X"C0",X"01",X"27",X"C4",
		X"81",X"0F",X"C8",X"81",X"07",X"C8",X"49",X"0F",X"CC",X"99",X"08",X"D4",X"01",X"29",X"D6",X"01",
		X"25",X"DA",X"81",X"0B",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"6A",
		X"22",X"00",X"4C",X"26",X"00",X"25",X"28",X"00",X"45",X"2A",X"00",X"45",X"2C",X"00",X"25",X"32",
		X"98",X"0A",X"38",X"00",X"2F",X"3A",X"80",X"06",X"3E",X"00",X"4A",X"46",X"00",X"45",X"48",X"00",
		X"45",X"4A",X"00",X"25",X"4A",X"80",X"0D",X"52",X"00",X"2F",X"54",X"30",X"0B",X"58",X"80",X"08",
		X"5E",X"00",X"28",X"5E",X"00",X"2D",X"64",X"00",X"25",X"64",X"00",X"2A",X"64",X"00",X"2F",X"6C",
		X"00",X"29",X"70",X"00",X"2D",X"72",X"80",X"06",X"7A",X"00",X"25",X"7C",X"48",X"0B",X"80",X"00",
		X"27",X"84",X"98",X"0A",X"8C",X"80",X"07",X"90",X"00",X"27",X"92",X"00",X"2F",X"94",X"30",X"0B",
		X"9A",X"00",X"25",X"9E",X"00",X"2A",X"A4",X"00",X"68",X"A6",X"00",X"68",X"AE",X"60",X"06",X"AE",
		X"00",X"2F",X"B2",X"00",X"29",X"B8",X"00",X"25",X"BA",X"00",X"2D",X"C0",X"00",X"2D",X"C2",X"00",
		X"2B",X"C4",X"00",X"29",X"CA",X"00",X"2F",X"CE",X"00",X"29",X"D0",X"00",X"29",X"D2",X"00",X"27",
		X"D4",X"00",X"25",X"D6",X"00",X"2F",X"D8",X"00",X"4D",X"DA",X"80",X"08",X"DE",X"00",X"28",X"E4",
		X"00",X"2B",X"EA",X"98",X"06",X"EA",X"00",X"2F",X"F0",X"80",X"0B",X"F4",X"00",X"68",X"FC",X"00",
		X"2A",X"FC",X"00",X"2F",X"06",X"01",X"25",X"06",X"01",X"2A",X"08",X"81",X"0E",X"10",X"01",X"89",
		X"12",X"49",X"06",X"12",X"01",X"6B",X"14",X"01",X"4D",X"16",X"01",X"2F",X"1A",X"01",X"27",X"1C",
		X"01",X"47",X"1E",X"01",X"67",X"20",X"01",X"67",X"22",X"01",X"47",X"24",X"01",X"27",X"26",X"61",
		X"0E",X"2C",X"99",X"0B",X"30",X"01",X"28",X"34",X"01",X"2F",X"3A",X"01",X"65",X"3C",X"01",X"65",
		X"3E",X"01",X"45",X"40",X"01",X"25",X"42",X"81",X"0D",X"48",X"81",X"0B",X"4C",X"01",X"4A",X"4E",
		X"31",X"06",X"4E",X"01",X"2C",X"52",X"01",X"2F",X"58",X"01",X"27",X"58",X"01",X"2D",X"5A",X"01",
		X"25",X"5A",X"01",X"2F",X"62",X"01",X"68",X"64",X"01",X"2A",X"6C",X"01",X"65",X"70",X"81",X"0B",
		X"74",X"01",X"89",X"7A",X"81",X"06",X"7E",X"01",X"29",X"80",X"01",X"48",X"82",X"01",X"28",X"84",
		X"01",X"29",X"86",X"01",X"2A",X"88",X"01",X"2B",X"8A",X"01",X"2C",X"8C",X"01",X"2C",X"8E",X"01",
		X"2C",X"90",X"01",X"2C",X"90",X"81",X"0F",X"92",X"01",X"27",X"92",X"01",X"2C",X"94",X"01",X"26",
		X"94",X"01",X"2D",X"9C",X"01",X"48",X"9C",X"01",X"2F",X"A0",X"99",X"06",X"A6",X"01",X"2C",X"AC",
		X"01",X"27",X"B0",X"01",X"2F",X"B2",X"61",X"08",X"B2",X"01",X"4D",X"B4",X"01",X"4D",X"BA",X"01",
		X"25",X"BC",X"01",X"45",X"BC",X"01",X"2C",X"BE",X"01",X"45",X"C4",X"01",X"2A",X"C8",X"99",X"0C",
		X"CC",X"01",X"45",X"CE",X"01",X"25",X"D0",X"61",X"0A",X"D8",X"01",X"25",X"D8",X"01",X"29",X"DA",
		X"81",X"0D",X"DE",X"01",X"49",X"DE",X"01",X"2F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"20",X"00",X"6A",X"22",X"00",X"4C",X"26",X"00",X"25",X"26",X"00",X"45",
		X"2A",X"00",X"45",X"2C",X"00",X"25",X"30",X"00",X"29",X"32",X"00",X"2A",X"34",X"00",X"2B",X"3C",
		X"80",X"07",X"3C",X"00",X"2F",X"40",X"98",X"07",X"48",X"00",X"25",X"4A",X"00",X"2B",X"4C",X"00",
		X"2C",X"4E",X"00",X"2D",X"54",X"00",X"26",X"54",X"48",X"0B",X"54",X"00",X"2F",X"56",X"00",X"27",
		X"58",X"00",X"28",X"5A",X"00",X"26",X"5C",X"00",X"25",X"62",X"80",X"0C",X"66",X"00",X"68",X"68",
		X"00",X"49",X"6A",X"00",X"2A",X"72",X"30",X"0C",X"72",X"00",X"2F",X"74",X"00",X"28",X"76",X"00",
		X"29",X"78",X"00",X"2A",X"7A",X"00",X"2B",X"7C",X"00",X"2C",X"7E",X"00",X"26",X"82",X"00",X"2F",
		X"86",X"00",X"28",X"8C",X"00",X"2B",X"90",X"00",X"2F",X"92",X"00",X"4D",X"96",X"80",X"08",X"98",
		X"00",X"26",X"9A",X"00",X"26",X"9C",X"00",X"25",X"9E",X"80",X"0D",X"A4",X"00",X"46",X"A4",X"80",
		X"0D",X"AC",X"80",X"08",X"AE",X"00",X"4C",X"B4",X"80",X"0D",X"B8",X"00",X"2A",X"BE",X"80",X"07",
		X"C2",X"00",X"46",X"C4",X"80",X"0D",X"CC",X"00",X"2A",X"CC",X"60",X"0D",X"D0",X"80",X"06",X"D6",
		X"00",X"4C",X"DC",X"80",X"08",X"E0",X"00",X"2A",X"E2",X"80",X"0E",X"EA",X"00",X"46",X"F0",X"80",
		X"0A",X"F4",X"00",X"2A",X"FC",X"80",X"06",X"FE",X"00",X"4C",X"06",X"81",X"0C",X"08",X"01",X"2A",
		X"0E",X"81",X"06",X"12",X"01",X"46",X"12",X"61",X"0D",X"1C",X"01",X"28",X"1C",X"31",X"0C",X"26",
		X"49",X"07",X"26",X"01",X"2C",X"2E",X"01",X"2F",X"30",X"01",X"26",X"30",X"31",X"0B",X"38",X"49",
		X"07",X"38",X"01",X"2D",X"42",X"31",X"0C",X"44",X"01",X"26",X"4A",X"01",X"2F",X"52",X"01",X"29",
		X"52",X"01",X"2E",X"56",X"81",X"06",X"58",X"01",X"27",X"58",X"01",X"2C",X"5E",X"01",X"29",X"5E",
		X"01",X"2E",X"62",X"01",X"25",X"66",X"01",X"2D",X"68",X"01",X"29",X"6C",X"01",X"25",X"6E",X"01",
		X"45",X"72",X"99",X"0B",X"7A",X"01",X"29",X"7C",X"01",X"29",X"80",X"01",X"29",X"84",X"01",X"29",
		X"88",X"01",X"29",X"8A",X"61",X"0C",X"8E",X"01",X"29",X"92",X"01",X"29",X"94",X"61",X"0E",X"96",
		X"01",X"29",X"98",X"61",X"06",X"9A",X"01",X"29",X"9E",X"99",X"06",X"A6",X"01",X"27",X"A8",X"81",
		X"06",X"AE",X"61",X"0E",X"B0",X"01",X"49",X"B6",X"81",X"0E",X"B8",X"01",X"27",X"B8",X"01",X"2D",
		X"BE",X"01",X"2A",X"C0",X"01",X"2A",X"C0",X"81",X"0D",X"C4",X"01",X"25",X"C6",X"01",X"45",X"C6",
		X"01",X"2D",X"C8",X"01",X"25",X"C8",X"01",X"2D",X"CA",X"01",X"2C",X"CC",X"01",X"2B",X"D2",X"01",
		X"27",X"D4",X"01",X"29",X"D4",X"01",X"2F",X"D6",X"81",X"0C",X"C2",X"01",X"2F",X"DA",X"01",X"27",
		X"DA",X"01",X"2C",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"20",
		X"00",X"6A",X"22",X"00",X"4C",X"26",X"00",X"25",X"28",X"00",X"45",X"2A",X"00",X"45",X"2C",X"00",
		X"25",X"30",X"00",X"2F",X"32",X"00",X"4D",X"34",X"00",X"6B",X"36",X"80",X"06",X"36",X"00",X"89",
		X"38",X"00",X"6B",X"3A",X"00",X"4D",X"3C",X"00",X"2F",X"3E",X"00",X"28",X"40",X"00",X"29",X"42",
		X"00",X"2A",X"44",X"80",X"0D",X"46",X"00",X"25",X"48",X"00",X"45",X"4E",X"00",X"2A",X"50",X"80",
		X"0E",X"52",X"00",X"2A",X"56",X"00",X"2A",X"5C",X"80",X"06",X"5E",X"00",X"2A",X"62",X"00",X"2A",
		X"64",X"48",X"06",X"66",X"00",X"2A",X"6A",X"00",X"2C",X"6C",X"00",X"26",X"6E",X"00",X"25",X"76",
		X"00",X"48",X"76",X"80",X"0E",X"7A",X"00",X"2A",X"7E",X"00",X"25",X"7E",X"00",X"2A",X"82",X"00",
		X"2A",X"8A",X"80",X"06",X"8A",X"00",X"2A",X"8E",X"00",X"2A",X"92",X"00",X"2C",X"94",X"00",X"2F",
		X"96",X"80",X"07",X"9A",X"00",X"25",X"9C",X"98",X"07",X"9E",X"60",X"0D",X"A2",X"00",X"2A",X"A4",
		X"00",X"4A",X"A4",X"80",X"0F",X"AA",X"00",X"2F",X"AE",X"00",X"25",X"B0",X"00",X"45",X"B2",X"00",
		X"25",X"B2",X"00",X"2F",X"B4",X"00",X"4D",X"B6",X"00",X"89",X"B8",X"00",X"6B",X"BA",X"00",X"4D",
		X"BC",X"00",X"25",X"BC",X"00",X"2F",X"C2",X"98",X"0A",X"C8",X"00",X"25",X"CA",X"00",X"45",X"CC",
		X"00",X"45",X"CE",X"00",X"45",X"CE",X"00",X"2C",X"D0",X"00",X"25",X"D6",X"00",X"2A",X"D6",X"00",
		X"2F",X"D8",X"00",X"25",X"DC",X"00",X"45",X"DE",X"00",X"2C",X"E2",X"00",X"2D",X"E6",X"00",X"29",
		X"EA",X"00",X"25",X"EA",X"80",X"0B",X"EC",X"00",X"45",X"EE",X"00",X"65",X"F0",X"00",X"65",X"F2",
		X"00",X"65",X"F4",X"00",X"65",X"F6",X"00",X"45",X"F6",X"00",X"2F",X"F8",X"00",X"25",X"F8",X"00",
		X"4D",X"FA",X"00",X"6B",X"FC",X"00",X"6B",X"FE",X"00",X"6B",X"00",X"01",X"6B",X"02",X"81",X"06",
		X"02",X"01",X"4D",X"04",X"01",X"2F",X"06",X"01",X"29",X"08",X"01",X"48",X"0A",X"01",X"48",X"0C",
		X"01",X"67",X"0E",X"01",X"67",X"10",X"01",X"67",X"12",X"01",X"48",X"14",X"01",X"29",X"18",X"01",
		X"25",X"1A",X"01",X"25",X"1A",X"99",X"0C",X"1C",X"01",X"25",X"1E",X"01",X"45",X"20",X"01",X"45",
		X"22",X"01",X"45",X"22",X"49",X"0D",X"24",X"01",X"65",X"26",X"01",X"65",X"28",X"01",X"85",X"2A",
		X"01",X"65",X"2C",X"01",X"65",X"2E",X"01",X"45",X"2E",X"01",X"2F",X"30",X"01",X"25",X"30",X"01",
		X"4D",X"32",X"01",X"6B",X"34",X"01",X"4D",X"36",X"01",X"2F",X"3A",X"01",X"25",X"3C",X"01",X"45",
		X"3C",X"01",X"4D",X"3E",X"01",X"25",X"3E",X"01",X"2F",X"44",X"01",X"26",X"48",X"61",X"0C",X"4E",
		X"61",X"07",X"50",X"01",X"2C",X"56",X"61",X"0C",X"5C",X"01",X"28",X"5E",X"61",X"0E",X"62",X"99",
		X"09",X"64",X"61",X"06",X"6C",X"61",X"0B",X"6C",X"01",X"2F",X"6E",X"01",X"26",X"74",X"61",X"06",
		X"76",X"01",X"2C",X"7C",X"61",X"0E",X"7E",X"01",X"2A",X"82",X"61",X"07",X"88",X"01",X"25",X"88",
		X"01",X"2F",X"8A",X"01",X"45",X"8A",X"01",X"4D",X"8C",X"01",X"25",X"8C",X"01",X"2F",X"94",X"81",
		X"08",X"98",X"31",X"0D",X"9E",X"49",X"07",X"A6",X"31",X"0B",X"AC",X"01",X"2D",X"AE",X"01",X"25",
		X"B2",X"99",X"07",X"B2",X"49",X"0D",X"B8",X"49",X"0B",X"BC",X"01",X"27",X"C0",X"01",X"2F",X"C2",
		X"31",X"07",X"C2",X"01",X"4D",X"C4",X"01",X"2F",X"CA",X"01",X"26",X"CA",X"49",X"0D",X"D0",X"61",
		X"07",X"D0",X"01",X"2C",X"D6",X"61",X"0B",X"C2",X"01",X"2F",X"D8",X"01",X"25",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"6A",X"22",X"00",X"4C",X"26",
		X"00",X"25",X"28",X"00",X"45",X"2A",X"00",X"45",X"2C",X"00",X"25",X"32",X"00",X"2F",X"36",X"00",
		X"4D",X"38",X"00",X"29",X"38",X"00",X"2F",X"40",X"98",X"05",X"40",X"00",X"2C",X"42",X"00",X"2D",
		X"44",X"00",X"2E",X"46",X"80",X"09",X"46",X"00",X"2F",X"4A",X"00",X"29",X"4C",X"00",X"29",X"4E",
		X"00",X"2A",X"4E",X"00",X"2F",X"50",X"00",X"2A",X"54",X"00",X"25",X"56",X"00",X"25",X"58",X"00",
		X"2F",X"5A",X"80",X"0A",X"5A",X"00",X"2E",X"5E",X"00",X"28",X"62",X"00",X"2C",X"66",X"98",X"07",
		X"6A",X"00",X"2F",X"6E",X"00",X"25",X"74",X"00",X"28",X"7A",X"00",X"25",X"7E",X"00",X"2F",X"80",
		X"00",X"28",X"84",X"80",X"0B",X"86",X"00",X"2C",X"88",X"00",X"2A",X"8E",X"00",X"25",X"90",X"00",
		X"45",X"90",X"98",X"09",X"90",X"80",X"0F",X"92",X"00",X"25",X"98",X"00",X"2F",X"9C",X"00",X"2B",
		X"9E",X"80",X"06",X"A2",X"00",X"28",X"A2",X"00",X"2D",X"A8",X"00",X"25",X"A8",X"00",X"2F",X"AE",
		X"00",X"27",X"B2",X"00",X"2C",X"B6",X"00",X"29",X"B8",X"00",X"2F",X"BA",X"48",X"0C",X"BC",X"00",
		X"25",X"C4",X"98",X"0C",X"C6",X"00",X"28",X"CC",X"00",X"26",X"CC",X"00",X"2F",X"D0",X"00",X"2A",
		X"D6",X"30",X"0F",X"D8",X"00",X"49",X"DC",X"00",X"25",X"DE",X"00",X"2F",X"E0",X"00",X"2F",X"E4",
		X"00",X"27",X"E8",X"00",X"2D",X"EC",X"00",X"29",X"EE",X"00",X"2B",X"F2",X"00",X"25",X"F2",X"00",
		X"2F",X"F4",X"80",X"0A",X"F8",X"00",X"27",X"FA",X"00",X"2C",X"FE",X"00",X"25",X"FE",X"98",X"09",
		X"FE",X"80",X"0F",X"04",X"01",X"2F",X"08",X"01",X"28",X"0C",X"01",X"2C",X"10",X"01",X"25",X"12",
		X"49",X"0A",X"14",X"01",X"2F",X"16",X"01",X"27",X"1A",X"61",X"0C",X"20",X"61",X"08",X"26",X"31",
		X"0C",X"2A",X"01",X"68",X"30",X"01",X"25",X"30",X"01",X"2F",X"34",X"01",X"2A",X"34",X"81",X"0F",
		X"38",X"01",X"25",X"38",X"01",X"2F",X"3E",X"01",X"28",X"3E",X"01",X"2C",X"40",X"81",X"0F",X"44",
		X"01",X"25",X"44",X"01",X"2F",X"48",X"81",X"05",X"48",X"01",X"2A",X"4C",X"01",X"25",X"4C",X"01",
		X"2F",X"52",X"01",X"28",X"52",X"01",X"2C",X"54",X"81",X"0F",X"58",X"01",X"25",X"58",X"01",X"2F",
		X"5C",X"01",X"2A",X"60",X"01",X"25",X"60",X"01",X"2F",X"62",X"81",X"08",X"66",X"01",X"2A",X"6C",
		X"01",X"25",X"6C",X"99",X"0B",X"74",X"01",X"25",X"74",X"81",X"09",X"76",X"01",X"45",X"80",X"81",
		X"07",X"80",X"01",X"2B",X"84",X"01",X"2B",X"88",X"81",X"06",X"88",X"01",X"2B",X"8C",X"01",X"2B",
		X"90",X"01",X"2B",X"94",X"01",X"2B",X"98",X"01",X"2B",X"9C",X"01",X"2B",X"A0",X"01",X"29",X"A4",
		X"01",X"26",X"AC",X"61",X"07",X"AE",X"99",X"0A",X"B2",X"01",X"25",X"B4",X"01",X"25",X"B4",X"01",
		X"2D",X"B6",X"01",X"45",X"B8",X"01",X"65",X"BA",X"01",X"85",X"BC",X"01",X"65",X"BE",X"01",X"45",
		X"BE",X"01",X"2F",X"C0",X"01",X"45",X"C0",X"01",X"4D",X"C2",X"01",X"45",X"C2",X"01",X"2F",X"C4",
		X"01",X"45",X"C4",X"01",X"2F",X"C6",X"01",X"45",X"C8",X"01",X"85",X"CA",X"01",X"65",X"CC",X"01",
		X"45",X"CC",X"01",X"2F",X"CE",X"01",X"25",X"CE",X"01",X"4D",X"D0",X"01",X"2F",X"D4",X"01",X"2A",
		X"D8",X"61",X"07",X"DA",X"01",X"2F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"20",X"00",X"6A",X"22",X"00",X"4C",X"26",X"00",X"25",X"28",X"00",X"45",X"2A",X"00",
		X"45",X"2C",X"00",X"25",X"34",X"00",X"2B",X"36",X"00",X"49",X"38",X"00",X"49",X"3A",X"00",X"49",
		X"3C",X"00",X"2B",X"3C",X"30",X"0E",X"40",X"00",X"25",X"40",X"80",X"08",X"40",X"00",X"6B",X"42",
		X"00",X"25",X"42",X"00",X"4D",X"44",X"00",X"45",X"44",X"00",X"2F",X"46",X"00",X"65",X"46",X"00",
		X"2F",X"48",X"00",X"65",X"48",X"00",X"2F",X"4A",X"00",X"45",X"4A",X"80",X"0C",X"4A",X"00",X"2F",
		X"4C",X"00",X"25",X"4C",X"00",X"4D",X"4E",X"00",X"25",X"4E",X"00",X"6B",X"50",X"00",X"6B",X"52",
		X"00",X"6B",X"54",X"80",X"07",X"54",X"00",X"4D",X"56",X"00",X"2F",X"5A",X"00",X"29",X"5C",X"00",
		X"29",X"5E",X"80",X"07",X"5E",X"00",X"29",X"60",X"00",X"2A",X"62",X"00",X"2B",X"64",X"00",X"25",
		X"64",X"00",X"2C",X"66",X"00",X"26",X"66",X"00",X"2D",X"68",X"00",X"28",X"68",X"80",X"0B",X"68",
		X"00",X"2F",X"6E",X"00",X"2B",X"70",X"00",X"2B",X"72",X"98",X"05",X"72",X"80",X"0E",X"74",X"00",
		X"2A",X"78",X"00",X"28",X"78",X"00",X"2F",X"7A",X"00",X"27",X"7A",X"00",X"2E",X"7C",X"80",X"0A",
		X"7E",X"00",X"26",X"80",X"00",X"25",X"80",X"00",X"2C",X"82",X"00",X"25",X"84",X"00",X"25",X"84",
		X"00",X"2B",X"86",X"00",X"25",X"86",X"80",X"08",X"86",X"00",X"2B",X"8A",X"00",X"2B",X"8C",X"00",
		X"25",X"8C",X"00",X"2B",X"8E",X"00",X"2C",X"90",X"00",X"26",X"90",X"80",X"09",X"90",X"00",X"2C",
		X"92",X"00",X"4D",X"94",X"00",X"27",X"94",X"00",X"2F",X"98",X"00",X"2A",X"98",X"00",X"2F",X"9A",
		X"00",X"2A",X"9A",X"80",X"0C",X"9C",X"00",X"2A",X"9E",X"00",X"2A",X"A0",X"00",X"2A",X"A2",X"00",
		X"2A",X"A2",X"80",X"0D",X"AA",X"00",X"25",X"AA",X"00",X"2A",X"AC",X"00",X"25",X"AC",X"00",X"29",
		X"AE",X"00",X"25",X"AE",X"00",X"29",X"B0",X"00",X"25",X"B0",X"00",X"29",X"B2",X"00",X"25",X"B2",
		X"00",X"29",X"B4",X"00",X"25",X"B4",X"00",X"29",X"B6",X"00",X"25",X"B6",X"00",X"29",X"B8",X"00",
		X"25",X"B8",X"80",X"07",X"B8",X"00",X"29",X"BC",X"00",X"2F",X"C0",X"00",X"26",X"C2",X"00",X"26",
		X"C2",X"98",X"0B",X"D0",X"00",X"2C",X"D2",X"00",X"2B",X"D4",X"00",X"48",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"21",X"32",X"80",X"CB",X"7E",X"20",X"20",X"CB",X"FE",X"3E",X"E4",X"11",X"A1",X"90",
		X"01",X"18",X"00",X"00",X"00",X"00",X"11",X"A1",X"90",X"3E",X"08",X"01",X"01",X"18",X"00",X"00",
		X"00",X"21",X"00",X"03",X"22",X"1B",X"80",X"18",X"7F",X"21",X"36",X"80",X"CB",X"76",X"C0",X"3A",
		X"30",X"80",X"FE",X"06",X"20",X"05",X"21",X"32",X"80",X"CB",X"EE",X"2A",X"30",X"80",X"ED",X"5B",
		X"33",X"80",X"19",X"22",X"33",X"80",X"11",X"03",X"00",X"B7",X"ED",X"52",X"28",X"02",X"38",X"58",
		X"2A",X"1B",X"80",X"00",X"22",X"1B",X"80",X"11",X"C0",X"00",X"B7",X"ED",X"52",X"20",X"0D",X"21",
		X"32",X"80",X"CB",X"6E",X"20",X"06",X"01",X"0D",X"01",X"CD",X"75",X"48",X"2A",X"1B",X"80",X"7D",
		X"0F",X"0F",X"E6",X"07",X"C6",X"DC",X"F5",X"3E",X"03",X"A4",X"67",X"3E",X"E0",X"A5",X"6F",X"01",
		X"A1",X"90",X"09",X"F1",X"00",X"2A",X"1B",X"80",X"7C",X"B5",X"20",X"10",X"21",X"36",X"80",X"CB",
		X"F6",X"21",X"23",X"80",X"CB",X"5E",X"C0",X"21",X"16",X"80",X"CB",X"DE",X"2A",X"33",X"80",X"11",
		X"03",X"00",X"B7",X"ED",X"52",X"22",X"33",X"80",X"3E",X"0E",X"EF",X"C9",X"21",X"30",X"80",X"CB",
		X"7E",X"20",X"24",X"CB",X"FE",X"2A",X"21",X"80",X"22",X"31",X"80",X"3E",X"C0",X"32",X"36",X"80",
		X"11",X"A2",X"90",X"01",X"18",X"00",X"3E",X"E4",X"CD",X"13",X"05",X"11",X"A3",X"90",X"01",X"01",
		X"18",X"3E",X"09",X"CD",X"32",X"05",X"C9",X"3A",X"36",X"80",X"B7",X"20",X"27",X"21",X"23",X"80",
		X"CB",X"DE",X"AF",X"32",X"A1",X"81",X"32",X"A9",X"81",X"32",X"B1",X"81",X"32",X"9F",X"81",X"3E",
		X"07",X"D3",X"08",X"3E",X"3F",X"32",X"A0",X"81",X"D3",X"09",X"01",X"03",X"03",X"CD",X"75",X"48",
		X"3E",X"0D",X"D7",X"C9",X"2A",X"21",X"80",X"ED",X"5B",X"33",X"80",X"44",X"4D",X"ED",X"52",X"C8",
		X"38",X"16",X"3E",X"07",X"BD",X"30",X"11",X"ED",X"43",X"33",X"80",X"21",X"14",X"80",X"CB",X"46",
		X"20",X"06",X"3E",X"0F",X"21",X"01",X"00",X"E7",X"ED",X"5B",X"31",X"80",X"2A",X"21",X"80",X"22",
		X"31",X"80",X"01",X"1C",X"00",X"B7",X"ED",X"42",X"30",X"05",X"21",X"14",X"80",X"CB",X"C6",X"2A",
		X"31",X"80",X"B7",X"ED",X"52",X"C8",X"21",X"35",X"80",X"38",X"03",X"34",X"18",X"01",X"35",X"3E",
		X"14",X"86",X"20",X"12",X"77",X"21",X"36",X"80",X"34",X"7E",X"E6",X"07",X"20",X"13",X"3E",X"E4",
		X"F5",X"7E",X"D6",X"08",X"18",X"12",X"FE",X"28",X"C0",X"AF",X"32",X"35",X"80",X"21",X"36",X"80",
		X"35",X"3E",X"07",X"A6",X"C6",X"DC",X"F5",X"7E",X"E6",X"F8",X"6F",X"26",X"00",X"29",X"29",X"11",
		X"A2",X"90",X"19",X"F1",X"77",X"EB",X"01",X"01",X"01",X"3E",X"09",X"CD",X"32",X"05",X"C9",X"21",
		X"32",X"80",X"CB",X"46",X"20",X"07",X"CB",X"C6",X"3A",X"2F",X"80",X"EF",X"C9",X"C3",X"5C",X"52",
		X"00",X"CB",X"CE",X"2A",X"30",X"80",X"22",X"34",X"80",X"21",X"07",X"27",X"22",X"36",X"80",X"3A",
		X"21",X"80",X"32",X"38",X"80",X"2E",X"02",X"CD",X"54",X"01",X"38",X"0E",X"2A",X"34",X"80",X"ED",
		X"4B",X"36",X"80",X"11",X"65",X"35",X"CD",X"92",X"01",X"C9",X"3E",X"0C",X"D7",X"C9",X"3A",X"33",
		X"80",X"E6",X"03",X"20",X"27",X"21",X"32",X"80",X"CB",X"6E",X"20",X"20",X"2A",X"34",X"80",X"11",
		X"04",X"04",X"19",X"01",X"08",X"18",X"CD",X"D0",X"3E",X"30",X"11",X"C3",X"18",X"52",X"CB",X"EE",
		X"3E",X"0E",X"21",X"00",X"01",X"E7",X"01",X"08",X"01",X"CD",X"75",X"48",X"21",X"33",X"80",X"34",
		X"7E",X"E6",X"03",X"21",X"32",X"80",X"20",X"04",X"CB",X"DE",X"18",X"02",X"CB",X"9E",X"CD",X"70",
		X"43",X"21",X"32",X"80",X"CB",X"76",X"C2",X"36",X"35",X"21",X"34",X"80",X"3E",X"50",X"BE",X"38",
		X"13",X"21",X"32",X"80",X"CB",X"F6",X"3A",X"30",X"80",X"ED",X"44",X"21",X"34",X"80",X"86",X"28",
		X"99",X"3D",X"28",X"96",X"3A",X"33",X"80",X"E6",X"0F",X"C2",X"C5",X"34",X"21",X"3D",X"80",X"34",
		X"7E",X"E6",X"03",X"4F",X"06",X"00",X"21",X"69",X"35",X"09",X"3E",X"9C",X"86",X"0F",X"0F",X"32",
		X"37",X"80",X"C3",X"C5",X"34",X"00",X"00",X"00",X"10",X"00",X"08",X"10",X"18",X"21",X"32",X"80",
		X"CB",X"5E",X"20",X"4B",X"CB",X"DE",X"01",X"00",X"03",X"CD",X"75",X"48",X"21",X"00",X"00",X"22",
		X"1D",X"80",X"22",X"21",X"80",X"21",X"18",X"00",X"22",X"1F",X"80",X"3E",X"48",X"32",X"1D",X"80",
		X"CD",X"EA",X"38",X"3E",X"20",X"32",X"39",X"80",X"3E",X"02",X"11",X"BE",X"39",X"CD",X"51",X"39",
		X"3E",X"20",X"32",X"39",X"80",X"32",X"3A",X"80",X"AF",X"32",X"2D",X"80",X"32",X"2A",X"80",X"21",
		X"16",X"80",X"CB",X"76",X"21",X"19",X"80",X"28",X"01",X"23",X"35",X"CD",X"DC",X"0C",X"C9",X"2A",
		X"21",X"80",X"11",X"10",X"01",X"B7",X"ED",X"52",X"38",X"05",X"21",X"14",X"80",X"CB",X"86",X"21",
		X"16",X"80",X"CB",X"5E",X"28",X"23",X"21",X"3E",X"80",X"CB",X"56",X"20",X"36",X"CB",X"D6",X"AF",
		X"32",X"9F",X"81",X"32",X"A1",X"81",X"32",X"A9",X"81",X"32",X"B1",X"81",X"3E",X"07",X"D3",X"08",
		X"3E",X"3F",X"32",X"A0",X"81",X"D3",X"09",X"18",X"1A",X"21",X"3E",X"80",X"CB",X"5E",X"20",X"13",
		X"3A",X"9F",X"81",X"B7",X"20",X"0D",X"01",X"06",X"02",X"CD",X"75",X"48",X"38",X"05",X"21",X"3E",
		X"80",X"CB",X"DE",X"21",X"14",X"80",X"CB",X"56",X"28",X"0F",X"3A",X"23",X"80",X"E6",X"FC",X"CB",
		X"D7",X"32",X"23",X"80",X"21",X"32",X"80",X"CB",X"EE",X"21",X"23",X"80",X"CB",X"5E",X"28",X"23",
		X"CB",X"9E",X"3E",X"FF",X"11",X"A5",X"88",X"01",X"16",X"00",X"CD",X"06",X"05",X"3E",X"0F",X"21",
		X"00",X"00",X"E7",X"3E",X"01",X"D7",X"21",X"16",X"80",X"CB",X"76",X"21",X"19",X"80",X"28",X"01",
		X"23",X"34",X"C9",X"21",X"16",X"80",X"CB",X"5E",X"C2",X"75",X"37",X"21",X"32",X"80",X"CB",X"7E",
		X"C2",X"ED",X"37",X"21",X"33",X"80",X"7E",X"E6",X"03",X"20",X"1A",X"2B",X"CB",X"6E",X"CC",X"1B",
		X"02",X"21",X"14",X"80",X"CB",X"46",X"20",X"0D",X"3A",X"33",X"80",X"E6",X"04",X"20",X"06",X"3E",
		X"0E",X"21",X"01",X"00",X"E7",X"21",X"23",X"80",X"CB",X"56",X"11",X"A7",X"3C",X"21",X"93",X"3C",
		X"20",X"06",X"11",X"F2",X"3C",X"21",X"9D",X"3C",X"06",X"04",X"3A",X"1F",X"80",X"BE",X"30",X"04",
		X"23",X"23",X"10",X"F9",X"06",X"00",X"23",X"4E",X"EB",X"09",X"3A",X"2D",X"80",X"4F",X"87",X"81",
		X"4F",X"09",X"EB",X"CD",X"60",X"3C",X"B7",X"28",X"05",X"21",X"3E",X"80",X"CB",X"FE",X"2A",X"21",
		X"80",X"06",X"00",X"CB",X"7F",X"28",X"01",X"05",X"4F",X"09",X"22",X"21",X"80",X"13",X"CD",X"60",
		X"3C",X"B7",X"28",X"05",X"21",X"3E",X"80",X"CB",X"FE",X"21",X"1F",X"80",X"86",X"77",X"13",X"CD",
		X"60",X"3C",X"B7",X"28",X"05",X"21",X"3E",X"80",X"CB",X"FE",X"21",X"1D",X"80",X"86",X"77",X"21",
		X"3E",X"80",X"CB",X"7E",X"28",X"0C",X"CB",X"BE",X"3A",X"33",X"80",X"E6",X"03",X"20",X"03",X"CD",
		X"16",X"3B",X"21",X"23",X"80",X"CB",X"56",X"28",X"12",X"CB",X"4E",X"28",X"05",X"CD",X"34",X"39",
		X"18",X"0C",X"CB",X"46",X"28",X"05",X"CD",X"29",X"39",X"18",X"03",X"CD",X"0F",X"39",X"11",X"BE",
		X"39",X"CD",X"51",X"39",X"21",X"23",X"80",X"CB",X"56",X"28",X"0B",X"3A",X"2D",X"80",X"11",X"B4",
		X"39",X"CD",X"80",X"39",X"18",X"0B",X"3E",X"FF",X"11",X"A5",X"88",X"01",X"16",X"00",X"CD",X"06",
		X"05",X"CD",X"EA",X"38",X"21",X"16",X"80",X"CB",X"4E",X"28",X"25",X"21",X"32",X"80",X"CB",X"FE",
		X"3E",X"FF",X"11",X"A5",X"88",X"01",X"16",X"00",X"CD",X"06",X"05",X"AF",X"32",X"33",X"80",X"3A",
		X"23",X"80",X"E6",X"F8",X"32",X"23",X"80",X"3A",X"32",X"80",X"E6",X"F8",X"32",X"32",X"80",X"C9",
		X"21",X"33",X"80",X"35",X"C9",X"3E",X"FF",X"11",X"A5",X"88",X"01",X"16",X"00",X"CD",X"06",X"05",
		X"21",X"3E",X"80",X"CB",X"66",X"20",X"08",X"CB",X"E6",X"01",X"08",X"01",X"CD",X"75",X"48",X"21",
		X"31",X"80",X"CB",X"7E",X"20",X"0D",X"21",X"33",X"80",X"34",X"7E",X"E6",X"0F",X"C0",X"21",X"31",
		X"80",X"CB",X"FE",X"21",X"3E",X"80",X"CB",X"6E",X"20",X"08",X"CB",X"EE",X"01",X"09",X"01",X"CD",
		X"75",X"48",X"3A",X"36",X"80",X"E6",X"E0",X"07",X"07",X"07",X"21",X"3A",X"80",X"BE",X"28",X"06",
		X"11",X"12",X"3A",X"CD",X"56",X"39",X"06",X"60",X"3A",X"36",X"80",X"B8",X"20",X"1A",X"21",X"14",
		X"80",X"CB",X"F6",X"3E",X"01",X"D7",X"21",X"00",X"88",X"11",X"01",X"88",X"01",X"FF",X"00",X"36",
		X"FF",X"ED",X"B0",X"21",X"32",X"00",X"F7",X"C9",X"21",X"36",X"80",X"34",X"C9",X"CD",X"1B",X"02",
		X"3A",X"34",X"80",X"E6",X"03",X"20",X"06",X"3E",X"0E",X"21",X"02",X"00",X"E7",X"21",X"34",X"80",
		X"34",X"21",X"32",X"80",X"CB",X"76",X"20",X"6B",X"CD",X"EA",X"38",X"11",X"BE",X"39",X"3E",X"02",
		X"CD",X"51",X"39",X"ED",X"5B",X"21",X"80",X"2A",X"1F",X"80",X"19",X"ED",X"5B",X"26",X"80",X"B7",
		X"ED",X"52",X"28",X"12",X"30",X"09",X"2A",X"21",X"80",X"23",X"22",X"21",X"80",X"18",X"07",X"2A",
		X"21",X"80",X"2B",X"22",X"21",X"80",X"ED",X"5B",X"24",X"80",X"2A",X"1D",X"80",X"B7",X"ED",X"52",
		X"28",X"0C",X"30",X"06",X"21",X"1D",X"80",X"34",X"18",X"04",X"21",X"1D",X"80",X"35",X"2A",X"24",
		X"80",X"ED",X"5B",X"1D",X"80",X"B7",X"ED",X"52",X"C0",X"ED",X"5B",X"26",X"80",X"2A",X"1F",X"80",
		X"ED",X"4B",X"21",X"80",X"09",X"B7",X"ED",X"52",X"C0",X"21",X"32",X"80",X"CB",X"F6",X"AF",X"32",
		X"34",X"80",X"C9",X"3A",X"34",X"80",X"E6",X"78",X"0F",X"0F",X"0F",X"32",X"37",X"80",X"21",X"34",
		X"80",X"34",X"21",X"30",X"80",X"CB",X"66",X"20",X"06",X"FE",X"0F",X"20",X"40",X"CB",X"E6",X"C6",
		X"02",X"E6",X"0F",X"FE",X"05",X"30",X"36",X"3A",X"23",X"80",X"E6",X"04",X"28",X"2F",X"47",X"3A",
		X"32",X"80",X"E6",X"04",X"B8",X"28",X"26",X"21",X"32",X"80",X"CB",X"BE",X"CB",X"B6",X"21",X"16",
		X"80",X"CB",X"8E",X"AF",X"32",X"34",X"80",X"32",X"37",X"80",X"32",X"2D",X"80",X"21",X"23",X"80",
		X"CB",X"EE",X"3E",X"20",X"32",X"39",X"80",X"21",X"30",X"80",X"CB",X"A6",X"C9",X"21",X"23",X"80",
		X"CB",X"56",X"20",X"07",X"21",X"32",X"80",X"CB",X"96",X"18",X"05",X"21",X"32",X"80",X"CB",X"D6",
		X"3A",X"37",X"80",X"11",X"D2",X"39",X"CD",X"51",X"39",X"C9",X"3A",X"1D",X"80",X"C6",X"68",X"21",
		X"00",X"B0",X"CB",X"66",X"20",X"07",X"21",X"16",X"80",X"CB",X"76",X"20",X"0E",X"ED",X"44",X"32",
		X"DF",X"98",X"3A",X"1F",X"80",X"D6",X"20",X"32",X"DE",X"98",X"C9",X"C6",X"90",X"18",X"F0",X"3A",
		X"33",X"80",X"E6",X"01",X"21",X"39",X"80",X"20",X"27",X"7E",X"FE",X"20",X"38",X"05",X"20",X"06",
		X"3E",X"02",X"C9",X"34",X"18",X"1A",X"35",X"18",X"17",X"21",X"39",X"80",X"7E",X"B7",X"20",X"01",
		X"C9",X"35",X"18",X"0C",X"21",X"39",X"80",X"7E",X"FE",X"40",X"20",X"03",X"3E",X"04",X"C9",X"34",
		X"3E",X"07",X"86",X"4F",X"3E",X"01",X"FE",X"10",X"28",X"05",X"07",X"CB",X"19",X"18",X"F7",X"79",
		X"C9",X"21",X"2D",X"80",X"BE",X"C8",X"77",X"26",X"00",X"6F",X"29",X"29",X"19",X"5E",X"23",X"56",
		X"23",X"7E",X"21",X"00",X"B0",X"CB",X"66",X"20",X"09",X"21",X"16",X"80",X"CB",X"76",X"28",X"02",
		X"EE",X"10",X"EB",X"32",X"DD",X"98",X"C3",X"00",X"51",X"01",X"04",X"04",X"CD",X"DB",X"04",X"C9",
		X"21",X"23",X"80",X"CB",X"56",X"C8",X"26",X"00",X"6F",X"29",X"19",X"5E",X"23",X"56",X"EB",X"3A",
		X"3B",X"80",X"E6",X"03",X"20",X"19",X"3A",X"3B",X"80",X"CB",X"5F",X"20",X"09",X"11",X"3C",X"00",
		X"19",X"3E",X"10",X"32",X"3B",X"80",X"11",X"A5",X"88",X"01",X"06",X"02",X"CD",X"DB",X"04",X"21",
		X"3B",X"80",X"35",X"C9",X"9E",X"3A",X"AA",X"3A",X"B6",X"3A",X"C2",X"3A",X"CE",X"3A",X"3E",X"3A",
		X"00",X"00",X"4E",X"3A",X"00",X"00",X"5E",X"3A",X"00",X"00",X"4E",X"3A",X"10",X"00",X"3E",X"3A",
		X"10",X"00",X"5E",X"3A",X"00",X"00",X"4E",X"3A",X"10",X"00",X"3E",X"3A",X"10",X"00",X"2E",X"3A",
		X"10",X"00",X"1E",X"3A",X"10",X"00",X"2E",X"3A",X"30",X"00",X"3E",X"3A",X"30",X"00",X"4E",X"3A",
		X"30",X"00",X"5E",X"3A",X"20",X"00",X"4E",X"3A",X"20",X"00",X"3E",X"3A",X"20",X"00",X"2E",X"3A",
		X"20",X"00",X"1E",X"3A",X"00",X"00",X"2E",X"3A",X"00",X"00",X"3E",X"3A",X"00",X"00",X"4E",X"3A",
		X"00",X"00",X"6E",X"3A",X"00",X"00",X"7E",X"3A",X"00",X"00",X"8E",X"3A",X"00",X"00",X"00",X"01",
		X"02",X"03",X"04",X"05",X"06",X"07",X"08",X"09",X"0A",X"0B",X"0C",X"0D",X"0E",X"0F",X"10",X"11",
		X"12",X"13",X"14",X"15",X"16",X"17",X"18",X"19",X"1A",X"1B",X"1C",X"1D",X"1E",X"1F",X"20",X"21",
		X"22",X"23",X"24",X"25",X"26",X"27",X"28",X"29",X"2A",X"2B",X"2C",X"2D",X"2E",X"2F",X"30",X"31",
		X"32",X"33",X"34",X"35",X"36",X"37",X"38",X"39",X"3A",X"3B",X"3C",X"3D",X"3E",X"3F",X"40",X"41",
		X"42",X"43",X"44",X"45",X"46",X"47",X"48",X"49",X"4A",X"4B",X"4C",X"4D",X"4E",X"4F",X"50",X"51",
		X"52",X"53",X"54",X"55",X"56",X"57",X"58",X"59",X"5A",X"5B",X"5C",X"5D",X"5E",X"5F",X"60",X"61",
		X"62",X"63",X"64",X"65",X"66",X"67",X"68",X"69",X"6A",X"6B",X"6C",X"6D",X"6E",X"6F",X"70",X"71",
		X"72",X"73",X"74",X"75",X"76",X"77",X"78",X"79",X"7A",X"7B",X"7C",X"7D",X"7E",X"7F",X"80",X"81",
		X"82",X"83",X"84",X"85",X"86",X"87",X"88",X"89",X"8A",X"8B",X"8C",X"8D",X"8E",X"8F",X"90",X"91",
		X"92",X"93",X"94",X"95",X"96",X"97",X"98",X"99",X"9A",X"9B",X"9C",X"9D",X"9E",X"9F",X"A0",X"A1",
		X"A2",X"A3",X"A4",X"A5",X"A6",X"A7",X"A8",X"A9",X"AA",X"AB",X"AC",X"AD",X"AE",X"AF",X"B0",X"B1",
		X"B2",X"B3",X"B4",X"B5",X"B6",X"B7",X"B8",X"B9",X"BA",X"BB",X"BC",X"BD",X"BE",X"BF",X"C0",X"C1",
		X"C2",X"C3",X"C4",X"C5",X"C6",X"C7",X"C8",X"C9",X"CA",X"CB",X"CC",X"CD",X"CE",X"CF",X"D0",X"D1",
		X"D2",X"D3",X"D4",X"D5",X"D6",X"D7",X"D8",X"D9",X"DA",X"DB",X"DC",X"DD",X"DE",X"DF",X"E0",X"E1",
		X"E2",X"E3",X"E4",X"E5",X"E6",X"E7",X"E8",X"E9",X"EA",X"EB",X"EC",X"ED",X"EE",X"EF",X"F0",X"F1",
		X"F2",X"F3",X"F4",X"F5",X"F6",X"F7",X"3A",X"2D",X"80",X"B7",X"20",X"4C",X"21",X"1D",X"80",X"46",
		X"21",X"1F",X"80",X"6E",X"3E",X"08",X"80",X"67",X"3E",X"10",X"85",X"6F",X"01",X"06",X"06",X"CD",
		X"D9",X"41",X"DA",X"5A",X"3C",X"21",X"1D",X"80",X"46",X"21",X"1F",X"80",X"6E",X"3E",X"0E",X"80",
		X"67",X"3E",X"0F",X"85",X"6F",X"01",X"06",X"05",X"CD",X"D9",X"41",X"DA",X"5A",X"3C",X"21",X"1D",
		X"80",X"66",X"3A",X"1F",X"80",X"6F",X"3E",X"10",X"84",X"67",X"3E",X"08",X"85",X"6F",X"01",X"09",
		X"07",X"CD",X"D9",X"41",X"DA",X"5A",X"3C",X"C9",X"FE",X"01",X"20",X"46",X"21",X"1D",X"80",X"66",
		X"3A",X"1F",X"80",X"C6",X"10",X"6F",X"3E",X"09",X"84",X"67",X"01",X"07",X"08",X"CD",X"D9",X"41",
		X"DA",X"5A",X"3C",X"21",X"1D",X"80",X"66",X"3A",X"1F",X"80",X"C6",X"0E",X"6F",X"3E",X"0B",X"84",
		X"67",X"01",X"09",X"07",X"CD",X"D9",X"41",X"DA",X"5A",X"3C",X"21",X"1D",X"80",X"66",X"3A",X"1F",
		X"80",X"C6",X"04",X"6F",X"3E",X"0E",X"84",X"67",X"01",X"0A",X"09",X"CD",X"D9",X"41",X"DA",X"5A",
		X"3C",X"C9",X"FE",X"02",X"20",X"28",X"3A",X"1D",X"80",X"C6",X"0B",X"67",X"3A",X"1F",X"80",X"6F",
		X"01",X"0A",X"16",X"CD",X"D9",X"41",X"DA",X"5A",X"3C",X"3A",X"1D",X"80",X"C6",X"0D",X"67",X"3A",
		X"1F",X"80",X"C6",X"16",X"6F",X"01",X"06",X"08",X"CD",X"D9",X"41",X"38",X"7D",X"C9",X"FE",X"03",
		X"20",X"3D",X"3A",X"1D",X"80",X"C6",X"08",X"67",X"3A",X"1F",X"80",X"C6",X"04",X"6F",X"01",X"0A",
		X"09",X"CD",X"D9",X"41",X"38",X"64",X"3A",X"1D",X"80",X"C6",X"0C",X"67",X"3A",X"1F",X"80",X"C6",
		X"0E",X"6F",X"01",X"09",X"07",X"CD",X"D9",X"41",X"38",X"50",X"3A",X"1D",X"80",X"C6",X"11",X"67",
		X"3A",X"1F",X"80",X"C6",X"15",X"6F",X"01",X"06",X"08",X"CD",X"D9",X"41",X"38",X"3C",X"C9",X"3A",
		X"1D",X"80",X"C6",X"06",X"67",X"3A",X"1F",X"80",X"C6",X"08",X"6F",X"01",X"0B",X"07",X"CD",X"D9",
		X"41",X"38",X"27",X"3A",X"1D",X"80",X"C6",X"0B",X"67",X"3A",X"1F",X"80",X"C6",X"0F",X"6F",X"01",
		X"07",X"04",X"CD",X"D9",X"41",X"38",X"13",X"3A",X"1D",X"80",X"C6",X"12",X"67",X"3A",X"1F",X"80",
		X"C6",X"10",X"6F",X"01",X"06",X"07",X"CD",X"D9",X"41",X"D0",X"21",X"16",X"80",X"CB",X"DE",X"C9",
		X"1A",X"B7",X"C8",X"21",X"33",X"80",X"CB",X"6F",X"20",X"1A",X"E6",X"0F",X"A6",X"3E",X"00",X"C0",
		X"1A",X"FE",X"C3",X"20",X"15",X"21",X"23",X"80",X"7E",X"E6",X"03",X"C8",X"3E",X"01",X"CB",X"4E",
		X"C0",X"3E",X"FF",X"C9",X"E6",X"0F",X"A6",X"3E",X"00",X"C8",X"1A",X"CB",X"7F",X"3E",X"01",X"C0",
		X"3E",X"FF",X"C9",X"40",X"00",X"38",X"0F",X"30",X"1E",X"20",X"2D",X"00",X"3C",X"38",X"00",X"30",
		X"0F",X"20",X"1E",X"19",X"2D",X"18",X"3C",X"81",X"00",X"41",X"A3",X"00",X"43",X"80",X"00",X"00",
		X"A3",X"00",X"83",X"81",X"00",X"81",X"81",X"83",X"41",X"A3",X"83",X"43",X"80",X"83",X"00",X"A3",
		X"83",X"83",X"81",X"83",X"81",X"83",X"83",X"41",X"81",X"83",X"43",X"81",X"83",X"00",X"81",X"83",
		X"83",X"83",X"83",X"81",X"87",X"83",X"43",X"83",X"83",X"47",X"83",X"83",X"00",X"83",X"83",X"87",
		X"87",X"83",X"83",X"00",X"83",X"47",X"00",X"83",X"4F",X"00",X"83",X"00",X"00",X"83",X"8F",X"00",
		X"83",X"87",X"83",X"47",X"47",X"81",X"47",X"4F",X"81",X"47",X"C3",X"81",X"47",X"8F",X"83",X"47",
		X"87",X"87",X"43",X"43",X"83",X"43",X"47",X"83",X"43",X"C3",X"83",X"43",X"87",X"87",X"43",X"8F",
		X"00",X"43",X"43",X"00",X"43",X"47",X"00",X"43",X"C3",X"00",X"43",X"87",X"00",X"43",X"83",X"00",
		X"43",X"47",X"00",X"43",X"4F",X"00",X"43",X"00",X"00",X"43",X"8F",X"00",X"43",X"87",X"43",X"00",
		X"00",X"43",X"00",X"00",X"43",X"00",X"00",X"43",X"00",X"00",X"43",X"00",X"00",X"21",X"39",X"80",
		X"CB",X"66",X"20",X"46",X"CB",X"7E",X"20",X"07",X"CB",X"FE",X"3A",X"2F",X"80",X"EF",X"C9",X"CB",
		X"E6",X"21",X"1D",X"06",X"22",X"34",X"80",X"2A",X"30",X"80",X"22",X"32",X"80",X"7C",X"B7",X"20",
		X"05",X"21",X"39",X"80",X"CB",X"DE",X"AF",X"11",X"AB",X"3E",X"CD",X"15",X"42",X"21",X"01",X"06",
		X"CD",X"54",X"01",X"DA",X"33",X"3E",X"2A",X"32",X"80",X"ED",X"4B",X"34",X"80",X"11",X"72",X"3E",
		X"CD",X"92",X"01",X"3A",X"21",X"80",X"32",X"37",X"80",X"C9",X"21",X"39",X"80",X"CB",X"56",X"C2",
		X"12",X"3E",X"3A",X"32",X"80",X"D6",X"D0",X"30",X"05",X"21",X"39",X"80",X"CB",X"CE",X"2A",X"32",
		X"80",X"11",X"03",X"03",X"19",X"01",X"0A",X"0A",X"CD",X"D0",X"3E",X"30",X"07",X"21",X"16",X"80",
		X"CB",X"DE",X"18",X"7F",X"21",X"38",X"80",X"34",X"7E",X"E6",X"03",X"20",X"7F",X"3E",X"01",X"11",
		X"AB",X"3E",X"CD",X"15",X"42",X"B7",X"C8",X"4F",X"CB",X"41",X"28",X"10",X"CD",X"74",X"3E",X"21",
		X"39",X"80",X"CB",X"4E",X"28",X"06",X"B7",X"28",X"5A",X"3C",X"28",X"57",X"CB",X"49",X"28",X"19",
		X"CD",X"91",X"3E",X"2A",X"32",X"80",X"11",X"03",X"03",X"19",X"01",X"0A",X"0A",X"CD",X"D9",X"41",
		X"38",X"07",X"21",X"39",X"80",X"CB",X"D6",X"18",X"19",X"CB",X"51",X"CA",X"6D",X"3D",X"CD",X"9F",
		X"3E",X"21",X"39",X"80",X"CB",X"4E",X"CA",X"6D",X"3D",X"B7",X"28",X"27",X"3C",X"28",X"24",X"C3",
		X"6D",X"3D",X"21",X"36",X"80",X"34",X"46",X"3E",X"10",X"B8",X"38",X"17",X"78",X"E6",X"03",X"28",
		X"08",X"3E",X"0A",X"32",X"35",X"80",X"C3",X"6D",X"3D",X"3E",X"0A",X"CB",X"F7",X"32",X"35",X"80",
		X"C3",X"6D",X"3D",X"AF",X"32",X"39",X"80",X"3A",X"2F",X"80",X"D7",X"C9",X"21",X"3A",X"80",X"34",
		X"7E",X"E6",X"0C",X"20",X"08",X"3E",X"06",X"32",X"35",X"80",X"C3",X"6D",X"3D",X"FE",X"04",X"20",
		X"08",X"3E",X"07",X"32",X"35",X"80",X"C3",X"6D",X"3D",X"FE",X"08",X"20",X"08",X"3E",X"08",X"32",
		X"35",X"80",X"C3",X"6D",X"3D",X"FE",X"0C",X"C2",X"6D",X"3D",X"3E",X"09",X"32",X"35",X"80",X"C3",
		X"6D",X"3D",X"00",X"00",X"3A",X"21",X"80",X"47",X"3A",X"37",X"80",X"21",X"32",X"80",X"90",X"78",
		X"32",X"37",X"80",X"38",X"03",X"35",X"18",X"01",X"34",X"46",X"3A",X"30",X"80",X"ED",X"44",X"80",
		X"C9",X"21",X"33",X"80",X"3A",X"39",X"80",X"CB",X"5F",X"28",X"02",X"34",X"C9",X"35",X"C9",X"21",
		X"32",X"80",X"35",X"46",X"3A",X"30",X"80",X"ED",X"44",X"80",X"C9",X"B3",X"3E",X"C3",X"3E",X"B3",
		X"3E",X"C3",X"3E",X"F4",X"F5",X"F4",X"F5",X"F6",X"F6",X"F7",X"F7",X"F7",X"F7",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"F4",X"F4",X"F7",X"F4",X"F5",X"F4",X"F5",X"F6",X"F7",X"FF",X"FF",X"FF",X"FF",
		X"3A",X"2D",X"80",X"FE",X"05",X"38",X"02",X"3E",X"02",X"57",X"87",X"87",X"82",X"87",X"5F",X"16",
		X"00",X"FD",X"21",X"36",X"3F",X"FD",X"19",X"3A",X"1D",X"80",X"FD",X"86",X"00",X"57",X"3A",X"1F",
		X"80",X"FD",X"86",X"01",X"95",X"30",X"0B",X"ED",X"44",X"FD",X"BE",X"02",X"30",X"20",X"1E",X"01",
		X"18",X"05",X"B8",X"30",X"19",X"1E",X"01",X"7A",X"94",X"30",X"09",X"ED",X"44",X"FD",X"BE",X"03",
		X"30",X"0C",X"18",X"03",X"B9",X"30",X"07",X"3E",X"01",X"A3",X"28",X"02",X"37",X"C9",X"FD",X"7E",
		X"04",X"B7",X"C8",X"3A",X"2D",X"80",X"FE",X"05",X"38",X"02",X"3E",X"02",X"57",X"87",X"87",X"82",
		X"87",X"C6",X"05",X"5F",X"18",X"A9",X"06",X"0E",X"0B",X"0A",X"01",X"0E",X"06",X"0A",X"0B",X"00",
		X"08",X"0A",X"10",X"07",X"01",X"0D",X"02",X"11",X"08",X"00",X"08",X"02",X"14",X"0C",X"01",X"0B",
		X"16",X"07",X"06",X"00",X"05",X"02",X"11",X"08",X"01",X"0D",X"0A",X"10",X"07",X"00",X"03",X"06",
		X"0A",X"0B",X"01",X"0C",X"0E",X"0B",X"0A",X"00",X"3A",X"00",X"B8",X"21",X"32",X"80",X"CB",X"66",
		X"C2",X"B1",X"3F",X"CB",X"E6",X"3A",X"14",X"80",X"CB",X"7F",X"20",X"31",X"21",X"14",X"80",X"CB",
		X"4E",X"20",X"2A",X"CB",X"CE",X"11",X"BA",X"90",X"AF",X"01",X"06",X"00",X"CD",X"06",X"05",X"3A",
		X"16",X"80",X"CB",X"7F",X"20",X"0D",X"11",X"3A",X"91",X"3E",X"24",X"01",X"06",X"00",X"CD",X"06",
		X"05",X"18",X"0A",X"11",X"3A",X"91",X"AF",X"01",X"06",X"00",X"CD",X"06",X"05",X"3E",X"0F",X"EF",
		X"C9",X"3A",X"14",X"80",X"CB",X"7F",X"20",X"F5",X"21",X"32",X"80",X"CB",X"46",X"C2",X"A0",X"40",
		X"2A",X"30",X"80",X"7C",X"B5",X"CA",X"7B",X"40",X"3A",X"16",X"80",X"CB",X"77",X"20",X"0E",X"11",
		X"BE",X"90",X"CD",X"36",X"41",X"21",X"BA",X"90",X"3A",X"2B",X"80",X"18",X"0C",X"11",X"3E",X"91",
		X"CD",X"36",X"41",X"21",X"3A",X"91",X"3A",X"2C",X"80",X"F5",X"E5",X"CD",X"60",X"41",X"E1",X"F1",
		X"B7",X"20",X"21",X"E5",X"11",X"BA",X"92",X"CD",X"28",X"05",X"E1",X"D2",X"71",X"40",X"11",X"BA",
		X"92",X"CD",X"05",X"41",X"0E",X"04",X"3E",X"24",X"11",X"9B",X"92",X"CD",X"06",X"05",X"CD",X"21",
		X"41",X"C3",X"71",X"40",X"FE",X"01",X"20",X"28",X"E5",X"11",X"BA",X"92",X"CD",X"05",X"41",X"E1",
		X"11",X"3A",X"92",X"CD",X"28",X"05",X"D2",X"71",X"40",X"21",X"3A",X"92",X"11",X"BA",X"92",X"CD",
		X"10",X"41",X"21",X"1B",X"92",X"11",X"9B",X"92",X"CD",X"14",X"41",X"CD",X"21",X"41",X"18",X"31",
		X"FE",X"02",X"20",X"27",X"E5",X"11",X"3A",X"92",X"CD",X"05",X"41",X"E1",X"11",X"BA",X"91",X"CD",
		X"28",X"05",X"30",X"1D",X"21",X"BA",X"91",X"11",X"3A",X"92",X"CD",X"10",X"41",X"21",X"9B",X"91",
		X"11",X"1B",X"92",X"CD",X"14",X"41",X"CD",X"21",X"41",X"18",X"06",X"11",X"BA",X"91",X"CD",X"05",
		X"41",X"21",X"32",X"80",X"CB",X"46",X"C0",X"3E",X"0F",X"EF",X"C9",X"C3",X"2C",X"52",X"00",X"00",
		X"3E",X"23",X"CD",X"12",X"0D",X"3E",X"24",X"01",X"0F",X"00",X"11",X"48",X"91",X"CD",X"06",X"05",
		X"3E",X"24",X"01",X"13",X"00",X"11",X"86",X"91",X"CD",X"06",X"05",X"21",X"32",X"80",X"CB",X"C6",
		X"2A",X"1B",X"80",X"EB",X"21",X"32",X"80",X"CB",X"76",X"20",X"06",X"CB",X"F6",X"ED",X"53",X"35",
		X"80",X"7B",X"B2",X"20",X"22",X"11",X"80",X"00",X"B7",X"2A",X"35",X"80",X"ED",X"52",X"30",X"05",
		X"21",X"18",X"01",X"18",X"03",X"21",X"50",X"00",X"F7",X"21",X"14",X"80",X"CB",X"EE",X"21",X"16",
		X"80",X"CB",X"86",X"3E",X"0F",X"D7",X"C9",X"3E",X"0E",X"21",X"03",X"00",X"E7",X"21",X"34",X"80",
		X"7E",X"34",X"E6",X"01",X"C0",X"21",X"17",X"80",X"3A",X"16",X"80",X"CB",X"77",X"28",X"01",X"23",
		X"7E",X"FE",X"0A",X"38",X"02",X"3E",X"0A",X"21",X"56",X"41",X"3D",X"5F",X"16",X"00",X"19",X"6E",
		X"26",X"00",X"C3",X"C8",X"3F",X"01",X"05",X"00",X"18",X"03",X"01",X"04",X"00",X"ED",X"B0",X"C9",
		X"06",X"05",X"18",X"02",X"06",X"04",X"4E",X"1A",X"77",X"EB",X"71",X"EB",X"23",X"13",X"10",X"F6",
		X"C9",X"3A",X"16",X"80",X"21",X"2B",X"80",X"11",X"2C",X"80",X"CB",X"77",X"28",X"01",X"EB",X"34",
		X"1A",X"BE",X"C0",X"EB",X"35",X"C9",X"01",X"00",X"05",X"EB",X"3E",X"0F",X"A3",X"81",X"0E",X"00",
		X"86",X"77",X"C6",X"F6",X"30",X"02",X"77",X"0C",X"2B",X"3E",X"04",X"B7",X"CB",X"1A",X"CB",X"1B",
		X"3D",X"20",X"F8",X"10",X"E5",X"C9",X"01",X"01",X"02",X"02",X"03",X"04",X"05",X"07",X"07",X"10",
		X"EB",X"01",X"2E",X"80",X"0A",X"21",X"16",X"80",X"CB",X"76",X"20",X"09",X"CB",X"7F",X"C0",X"CB",
		X"77",X"28",X"09",X"18",X"18",X"CB",X"6F",X"C0",X"CB",X"67",X"20",X"11",X"21",X"CF",X"41",X"EB",
		X"01",X"00",X"B0",X"0A",X"CB",X"5F",X"28",X"09",X"11",X"D4",X"41",X"18",X"04",X"21",X"CA",X"41",
		X"EB",X"CD",X"28",X"05",X"D0",X"01",X"0A",X"01",X"CD",X"75",X"48",X"21",X"19",X"80",X"3A",X"16",
		X"80",X"CB",X"77",X"20",X"11",X"34",X"CD",X"DC",X"0C",X"21",X"2E",X"80",X"CB",X"76",X"20",X"03",
		X"CB",X"F6",X"C9",X"CB",X"FE",X"C9",X"21",X"1A",X"80",X"34",X"CD",X"DC",X"0C",X"21",X"2E",X"80",
		X"CB",X"66",X"20",X"03",X"CB",X"E6",X"C9",X"CB",X"EE",X"C9",X"01",X"00",X"00",X"00",X"00",X"00",
		X"02",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"7C",X"E6",X"07",X"81",X"C6",X"07",X"E6",
		X"F8",X"0F",X"0F",X"0F",X"4F",X"7D",X"80",X"47",X"E5",X"C5",X"CD",X"F8",X"41",X"C1",X"E1",X"D8",
		X"7D",X"C6",X"08",X"6F",X"B8",X"38",X"F1",X"C9",X"3A",X"21",X"80",X"85",X"6F",X"CD",X"46",X"46",
		X"1A",X"FE",X"35",X"28",X"0B",X"FE",X"86",X"30",X"07",X"FE",X"5C",X"D8",X"FE",X"9C",X"3F",X"D8",
		X"13",X"0D",X"20",X"EC",X"C9",X"B7",X"20",X"0E",X"ED",X"5F",X"E6",X"03",X"11",X"3C",X"80",X"12",
		X"AF",X"13",X"12",X"13",X"12",X"C9",X"42",X"4B",X"2A",X"3C",X"80",X"26",X"00",X"29",X"19",X"5E",
		X"23",X"56",X"EB",X"ED",X"5B",X"3D",X"80",X"16",X"00",X"19",X"3A",X"3E",X"80",X"B7",X"28",X"08",
		X"3D",X"32",X"3E",X"80",X"7E",X"E6",X"0F",X"C9",X"7E",X"FE",X"FF",X"28",X"12",X"E6",X"F0",X"0F",
		X"0F",X"0F",X"0F",X"32",X"3E",X"80",X"23",X"11",X"3D",X"80",X"1A",X"3C",X"12",X"18",X"C7",X"21",
		X"3D",X"80",X"36",X"00",X"23",X"36",X"00",X"50",X"59",X"18",X"BB",X"3A",X"00",X"B8",X"21",X"16",
		X"80",X"CB",X"5E",X"C0",X"21",X"32",X"80",X"CB",X"46",X"20",X"30",X"CB",X"C6",X"21",X"37",X"80",
		X"3A",X"2F",X"80",X"E6",X"1F",X"FE",X"09",X"28",X"16",X"3E",X"04",X"32",X"36",X"80",X"36",X"0F",
		X"ED",X"5F",X"CB",X"47",X"28",X"10",X"3E",X"05",X"32",X"36",X"80",X"36",X"13",X"18",X"07",X"3E",
		X"03",X"32",X"36",X"80",X"36",X"0B",X"3A",X"2F",X"80",X"EF",X"C9",X"CB",X"4E",X"20",X"26",X"CB",
		X"CE",X"AF",X"32",X"33",X"80",X"3A",X"21",X"80",X"32",X"38",X"80",X"21",X"02",X"07",X"CD",X"54",
		X"01",X"DA",X"5C",X"43",X"11",X"61",X"43",X"2A",X"30",X"80",X"22",X"34",X"80",X"ED",X"4B",X"36",
		X"80",X"CD",X"92",X"01",X"C9",X"21",X"33",X"80",X"34",X"7E",X"21",X"32",X"80",X"CB",X"9E",X"E6",
		X"07",X"20",X"02",X"CB",X"DE",X"21",X"02",X"07",X"CD",X"54",X"01",X"DA",X"5C",X"43",X"2A",X"34",
		X"80",X"CD",X"70",X"43",X"11",X"61",X"43",X"ED",X"4B",X"36",X"80",X"3A",X"39",X"80",X"B7",X"28",
		X"11",X"11",X"65",X"43",X"3A",X"39",X"80",X"04",X"04",X"FE",X"01",X"28",X"05",X"CB",X"F0",X"11",
		X"69",X"43",X"2A",X"34",X"80",X"CD",X"92",X"01",X"3A",X"33",X"80",X"E6",X"03",X"20",X"33",X"2A",
		X"34",X"80",X"11",X"04",X"04",X"19",X"01",X"08",X"0C",X"CD",X"D0",X"3E",X"38",X"1E",X"21",X"6D",
		X"43",X"3A",X"39",X"80",X"5F",X"16",X"00",X"19",X"7E",X"2A",X"34",X"80",X"84",X"C6",X"04",X"67",
		X"7D",X"C6",X"10",X"6F",X"01",X"08",X"0C",X"CD",X"D0",X"3E",X"30",X"06",X"21",X"16",X"80",X"CB",
		X"DE",X"C9",X"3A",X"34",X"80",X"C6",X"1E",X"B7",X"28",X"02",X"3D",X"C0",X"3A",X"2F",X"80",X"D7",
		X"C9",X"00",X"00",X"00",X"10",X"00",X"00",X"04",X"10",X"00",X"00",X"FC",X"10",X"00",X"04",X"FC",
		X"21",X"38",X"80",X"46",X"3A",X"21",X"80",X"77",X"4F",X"78",X"91",X"21",X"34",X"80",X"86",X"77",
		X"3A",X"32",X"80",X"CB",X"5F",X"C8",X"CB",X"57",X"20",X"06",X"21",X"34",X"80",X"35",X"18",X"5C",
		X"3A",X"35",X"80",X"C6",X"08",X"47",X"3A",X"28",X"80",X"C6",X"08",X"4F",X"3A",X"29",X"80",X"91",
		X"E6",X"FE",X"0F",X"21",X"32",X"80",X"CB",X"E6",X"81",X"B8",X"28",X"4E",X"CB",X"A6",X"3A",X"3A",
		X"80",X"B8",X"28",X"46",X"01",X"08",X"10",X"3A",X"39",X"80",X"FE",X"01",X"20",X"17",X"2A",X"34",
		X"80",X"11",X"00",X"F8",X"19",X"CD",X"D9",X"41",X"30",X"06",X"3E",X"02",X"32",X"39",X"80",X"C9",
		X"21",X"35",X"80",X"35",X"C9",X"2A",X"34",X"80",X"11",X"00",X"10",X"19",X"CD",X"D9",X"41",X"30",
		X"06",X"3E",X"01",X"32",X"39",X"80",X"C9",X"21",X"35",X"80",X"34",X"C9",X"21",X"3B",X"80",X"34",
		X"7E",X"E6",X"1F",X"28",X"05",X"3A",X"39",X"80",X"18",X"09",X"ED",X"5F",X"E6",X"03",X"FE",X"03",
		X"20",X"01",X"AF",X"06",X"03",X"32",X"39",X"80",X"4F",X"87",X"87",X"81",X"5F",X"16",X"00",X"21",
		X"BE",X"44",X"19",X"C5",X"E5",X"46",X"23",X"4E",X"23",X"7E",X"23",X"66",X"6F",X"3A",X"34",X"80",
		X"85",X"6F",X"3A",X"35",X"80",X"84",X"67",X"CD",X"D9",X"41",X"D1",X"C1",X"30",X"70",X"3A",X"39",
		X"80",X"3C",X"FE",X"03",X"20",X"01",X"AF",X"32",X"39",X"80",X"10",X"CC",X"21",X"32",X"80",X"CB",
		X"D6",X"CB",X"66",X"20",X"49",X"3A",X"28",X"80",X"C6",X"08",X"47",X"3A",X"29",X"80",X"90",X"E6",
		X"FC",X"0F",X"0F",X"4F",X"80",X"57",X"3A",X"35",X"80",X"C6",X"08",X"5F",X"92",X"28",X"10",X"38",
		X"0E",X"79",X"87",X"81",X"47",X"7B",X"90",X"30",X"14",X"ED",X"5F",X"CB",X"5F",X"20",X"0E",X"79",
		X"87",X"81",X"32",X"3A",X"80",X"21",X"35",X"80",X"34",X"3E",X"02",X"18",X"0A",X"79",X"32",X"3A",
		X"80",X"21",X"35",X"80",X"35",X"3E",X"01",X"32",X"39",X"80",X"32",X"3C",X"80",X"C9",X"3A",X"3C",
		X"80",X"32",X"39",X"80",X"21",X"35",X"80",X"FE",X"01",X"20",X"01",X"35",X"34",X"C9",X"21",X"32",
		X"80",X"CB",X"96",X"CB",X"A6",X"3E",X"04",X"83",X"5F",X"3E",X"00",X"8A",X"57",X"1A",X"32",X"39",
		X"80",X"B7",X"C8",X"21",X"35",X"80",X"FE",X"01",X"20",X"02",X"35",X"C9",X"34",X"C9",X"18",X"10",
		X"F0",X"00",X"00",X"18",X"08",X"F0",X"F8",X"01",X"18",X"08",X"F0",X"10",X"02",X"3A",X"00",X"B8",
		X"21",X"16",X"80",X"CB",X"5E",X"C0",X"21",X"32",X"80",X"CB",X"46",X"20",X"07",X"CB",X"C6",X"3A",
		X"2F",X"80",X"EF",X"C9",X"CB",X"4E",X"20",X"2A",X"CB",X"CE",X"AF",X"32",X"33",X"80",X"21",X"01",
		X"05",X"CD",X"54",X"01",X"DA",X"F3",X"45",X"06",X"03",X"0E",X"1C",X"ED",X"43",X"36",X"80",X"3A",
		X"21",X"80",X"32",X"38",X"80",X"2A",X"30",X"80",X"22",X"34",X"80",X"11",X"6C",X"46",X"CD",X"92",
		X"01",X"C9",X"CB",X"6E",X"C2",X"09",X"46",X"CB",X"76",X"C2",X"13",X"46",X"21",X"33",X"80",X"34",
		X"7E",X"21",X"32",X"80",X"CB",X"9E",X"E6",X"07",X"20",X"02",X"CB",X"DE",X"21",X"01",X"05",X"CD",
		X"54",X"01",X"DA",X"F3",X"45",X"CD",X"70",X"43",X"CD",X"33",X"46",X"11",X"6C",X"46",X"2A",X"34",
		X"80",X"ED",X"4B",X"36",X"80",X"CD",X"92",X"01",X"3A",X"33",X"80",X"E6",X"03",X"C2",X"E9",X"45",
		X"2A",X"34",X"80",X"11",X"02",X"01",X"19",X"01",X"0C",X"0E",X"CD",X"D0",X"3E",X"D2",X"E9",X"45",
		X"3A",X"2D",X"80",X"FE",X"02",X"20",X"2F",X"3A",X"1F",X"80",X"C6",X"18",X"47",X"3A",X"34",X"80",
		X"90",X"38",X"23",X"3A",X"35",X"80",X"C6",X"08",X"47",X"3A",X"1D",X"80",X"C6",X"0C",X"B8",X"30",
		X"15",X"C6",X"06",X"B8",X"38",X"10",X"01",X"0C",X"01",X"CD",X"75",X"48",X"21",X"32",X"80",X"CB",
		X"F6",X"AF",X"32",X"2A",X"80",X"C9",X"21",X"32",X"80",X"CB",X"EE",X"CD",X"FD",X"01",X"01",X"0B",
		X"01",X"CD",X"75",X"48",X"AF",X"32",X"33",X"80",X"3A",X"2A",X"80",X"3C",X"FE",X"0A",X"30",X"09",
		X"07",X"07",X"07",X"07",X"6F",X"26",X"00",X"18",X"04",X"26",X"01",X"2E",X"00",X"3E",X"0F",X"E7",
		X"3A",X"34",X"80",X"2A",X"21",X"80",X"85",X"6F",X"3A",X"35",X"80",X"67",X"CD",X"46",X"46",X"3E",
		X"86",X"21",X"2A",X"80",X"86",X"3C",X"12",X"13",X"3E",X"86",X"12",X"21",X"2A",X"80",X"7E",X"FE",
		X"09",X"30",X"01",X"34",X"AF",X"32",X"33",X"80",X"C9",X"3A",X"34",X"80",X"C6",X"10",X"B7",X"28",
		X"02",X"3D",X"C0",X"3A",X"32",X"80",X"CB",X"77",X"20",X"06",X"3E",X"0E",X"21",X"20",X"00",X"E7",
		X"AF",X"32",X"2A",X"80",X"3A",X"2F",X"80",X"D7",X"C9",X"21",X"33",X"80",X"34",X"7E",X"FE",X"40",
		X"28",X"F2",X"C9",X"21",X"01",X"05",X"CD",X"54",X"01",X"38",X"D8",X"21",X"35",X"80",X"56",X"2B",
		X"7E",X"3D",X"32",X"34",X"80",X"5F",X"EB",X"0E",X"1C",X"06",X"05",X"11",X"6C",X"46",X"CD",X"92",
		X"01",X"18",X"B6",X"21",X"3D",X"80",X"34",X"7E",X"E6",X"0F",X"C0",X"21",X"37",X"80",X"34",X"7E",
		X"FE",X"05",X"C0",X"36",X"03",X"C9",X"7D",X"C6",X"18",X"ED",X"44",X"E6",X"F8",X"5F",X"16",X"00",
		X"CB",X"13",X"CB",X"12",X"CB",X"13",X"CB",X"12",X"7A",X"E6",X"03",X"57",X"7C",X"C6",X"20",X"E6",
		X"F8",X"0F",X"0F",X"0F",X"B3",X"5F",X"21",X"00",X"90",X"19",X"EB",X"C9",X"00",X"00",X"3A",X"00",
		X"B8",X"21",X"32",X"80",X"CB",X"7E",X"20",X"11",X"CB",X"FE",X"3E",X"13",X"EF",X"21",X"23",X"80",
		X"CB",X"AE",X"2A",X"21",X"80",X"22",X"37",X"80",X"C9",X"CB",X"76",X"20",X"3F",X"CB",X"F6",X"21",
		X"16",X"80",X"CB",X"D6",X"21",X"36",X"80",X"36",X"00",X"2A",X"31",X"80",X"26",X"00",X"22",X"24",
		X"80",X"2A",X"30",X"80",X"26",X"00",X"ED",X"5B",X"37",X"80",X"19",X"22",X"26",X"80",X"22",X"37",
		X"80",X"3A",X"24",X"80",X"67",X"CD",X"46",X"46",X"D5",X"21",X"A8",X"47",X"01",X"04",X"01",X"CD",
		X"C5",X"04",X"D1",X"3E",X"06",X"01",X"04",X"01",X"CD",X"32",X"05",X"C9",X"21",X"34",X"80",X"34",
		X"7E",X"E6",X"03",X"C0",X"CD",X"26",X"47",X"28",X"36",X"21",X"16",X"80",X"CB",X"8E",X"21",X"23",
		X"80",X"CB",X"6E",X"20",X"1B",X"2A",X"26",X"80",X"ED",X"5B",X"21",X"80",X"B7",X"ED",X"52",X"3A",
		X"24",X"80",X"67",X"01",X"20",X"20",X"CD",X"D0",X"3E",X"30",X"05",X"21",X"16",X"80",X"CB",X"CE",
		X"21",X"35",X"80",X"34",X"7E",X"E6",X"01",X"C0",X"23",X"34",X"7E",X"E6",X"03",X"77",X"C9",X"3E",
		X"13",X"D7",X"21",X"16",X"80",X"CB",X"96",X"21",X"23",X"80",X"CB",X"AE",X"21",X"00",X"00",X"22",
		X"24",X"80",X"22",X"26",X"80",X"C9",X"21",X"33",X"80",X"36",X"00",X"21",X"33",X"80",X"7E",X"CB",
		X"BF",X"6F",X"26",X"00",X"29",X"29",X"29",X"ED",X"5B",X"37",X"80",X"19",X"ED",X"5B",X"21",X"80",
		X"EB",X"01",X"10",X"00",X"B7",X"ED",X"42",X"B7",X"ED",X"52",X"30",X"23",X"2A",X"21",X"80",X"01",
		X"E8",X"00",X"09",X"ED",X"52",X"38",X"18",X"CD",X"7D",X"47",X"D5",X"01",X"04",X"01",X"CD",X"C5",
		X"04",X"D1",X"3E",X"06",X"01",X"04",X"01",X"CD",X"32",X"05",X"21",X"33",X"80",X"CB",X"FE",X"21",
		X"33",X"80",X"34",X"7E",X"CB",X"BF",X"FE",X"04",X"20",X"B1",X"CB",X"7E",X"C9",X"6B",X"3A",X"24",
		X"80",X"67",X"CD",X"46",X"46",X"D5",X"3A",X"36",X"80",X"11",X"A0",X"47",X"26",X"00",X"6F",X"29",
		X"19",X"5E",X"23",X"56",X"2A",X"33",X"80",X"CB",X"BD",X"26",X"00",X"29",X"29",X"19",X"D1",X"C9",
		X"A8",X"47",X"B8",X"47",X"C7",X"47",X"D7",X"47",X"5C",X"5D",X"5E",X"5F",X"60",X"61",X"62",X"63",
		X"64",X"65",X"66",X"67",X"68",X"69",X"6A",X"6B",X"6C",X"6D",X"6E",X"6F",X"70",X"71",X"72",X"73",
		X"74",X"75",X"76",X"77",X"78",X"7A",X"7B",X"7C",X"7D",X"7E",X"7F",X"80",X"81",X"82",X"83",X"84",
		X"85",X"86",X"87",X"88",X"89",X"8A",X"8B",X"8C",X"8D",X"8E",X"8F",X"90",X"91",X"92",X"93",X"94",
		X"95",X"96",X"97",X"98",X"99",X"9A",X"9B",X"DD",X"21",X"A1",X"81",X"DD",X"CB",X"00",X"7E",X"C4",
		X"09",X"48",X"DD",X"21",X"A9",X"81",X"DD",X"CB",X"00",X"7E",X"C4",X"09",X"48",X"DD",X"21",X"B1",
		X"81",X"DD",X"CB",X"00",X"7E",X"C4",X"09",X"48",X"C9",X"DD",X"7E",X"02",X"B7",X"28",X"04",X"DD",
		X"35",X"02",X"C9",X"DD",X"7E",X"03",X"DD",X"77",X"02",X"DD",X"7E",X"04",X"B7",X"28",X"04",X"DD",
		X"35",X"04",X"C9",X"DD",X"6E",X"06",X"DD",X"66",X"07",X"06",X"00",X"DD",X"4E",X"05",X"09",X"7E",
		X"FE",X"FF",X"20",X"1B",X"DD",X"CB",X"00",X"6E",X"20",X"0C",X"DD",X"CB",X"00",X"76",X"28",X"06",
		X"DD",X"36",X"05",X"00",X"18",X"DD",X"DD",X"36",X"00",X"00",X"21",X"9F",X"81",X"35",X"C9",X"0F",
		X"0F",X"0F",X"0F",X"E6",X"0F",X"DD",X"77",X"04",X"7E",X"E6",X"0F",X"07",X"01",X"EE",X"49",X"EB",
		X"26",X"00",X"6F",X"09",X"4E",X"23",X"46",X"60",X"69",X"01",X"72",X"48",X"C5",X"13",X"DD",X"34",
		X"05",X"E9",X"38",X"AF",X"C9",X"21",X"14",X"80",X"CB",X"7E",X"C0",X"C5",X"79",X"CD",X"85",X"48",
		X"C1",X"0C",X"10",X"F1",X"C9",X"21",X"A1",X"81",X"11",X"08",X"00",X"06",X"03",X"4F",X"E6",X"7F",
		X"CB",X"79",X"20",X"42",X"3A",X"9F",X"81",X"3C",X"FE",X"04",X"3F",X"D8",X"32",X"9F",X"81",X"AF",
		X"BE",X"28",X"05",X"19",X"10",X"FA",X"37",X"C9",X"E5",X"05",X"70",X"23",X"71",X"EB",X"69",X"67",
		X"47",X"29",X"09",X"01",X"C4",X"49",X"09",X"EB",X"1A",X"CB",X"47",X"28",X"04",X"2B",X"CB",X"F6",
		X"23",X"AF",X"23",X"77",X"23",X"77",X"23",X"77",X"23",X"77",X"23",X"13",X"1A",X"77",X"23",X"13",
		X"1A",X"77",X"E1",X"CB",X"FE",X"C9",X"23",X"4F",X"7E",X"B9",X"28",X"05",X"19",X"10",X"F9",X"37",
		X"C9",X"2B",X"CB",X"EE",X"C9",X"37",X"C9",X"DD",X"7E",X"00",X"E6",X"03",X"07",X"D3",X"08",X"47",
		X"1A",X"D3",X"09",X"04",X"78",X"D3",X"08",X"13",X"1A",X"D3",X"09",X"DD",X"34",X"05",X"DD",X"34",
		X"05",X"37",X"C9",X"DD",X"7E",X"00",X"E6",X"03",X"C6",X"08",X"D3",X"08",X"1A",X"D3",X"09",X"DD",
		X"34",X"05",X"37",X"C9",X"3E",X"0B",X"D3",X"08",X"1A",X"D3",X"09",X"13",X"3E",X"0C",X"D3",X"08",
		X"1A",X"D3",X"09",X"DD",X"34",X"05",X"DD",X"34",X"05",X"37",X"C9",X"3E",X"0D",X"D3",X"08",X"1A",
		X"D3",X"09",X"DD",X"34",X"05",X"37",X"C9",X"3E",X"07",X"D3",X"08",X"DD",X"7E",X"00",X"E6",X"03",
		X"3C",X"47",X"3E",X"80",X"07",X"10",X"FD",X"21",X"A0",X"81",X"B6",X"77",X"D3",X"09",X"B7",X"C9",
		X"1A",X"DD",X"77",X"03",X"DD",X"34",X"05",X"37",X"C9",X"3E",X"07",X"D3",X"08",X"DD",X"7E",X"00",
		X"E6",X"03",X"3C",X"47",X"3E",X"80",X"07",X"10",X"FD",X"21",X"A0",X"81",X"2F",X"A6",X"77",X"D3",
		X"09",X"B7",X"C9",X"1A",X"07",X"21",X"21",X"4E",X"16",X"00",X"5F",X"19",X"EB",X"CD",X"E7",X"48",
		X"DD",X"35",X"05",X"18",X"D4",X"3E",X"07",X"D3",X"08",X"DD",X"7E",X"00",X"E6",X"03",X"3C",X"47",
		X"3E",X"04",X"07",X"10",X"FD",X"21",X"A0",X"81",X"2F",X"A6",X"77",X"D3",X"09",X"B7",X"C9",X"3E",
		X"07",X"D3",X"08",X"DD",X"7E",X"00",X"E6",X"03",X"3C",X"47",X"3E",X"04",X"07",X"10",X"FD",X"21",
		X"A0",X"81",X"B6",X"77",X"D3",X"09",X"B7",X"C9",X"3E",X"06",X"D3",X"08",X"1A",X"D3",X"09",X"DD",
		X"34",X"05",X"37",X"C9",X"00",X"0C",X"4A",X"00",X"6F",X"4A",X"00",X"AD",X"4A",X"00",X"E2",X"4A",
		X"00",X"22",X"4B",X"00",X"61",X"4B",X"01",X"A0",X"4B",X"01",X"89",X"4C",X"00",X"48",X"4D",X"00",
		X"9C",X"4D",X"00",X"BE",X"4D",X"00",X"D8",X"4D",X"00",X"EA",X"4D",X"00",X"10",X"4E",X"E5",X"48",
		X"E7",X"48",X"03",X"49",X"37",X"49",X"50",X"49",X"14",X"49",X"2B",X"49",X"59",X"49",X"73",X"49",
		X"85",X"49",X"9F",X"49",X"B8",X"49",X"E5",X"48",X"E5",X"48",X"E5",X"48",X"04",X"02",X"02",X"0B",
		X"28",X"05",X"03",X"28",X"05",X"03",X"18",X"05",X"18",X"04",X"18",X"05",X"18",X"07",X"28",X"09",
		X"03",X"28",X"09",X"03",X"18",X"09",X"18",X"07",X"18",X"09",X"18",X"0A",X"28",X"0C",X"03",X"28",
		X"0C",X"03",X"18",X"0C",X"18",X"0B",X"18",X"0C",X"18",X"11",X"78",X"0C",X"33",X"00",X"28",X"0C",
		X"03",X"28",X"0E",X"03",X"28",X"0C",X"03",X"28",X"0A",X"03",X"28",X"09",X"03",X"28",X"07",X"03",
		X"28",X"05",X"03",X"28",X"04",X"03",X"28",X"05",X"03",X"28",X"07",X"03",X"08",X"09",X"03",X"08",
		X"0A",X"03",X"28",X"09",X"03",X"28",X"07",X"03",X"78",X"05",X"73",X"00",X"02",X"00",X"FF",X"04",
		X"02",X"02",X"0C",X"68",X"05",X"03",X"68",X"00",X"03",X"68",X"09",X"03",X"68",X"05",X"43",X"28",
		X"00",X"03",X"68",X"05",X"03",X"08",X"05",X"03",X"08",X"05",X"03",X"28",X"04",X"03",X"28",X"02",
		X"03",X"28",X"00",X"03",X"68",X"0A",X"03",X"68",X"07",X"03",X"68",X"04",X"03",X"68",X"00",X"03",
		X"68",X"07",X"03",X"68",X"00",X"03",X"68",X"05",X"03",X"02",X"00",X"73",X"FF",X"04",X"02",X"02",
		X"09",X"33",X"08",X"11",X"63",X"08",X"11",X"63",X"08",X"11",X"63",X"08",X"11",X"63",X"08",X"11",
		X"63",X"08",X"11",X"63",X"08",X"11",X"63",X"08",X"11",X"63",X"08",X"11",X"63",X"08",X"11",X"63",
		X"08",X"11",X"63",X"08",X"11",X"63",X"08",X"11",X"63",X"08",X"11",X"23",X"08",X"11",X"02",X"00",
		X"43",X"FF",X"04",X"02",X"02",X"0C",X"88",X"0C",X"03",X"08",X"0C",X"03",X"08",X"0C",X"03",X"28",
		X"0C",X"03",X"28",X"07",X"03",X"28",X"04",X"03",X"28",X"07",X"03",X"28",X"0C",X"03",X"28",X"07",
		X"03",X"28",X"0C",X"03",X"28",X"10",X"03",X"68",X"0C",X"03",X"48",X"13",X"03",X"08",X"13",X"03",
		X"E8",X"13",X"03",X"A8",X"10",X"03",X"28",X"07",X"03",X"E8",X"0C",X"38",X"0C",X"02",X"00",X"B3",
		X"00",X"FF",X"04",X"02",X"02",X"0C",X"88",X"07",X"03",X"08",X"07",X"03",X"08",X"07",X"03",X"28",
		X"07",X"03",X"28",X"04",X"03",X"28",X"04",X"03",X"28",X"07",X"03",X"28",X"07",X"03",X"28",X"04",
		X"03",X"28",X"07",X"03",X"28",X"0C",X"03",X"68",X"07",X"03",X"48",X"10",X"03",X"08",X"10",X"03",
		X"E8",X"10",X"03",X"A8",X"0C",X"03",X"28",X"07",X"03",X"E8",X"07",X"38",X"07",X"02",X"00",X"B3",
		X"FF",X"04",X"02",X"02",X"0C",X"88",X"04",X"03",X"08",X"04",X"03",X"08",X"04",X"03",X"28",X"04",
		X"03",X"28",X"00",X"03",X"28",X"00",X"03",X"28",X"04",X"03",X"28",X"04",X"03",X"28",X"00",X"03",
		X"28",X"04",X"03",X"28",X"07",X"03",X"68",X"04",X"03",X"48",X"0C",X"03",X"08",X"0C",X"03",X"E8",
		X"0C",X"03",X"A8",X"07",X"03",X"28",X"04",X"03",X"E8",X"00",X"38",X"00",X"02",X"00",X"B3",X"FF",
		X"04",X"05",X"02",X"08",X"08",X"0C",X"08",X"10",X"08",X"13",X"08",X"10",X"08",X"13",X"03",X"08",
		X"18",X"03",X"08",X"17",X"03",X"08",X"15",X"03",X"08",X"13",X"03",X"08",X"11",X"03",X"08",X"10",
		X"08",X"11",X"08",X"13",X"08",X"10",X"08",X"11",X"08",X"0E",X"08",X"10",X"08",X"0C",X"08",X"0B",
		X"08",X"0E",X"08",X"13",X"08",X"17",X"08",X"13",X"08",X"11",X"08",X"10",X"08",X"0E",X"08",X"0C",
		X"08",X"10",X"08",X"13",X"08",X"10",X"08",X"13",X"03",X"08",X"18",X"03",X"08",X"17",X"03",X"08",
		X"15",X"03",X"08",X"13",X"03",X"08",X"11",X"03",X"08",X"10",X"08",X"11",X"08",X"13",X"08",X"10",
		X"08",X"11",X"08",X"0E",X"08",X"10",X"08",X"0C",X"08",X"0E",X"08",X"13",X"08",X"17",X"08",X"13",
		X"28",X"18",X"03",X"08",X"15",X"08",X"17",X"08",X"18",X"08",X"15",X"08",X"17",X"08",X"15",X"08",
		X"13",X"08",X"11",X"08",X"13",X"08",X"15",X"08",X"17",X"08",X"13",X"08",X"15",X"08",X"13",X"08",
		X"11",X"08",X"10",X"08",X"11",X"08",X"13",X"08",X"15",X"08",X"11",X"08",X"13",X"08",X"11",X"08",
		X"10",X"08",X"0E",X"08",X"11",X"08",X"0E",X"08",X"11",X"08",X"15",X"08",X"13",X"08",X"11",X"08",
		X"10",X"08",X"0E",X"08",X"0C",X"08",X"10",X"08",X"13",X"08",X"10",X"08",X"13",X"03",X"08",X"18",
		X"03",X"08",X"17",X"03",X"08",X"15",X"03",X"08",X"13",X"03",X"08",X"11",X"03",X"08",X"10",X"08",
		X"11",X"08",X"13",X"08",X"10",X"08",X"11",X"08",X"0E",X"08",X"10",X"08",X"0C",X"08",X"0B",X"08",
		X"0E",X"08",X"13",X"08",X"17",X"28",X"18",X"03",X"FF",X"04",X"05",X"02",X"08",X"08",X"00",X"03",
		X"08",X"07",X"03",X"08",X"00",X"03",X"08",X"07",X"03",X"08",X"00",X"03",X"08",X"07",X"03",X"08",
		X"00",X"03",X"08",X"07",X"03",X"08",X"02",X"03",X"08",X"05",X"03",X"08",X"02",X"03",X"08",X"05",
		X"03",X"08",X"02",X"03",X"08",X"05",X"03",X"08",X"07",X"03",X"08",X"02",X"03",X"08",X"00",X"03",
		X"08",X"07",X"03",X"08",X"00",X"03",X"08",X"07",X"03",X"08",X"00",X"03",X"08",X"07",X"03",X"08",
		X"00",X"03",X"08",X"07",X"03",X"08",X"05",X"03",X"08",X"02",X"03",X"08",X"05",X"03",X"08",X"02",
		X"03",X"08",X"07",X"03",X"08",X"07",X"03",X"28",X"00",X"03",X"08",X"09",X"03",X"08",X"05",X"03",
		X"08",X"09",X"03",X"08",X"05",X"03",X"08",X"07",X"03",X"08",X"04",X"03",X"08",X"07",X"03",X"08",
		X"04",X"03",X"08",X"09",X"03",X"08",X"05",X"03",X"08",X"09",X"03",X"08",X"05",X"03",X"08",X"07",
		X"03",X"08",X"05",X"03",X"08",X"04",X"03",X"08",X"02",X"03",X"08",X"00",X"03",X"08",X"07",X"03",
		X"08",X"00",X"03",X"08",X"07",X"03",X"08",X"00",X"03",X"08",X"07",X"03",X"08",X"00",X"03",X"08",
		X"07",X"03",X"08",X"05",X"03",X"08",X"02",X"03",X"08",X"05",X"03",X"08",X"02",X"03",X"08",X"07",
		X"03",X"08",X"07",X"03",X"28",X"00",X"03",X"FF",X"04",X"01",X"02",X"0C",X"01",X"8E",X"01",X"27",
		X"01",X"C6",X"00",X"27",X"01",X"9F",X"00",X"27",X"01",X"49",X"00",X"27",X"01",X"4C",X"00",X"27",
		X"01",X"51",X"00",X"27",X"01",X"56",X"00",X"37",X"02",X"0A",X"01",X"5E",X"00",X"37",X"02",X"09",
		X"01",X"68",X"00",X"37",X"02",X"08",X"01",X"79",X"00",X"37",X"01",X"99",X"00",X"37",X"02",X"07",
		X"01",X"F2",X"00",X"37",X"02",X"06",X"01",X"1D",X"01",X"37",X"02",X"05",X"01",X"3C",X"01",X"37",
		X"02",X"03",X"01",X"65",X"01",X"37",X"01",X"9E",X"01",X"37",X"03",X"FF",X"04",X"05",X"02",X"0C",
		X"07",X"61",X"63",X"00",X"61",X"6B",X"00",X"61",X"75",X"00",X"61",X"7F",X"00",X"61",X"8E",X"00",
		X"61",X"7F",X"00",X"61",X"75",X"00",X"61",X"6B",X"00",X"61",X"63",X"00",X"33",X"FF",X"04",X"02",
		X"02",X"0C",X"08",X"0C",X"08",X"10",X"08",X"13",X"08",X"10",X"08",X"13",X"08",X"10",X"08",X"13",
		X"08",X"10",X"38",X"0A",X"02",X"00",X"63",X"FF",X"04",X"00",X"02",X"0C",X"18",X"12",X"18",X"13",
		X"18",X"14",X"18",X"16",X"38",X"17",X"02",X"00",X"73",X"FF",X"04",X"01",X"02",X"0A",X"68",X"09",
		X"03",X"48",X"09",X"03",X"08",X"09",X"03",X"68",X"09",X"03",X"48",X"0C",X"03",X"08",X"0B",X"03",
		X"48",X"0B",X"03",X"08",X"09",X"03",X"48",X"09",X"03",X"08",X"08",X"03",X"68",X"09",X"03",X"FF",
		X"02",X"0C",X"04",X"05",X"58",X"15",X"23",X"58",X"15",X"23",X"58",X"15",X"23",X"58",X"15",X"23",
		X"FF",X"4E",X"01",X"3C",X"01",X"2A",X"01",X"19",X"01",X"09",X"01",X"FB",X"00",X"EC",X"00",X"DF",
		X"00",X"D3",X"00",X"C7",X"00",X"BC",X"00",X"B1",X"00",X"A7",X"00",X"9E",X"00",X"95",X"00",X"8D",
		X"00",X"85",X"00",X"7D",X"00",X"76",X"00",X"70",X"00",X"69",X"00",X"63",X"00",X"5E",X"00",X"59",
		X"00",X"54",X"00",X"01",X"00",X"00",X"3A",X"00",X"B8",X"E5",X"E1",X"E5",X"E1",X"10",X"FA",X"0D",
		X"20",X"F4",X"C3",X"D1",X"02",X"E2",X"E3",X"E4",X"E5",X"E6",X"E7",X"E8",X"E9",X"EA",X"EB",X"EC",
		X"ED",X"EE",X"EF",X"F0",X"F1",X"F2",X"F3",X"F4",X"F5",X"F6",X"F7",X"3A",X"2D",X"80",X"B7",X"20",
		X"4C",X"21",X"1D",X"80",X"46",X"21",X"1F",X"80",X"6E",X"3E",X"08",X"80",X"67",X"3E",X"10",X"85",
		X"6F",X"01",X"06",X"06",X"CD",X"D9",X"41",X"DA",X"5A",X"3C",X"21",X"1D",X"80",X"46",X"21",X"1F",
		X"80",X"6E",X"3E",X"0E",X"80",X"67",X"3E",X"0F",X"85",X"6F",X"01",X"06",X"05",X"CD",X"D9",X"41",
		X"DA",X"5A",X"3C",X"21",X"1D",X"80",X"66",X"3A",X"1F",X"80",X"6F",X"3E",X"10",X"84",X"67",X"3E",
		X"08",X"85",X"6F",X"01",X"09",X"07",X"CD",X"D9",X"41",X"DA",X"5A",X"3C",X"C9",X"FE",X"01",X"20",
		X"46",X"21",X"1D",X"80",X"66",X"3A",X"1F",X"80",X"C6",X"10",X"6F",X"3E",X"09",X"84",X"67",X"01",
		X"07",X"08",X"CD",X"D9",X"41",X"DA",X"5A",X"3C",X"21",X"1D",X"80",X"66",X"3A",X"1F",X"80",X"C6",
		X"0E",X"6F",X"3E",X"0B",X"84",X"67",X"01",X"09",X"07",X"CD",X"D9",X"41",X"DA",X"5A",X"3C",X"21",
		X"1D",X"80",X"66",X"3A",X"1F",X"80",X"C6",X"04",X"6F",X"3E",X"0E",X"84",X"67",X"01",X"0A",X"09",
		X"CD",X"D9",X"41",X"DA",X"5A",X"3C",X"C9",X"FE",X"02",X"20",X"28",X"3A",X"1D",X"80",X"C6",X"0B",
		X"67",X"3A",X"1F",X"80",X"6F",X"01",X"0A",X"16",X"CD",X"D9",X"41",X"DA",X"5A",X"3C",X"3A",X"1D",
		X"80",X"C6",X"0D",X"67",X"3A",X"1F",X"80",X"C6",X"16",X"6F",X"01",X"06",X"08",X"CD",X"D9",X"41",
		X"38",X"7D",X"C9",X"FE",X"03",X"20",X"3D",X"3A",X"1D",X"80",X"C6",X"08",X"67",X"3A",X"1F",X"80",
		X"C6",X"04",X"6F",X"01",X"0A",X"09",X"CD",X"D9",X"41",X"38",X"64",X"3A",X"1D",X"80",X"C6",X"0C",
		X"67",X"3A",X"1F",X"80",X"C6",X"0E",X"6F",X"01",X"09",X"07",X"CD",X"D9",X"41",X"38",X"50",X"3A",
		X"1D",X"80",X"C6",X"11",X"67",X"3A",X"1F",X"80",X"C6",X"15",X"6F",X"01",X"06",X"08",X"CD",X"D9",
		X"41",X"38",X"3C",X"C9",X"3A",X"1D",X"80",X"C6",X"06",X"67",X"3A",X"1F",X"80",X"C6",X"08",X"6F",
		X"01",X"0B",X"07",X"CD",X"D9",X"41",X"38",X"27",X"3A",X"1D",X"80",X"C6",X"0B",X"67",X"3A",X"1F",
		X"80",X"C6",X"0F",X"6F",X"01",X"07",X"04",X"CD",X"D9",X"41",X"38",X"13",X"3A",X"1D",X"80",X"C6",
		X"12",X"67",X"3A",X"1F",X"80",X"C6",X"10",X"6F",X"01",X"06",X"07",X"CD",X"D9",X"41",X"D0",X"21",
		X"16",X"80",X"CB",X"DE",X"C9",X"1A",X"B7",X"C8",X"21",X"33",X"80",X"CB",X"6F",X"20",X"1A",X"E6",
		X"0F",X"A6",X"3E",X"00",X"C0",X"1A",X"FE",X"C3",X"20",X"15",X"21",X"23",X"80",X"7E",X"E6",X"03",
		X"C8",X"3E",X"01",X"CB",X"4E",X"C0",X"3E",X"FF",X"C9",X"E6",X"0F",X"A6",X"3E",X"00",X"C8",X"1A",
		X"CB",X"7F",X"3E",X"01",X"C0",X"3E",X"FF",X"C9",X"40",X"00",X"38",X"0F",X"30",X"1E",X"20",X"2D",
		X"F5",X"E5",X"D5",X"C5",X"11",X"5A",X"50",X"6F",X"26",X"00",X"29",X"29",X"19",X"7E",X"32",X"00",
		X"A8",X"23",X"3E",X"00",X"32",X"07",X"A0",X"3E",X"07",X"D3",X"08",X"3E",X"C0",X"D3",X"09",X"3E",
		X"0E",X"D3",X"08",X"7E",X"D3",X"09",X"23",X"3E",X"0F",X"D3",X"08",X"7E",X"D3",X"09",X"23",X"7E",
		X"32",X"00",X"B0",X"3E",X"FF",X"32",X"04",X"A0",X"3E",X"00",X"32",X"04",X"A0",X"CD",X"4A",X"50",
		X"3E",X"FF",X"32",X"04",X"A0",X"C1",X"D1",X"E1",X"F1",X"C9",X"06",X"01",X"21",X"10",X"00",X"2B",
		X"3A",X"00",X"B8",X"7C",X"B5",X"20",X"F8",X"10",X"F3",X"C9",X"40",X"00",X"7F",X"FF",X"50",X"10",
		X"7F",X"FF",X"80",X"28",X"7F",X"FF",X"30",X"40",X"7F",X"FF",X"80",X"4D",X"7F",X"FF",X"40",X"58",
		X"7F",X"FF",X"60",X"68",X"7F",X"FF",X"C0",X"70",X"7F",X"FF",X"30",X"80",X"7F",X"FF",X"80",X"C0",
		X"7F",X"FF",X"80",X"70",X"7F",X"FF",X"80",X"70",X"7F",X"FF",X"C9",X"3A",X"A1",X"81",X"FE",X"00",
		X"20",X"02",X"F1",X"C9",X"F1",X"CD",X"00",X"50",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F5",X"11",X"66",X"88",X"1A",X"FE",X"10",X"20",X"10",X"3A",X"00",X"83",X"B7",X"20",X"0E",X"3E",
		X"00",X"CD",X"8A",X"50",X"3E",X"0A",X"32",X"00",X"83",X"F1",X"C3",X"79",X"39",X"3A",X"00",X"83",
		X"3D",X"18",X"F3",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"CD",X"13",X"05",X"F5",X"E5",X"21",X"80",X"90",X"36",X"10",X"23",X"36",X"18",X"23",X"36",X"0A",
		X"23",X"36",X"15",X"E1",X"F1",X"C3",X"37",X"52",X"E5",X"21",X"00",X"00",X"22",X"1B",X"80",X"E1",
		X"C3",X"52",X"52",X"E5",X"21",X"00",X"00",X"22",X"1B",X"80",X"E1",X"C9",X"3E",X"22",X"CD",X"12",
		X"0D",X"CD",X"23",X"52",X"C3",X"79",X"52",X"E5",X"21",X"1B",X"92",X"36",X"0C",X"23",X"36",X"18",
		X"23",X"36",X"17",X"21",X"9B",X"92",X"36",X"15",X"23",X"36",X"1D",X"23",X"36",X"0D",X"E1",X"C3",
		X"CA",X"06",X"F5",X"3E",X"00",X"CD",X"8A",X"50",X"F1",X"C3",X"FE",X"34",X"F5",X"3A",X"00",X"83",
		X"B7",X"20",X"13",X"3E",X"02",X"CD",X"8A",X"50",X"3E",X"0A",X"32",X"00",X"83",X"F1",X"CB",X"4E",
		X"C2",X"DE",X"34",X"C3",X"B1",X"34",X"3D",X"18",X"F1",X"CD",X"D0",X"52",X"C3",X"80",X"40",X"00",
		X"F5",X"E5",X"D5",X"C5",X"3E",X"91",X"21",X"A6",X"90",X"06",X"04",X"0E",X"13",X"77",X"23",X"3C",
		X"0D",X"20",X"FA",X"11",X"0D",X"00",X"19",X"00",X"10",X"F1",X"21",X"86",X"9C",X"06",X"05",X"0E",
		X"13",X"36",X"12",X"23",X"0D",X"20",X"FA",X"11",X"0D",X"00",X"19",X"00",X"10",X"F1",X"C1",X"D1",
		X"E1",X"F1",X"C9",X"F5",X"E5",X"D5",X"C5",X"21",X"64",X"90",X"06",X"07",X"0E",X"16",X"36",X"35",
		X"23",X"0D",X"20",X"FA",X"11",X"0A",X"00",X"19",X"10",X"F2",X"C1",X"D1",X"E1",X"F1",X"C9",X"00",
		X"CD",X"B3",X"52",X"CD",X"80",X"52",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3E",X"09",X"CD",X"8A",X"50",X"CD",X"10",X"57",X"00",X"00",X"00",X"C3",X"00",X"57",X"00",X"00",
		X"F5",X"E5",X"D5",X"C5",X"06",X"01",X"21",X"00",X"00",X"23",X"3A",X"00",X"B8",X"3E",X"FF",X"BC",
		X"00",X"00",X"00",X"20",X"F4",X"10",X"EF",X"C1",X"D1",X"E1",X"F1",X"C9",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
