library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity rom_sprite_l is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of rom_sprite_l is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"35",X"00",X"AA",X"02",X"AA",X"0A",X"AA",X"0B",X"E9",
		X"00",X"00",X"40",X"00",X"40",X"00",X"5C",X"00",X"AA",X"00",X"AA",X"80",X"AA",X"A0",X"6B",X"E0",
		X"0B",X"E5",X"0A",X"A5",X"0A",X"E9",X"02",X"AA",X"02",X"A6",X"00",X"AA",X"00",X"0A",X"00",X"00",
		X"5B",X"E0",X"5A",X"A0",X"6B",X"A0",X"AA",X"80",X"9A",X"80",X"AA",X"00",X"A0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"04",X"00",X"01",X"00",X"35",X"00",X"AA",X"02",X"AA",X"0A",X"AA",X"0B",X"EB",
		X"00",X"00",X"10",X"00",X"40",X"00",X"5C",X"00",X"AA",X"00",X"AA",X"80",X"AA",X"A0",X"EB",X"E0",
		X"0B",X"EF",X"0A",X"AF",X"0A",X"6B",X"02",X"AA",X"02",X"AE",X"00",X"AA",X"00",X"0A",X"00",X"00",
		X"FB",X"E0",X"FA",X"A0",X"E9",X"A0",X"AA",X"80",X"BA",X"80",X"AA",X"00",X"A0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"14",X"00",X"01",X"00",X"35",X"00",X"AA",X"02",X"AA",X"0A",X"AA",X"09",X"6B",
		X"00",X"00",X"14",X"00",X"40",X"00",X"5C",X"00",X"AA",X"00",X"AA",X"80",X"AA",X"A0",X"E9",X"60",
		X"09",X"6F",X"0A",X"AF",X"0A",X"EB",X"02",X"AA",X"02",X"AE",X"00",X"AA",X"00",X"0A",X"00",X"00",
		X"F9",X"60",X"FA",X"A0",X"EB",X"A0",X"AA",X"80",X"BA",X"80",X"AA",X"00",X"A0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"2A",X"02",X"AB",X"0A",X"BB",X"0A",X"AA",X"29",X"A5",X"2A",X"95",
		X"00",X"00",X"00",X"00",X"A0",X"00",X"E8",X"00",X"EA",X"00",X"AA",X"C0",X"AA",X"40",X"6A",X"54",
		X"2A",X"95",X"29",X"A5",X"0A",X"AA",X"0A",X"BB",X"02",X"AB",X"00",X"2A",X"00",X"00",X"00",X"00",
		X"6A",X"54",X"AA",X"40",X"AA",X"C0",X"EA",X"00",X"E8",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"2A",X"02",X"AB",X"0A",X"9B",X"0A",X"AA",X"2B",X"AF",X"2A",X"BF",
		X"00",X"00",X"00",X"00",X"A0",X"00",X"E8",X"00",X"EA",X"00",X"AA",X"C0",X"AA",X"44",X"EA",X"50",
		X"2A",X"BF",X"2B",X"AF",X"0A",X"AA",X"0A",X"9B",X"02",X"AB",X"00",X"2A",X"00",X"00",X"00",X"00",
		X"EA",X"50",X"AA",X"44",X"AA",X"C0",X"EA",X"00",X"E8",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"2A",X"02",X"A9",X"0A",X"B9",X"0A",X"AA",X"2B",X"AF",X"2A",X"BF",
		X"00",X"00",X"00",X"00",X"A0",X"00",X"68",X"00",X"6A",X"00",X"AA",X"C4",X"AA",X"44",X"EA",X"50",
		X"2A",X"BF",X"2B",X"AF",X"0A",X"AA",X"0A",X"B9",X"02",X"A9",X"00",X"2A",X"00",X"00",X"00",X"00",
		X"EA",X"50",X"AA",X"44",X"AA",X"C4",X"6A",X"00",X"68",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"28",X"00",X"80",X"00",X"88",X"04",X"A1",X"04",X"35",X"04",X"AA",X"02",X"AA",X"0A",X"AE",
		X"28",X"00",X"02",X"00",X"22",X"00",X"48",X"10",X"5C",X"10",X"AA",X"10",X"AA",X"80",X"BA",X"A0",
		X"0A",X"AA",X"0A",X"AE",X"0A",X"AA",X"06",X"AE",X"06",X"AA",X"00",X"AE",X"00",X"0A",X"00",X"00",
		X"AA",X"A0",X"BA",X"A0",X"AA",X"A0",X"BA",X"90",X"AA",X"90",X"BA",X"00",X"A0",X"00",X"00",X"00",
		X"00",X"F0",X"02",X"00",X"02",X"30",X"00",X"81",X"04",X"B5",X"04",X"AA",X"02",X"AA",X"0A",X"AE",
		X"0F",X"00",X"00",X"80",X"0C",X"80",X"42",X"80",X"5E",X"10",X"AA",X"10",X"AA",X"80",X"BA",X"A0",
		X"0A",X"AA",X"0A",X"AE",X"0A",X"AA",X"02",X"AE",X"06",X"AA",X"04",X"AE",X"00",X"0A",X"00",X"00",
		X"AA",X"A0",X"BA",X"A0",X"AA",X"A0",X"BA",X"80",X"AA",X"90",X"BA",X"10",X"A0",X"00",X"00",X"00",
		X"02",X"80",X"08",X"00",X"08",X"C0",X"0A",X"01",X"02",X"35",X"04",X"AA",X"06",X"AA",X"0A",X"AE",
		X"02",X"80",X"00",X"20",X"03",X"20",X"40",X"A0",X"5C",X"80",X"AA",X"10",X"AA",X"90",X"BA",X"A0",
		X"0A",X"AA",X"0A",X"AE",X"0A",X"AA",X"02",X"AE",X"06",X"AA",X"04",X"AE",X"04",X"0A",X"00",X"00",
		X"AA",X"A0",X"BA",X"A0",X"AA",X"A0",X"BA",X"80",X"AA",X"90",X"BA",X"10",X"A0",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"6A",X"02",X"AA",X"0A",X"AA",X"0A",X"AA",X"2E",X"EE",X"2A",X"AA",
		X"00",X"00",X"00",X"00",X"85",X"40",X"A0",X"00",X"A8",X"A8",X"AB",X"82",X"E9",X"22",X"A9",X"40",
		X"2A",X"AA",X"2E",X"EE",X"0A",X"AA",X"0A",X"AA",X"02",X"AA",X"01",X"6A",X"00",X"00",X"00",X"00",
		X"A9",X"40",X"E9",X"22",X"AB",X"82",X"A8",X"28",X"A0",X"00",X"85",X"40",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"05",X"2A",X"02",X"AA",X"0A",X"AA",X"0A",X"AA",X"2E",X"EE",X"2A",X"AA",
		X"00",X"00",X"00",X"00",X"85",X"00",X"A0",X"28",X"AA",X"83",X"AB",X"33",X"E9",X"00",X"A9",X"40",
		X"2A",X"AA",X"2E",X"EE",X"0A",X"AA",X"0A",X"AA",X"02",X"AA",X"05",X"2A",X"00",X"00",X"00",X"00",
		X"A9",X"40",X"E9",X"00",X"AB",X"33",X"AA",X"83",X"A0",X"A8",X"85",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"15",X"2A",X"02",X"AA",X"0A",X"AA",X"0A",X"AA",X"2E",X"EE",X"2A",X"AA",
		X"00",X"00",X"00",X"00",X"94",X"A8",X"A2",X"82",X"A8",X"32",X"AB",X"00",X"E9",X"00",X"A9",X"40",
		X"2A",X"AA",X"2E",X"EE",X"0A",X"AA",X"0A",X"AA",X"02",X"AA",X"15",X"2A",X"00",X"00",X"00",X"00",
		X"A9",X"40",X"E9",X"00",X"AB",X"00",X"A8",X"32",X"A2",X"82",X"94",X"A8",X"00",X"00",X"00",X"00",
		X"03",X"F0",X"0C",X"3C",X"0C",X"3E",X"0F",X"FE",X"03",X"FA",X"00",X"A9",X"00",X"2A",X"00",X"09",
		X"0F",X"C0",X"30",X"F0",X"B0",X"F0",X"BF",X"F0",X"AF",X"C0",X"6A",X"00",X"A8",X"00",X"60",X"00",
		X"00",X"0A",X"00",X"09",X"00",X"5A",X"01",X"09",X"00",X"1A",X"00",X"49",X"01",X"02",X"00",X"00",
		X"A0",X"00",X"60",X"00",X"A5",X"00",X"60",X"40",X"A4",X"00",X"61",X"00",X"80",X"40",X"00",X"00",
		X"03",X"F0",X"0F",X"0C",X"0F",X"0E",X"0F",X"FE",X"03",X"FA",X"00",X"A9",X"02",X"AA",X"02",X"95",
		X"0F",X"C0",X"3C",X"30",X"BC",X"30",X"BF",X"F0",X"AF",X"C0",X"6A",X"00",X"AA",X"80",X"56",X"80",
		X"00",X"AA",X"04",X"95",X"01",X"AA",X"00",X"29",X"00",X"4A",X"05",X"09",X"00",X"02",X"00",X"00",
		X"AA",X"00",X"56",X"10",X"AA",X"40",X"68",X"00",X"A1",X"00",X"60",X"50",X"80",X"00",X"00",X"00",
		X"03",X"F0",X"0F",X"FC",X"0C",X"02",X"0F",X"FE",X"03",X"FA",X"00",X"A9",X"00",X"2A",X"00",X"09",
		X"0F",X"C0",X"3F",X"F0",X"80",X"30",X"BF",X"F0",X"AF",X"C0",X"6A",X"00",X"A8",X"00",X"60",X"00",
		X"04",X"2A",X"01",X"25",X"00",X"AA",X"04",X"95",X"01",X"AA",X"00",X"29",X"00",X"0A",X"00",X"00",
		X"A8",X"10",X"58",X"40",X"AA",X"00",X"56",X"10",X"AA",X"40",X"68",X"00",X"A0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"40",X"04",X"10",X"01",X"10",X"0A",X"AA",X"26",X"66",
		X"00",X"00",X"00",X"00",X"00",X"FC",X"03",X"C3",X"0B",X"C3",X"2B",X"FF",X"AA",X"FC",X"66",X"A0",
		X"26",X"66",X"0A",X"AA",X"01",X"10",X"04",X"10",X"10",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"A0",X"AA",X"FC",X"2B",X"C3",X"0B",X"C3",X"03",X"FF",X"00",X"FC",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"04",X"04",X"10",X"01",X"2A",X"00",X"A6",X"0A",X"A6",X"26",X"66",
		X"00",X"00",X"00",X"00",X"00",X"FC",X"A3",X"FF",X"AB",X"C3",X"6B",X"C3",X"6A",X"FC",X"66",X"A0",
		X"26",X"66",X"0A",X"A6",X"00",X"A6",X"01",X"2A",X"04",X"10",X"04",X"04",X"00",X"00",X"00",X"00",
		X"66",X"A0",X"6A",X"FC",X"6B",X"FF",X"AB",X"C3",X"A3",X"C3",X"00",X"FC",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"41",X"01",X"04",X"02",X"A0",X"0A",X"6A",X"2A",X"66",X"26",X"66",
		X"00",X"00",X"00",X"00",X"00",X"FC",X"03",X"CF",X"0B",X"CF",X"2B",X"CF",X"AA",X"CC",X"66",X"A0",
		X"26",X"66",X"2A",X"66",X"0A",X"6A",X"02",X"A0",X"01",X"04",X"00",X"41",X"00",X"00",X"00",X"00",
		X"66",X"A0",X"AA",X"CC",X"2B",X"CF",X"0B",X"CF",X"03",X"CF",X"00",X"FC",X"00",X"00",X"00",X"00",
		X"00",X"28",X"00",X"20",X"00",X"20",X"00",X"08",X"00",X"FE",X"00",X"3E",X"0C",X"3E",X"0F",X"FE",
		X"28",X"00",X"08",X"00",X"08",X"00",X"20",X"00",X"BF",X"00",X"83",X"C0",X"83",X"F0",X"BF",X"F0",
		X"00",X"2A",X"02",X"55",X"08",X"AA",X"08",X"55",X"00",X"2A",X"00",X"85",X"02",X"02",X"00",X"00",
		X"A8",X"00",X"55",X"80",X"AA",X"20",X"55",X"20",X"A8",X"00",X"52",X"00",X"80",X"80",X"00",X"00",
		X"00",X"A0",X"00",X"80",X"00",X"A0",X"00",X"08",X"00",X"FE",X"03",X"C2",X"0F",X"C2",X"0F",X"FE",
		X"0A",X"00",X"02",X"00",X"0A",X"00",X"20",X"00",X"BF",X"00",X"83",X"C0",X"83",X"F0",X"BF",X"F0",
		X"00",X"2A",X"00",X"05",X"02",X"2A",X"08",X"55",X"00",X"AA",X"02",X"55",X"08",X"2A",X"00",X"00",
		X"A8",X"00",X"50",X"00",X"A8",X"80",X"55",X"20",X"AA",X"00",X"55",X"80",X"A8",X"20",X"00",X"00",
		X"02",X"00",X"02",X"00",X"00",X"A0",X"00",X"08",X"00",X"FE",X"03",X"C2",X"0F",X"C2",X"0F",X"FE",
		X"00",X"80",X"00",X"80",X"0A",X"00",X"20",X"00",X"BF",X"00",X"BC",X"00",X"BC",X"30",X"BF",X"F0",
		X"00",X"2A",X"08",X"95",X"02",X"2A",X"00",X"05",X"02",X"8A",X"00",X"25",X"00",X"02",X"00",X"00",
		X"A8",X"00",X"56",X"20",X"A8",X"80",X"50",X"00",X"A2",X"80",X"58",X"00",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"A0",X"20",X"08",X"08",X"64",X"02",X"66",X"06",X"66",X"26",X"66",
		X"00",X"00",X"00",X"00",X"F0",X"00",X"C0",X"00",X"C3",X"00",X"FF",X"2A",X"FF",X"82",X"AA",X"00",
		X"26",X"66",X"06",X"66",X"02",X"66",X"08",X"64",X"20",X"08",X"00",X"A0",X"00",X"00",X"00",X"00",
		X"AA",X"00",X"C3",X"82",X"C3",X"2A",X"FF",X"00",X"FC",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"20",X"80",X"08",X"20",X"06",X"40",X"26",X"62",X"26",X"66",X"26",X"66",
		X"00",X"00",X"00",X"00",X"F0",X"00",X"FC",X"00",X"FF",X"2A",X"C3",X"22",X"C3",X"80",X"AA",X"00",
		X"26",X"66",X"26",X"66",X"26",X"62",X"06",X"40",X"08",X"20",X"20",X"80",X"00",X"00",X"00",X"00",
		X"AA",X"00",X"C3",X"80",X"C3",X"22",X"FF",X"2A",X"FC",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"08",X"02",X"20",X"02",X"08",X"08",X"26",X"06",X"66",X"26",X"66",
		X"00",X"00",X"00",X"00",X"F0",X"00",X"FC",X"0A",X"FF",X"20",X"C3",X"20",X"C3",X"80",X"AA",X"00",
		X"26",X"66",X"06",X"66",X"08",X"26",X"02",X"08",X"02",X"20",X"00",X"08",X"00",X"00",X"00",X"00",
		X"AA",X"00",X"FF",X"80",X"FF",X"20",X"C3",X"20",X"C0",X"0A",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"43",X"01",X"50",X"05",X"10",X"04",X"10",X"00",X"12",X"00",X"4A",X"00",X"6A",
		X"14",X"00",X"AA",X"C0",X"AA",X"00",X"28",X"00",X"A8",X"40",X"A0",X"50",X"A1",X"10",X"A9",X"10",
		X"00",X"AE",X"00",X"AA",X"05",X"AE",X"04",X"2A",X"04",X"2E",X"00",X"0A",X"00",X"02",X"00",X"00",
		X"BA",X"00",X"AA",X"00",X"BA",X"50",X"A8",X"10",X"B8",X"10",X"A0",X"00",X"80",X"00",X"00",X"00",
		X"00",X"01",X"00",X"3A",X"01",X"0A",X"05",X"42",X"04",X"42",X"04",X"12",X"00",X"1A",X"00",X"2A",
		X"40",X"00",X"AC",X"00",X"A0",X"40",X"81",X"50",X"81",X"10",X"84",X"10",X"A4",X"00",X"A8",X"00",
		X"00",X"AE",X"00",X"AA",X"00",X"AE",X"01",X"AA",X"04",X"BA",X"04",X"28",X"01",X"20",X"00",X"00",
		X"BA",X"00",X"AA",X"00",X"BA",X"00",X"AA",X"40",X"AE",X"10",X"28",X"10",X"08",X"40",X"00",X"00",
		X"00",X"14",X"03",X"AA",X"00",X"AA",X"00",X"28",X"01",X"2A",X"05",X"0A",X"04",X"4A",X"04",X"6A",
		X"00",X"00",X"C1",X"00",X"05",X"40",X"04",X"50",X"04",X"10",X"84",X"00",X"A1",X"00",X"A9",X"00",
		X"00",X"AE",X"00",X"AA",X"00",X"AE",X"01",X"2A",X"04",X"2E",X"01",X"0A",X"00",X"42",X"00",X"00",
		X"BA",X"00",X"AA",X"00",X"BA",X"00",X"A8",X"40",X"B8",X"10",X"A0",X"40",X"81",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"50",X"00",X"10",X"00",X"2A",X"02",X"AA",X"0B",X"BB",X"2A",X"AA",
		X"00",X"00",X"00",X"00",X"01",X"40",X"00",X"50",X"50",X"14",X"85",X"50",X"A0",X"00",X"A8",X"0C",
		X"2A",X"AA",X"0B",X"BB",X"02",X"AA",X"00",X"2A",X"00",X"10",X"01",X"50",X"00",X"00",X"00",X"00",
		X"AA",X"28",X"AA",X"A9",X"82",X"A9",X"50",X"28",X"05",X"0C",X"54",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"05",X"00",X"10",X"40",X"02",X"AA",X"2B",X"AA",X"0A",X"BB",X"02",X"AA",
		X"00",X"00",X"00",X"00",X"05",X"40",X"00",X"50",X"01",X"40",X"94",X"0C",X"A0",X"28",X"AA",X"A9",
		X"02",X"AA",X"0A",X"BB",X"2B",X"AA",X"02",X"AA",X"10",X"40",X"05",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"A9",X"A0",X"28",X"94",X"0C",X"01",X"40",X"00",X"50",X"05",X"40",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"04",X"40",X"10",X"2A",X"02",X"AA",X"0B",X"BB",X"2A",X"AA",
		X"00",X"00",X"00",X"00",X"54",X"00",X"05",X"0C",X"50",X"28",X"82",X"A9",X"AA",X"A9",X"AA",X"28",
		X"2A",X"AA",X"0B",X"BB",X"02",X"AA",X"10",X"2A",X"04",X"40",X"01",X"00",X"00",X"00",X"00",X"00",
		X"A8",X"0C",X"A0",X"00",X"85",X"50",X"50",X"14",X"00",X"50",X"01",X"40",X"00",X"00",X"00",X"00",
		X"00",X"08",X"00",X"0A",X"04",X"02",X"04",X"0E",X"04",X"2A",X"01",X"AA",X"02",X"AA",X"0A",X"AA",
		X"20",X"00",X"A0",X"00",X"80",X"10",X"B0",X"10",X"A8",X"10",X"AA",X"40",X"AA",X"80",X"AA",X"A0",
		X"03",X"FF",X"0A",X"AA",X"0A",X"AA",X"02",X"AA",X"04",X"AA",X"04",X"2A",X"01",X"0A",X"00",X"00",
		X"FF",X"C0",X"AA",X"A0",X"AA",X"A0",X"AA",X"80",X"AA",X"10",X"A8",X"10",X"A0",X"40",X"00",X"00",
		X"00",X"80",X"00",X"AA",X"00",X"02",X"01",X"0E",X"04",X"2A",X"01",X"AA",X"02",X"AA",X"0A",X"AA",
		X"02",X"00",X"AA",X"00",X"80",X"00",X"B0",X"40",X"A8",X"10",X"AA",X"40",X"AA",X"80",X"AA",X"A0",
		X"03",X"FF",X"0A",X"AA",X"0A",X"AA",X"02",X"AB",X"02",X"AB",X"04",X"AB",X"04",X"28",X"00",X"00",
		X"FF",X"C0",X"AA",X"A0",X"AA",X"A0",X"EA",X"80",X"EA",X"80",X"EA",X"10",X"28",X"10",X"00",X"00",
		X"08",X"00",X"0A",X"AA",X"00",X"02",X"04",X"0E",X"04",X"2A",X"04",X"AA",X"02",X"AA",X"0A",X"AA",
		X"00",X"20",X"AA",X"A0",X"80",X"00",X"B0",X"10",X"A8",X"10",X"AA",X"10",X"AA",X"80",X"AA",X"A0",
		X"03",X"FF",X"0A",X"AB",X"0A",X"AB",X"0A",X"AB",X"0A",X"AF",X"02",X"AF",X"04",X"A0",X"00",X"00",
		X"FF",X"C0",X"EA",X"A0",X"EA",X"A0",X"EA",X"A0",X"FA",X"A0",X"FA",X"80",X"0A",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"05",X"28",X"10",X"AB",X"02",X"AB",X"0A",X"AB",X"2A",X"AB",X"2A",X"AB",
		X"00",X"00",X"00",X"00",X"81",X"50",X"A4",X"00",X"A8",X"00",X"AA",X"00",X"AA",X"CA",X"AA",X"A8",
		X"2A",X"AB",X"2A",X"AB",X"0A",X"AB",X"02",X"AB",X"10",X"AB",X"05",X"28",X"00",X"00",X"00",X"00",
		X"AA",X"A8",X"AA",X"CA",X"AA",X"00",X"A8",X"00",X"A4",X"00",X"81",X"50",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"14",X"28",X"02",X"AB",X"0A",X"AB",X"2A",X"AB",X"2A",X"AB",X"0F",X"EB",
		X"00",X"00",X"00",X"00",X"81",X"00",X"A4",X"40",X"A8",X"0A",X"AA",X"08",X"AA",X"C8",X"AA",X"A8",
		X"0F",X"EB",X"2A",X"AB",X"2A",X"AB",X"0A",X"AB",X"02",X"AB",X"14",X"28",X"00",X"00",X"00",X"00",
		X"AA",X"A8",X"AA",X"C8",X"AA",X"08",X"A8",X"0A",X"A4",X"40",X"81",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"12",X"A8",X"0A",X"AB",X"2A",X"AB",X"2A",X"AB",X"0F",X"AB",X"0F",X"FF",
		X"00",X"00",X"00",X"00",X"85",X"4A",X"A0",X"08",X"A8",X"08",X"AA",X"08",X"AA",X"C8",X"AA",X"A8",
		X"0F",X"FF",X"0F",X"AB",X"2A",X"AB",X"2A",X"AB",X"0A",X"AB",X"12",X"A8",X"00",X"00",X"00",X"00",
		X"AA",X"A8",X"AA",X"C8",X"AA",X"08",X"A8",X"08",X"A0",X"08",X"85",X"4A",X"00",X"00",X"00",X"00",
		X"02",X"A3",X"00",X"0F",X"00",X"02",X"00",X"CA",X"03",X"1A",X"0C",X"16",X"0C",X"17",X"00",X"16",
		X"CA",X"80",X"F0",X"00",X"80",X"00",X"A3",X"00",X"A4",X"C0",X"94",X"30",X"D4",X"30",X"94",X"00",
		X"00",X"57",X"00",X"56",X"00",X"57",X"00",X"56",X"00",X"57",X"00",X"54",X"00",X"14",X"00",X"00",
		X"D5",X"00",X"95",X"00",X"D5",X"00",X"95",X"00",X"D5",X"00",X"15",X"00",X"14",X"00",X"00",X"00",
		X"00",X"A3",X"00",X"0F",X"0C",X"02",X"0C",X"CA",X"03",X"1A",X"00",X"56",X"00",X"57",X"01",X"5A",
		X"CA",X"00",X"F0",X"00",X"80",X"30",X"A3",X"30",X"A4",X"C0",X"95",X"00",X"D5",X"00",X"A5",X"40",
		X"01",X"5F",X"05",X"5A",X"05",X"5F",X"05",X"4A",X"05",X"43",X"05",X"00",X"04",X"00",X"00",X"00",
		X"F5",X"40",X"A5",X"50",X"F5",X"50",X"A1",X"50",X"C1",X"50",X"00",X"50",X"00",X"10",X"00",X"00",
		X"00",X"23",X"0C",X"8F",X"0C",X"02",X"03",X"CA",X"00",X"1A",X"01",X"56",X"01",X"57",X"05",X"52",
		X"C8",X"00",X"F2",X"30",X"80",X"30",X"A3",X"C0",X"A4",X"00",X"95",X"40",X"D5",X"40",X"85",X"50",
		X"05",X"5F",X"05",X"4A",X"05",X"7F",X"05",X"2A",X"05",X"3F",X"04",X"0A",X"00",X"03",X"00",X"00",
		X"F5",X"50",X"A1",X"50",X"FD",X"50",X"A8",X"50",X"FC",X"50",X"A0",X"10",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"55",X"15",X"55",X"15",X"55",X"03",X"BB",
		X"00",X"00",X"00",X"00",X"3C",X"00",X"03",X"02",X"00",X"C2",X"55",X"02",X"56",X"8C",X"BA",X"AF",
		X"03",X"BB",X"15",X"55",X"15",X"55",X"05",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"BA",X"AF",X"56",X"8C",X"55",X"02",X"00",X"C2",X"03",X"02",X"3C",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"15",X"54",X"05",X"55",X"01",X"55",X"00",X"15",X"00",X"BB",X"03",X"BB",
		X"00",X"00",X"00",X"00",X"00",X"F0",X"43",X"00",X"54",X"C2",X"55",X"02",X"96",X"8C",X"BA",X"AF",
		X"03",X"BB",X"00",X"BB",X"00",X"15",X"01",X"55",X"05",X"55",X"15",X"54",X"00",X"00",X"00",X"00",
		X"BA",X"AF",X"96",X"8C",X"55",X"02",X"54",X"C2",X"43",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"05",X"55",X"01",X"55",X"00",X"15",X"03",X"B1",X"0B",X"BB",X"3B",X"BB",
		X"00",X"00",X"00",X"00",X"40",X"3C",X"54",X"C0",X"54",X"C8",X"55",X"02",X"16",X"8C",X"BA",X"AF",
		X"3B",X"BB",X"0B",X"BB",X"03",X"B1",X"00",X"15",X"01",X"55",X"05",X"55",X"00",X"00",X"00",X"00",
		X"BA",X"AF",X"16",X"8C",X"55",X"02",X"54",X"C8",X"54",X"C0",X"40",X"3C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"02",X"A0",X"0A",X"A8",X"0B",X"C2",X"0B",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"0A",X"80",X"2A",X"A0",X"BC",X"20",X"BC",X"20",
		X"0B",X"FE",X"0A",X"FE",X"0A",X"AA",X"09",X"40",X"05",X"88",X"0A",X"64",X"01",X"A0",X"00",X"00",
		X"BF",X"E0",X"BF",X"A0",X"AA",X"A0",X"01",X"60",X"22",X"50",X"19",X"A0",X"0A",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"02",X"A0",X"0A",X"A8",X"0B",X"FE",X"0B",X"0E",X"0B",X"0E",
		X"00",X"00",X"00",X"00",X"02",X"00",X"0A",X"80",X"2A",X"A0",X"BF",X"E0",X"B0",X"E0",X"B0",X"E0",
		X"0A",X"FE",X"0A",X"AA",X"05",X"50",X"0A",X"80",X"05",X"40",X"02",X"90",X"00",X"58",X"00",X"00",
		X"BF",X"A0",X"AA",X"A0",X"05",X"50",X"02",X"A0",X"01",X"50",X"06",X"80",X"25",X"00",X"00",X"00",
		X"00",X"80",X"02",X"A0",X"0A",X"A8",X"08",X"3E",X"08",X"3E",X"0B",X"FE",X"0A",X"FE",X"0A",X"AA",
		X"02",X"00",X"0A",X"80",X"2A",X"A0",X"83",X"E0",X"83",X"E0",X"BF",X"E0",X"BF",X"A0",X"AA",X"A0",
		X"05",X"54",X"0A",X"A8",X"01",X"54",X"02",X"A8",X"00",X"54",X"00",X"28",X"00",X"04",X"00",X"00",
		X"15",X"50",X"2A",X"A0",X"15",X"40",X"2A",X"80",X"15",X"00",X"28",X"00",X"10",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"09",X"AA",X"19",X"6B",X"26",X"6F",X"28",X"2F",X"06",X"2F",X"00",X"2A",
		X"00",X"00",X"00",X"00",X"A8",X"00",X"FA",X"00",X"FA",X"80",X"0A",X"00",X"08",X"00",X"A0",X"00",
		X"00",X"2A",X"06",X"2F",X"28",X"2F",X"26",X"6F",X"19",X"6B",X"09",X"AA",X"00",X"00",X"00",X"00",
		X"A0",X"00",X"F8",X"00",X"FA",X"00",X"0A",X"80",X"0A",X"00",X"A8",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"9A",X"09",X"9A",X"19",X"9B",X"14",X"1B",X"20",X"0B",X"00",X"0A",
		X"00",X"00",X"00",X"00",X"AA",X"00",X"FE",X"80",X"0E",X"A0",X"0E",X"80",X"FE",X"00",X"A8",X"00",
		X"00",X"0A",X"20",X"0B",X"14",X"1B",X"19",X"9B",X"09",X"9A",X"01",X"9A",X"00",X"00",X"00",X"00",
		X"A8",X"00",X"FE",X"00",X"0E",X"80",X"0E",X"A0",X"FE",X"80",X"AA",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"99",X"01",X"99",X"09",X"99",X"19",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"AA",X"A0",X"AC",X"28",X"BC",X"2A",X"BF",X"E8",X"BF",X"E0",X"AA",X"80",
		X"00",X"00",X"19",X"99",X"09",X"99",X"01",X"99",X"00",X"99",X"00",X"09",X"00",X"00",X"00",X"00",
		X"AA",X"80",X"BC",X"20",X"BC",X"28",X"BF",X"EA",X"AF",X"E8",X"AA",X"A0",X"00",X"00",X"00",X"00",
		X"00",X"E0",X"03",X"F2",X"02",X"D4",X"00",X"55",X"02",X"15",X"08",X"25",X"00",X"81",X"00",X"08",
		X"80",X"00",X"08",X"00",X"20",X"00",X"80",X"80",X"42",X"00",X"58",X"00",X"54",X"A0",X"56",X"00",
		X"00",X"20",X"00",X"00",X"00",X"A1",X"00",X"05",X"00",X"95",X"02",X"15",X"00",X"04",X"00",X"00",
		X"54",X"00",X"54",X"A0",X"56",X"00",X"50",X"00",X"4A",X"00",X"80",X"80",X"20",X"00",X"00",X"00",
		X"00",X"03",X"02",X"0B",X"08",X"8F",X"00",X"25",X"02",X"05",X"08",X"85",X"00",X"25",X"02",X"05",
		X"C0",X"00",X"E0",X"80",X"F2",X"20",X"58",X"00",X"50",X"80",X"52",X"20",X"58",X"00",X"50",X"80",
		X"08",X"85",X"00",X"25",X"02",X"05",X"08",X"85",X"00",X"25",X"00",X"05",X"00",X"01",X"00",X"00",
		X"52",X"20",X"58",X"00",X"50",X"80",X"52",X"20",X"58",X"00",X"50",X"00",X"80",X"00",X"00",X"00",
		X"00",X"02",X"00",X"20",X"00",X"08",X"02",X"02",X"00",X"81",X"00",X"25",X"0A",X"15",X"00",X"95",
		X"0B",X"00",X"8F",X"C0",X"17",X"80",X"55",X"00",X"54",X"80",X"58",X"20",X"42",X"00",X"20",X"00",
		X"00",X"15",X"0A",X"15",X"00",X"95",X"00",X"05",X"00",X"A1",X"02",X"02",X"00",X"08",X"00",X"00",
		X"08",X"00",X"00",X"00",X"4A",X"00",X"50",X"00",X"56",X"00",X"54",X"80",X"10",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"02",X"20",X"05",X"22",X"15",X"40",X"05",X"50",
		X"00",X"00",X"00",X"00",X"08",X"00",X"02",X"2C",X"20",X"7F",X"09",X"5E",X"85",X"50",X"15",X"48",
		X"09",X"55",X"20",X"55",X"02",X"15",X"02",X"20",X"08",X"08",X"00",X"08",X"00",X"00",X"00",X"00",
		X"55",X"82",X"54",X"20",X"58",X"08",X"82",X"00",X"20",X"80",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"82",X"00",X"20",X"00",X"82",X"02",X"08",X"05",X"55",X"15",X"55",
		X"00",X"00",X"00",X"00",X"08",X"20",X"82",X"08",X"08",X"20",X"20",X"80",X"55",X"78",X"55",X"7F",
		X"15",X"55",X"05",X"55",X"02",X"08",X"00",X"82",X"00",X"20",X"00",X"82",X"00",X"00",X"00",X"00",
		X"55",X"7F",X"55",X"78",X"20",X"80",X"08",X"20",X"82",X"08",X"08",X"20",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"08",X"02",X"20",X"02",X"15",X"20",X"55",X"09",X"55",
		X"00",X"00",X"00",X"00",X"20",X"00",X"20",X"80",X"82",X"00",X"58",X"08",X"54",X"20",X"55",X"82",
		X"05",X"50",X"15",X"40",X"05",X"22",X"02",X"20",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"15",X"48",X"85",X"50",X"09",X"5E",X"20",X"7F",X"02",X"2C",X"08",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"30",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"30",
		X"00",X"00",X"00",X"00",X"F0",X"00",X"0C",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",X"0C",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"30",X"00",X"3F",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"FC",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"30",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"30",
		X"00",X"00",X"00",X"00",X"F0",X"00",X"0C",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",X"0C",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"30",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"00",X"00",X"00",X"3C",X"00",X"CC",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"30",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"30",
		X"00",X"00",X"00",X"00",X"F0",X"00",X"0C",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",X"0C",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"30",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"00",X"00",X"00",X"30",X"00",X"CC",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"AA",X"02",X"AA",X"02",X"AA",X"0A",X"AA",X"0A",X"AA",
		X"00",X"00",X"00",X"00",X"A0",X"00",X"A8",X"00",X"AA",X"00",X"AA",X"80",X"AA",X"88",X"AA",X"A0",
		X"0A",X"AA",X"0A",X"AA",X"02",X"AA",X"02",X"AA",X"00",X"AA",X"00",X"0A",X"00",X"00",X"00",X"00",
		X"AA",X"A0",X"AA",X"88",X"AA",X"80",X"AA",X"00",X"A8",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"AA",X"02",X"AA",X"02",X"AA",X"0A",X"AA",X"0A",X"AA",
		X"00",X"00",X"00",X"00",X"A0",X"00",X"AA",X"00",X"AA",X"80",X"AA",X"80",X"AA",X"A0",X"AA",X"A0",
		X"0A",X"AA",X"0A",X"AA",X"02",X"AA",X"02",X"AA",X"00",X"AA",X"00",X"0A",X"00",X"00",X"00",X"00",
		X"AA",X"A0",X"AA",X"A0",X"AA",X"80",X"AA",X"80",X"AA",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"2A",X"00",X"AA",X"02",X"AA",X"02",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"A8",X"00",X"AA",X"00",X"AA",X"80",X"AA",X"80",
		X"02",X"AA",X"02",X"AA",X"00",X"AA",X"00",X"2A",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"80",X"AA",X"80",X"AA",X"00",X"A8",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"2A",X"00",X"AA",X"00",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"A8",X"00",X"AA",X"00",X"AA",X"00",
		X"00",X"AA",X"00",X"AA",X"00",X"2A",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"00",X"AA",X"00",X"A8",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"0A",X"00",X"2A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"A0",X"00",X"A8",X"00",
		X"00",X"2A",X"00",X"0A",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A8",X"00",X"A0",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"0A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"A0",X"00",
		X"00",X"0A",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A0",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",
		X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
