library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity skyskip_sp_bits_3 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of skyskip_sp_bits_3 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FD",X"F9",X"7A",X"9C",X"80",X"40",X"E0",X"C0",X"80",X"80",X"CC",X"DC",X"FC",X"F4",
		X"F4",X"F4",X"F4",X"FC",X"F8",X"E0",X"C0",X"C0",X"E0",X"E0",X"F8",X"FE",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"DF",X"8F",X"0F",X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
		X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"02",X"04",X"04",X"00",X"00",X"00",
		X"01",X"01",X"01",X"01",X"01",X"81",X"42",X"E3",X"E3",X"80",X"C0",X"E1",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FC",X"78",X"B1",
		X"02",X"00",X"00",X"0E",X"1F",X"38",X"30",X"30",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"C0",X"70",X"1F",X"07",X"03",X"00",X"00",X"00",X"06",X"0F",X"3E",
		X"0F",X"0F",X"0F",X"0F",X"07",X"01",X"01",X"01",X"02",X"03",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"18",X"38",X"78",X"78",X"7C",X"7C",X"7C",X"72",X"3F",X"1F",X"0C",X"00",X"0F",X"00",
		X"00",X"E0",X"40",X"03",X"07",X"0F",X"1F",X"1B",X"1B",X"17",X"07",X"07",X"01",X"08",X"04",X"04",
		X"0C",X"00",X"01",X"0F",X"0F",X"0F",X"07",X"07",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"1F",X"0F",X"0F",X"0F",X"0F",X"9F",X"9F",X"DF",
		X"4F",X"67",X"67",X"63",X"ED",X"DF",X"FF",X"FF",X"FF",X"FE",X"FE",X"7C",X"78",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"03",X"06",X"0D",X"1B",X"17",X"37",X"2F",X"2F",X"27",X"33",X"1F",X"0E",
		X"F8",X"F0",X"F0",X"60",X"20",X"00",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"E0",X"E7",X"C1",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"9C",X"EF",X"EF",X"EF",X"DF",X"DF",X"BF",X"8F",X"07",X"07",X"07",X"8F",X"FF",X"7D",X"F9",X"F8",
		X"E0",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"83",X"80",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"83",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"78",X"78",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"02",X"02",X"05",X"00",X"00",
		X"0F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"1F",X"0F",X"03",
		X"00",X"00",X"80",X"C0",X"E0",X"E0",X"E0",X"E0",X"E0",X"C1",X"81",X"01",X"01",X"02",X"06",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"81",X"81",X"81",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"F7",X"F7",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"3F",X"3F",X"3F",X"3F",X"3F",X"38",
		X"04",X"1C",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CF",X"00",X"40",X"48",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"79",X"08",X"10",X"21",X"41",X"78",X"00",X"00",X"21",X"21",X"00",
		X"00",X"02",X"02",X"02",X"09",X"1C",X"3E",X"3F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"3F",X"DF",X"7F",X"3F",X"3F",X"1F",X"1F",X"1F",X"3F",X"3F",
		X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"3F",X"3F",X"3F",X"1F",X"1F",X"0F",X"07",X"4F",X"7F",
		X"7F",X"FF",X"FF",X"7F",X"3F",X"1F",X"0F",X"07",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"3F",X"1F",X"1F",X"1F",X"1F",X"3F",X"3F",X"7F",X"FF",X"FF",X"7F",X"3F",X"1F",X"0F",X"07",
		X"01",X"10",X"80",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"3F",X"3F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"7F",X"73",X"00",X"00",X"04",X"04",X"00",
		X"60",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F9",X"F9",X"FF",X"FF",X"FF",X"3E",X"0F",X"0F",
		X"83",X"89",X"C7",X"E3",X"FB",X"FF",X"FF",X"FF",X"FF",X"F9",X"FB",X"3F",X"07",X"07",X"03",X"03",
		X"3C",X"FC",X"FC",X"FC",X"F8",X"F8",X"F0",X"F0",X"E0",X"E0",X"F0",X"F8",X"FC",X"EC",X"C0",X"C0",
		X"60",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F8",X"F8",X"FC",X"7C",X"7E",X"3E",X"3E",
		X"60",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"78",X"78",X"3C",X"3C",X"3E",X"3E",X"0F",X"03",
		X"DE",X"CE",X"FE",X"FE",X"FE",X"FC",X"F8",X"F0",X"F0",X"E0",X"C0",X"00",X"00",X"80",X"80",X"80",
		X"83",X"89",X"C7",X"E3",X"FB",X"FF",X"FF",X"FF",X"FF",X"F9",X"FB",X"3F",X"87",X"87",X"83",X"83",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B3",X"B3",X"B3",X"B3",X"00",X"00",X"00",
		X"02",X"80",X"00",X"00",X"00",X"00",X"03",X"03",X"03",X"03",X"03",X"07",X"1F",X"1F",X"0E",X"06",
		X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"03",X"07",X"3F",X"7F",X"7E",X"7C",X"FC",X"F8",
		X"F1",X"F3",X"FF",X"FF",X"FF",X"FF",X"FB",X"FD",X"FE",X"FF",X"FE",X"FE",X"FE",X"7D",X"39",X"01",
		X"F1",X"F3",X"FF",X"FF",X"FF",X"FE",X"E1",X"E0",X"C1",X"81",X"03",X"03",X"03",X"20",X"A0",X"F4",
		X"F1",X"F3",X"FF",X"FF",X"FF",X"FF",X"FB",X"FD",X"FE",X"FF",X"FE",X"FE",X"FE",X"FC",X"38",X"00",
		X"0F",X"1F",X"1F",X"D7",X"93",X"1B",X"3E",X"AE",X"EE",X"EB",X"63",X"C7",X"0F",X"0F",X"0F",X"07",
		X"00",X"00",X"00",X"C0",X"80",X"10",X"30",X"B0",X"F0",X"F1",X"63",X"C7",X"0F",X"0F",X"07",X"07",
		X"0C",X"07",X"F7",X"F3",X"9F",X"90",X"61",X"03",X"03",X"07",X"07",X"0F",X"0E",X"06",X"03",X"01",
		X"03",X"00",X"F8",X"F8",X"9C",X"90",X"71",X"03",X"03",X"07",X"07",X"0F",X"0E",X"06",X"03",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"1F",X"3F",X"3C",X"78",X"7C",X"6C",X"48",
		X"41",X"40",X"60",X"30",X"1C",X"0F",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"1D",X"7F",X"7F",X"BF",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7E",X"7E",X"3F",X"3E",X"3E",X"3E",X"3C",X"3C",X"3C",X"7C",X"7C",X"7C",X"FE",X"FE",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"7F",X"3F",X"7F",X"3F",X"7F",X"5E",X"4C",X"C0",X"C0",X"90",X"10",X"10",X"90",
		X"FF",X"FF",X"FF",X"7F",X"3F",X"7F",X"3F",X"7F",X"5F",X"4F",X"C7",X"C3",X"93",X"13",X"10",X"90",
		X"C0",X"E0",X"E0",X"E0",X"E0",X"E0",X"C0",X"80",X"01",X"03",X"02",X"02",X"02",X"03",X"01",X"01",
		X"C0",X"E0",X"E0",X"E0",X"E0",X"E2",X"CE",X"99",X"37",X"6F",X"5F",X"5E",X"6E",X"3C",X"18",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"3F",X"7E",X"F8",X"F8",X"F0",X"E0",X"E0",X"E0",
		X"E0",X"C0",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"80",X"81",X"E1",X"C0",X"82",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"60",X"F1",X"F2",X"60",X"00",X"00",X"07",X"0F",X"1F",X"12",X"12",X"02",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"0F",X"0F",X"1F",X"1F",X"00",X"00",
		X"0F",X"1F",X"3F",X"3F",X"3F",X"3F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"3F",X"1F",X"00",X"00",
		X"00",X"00",X"00",X"0E",X"0E",X"0E",X"0C",X"0C",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"01",X"02",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"03",X"03",X"03",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"05",X"05",X"05",X"04",X"16",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"0F",X"0F",X"0F",X"07",X"03",X"00",
		X"10",X"10",X"08",X"00",X"00",X"00",X"0E",X"1F",X"3F",X"3F",X"3F",X"3F",X"1F",X"0E",X"00",X"00",
		X"10",X"10",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"3E",X"7F",X"7F",X"7F",X"7F",X"3E",X"1C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"7F",X"FF",X"FF",X"FF",X"FB",X"FB",X"FE",X"EE",X"0E",X"0F",X"1F",X"0F",X"07",X"07",
		X"00",X"00",X"C0",X"E0",X"F0",X"F0",X"F0",X"F8",X"FC",X"FC",X"FF",X"FF",X"FE",X"FC",X"FC",X"F8",
		X"07",X"03",X"03",X"01",X"00",X"00",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"E0",X"E7",X"E1",X"C0",
		X"F8",X"F0",X"F0",X"60",X"21",X"01",X"81",X"C0",X"C0",X"C0",X"C0",X"C0",X"E0",X"E7",X"C1",X"80",
		X"87",X"0D",X"1D",X"38",X"DD",X"DD",X"9D",X"1F",X"07",X"00",X"06",X"0C",X"1F",X"1F",X"03",X"13",
		X"00",X"00",X"61",X"27",X"18",X"18",X"00",X"00",X"00",X"00",X"06",X"0C",X"1E",X"1F",X"03",X"13",
		X"1E",X"1E",X"00",X"01",X"0F",X"1F",X"3F",X"17",X"07",X"06",X"02",X"02",X"01",X"00",X"00",X"00",
		X"28",X"2E",X"00",X"01",X"07",X"07",X"1F",X"1F",X"37",X"2D",X"09",X"00",X"00",X"00",X"00",X"00",
		X"2E",X"2E",X"00",X"01",X"0F",X"1F",X"3F",X"7F",X"9F",X"38",X"20",X"40",X"00",X"00",X"00",X"00",
		X"00",X"00",X"07",X"0F",X"0F",X"0F",X"0F",X"07",X"09",X"3C",X"7F",X"FF",X"FF",X"7F",X"B1",X"D0",
		X"1F",X"1F",X"1F",X"1F",X"0F",X"07",X"00",X"01",X"03",X"1F",X"3F",X"3F",X"3F",X"7F",X"FF",X"FF",
		X"E8",X"F0",X"F0",X"82",X"81",X"81",X"89",X"C9",X"FF",X"F7",X"74",X"14",X"0F",X"0F",X"0F",X"0F",
		X"FF",X"E7",X"93",X"09",X"01",X"E8",X"E6",X"07",X"C3",X"07",X"0F",X"9F",X"7F",X"0F",X"0F",X"0F",
		X"0F",X"1F",X"1F",X"1F",X"2F",X"2F",X"2F",X"EF",X"FF",X"7F",X"7F",X"7F",X"FB",X"F8",X"F0",X"F0",
		X"0F",X"17",X"17",X"17",X"1B",X"3B",X"3B",X"7F",X"7F",X"FF",X"7F",X"7F",X"7F",X"FB",X"F1",X"E0",
		X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"F8",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FC",X"F8",X"E0",X"80",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"F3",X"E7",X"EF",X"C3",X"80",X"00",X"00",
		X"0F",X"9F",X"FF",X"FE",X"FD",X"FB",X"F3",X"F7",X"F7",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"CF",X"EF",X"F7",X"FF",X"7F",X"7F",X"7F",X"7F",X"7F",X"3F",X"3F",X"1F",X"0F",X"0F",X"07",X"01",
		X"00",X"07",X"0F",X"1F",X"3F",X"7F",X"7F",X"7F",X"7F",X"3F",X"3F",X"3F",X"1F",X"0F",X"07",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"07",X"1F",X"7F",X"FF",X"7F",X"FF",X"7F",X"FF",X"07",X"00",X"01",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"E0",X"DF",X"DF",X"E3",X"FD",X"FD",X"ED",X"FD",X"FD",X"FD",X"FD",X"FE",X"FF",X"FF",
		X"FF",X"FF",X"07",X"FB",X"FB",X"DB",X"DB",X"FB",X"FB",X"DB",X"DB",X"FB",X"FB",X"07",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"7F",X"BF",X"BF",X"BD",X"BD",X"BF",X"BF",X"B8",X"BB",X"BB",X"7C",X"FF",X"FF",
		X"FF",X"C0",X"C0",X"CF",X"CF",X"CF",X"FF",X"FF",X"3F",X"1F",X"0F",X"07",X"03",X"03",X"03",X"03",
		X"00",X"00",X"01",X"1F",X"27",X"66",X"FE",X"FC",X"FC",X"78",X"70",X"B8",X"DC",X"DC",X"7E",X"3E",
		X"1F",X"3F",X"3F",X"7F",X"3F",X"1F",X"0F",X"16",X"46",X"67",X"76",X"76",X"7E",X"3E",X"1C",X"08",
		X"FE",X"FC",X"FF",X"67",X"0F",X"0E",X"1E",X"1C",X"1C",X"18",X"90",X"D8",X"DC",X"FC",X"7E",X"1E",
		X"1F",X"3F",X"3F",X"7F",X"3F",X"1F",X"0F",X"16",X"06",X"07",X"06",X"66",X"FE",X"FE",X"7E",X"1C",
		X"F8",X"3C",X"38",X"3F",X"3F",X"7F",X"7E",X"7F",X"7C",X"78",X"78",X"78",X"7C",X"7F",X"7E",X"76",
		X"6F",X"6B",X"79",X"FE",X"FF",X"FF",X"FF",X"DF",X"DF",X"5E",X"5F",X"CF",X"EF",X"ED",X"AD",X"06",
		X"FC",X"7C",X"3C",X"3F",X"7F",X"7F",X"7E",X"7F",X"7C",X"78",X"F8",X"F8",X"FC",X"FF",X"FE",X"76",
		X"6F",X"6B",X"79",X"3E",X"3F",X"3F",X"3F",X"1F",X"1F",X"1E",X"1F",X"0F",X"0D",X"0D",X"0F",X"06",
		X"7C",X"1E",X"06",X"04",X"05",X"47",X"EE",X"6E",X"7C",X"D8",X"B8",X"30",X"20",X"40",X"40",X"40",
		X"40",X"60",X"61",X"73",X"3F",X"3F",X"3F",X"1D",X"1D",X"0F",X"02",X"00",X"00",X"00",X"00",X"00",
		X"7C",X"1E",X"06",X"04",X"05",X"07",X"0E",X"0E",X"1C",X"18",X"38",X"30",X"20",X"40",X"40",X"40",
		X"40",X"60",X"61",X"73",X"3F",X"3F",X"3F",X"1F",X"1D",X"0F",X"02",X"00",X"00",X"00",X"00",X"00",
		X"1E",X"1F",X"1F",X"1F",X"00",X"00",X"02",X"07",X"07",X"05",X"05",X"02",X"00",X"00",X"00",X"00",
		X"7E",X"7E",X"32",X"00",X"1F",X"1F",X"1C",X"1E",X"1F",X"18",X"10",X"10",X"D0",X"F0",X"78",X"3C",
		X"1E",X"00",X"00",X"02",X"07",X"07",X"05",X"05",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"38",X"78",X"F8",X"E0",X"C0",X"1F",X"1F",X"1C",X"1E",X"1F",X"18",X"10",X"30",X"70",X"F0",X"D8",
		X"1C",X"1E",X"1F",X"1F",X"00",X"00",X"02",X"07",X"07",X"05",X"05",X"02",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"07",X"0E",X"0E",X"1E",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"03",X"02",X"02",X"02",X"01",X"00",X"30",X"78",X"38",X"78",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"02",X"00",X"00",X"02",X"09",X"05",X"02",X"02",X"30",X"78",X"38",X"78",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"3C",X"3C",X"3C",X"18",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"07",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"03",X"01",X"03",X"03",X"01",X"00",X"01",X"03",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"0F",X"1F",X"0F",X"00",X"10",X"18",X"0C",X"0F",X"07",X"02",X"00",X"00",
		X"00",X"00",X"00",X"01",X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"03",X"01",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"07",X"03",X"02",X"06",X"05",X"05",X"01",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"7E",X"7E",X"FF",X"FF",X"FD",X"FC",X"F8",X"7C",X"0E",X"07",
		X"00",X"00",X"00",X"00",X"07",X"3E",X"7E",X"7F",X"FF",X"FF",X"7F",X"3E",X"1C",X"0E",X"07",X"03",
		X"01",X"03",X"01",X"03",X"01",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"41",X"C3",X"67",X"7F",X"7F",X"3F",X"3F",X"1F",X"0F",X"03",
		X"40",X"C0",X"61",X"73",X"3F",X"3F",X"1F",X"0F",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"1B",X"1F",X"0F",X"0F",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"39",X"39",X"4F",X"4F",X"7F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"00",X"00",X"00",
		X"1F",X"27",X"27",X"7C",X"7C",X"7F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"00",
		X"1F",X"39",X"39",X"4F",X"4F",X"7F",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"00",X"0F",X"00",X"07",X"00",X"07",X"00",X"30",X"00",X"7C",X"00",X"3C",X"00",
		X"2A",X"00",X"7F",X"00",X"3F",X"00",X"0F",X"00",X"03",X"00",X"E0",X"00",X"FE",X"00",X"FE",X"00",
		X"FC",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"35",X"00",X"7F",X"00",X"3F",X"00",X"1F",X"00",X"07",X"00",X"FC",X"00",X"FE",X"00",X"7E",X"00",
		X"AA",X"00",X"FF",X"00",X"7F",X"00",X"BF",X"00",X"BF",X"00",X"DF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"7F",X"00",X"01",X"00",X"81",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"3C",X"00",X"0C",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"C0",X"C0",X"E0",X"60",X"70",X"30",X"3C",X"1E",X"0F",X"07",X"00",X"10",X"00",X"38",X"00",
		X"03",X"07",X"07",X"07",X"03",X"03",X"80",X"81",X"83",X"83",X"C1",X"C1",X"E0",X"F0",X"FC",X"FF",
		X"FF",X"7F",X"7F",X"1F",X"83",X"E1",X"60",X"30",X"30",X"18",X"1C",X"1E",X"0F",X"07",X"00",X"00",
		X"3C",X"00",X"3E",X"00",X"1F",X"00",X"1F",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"60",X"E0",X"F0",X"78",X"1C",X"06",X"06",X"0E",X"0E",X"0F",X"0F",X"07",X"07",X"03",X"81",
		X"F8",X"F8",X"F8",X"FC",X"FC",X"FE",X"FE",X"FE",X"7F",X"7F",X"7F",X"3F",X"1F",X"1F",X"1F",X"1F",
		X"0F",X"0F",X"07",X"C1",X"FF",X"FF",X"FF",X"FF",X"F7",X"E7",X"03",X"03",X"01",X"00",X"00",X"00",
		X"00",X"C0",X"00",X"C0",X"00",X"60",X"00",X"78",X"00",X"3E",X"00",X"07",X"00",X"00",X"00",X"00",
		X"FF",X"0F",X"E3",X"E3",X"F1",X"71",X"70",X"78",X"38",X"3C",X"1F",X"0F",X"07",X"01",X"00",X"00",
		X"FF",X"FF",X"FE",X"FC",X"FC",X"78",X"78",X"30",X"01",X"01",X"01",X"03",X"03",X"03",X"03",X"43",
		X"00",X"00",X"00",X"00",X"80",X"E0",X"FC",X"FE",X"FE",X"FC",X"FC",X"FC",X"F0",X"00",X"00",X"00",
		X"63",X"E3",X"E1",X"E1",X"F1",X"F1",X"F1",X"F0",X"F8",X"78",X"7C",X"3C",X"3F",X"1F",X"07",X"01",
		X"3F",X"0F",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"87",X"87",X"87",X"C3",X"C3",X"E3",X"61",X"71",X"71",X"38",X"3C",X"1F",X"0F",X"87",X"C3",X"E0",
		X"F0",X"7C",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"C6",X"C6",X"C6",X"C6",X"C6",X"C6",X"C6",X"C6",X"C6",X"C6",X"C6",X"DE",X"CE",X"DE",X"C6",
		X"FF",X"C6",X"C6",X"C6",X"C6",X"C6",X"C6",X"CE",X"CF",X"DE",X"C6",X"C6",X"C6",X"C6",X"C6",X"C6",
		X"C6",X"C6",X"C6",X"C6",X"C6",X"C6",X"C6",X"C6",X"C6",X"C6",X"C6",X"C6",X"C6",X"C6",X"C6",X"FF",
		X"C6",X"C6",X"C6",X"C6",X"C6",X"C6",X"C6",X"DE",X"FE",X"FE",X"FE",X"DE",X"C6",X"C6",X"C6",X"FF",
		X"00",X"00",X"00",X"18",X"18",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"09",X"0C",
		X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"C6",X"C6",X"C6",X"C7",X"DE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FE",X"DE",X"DE",X"CF",X"C7",
		X"FF",X"C6",X"C6",X"C6",X"C6",X"CE",X"FE",X"FE",X"FF",X"FF",X"F9",X"F8",X"F8",X"FC",X"FE",X"DF",
		X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",
		X"01",X"03",X"01",X"03",X"01",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F8",X"78",X"0C",X"0E",X"0E",X"07",X"87",X"83",X"C1",X"C0",X"E0",X"F0",X"7C",X"3F",
		X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"1F",X"07",X"01",X"00",X"04",X"06",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"0F",X"1F",X"3F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"3F",X"1F",X"0F",X"03",
		X"03",X"0F",X"1F",X"3F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"3F",X"1F",X"0F",X"03",
		X"00",X"70",X"70",X"70",X"0C",X"0C",X"02",X"00",X"00",X"02",X"0C",X"0C",X"70",X"70",X"70",X"00",
		X"17",X"7F",X"7F",X"B9",X"3B",X"77",X"7F",X"3F",X"9B",X"0F",X"1B",X"1D",X"9E",X"9F",X"4F",X"2F",
		X"00",X"01",X"03",X"01",X"00",X"10",X"08",X"08",X"09",X"0A",X"0C",X"04",X"02",X"01",X"00",X"00",
		X"00",X"00",X"00",X"40",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"20",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"1F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"1F",X"3F",X"3F",X"3F",X"3F",X"2F",X"3F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"20",X"40",X"90",X"E0",X"E0",X"FA",X"FE",X"FF",X"FE",X"FC",X"FC",X"FE",X"FF",X"FF",X"FF",
		X"40",X"80",X"00",X"90",X"E0",X"E0",X"F8",X"FE",X"FE",X"FE",X"FC",X"FC",X"FE",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"7F",X"1F",X"07",X"01",X"00",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"02",X"01",X"00",X"06",X"66",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"02",X"06",X"66",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"7F",X"FF",X"FF",X"FF",X"0F",X"17",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"01",X"03",X"01",X"01",X"01",X"03",X"07",X"17",X"07",X"0B",X"03",X"07",X"0E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"07",X"0A",X"1A",X"13",X"1F",X"4F",X"27",X"27",X"1F",X"7C",X"F9",X"F7",
		X"00",X"00",X"00",X"0F",X"07",X"0A",X"1A",X"13",X"1F",X"4F",X"27",X"27",X"1F",X"7C",X"F9",X"7F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"3F",X"3F",X"1F",X"1F",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"3F",X"3F",X"1F",X"1F",X"0F",
		X"00",X"00",X"20",X"33",X"1F",X"03",X"03",X"0D",X"01",X"01",X"07",X"0E",X"0E",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"02",X"02",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"02",X"02",X"02",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"18",X"38",X"78",X"F8",X"F0",X"F0",X"E0",X"F0",X"F8",X"F8",X"F0",X"F0",X"E0",X"E0",X"C0",X"C0",
		X"00",X"01",X"01",X"00",X"01",X"01",X"03",X"23",X"13",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"01",X"00",X"01",X"01",X"03",X"03",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"C0",X"80",X"88",X"88",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"07",X"01",X"01",X"00",
		X"00",X"00",X"00",X"01",X"3F",X"7E",X"FF",X"FF",X"FF",X"FF",X"DF",X"8E",X"04",X"00",X"00",X"00",
		X"00",X"80",X"D0",X"D0",X"C8",X"C8",X"20",X"20",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"41",X"23",X"03",X"03",X"05",X"04",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"03",X"03",X"0A",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"07",X"03",X"41",X"40",X"00",X"01",X"4B",X"1B",X"1B",X"1B",X"2D",X"0D",X"0D",
		X"00",X"00",X"03",X"07",X"03",X"01",X"00",X"00",X"01",X"8B",X"1B",X"9B",X"1B",X"2D",X"0D",X"0D",
		X"00",X"00",X"00",X"00",X"00",X"07",X"FF",X"FF",X"7F",X"1E",X"1F",X"3F",X"FF",X"FF",X"C3",X"C1",
		X"B9",X"70",X"F4",X"54",X"28",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0D",X"06",X"06",X"06",X"16",X"0F",X"03",X"08",X"00",X"00",X"04",X"04",X"00",X"00",X"00",X"00",
		X"0D",X"06",X"06",X"06",X"0E",X"27",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"20",X"20",X"00",X"00",X"00",X"10",X"02",X"06",X"06",X"06",X"06",X"06",X"06",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"06",X"26",X"06",X"26",X"06",X"06",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"F0",X"FC",X"7F",X"1F",X"3F",X"FF",X"FF",
		X"0F",X"0F",X"03",X"01",X"39",X"79",X"F1",X"54",X"24",X"58",X"20",X"00",X"00",X"00",X"00",X"00",
		X"06",X"06",X"06",X"06",X"06",X"02",X"10",X"08",X"08",X"00",X"20",X"20",X"00",X"03",X"01",X"00",
		X"06",X"0E",X"06",X"26",X"06",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"01",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
