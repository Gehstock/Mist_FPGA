library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity power_surge_prog is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of power_surge_prog is
	type rom is array(0 to  24575) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"F3",X"C3",X"00",X"30",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"08",X"D9",X"DD",X"E5",X"FD",X"E5",X"3E",X"01",X"32",X"00",
		X"C2",X"3A",X"A9",X"A8",X"FE",X"FF",X"20",X"05",X"3E",X"00",X"32",X"A9",X"A8",X"3A",X"A9",X"A8",
		X"E6",X"0F",X"32",X"A9",X"A8",X"3A",X"F5",X"A8",X"3C",X"32",X"F5",X"A8",X"E6",X"01",X"CA",X"DF",
		X"00",X"3A",X"F3",X"A8",X"FE",X"00",X"C2",X"B2",X"00",X"21",X"40",X"B0",X"11",X"10",X"B0",X"01",
		X"2F",X"00",X"ED",X"B0",X"21",X"40",X"B4",X"11",X"10",X"B4",X"01",X"2F",X"00",X"ED",X"B0",X"C3",
		X"DE",X"00",X"21",X"40",X"B0",X"11",X"10",X"B0",X"01",X"F0",X"18",X"7E",X"2F",X"D6",X"10",X"12",
		X"23",X"13",X"ED",X"A0",X"10",X"F5",X"21",X"40",X"B4",X"11",X"10",X"B4",X"01",X"F0",X"18",X"7E",
		X"EE",X"C0",X"12",X"23",X"13",X"7E",X"2F",X"D6",X"10",X"12",X"23",X"13",X"10",X"F1",X"00",X"3A",
		X"00",X"C3",X"E6",X"01",X"20",X"06",X"CD",X"19",X"01",X"C3",X"F1",X"00",X"3E",X"00",X"32",X"F6",
		X"A8",X"3A",X"00",X"C3",X"E6",X"02",X"20",X"06",X"CC",X"45",X"01",X"C3",X"03",X"01",X"3E",X"00",
		X"32",X"F7",X"A8",X"3A",X"04",X"60",X"E6",X"80",X"C8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FD",X"E1",X"DD",X"E1",X"D9",X"08",X"ED",X"45",X"3A",X"F6",X"A8",X"FE",X"00",X"28",X"01",
		X"C9",X"3E",X"01",X"CD",X"71",X"01",X"3E",X"40",X"32",X"F6",X"A8",X"21",X"FD",X"A8",X"35",X"C0",
		X"3A",X"B9",X"A8",X"47",X"3A",X"A9",X"A8",X"80",X"32",X"A9",X"A8",X"CD",X"44",X"4C",X"3A",X"B8",
		X"A8",X"32",X"FD",X"A8",X"C9",X"3A",X"F7",X"A8",X"FE",X"00",X"28",X"01",X"C9",X"3E",X"01",X"CD",
		X"71",X"01",X"3E",X"40",X"32",X"F7",X"A8",X"21",X"FE",X"A8",X"35",X"C0",X"3A",X"BB",X"A8",X"47",
		X"3A",X"A9",X"A8",X"80",X"32",X"A9",X"A8",X"CD",X"44",X"4C",X"3A",X"BA",X"A8",X"32",X"FE",X"A8",
		X"C9",X"32",X"00",X"C0",X"3E",X"FF",X"32",X"04",X"C3",X"3E",X"00",X"32",X"04",X"C3",X"C9",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C1",X"C2",X"00",X"00",X"00",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"2B",X"2B",X"2B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C3",X"C4",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"2B",X"2B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"19",X"11",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"1A",X"00",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"19",X"11",X"1A",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"00",X"00",X"00",X"28",X"27",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"19",X"11",X"24",
		X"0B",X"0B",X"0B",X"0B",X"07",X"07",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"00",X"2E",X"30",X"00",X"00",X"2D",X"2F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0B",X"0B",X"CF",X"CF",X"0B",X"0B",X"CF",X"CF",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"11",X"31",X"34",X"32",X"19",X"31",X"35",X"33",X"04",X"00",X"00",X"00",X"05",X"00",X"00",X"00",
		X"0B",X"0F",X"02",X"02",X"0B",X"0F",X"02",X"02",X"07",X"0B",X"0B",X"0B",X"07",X"0B",X"0B",X"0B",
		X"00",X"00",X"00",X"00",X"11",X"11",X"14",X"11",X"00",X"00",X"10",X"00",X"23",X"11",X"17",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"00",X"10",X"00",X"11",X"36",X"37",X"00",X"00",X"38",X"39",X"00",X"00",X"10",X"00",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0F",X"0F",X"0B",X"0B",X"0F",X"0F",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"21",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"18",X"11",X"11",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"14",X"11",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"12",X"11",X"11",X"11",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"10",X"00",X"0B",X"00",X"10",X"00",X"0C",X"51",X"10",X"00",X"00",X"00",X"12",X"11",X"1A",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"00",X"19",X"11",X"2E",X"30",X"08",X"00",X"2D",X"2F",X"10",X"00",X"00",X"00",X"18",X"11",
		X"0B",X"0B",X"0B",X"0B",X"CF",X"CF",X"0B",X"0B",X"CF",X"CF",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"11",X"17",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"11",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"00",X"10",X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"10",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"10",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"11",X"11",X"15",X"00",X"00",X"00",X"10",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"10",X"00",X"00",X"00",X"13",X"11",X"11",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"00",X"00",X"00",X"11",X"14",X"11",X"11",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"10",X"00",X"00",X"11",X"16",X"11",X"11",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"2E",X"30",X"08",X"00",X"2D",X"2F",X"10",X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"22",
		X"0B",X"CF",X"CF",X"0B",X"0B",X"CF",X"CF",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"22",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"13",X"11",X"1A",X"00",X"10",X"00",X"54",X"00",X"13",X"11",X"17",X"00",X"10",X"00",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"03",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"21",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"21",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"18",X"11",X"11",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"10",X"00",X"00",X"00",X"18",X"11",X"11",X"00",X"00",X"00",X"00",X"11",X"11",X"1A",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"00",X"00",X"10",X"11",X"11",X"11",X"12",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"00",X"10",X"00",X"11",X"11",X"15",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"00",X"00",X"00",X"11",X"24",X"23",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"10",X"00",X"00",X"11",X"16",X"11",X"11",X"00",X"21",X"00",X"00",X"00",X"22",X"00",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"00",X"00",X"00",X"28",X"27",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0B",X"0B",X"0B",X"0B",X"07",X"07",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"2E",X"30",X"08",X"00",X"2D",X"2F",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",
		X"CF",X"CF",X"0B",X"0B",X"CF",X"CF",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"10",X"00",X"00",X"00",X"18",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"14",X"00",X"00",X"00",X"25",X"00",X"00",X"00",X"26",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"07",X"0B",X"0B",X"0B",X"07",
		X"00",X"10",X"00",X"00",X"11",X"12",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"00",X"10",X"00",X"11",X"11",X"17",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"19",X"11",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"00",X"00",X"00",X"11",X"11",X"1A",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"00",X"00",X"00",X"28",X"27",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"19",X"11",X"11",
		X"0B",X"0B",X"0B",X"0B",X"07",X"07",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"11",X"00",X"00",X"00",X"00",X"11",X"24",X"23",X"11",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"00",X"00",X"00",X"11",X"14",X"11",X"11",X"00",X"10",X"00",X"00",X"11",X"15",X"00",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"10",X"00",X"00",X"00",X"12",X"11",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"00",X"10",X"00",X"11",X"11",X"16",X"11",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"00",X"0B",X"00",X"1A",X"00",X"0C",X"51",X"18",X"11",X"1A",X"00",X"00",X"00",X"10",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"00",X"00",X"00",X"31",X"28",X"27",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"07",X"07",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"00",X"10",X"00",X"24",X"23",X"17",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"22",X"00",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"10",X"00",X"00",X"11",X"12",X"14",X"11",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"10",X"00",X"00",X"00",X"12",X"11",X"1A",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"13",X"11",X"11",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"11",X"11",X"1A",X"00",X"2E",X"30",X"08",X"00",X"2D",X"2F",X"18",X"11",X"00",X"00",X"00",X"00",
		X"0B",X"0B",X"0B",X"0B",X"CF",X"CF",X"0B",X"0B",X"CF",X"CF",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"11",X"12",X"28",X"27",X"00",X"00",X"00",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"07",X"07",X"0B",X"0B",X"0B",X"0B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"24",X"23",X"11",X"00",X"00",X"00",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"00",X"18",X"11",X"00",X"00",X"00",X"00",X"11",X"24",X"23",X"11",X"00",X"00",X"00",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"11",X"11",X"1A",X"00",X"00",X"00",X"10",X"00",X"11",X"11",X"12",X"11",X"00",X"00",X"00",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"00",X"00",X"00",X"14",X"24",X"23",X"11",X"18",X"11",X"11",X"11",X"00",X"00",X"00",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"00",X"00",X"00",X"11",X"24",X"23",X"14",X"11",X"11",X"11",X"17",X"00",X"00",X"00",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"11",X"1A",X"00",X"50",X"00",X"0B",X"00",X"10",X"00",X"0C",X"11",X"17",X"00",X"00",X"00",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"00",X"00",X"00",X"11",X"11",X"14",X"11",X"00",X"00",X"04",X"00",X"00",X"00",X"05",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"07",X"0B",X"0B",X"0B",X"07",X"0B",
		X"00",X"00",X"00",X"10",X"28",X"27",X"11",X"16",X"00",X"00",X"00",X"10",X"00",X"19",X"11",X"17",
		X"0B",X"0B",X"0B",X"0B",X"07",X"07",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"00",X"13",X"11",X"00",X"00",X"21",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"10",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"24",X"23",X"11",X"1A",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"18",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"00",X"0B",X"00",X"00",X"00",X"0C",X"51",X"00",X"00",X"00",X"00",X"24",X"23",X"1A",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"10",X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"10",X"00",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"10",X"2E",X"30",X"00",X"10",X"2D",X"2F",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",
		X"0B",X"0B",X"CF",X"CF",X"0B",X"0B",X"CF",X"CF",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"13",X"11",X"00",X"00",X"10",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"1A",X"00",X"00",X"00",X"10",X"00",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"10",X"00",X"00",X"11",X"12",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"19",X"11",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"10",X"00",X"00",X"00",X"12",X"11",X"11",X"11",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"11",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"00",X"10",X"00",X"11",X"11",X"15",X"00",X"00",X"00",X"10",X"00",X"11",X"11",X"15",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"00",X"10",X"00",X"00",X"00",X"13",X"11",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"10",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"18",X"11",X"11",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"07",X"0B",X"0B",X"0B",X"07",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"24",X"23",X"11",X"24",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"23",X"11",X"17",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"13",X"11",X"11",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"11",X"11",X"11",X"41",X"00",X"3A",X"3C",X"02",X"00",X"3B",X"3D",X"02",X"00",X"00",X"00",X"02",
		X"0B",X"0B",X"0B",X"1A",X"0B",X"82",X"83",X"1A",X"0B",X"82",X"83",X"1A",X"0B",X"0B",X"0B",X"1A",
		X"41",X"47",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"19",X"11",X"11",X"02",X"10",X"02",X"02",
		X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"3E",X"3F",X"3F",X"3E",X"02",X"02",X"02",X"02",X"11",X"24",X"23",X"11",X"02",X"02",X"02",X"02",
		X"EA",X"EA",X"6A",X"6A",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"02",X"02",X"48",X"41",X"02",X"02",X"02",X"02",X"11",X"11",X"1A",X"02",X"02",X"02",X"10",X"02",
		X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"41",X"11",X"11",X"11",X"02",X"3C",X"3A",X"00",X"02",X"3D",X"3B",X"00",X"02",X"00",X"00",X"00",
		X"1A",X"0B",X"0B",X"0B",X"1A",X"03",X"02",X"0B",X"1A",X"03",X"02",X"0B",X"1A",X"0B",X"0B",X"0B",
		X"11",X"11",X"15",X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"10",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"00",X"00",X"02",X"09",X"3A",X"3C",X"11",X"0A",X"3B",X"3D",X"02",X"00",X"00",X"00",X"02",
		X"0B",X"0B",X"0B",X"1A",X"0B",X"82",X"83",X"22",X"0B",X"82",X"83",X"1A",X"0B",X"0B",X"0B",X"1A",
		X"00",X"00",X"00",X"02",X"00",X"3A",X"3C",X"02",X"00",X"3B",X"3D",X"02",X"00",X"00",X"00",X"02",
		X"0B",X"0B",X"0B",X"1A",X"0B",X"82",X"83",X"1A",X"0B",X"82",X"83",X"1A",X"0B",X"0B",X"0B",X"1A",
		X"02",X"00",X"00",X"00",X"11",X"3C",X"3A",X"09",X"02",X"3D",X"3B",X"0A",X"02",X"00",X"00",X"00",
		X"1A",X"0B",X"0B",X"0B",X"22",X"03",X"02",X"8B",X"1A",X"03",X"02",X"8B",X"1A",X"0B",X"0B",X"0B",
		X"02",X"00",X"00",X"00",X"02",X"3C",X"3A",X"00",X"02",X"3D",X"3B",X"00",X"02",X"00",X"00",X"00",
		X"1A",X"0B",X"0B",X"0B",X"1A",X"03",X"02",X"0B",X"1A",X"03",X"02",X"0B",X"1A",X"0B",X"0B",X"0B",
		X"00",X"00",X"00",X"00",X"06",X"07",X"1A",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",
		X"0B",X"0B",X"0B",X"0B",X"07",X"07",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"00",X"10",X"00",X"11",X"11",X"16",X"11",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"10",X"00",X"00",X"11",X"16",X"11",X"11",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"19",X"11",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"00",X"00",X"00",X"11",X"11",X"14",X"11",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"00",X"00",X"00",X"11",X"1A",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"10",X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"10",X"00",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"10",X"00",X"00",X"11",X"17",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"00",X"10",X"00",X"11",X"11",X"12",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"02",X"10",X"02",X"02",X"11",X"16",X"11",X"11",X"02",X"10",X"02",X"02",X"02",X"10",X"02",X"02",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"02",X"02",X"02",X"02",X"24",X"23",X"14",X"11",X"02",X"02",X"10",X"02",X"02",X"02",X"13",X"11",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"02",X"02",X"10",X"02",X"24",X"23",X"12",X"11",X"02",X"02",X"02",X"02",X"28",X"27",X"1A",X"02",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"2A",X"2A",X"22",X"22",
		X"02",X"10",X"02",X"02",X"02",X"13",X"28",X"27",X"02",X"10",X"02",X"02",X"02",X"10",X"02",X"02",
		X"22",X"22",X"22",X"22",X"22",X"22",X"2A",X"2A",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"02",X"02",X"10",X"02",X"11",X"36",X"37",X"02",X"02",X"38",X"39",X"02",X"02",X"10",X"02",X"02",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"02",X"02",X"10",X"02",X"02",X"02",X"21",X"02",X"02",X"02",X"22",X"02",X"02",X"02",X"10",X"02",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"02",X"10",X"02",X"02",X"02",X"13",X"24",X"23",X"02",X"18",X"28",X"27",X"02",X"02",X"02",X"02",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"2A",X"2A",X"22",X"22",X"22",X"22",
		X"02",X"10",X"02",X"02",X"11",X"16",X"11",X"11",X"11",X"17",X"02",X"02",X"02",X"02",X"02",X"02",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"02",X"02",X"10",X"02",X"24",X"23",X"12",X"11",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"02",X"10",X"02",X"19",X"11",X"16",X"11",X"12",X"02",X"10",X"02",X"02",X"02",X"10",X"02",X"02",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"11",X"11",X"11",X"11",X"11",X"11",X"14",X"11",X"02",X"02",X"21",X"02",X"02",X"02",X"22",X"02",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"1A",X"02",X"10",X"02",X"16",X"11",X"16",X"11",X"21",X"02",X"10",X"02",X"22",X"02",X"10",X"02",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"10",X"02",X"10",X"02",X"13",X"11",X"15",X"02",X"10",X"02",X"10",X"02",X"25",X"02",X"10",X"02",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"2A",X"22",X"22",X"22",
		X"02",X"10",X"02",X"02",X"02",X"13",X"24",X"23",X"02",X"10",X"02",X"02",X"02",X"18",X"11",X"11",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"02",X"10",X"02",X"02",X"11",X"12",X"11",X"11",X"02",X"02",X"02",X"02",X"11",X"24",X"23",X"11",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"26",X"02",X"10",X"02",X"17",X"02",X"13",X"11",X"02",X"02",X"10",X"02",X"11",X"11",X"17",X"02",
		X"2A",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"19",X"1A",X"00",X"50",X"10",X"0B",X"00",X"10",X"10",X"0C",X"11",X"17",X"10",X"00",X"00",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"18",X"11",X"1A",X"00",X"28",X"27",X"16",X"11",X"00",X"00",X"10",X"00",X"00",X"19",X"17",X"00",
		X"0B",X"0B",X"0B",X"0B",X"07",X"07",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"10",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"10",X"00",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"07",X"0B",X"0B",X"0B",X"07",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"10",X"00",X"00",X"00",X"18",X"11",X"14",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"2E",X"30",X"08",X"00",X"2D",X"2F",X"10",X"00",X"00",X"00",X"18",X"00",X"00",X"00",X"00",
		X"0B",X"CF",X"CF",X"0B",X"0B",X"CF",X"CF",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"11",X"00",X"00",X"00",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"24",X"23",X"11",X"00",X"00",X"00",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"06",X"07",X"00",X"00",X"00",X"00",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"07",X"07",X"0B",X"0B",X"0B",X"0B",
		X"00",X"31",X"34",X"32",X"19",X"31",X"35",X"33",X"17",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0B",X"0F",X"02",X"02",X"0B",X"0F",X"02",X"02",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"02",X"04",X"02",X"02",X"02",X"05",X"02",X"02",X"19",X"12",X"11",X"24",X"10",X"02",X"02",X"02",
		X"22",X"2A",X"22",X"22",X"22",X"2A",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"02",X"04",X"19",X"11",X"02",X"05",X"13",X"11",X"23",X"17",X"13",X"11",X"02",X"02",X"13",X"11",
		X"22",X"2A",X"22",X"22",X"22",X"2A",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"11",X"11",X"11",X"1A",X"11",X"11",X"1A",X"10",X"11",X"1A",X"10",X"10",X"1A",X"10",X"10",X"10",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"19",X"28",X"27",X"1A",X"10",X"19",X"1A",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"22",X"2A",X"2A",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"10",X"02",X"02",X"02",X"16",X"11",X"28",X"27",X"10",X"02",X"02",X"02",X"10",X"02",X"02",X"02",
		X"22",X"22",X"22",X"22",X"22",X"22",X"2A",X"2A",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"21",X"21",X"21",X"21",X"22",X"22",X"22",X"22",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"18",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"10",X"21",X"21",X"10",X"10",X"22",X"22",X"10",X"10",X"10",X"10",X"10",X"17",X"10",X"10",X"10",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"10",X"02",X"02",X"02",X"10",X"02",X"02",X"02",X"10",X"02",X"02",X"02",X"10",X"02",X"02",X"02",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"02",X"18",X"11",X"11",X"02",X"02",X"02",X"02",X"02",X"02",X"19",X"11",X"02",X"02",X"10",X"02",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"12",X"15",X"18",X"11",X"02",X"18",X"11",X"28",X"11",X"11",X"11",X"11",X"19",X"11",X"11",X"24",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"2A",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"11",X"17",X"10",X"10",X"27",X"11",X"15",X"10",X"11",X"11",X"15",X"10",X"23",X"11",X"15",X"10",
		X"22",X"22",X"22",X"22",X"2A",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"10",X"02",X"02",X"02",X"13",X"11",X"28",X"27",X"13",X"11",X"1A",X"02",X"13",X"1A",X"10",X"02",
		X"22",X"22",X"22",X"22",X"22",X"22",X"2A",X"2A",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"10",X"02",X"02",X"02",X"10",X"02",X"02",X"19",X"04",X"02",X"02",X"04",X"05",X"02",X"02",X"05",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"2A",X"22",X"22",X"2A",X"2A",X"22",X"22",X"2A",
		X"02",X"02",X"10",X"10",X"11",X"11",X"15",X"10",X"02",X"02",X"04",X"10",X"02",X"02",X"05",X"10",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"2A",X"22",X"22",X"22",X"2A",X"22",
		X"21",X"21",X"21",X"02",X"22",X"22",X"22",X"02",X"10",X"10",X"18",X"11",X"10",X"18",X"11",X"11",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"02",X"04",X"02",X"02",X"02",X"05",X"02",X"02",X"11",X"17",X"02",X"02",X"11",X"24",X"23",X"11",
		X"22",X"2A",X"22",X"22",X"22",X"2A",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"10",X"02",X"02",X"10",X"10",X"02",X"02",X"13",X"10",X"02",X"02",X"10",X"17",X"02",X"02",X"13",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"02",X"02",X"10",X"10",X"24",X"23",X"15",X"10",X"02",X"02",X"10",X"10",X"24",X"23",X"15",X"10",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"10",X"02",X"02",X"02",X"15",X"02",X"02",X"02",X"10",X"02",X"02",X"02",X"18",X"11",X"24",X"23",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"02",X"02",X"02",X"02",X"02",X"02",X"19",X"11",X"02",X"02",X"10",X"02",X"11",X"11",X"12",X"11",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"02",X"02",X"02",X"10",X"11",X"11",X"11",X"12",X"02",X"02",X"02",X"02",X"11",X"11",X"11",X"11",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"02",X"02",X"10",X"10",X"24",X"23",X"17",X"10",X"02",X"02",X"02",X"10",X"11",X"11",X"11",X"17",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"02",X"02",X"3E",X"3F",X"02",X"02",X"02",X"02",X"11",X"11",X"14",X"11",X"02",X"02",X"10",X"02",
		X"22",X"22",X"EA",X"EA",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"3F",X"3E",X"48",X"41",X"02",X"02",X"02",X"02",X"11",X"24",X"23",X"11",X"02",X"02",X"02",X"02",
		X"6A",X"6A",X"1A",X"1A",X"32",X"32",X"32",X"32",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"41",X"41",X"41",X"41",X"02",X"02",X"02",X"02",X"11",X"11",X"1A",X"02",X"02",X"02",X"10",X"02",
		X"1A",X"1A",X"1A",X"1A",X"32",X"32",X"32",X"32",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"41",X"11",X"17",X"00",X"02",X"3C",X"3A",X"00",X"02",X"3D",X"3B",X"00",X"02",X"00",X"00",X"00",
		X"1A",X"0B",X"0B",X"0B",X"1A",X"03",X"02",X"0B",X"1A",X"03",X"02",X"0B",X"1A",X"0B",X"0B",X"0B",
		X"10",X"10",X"10",X"02",X"18",X"12",X"12",X"11",X"02",X"19",X"11",X"11",X"02",X"10",X"02",X"02",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"00",X"10",X"00",X"00",X"00",X"18",X"11",X"1A",X"00",X"00",X"00",X"25",X"00",X"00",X"00",X"26",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"07",X"0B",X"0B",X"0B",X"07",
		X"02",X"10",X"02",X"02",X"14",X"12",X"28",X"27",X"10",X"02",X"02",X"02",X"10",X"02",X"02",X"02",
		X"22",X"22",X"22",X"22",X"22",X"22",X"2A",X"2A",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"02",X"02",X"02",X"02",X"02",X"19",X"11",X"11",X"02",X"10",X"02",X"02",X"02",X"10",X"02",X"02",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"02",X"02",X"10",X"02",X"11",X"11",X"17",X"02",X"19",X"24",X"23",X"1A",X"10",X"02",X"02",X"10",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"10",X"02",X"02",X"02",X"10",X"02",X"02",X"02",X"13",X"11",X"11",X"24",X"10",X"02",X"02",X"02",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"11",X"12",X"11",X"11",X"11",X"24",X"23",X"11",X"11",X"11",X"11",X"11",X"1A",X"02",X"02",X"02",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"17",X"02",X"02",X"10",X"11",X"11",X"11",X"15",X"11",X"11",X"1A",X"10",X"02",X"02",X"10",X"10",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"02",X"10",X"02",X"02",X"11",X"12",X"1A",X"02",X"11",X"1A",X"10",X"02",X"02",X"10",X"18",X"11",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"10",X"02",X"02",X"10",X"18",X"11",X"11",X"16",X"02",X"02",X"02",X"10",X"11",X"24",X"23",X"12",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"02",X"02",X"10",X"10",X"24",X"23",X"17",X"10",X"02",X"02",X"02",X"10",X"11",X"11",X"11",X"17",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0C",X"A0",X"00",X"01",X"01",X"01",X"01",X"04",X"01",X"08",X"05",X"FF",X"FF",X"FF",X"FF",X"00",
		X"01",X"02",X"03",X"06",X"07",X"04",X"05",X"08",X"09",X"0A",X"0B",X"0C",X"0D",X"1A",X"5F",X"5E",
		X"60",X"5D",X"61",X"50",X"14",X"09",X"62",X"11",X"11",X"1A",X"11",X"0E",X"25",X"5E",X"64",X"5D",
		X"63",X"50",X"14",X"21",X"22",X"23",X"09",X"1B",X"24",X"25",X"26",X"27",X"21",X"27",X"15",X"28",
		X"0C",X"A0",X"00",X"02",X"02",X"02",X"02",X"04",X"01",X"08",X"05",X"FF",X"FF",X"FF",X"FF",X"1B",
		X"1B",X"06",X"07",X"29",X"21",X"2A",X"2B",X"2C",X"2D",X"2E",X"2F",X"21",X"30",X"51",X"52",X"53",
		X"54",X"55",X"56",X"57",X"14",X"58",X"65",X"66",X"67",X"5A",X"28",X"45",X"59",X"68",X"69",X"6A",
		X"5B",X"1B",X"1A",X"59",X"6B",X"6C",X"6D",X"5A",X"2A",X"25",X"26",X"15",X"21",X"15",X"15",X"28",
		X"0C",X"A0",X"00",X"04",X"03",X"03",X"03",X"04",X"01",X"08",X"05",X"FF",X"FF",X"FF",X"FF",X"3E",
		X"3F",X"29",X"21",X"40",X"15",X"2A",X"41",X"15",X"09",X"1B",X"42",X"43",X"44",X"45",X"1B",X"46",
		X"07",X"47",X"48",X"11",X"14",X"21",X"49",X"4A",X"4B",X"1A",X"11",X"14",X"23",X"09",X"1B",X"4C",
		X"27",X"20",X"1A",X"1B",X"4D",X"4E",X"4F",X"1B",X"50",X"25",X"26",X"15",X"21",X"15",X"15",X"28",
		X"0C",X"A0",X"00",X"04",X"04",X"04",X"04",X"04",X"01",X"08",X"05",X"FF",X"FF",X"FF",X"FF",X"1B",
		X"1B",X"06",X"07",X"29",X"21",X"2A",X"2B",X"2C",X"2D",X"2E",X"2F",X"21",X"30",X"1A",X"1B",X"14",
		X"23",X"09",X"31",X"32",X"33",X"1B",X"33",X"1B",X"33",X"06",X"07",X"0E",X"1B",X"14",X"21",X"34",
		X"15",X"35",X"36",X"37",X"38",X"39",X"3A",X"3B",X"13",X"25",X"26",X"15",X"3C",X"3D",X"15",X"28",
		X"0C",X"A0",X"00",X"05",X"05",X"05",X"05",X"04",X"01",X"08",X"05",X"FF",X"FF",X"FF",X"FF",X"1B",
		X"1B",X"02",X"03",X"06",X"07",X"04",X"05",X"08",X"09",X"0A",X"0B",X"0C",X"0D",X"51",X"52",X"53",
		X"54",X"55",X"56",X"57",X"14",X"58",X"6E",X"6F",X"70",X"5A",X"28",X"45",X"59",X"68",X"69",X"71",
		X"5B",X"1B",X"1A",X"59",X"72",X"73",X"74",X"5A",X"5C",X"25",X"26",X"15",X"3C",X"3D",X"15",X"28",
		X"0C",X"A0",X"00",X"06",X"06",X"06",X"06",X"04",X"01",X"08",X"05",X"FF",X"FF",X"FF",X"FF",X"1B",
		X"1B",X"06",X"07",X"29",X"21",X"2A",X"2B",X"2C",X"2D",X"2E",X"2F",X"21",X"30",X"0E",X"0F",X"10",
		X"03",X"11",X"12",X"13",X"14",X"15",X"16",X"17",X"09",X"18",X"19",X"1A",X"1B",X"1C",X"1D",X"1E",
		X"1F",X"20",X"14",X"21",X"22",X"23",X"09",X"1B",X"24",X"25",X"26",X"27",X"21",X"27",X"15",X"28",
		X"0C",X"A0",X"00",X"07",X"07",X"07",X"07",X"04",X"01",X"08",X"05",X"FF",X"FF",X"FF",X"FF",X"75",
		X"59",X"7E",X"7F",X"80",X"81",X"5B",X"76",X"58",X"82",X"69",X"83",X"84",X"5B",X"77",X"59",X"85",
		X"86",X"87",X"88",X"5B",X"1A",X"59",X"89",X"69",X"8A",X"8B",X"5B",X"45",X"59",X"8C",X"8D",X"8E",
		X"8F",X"5B",X"78",X"58",X"90",X"91",X"92",X"93",X"5B",X"79",X"7A",X"7B",X"7B",X"7B",X"7C",X"7D",
		X"0C",X"A0",X"00",X"08",X"08",X"08",X"08",X"04",X"01",X"08",X"05",X"FF",X"FF",X"FF",X"FF",X"1B",
		X"1B",X"02",X"03",X"06",X"07",X"04",X"05",X"08",X"09",X"0A",X"0B",X"0C",X"0D",X"51",X"52",X"53",
		X"94",X"95",X"96",X"97",X"14",X"58",X"9A",X"69",X"9B",X"9C",X"5B",X"45",X"59",X"9D",X"7F",X"9E",
		X"9F",X"5B",X"1A",X"59",X"89",X"69",X"8A",X"8B",X"5B",X"99",X"59",X"98",X"A0",X"A1",X"A2",X"5B",
		X"0C",X"A0",X"00",X"09",X"09",X"09",X"09",X"04",X"01",X"08",X"05",X"FF",X"FF",X"FF",X"FF",X"3E",
		X"3F",X"29",X"21",X"40",X"15",X"2A",X"41",X"15",X"09",X"1B",X"42",X"43",X"44",X"45",X"1B",X"46",
		X"07",X"47",X"48",X"11",X"14",X"21",X"49",X"4A",X"4B",X"1A",X"11",X"14",X"23",X"09",X"1B",X"4C",
		X"27",X"20",X"36",X"37",X"38",X"39",X"3A",X"3B",X"13",X"25",X"26",X"15",X"3C",X"3D",X"15",X"28",
		X"0C",X"A0",X"00",X"01",X"01",X"01",X"01",X"04",X"01",X"08",X"05",X"FF",X"FF",X"FF",X"FF",X"1B",
		X"1B",X"06",X"07",X"29",X"21",X"2A",X"2B",X"2C",X"2D",X"2E",X"2F",X"21",X"30",X"45",X"1B",X"46",
		X"07",X"47",X"48",X"11",X"14",X"21",X"49",X"4A",X"4B",X"1A",X"11",X"14",X"23",X"09",X"1B",X"4C",
		X"27",X"20",X"36",X"37",X"38",X"39",X"3A",X"3B",X"13",X"25",X"26",X"15",X"3C",X"3D",X"15",X"28",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"31",X"40",X"A0",X"C3",X"19",X"32",X"CD",X"EA",X"3D",X"CD",X"4A",X"3E",X"CD",X"59",X"3D",X"CD",
		X"76",X"3C",X"CD",X"BA",X"3C",X"CD",X"50",X"41",X"CD",X"F5",X"37",X"3E",X"05",X"32",X"10",X"A8",
		X"06",X"14",X"C5",X"CD",X"1D",X"38",X"01",X"00",X"08",X"0D",X"20",X"FD",X"10",X"FB",X"C1",X"10",
		X"F1",X"3A",X"C1",X"A8",X"FE",X"02",X"20",X"13",X"21",X"10",X"32",X"06",X"2C",X"11",X"A9",X"A7",
		X"CD",X"DB",X"36",X"3A",X"9A",X"A8",X"C6",X"B0",X"32",X"E9",X"A6",X"21",X"04",X"32",X"06",X"2C",
		X"11",X"AB",X"A7",X"CD",X"DB",X"36",X"21",X"0C",X"32",X"06",X"2C",X"11",X"6D",X"A7",X"CD",X"DB",
		X"36",X"01",X"00",X"F0",X"0D",X"20",X"FD",X"10",X"FB",X"21",X"F0",X"31",X"11",X"40",X"B0",X"01",
		X"0A",X"00",X"ED",X"B0",X"21",X"FA",X"31",X"11",X"40",X"B4",X"01",X"0A",X"00",X"ED",X"B0",X"3E",
		X"02",X"32",X"10",X"A8",X"DD",X"21",X"41",X"B4",X"06",X"05",X"DD",X"35",X"00",X"DD",X"23",X"DD",
		X"23",X"10",X"F7",X"01",X"00",X"0C",X"0D",X"20",X"FD",X"10",X"FB",X"3A",X"45",X"B0",X"FE",X"FF",
		X"28",X"1D",X"3A",X"10",X"A8",X"3D",X"32",X"10",X"A8",X"20",X"14",X"3E",X"04",X"32",X"10",X"A8",
		X"3A",X"45",X"B0",X"06",X"13",X"FE",X"13",X"20",X"02",X"06",X"16",X"78",X"32",X"45",X"B0",X"3A",
		X"41",X"B4",X"FE",X"E8",X"CC",X"DF",X"30",X"FE",X"D8",X"CC",X"E5",X"30",X"FE",X"C8",X"CC",X"EB",
		X"30",X"FE",X"B8",X"CC",X"F1",X"30",X"FE",X"A0",X"CA",X"F7",X"30",X"C3",X"84",X"30",X"C9",X"3E",
		X"12",X"32",X"43",X"B0",X"C9",X"3E",X"13",X"32",X"45",X"B0",X"C9",X"3E",X"14",X"32",X"47",X"B0",
		X"C9",X"3E",X"15",X"32",X"49",X"B0",X"C9",X"CD",X"F1",X"49",X"3E",X"01",X"32",X"98",X"A8",X"3E",
		X"01",X"32",X"09",X"A8",X"3E",X"BC",X"32",X"52",X"B0",X"32",X"54",X"B0",X"3E",X"02",X"32",X"52",
		X"B4",X"32",X"54",X"B4",X"3E",X"90",X"32",X"53",X"B4",X"3E",X"A0",X"32",X"55",X"B4",X"3E",X"90",
		X"32",X"53",X"B0",X"3E",X"91",X"32",X"55",X"B0",X"3E",X"17",X"32",X"45",X"B0",X"01",X"00",X"20",
		X"0D",X"20",X"FD",X"10",X"FB",X"3A",X"53",X"B0",X"3C",X"3C",X"FE",X"98",X"28",X"0E",X"32",X"53",
		X"B0",X"3A",X"55",X"B0",X"3C",X"3C",X"32",X"55",X"B0",X"C3",X"2D",X"31",X"3E",X"FF",X"32",X"53",
		X"B0",X"32",X"55",X"B0",X"3E",X"96",X"32",X"51",X"B4",X"3E",X"BC",X"32",X"50",X"B0",X"3E",X"02",
		X"32",X"50",X"B4",X"CD",X"50",X"46",X"DD",X"21",X"41",X"B4",X"06",X"05",X"DD",X"34",X"00",X"DD",
		X"23",X"DD",X"23",X"10",X"F7",X"01",X"00",X"0C",X"0D",X"20",X"FD",X"10",X"FB",X"3A",X"45",X"B0",
		X"FE",X"FF",X"28",X"06",X"06",X"17",X"78",X"32",X"45",X"B0",X"CD",X"50",X"46",X"3A",X"41",X"B4",
		X"FE",X"E8",X"CC",X"AD",X"31",X"FE",X"D8",X"CC",X"B3",X"31",X"FE",X"C8",X"CC",X"B9",X"31",X"FE",
		X"B8",X"CC",X"BF",X"31",X"FE",X"F4",X"CA",X"C5",X"31",X"C3",X"66",X"31",X"C9",X"3E",X"FF",X"32",
		X"43",X"B0",X"C9",X"3E",X"FF",X"32",X"45",X"B0",X"C9",X"3E",X"FF",X"32",X"47",X"B0",X"C9",X"3E",
		X"FF",X"32",X"49",X"B0",X"C9",X"06",X"08",X"C5",X"CD",X"1D",X"38",X"3A",X"51",X"B4",X"C6",X"08",
		X"32",X"51",X"B4",X"01",X"00",X"18",X"0D",X"20",X"FD",X"10",X"FB",X"C1",X"10",X"E9",X"06",X"40",
		X"C5",X"01",X"00",X"10",X"0D",X"20",X"FD",X"10",X"FB",X"CD",X"50",X"46",X"C1",X"10",X"F1",X"C9",
		X"BC",X"11",X"BC",X"FF",X"BC",X"FF",X"BC",X"FF",X"BC",X"FF",X"8C",X"F0",X"8C",X"00",X"82",X"10",
		X"90",X"20",X"90",X"30",X"10",X"15",X"0C",X"13",X"09",X"0E",X"07",X"FF",X"0E",X"0F",X"17",X"FF",
		X"10",X"0C",X"01",X"19",X"05",X"12",X"20",X"20",X"FF",X"00",X"31",X"40",X"A0",X"3E",X"00",X"32",
		X"F4",X"A8",X"3E",X"00",X"CD",X"D4",X"49",X"3E",X"00",X"32",X"F3",X"A8",X"CD",X"3C",X"4A",X"3E",
		X"00",X"32",X"F0",X"A8",X"32",X"F6",X"A8",X"32",X"F7",X"A8",X"3E",X"00",X"32",X"A9",X"A8",X"3E",
		X"30",X"32",X"C5",X"A8",X"32",X"C6",X"A8",X"21",X"2A",X"36",X"11",X"80",X"B0",X"01",X"4F",X"00",
		X"ED",X"B0",X"21",X"70",X"B0",X"11",X"71",X"B0",X"36",X"20",X"01",X"0F",X"00",X"ED",X"B0",X"21",
		X"7A",X"36",X"11",X"6C",X"A8",X"01",X"06",X"00",X"ED",X"B0",X"CD",X"BE",X"36",X"3E",X"00",X"32",
		X"02",X"C3",X"32",X"F3",X"A8",X"CD",X"E7",X"4C",X"CD",X"27",X"40",X"CD",X"29",X"4C",X"CD",X"D1",
		X"36",X"CD",X"97",X"49",X"3E",X"00",X"32",X"F4",X"A8",X"CD",X"44",X"4C",X"CD",X"F3",X"4E",X"32",
		X"C1",X"A8",X"FE",X"01",X"CA",X"89",X"34",X"C3",X"9A",X"32",X"3A",X"CE",X"A8",X"32",X"E0",X"A8",
		X"32",X"E8",X"A8",X"3E",X"00",X"32",X"E2",X"A8",X"32",X"EA",X"A8",X"32",X"E3",X"A8",X"32",X"EB",
		X"A8",X"32",X"E4",X"A8",X"32",X"EC",X"A8",X"3A",X"C2",X"A8",X"32",X"E1",X"A8",X"32",X"E9",X"A8",
		X"21",X"60",X"A8",X"11",X"61",X"A8",X"36",X"20",X"21",X"60",X"A8",X"11",X"61",X"A8",X"01",X"0B",
		X"00",X"ED",X"B0",X"3E",X"30",X"32",X"65",X"A8",X"32",X"6B",X"A8",X"C3",X"DE",X"32",X"3A",X"E4",
		X"A8",X"FE",X"FF",X"CA",X"1E",X"33",X"3E",X"01",X"32",X"9A",X"A8",X"3A",X"E0",X"A8",X"32",X"CF",
		X"A8",X"3A",X"E1",X"A8",X"32",X"9B",X"A8",X"3A",X"E2",X"A8",X"32",X"C0",X"A8",X"3A",X"E3",X"A8",
		X"32",X"9E",X"A8",X"CD",X"6B",X"33",X"3A",X"CF",X"A8",X"32",X"E0",X"A8",X"3A",X"9B",X"A8",X"32",
		X"E1",X"A8",X"3A",X"C0",X"A8",X"32",X"E2",X"A8",X"3A",X"9E",X"A8",X"32",X"E3",X"A8",X"3A",X"EC",
		X"A8",X"FE",X"FF",X"20",X"0B",X"3A",X"E4",X"A8",X"FE",X"FF",X"C2",X"DE",X"32",X"C3",X"6D",X"32",
		X"3E",X"02",X"32",X"9A",X"A8",X"3A",X"E8",X"A8",X"32",X"CF",X"A8",X"3A",X"E9",X"A8",X"32",X"9B",
		X"A8",X"3A",X"EA",X"A8",X"32",X"C0",X"A8",X"3A",X"EB",X"A8",X"32",X"9E",X"A8",X"CD",X"6B",X"33",
		X"3A",X"CF",X"A8",X"32",X"E8",X"A8",X"3A",X"9B",X"A8",X"32",X"E9",X"A8",X"3A",X"C0",X"A8",X"32",
		X"EA",X"A8",X"3A",X"9E",X"A8",X"32",X"EB",X"A8",X"C3",X"DE",X"32",X"CD",X"FC",X"4F",X"CD",X"E7",
		X"4C",X"CD",X"81",X"36",X"3E",X"00",X"32",X"F4",X"A8",X"CD",X"E7",X"4C",X"CD",X"B7",X"35",X"FE",
		X"FF",X"CA",X"F0",X"33",X"32",X"C0",X"A8",X"C5",X"3A",X"CF",X"A8",X"3C",X"32",X"CF",X"A8",X"CD",
		X"CA",X"4D",X"C1",X"78",X"FE",X"01",X"20",X"06",X"CD",X"4D",X"39",X"C3",X"B5",X"33",X"FE",X"03",
		X"20",X"06",X"CD",X"7F",X"39",X"C3",X"B5",X"33",X"FE",X"00",X"20",X"06",X"CD",X"E3",X"39",X"C3",
		X"B5",X"33",X"CD",X"B1",X"39",X"CD",X"09",X"41",X"CD",X"98",X"4E",X"CD",X"AF",X"4E",X"21",X"B1",
		X"35",X"11",X"4E",X"A6",X"06",X"21",X"CD",X"DB",X"36",X"21",X"81",X"34",X"11",X"6C",X"A6",X"06",
		X"21",X"CD",X"DB",X"36",X"3A",X"9A",X"A8",X"C6",X"B0",X"32",X"AC",X"A5",X"3E",X"05",X"01",X"00",
		X"00",X"0D",X"20",X"FD",X"05",X"20",X"FA",X"3D",X"20",X"F7",X"CD",X"D6",X"4E",X"C3",X"74",X"33",
		X"3E",X"00",X"CD",X"D4",X"49",X"CD",X"19",X"4A",X"3E",X"01",X"32",X"81",X"A8",X"2A",X"50",X"B0",
		X"26",X"90",X"22",X"52",X"B0",X"24",X"22",X"54",X"B0",X"2A",X"50",X"B4",X"7C",X"D6",X"08",X"67",
		X"22",X"52",X"B4",X"7C",X"C6",X"10",X"67",X"22",X"54",X"B4",X"3E",X"04",X"32",X"1B",X"A8",X"3E",
		X"FF",X"32",X"51",X"B0",X"32",X"50",X"B0",X"CD",X"03",X"36",X"3A",X"1B",X"A8",X"FE",X"00",X"20",
		X"F6",X"01",X"00",X"09",X"C5",X"CD",X"03",X"36",X"C1",X"0D",X"20",X"F8",X"10",X"F6",X"3E",X"00",
		X"32",X"81",X"A8",X"3E",X"03",X"32",X"93",X"A8",X"3A",X"9B",X"A8",X"3D",X"FE",X"FF",X"20",X"2D",
		X"CD",X"12",X"52",X"FE",X"FF",X"20",X"10",X"21",X"E4",X"A8",X"3A",X"9A",X"A8",X"FE",X"01",X"28",
		X"03",X"21",X"EC",X"A8",X"36",X"FF",X"C9",X"DD",X"21",X"E0",X"A8",X"3A",X"9A",X"A8",X"FE",X"01",
		X"28",X"04",X"DD",X"21",X"E8",X"A8",X"3A",X"C2",X"A8",X"DD",X"77",X"01",X"C9",X"32",X"9B",X"A8",
		X"C9",X"10",X"0C",X"01",X"19",X"05",X"12",X"20",X"FF",X"3A",X"CE",X"A8",X"32",X"CF",X"A8",X"3E",
		X"00",X"32",X"C0",X"A8",X"32",X"9E",X"A8",X"3A",X"C2",X"A8",X"32",X"9B",X"A8",X"21",X"60",X"A8",
		X"11",X"61",X"A8",X"36",X"20",X"21",X"60",X"A8",X"11",X"61",X"A8",X"01",X"0B",X"00",X"ED",X"B0",
		X"3E",X"30",X"32",X"65",X"A8",X"32",X"6B",X"A8",X"3E",X"03",X"32",X"93",X"A8",X"C3",X"C0",X"34",
		X"3E",X"00",X"32",X"02",X"C3",X"32",X"F3",X"A8",X"3E",X"01",X"32",X"9A",X"A8",X"CD",X"E7",X"4C",
		X"CD",X"81",X"36",X"CD",X"E7",X"4C",X"CD",X"B7",X"35",X"FE",X"FF",X"CA",X"37",X"35",X"32",X"C0",
		X"A8",X"C5",X"3A",X"CF",X"A8",X"3C",X"32",X"CF",X"A8",X"CD",X"CA",X"4D",X"C1",X"78",X"FE",X"01",
		X"20",X"06",X"CD",X"4D",X"39",X"C3",X"0F",X"35",X"FE",X"03",X"20",X"06",X"CD",X"7F",X"39",X"C3",
		X"0F",X"35",X"FE",X"00",X"20",X"06",X"CD",X"E3",X"39",X"C3",X"0F",X"35",X"CD",X"B1",X"39",X"CD",
		X"09",X"41",X"CD",X"98",X"4E",X"CD",X"AF",X"4E",X"21",X"B1",X"35",X"11",X"4D",X"A6",X"06",X"21",
		X"CD",X"DB",X"36",X"3E",X"05",X"01",X"00",X"00",X"0D",X"20",X"FD",X"05",X"20",X"FA",X"3D",X"20",
		X"F7",X"CD",X"D6",X"4E",X"C3",X"D3",X"34",X"3E",X"00",X"CD",X"D4",X"49",X"CD",X"19",X"4A",X"3E",
		X"01",X"32",X"81",X"A8",X"2A",X"50",X"B0",X"26",X"90",X"22",X"52",X"B0",X"24",X"22",X"54",X"B0",
		X"2A",X"50",X"B4",X"7C",X"D6",X"08",X"67",X"22",X"52",X"B4",X"7C",X"C6",X"10",X"67",X"22",X"54",
		X"B4",X"3E",X"04",X"32",X"1B",X"A8",X"3E",X"FF",X"32",X"51",X"B0",X"32",X"50",X"B0",X"CD",X"03",
		X"36",X"3A",X"1B",X"A8",X"FE",X"00",X"20",X"F6",X"01",X"00",X"09",X"C5",X"CD",X"03",X"36",X"C1",
		X"0D",X"20",X"F8",X"10",X"F6",X"3E",X"00",X"32",X"81",X"A8",X"3E",X"03",X"32",X"93",X"A8",X"3A",
		X"9B",X"A8",X"3D",X"FE",X"FF",X"20",X"11",X"CD",X"12",X"52",X"FE",X"FF",X"CA",X"6D",X"32",X"3A",
		X"C2",X"A8",X"32",X"9B",X"A8",X"C3",X"C0",X"34",X"32",X"9B",X"A8",X"CD",X"FC",X"4F",X"C3",X"C0",
		X"34",X"12",X"05",X"01",X"04",X"19",X"FF",X"CD",X"9E",X"54",X"CD",X"EB",X"47",X"CD",X"7D",X"46",
		X"CD",X"DB",X"54",X"CD",X"BE",X"3E",X"CD",X"03",X"44",X"CD",X"03",X"44",X"CD",X"03",X"44",X"CD",
		X"A5",X"42",X"CD",X"34",X"42",X"3A",X"8C",X"A8",X"FE",X"FF",X"C8",X"3A",X"8E",X"A8",X"E6",X"FC",
		X"FE",X"50",X"20",X"0D",X"3A",X"8E",X"A8",X"E6",X"03",X"47",X"C6",X"B0",X"6F",X"26",X"A8",X"7E",
		X"C9",X"21",X"92",X"A8",X"35",X"20",X"C0",X"3E",X"08",X"77",X"CD",X"E6",X"53",X"CD",X"AA",X"43",
		X"C3",X"B7",X"35",X"CD",X"9E",X"54",X"CD",X"DB",X"54",X"CD",X"BE",X"3E",X"CD",X"03",X"44",X"CD",
		X"03",X"44",X"CD",X"03",X"44",X"CD",X"A5",X"42",X"CD",X"34",X"42",X"21",X"92",X"A8",X"35",X"C0",
		X"3E",X"08",X"77",X"CD",X"E6",X"53",X"CD",X"AA",X"43",X"C9",X"31",X"2E",X"20",X"01",X"01",X"01",
		X"20",X"20",X"32",X"35",X"30",X"30",X"30",X"20",X"20",X"20",X"32",X"2E",X"20",X"02",X"02",X"02",
		X"20",X"20",X"32",X"30",X"30",X"30",X"30",X"20",X"20",X"20",X"33",X"2E",X"20",X"03",X"03",X"03",
		X"20",X"20",X"31",X"35",X"30",X"30",X"30",X"20",X"20",X"20",X"34",X"2E",X"20",X"04",X"04",X"04",
		X"20",X"20",X"31",X"30",X"30",X"30",X"30",X"20",X"20",X"20",X"35",X"2E",X"20",X"05",X"05",X"05",
		X"20",X"20",X"20",X"35",X"30",X"30",X"30",X"20",X"20",X"20",X"20",X"32",X"35",X"30",X"30",X"30",
		X"30",X"CD",X"9A",X"4C",X"CD",X"29",X"4C",X"CD",X"06",X"30",X"CD",X"09",X"41",X"3A",X"18",X"A8",
		X"E6",X"1F",X"6F",X"26",X"00",X"11",X"9E",X"36",X"19",X"7E",X"32",X"87",X"A8",X"C9",X"04",X"05",
		X"05",X"06",X"06",X"06",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",
		X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"21",X"60",
		X"A8",X"11",X"61",X"A8",X"01",X"0B",X"00",X"ED",X"B0",X"3E",X"30",X"32",X"65",X"A8",X"32",X"6B",
		X"A8",X"CD",X"EA",X"3D",X"CD",X"4A",X"3E",X"CD",X"44",X"4C",X"C9",X"EB",X"E5",X"DD",X"E1",X"C5",
		X"01",X"00",X"FC",X"09",X"C1",X"E5",X"FD",X"E1",X"EB",X"7E",X"F6",X"80",X"DD",X"77",X"00",X"78",
		X"FD",X"77",X"00",X"11",X"E0",X"FF",X"DD",X"19",X"FD",X"19",X"23",X"7E",X"FE",X"FF",X"20",X"E9",
		X"C9",X"CD",X"23",X"4A",X"21",X"02",X"A9",X"22",X"D0",X"A8",X"21",X"82",X"AC",X"22",X"D2",X"A8",
		X"C9",X"21",X"43",X"A4",X"22",X"D4",X"A8",X"21",X"43",X"A0",X"22",X"D6",X"A8",X"06",X"1C",X"C5",
		X"2A",X"D4",X"A8",X"E5",X"D1",X"1B",X"01",X"1C",X"00",X"ED",X"B0",X"2A",X"D6",X"A8",X"E5",X"D1",
		X"1B",X"01",X"1C",X"00",X"ED",X"B0",X"11",X"20",X"00",X"2A",X"D4",X"A8",X"19",X"22",X"D4",X"A8",
		X"2A",X"D6",X"A8",X"19",X"22",X"D6",X"A8",X"C1",X"10",X"D5",X"06",X"1C",X"DD",X"2A",X"D0",X"A8",
		X"FD",X"2A",X"D2",X"A8",X"21",X"5D",X"A4",X"11",X"5D",X"A0",X"C5",X"DD",X"7E",X"00",X"77",X"FD",
		X"7E",X"00",X"12",X"01",X"20",X"00",X"DD",X"09",X"FD",X"09",X"09",X"E5",X"EB",X"09",X"EB",X"E1",
		X"C1",X"10",X"E7",X"21",X"D0",X"A8",X"34",X"23",X"23",X"34",X"C9",X"CD",X"23",X"4A",X"21",X"1D",
		X"A9",X"22",X"D0",X"A8",X"21",X"9D",X"AC",X"22",X"D2",X"A8",X"C9",X"21",X"5D",X"A4",X"22",X"D4",
		X"A8",X"21",X"5D",X"A0",X"22",X"D6",X"A8",X"06",X"1C",X"C5",X"2A",X"D4",X"A8",X"E5",X"D1",X"2B",
		X"01",X"1B",X"00",X"ED",X"B8",X"2A",X"D6",X"A8",X"E5",X"D1",X"2B",X"01",X"1B",X"00",X"ED",X"B8",
		X"11",X"20",X"00",X"2A",X"D4",X"A8",X"19",X"22",X"D4",X"A8",X"2A",X"D6",X"A8",X"19",X"22",X"D6",
		X"A8",X"C1",X"10",X"D5",X"06",X"1C",X"DD",X"2A",X"D0",X"A8",X"FD",X"2A",X"D2",X"A8",X"21",X"42",
		X"A4",X"11",X"42",X"A0",X"C5",X"DD",X"7E",X"00",X"77",X"FD",X"7E",X"00",X"12",X"01",X"20",X"00",
		X"DD",X"09",X"FD",X"09",X"09",X"E5",X"EB",X"09",X"EB",X"E1",X"C1",X"10",X"E7",X"21",X"D0",X"A8",
		X"35",X"23",X"23",X"35",X"C9",X"CD",X"23",X"4A",X"21",X"82",X"A7",X"22",X"D0",X"A8",X"21",X"A2",
		X"A7",X"22",X"D2",X"A8",X"21",X"82",X"A3",X"22",X"D4",X"A8",X"21",X"A2",X"A3",X"22",X"D6",X"A8",
		X"21",X"62",X"AC",X"22",X"D8",X"A8",X"21",X"E2",X"AF",X"22",X"DA",X"A8",X"C9",X"21",X"82",X"A7",
		X"22",X"D0",X"A8",X"21",X"A2",X"A7",X"22",X"D2",X"A8",X"21",X"82",X"A3",X"22",X"D4",X"A8",X"21",
		X"A2",X"A3",X"22",X"D6",X"A8",X"3E",X"1B",X"32",X"DC",X"A8",X"2A",X"D0",X"A8",X"EB",X"2A",X"D2",
		X"A8",X"EB",X"01",X"1C",X"00",X"ED",X"B0",X"2A",X"D4",X"A8",X"EB",X"2A",X"D6",X"A8",X"EB",X"01",
		X"1C",X"00",X"ED",X"B0",X"11",X"E0",X"FF",X"2A",X"D0",X"A8",X"19",X"22",X"D0",X"A8",X"2A",X"D2",
		X"A8",X"19",X"22",X"D2",X"A8",X"2A",X"D4",X"A8",X"19",X"22",X"D4",X"A8",X"2A",X"D6",X"A8",X"19",
		X"22",X"D6",X"A8",X"21",X"DC",X"A8",X"35",X"20",X"C1",X"2A",X"D8",X"A8",X"11",X"42",X"A4",X"01",
		X"1C",X"00",X"ED",X"B0",X"2A",X"DA",X"A8",X"11",X"42",X"A0",X"01",X"1C",X"00",X"ED",X"B0",X"11",
		X"E0",X"FF",X"2A",X"D8",X"A8",X"19",X"22",X"D8",X"A8",X"2A",X"DA",X"A8",X"19",X"22",X"DA",X"A8",
		X"C9",X"CD",X"23",X"4A",X"21",X"62",X"A4",X"22",X"D0",X"A8",X"21",X"42",X"A4",X"22",X"D2",X"A8",
		X"21",X"62",X"A0",X"22",X"D4",X"A8",X"21",X"42",X"A0",X"22",X"D6",X"A8",X"21",X"02",X"A9",X"22",
		X"D8",X"A8",X"21",X"82",X"AC",X"22",X"DA",X"A8",X"C9",X"21",X"62",X"A4",X"22",X"D0",X"A8",X"21",
		X"42",X"A4",X"22",X"D2",X"A8",X"21",X"62",X"A0",X"22",X"D4",X"A8",X"21",X"42",X"A0",X"22",X"D6",
		X"A8",X"3E",X"1B",X"32",X"DC",X"A8",X"2A",X"D0",X"A8",X"EB",X"2A",X"D2",X"A8",X"EB",X"01",X"1C",
		X"00",X"ED",X"B0",X"2A",X"D4",X"A8",X"EB",X"2A",X"D6",X"A8",X"EB",X"01",X"1C",X"00",X"ED",X"B0",
		X"11",X"20",X"00",X"2A",X"D0",X"A8",X"19",X"22",X"D0",X"A8",X"2A",X"D2",X"A8",X"19",X"22",X"D2",
		X"A8",X"2A",X"D4",X"A8",X"19",X"22",X"D4",X"A8",X"2A",X"D6",X"A8",X"19",X"22",X"D6",X"A8",X"21",
		X"DC",X"A8",X"35",X"20",X"C1",X"2A",X"D8",X"A8",X"11",X"A2",X"A7",X"01",X"1C",X"00",X"ED",X"B0",
		X"2A",X"DA",X"A8",X"11",X"A2",X"A3",X"01",X"1C",X"00",X"ED",X"B0",X"11",X"20",X"00",X"2A",X"D8",
		X"A8",X"19",X"22",X"D8",X"A8",X"2A",X"DA",X"A8",X"19",X"22",X"DA",X"A8",X"C9",X"CD",X"50",X"41",
		X"2A",X"50",X"B0",X"E5",X"2A",X"50",X"B4",X"E5",X"CD",X"29",X"4C",X"CD",X"F5",X"37",X"06",X"1C",
		X"C5",X"CD",X"1D",X"38",X"01",X"00",X"08",X"0D",X"20",X"FD",X"10",X"FB",X"C1",X"10",X"F1",X"E1",
		X"26",X"D0",X"22",X"50",X"B4",X"E1",X"22",X"50",X"B0",X"3E",X"01",X"32",X"09",X"A8",X"C9",X"CD",
		X"50",X"41",X"2A",X"50",X"B0",X"E5",X"2A",X"50",X"B4",X"E5",X"CD",X"29",X"4C",X"CD",X"A1",X"38",
		X"06",X"1C",X"C5",X"CD",X"C9",X"38",X"01",X"00",X"08",X"0D",X"20",X"FD",X"10",X"FB",X"C1",X"10",
		X"F1",X"E1",X"26",X"10",X"22",X"50",X"B4",X"E1",X"22",X"50",X"B0",X"3E",X"03",X"32",X"09",X"A8",
		X"C9",X"CD",X"50",X"41",X"2A",X"50",X"B0",X"E5",X"2A",X"50",X"B4",X"E5",X"CD",X"29",X"4C",X"CD",
		X"01",X"37",X"06",X"1C",X"C5",X"CD",X"11",X"37",X"01",X"00",X"08",X"0D",X"20",X"FD",X"10",X"FB",
		X"C1",X"10",X"F1",X"E1",X"22",X"50",X"B4",X"E1",X"2E",X"D0",X"22",X"50",X"B0",X"3E",X"02",X"32",
		X"09",X"A8",X"C9",X"CD",X"50",X"41",X"2A",X"50",X"B0",X"E5",X"2A",X"50",X"B4",X"E5",X"CD",X"29",
		X"4C",X"CD",X"7B",X"37",X"06",X"1C",X"C5",X"CD",X"8B",X"37",X"01",X"00",X"08",X"0D",X"20",X"FD",
		X"10",X"FB",X"C1",X"10",X"F1",X"E1",X"22",X"50",X"B4",X"E1",X"2E",X"19",X"22",X"50",X"B0",X"3E",
		X"00",X"32",X"09",X"A8",X"C9",X"00",X"00",X"01",X"FF",X"01",X"4B",X"00",X"86",X"01",X"2D",X"09",
		X"12",X"08",X"8B",X"00",X"00",X"08",X"08",X"09",X"0A",X"01",X"21",X"11",X"03",X"10",X"11",X"00",
		X"FF",X"00",X"19",X"04",X"FF",X"04",X"BF",X"00",X"0E",X"01",X"52",X"00",X"4C",X"01",X"95",X"00",
		X"0C",X"04",X"66",X"00",X"21",X"04",X"D6",X"00",X"1A",X"08",X"47",X"00",X"00",X"08",X"18",X"00",
		X"05",X"02",X"FF",X"02",X"91",X"04",X"62",X"00",X"37",X"02",X"59",X"00",X"FF",X"00",X"99",X"01",
		X"25",X"09",X"00",X"08",X"3D",X"09",X"00",X"01",X"FF",X"01",X"75",X"00",X"2F",X"04",X"5B",X"00",
		X"FF",X"00",X"D6",X"08",X"2C",X"00",X"0D",X"02",X"41",X"00",X"0F",X"10",X"13",X"00",X"FF",X"00",
		X"7C",X"04",X"6A",X"00",X"1E",X"01",X"51",X"00",X"FF",X"00",X"48",X"08",X"19",X"09",X"01",X"01",
		X"26",X"09",X"01",X"08",X"55",X"09",X"08",X"01",X"FF",X"01",X"78",X"00",X"5A",X"04",X"3A",X"00",
		X"7D",X"01",X"FF",X"01",X"1B",X"00",X"B1",X"02",X"2E",X"00",X"1B",X"10",X"13",X"00",X"EC",X"08",
		X"6B",X"00",X"1D",X"01",X"75",X"00",X"1E",X"08",X"6B",X"00",X"2C",X"02",X"75",X"0A",X"03",X"08",
		X"5A",X"0A",X"00",X"02",X"A1",X"0A",X"34",X"08",X"1D",X"00",X"06",X"10",X"0F",X"00",X"F5",X"04",
		X"FF",X"04",X"FF",X"04",X"6C",X"3E",X"30",X"32",X"1D",X"A8",X"32",X"1E",X"A8",X"32",X"1F",X"A8",
		X"3A",X"CE",X"A8",X"32",X"E0",X"A8",X"32",X"E8",X"A8",X"3E",X"00",X"32",X"E2",X"A8",X"32",X"EA",
		X"A8",X"32",X"E3",X"A8",X"32",X"EB",X"A8",X"32",X"E4",X"A8",X"32",X"EC",X"A8",X"3A",X"C2",X"A8",
		X"32",X"E1",X"A8",X"32",X"E9",X"A8",X"3E",X"01",X"32",X"9A",X"A8",X"3A",X"E0",X"A8",X"32",X"CF",
		X"A8",X"3A",X"E1",X"A8",X"3E",X"00",X"32",X"9B",X"A8",X"3E",X"C0",X"32",X"85",X"A8",X"3A",X"E2",
		X"A8",X"32",X"C0",X"A8",X"3A",X"E3",X"A8",X"32",X"9E",X"A8",X"CD",X"E7",X"4C",X"3E",X"02",X"32",
		X"C0",X"A8",X"CD",X"81",X"36",X"21",X"15",X"3A",X"22",X"F8",X"A8",X"7E",X"32",X"FA",X"A8",X"23",
		X"7E",X"23",X"32",X"FB",X"A8",X"3E",X"00",X"32",X"FC",X"A8",X"3E",X"03",X"32",X"93",X"A8",X"CD",
		X"9E",X"54",X"CD",X"A7",X"3B",X"CD",X"7D",X"46",X"CD",X"DB",X"54",X"CD",X"BE",X"3E",X"CD",X"03",
		X"44",X"CD",X"03",X"44",X"CD",X"03",X"44",X"CD",X"A5",X"42",X"CD",X"34",X"42",X"3A",X"FC",X"A8",
		X"FE",X"C0",X"C8",X"3A",X"A9",X"A8",X"FE",X"00",X"C0",X"3A",X"8C",X"A8",X"FE",X"FF",X"C8",X"3A",
		X"8E",X"A8",X"E6",X"FC",X"FE",X"50",X"20",X"0D",X"3A",X"8E",X"A8",X"E6",X"03",X"47",X"C6",X"B0",
		X"6F",X"26",X"A8",X"7E",X"C9",X"21",X"92",X"A8",X"35",X"20",X"B4",X"3E",X"08",X"77",X"CD",X"E6",
		X"53",X"CD",X"AA",X"43",X"C3",X"4F",X"3B",X"21",X"0A",X"A8",X"06",X"06",X"36",X"00",X"23",X"10",
		X"FB",X"3A",X"FA",X"A8",X"21",X"0F",X"A8",X"06",X"05",X"CB",X"3F",X"CB",X"16",X"2B",X"10",X"F9",
		X"3A",X"FB",X"A8",X"3D",X"32",X"FB",X"A8",X"FE",X"00",X"C0",X"2A",X"F8",X"A8",X"7E",X"32",X"FA",
		X"A8",X"23",X"7E",X"32",X"FB",X"A8",X"23",X"22",X"F8",X"A8",X"3A",X"FC",X"A8",X"3C",X"32",X"FC",
		X"A8",X"C9",X"E5",X"D5",X"C5",X"DD",X"E5",X"FD",X"E5",X"47",X"3A",X"F4",X"A8",X"FE",X"00",X"20",
		X"17",X"3A",X"9A",X"A8",X"DD",X"21",X"64",X"A8",X"FE",X"01",X"28",X"04",X"DD",X"21",X"6A",X"A8",
		X"CD",X"10",X"3C",X"10",X"FB",X"CD",X"4A",X"3E",X"FD",X"E1",X"DD",X"E1",X"C1",X"D1",X"E1",X"C9",
		X"DD",X"E5",X"DD",X"7E",X"00",X"FE",X"20",X"20",X"02",X"3E",X"30",X"3C",X"FE",X"3A",X"28",X"09",
		X"DD",X"77",X"00",X"DD",X"E1",X"CD",X"33",X"3C",X"C9",X"3E",X"30",X"DD",X"77",X"00",X"DD",X"2B",
		X"C3",X"12",X"3C",X"E5",X"D5",X"C5",X"DD",X"E5",X"E1",X"11",X"69",X"3C",X"3A",X"CD",X"A8",X"FE",
		X"00",X"28",X"03",X"11",X"6F",X"3C",X"2B",X"2B",X"2B",X"06",X"04",X"1A",X"BE",X"28",X"04",X"C1",
		X"D1",X"E1",X"C9",X"13",X"23",X"10",X"F4",X"3A",X"9B",X"A8",X"FE",X"05",X"28",X"07",X"3C",X"32",
		X"9B",X"A8",X"CD",X"BA",X"3C",X"C1",X"D1",X"E1",X"C9",X"35",X"30",X"30",X"30",X"30",X"30",X"30",
		X"30",X"30",X"30",X"30",X"30",X"30",X"3A",X"00",X"C2",X"E6",X"10",X"20",X"05",X"3E",X"0F",X"32",
		X"93",X"A8",X"DD",X"21",X"FE",X"A4",X"FD",X"21",X"FE",X"A0",X"11",X"E0",X"FF",X"3A",X"93",X"A8",
		X"47",X"0E",X"00",X"78",X"FE",X"00",X"28",X"0D",X"3E",X"88",X"DD",X"77",X"00",X"3E",X"10",X"FD",
		X"77",X"00",X"05",X"18",X"0A",X"3E",X"00",X"DD",X"77",X"00",X"3E",X"10",X"FD",X"77",X"00",X"DD",
		X"19",X"FD",X"19",X"0C",X"79",X"FE",X"05",X"20",X"DA",X"C9",X"DD",X"21",X"BF",X"A7",X"FD",X"21",
		X"BF",X"A3",X"11",X"E0",X"FF",X"3A",X"9B",X"A8",X"47",X"0E",X"00",X"78",X"FE",X"00",X"28",X"0D",
		X"3E",X"84",X"DD",X"77",X"00",X"3E",X"14",X"FD",X"77",X"00",X"05",X"18",X"0A",X"3E",X"00",X"DD",
		X"77",X"00",X"3E",X"14",X"FD",X"77",X"00",X"DD",X"19",X"FD",X"19",X"0C",X"79",X"FE",X"05",X"20",
		X"DA",X"C9",X"C6",X"20",X"6F",X"CB",X"25",X"26",X"B0",X"7E",X"57",X"26",X"B4",X"2C",X"7E",X"5F",
		X"78",X"C6",X"20",X"47",X"68",X"CB",X"25",X"26",X"B0",X"7E",X"47",X"26",X"B4",X"2C",X"7E",X"4F",
		X"7A",X"D6",X"04",X"B8",X"30",X"15",X"7A",X"C6",X"04",X"B8",X"38",X"0F",X"7B",X"D6",X"04",X"B9",
		X"30",X"09",X"7B",X"C6",X"04",X"B9",X"38",X"03",X"3E",X"00",X"C9",X"7A",X"D6",X"06",X"B8",X"30",
		X"15",X"7A",X"C6",X"06",X"B8",X"38",X"0F",X"7B",X"D6",X"06",X"B9",X"30",X"09",X"7B",X"C6",X"06",
		X"B9",X"38",X"03",X"3E",X"01",X"C9",X"3E",X"FF",X"C9",X"10",X"10",X"10",X"10",X"1C",X"1C",X"1C",
		X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"E5",X"C5",X"D5",X"DD",X"E5",X"DD",X"21",
		X"49",X"3D",X"21",X"1E",X"A3",X"06",X"10",X"11",X"E0",X"FF",X"DD",X"7E",X"00",X"77",X"19",X"DD",
		X"23",X"10",X"F7",X"3A",X"85",X"A8",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"DD",X"21",
		X"1E",X"A7",X"4F",X"06",X"10",X"11",X"E0",X"FF",X"79",X"FE",X"00",X"28",X"0C",X"3E",X"80",X"DD",
		X"77",X"00",X"DD",X"19",X"05",X"0D",X"C3",X"88",X"3D",X"3A",X"85",X"A8",X"E6",X"0F",X"CB",X"3F",
		X"CB",X"3F",X"FE",X"00",X"28",X"10",X"EE",X"03",X"C6",X"80",X"FE",X"84",X"20",X"02",X"3E",X"85",
		X"DD",X"77",X"00",X"DD",X"19",X"05",X"78",X"FE",X"00",X"28",X"0F",X"FE",X"FF",X"28",X"0B",X"3E",
		X"85",X"DD",X"77",X"00",X"DD",X"19",X"05",X"C3",X"B6",X"3D",X"06",X"02",X"3A",X"85",X"A8",X"E6",
		X"E0",X"FE",X"E0",X"28",X"0B",X"06",X"01",X"3A",X"85",X"A8",X"E6",X"E0",X"20",X"02",X"06",X"00",
		X"78",X"32",X"86",X"A8",X"DD",X"E1",X"D1",X"C1",X"E1",X"C9",X"DD",X"21",X"A0",X"A7",X"FD",X"21",
		X"A0",X"A3",X"21",X"12",X"3E",X"11",X"2E",X"3E",X"06",X"1C",X"7E",X"F6",X"80",X"DD",X"77",X"00",
		X"1A",X"FD",X"77",X"00",X"D5",X"11",X"E0",X"FF",X"DD",X"19",X"FD",X"19",X"D1",X"13",X"23",X"10",
		X"E9",X"C9",X"20",X"10",X"0C",X"01",X"19",X"05",X"12",X"31",X"20",X"20",X"08",X"09",X"20",X"13",
		X"03",X"0F",X"12",X"05",X"20",X"20",X"10",X"0C",X"01",X"19",X"05",X"12",X"32",X"20",X"2C",X"2C",
		X"2C",X"2C",X"2C",X"2C",X"2C",X"2C",X"2C",X"2C",X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"24",
		X"2C",X"2C",X"2C",X"2C",X"2C",X"2C",X"2C",X"2C",X"2C",X"2C",X"DD",X"21",X"81",X"A7",X"FD",X"21",
		X"81",X"A3",X"21",X"60",X"A8",X"06",X"06",X"11",X"E0",X"FF",X"7E",X"F6",X"80",X"DD",X"77",X"00",
		X"3A",X"82",X"A8",X"FD",X"77",X"00",X"DD",X"19",X"FD",X"19",X"23",X"10",X"ED",X"DD",X"21",X"21",
		X"A5",X"FD",X"21",X"21",X"A1",X"21",X"66",X"A8",X"06",X"06",X"7E",X"F6",X"80",X"DD",X"77",X"00",
		X"3A",X"83",X"A8",X"FD",X"77",X"00",X"DD",X"19",X"FD",X"19",X"23",X"10",X"ED",X"DD",X"21",X"41",
		X"A6",X"FD",X"21",X"41",X"A2",X"21",X"6C",X"A8",X"06",X"06",X"7E",X"F6",X"80",X"DD",X"77",X"00",
		X"3A",X"84",X"A8",X"FD",X"77",X"00",X"DD",X"19",X"FD",X"19",X"23",X"10",X"ED",X"C9",X"34",X"20",
		X"24",X"28",X"2C",X"34",X"30",X"30",X"34",X"2C",X"28",X"24",X"20",X"34",X"34",X"34",X"21",X"C9",
		X"A8",X"35",X"20",X"2B",X"3E",X"07",X"77",X"2B",X"35",X"20",X"24",X"3E",X"30",X"77",X"2B",X"35",
		X"20",X"1D",X"3E",X"08",X"77",X"3A",X"18",X"A8",X"3C",X"FE",X"20",X"20",X"02",X"3E",X"1F",X"32",
		X"18",X"A8",X"3A",X"87",X"A8",X"3C",X"FE",X"08",X"20",X"02",X"3E",X"07",X"32",X"87",X"A8",X"21",
		X"1C",X"A8",X"35",X"C0",X"3A",X"86",X"A8",X"FE",X"02",X"20",X"21",X"3A",X"00",X"A8",X"3C",X"32",
		X"00",X"A8",X"E6",X"07",X"6F",X"26",X"00",X"11",X"AE",X"3E",X"19",X"46",X"21",X"82",X"A8",X"3A",
		X"9A",X"A8",X"FE",X"01",X"28",X"03",X"21",X"83",X"A8",X"70",X"18",X"08",X"3E",X"34",X"32",X"82",
		X"A8",X"32",X"83",X"A8",X"CD",X"4A",X"3E",X"3E",X"40",X"32",X"1C",X"A8",X"3A",X"1B",X"A8",X"FE",
		X"00",X"20",X"07",X"3A",X"8F",X"A8",X"FE",X"00",X"28",X"23",X"3A",X"53",X"B0",X"3C",X"3C",X"FE",
		X"98",X"20",X"13",X"3E",X"FF",X"32",X"53",X"B0",X"32",X"55",X"B0",X"3E",X"00",X"32",X"1B",X"A8",
		X"32",X"8F",X"A8",X"C3",X"5D",X"3F",X"32",X"53",X"B0",X"3C",X"32",X"55",X"B0",X"21",X"8B",X"A8",
		X"7E",X"FE",X"00",X"28",X"10",X"3A",X"57",X"B0",X"3C",X"FE",X"A0",X"20",X"05",X"3E",X"00",X"77",
		X"3E",X"FF",X"32",X"57",X"B0",X"3A",X"8D",X"A8",X"FE",X"00",X"28",X"15",X"3A",X"59",X"B0",X"3D",
		X"FE",X"97",X"20",X"07",X"3E",X"00",X"32",X"8D",X"A8",X"3E",X"FF",X"32",X"59",X"B0",X"32",X"5B",
		X"B0",X"3A",X"96",X"A8",X"FE",X"00",X"28",X"12",X"3A",X"61",X"B0",X"3C",X"FE",X"A0",X"20",X"07",
		X"3E",X"00",X"32",X"96",X"A8",X"3E",X"FF",X"32",X"61",X"B0",X"3A",X"99",X"A8",X"FE",X"00",X"28",
		X"17",X"3D",X"28",X"0F",X"32",X"99",X"A8",X"3A",X"62",X"B4",X"EE",X"02",X"F6",X"80",X"32",X"62",
		X"B4",X"18",X"05",X"3E",X"FF",X"32",X"63",X"B0",X"3A",X"B4",X"A8",X"FE",X"00",X"28",X"41",X"E6",
		X"E0",X"20",X"0C",X"3A",X"B4",X"A8",X"CB",X"3F",X"E6",X"01",X"C6",X"0F",X"32",X"65",X"B0",X"3A",
		X"B4",X"A8",X"3D",X"32",X"B4",X"A8",X"20",X"28",X"3E",X"FF",X"32",X"65",X"B0",X"DD",X"21",X"20",
		X"A8",X"06",X"00",X"11",X"40",X"B4",X"DD",X"7E",X"00",X"FE",X"02",X"20",X"08",X"3E",X"02",X"12",
		X"3E",X"01",X"DD",X"77",X"00",X"13",X"13",X"D5",X"11",X"08",X"00",X"DD",X"19",X"D1",X"10",X"E6",
		X"21",X"B6",X"A8",X"34",X"20",X"10",X"3A",X"B6",X"A8",X"77",X"21",X"89",X"A8",X"34",X"7E",X"FE",
		X"21",X"20",X"03",X"3E",X"20",X"77",X"C9",X"DD",X"21",X"A0",X"A7",X"FD",X"21",X"A0",X"A3",X"CD",
		X"3A",X"40",X"DD",X"21",X"BE",X"A7",X"FD",X"21",X"BE",X"A3",X"11",X"E0",X"FF",X"DD",X"E5",X"FD",
		X"E5",X"3E",X"20",X"06",X"1C",X"DD",X"77",X"00",X"FD",X"77",X"00",X"DD",X"19",X"FD",X"19",X"10",
		X"F4",X"FD",X"E1",X"DD",X"E1",X"FD",X"23",X"DD",X"23",X"06",X"1C",X"DD",X"77",X"00",X"FD",X"77",
		X"00",X"DD",X"19",X"FD",X"19",X"10",X"F4",X"C9",X"D5",X"C5",X"78",X"2F",X"CB",X"3F",X"CB",X"3F",
		X"CB",X"3F",X"3D",X"47",X"69",X"CB",X"3D",X"CB",X"3D",X"CB",X"3D",X"2D",X"26",X"00",X"3E",X"05",
		X"CB",X"25",X"CB",X"14",X"3D",X"20",X"F9",X"11",X"40",X"A4",X"19",X"48",X"06",X"00",X"09",X"7E",
		X"C1",X"D1",X"C9",X"E5",X"2A",X"1E",X"A8",X"3A",X"1D",X"A8",X"86",X"32",X"1D",X"A8",X"23",X"26",
		X"30",X"22",X"1E",X"A8",X"E1",X"C9",X"D5",X"E5",X"6F",X"26",X"00",X"11",X"B3",X"40",X"19",X"7E",
		X"E1",X"D1",X"C9",X"0C",X"00",X"00",X"00",X"03",X"02",X"08",X"0C",X"03",X"0C",X"0C",X"01",X"02",
		X"03",X"05",X"00",X"03",X"0C",X"0D",X"07",X"0E",X"0B",X"0F",X"09",X"05",X"06",X"0A",X"00",X"03",
		X"03",X"0C",X"0C",X"00",X"03",X"03",X"0C",X"0C",X"01",X"03",X"04",X"0C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"FF",X"FF",X"FF",X"FF",X"0E",X"09",X"02",X"00",X"0C",X"0C",X"0C",
		X"0C",X"FF",X"FF",X"03",X"0C",X"0D",X"07",X"0E",X"0B",X"0F",X"09",X"05",X"06",X"0A",X"00",X"00",
		X"00",X"00",X"00",X"01",X"04",X"02",X"08",X"03",X"03",X"DD",X"21",X"14",X"A8",X"3E",X"FF",X"DD",
		X"77",X"00",X"DD",X"77",X"01",X"DD",X"77",X"02",X"DD",X"77",X"03",X"21",X"42",X"A4",X"16",X"10",
		X"06",X"1C",X"1E",X"F0",X"3E",X"35",X"BE",X"28",X"14",X"23",X"7B",X"D6",X"08",X"5F",X"10",X"F4",
		X"23",X"23",X"23",X"23",X"7A",X"C6",X"08",X"57",X"FE",X"E0",X"20",X"E4",X"C9",X"7A",X"C6",X"04",
		X"DD",X"77",X"01",X"7B",X"D6",X"0C",X"DD",X"77",X"00",X"DD",X"23",X"DD",X"23",X"C3",X"29",X"41",
		X"3A",X"C0",X"A8",X"6F",X"26",X"00",X"06",X"06",X"CB",X"25",X"CB",X"14",X"10",X"FA",X"11",X"00",
		X"2C",X"19",X"7E",X"32",X"9C",X"A8",X"23",X"7E",X"32",X"9D",X"A8",X"23",X"7E",X"32",X"9E",X"A8",
		X"23",X"7E",X"32",X"B0",X"A8",X"23",X"7E",X"32",X"B1",X"A8",X"23",X"7E",X"32",X"B2",X"A8",X"23",
		X"7E",X"32",X"B3",X"A8",X"23",X"7E",X"32",X"88",X"A8",X"23",X"7E",X"32",X"B5",X"A8",X"23",X"7E",
		X"32",X"9F",X"A8",X"32",X"04",X"A8",X"32",X"05",X"A8",X"23",X"7E",X"32",X"87",X"A8",X"23",X"23",
		X"23",X"23",X"23",X"11",X"62",X"AC",X"3E",X"07",X"32",X"12",X"A8",X"3E",X"07",X"32",X"13",X"A8",
		X"7E",X"E5",X"D5",X"D5",X"E1",X"CD",X"D9",X"41",X"E1",X"D1",X"01",X"80",X"FF",X"09",X"EB",X"23",
		X"3A",X"13",X"A8",X"3D",X"32",X"13",X"A8",X"20",X"E7",X"EB",X"01",X"84",X"03",X"09",X"EB",X"3A",
		X"12",X"A8",X"3D",X"32",X"12",X"A8",X"20",X"D3",X"C9",X"C5",X"D5",X"E5",X"DD",X"E5",X"E5",X"4F",
		X"06",X"00",X"3E",X"05",X"CB",X"21",X"CB",X"10",X"3D",X"20",X"F9",X"21",X"00",X"10",X"09",X"E5",
		X"DD",X"E1",X"E1",X"E5",X"11",X"80",X"03",X"19",X"EB",X"E1",X"3E",X"04",X"32",X"11",X"A8",X"3E",
		X"04",X"32",X"10",X"A8",X"01",X"E0",X"FF",X"DD",X"7E",X"00",X"77",X"DD",X"7E",X"10",X"12",X"09",
		X"EB",X"09",X"EB",X"DD",X"23",X"3A",X"10",X"A8",X"3D",X"32",X"10",X"A8",X"20",X"E9",X"01",X"81",
		X"00",X"09",X"EB",X"09",X"EB",X"3A",X"11",X"A8",X"3D",X"32",X"11",X"A8",X"20",X"D1",X"DD",X"E1",
		X"E1",X"D1",X"C1",X"C9",X"3A",X"0B",X"A8",X"FE",X"00",X"28",X"0E",X"3A",X"F0",X"A8",X"FE",X"01",
		X"C8",X"3E",X"01",X"32",X"F0",X"A8",X"C3",X"55",X"42",X"3A",X"F0",X"A8",X"FE",X"00",X"C8",X"3E",
		X"00",X"32",X"F0",X"A8",X"C9",X"3A",X"A0",X"A8",X"FE",X"00",X"C0",X"3A",X"93",X"A8",X"FE",X"00",
		X"C8",X"3D",X"32",X"93",X"A8",X"CD",X"76",X"3C",X"DD",X"21",X"A0",X"A8",X"3E",X"20",X"DD",X"77",
		X"00",X"3A",X"09",X"A8",X"DD",X"77",X"01",X"2A",X"50",X"B0",X"CD",X"8C",X"42",X"61",X"22",X"5E",
		X"B0",X"2A",X"50",X"B4",X"78",X"F6",X"05",X"6F",X"22",X"5E",X"B4",X"C9",X"3A",X"A1",X"A8",X"01",
		X"0B",X"40",X"FE",X"00",X"C8",X"01",X"05",X"80",X"FE",X"01",X"C8",X"01",X"0B",X"00",X"FE",X"02",
		X"C8",X"01",X"05",X"00",X"C9",X"21",X"97",X"A8",X"35",X"C0",X"3E",X"04",X"77",X"DD",X"21",X"A0",
		X"A8",X"DD",X"7E",X"00",X"FE",X"00",X"C8",X"3A",X"5F",X"B0",X"3C",X"06",X"05",X"FE",X"09",X"28",
		X"07",X"06",X"0B",X"FE",X"0F",X"28",X"01",X"47",X"78",X"32",X"5F",X"B0",X"DD",X"7E",X"00",X"FE",
		X"01",X"28",X"05",X"DD",X"35",X"00",X"18",X"26",X"DD",X"E5",X"3E",X"08",X"06",X"0F",X"CD",X"F2",
		X"3C",X"DD",X"E1",X"FE",X"FF",X"28",X"17",X"3E",X"FF",X"32",X"5F",X"B0",X"21",X"93",X"A8",X"34",
		X"CD",X"76",X"3C",X"3E",X"00",X"32",X"A0",X"A8",X"3E",X"01",X"CD",X"E2",X"3B",X"C9",X"21",X"5E",
		X"B0",X"11",X"5F",X"B4",X"DD",X"E5",X"3A",X"A1",X"A8",X"F5",X"CD",X"3A",X"55",X"F1",X"47",X"3A",
		X"A1",X"A8",X"B8",X"28",X"0D",X"CD",X"8C",X"42",X"78",X"F6",X"05",X"32",X"5E",X"B4",X"79",X"32",
		X"5F",X"B0",X"DD",X"E1",X"3A",X"91",X"A8",X"FE",X"FF",X"28",X"7E",X"3A",X"90",X"A8",X"FE",X"21",
		X"28",X"22",X"FE",X"24",X"20",X"73",X"3A",X"5E",X"B0",X"32",X"60",X"B0",X"3A",X"5F",X"B4",X"D6",
		X"04",X"32",X"61",X"B4",X"2A",X"94",X"A8",X"3E",X"1F",X"77",X"11",X"E0",X"FF",X"19",X"3E",X"1E",
		X"77",X"C3",X"6E",X"43",X"3A",X"5E",X"B0",X"D6",X"04",X"32",X"60",X"B0",X"3A",X"5F",X"B4",X"C6",
		X"04",X"32",X"61",X"B4",X"2A",X"94",X"A8",X"3E",X"1C",X"77",X"3E",X"1D",X"23",X"77",X"3E",X"9C",
		X"32",X"61",X"B0",X"3E",X"09",X"32",X"60",X"B4",X"3E",X"04",X"32",X"96",X"A8",X"CD",X"0F",X"4A",
		X"2A",X"5E",X"B0",X"7D",X"C6",X"10",X"6F",X"26",X"0A",X"22",X"62",X"B0",X"2A",X"5E",X"B4",X"2E",
		X"03",X"22",X"62",X"B4",X"3E",X"20",X"32",X"99",X"A8",X"3E",X"32",X"CD",X"E2",X"3B",X"3E",X"00",
		X"32",X"A0",X"A8",X"3E",X"FF",X"32",X"5F",X"B0",X"C9",X"C9",X"3A",X"78",X"A8",X"FE",X"00",X"C8",
		X"3E",X"0E",X"06",X"08",X"CD",X"F2",X"3C",X"FE",X"FF",X"C8",X"2A",X"5C",X"B0",X"7D",X"C6",X"08",
		X"6F",X"26",X"09",X"22",X"62",X"B0",X"2A",X"5C",X"B4",X"2E",X"03",X"22",X"62",X"B4",X"3E",X"20",
		X"32",X"99",X"A8",X"3E",X"0A",X"CD",X"E2",X"3B",X"3A",X"7B",X"A8",X"06",X"40",X"3A",X"85",X"A8",
		X"80",X"30",X"02",X"3E",X"FF",X"32",X"85",X"A8",X"CD",X"59",X"3D",X"3E",X"FF",X"32",X"5D",X"B0",
		X"3E",X"00",X"32",X"78",X"A8",X"3A",X"93",X"A8",X"3C",X"32",X"93",X"A8",X"CD",X"76",X"3C",X"CD",
		X"32",X"4A",X"C9",X"DD",X"21",X"78",X"A8",X"DD",X"7E",X"00",X"FE",X"00",X"C8",X"21",X"5C",X"B0",
		X"11",X"5D",X"B4",X"CD",X"2B",X"55",X"3A",X"F2",X"A8",X"3D",X"32",X"F2",X"A8",X"FE",X"00",X"20",
		X"2B",X"3E",X"03",X"32",X"F2",X"A8",X"3A",X"5C",X"B4",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",
		X"3F",X"CB",X"3F",X"CB",X"3F",X"3C",X"CB",X"27",X"CB",X"27",X"CB",X"27",X"CB",X"27",X"CB",X"27",
		X"CB",X"27",X"F6",X"39",X"32",X"5C",X"B4",X"3E",X"04",X"32",X"5D",X"B0",X"3A",X"91",X"A8",X"FE",
		X"FF",X"C8",X"3A",X"90",X"A8",X"FE",X"21",X"28",X"05",X"FE",X"24",X"28",X"01",X"C9",X"DD",X"21",
		X"78",X"A8",X"3E",X"FD",X"DD",X"86",X"03",X"30",X"04",X"DD",X"77",X"03",X"C9",X"3E",X"00",X"DD",
		X"77",X"00",X"3E",X"FF",X"32",X"5D",X"B0",X"C9",X"E5",X"D5",X"C5",X"DD",X"E5",X"FD",X"E5",X"7E",
		X"E6",X"07",X"FE",X"04",X"C2",X"2D",X"45",X"1A",X"E6",X"07",X"FE",X"04",X"C2",X"2D",X"45",X"46",
		X"1A",X"4F",X"CD",X"68",X"40",X"32",X"8E",X"A8",X"23",X"7E",X"2B",X"FE",X"0B",X"CA",X"35",X"45",
		X"7E",X"FE",X"36",X"CA",X"7D",X"45",X"FE",X"08",X"20",X"51",X"3A",X"8B",X"A8",X"FE",X"00",X"C2",
		X"2D",X"45",X"3A",X"89",X"A8",X"E6",X"F8",X"CA",X"2D",X"45",X"3E",X"01",X"CD",X"E2",X"3B",X"3A",
		X"89",X"A8",X"47",X"3A",X"85",X"A8",X"80",X"30",X"02",X"3E",X"FF",X"32",X"85",X"A8",X"3E",X"00",
		X"32",X"89",X"A8",X"CD",X"05",X"4A",X"3E",X"04",X"32",X"8B",X"A8",X"3A",X"50",X"B0",X"D6",X"02",
		X"32",X"56",X"B0",X"3E",X"9C",X"32",X"57",X"B0",X"3A",X"51",X"B4",X"C6",X"08",X"32",X"57",X"B4",
		X"3E",X"09",X"32",X"56",X"B4",X"CD",X"59",X"3D",X"C3",X"2D",X"45",X"FE",X"21",X"28",X"09",X"FE",
		X"54",X"CA",X"14",X"46",X"FE",X"24",X"20",X"25",X"CD",X"00",X"4A",X"3E",X"01",X"CD",X"E2",X"3B",
		X"3E",X"04",X"32",X"8A",X"A8",X"3A",X"88",X"A8",X"2F",X"47",X"3A",X"85",X"A8",X"80",X"38",X"07",
		X"3E",X"FF",X"32",X"8C",X"A8",X"3E",X"00",X"32",X"85",X"A8",X"CD",X"59",X"3D",X"FD",X"E1",X"DD",
		X"E1",X"C1",X"D1",X"E1",X"C9",X"3A",X"86",X"A8",X"FE",X"02",X"20",X"F1",X"23",X"3E",X"0D",X"77",
		X"23",X"3E",X"0E",X"77",X"3A",X"50",X"B0",X"D6",X"04",X"32",X"58",X"B0",X"D6",X"10",X"32",X"5A",
		X"B0",X"3A",X"51",X"B4",X"32",X"59",X"B4",X"32",X"5B",X"B4",X"3E",X"09",X"32",X"58",X"B4",X"32",
		X"5A",X"B4",X"3E",X"9B",X"32",X"59",X"B0",X"32",X"5B",X"B0",X"3E",X"04",X"32",X"8D",X"A8",X"3E",
		X"64",X"CD",X"E2",X"3B",X"CD",X"9D",X"4D",X"CD",X"59",X"3D",X"C3",X"2D",X"45",X"3A",X"78",X"A8",
		X"FE",X"00",X"C2",X"2D",X"45",X"3E",X"05",X"CD",X"E2",X"3B",X"DD",X"21",X"78",X"A8",X"3E",X"01",
		X"DD",X"77",X"00",X"3E",X"08",X"DD",X"77",X"02",X"3E",X"20",X"DD",X"77",X"03",X"3E",X"01",X"DD",
		X"77",X"04",X"DD",X"77",X"05",X"CD",X"FB",X"49",X"CD",X"93",X"40",X"E6",X"01",X"28",X"16",X"3E",
		X"02",X"DD",X"77",X"01",X"3A",X"50",X"B0",X"D6",X"0F",X"32",X"5C",X"B0",X"3A",X"51",X"B4",X"32",
		X"5D",X"B4",X"C3",X"DA",X"45",X"3E",X"00",X"DD",X"77",X"01",X"3A",X"50",X"B0",X"C6",X"08",X"32",
		X"5C",X"B0",X"3A",X"51",X"B4",X"D6",X"08",X"32",X"5D",X"B4",X"3E",X"0F",X"32",X"5C",X"B4",X"3E",
		X"C0",X"32",X"5D",X"B0",X"3A",X"50",X"B0",X"32",X"52",X"B0",X"32",X"54",X"B0",X"3A",X"51",X"B4",
		X"D6",X"08",X"32",X"55",X"B4",X"D6",X"10",X"32",X"53",X"B4",X"3E",X"09",X"32",X"52",X"B4",X"32",
		X"54",X"B4",X"3E",X"90",X"32",X"53",X"B0",X"3E",X"91",X"32",X"55",X"B0",X"3E",X"04",X"32",X"8F",
		X"A8",X"C3",X"2D",X"45",X"CD",X"37",X"4A",X"3E",X"55",X"77",X"3E",X"80",X"32",X"B4",X"A8",X"2A",
		X"50",X"B0",X"26",X"0F",X"2D",X"22",X"64",X"B0",X"2A",X"50",X"B4",X"24",X"22",X"64",X"B4",X"3E",
		X"0F",X"CD",X"E2",X"3B",X"DD",X"21",X"20",X"A8",X"06",X"08",X"11",X"08",X"00",X"DD",X"7E",X"00",
		X"FE",X"00",X"28",X"05",X"3E",X"02",X"DD",X"77",X"00",X"DD",X"19",X"10",X"F0",X"C3",X"2D",X"45",
		X"3A",X"98",X"A8",X"3D",X"32",X"98",X"A8",X"20",X"20",X"3A",X"86",X"A8",X"CB",X"27",X"EE",X"FF",
		X"E6",X"07",X"32",X"98",X"A8",X"3A",X"51",X"B0",X"06",X"99",X"FE",X"99",X"20",X"02",X"06",X"9A",
		X"78",X"32",X"51",X"B0",X"3E",X"02",X"32",X"50",X"B4",X"3E",X"02",X"77",X"C9",X"21",X"08",X"A8",
		X"35",X"28",X"01",X"C9",X"3A",X"BE",X"A8",X"3D",X"32",X"BE",X"A8",X"20",X"11",X"3E",X"50",X"32",
		X"BE",X"A8",X"3A",X"86",X"A8",X"FE",X"02",X"20",X"05",X"3E",X"02",X"CD",X"D4",X"49",X"3A",X"98",
		X"A8",X"3D",X"32",X"98",X"A8",X"20",X"20",X"3A",X"86",X"A8",X"CB",X"27",X"EE",X"FF",X"E6",X"07",
		X"32",X"98",X"A8",X"3A",X"51",X"B0",X"06",X"99",X"FE",X"99",X"20",X"02",X"06",X"9A",X"78",X"32",
		X"51",X"B0",X"3E",X"02",X"32",X"50",X"B4",X"3E",X"08",X"77",X"21",X"50",X"B0",X"11",X"51",X"B4",
		X"3A",X"80",X"A8",X"FE",X"00",X"20",X"05",X"3E",X"01",X"32",X"F1",X"A8",X"3A",X"80",X"A8",X"FE",
		X"00",X"C4",X"95",X"48",X"3A",X"F1",X"A8",X"FE",X"00",X"C8",X"3A",X"09",X"A8",X"FE",X"00",X"20",
		X"04",X"34",X"C3",X"0A",X"47",X"FE",X"01",X"20",X"06",X"1A",X"3D",X"12",X"C3",X"0A",X"47",X"FE",
		X"02",X"20",X"04",X"35",X"C3",X"0A",X"47",X"1A",X"3C",X"12",X"CD",X"78",X"44",X"7E",X"E6",X"07",
		X"32",X"10",X"A8",X"1A",X"E6",X"07",X"32",X"11",X"A8",X"46",X"1A",X"4F",X"CD",X"68",X"40",X"CD",
		X"A6",X"40",X"47",X"3A",X"0C",X"A8",X"FE",X"00",X"28",X"0A",X"78",X"E6",X"01",X"28",X"05",X"3E",
		X"00",X"C3",X"A1",X"47",X"3A",X"0D",X"A8",X"FE",X"00",X"28",X"0A",X"78",X"E6",X"02",X"28",X"05",
		X"3E",X"02",X"C3",X"A1",X"47",X"3A",X"0E",X"A8",X"FE",X"00",X"28",X"0A",X"78",X"E6",X"08",X"28",
		X"05",X"3E",X"03",X"C3",X"A1",X"47",X"3A",X"0F",X"A8",X"FE",X"00",X"28",X"0A",X"78",X"E6",X"04",
		X"28",X"05",X"3E",X"01",X"C3",X"A1",X"47",X"50",X"3A",X"09",X"A8",X"5F",X"01",X"15",X"56",X"6B",
		X"26",X"00",X"09",X"7E",X"A2",X"C0",X"7B",X"3C",X"E6",X"03",X"6F",X"26",X"00",X"09",X"7E",X"A2",
		X"28",X"07",X"7B",X"3C",X"E6",X"03",X"C3",X"A1",X"47",X"7B",X"3D",X"E6",X"03",X"6F",X"26",X"00",
		X"09",X"7E",X"A2",X"28",X"07",X"7B",X"3D",X"E6",X"03",X"C3",X"A1",X"47",X"7B",X"3C",X"3C",X"E6",
		X"03",X"47",X"3A",X"09",X"A8",X"B8",X"C8",X"E6",X"01",X"28",X"0A",X"78",X"E6",X"01",X"28",X"0A",
		X"78",X"32",X"09",X"A8",X"C9",X"78",X"E6",X"01",X"28",X"F6",X"3A",X"10",X"A8",X"FE",X"04",X"C0",
		X"3A",X"11",X"A8",X"FE",X"04",X"C0",X"78",X"32",X"09",X"A8",X"3A",X"51",X"B4",X"E6",X"FC",X"F6",
		X"04",X"32",X"51",X"B4",X"3A",X"50",X"B0",X"E6",X"FC",X"F6",X"04",X"32",X"50",X"B0",X"C9",X"C5",
		X"01",X"00",X"01",X"0D",X"20",X"FD",X"05",X"20",X"FA",X"C1",X"C9",X"E5",X"DD",X"E5",X"21",X"0A",
		X"A8",X"06",X"06",X"36",X"00",X"23",X"10",X"FB",X"3E",X"00",X"32",X"01",X"A8",X"32",X"02",X"A8",
		X"3A",X"00",X"C3",X"E6",X"08",X"20",X"05",X"3E",X"01",X"32",X"01",X"A8",X"3A",X"00",X"C3",X"E6",
		X"10",X"20",X"05",X"3E",X"01",X"32",X"02",X"A8",X"3A",X"CB",X"A8",X"FE",X"00",X"CA",X"2B",X"48",
		X"3A",X"9A",X"A8",X"FE",X"01",X"CA",X"2B",X"48",X"C3",X"60",X"48",X"DD",X"21",X"0A",X"A8",X"3A",
		X"20",X"C3",X"CB",X"3F",X"38",X"03",X"DD",X"34",X"04",X"CB",X"3F",X"38",X"03",X"DD",X"34",X"05",
		X"CB",X"3F",X"38",X"03",X"DD",X"34",X"02",X"CB",X"3F",X"38",X"03",X"DD",X"34",X"03",X"CB",X"3F",
		X"38",X"03",X"DD",X"34",X"01",X"CB",X"3F",X"38",X"03",X"DD",X"34",X"01",X"DD",X"E1",X"E1",X"C9",
		X"DD",X"21",X"0A",X"A8",X"3A",X"40",X"C3",X"CB",X"3F",X"38",X"03",X"DD",X"34",X"04",X"CB",X"3F",
		X"38",X"03",X"DD",X"34",X"05",X"CB",X"3F",X"38",X"03",X"DD",X"34",X"02",X"CB",X"3F",X"38",X"03",
		X"DD",X"34",X"03",X"CB",X"3F",X"38",X"03",X"DD",X"34",X"01",X"CB",X"3F",X"38",X"03",X"DD",X"34",
		X"01",X"DD",X"E1",X"E1",X"C9",X"E5",X"D5",X"C5",X"CD",X"9F",X"48",X"C1",X"D1",X"E1",X"C9",X"E5",
		X"21",X"0C",X"A8",X"7E",X"23",X"86",X"23",X"86",X"23",X"86",X"E1",X"FE",X"00",X"C2",X"FC",X"48",
		X"7E",X"E6",X"07",X"FE",X"04",X"C0",X"1A",X"E6",X"07",X"FE",X"04",X"C0",X"46",X"1A",X"4F",X"CD",
		X"68",X"40",X"CD",X"A6",X"40",X"47",X"3A",X"09",X"A8",X"3C",X"E6",X"03",X"6F",X"26",X"00",X"11",
		X"15",X"56",X"19",X"7E",X"A0",X"28",X"06",X"3E",X"00",X"32",X"F1",X"A8",X"C9",X"3A",X"09",X"A8",
		X"3D",X"E6",X"03",X"6F",X"26",X"00",X"19",X"7E",X"A0",X"20",X"EC",X"3A",X"09",X"A8",X"6F",X"26",
		X"00",X"19",X"7E",X"A0",X"28",X"E1",X"3E",X"01",X"32",X"F1",X"A8",X"C9",X"E5",X"D5",X"7E",X"E6",
		X"07",X"FE",X"04",X"20",X"0A",X"1A",X"E6",X"07",X"FE",X"04",X"20",X"03",X"CD",X"BC",X"48",X"D1",
		X"E1",X"46",X"1A",X"4F",X"E5",X"D5",X"CD",X"68",X"40",X"CD",X"A6",X"40",X"D1",X"E1",X"47",X"3A",
		X"0C",X"A8",X"FE",X"00",X"28",X"16",X"78",X"E6",X"01",X"28",X"11",X"3E",X"00",X"32",X"09",X"A8",
		X"3E",X"01",X"32",X"F1",X"A8",X"1A",X"E6",X"FC",X"F6",X"04",X"12",X"C9",X"3A",X"0D",X"A8",X"FE",
		X"00",X"28",X"16",X"78",X"E6",X"02",X"28",X"11",X"3E",X"02",X"32",X"09",X"A8",X"3E",X"01",X"32",
		X"F1",X"A8",X"1A",X"E6",X"FC",X"F6",X"04",X"12",X"C9",X"3A",X"0E",X"A8",X"FE",X"00",X"28",X"16",
		X"78",X"E6",X"08",X"28",X"11",X"3E",X"03",X"32",X"09",X"A8",X"3E",X"01",X"32",X"F1",X"A8",X"7E",
		X"E6",X"FC",X"F6",X"04",X"77",X"C9",X"3A",X"0F",X"A8",X"FE",X"00",X"C8",X"78",X"E6",X"04",X"C8",
		X"3E",X"01",X"32",X"09",X"A8",X"3E",X"01",X"32",X"F1",X"A8",X"7E",X"E6",X"FC",X"F6",X"04",X"77",
		X"C9",X"21",X"20",X"A6",X"34",X"C9",X"C9",X"CD",X"79",X"4B",X"3A",X"A9",X"A8",X"FE",X"00",X"C0",
		X"CD",X"EB",X"47",X"3A",X"0B",X"A8",X"FE",X"00",X"C0",X"CD",X"C2",X"49",X"3A",X"A9",X"A8",X"FE",
		X"00",X"C0",X"3E",X"01",X"32",X"F4",X"A8",X"CD",X"D5",X"3A",X"3E",X"00",X"32",X"F4",X"A8",X"C3",
		X"97",X"49",X"16",X"40",X"0D",X"20",X"FD",X"3A",X"A9",X"A8",X"FE",X"00",X"C0",X"05",X"20",X"F4",
		X"15",X"20",X"F1",X"C9",X"F5",X"3A",X"F4",X"A8",X"FE",X"00",X"20",X"04",X"F1",X"C3",X"E3",X"49",
		X"F1",X"3E",X"00",X"32",X"00",X"C0",X"3E",X"FF",X"32",X"04",X"C3",X"3E",X"00",X"32",X"04",X"C3",
		X"C9",X"3E",X"4D",X"C3",X"D4",X"49",X"3E",X"4A",X"C3",X"D4",X"49",X"3E",X"09",X"C3",X"D4",X"49",
		X"3E",X"55",X"C3",X"D4",X"49",X"3E",X"4F",X"C3",X"D4",X"49",X"3E",X"47",X"C3",X"D4",X"49",X"3E",
		X"49",X"C3",X"D4",X"49",X"3E",X"47",X"C3",X"D4",X"49",X"3E",X"09",X"C3",X"D4",X"49",X"3E",X"10",
		X"C3",X"D4",X"49",X"3E",X"15",X"C3",X"D4",X"49",X"3E",X"4C",X"C3",X"D4",X"49",X"3E",X"4F",X"C3",
		X"D4",X"49",X"3E",X"4C",X"C3",X"D4",X"49",X"3E",X"02",X"C3",X"D4",X"49",X"21",X"60",X"A8",X"11",
		X"61",X"A8",X"01",X"0B",X"00",X"36",X"20",X"ED",X"B0",X"3A",X"00",X"C2",X"06",X"00",X"E6",X"80",
		X"20",X"01",X"04",X"78",X"32",X"80",X"A8",X"3A",X"00",X"C2",X"06",X"00",X"E6",X"40",X"20",X"01",
		X"04",X"78",X"32",X"CD",X"A8",X"3A",X"60",X"C3",X"06",X"00",X"E6",X"80",X"20",X"01",X"04",X"78",
		X"32",X"CB",X"A8",X"3A",X"60",X"C3",X"06",X"00",X"E6",X"40",X"28",X"01",X"04",X"78",X"32",X"CC",
		X"A8",X"3A",X"60",X"C3",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"E6",X"03",X"EE",X"03",
		X"C6",X"02",X"32",X"C2",X"A8",X"3A",X"60",X"C3",X"06",X"40",X"E6",X"08",X"28",X"02",X"06",X"60",
		X"78",X"32",X"CA",X"A8",X"3A",X"60",X"C3",X"E6",X"07",X"EE",X"07",X"32",X"CE",X"A8",X"3A",X"00",
		X"C2",X"E6",X"03",X"EE",X"03",X"6F",X"26",X"00",X"11",X"F3",X"4A",X"19",X"7E",X"32",X"B8",X"A8",
		X"11",X"08",X"00",X"19",X"7E",X"32",X"B9",X"A8",X"3A",X"00",X"C2",X"CB",X"3F",X"CB",X"3F",X"E6",
		X"03",X"EE",X"03",X"6F",X"26",X"00",X"11",X"F3",X"4A",X"19",X"7E",X"32",X"BA",X"A8",X"11",X"08",
		X"00",X"19",X"7E",X"32",X"BB",X"A8",X"3A",X"B8",X"A8",X"32",X"FD",X"A8",X"3A",X"BA",X"A8",X"32",
		X"FE",X"A8",X"C9",X"01",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"03",X"05",X"01",
		X"01",X"01",X"01",X"C8",X"18",X"C8",X"1A",X"C8",X"1B",X"C8",X"1D",X"C8",X"1F",X"C8",X"21",X"C8",
		X"23",X"C8",X"1F",X"C8",X"25",X"C8",X"1D",X"B8",X"19",X"B8",X"1A",X"B8",X"1C",X"B8",X"1E",X"B8",
		X"20",X"B8",X"22",X"B8",X"24",X"B8",X"20",X"B8",X"26",X"B8",X"1E",X"82",X"C8",X"82",X"B8",X"82",
		X"A8",X"82",X"98",X"82",X"88",X"82",X"68",X"82",X"58",X"82",X"48",X"82",X"38",X"82",X"28",X"82",
		X"C8",X"C2",X"B8",X"82",X"A8",X"82",X"98",X"82",X"88",X"82",X"68",X"82",X"58",X"82",X"48",X"82",
		X"38",X"82",X"28",X"09",X"A6",X"20",X"20",X"20",X"FF",X"CD",X"A6",X"30",X"02",X"12",X"09",X"07",
		X"08",X"14",X"20",X"13",X"10",X"01",X"12",X"0B",X"13",X"FF",X"5A",X"A6",X"20",X"D0",X"20",X"CD",
		X"CE",X"CF",X"CF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CD",X"29",X"4C",X"CD",X"04",X"4C",X"21",
		X"5E",X"A4",X"11",X"20",X"00",X"06",X"18",X"36",X"00",X"19",X"10",X"FB",X"CD",X"9A",X"4C",X"21",
		X"03",X"4B",X"11",X"40",X"B0",X"01",X"28",X"00",X"ED",X"B0",X"21",X"2B",X"4B",X"11",X"40",X"B4",
		X"01",X"28",X"00",X"ED",X"B0",X"21",X"53",X"4B",X"5E",X"23",X"56",X"23",X"46",X"23",X"CD",X"DB",
		X"36",X"23",X"7E",X"FE",X"FF",X"20",X"F1",X"CD",X"BB",X"4B",X"C9",X"3E",X"FF",X"32",X"8F",X"B0",
		X"32",X"9F",X"B0",X"32",X"AF",X"B0",X"32",X"BF",X"B0",X"32",X"CF",X"B0",X"21",X"80",X"B0",X"11",
		X"CF",X"A6",X"06",X"34",X"CD",X"DB",X"36",X"21",X"90",X"B0",X"11",X"D1",X"A6",X"06",X"2C",X"CD",
		X"DB",X"36",X"21",X"A0",X"B0",X"11",X"D3",X"A6",X"06",X"2C",X"CD",X"DB",X"36",X"21",X"B0",X"B0",
		X"11",X"D5",X"A6",X"06",X"2C",X"CD",X"DB",X"36",X"21",X"C0",X"B0",X"11",X"D7",X"A6",X"06",X"2C",
		X"CD",X"DB",X"36",X"C9",X"21",X"00",X"A9",X"11",X"01",X"A9",X"36",X"20",X"01",X"FF",X"06",X"ED",
		X"B0",X"CD",X"29",X"4C",X"CD",X"F5",X"37",X"06",X"1C",X"C5",X"CD",X"1D",X"38",X"01",X"00",X"10",
		X"0D",X"20",X"FD",X"10",X"FB",X"C1",X"10",X"F1",X"C9",X"21",X"40",X"B0",X"11",X"41",X"B0",X"01",
		X"3F",X"00",X"36",X"FF",X"ED",X"B0",X"21",X"40",X"B4",X"11",X"41",X"B4",X"01",X"3F",X"00",X"36",
		X"FF",X"ED",X"B0",X"C9",X"3A",X"A9",X"A8",X"47",X"3E",X"30",X"32",X"C5",X"A8",X"32",X"C6",X"A8",
		X"78",X"FE",X"00",X"28",X"19",X"3A",X"C6",X"A8",X"3C",X"32",X"C6",X"A8",X"FE",X"3A",X"20",X"0C",
		X"3E",X"30",X"32",X"C6",X"A8",X"3A",X"C5",X"A8",X"3C",X"32",X"C5",X"A8",X"10",X"E7",X"21",X"92",
		X"4C",X"11",X"9F",X"A5",X"06",X"30",X"CD",X"DB",X"36",X"3A",X"C5",X"A8",X"F6",X"80",X"32",X"9F",
		X"A4",X"3A",X"C6",X"A8",X"F6",X"80",X"32",X"7F",X"A4",X"3E",X"30",X"32",X"9F",X"A0",X"32",X"7F",
		X"A0",X"C9",X"03",X"12",X"05",X"04",X"09",X"14",X"13",X"FF",X"DD",X"21",X"A2",X"A7",X"FD",X"21",
		X"A2",X"A3",X"11",X"E0",X"FF",X"0E",X"1C",X"DD",X"E5",X"FD",X"E5",X"3E",X"20",X"06",X"1C",X"DD",
		X"77",X"00",X"FD",X"77",X"00",X"DD",X"19",X"FD",X"19",X"10",X"F4",X"FD",X"E1",X"DD",X"E1",X"FD",
		X"23",X"DD",X"23",X"0D",X"20",X"E1",X"C9",X"04",X"04",X"A0",X"00",X"05",X"06",X"80",X"00",X"06",
		X"07",X"70",X"00",X"07",X"08",X"60",X"00",X"08",X"10",X"20",X"00",X"08",X"10",X"20",X"00",X"08",
		X"10",X"20",X"00",X"08",X"20",X"20",X"00",X"3E",X"00",X"32",X"07",X"A8",X"3A",X"9E",X"A8",X"47",
		X"3A",X"CE",X"A8",X"80",X"47",X"3A",X"CF",X"A8",X"80",X"32",X"18",X"A8",X"6F",X"CB",X"3D",X"CB",
		X"3D",X"CB",X"25",X"CB",X"25",X"26",X"00",X"11",X"C7",X"4C",X"19",X"7E",X"32",X"87",X"A8",X"23",
		X"7E",X"32",X"88",X"A8",X"23",X"7E",X"32",X"9F",X"A8",X"3E",X"01",X"32",X"06",X"A8",X"32",X"07",
		X"A8",X"32",X"08",X"A8",X"32",X"1C",X"A8",X"32",X"92",X"A8",X"32",X"98",X"A8",X"32",X"B6",X"A8",
		X"3E",X"00",X"32",X"8C",X"A8",X"32",X"8E",X"A8",X"32",X"1B",X"A8",X"32",X"81",X"A8",X"32",X"8B",
		X"A8",X"32",X"8D",X"A8",X"32",X"8F",X"A8",X"32",X"96",X"A8",X"32",X"99",X"A8",X"32",X"B4",X"A8",
		X"32",X"78",X"A8",X"32",X"A0",X"A8",X"32",X"20",X"A8",X"32",X"28",X"A8",X"32",X"30",X"A8",X"32",
		X"38",X"A8",X"32",X"40",X"A8",X"32",X"48",X"A8",X"32",X"50",X"A8",X"32",X"58",X"A8",X"CD",X"93",
		X"40",X"E6",X"0F",X"32",X"89",X"A8",X"3E",X"34",X"32",X"82",X"A8",X"32",X"83",X"A8",X"3E",X"30",
		X"32",X"84",X"A8",X"3A",X"CA",X"A8",X"32",X"85",X"A8",X"CD",X"59",X"3D",X"CD",X"76",X"3C",X"3E",
		X"F0",X"32",X"C7",X"A8",X"3E",X"00",X"32",X"C8",X"A8",X"32",X"C9",X"A8",X"C9",X"CD",X"0A",X"4A",
		X"06",X"20",X"21",X"42",X"A0",X"0E",X"1C",X"16",X"1C",X"7E",X"EE",X"0D",X"77",X"23",X"15",X"20",
		X"F8",X"23",X"23",X"23",X"23",X"0D",X"20",X"EF",X"C5",X"01",X"00",X"08",X"0D",X"20",X"FD",X"10",
		X"FB",X"C1",X"10",X"DE",X"3E",X"40",X"32",X"85",X"A8",X"C9",X"2A",X"50",X"B0",X"E5",X"2A",X"50",
		X"B4",X"E5",X"CD",X"29",X"4C",X"E1",X"22",X"50",X"B4",X"E1",X"22",X"50",X"B0",X"CD",X"98",X"4E",
		X"CD",X"AF",X"4E",X"3E",X"00",X"32",X"F4",X"A8",X"21",X"8B",X"4E",X"11",X"4C",X"A6",X"06",X"35",
		X"CD",X"DB",X"36",X"21",X"91",X"4E",X"11",X"6E",X"A6",X"06",X"2D",X"CD",X"DB",X"36",X"3E",X"05",
		X"01",X"00",X"00",X"0D",X"20",X"FD",X"05",X"20",X"FA",X"3D",X"20",X"F7",X"3E",X"00",X"CD",X"D4",
		X"49",X"3A",X"C7",X"A8",X"C6",X"0A",X"47",X"CD",X"5C",X"4E",X"10",X"FB",X"3E",X"02",X"01",X"00",
		X"00",X"0D",X"20",X"FD",X"05",X"20",X"FA",X"3D",X"20",X"F7",X"3A",X"C7",X"A8",X"C6",X"0A",X"47",
		X"3E",X"00",X"32",X"F4",X"A8",X"C5",X"3E",X"01",X"CD",X"E2",X"3B",X"CD",X"4A",X"3E",X"01",X"00",
		X"02",X"0D",X"20",X"FD",X"05",X"20",X"FA",X"C1",X"10",X"EB",X"3E",X"04",X"01",X"00",X"00",X"0D",
		X"20",X"FD",X"05",X"20",X"FA",X"3D",X"20",X"F7",X"CD",X"D6",X"4E",X"C9",X"CD",X"1E",X"4A",X"11",
		X"00",X"10",X"1D",X"20",X"FD",X"15",X"20",X"FA",X"DD",X"21",X"EE",X"A5",X"DD",X"7E",X"00",X"FE",
		X"A0",X"20",X"02",X"3E",X"B0",X"3C",X"FE",X"BA",X"28",X"04",X"DD",X"77",X"00",X"C9",X"3E",X"B0",
		X"DD",X"77",X"00",X"11",X"20",X"00",X"DD",X"19",X"C3",X"6C",X"4E",X"02",X"0F",X"0E",X"15",X"13",
		X"FF",X"20",X"20",X"20",X"20",X"20",X"30",X"FF",X"21",X"40",X"A4",X"11",X"00",X"A9",X"01",X"80",
		X"03",X"ED",X"B0",X"21",X"40",X"A0",X"11",X"80",X"AC",X"01",X"80",X"03",X"ED",X"B0",X"C9",X"DD",
		X"21",X"EB",X"A6",X"FD",X"21",X"EB",X"A2",X"06",X"10",X"0E",X"05",X"3E",X"20",X"DD",X"77",X"00",
		X"3E",X"25",X"FD",X"77",X"00",X"DD",X"23",X"FD",X"23",X"0D",X"20",X"EF",X"11",X"DB",X"FF",X"DD",
		X"19",X"FD",X"19",X"10",X"E4",X"C9",X"21",X"00",X"A9",X"11",X"40",X"A4",X"01",X"78",X"03",X"ED",
		X"B0",X"CD",X"4A",X"3E",X"21",X"80",X"AC",X"11",X"40",X"A0",X"01",X"78",X"03",X"ED",X"B0",X"CD",
		X"4A",X"3E",X"C9",X"CD",X"29",X"4C",X"CD",X"9A",X"4C",X"21",X"03",X"4B",X"11",X"40",X"B0",X"01",
		X"28",X"00",X"ED",X"B0",X"21",X"2B",X"4B",X"11",X"40",X"B4",X"01",X"28",X"00",X"ED",X"B0",X"21",
		X"9D",X"4F",X"5E",X"23",X"56",X"23",X"46",X"23",X"CD",X"DB",X"36",X"23",X"7E",X"FE",X"FF",X"20",
		X"F1",X"CD",X"EB",X"47",X"3A",X"01",X"A8",X"FE",X"00",X"28",X"0D",X"3A",X"A9",X"A8",X"3D",X"32",
		X"A9",X"A8",X"CD",X"44",X"4C",X"3E",X"01",X"C9",X"3A",X"A9",X"A8",X"FE",X"01",X"CA",X"21",X"4F",
		X"C3",X"43",X"4F",X"CD",X"29",X"4C",X"CD",X"9A",X"4C",X"21",X"03",X"4B",X"11",X"40",X"B0",X"01",
		X"28",X"00",X"ED",X"B0",X"21",X"2B",X"4B",X"11",X"40",X"B4",X"01",X"28",X"00",X"ED",X"B0",X"21",
		X"CB",X"4F",X"5E",X"23",X"56",X"23",X"46",X"23",X"CD",X"DB",X"36",X"23",X"7E",X"FE",X"FF",X"20",
		X"F1",X"CD",X"EB",X"47",X"3A",X"01",X"A8",X"FE",X"00",X"28",X"0D",X"3A",X"A9",X"A8",X"3D",X"32",
		X"A9",X"A8",X"CD",X"44",X"4C",X"3E",X"01",X"C9",X"3A",X"02",X"A8",X"FE",X"00",X"28",X"E2",X"3A",
		X"A9",X"A8",X"3D",X"3D",X"32",X"A9",X"A8",X"CD",X"44",X"4C",X"3E",X"02",X"C9",X"09",X"A6",X"20",
		X"20",X"20",X"FF",X"4F",X"A7",X"30",X"10",X"12",X"05",X"13",X"13",X"20",X"0F",X"0E",X"05",X"20",
		X"10",X"0C",X"01",X"19",X"05",X"12",X"20",X"0F",X"0E",X"0C",X"19",X"FF",X"5A",X"A6",X"20",X"D0",
		X"20",X"CD",X"CE",X"CF",X"CF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"09",X"A6",X"20",X"20",X"20",
		X"FF",X"6F",X"A7",X"30",X"10",X"12",X"05",X"13",X"13",X"20",X"0F",X"0E",X"05",X"20",X"0F",X"12",
		X"20",X"14",X"17",X"0F",X"20",X"10",X"0C",X"01",X"19",X"05",X"12",X"13",X"FF",X"5A",X"A6",X"20",
		X"D0",X"20",X"CD",X"CE",X"CF",X"CF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CD",X"29",X"4C",X"CD",
		X"04",X"4C",X"CD",X"BA",X"3C",X"3A",X"9A",X"A8",X"FE",X"02",X"20",X"11",X"3A",X"CB",X"A8",X"FE",
		X"00",X"28",X"0A",X"3E",X"FF",X"32",X"02",X"C3",X"32",X"F3",X"A8",X"18",X"08",X"3E",X"00",X"32",
		X"02",X"C3",X"32",X"F3",X"A8",X"3A",X"9B",X"A8",X"C6",X"B0",X"32",X"CE",X"A6",X"3E",X"30",X"32",
		X"CE",X"A2",X"21",X"66",X"50",X"11",X"8E",X"A6",X"06",X"30",X"CD",X"DB",X"36",X"3A",X"C1",X"A8",
		X"FE",X"02",X"20",X"13",X"21",X"72",X"50",X"11",X"6C",X"A6",X"06",X"30",X"CD",X"DB",X"36",X"3A",
		X"9A",X"A8",X"C6",X"B0",X"32",X"AC",X"A5",X"3E",X"06",X"01",X"00",X"00",X"0D",X"20",X"FD",X"05",
		X"20",X"FA",X"3D",X"20",X"F7",X"C9",X"13",X"10",X"01",X"12",X"0B",X"13",X"20",X"0C",X"05",X"06",
		X"14",X"FF",X"10",X"0C",X"01",X"19",X"05",X"12",X"20",X"FF",X"06",X"00",X"11",X"87",X"B0",X"CD",
		X"74",X"51",X"FE",X"00",X"28",X"2D",X"11",X"97",X"B0",X"04",X"CD",X"74",X"51",X"FE",X"00",X"28",
		X"22",X"11",X"A7",X"B0",X"04",X"CD",X"74",X"51",X"FE",X"00",X"28",X"17",X"11",X"B7",X"B0",X"04",
		X"CD",X"74",X"51",X"FE",X"00",X"28",X"0C",X"11",X"C7",X"B0",X"04",X"CD",X"74",X"51",X"FE",X"00",
		X"28",X"01",X"C9",X"E5",X"C5",X"E5",X"48",X"06",X"00",X"CB",X"21",X"CB",X"21",X"CB",X"21",X"21",
		X"39",X"51",X"09",X"E5",X"DD",X"E1",X"21",X"C0",X"B0",X"11",X"D0",X"B0",X"DD",X"46",X"06",X"DD",
		X"4E",X"07",X"ED",X"B8",X"3E",X"32",X"32",X"90",X"B0",X"3C",X"32",X"A0",X"B0",X"3C",X"32",X"B0",
		X"B0",X"3C",X"32",X"C0",X"B0",X"E1",X"DD",X"56",X"00",X"DD",X"5E",X"01",X"01",X"06",X"00",X"ED",
		X"B0",X"DD",X"66",X"02",X"DD",X"6E",X"03",X"36",X"20",X"23",X"36",X"20",X"23",X"36",X"20",X"DD",
		X"E5",X"CD",X"BB",X"4B",X"21",X"61",X"51",X"11",X"29",X"A7",X"06",X"30",X"CD",X"DB",X"36",X"DD",
		X"E1",X"DD",X"66",X"04",X"DD",X"6E",X"05",X"DD",X"56",X"02",X"DD",X"5E",X"03",X"CD",X"A3",X"51",
		X"C1",X"E1",X"78",X"FE",X"00",X"CC",X"8C",X"52",X"3E",X"2E",X"32",X"81",X"B0",X"3E",X"20",X"32",
		X"82",X"B0",X"32",X"86",X"B0",X"32",X"8E",X"B0",X"C9",X"B0",X"87",X"B0",X"83",X"A6",X"6F",X"00",
		X"50",X"B0",X"97",X"B0",X"93",X"A6",X"71",X"00",X"40",X"B0",X"A7",X"B0",X"A3",X"A6",X"73",X"00",
		X"30",X"B0",X"B7",X"B0",X"B3",X"A6",X"75",X"00",X"20",X"B0",X"C7",X"B0",X"C3",X"A6",X"77",X"00",
		X"10",X"05",X"0E",X"14",X"05",X"12",X"20",X"09",X"0E",X"20",X"19",X"0F",X"15",X"12",X"20",X"0E",
		X"01",X"0D",X"05",X"FF",X"E5",X"D5",X"C5",X"06",X"06",X"1A",X"BE",X"28",X"10",X"FE",X"20",X"28",
		X"1C",X"7E",X"FE",X"20",X"28",X"11",X"1A",X"BE",X"38",X"13",X"C3",X"97",X"51",X"23",X"13",X"10",
		X"E8",X"C1",X"D1",X"E1",X"3E",X"FF",X"C9",X"C1",X"D1",X"E1",X"3E",X"FF",X"C9",X"C1",X"D1",X"E1",
		X"3E",X"00",X"C9",X"7C",X"E6",X"FB",X"47",X"4D",X"3E",X"03",X"32",X"10",X"A8",X"0A",X"EE",X"01",
		X"02",X"CD",X"81",X"52",X"0A",X"EE",X"01",X"02",X"C5",X"CD",X"EB",X"47",X"C1",X"3A",X"0B",X"A8",
		X"FE",X"00",X"20",X"21",X"3A",X"0E",X"A8",X"FE",X"00",X"28",X"09",X"7E",X"3D",X"E6",X"1F",X"F6",
		X"80",X"77",X"18",X"D9",X"3A",X"0F",X"A8",X"FE",X"00",X"28",X"D2",X"7E",X"3C",X"E6",X"1F",X"F6",
		X"80",X"77",X"C3",X"AD",X"51",X"7E",X"E6",X"7F",X"12",X"13",X"D5",X"11",X"E0",X"FF",X"19",X"E5",
		X"21",X"E0",X"FF",X"09",X"E5",X"C1",X"E1",X"D1",X"CD",X"81",X"52",X"CD",X"81",X"52",X"CD",X"81",
		X"52",X"CD",X"81",X"52",X"CD",X"81",X"52",X"3A",X"10",X"A8",X"3D",X"32",X"10",X"A8",X"C2",X"AD",
		X"51",X"C9",X"CD",X"29",X"4C",X"CD",X"04",X"4C",X"21",X"6E",X"52",X"11",X"8F",X"A6",X"06",X"30",
		X"CD",X"DB",X"36",X"3A",X"C1",X"A8",X"FE",X"02",X"20",X"13",X"21",X"78",X"52",X"11",X"71",X"A6",
		X"06",X"30",X"CD",X"DB",X"36",X"3A",X"9A",X"A8",X"C6",X"B0",X"32",X"B1",X"A5",X"3E",X"04",X"01",
		X"00",X"00",X"0D",X"20",X"FD",X"05",X"20",X"FA",X"3D",X"20",X"F7",X"CD",X"04",X"4C",X"3A",X"CC",
		X"A8",X"FE",X"01",X"20",X"03",X"C3",X"D0",X"52",X"CD",X"04",X"4C",X"21",X"60",X"A8",X"3A",X"9A",
		X"A8",X"FE",X"01",X"28",X"03",X"21",X"66",X"A8",X"CD",X"7A",X"50",X"3E",X"FF",X"C9",X"07",X"01",
		X"0D",X"05",X"20",X"0F",X"16",X"05",X"12",X"FF",X"10",X"0C",X"01",X"19",X"05",X"12",X"20",X"20",
		X"FF",X"C5",X"01",X"00",X"40",X"0D",X"20",X"FD",X"10",X"FB",X"C1",X"C9",X"C5",X"11",X"6C",X"A8",
		X"01",X"06",X"00",X"ED",X"B0",X"C1",X"C9",X"03",X"0F",X"0E",X"14",X"09",X"0E",X"15",X"05",X"FF",
		X"10",X"0C",X"01",X"19",X"FF",X"19",X"05",X"13",X"FF",X"0E",X"0F",X"20",X"FF",X"10",X"12",X"05",
		X"13",X"13",X"20",X"06",X"09",X"12",X"05",X"FF",X"21",X"A9",X"52",X"11",X"2B",X"A6",X"06",X"30",
		X"CD",X"DB",X"36",X"C9",X"21",X"A5",X"52",X"11",X"2B",X"A6",X"06",X"30",X"CD",X"DB",X"36",X"C9",
		X"21",X"97",X"52",X"11",X"86",X"A6",X"06",X"2C",X"CD",X"DB",X"36",X"21",X"A0",X"52",X"11",X"48",
		X"A6",X"06",X"2C",X"CD",X"DB",X"36",X"21",X"AD",X"52",X"11",X"B3",X"A6",X"06",X"2C",X"CD",X"DB",
		X"36",X"CD",X"C4",X"52",X"3E",X"00",X"32",X"10",X"A8",X"3E",X"20",X"32",X"10",X"A2",X"3E",X"B9",
		X"32",X"10",X"A6",X"3E",X"0C",X"32",X"11",X"A8",X"06",X"68",X"0D",X"20",X"FD",X"10",X"FB",X"CD",
		X"EB",X"47",X"3A",X"0F",X"A8",X"FE",X"00",X"C2",X"68",X"53",X"3A",X"0E",X"A8",X"FE",X"00",X"C2",
		X"68",X"53",X"3A",X"A9",X"A8",X"FE",X"00",X"28",X"18",X"3A",X"0B",X"A8",X"FE",X"00",X"28",X"11",
		X"3A",X"10",X"A8",X"FE",X"00",X"20",X"0A",X"21",X"A9",X"A8",X"35",X"CD",X"44",X"4C",X"3E",X"00",
		X"C9",X"3A",X"10",X"A8",X"FE",X"00",X"28",X"0A",X"3A",X"0B",X"A8",X"FE",X"00",X"28",X"03",X"C3",
		X"58",X"52",X"21",X"11",X"A8",X"35",X"C2",X"08",X"53",X"3A",X"10",X"A6",X"3D",X"FE",X"AF",X"CA",
		X"58",X"52",X"32",X"10",X"A6",X"C3",X"03",X"53",X"3A",X"10",X"A8",X"FE",X"00",X"20",X"0B",X"3E",
		X"01",X"32",X"10",X"A8",X"CD",X"B8",X"52",X"C3",X"22",X"53",X"3E",X"00",X"32",X"10",X"A8",X"CD",
		X"C4",X"52",X"C3",X"22",X"53",X"DD",X"E5",X"C5",X"D5",X"3A",X"A0",X"A8",X"FE",X"00",X"28",X"51",
		X"3E",X"00",X"DD",X"77",X"00",X"69",X"CB",X"25",X"26",X"B0",X"3E",X"FF",X"11",X"41",X"00",X"19",
		X"77",X"CD",X"14",X"4A",X"2A",X"5E",X"B0",X"26",X"09",X"22",X"62",X"B0",X"2A",X"5E",X"B4",X"2E",
		X"83",X"7C",X"C6",X"10",X"67",X"22",X"62",X"B4",X"3E",X"20",X"32",X"99",X"A8",X"3E",X"0A",X"CD",
		X"E2",X"3B",X"2A",X"5E",X"B0",X"26",X"9C",X"22",X"60",X"B0",X"2A",X"5E",X"B4",X"2E",X"09",X"22",
		X"60",X"B4",X"3E",X"04",X"32",X"96",X"A8",X"3E",X"FF",X"32",X"5F",X"B0",X"3E",X"00",X"32",X"A0",
		X"A8",X"D1",X"C1",X"DD",X"E1",X"C9",X"DD",X"21",X"20",X"A8",X"0E",X"00",X"DD",X"7E",X"00",X"FE",
		X"00",X"28",X"5F",X"C5",X"DD",X"E5",X"41",X"3E",X"0F",X"CD",X"F2",X"3C",X"DD",X"E1",X"C1",X"FE",
		X"00",X"CC",X"85",X"53",X"C5",X"DD",X"E5",X"41",X"3E",X"08",X"CD",X"F2",X"3C",X"DD",X"E1",X"C1",
		X"FE",X"00",X"20",X"3E",X"DD",X"7E",X"00",X"FE",X"02",X"20",X"06",X"CD",X"28",X"4A",X"C3",X"5E",
		X"54",X"CD",X"2D",X"4A",X"3E",X"05",X"CD",X"E2",X"3B",X"DD",X"7E",X"03",X"2F",X"47",X"3A",X"85",
		X"A8",X"80",X"38",X"07",X"3E",X"FF",X"32",X"8C",X"A8",X"3E",X"00",X"32",X"85",X"A8",X"CD",X"59",
		X"3D",X"3E",X"00",X"DD",X"77",X"00",X"69",X"CB",X"25",X"26",X"B0",X"3E",X"FF",X"11",X"41",X"00",
		X"19",X"77",X"11",X"08",X"00",X"DD",X"19",X"0C",X"79",X"FE",X"08",X"20",X"8F",X"C9",X"69",X"CB",
		X"25",X"26",X"B0",X"3E",X"FF",X"11",X"41",X"00",X"19",X"77",X"3E",X"32",X"CD",X"E2",X"3B",X"3E",
		X"00",X"DD",X"77",X"00",X"2A",X"50",X"B0",X"26",X"0A",X"22",X"62",X"B0",X"2A",X"50",X"B4",X"22",
		X"62",X"B4",X"3E",X"20",X"32",X"99",X"A8",X"DD",X"7E",X"03",X"CB",X"3F",X"47",X"3A",X"85",X"A8",
		X"80",X"30",X"02",X"3E",X"FF",X"32",X"85",X"A8",X"CD",X"59",X"3D",X"C3",X"52",X"54",X"3A",X"81",
		X"A8",X"FE",X"00",X"C0",X"21",X"03",X"A8",X"35",X"C0",X"3E",X"80",X"77",X"21",X"07",X"A8",X"35",
		X"20",X"13",X"3A",X"04",X"A8",X"77",X"2A",X"14",X"A8",X"22",X"19",X"A8",X"7C",X"FE",X"FF",X"28",
		X"04",X"CD",X"27",X"56",X"C9",X"21",X"06",X"A8",X"35",X"C0",X"3A",X"05",X"A8",X"77",X"2A",X"16",
		X"A8",X"22",X"19",X"A8",X"7C",X"FE",X"FF",X"C8",X"C3",X"27",X"56",X"21",X"40",X"B0",X"11",X"41",
		X"B4",X"DD",X"21",X"20",X"A8",X"06",X"08",X"DD",X"7E",X"00",X"FE",X"00",X"C4",X"FD",X"54",X"23",
		X"23",X"13",X"13",X"C5",X"01",X"08",X"00",X"DD",X"09",X"C1",X"10",X"EB",X"C9",X"FE",X"02",X"20",
		X"19",X"3A",X"B4",X"A8",X"E6",X"E0",X"20",X"0D",X"3A",X"B4",X"A8",X"CB",X"3F",X"E6",X"01",X"20",
		X"04",X"3E",X"02",X"18",X"02",X"3E",X"22",X"1B",X"12",X"13",X"DD",X"35",X"05",X"20",X"0C",X"3E",
		X"08",X"DD",X"77",X"05",X"23",X"7E",X"3C",X"E6",X"03",X"77",X"2B",X"3E",X"FF",X"32",X"91",X"A8",
		X"DD",X"35",X"04",X"C0",X"DD",X"7E",X"02",X"DD",X"77",X"04",X"DD",X"7E",X"01",X"FE",X"00",X"20",
		X"04",X"34",X"C3",X"5A",X"55",X"FE",X"01",X"20",X"06",X"1A",X"3D",X"12",X"C3",X"5A",X"55",X"FE",
		X"02",X"20",X"04",X"35",X"C3",X"5A",X"55",X"1A",X"3C",X"12",X"1A",X"E6",X"07",X"FE",X"04",X"C0",
		X"7E",X"E6",X"07",X"FE",X"04",X"C0",X"E5",X"C5",X"D5",X"DD",X"E5",X"46",X"1A",X"4F",X"CD",X"68",
		X"40",X"22",X"94",X"A8",X"3E",X"00",X"32",X"91",X"A8",X"7E",X"32",X"90",X"A8",X"CD",X"A6",X"40",
		X"DD",X"E1",X"DD",X"46",X"01",X"DD",X"E5",X"CD",X"93",X"55",X"DD",X"E1",X"DD",X"77",X"01",X"D1",
		X"C1",X"E1",X"C9",X"57",X"58",X"68",X"26",X"00",X"01",X"15",X"56",X"09",X"7E",X"A2",X"20",X"03",
		X"C3",X"C4",X"55",X"CD",X"93",X"40",X"E6",X"01",X"28",X"02",X"7B",X"C9",X"7B",X"3D",X"E6",X"03",
		X"6F",X"26",X"00",X"09",X"7E",X"A2",X"20",X"0C",X"7B",X"3C",X"E6",X"03",X"6F",X"26",X"00",X"09",
		X"7E",X"A2",X"28",X"E6",X"CD",X"93",X"40",X"E6",X"01",X"28",X"11",X"7B",X"3D",X"E6",X"03",X"6F",
		X"26",X"00",X"09",X"7E",X"A2",X"28",X"16",X"7B",X"3D",X"E6",X"03",X"C9",X"7B",X"3C",X"E6",X"03",
		X"6F",X"26",X"00",X"09",X"7E",X"A2",X"28",X"16",X"7B",X"3C",X"E6",X"03",X"C9",X"7B",X"3C",X"E6",
		X"03",X"6F",X"26",X"00",X"09",X"7E",X"A2",X"28",X"16",X"7B",X"3C",X"E6",X"03",X"C9",X"7B",X"3D",
		X"E6",X"03",X"6F",X"26",X"00",X"09",X"7E",X"A2",X"28",X"05",X"7B",X"3D",X"E6",X"03",X"C9",X"7B",
		X"3D",X"3D",X"E6",X"03",X"C9",X"01",X"04",X"02",X"08",X"21",X"20",X"A8",X"11",X"21",X"A8",X"36",
		X"00",X"01",X"3F",X"00",X"ED",X"B0",X"C9",X"E5",X"D5",X"C5",X"DD",X"E5",X"21",X"20",X"A8",X"0E",
		X"00",X"7E",X"FE",X"00",X"28",X"15",X"0C",X"11",X"08",X"00",X"19",X"3A",X"87",X"A8",X"47",X"79",
		X"B8",X"20",X"EE",X"3E",X"FF",X"DD",X"E1",X"C1",X"D1",X"E1",X"C9",X"CD",X"F6",X"49",X"E5",X"DD",
		X"E1",X"C5",X"3E",X"01",X"DD",X"77",X"00",X"3E",X"03",X"DD",X"77",X"01",X"3E",X"01",X"DD",X"77",
		X"04",X"DD",X"77",X"05",X"3A",X"18",X"A8",X"4F",X"06",X"00",X"CB",X"21",X"CB",X"10",X"21",X"D1",
		X"56",X"09",X"7E",X"DD",X"77",X"02",X"23",X"7E",X"DD",X"77",X"03",X"C1",X"CB",X"21",X"06",X"00",
		X"21",X"40",X"B0",X"09",X"E5",X"01",X"00",X"04",X"09",X"D1",X"3A",X"19",X"A8",X"12",X"3E",X"35",
		X"77",X"23",X"13",X"3A",X"1A",X"A8",X"77",X"3E",X"00",X"12",X"3A",X"19",X"A8",X"C6",X"04",X"32",
		X"52",X"B0",X"32",X"54",X"B0",X"3A",X"1A",X"A8",X"D6",X"14",X"32",X"53",X"B4",X"C6",X"10",X"32",
		X"55",X"B4",X"3E",X"09",X"32",X"52",X"B4",X"32",X"54",X"B4",X"3E",X"90",X"32",X"53",X"B0",X"3E",
		X"91",X"32",X"55",X"B0",X"3E",X"03",X"32",X"1B",X"A8",X"DD",X"E1",X"C1",X"D1",X"E1",X"3E",X"00",
		X"C9",X"18",X"20",X"18",X"20",X"14",X"28",X"14",X"30",X"10",X"30",X"10",X"30",X"0C",X"30",X"0C",
		X"40",X"0A",X"40",X"0A",X"40",X"08",X"40",X"08",X"40",X"08",X"40",X"08",X"40",X"08",X"40",X"08",
		X"40",X"04",X"40",X"04",X"40",X"04",X"40",X"04",X"40",X"04",X"40",X"04",X"40",X"04",X"40",X"04",
		X"40",X"0A",X"40",X"0A",X"40",X"0A",X"40",X"0A",X"40",X"08",X"40",X"08",X"40",X"08",X"40",X"08",
		X"40",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
