library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity cmd_snd_rom is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of cmd_snd_rom is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"F3",X"C3",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F5",X"DD",X"E5",X"E5",X"C5",X"D5",X"FD",X"E5",
		X"00",X"00",X"00",X"CD",X"46",X"01",X"CD",X"32",X"03",X"CD",X"F9",X"05",X"FD",X"E1",X"D1",X"C1",
		X"E1",X"DD",X"E1",X"F1",X"FB",X"ED",X"4D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"21",X"00",X"20",X"11",X"01",X"20",X"01",X"FF",X"03",X"36",X"00",X"ED",X"B0",X"31",X"FF",X"23",
		X"DD",X"21",X"67",X"06",X"0E",X"10",X"16",X"00",X"7A",X"DD",X"46",X"00",X"CD",X"57",X"06",X"DD",
		X"23",X"14",X"0D",X"C2",X"18",X"01",X"DD",X"21",X"67",X"06",X"16",X"00",X"0E",X"10",X"7A",X"DD",
		X"46",X"00",X"CD",X"5F",X"06",X"DD",X"23",X"14",X"0D",X"C2",X"2E",X"01",X"FB",X"00",X"CD",X"86",
		X"01",X"00",X"00",X"C3",X"3D",X"01",X"3E",X"0E",X"CD",X"49",X"06",X"CB",X"7F",X"C2",X"59",X"01",
		X"26",X"00",X"6F",X"22",X"00",X"20",X"C3",X"75",X"01",X"CB",X"BF",X"67",X"2E",X"00",X"CB",X"3C",
		X"CB",X"1D",X"CB",X"3C",X"CB",X"1D",X"CB",X"3C",X"CB",X"1D",X"CB",X"3C",X"CB",X"1D",X"CB",X"3C",
		X"CB",X"1D",X"22",X"00",X"20",X"DD",X"21",X"02",X"20",X"DD",X"34",X"07",X"DD",X"34",X"0F",X"DD",
		X"34",X"17",X"DD",X"34",X"2F",X"C9",X"ED",X"5B",X"00",X"20",X"21",X"00",X"00",X"22",X"00",X"20",
		X"CB",X"43",X"C2",X"F7",X"01",X"CB",X"3A",X"CB",X"1B",X"CB",X"43",X"C2",X"86",X"02",X"CB",X"3A",
		X"CB",X"1B",X"CB",X"43",X"C2",X"3C",X"02",X"3A",X"33",X"20",X"A7",X"C0",X"CB",X"3A",X"CB",X"1B",
		X"0E",X"07",X"DD",X"21",X"87",X"06",X"CB",X"43",X"C4",X"C8",X"02",X"CB",X"3A",X"CB",X"1B",X"DD",
		X"23",X"DD",X"23",X"DD",X"23",X"DD",X"23",X"0D",X"C2",X"B6",X"01",X"DD",X"21",X"02",X"20",X"CD",
		X"E8",X"01",X"DD",X"21",X"0A",X"20",X"CD",X"E8",X"01",X"DD",X"21",X"12",X"20",X"CD",X"E8",X"01",
		X"DD",X"21",X"2A",X"20",X"CD",X"E8",X"01",X"C9",X"DD",X"7E",X"07",X"FE",X"20",X"D8",X"DD",X"36",
		X"07",X"00",X"DD",X"36",X"00",X"0F",X"C9",X"3E",X"0F",X"32",X"02",X"20",X"32",X"0A",X"20",X"32",
		X"12",X"20",X"32",X"1A",X"20",X"32",X"22",X"20",X"32",X"2A",X"20",X"DD",X"21",X"67",X"06",X"0E",
		X"10",X"16",X"00",X"7A",X"DD",X"46",X"00",X"CD",X"57",X"06",X"DD",X"23",X"14",X"0D",X"C2",X"13",
		X"02",X"DD",X"21",X"67",X"06",X"16",X"00",X"0E",X"10",X"7A",X"DD",X"46",X"00",X"CD",X"5F",X"06",
		X"DD",X"23",X"14",X"0D",X"C2",X"29",X"02",X"AF",X"32",X"33",X"20",X"C9",X"AF",X"32",X"02",X"20",
		X"32",X"0A",X"20",X"32",X"12",X"20",X"32",X"1A",X"20",X"32",X"22",X"20",X"32",X"2A",X"20",X"3A",
		X"33",X"20",X"A7",X"C0",X"3E",X"FF",X"32",X"33",X"20",X"DD",X"21",X"77",X"06",X"16",X"00",X"0E",
		X"10",X"7A",X"DD",X"46",X"00",X"CD",X"57",X"06",X"DD",X"23",X"14",X"0D",X"C2",X"61",X"02",X"DD",
		X"21",X"67",X"06",X"16",X"00",X"0E",X"10",X"7A",X"DD",X"46",X"00",X"CD",X"5F",X"06",X"DD",X"23",
		X"14",X"0D",X"C2",X"77",X"02",X"C9",X"3A",X"1A",X"20",X"A7",X"C0",X"DD",X"21",X"1A",X"20",X"DD",
		X"36",X"00",X"FF",X"DD",X"36",X"01",X"01",X"DD",X"36",X"02",X"00",X"21",X"7A",X"08",X"DD",X"75",
		X"03",X"DD",X"74",X"04",X"DD",X"36",X"05",X"00",X"DD",X"21",X"22",X"20",X"DD",X"36",X"00",X"FF",
		X"DD",X"36",X"01",X"01",X"DD",X"36",X"02",X"00",X"21",X"C6",X"09",X"DD",X"75",X"03",X"DD",X"74",
		X"04",X"DD",X"36",X"05",X"01",X"C3",X"AC",X"01",X"DD",X"7E",X"02",X"FE",X"03",X"CA",X"E1",X"02",
		X"FE",X"00",X"CA",X"E8",X"02",X"FE",X"01",X"CA",X"EF",X"02",X"FD",X"21",X"12",X"20",X"C3",X"F3",
		X"02",X"FD",X"21",X"2A",X"20",X"C3",X"F3",X"02",X"FD",X"21",X"02",X"20",X"C3",X"F3",X"02",X"FD",
		X"21",X"0A",X"20",X"FD",X"7E",X"00",X"A7",X"CA",X"04",X"03",X"DD",X"7E",X"03",X"FD",X"BE",X"05",
		X"CA",X"2D",X"03",X"D0",X"FD",X"36",X"00",X"FF",X"FD",X"36",X"01",X"01",X"FD",X"36",X"02",X"00",
		X"FD",X"36",X"07",X"00",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"FD",X"75",X"03",X"FD",X"74",X"04",
		X"DD",X"7E",X"03",X"FD",X"77",X"05",X"DD",X"7E",X"02",X"FD",X"77",X"06",X"C9",X"FD",X"36",X"07",
		X"00",X"C9",X"CD",X"52",X"03",X"DD",X"21",X"2A",X"20",X"CD",X"32",X"04",X"DD",X"21",X"02",X"20",
		X"CD",X"32",X"04",X"DD",X"21",X"0A",X"20",X"CD",X"32",X"04",X"DD",X"21",X"12",X"20",X"CD",X"32",
		X"04",X"C9",X"3A",X"32",X"20",X"3C",X"32",X"32",X"20",X"FE",X"01",X"C0",X"AF",X"32",X"32",X"20",
		X"DD",X"21",X"1A",X"20",X"CD",X"6F",X"03",X"DD",X"21",X"22",X"20",X"CD",X"6F",X"03",X"C9",X"DD",
		X"7E",X"00",X"A7",X"C8",X"FE",X"0F",X"CA",X"08",X"04",X"DD",X"7E",X"01",X"3D",X"DD",X"77",X"01",
		X"C0",X"DD",X"6E",X"03",X"DD",X"66",X"04",X"DD",X"4E",X"02",X"DD",X"34",X"02",X"06",X"00",X"CB",
		X"21",X"CB",X"10",X"CB",X"21",X"CB",X"10",X"09",X"E5",X"FD",X"E1",X"FD",X"7E",X"00",X"FE",X"FF",
		X"CA",X"C2",X"03",X"DD",X"77",X"01",X"DD",X"7E",X"05",X"FE",X"00",X"CA",X"CB",X"03",X"FE",X"01",
		X"CA",X"DA",X"03",X"16",X"04",X"3E",X"07",X"CD",X"49",X"06",X"CB",X"97",X"CB",X"EF",X"4F",X"C3",
		X"E6",X"03",X"DD",X"36",X"02",X"00",X"DD",X"36",X"01",X"01",X"C9",X"16",X"00",X"3E",X"07",X"CD",
		X"49",X"06",X"CB",X"87",X"CB",X"DF",X"4F",X"C3",X"E6",X"03",X"16",X"02",X"3E",X"07",X"CD",X"49",
		X"06",X"CB",X"8F",X"CB",X"E7",X"4F",X"7A",X"FD",X"46",X"01",X"CD",X"57",X"06",X"7A",X"C6",X"01",
		X"FD",X"46",X"02",X"CD",X"57",X"06",X"7A",X"CB",X"3F",X"C6",X"08",X"FD",X"46",X"03",X"CD",X"57",
		X"06",X"3E",X"07",X"41",X"CD",X"57",X"06",X"C9",X"3E",X"07",X"CD",X"49",X"06",X"4F",X"DD",X"7E",
		X"05",X"FE",X"00",X"CA",X"20",X"04",X"FE",X"01",X"CA",X"25",X"04",X"CB",X"D1",X"C3",X"27",X"04",
		X"CB",X"C1",X"C3",X"27",X"04",X"CB",X"C9",X"3E",X"07",X"41",X"CD",X"57",X"06",X"DD",X"36",X"00",
		X"00",X"C9",X"DD",X"7E",X"00",X"A7",X"C8",X"FE",X"0F",X"CA",X"42",X"05",X"DD",X"7E",X"01",X"3D",
		X"DD",X"77",X"01",X"C0",X"DD",X"4E",X"02",X"DD",X"34",X"02",X"06",X"00",X"21",X"00",X"00",X"09",
		X"09",X"09",X"09",X"09",X"09",X"DD",X"4E",X"03",X"DD",X"46",X"04",X"09",X"E5",X"FD",X"E1",X"FD",
		X"7E",X"00",X"FE",X"FF",X"CA",X"9A",X"04",X"FE",X"FE",X"CA",X"9F",X"04",X"DD",X"77",X"01",X"FD",
		X"5E",X"01",X"3E",X"07",X"CD",X"50",X"06",X"47",X"DD",X"7E",X"06",X"FE",X"03",X"CA",X"8A",X"05",
		X"FE",X"00",X"CA",X"A8",X"04",X"FE",X"01",X"CA",X"B8",X"04",X"16",X"04",X"CB",X"4B",X"C4",X"DC",
		X"04",X"CB",X"53",X"C4",X"E1",X"04",X"48",X"C3",X"E6",X"04",X"DD",X"36",X"00",X"0F",X"C9",X"DD",
		X"36",X"02",X"00",X"DD",X"36",X"01",X"01",X"C9",X"16",X"00",X"CB",X"4B",X"C4",X"C8",X"04",X"CB",
		X"53",X"C4",X"CD",X"04",X"48",X"C3",X"E6",X"04",X"16",X"02",X"CB",X"4B",X"C4",X"D2",X"04",X"CB",
		X"53",X"C4",X"D7",X"04",X"48",X"C3",X"E6",X"04",X"CB",X"80",X"CB",X"D8",X"C9",X"CB",X"98",X"CB",
		X"C0",X"C9",X"CB",X"88",X"CB",X"E0",X"C9",X"CB",X"A0",X"CB",X"C8",X"C9",X"CB",X"90",X"CB",X"E8",
		X"C9",X"CB",X"A8",X"CB",X"D0",X"C9",X"CB",X"43",X"C2",X"15",X"05",X"7A",X"FD",X"46",X"02",X"CD",
		X"5F",X"06",X"7A",X"C6",X"01",X"FD",X"46",X"03",X"CD",X"5F",X"06",X"3E",X"06",X"FD",X"46",X"04",
		X"CD",X"5F",X"06",X"7A",X"CB",X"3F",X"C6",X"08",X"FD",X"46",X"05",X"CD",X"5F",X"06",X"3E",X"07",
		X"41",X"CD",X"5F",X"06",X"C9",X"3E",X"0B",X"FD",X"46",X"02",X"CD",X"5F",X"06",X"3E",X"0C",X"FD",
		X"46",X"03",X"CD",X"5F",X"06",X"3E",X"06",X"FD",X"46",X"04",X"CD",X"5F",X"06",X"7A",X"CB",X"3F",
		X"C6",X"08",X"06",X"10",X"CD",X"5F",X"06",X"3E",X"0D",X"FD",X"46",X"05",X"CD",X"5F",X"06",X"C3",
		X"0E",X"05",X"3E",X"07",X"CD",X"50",X"06",X"47",X"DD",X"7E",X"06",X"FE",X"03",X"CA",X"76",X"05",
		X"FE",X"00",X"CA",X"61",X"05",X"FE",X"01",X"CA",X"68",X"05",X"CB",X"D0",X"CB",X"E8",X"C3",X"6C",
		X"05",X"CB",X"C0",X"CB",X"D8",X"C3",X"6C",X"05",X"CB",X"C8",X"CB",X"D0",X"3E",X"07",X"CD",X"5F",
		X"06",X"AF",X"DD",X"77",X"00",X"C9",X"3E",X"07",X"CD",X"49",X"06",X"CB",X"D7",X"CB",X"EF",X"47",
		X"3E",X"07",X"CD",X"57",X"06",X"DD",X"36",X"00",X"00",X"C9",X"3E",X"07",X"CD",X"49",X"06",X"47",
		X"16",X"04",X"CB",X"4B",X"C4",X"DC",X"04",X"CB",X"53",X"C4",X"E1",X"04",X"48",X"CB",X"43",X"C2",
		X"CC",X"05",X"7A",X"FD",X"46",X"02",X"CD",X"57",X"06",X"7A",X"C6",X"01",X"FD",X"46",X"03",X"CD",
		X"57",X"06",X"3E",X"06",X"FD",X"46",X"04",X"CD",X"57",X"06",X"7A",X"CB",X"3F",X"C6",X"08",X"FD",
		X"46",X"05",X"CD",X"57",X"06",X"3E",X"07",X"41",X"CD",X"57",X"06",X"C9",X"3E",X"0B",X"FD",X"46",
		X"02",X"CD",X"57",X"06",X"3E",X"0C",X"FD",X"46",X"03",X"CD",X"57",X"06",X"3E",X"06",X"FD",X"46",
		X"04",X"CD",X"57",X"06",X"7A",X"CB",X"3F",X"C6",X"08",X"06",X"10",X"CD",X"57",X"06",X"3E",X"0D",
		X"FD",X"46",X"05",X"CD",X"57",X"06",X"C3",X"C5",X"05",X"3A",X"33",X"20",X"A7",X"C8",X"3D",X"32",
		X"33",X"20",X"FE",X"04",X"D0",X"AF",X"32",X"33",X"20",X"3A",X"1A",X"20",X"A7",X"C0",X"DD",X"21",
		X"1A",X"20",X"DD",X"36",X"00",X"FF",X"DD",X"36",X"01",X"01",X"DD",X"36",X"02",X"00",X"21",X"7A",
		X"08",X"DD",X"75",X"03",X"DD",X"74",X"04",X"DD",X"36",X"05",X"00",X"DD",X"21",X"22",X"20",X"DD",
		X"36",X"00",X"FF",X"DD",X"36",X"01",X"01",X"DD",X"36",X"02",X"00",X"21",X"C6",X"09",X"DD",X"75",
		X"03",X"DD",X"74",X"04",X"DD",X"36",X"05",X"01",X"C9",X"32",X"00",X"50",X"3A",X"00",X"40",X"C9",
		X"32",X"00",X"70",X"3A",X"00",X"60",X"C9",X"32",X"00",X"50",X"78",X"32",X"00",X"40",X"C9",X"32",
		X"00",X"70",X"78",X"32",X"00",X"60",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"37",X"10",
		X"00",X"00",X"00",X"60",X"09",X"00",X"00",X"A7",X"06",X"02",X"04",X"03",X"07",X"00",X"05",X"CB",
		X"06",X"03",X"06",X"FB",X"06",X"00",X"07",X"7C",X"07",X"01",X"08",X"0B",X"07",X"01",X"09",X"49",
		X"07",X"00",X"0A",X"49",X"07",X"00",X"0A",X"04",X"02",X"F0",X"00",X"00",X"0E",X"02",X"02",X"A0",
		X"00",X"00",X"0E",X"02",X"02",X"90",X"00",X"00",X"0E",X"02",X"02",X"80",X"00",X"00",X"0E",X"02",
		X"02",X"70",X"00",X"00",X"0E",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"02",X"02",X"F0",X"00",X"00",
		X"0E",X"02",X"02",X"00",X"00",X"00",X"00",X"02",X"02",X"F0",X"00",X"00",X"0E",X"02",X"02",X"00",
		X"00",X"00",X"0E",X"02",X"02",X"F0",X"00",X"00",X"0E",X"02",X"02",X"00",X"00",X"00",X"00",X"02",
		X"02",X"F0",X"00",X"00",X"0E",X"02",X"02",X"00",X"00",X"00",X"00",X"20",X"05",X"00",X"10",X"07",
		X"09",X"FF",X"FF",X"20",X"05",X"00",X"20",X"0F",X"09",X"0F",X"0F",X"02",X"02",X"00",X"02",X"00",
		X"0F",X"02",X"02",X"00",X"00",X"00",X"00",X"02",X"02",X"80",X"01",X"00",X"0F",X"02",X"02",X"40",
		X"01",X"00",X"0F",X"02",X"02",X"00",X"00",X"00",X"00",X"02",X"02",X"20",X"01",X"00",X"0F",X"02",
		X"02",X"00",X"00",X"00",X"00",X"02",X"00",X"10",X"00",X"00",X"0F",X"05",X"02",X"E0",X"00",X"00",
		X"0F",X"05",X"02",X"20",X"01",X"00",X"0F",X"FF",X"FF",X"05",X"02",X"00",X"02",X"00",X"0C",X"02",
		X"00",X"00",X"00",X"00",X"00",X"05",X"02",X"00",X"01",X"00",X"0C",X"02",X"00",X"00",X"00",X"00",
		X"00",X"05",X"02",X"00",X"02",X"00",X"0C",X"02",X"00",X"00",X"00",X"00",X"00",X"05",X"02",X"00",
		X"01",X"00",X"0C",X"02",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"08",X"02",X"00",X"01",
		X"00",X"0E",X"08",X"02",X"08",X"01",X"00",X"0E",X"08",X"02",X"10",X"01",X"00",X"0E",X"08",X"02",
		X"18",X"01",X"00",X"0E",X"08",X"02",X"20",X"01",X"00",X"0E",X"08",X"02",X"28",X"01",X"00",X"0E",
		X"08",X"02",X"30",X"01",X"00",X"0E",X"08",X"02",X"38",X"01",X"00",X"0E",X"08",X"02",X"40",X"01",
		X"00",X"0E",X"08",X"02",X"48",X"01",X"00",X"0E",X"08",X"02",X"50",X"01",X"00",X"0E",X"08",X"02",
		X"58",X"01",X"00",X"0E",X"08",X"02",X"60",X"01",X"00",X"0E",X"08",X"02",X"68",X"01",X"00",X"0E",
		X"08",X"02",X"70",X"01",X"00",X"0E",X"08",X"02",X"78",X"01",X"00",X"0E",X"08",X"02",X"80",X"01",
		X"00",X"0E",X"08",X"02",X"88",X"01",X"00",X"0E",X"08",X"02",X"90",X"01",X"00",X"0E",X"08",X"02",
		X"98",X"01",X"00",X"0E",X"08",X"02",X"A0",X"01",X"00",X"0E",X"08",X"02",X"A8",X"01",X"00",X"0E",
		X"08",X"02",X"B0",X"01",X"00",X"0E",X"08",X"02",X"B8",X"01",X"00",X"0E",X"08",X"02",X"C0",X"01",
		X"00",X"0E",X"08",X"02",X"C8",X"01",X"00",X"0E",X"08",X"02",X"D0",X"01",X"00",X"0E",X"08",X"02",
		X"D8",X"01",X"00",X"0E",X"08",X"02",X"E0",X"01",X"00",X"0E",X"08",X"02",X"E8",X"01",X"00",X"0E",
		X"08",X"02",X"F0",X"01",X"00",X"0E",X"08",X"02",X"F8",X"01",X"00",X"0E",X"08",X"02",X"00",X"02",
		X"00",X"0E",X"08",X"02",X"08",X"02",X"00",X"0E",X"08",X"02",X"10",X"02",X"00",X"0E",X"08",X"02",
		X"18",X"02",X"00",X"0E",X"08",X"02",X"20",X"02",X"00",X"0E",X"08",X"02",X"28",X"02",X"00",X"0E",
		X"08",X"02",X"30",X"02",X"00",X"0E",X"08",X"02",X"38",X"02",X"00",X"0E",X"08",X"02",X"40",X"02",
		X"00",X"0E",X"08",X"02",X"48",X"02",X"00",X"0E",X"FF",X"FF",X"0A",X"8F",X"00",X"09",X"02",X"01",
		X"00",X"00",X"0A",X"AA",X"00",X"09",X"26",X"01",X"00",X"00",X"0B",X"AA",X"00",X"09",X"01",X"01",
		X"00",X"00",X"0B",X"A0",X"00",X"09",X"01",X"01",X"00",X"00",X"0B",X"8F",X"00",X"09",X"01",X"01",
		X"00",X"00",X"0A",X"55",X"00",X"09",X"0E",X"01",X"00",X"00",X"0A",X"55",X"00",X"09",X"0E",X"01",
		X"00",X"00",X"23",X"6B",X"00",X"09",X"0D",X"01",X"00",X"00",X"0A",X"8F",X"00",X"09",X"02",X"01",
		X"00",X"00",X"0A",X"AA",X"00",X"09",X"26",X"01",X"00",X"00",X"0B",X"AA",X"00",X"09",X"01",X"01",
		X"00",X"00",X"0B",X"A0",X"00",X"09",X"01",X"01",X"00",X"00",X"0B",X"AA",X"00",X"09",X"01",X"01",
		X"00",X"00",X"0A",X"8F",X"00",X"09",X"0E",X"01",X"00",X"00",X"0A",X"8F",X"00",X"09",X"0E",X"01",
		X"00",X"00",X"23",X"A0",X"00",X"09",X"0D",X"01",X"00",X"00",X"0A",X"A0",X"00",X"09",X"02",X"01",
		X"00",X"00",X"0A",X"BE",X"00",X"09",X"26",X"01",X"00",X"00",X"0B",X"BE",X"00",X"09",X"01",X"01",
		X"00",X"00",X"0B",X"AA",X"00",X"09",X"01",X"01",X"00",X"00",X"0B",X"A0",X"00",X"09",X"01",X"01",
		X"00",X"00",X"0A",X"8F",X"00",X"09",X"02",X"01",X"00",X"00",X"0A",X"AA",X"00",X"09",X"26",X"01",
		X"00",X"00",X"0B",X"AA",X"00",X"09",X"01",X"01",X"00",X"00",X"0B",X"97",X"00",X"09",X"01",X"01",
		X"00",X"00",X"0B",X"AA",X"00",X"09",X"01",X"01",X"00",X"00",X"0B",X"BE",X"00",X"09",X"01",X"01",
		X"00",X"00",X"17",X"8F",X"00",X"09",X"01",X"01",X"00",X"00",X"0B",X"AA",X"00",X"09",X"01",X"01",
		X"00",X"00",X"0B",X"97",X"00",X"09",X"01",X"01",X"00",X"00",X"0A",X"BE",X"00",X"09",X"0E",X"01",
		X"00",X"00",X"0B",X"7F",X"00",X"09",X"01",X"01",X"00",X"00",X"11",X"8F",X"00",X"09",X"01",X"01",
		X"00",X"00",X"05",X"97",X"00",X"09",X"01",X"01",X"00",X"00",X"0B",X"8F",X"00",X"09",X"01",X"01",
		X"00",X"00",X"0B",X"7F",X"00",X"09",X"01",X"01",X"00",X"00",X"0B",X"8F",X"00",X"09",X"01",X"01",
		X"00",X"00",X"0B",X"A0",X"00",X"09",X"01",X"01",X"00",X"00",X"0B",X"AA",X"00",X"09",X"01",X"01",
		X"00",X"00",X"0B",X"BE",X"00",X"09",X"01",X"01",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"23",X"53",X"01",X"08",X"01",X"01",X"00",X"00",X"0B",X"AC",
		X"01",X"08",X"01",X"01",X"00",X"00",X"23",X"53",X"01",X"08",X"01",X"01",X"00",X"00",X"0B",X"AC",
		X"01",X"08",X"01",X"01",X"00",X"00",X"17",X"1D",X"01",X"08",X"01",X"01",X"00",X"00",X"17",X"53",
		X"01",X"08",X"01",X"01",X"00",X"00",X"17",X"AC",X"01",X"08",X"19",X"01",X"00",X"00",X"23",X"53",
		X"01",X"08",X"01",X"01",X"00",X"00",X"0B",X"7D",X"01",X"08",X"01",X"01",X"00",X"00",X"23",X"53",
		X"01",X"08",X"01",X"01",X"00",X"00",X"0B",X"7D",X"01",X"08",X"01",X"01",X"00",X"00",X"17",X"FE",
		X"00",X"08",X"01",X"01",X"00",X"00",X"17",X"40",X"01",X"08",X"01",X"01",X"00",X"00",X"17",X"AC",
		X"01",X"08",X"19",X"01",X"00",X"00",X"0B",X"40",X"01",X"08",X"07",X"01",X"00",X"00",X"05",X"AC",
		X"01",X"08",X"01",X"01",X"00",X"00",X"17",X"AC",X"01",X"08",X"01",X"01",X"00",X"00",X"0B",X"40",
		X"01",X"08",X"07",X"01",X"00",X"00",X"05",X"AC",X"01",X"08",X"01",X"01",X"00",X"00",X"17",X"AC",
		X"01",X"08",X"01",X"01",X"00",X"00",X"0B",X"1D",X"01",X"08",X"07",X"01",X"00",X"00",X"05",X"AC",
		X"01",X"08",X"01",X"01",X"00",X"00",X"17",X"AC",X"01",X"08",X"01",X"01",X"00",X"00",X"0B",X"1D",
		X"01",X"08",X"07",X"01",X"00",X"00",X"05",X"AC",X"01",X"08",X"01",X"01",X"00",X"00",X"17",X"AC",
		X"01",X"08",X"01",X"01",X"00",X"00",X"17",X"1D",X"01",X"08",X"01",X"01",X"00",X"00",X"11",X"1D",
		X"01",X"08",X"01",X"01",X"00",X"00",X"05",X"FE",X"00",X"08",X"01",X"01",X"00",X"00",X"0B",X"1D",
		X"01",X"08",X"01",X"01",X"00",X"00",X"0B",X"53",X"01",X"08",X"01",X"01",X"00",X"00",X"0B",X"AC",
		X"01",X"08",X"01",X"01",X"00",X"00",X"0B",X"53",X"01",X"08",X"01",X"01",X"00",X"00",X"05",X"1D",
		X"01",X"08",X"07",X"01",X"00",X"00",X"05",X"1D",X"01",X"08",X"01",X"01",X"00",X"00",X"05",X"FE",
		X"00",X"08",X"01",X"01",X"00",X"00",X"05",X"1D",X"01",X"08",X"07",X"01",X"00",X"00",X"05",X"1D",
		X"01",X"08",X"01",X"01",X"00",X"00",X"05",X"FE",X"00",X"08",X"01",X"01",X"00",X"00",X"23",X"1D",
		X"01",X"08",X"0D",X"01",X"00",X"00",X"FF",X"53",X"01",X"08",X"01",X"01",X"00",X"00",X"0B",X"1D",
		X"01",X"07",X"0D",X"01",X"00",X"00",X"11",X"1D",X"01",X"07",X"01",X"01",X"00",X"00",X"05",X"FE",
		X"00",X"0A",X"01",X"01",X"00",X"00",X"0B",X"1D",X"01",X"07",X"01",X"01",X"00",X"00",X"0B",X"53",
		X"01",X"07",X"01",X"01",X"00",X"00",X"0B",X"AC",X"01",X"07",X"01",X"01",X"00",X"00",X"0B",X"53",
		X"01",X"07",X"01",X"01",X"00",X"00",X"05",X"1D",X"01",X"07",X"07",X"01",X"00",X"00",X"05",X"1D",
		X"01",X"07",X"01",X"01",X"00",X"00",X"05",X"FE",X"00",X"0A",X"01",X"01",X"00",X"00",X"05",X"1D",
		X"01",X"07",X"07",X"01",X"00",X"00",X"05",X"1D",X"01",X"07",X"01",X"01",X"00",X"00",X"05",X"FE",
		X"00",X"0A",X"01",X"01",X"00",X"00",X"23",X"1D",X"01",X"07",X"0D",X"01",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
