`define BUILD_DATE "190227"
`define BUILD_TIME "185900"
