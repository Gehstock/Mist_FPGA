library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_8R is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_8R is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"04",X"40",X"54",X"01",X"10",X"26",X"16",X"01",X"08",X"12",X"55",X"07",X"25",X"11",X"4C",X"00",
		X"C0",X"0D",X"58",X"15",X"11",X"05",X"86",X"00",X"45",X"29",X"54",X"10",X"42",X"01",X"00",X"00",
		X"4C",X"05",X"01",X"54",X"00",X"14",X"A5",X"14",X"4B",X"15",X"80",X"54",X"E0",X"45",X"10",X"14",
		X"42",X"D5",X"43",X"14",X"11",X"00",X"C0",X"00",X"65",X"00",X"10",X"15",X"40",X"41",X"00",X"00",
		X"76",X"DA",X"F6",X"EC",X"68",X"F6",X"7C",X"F1",X"B5",X"08",X"D0",X"10",X"88",X"20",X"42",X"08",
		X"48",X"F8",X"ED",X"DA",X"79",X"ED",X"7F",X"A2",X"00",X"02",X"00",X"10",X"02",X"40",X"00",X"42",
		X"78",X"E8",X"74",X"F2",X"78",X"E0",X"76",X"B9",X"46",X"00",X"05",X"6E",X"7F",X"06",X"27",X"00",
		X"70",X"D8",X"F0",X"C1",X"70",X"E4",X"60",X"F1",X"00",X"0C",X"85",X"D7",X"76",X"5F",X"03",X"13",
		X"84",X"D4",X"8A",X"CA",X"9A",X"1D",X"B4",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"6D",X"A5",X"4A",X"CA",X"84",X"71",X"6E",X"AC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7E",X"F5",X"FE",X"F9",X"76",X"BD",X"79",X"FC",X"84",X"12",X"08",X"07",X"8B",X"40",X"81",X"80",
		X"76",X"B8",X"5E",X"B9",X"3C",X"F9",X"76",X"FA",X"09",X"C0",X"00",X"03",X"A1",X"8B",X"40",X"90",
		X"FF",X"FD",X"7E",X"3D",X"58",X"DE",X"EA",X"A5",X"71",X"F3",X"FB",X"BF",X"7F",X"1F",X"17",X"0B",
		X"C9",X"3B",X"7F",X"FF",X"FF",X"7F",X"02",X"01",X"BC",X"FF",X"FF",X"F6",X"FC",X"FC",X"F6",X"0F",
		X"0B",X"84",X"90",X"15",X"B0",X"FE",X"FF",X"BC",X"07",X"82",X"A0",X"E8",X"FC",X"DD",X"5D",X"7F",
		X"E8",X"18",X"DF",X"DF",X"0F",X"07",X"01",X"9B",X"0E",X"A5",X"FE",X"FA",X"D0",X"84",X"C2",X"E0",
		X"04",X"40",X"54",X"01",X"10",X"26",X"16",X"01",X"08",X"12",X"55",X"07",X"25",X"11",X"4C",X"00",
		X"C0",X"0D",X"58",X"15",X"11",X"55",X"C6",X"40",X"45",X"29",X"54",X"10",X"42",X"01",X"0C",X"D5",
		X"40",X"11",X"55",X"10",X"C4",X"60",X"05",X"46",X"05",X"80",X"05",X"17",X"05",X"40",X"00",X"04",
		X"11",X"11",X"0C",X"40",X"31",X"54",X"11",X"41",X"10",X"35",X"11",X"00",X"41",X"04",X"40",X"04",
		X"F2",X"9C",X"61",X"36",X"33",X"DB",X"53",X"87",X"D7",X"BE",X"F8",X"F8",X"F0",X"A0",X"E0",X"90",
		X"7E",X"AF",X"5D",X"BE",X"7F",X"FE",X"FC",X"F5",X"D4",X"80",X"00",X"90",X"40",X"01",X"20",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"FF",X"4A",X"A0",X"D4",X"94",X"08",X"40",X"E4",X"30",
		X"FC",X"FE",X"FC",X"F8",X"F9",X"F9",X"C9",X"C9",X"50",X"08",X"04",X"44",X"12",X"80",X"20",X"48",
		X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FF",X"FF",X"BF",X"BF",X"BF",X"3F",X"80",X"BF",
		X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"BF",X"BF",X"3F",X"80",X"BF",X"BF",X"BF",X"3F",
		X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",
		X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",
		X"C9",X"C9",X"C9",X"C9",X"C9",X"C9",X"C9",X"C9",X"40",X"A0",X"34",X"44",X"A8",X"30",X"3A",X"60",
		X"C9",X"C9",X"C9",X"C9",X"C9",X"C9",X"C9",X"C9",X"50",X"10",X"A8",X"34",X"60",X"10",X"08",X"50",
		X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FF",X"80",X"BF",X"BF",X"BF",X"3F",X"80",X"BF",X"BF",
		X"E7",X"E0",X"E1",X"E0",X"E1",X"E8",X"E8",X"E9",X"BF",X"BF",X"83",X"01",X"01",X"1F",X"7F",X"3F",
		X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FB",X"E8",X"E9",X"E0",X"E8",X"E0",X"E1",X"E9",X"BF",X"1F",X"0F",X"0F",X"01",X"01",X"1F",X"3F",
		X"FC",X"E0",X"E9",X"E8",X"E8",X"E8",X"E0",X"EC",X"3F",X"3F",X"1F",X"0F",X"0F",X"0F",X"8F",X"BF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",
		X"E3",X"E3",X"E3",X"E3",X"E3",X"E3",X"E3",X"FB",X"BF",X"BF",X"3F",X"80",X"BF",X"BF",X"BF",X"3F",
		X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"80",X"BF",X"BF",X"BF",X"3F",X"80",X"BF",X"BF",
		X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",
		X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"BF",X"3F",X"80",X"BF",X"BF",X"BF",X"3F",X"80",
		X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"BF",X"BF",X"BF",X"3F",X"80",X"BF",X"BF",X"BF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FC",X"FC",X"F8",X"F8",X"F8",X"F0",X"F0",
		X"FB",X"FB",X"7B",X"7B",X"44",X"44",X"5C",X"44",X"3F",X"80",X"BF",X"3F",X"3F",X"3F",X"00",X"00",
		X"5C",X"44",X"5C",X"44",X"5C",X"44",X"5C",X"44",X"00",X"BF",X"BF",X"BF",X"3F",X"3F",X"00",X"00",
		X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"E0",X"E0",X"E0",X"C0",X"C0",X"C0",X"80",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"80",X"80",X"00",X"00",X"00",X"80",X"C8",X"F0",
		X"5C",X"44",X"5C",X"44",X"5C",X"44",X"5C",X"44",X"00",X"BF",X"BF",X"BF",X"3F",X"3F",X"00",X"00",
		X"5C",X"44",X"5C",X"44",X"5C",X"44",X"5C",X"44",X"00",X"BF",X"BF",X"BF",X"3F",X"3F",X"00",X"00",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"FC",X"FC",X"FC",X"FE",X"FE",X"FE",X"FF",X"FF",X"40",X"30",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"80",X"80",X"80",X"C0",X"C4",X"F8",X"F8",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"D0",X"D8",X"C8",X"E8",X"E8",X"F8",X"F8",X"F8",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FC",X"FA",X"F9",X"FD",X"FD",X"FF",X"FF",
		X"5C",X"44",X"5C",X"44",X"5C",X"44",X"5C",X"44",X"00",X"BF",X"BF",X"BF",X"3F",X"3F",X"00",X"00",
		X"5C",X"44",X"5C",X"44",X"5C",X"44",X"5C",X"44",X"00",X"BF",X"BF",X"BF",X"3F",X"3F",X"7F",X"FF",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"36",X"F6",X"F6",X"FE",X"FF",X"FF",X"FD",X"FE",X"48",X"A8",X"58",X"54",X"08",X"A8",X"E0",X"C0",
		X"FE",X"FF",X"FF",X"FE",X"FF",X"FF",X"FE",X"FF",X"54",X"8C",X"84",X"94",X"52",X"A8",X"26",X"54",
		X"CE",X"CE",X"F6",X"36",X"36",X"36",X"36",X"36",X"20",X"82",X"56",X"44",X"40",X"A8",X"50",X"44",
		X"36",X"36",X"36",X"36",X"36",X"36",X"36",X"36",X"A0",X"F0",X"24",X"B0",X"78",X"A8",X"28",X"54",
		X"36",X"36",X"36",X"36",X"36",X"36",X"36",X"36",X"48",X"A0",X"50",X"50",X"28",X"A8",X"64",X"58",
		X"36",X"36",X"36",X"36",X"36",X"36",X"36",X"36",X"10",X"A8",X"20",X"78",X"70",X"B8",X"34",X"54",
		X"25",X"10",X"A4",X"01",X"00",X"11",X"00",X"08",X"BF",X"52",X"01",X"02",X"D0",X"32",X"0C",X"23",
		X"20",X"82",X"10",X"09",X"80",X"00",X"20",X"04",X"41",X"02",X"48",X"02",X"40",X"21",X"02",X"26",
		X"FF",X"11",X"00",X"48",X"91",X"00",X"00",X"50",X"FF",X"84",X"4C",X"84",X"02",X"00",X"A4",X"00",
		X"81",X"70",X"1C",X"27",X"54",X"10",X"00",X"28",X"8C",X"00",X"80",X"A2",X"C4",X"74",X"9E",X"83",
		X"DF",X"30",X"08",X"11",X"00",X"B0",X"14",X"80",X"D7",X"94",X"20",X"12",X"20",X"10",X"14",X"40",
		X"54",X"11",X"08",X"10",X"00",X"14",X"10",X"30",X"B1",X"10",X"40",X"90",X"08",X"15",X"00",X"30",
		X"FF",X"18",X"52",X"04",X"14",X"10",X"10",X"2A",X"28",X"04",X"00",X"44",X"40",X"00",X"00",X"20",
		X"10",X"02",X"08",X"92",X"30",X"18",X"10",X"90",X"00",X"24",X"04",X"90",X"10",X"00",X"00",X"62",
		X"00",X"02",X"00",X"0A",X"24",X"80",X"00",X"80",X"20",X"12",X"4A",X"28",X"8C",X"12",X"9A",X"43",
		X"01",X"08",X"12",X"00",X"A0",X"00",X"00",X"01",X"00",X"3A",X"80",X"10",X"53",X"02",X"29",X"0B",
		X"88",X"41",X"28",X"10",X"48",X"4D",X"02",X"08",X"84",X"04",X"80",X"00",X"0C",X"84",X"80",X"05",
		X"85",X"08",X"50",X"00",X"48",X"40",X"09",X"50",X"80",X"C0",X"A4",X"00",X"0C",X"04",X"0A",X"14",
		X"D0",X"30",X"1E",X"43",X"00",X"00",X"10",X"18",X"40",X"04",X"40",X"41",X"A0",X"70",X"08",X"47",
		X"40",X"88",X"10",X"14",X"21",X"91",X"04",X"30",X"03",X"D0",X"00",X"40",X"24",X"40",X"40",X"01",
		X"10",X"10",X"00",X"90",X"04",X"90",X"01",X"30",X"00",X"02",X"00",X"40",X"00",X"00",X"02",X"10",
		X"D0",X"70",X"34",X"37",X"01",X"12",X"90",X"30",X"00",X"08",X"00",X"02",X"80",X"10",X"00",X"48",
		X"08",X"00",X"20",X"00",X"44",X"80",X"00",X"02",X"80",X"02",X"44",X"20",X"52",X"00",X"09",X"83",
		X"00",X"00",X"00",X"08",X"20",X"00",X"82",X"80",X"00",X"44",X"00",X"02",X"02",X"10",X"81",X"06",
		X"64",X"88",X"04",X"40",X"08",X"48",X"04",X"02",X"08",X"86",X"01",X"44",X"80",X"04",X"44",X"80",
		X"48",X"88",X"00",X"00",X"4A",X"04",X"49",X"80",X"A4",X"10",X"0D",X"84",X"84",X"20",X"04",X"84",
		X"90",X"44",X"20",X"30",X"18",X"04",X"13",X"10",X"28",X"20",X"40",X"60",X"02",X"20",X"20",X"10",
		X"00",X"30",X"04",X"18",X"10",X"00",X"80",X"50",X"80",X"60",X"20",X"14",X"20",X"24",X"42",X"23",
		X"80",X"18",X"10",X"24",X"28",X"00",X"08",X"40",X"80",X"00",X"40",X"40",X"22",X"24",X"06",X"03",
		X"00",X"06",X"04",X"00",X"87",X"00",X"20",X"00",X"01",X"CC",X"97",X"43",X"B1",X"C6",X"4B",X"21",
		X"21",X"10",X"00",X"00",X"84",X"00",X"40",X"08",X"25",X"00",X"12",X"44",X"10",X"21",X"04",X"00",
		X"00",X"00",X"02",X"00",X"24",X"01",X"00",X"40",X"89",X"08",X"02",X"20",X"05",X"01",X"04",X"50",
		X"20",X"80",X"40",X"00",X"23",X"08",X"84",X"18",X"A4",X"00",X"14",X"82",X"00",X"84",X"04",X"00",
		X"02",X"20",X"00",X"20",X"00",X"C2",X"08",X"02",X"88",X"40",X"05",X"00",X"80",X"46",X"01",X"01",
		X"00",X"98",X"50",X"20",X"00",X"92",X"18",X"09",X"B0",X"00",X"40",X"60",X"02",X"20",X"50",X"08",
		X"14",X"10",X"22",X"41",X"10",X"08",X"10",X"00",X"20",X"22",X"60",X"01",X"80",X"E0",X"4A",X"A1",
		X"A0",X"01",X"00",X"80",X"02",X"40",X"00",X"00",X"8F",X"11",X"C3",X"4F",X"13",X"27",X"09",X"42",
		X"00",X"89",X"80",X"40",X"00",X"00",X"80",X"00",X"38",X"11",X"C7",X"1F",X"21",X"03",X"37",X"48",
		X"02",X"00",X"80",X"10",X"00",X"00",X"80",X"00",X"12",X"00",X"00",X"00",X"21",X"10",X"04",X"01",
		X"00",X"00",X"02",X"20",X"00",X"00",X"00",X"44",X"00",X"00",X"08",X"02",X"00",X"41",X"04",X"00",
		X"04",X"A4",X"00",X"02",X"10",X"04",X"00",X"20",X"40",X"22",X"84",X"90",X"04",X"10",X"94",X"08",
		X"0A",X"02",X"80",X"24",X"00",X"20",X"40",X"09",X"00",X"24",X"46",X"00",X"82",X"54",X"88",X"21",
		X"90",X"B2",X"00",X"14",X"88",X"01",X"10",X"12",X"20",X"10",X"2A",X"28",X"44",X"46",X"22",X"21",
		X"00",X"80",X"90",X"0C",X"14",X"13",X"00",X"30",X"10",X"20",X"B4",X"01",X"21",X"40",X"22",X"20",
		X"80",X"00",X"00",X"24",X"60",X"00",X"08",X"C0",X"83",X"C7",X"74",X"29",X"13",X"82",X"54",X"11",
		X"00",X"40",X"00",X"00",X"80",X"00",X"20",X"82",X"0F",X"27",X"48",X"07",X"13",X"29",X"6F",X"87",
		X"00",X"80",X"00",X"00",X"00",X"80",X"08",X"00",X"01",X"12",X"80",X"01",X"24",X"82",X"08",X"01",
		X"80",X"00",X"00",X"08",X"42",X"00",X"00",X"00",X"00",X"04",X"00",X"04",X"01",X"00",X"00",X"08",
		X"02",X"08",X"51",X"00",X"2A",X"02",X"00",X"90",X"64",X"02",X"14",X"20",X"86",X"08",X"81",X"14",
		X"00",X"02",X"40",X"0C",X"80",X"01",X"04",X"19",X"62",X"01",X"82",X"0A",X"84",X"10",X"05",X"92",
		X"14",X"A2",X"10",X"01",X"70",X"10",X"A0",X"01",X"A0",X"00",X"44",X"20",X"A0",X"08",X"30",X"20",
		X"14",X"40",X"10",X"00",X"00",X"11",X"70",X"08",X"28",X"12",X"04",X"80",X"2A",X"21",X"51",X"08",
		X"50",X"A0",X"00",X"50",X"89",X"20",X"02",X"52",X"0A",X"47",X"47",X"8B",X"11",X"0F",X"8C",X"51",
		X"81",X"18",X"20",X"80",X"50",X"20",X"10",X"60",X"0B",X"CF",X"8F",X"1B",X"35",X"42",X"05",X"1F",
		X"00",X"80",X"00",X"80",X"00",X"02",X"80",X"00",X"24",X"00",X"00",X"02",X"00",X"08",X"00",X"41",
		X"04",X"20",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"02",X"10",X"08",X"01",X"01",X"04",
		X"04",X"40",X"08",X"20",X"01",X"40",X"02",X"00",X"00",X"10",X"82",X"00",X"00",X"04",X"42",X"00",
		X"08",X"00",X"00",X"00",X"20",X"00",X"02",X"00",X"40",X"02",X"88",X"00",X"00",X"11",X"02",X"80",
		X"0A",X"90",X"01",X"80",X"50",X"00",X"00",X"22",X"23",X"10",X"22",X"04",X"48",X"A3",X"00",X"08",
		X"41",X"14",X"02",X"00",X"10",X"20",X"02",X"04",X"52",X"10",X"22",X"02",X"95",X"00",X"04",X"0A",
		X"84",X"20",X"40",X"92",X"A0",X"00",X"00",X"50",X"00",X"01",X"03",X"87",X"94",X"09",X"07",X"03",
		X"00",X"00",X"A0",X"40",X"00",X"04",X"10",X"A0",X"07",X"04",X"29",X"43",X"07",X"04",X"08",X"41",
		X"E4",X"C0",X"E4",X"C1",X"D0",X"E6",X"F6",X"C1",X"08",X"12",X"55",X"07",X"21",X"11",X"48",X"00",
		X"C0",X"CD",X"F8",X"D5",X"D1",X"F5",X"C6",X"C0",X"45",X"29",X"50",X"10",X"46",X"01",X"0C",X"D5",
		X"80",X"91",X"D5",X"D0",X"C4",X"80",X"85",X"86",X"05",X"80",X"05",X"14",X"05",X"40",X"00",X"04",
		X"D1",X"D1",X"8C",X"C0",X"B1",X"94",X"91",X"C1",X"10",X"35",X"11",X"00",X"41",X"04",X"40",X"04",
		X"C4",X"85",X"C1",X"F4",X"80",X"80",X"E5",X"D4",X"43",X"15",X"80",X"44",X"40",X"41",X"10",X"14",
		X"C2",X"C1",X"C1",X"94",X"D1",X"80",X"C5",X"D1",X"45",X"00",X"10",X"11",X"44",X"50",X"15",X"05",
		X"84",X"C0",X"D4",X"81",X"90",X"E6",X"D6",X"81",X"08",X"12",X"55",X"07",X"25",X"11",X"4C",X"00",
		X"C0",X"CD",X"D8",X"95",X"D1",X"85",X"C4",X"E0",X"45",X"29",X"54",X"10",X"42",X"01",X"04",X"00",
		X"80",X"13",X"94",X"49",X"62",X"38",X"34",X"C3",X"D0",X"E9",X"50",X"E0",X"70",X"13",X"A0",X"D0",
		X"A9",X"47",X"E0",X"8B",X"C7",X"71",X"C8",X"F6",X"61",X"C0",X"94",X"61",X"D8",X"89",X"24",X"E1",
		X"00",X"08",X"07",X"03",X"00",X"40",X"05",X"03",X"01",X"93",X"40",X"62",X"3D",X"D8",X"84",X"70",
		X"10",X"11",X"0E",X"04",X"01",X"13",X"0A",X"00",X"F9",X"10",X"21",X"D0",X"F1",X"09",X"78",X"98",
		X"10",X"09",X"07",X"02",X"08",X"5E",X"13",X"2A",X"40",X"39",X"9D",X"06",X"9C",X"79",X"04",X"48",
		X"C7",X"71",X"0E",X"04",X"01",X"1A",X"78",X"84",X"BA",X"15",X"40",X"C1",X"21",X"09",X"78",X"88",
		X"CC",X"3B",X"94",X"49",X"62",X"B8",X"34",X"C3",X"D0",X"E8",X"50",X"E0",X"71",X"10",X"A0",X"D0",
		X"A9",X"47",X"E0",X"8B",X"C7",X"71",X"C8",X"F6",X"61",X"C0",X"94",X"60",X"D8",X"89",X"24",X"E1",
		X"D6",X"2B",X"94",X"48",X"E1",X"CA",X"14",X"C0",X"C0",X"68",X"01",X"D3",X"E1",X"37",X"83",X"27",
		X"A7",X"49",X"E1",X"8F",X"93",X"00",X"8B",X"F6",X"05",X"CB",X"0F",X"45",X"83",X"83",X"20",X"E8",
		X"FF",X"FF",X"FF",X"FD",X"FD",X"F7",X"F8",X"FF",X"FF",X"FF",X"CF",X"AF",X"CB",X"47",X"83",X"47",
		X"FF",X"F8",X"F7",X"FD",X"FB",X"FE",X"FD",X"FF",X"43",X"E3",X"A3",X"47",X"87",X"CF",X"DB",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"DA",X"EC",X"FF",X"FF",X"FF",X"FF",X"FF",X"5F",X"7F",X"1F",
		X"FE",X"FA",X"C7",X"FD",X"FA",X"FD",X"F6",X"EF",X"3F",X"1F",X"1F",X"1F",X"3F",X"3F",X"7F",X"DF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"82",X"BA",X"AA",X"B2",X"A2",X"BE",X"80",X"FE",X"82",X"BA",X"AA",X"B2",X"A2",X"BE",X"80",
		X"FE",X"82",X"BA",X"AA",X"B2",X"A2",X"BE",X"80",X"FE",X"82",X"BA",X"AA",X"B2",X"A2",X"BE",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"82",X"12",X"52",X"50",X"50",X"C0",X"C1",X"85",X"D6",X"F3",X"D5",X"D2",X"56",X"77",X"6D",X"7A",
		X"85",X"D5",X"D3",X"D2",X"52",X"42",X"42",X"43",X"5D",X"74",X"EC",X"E9",X"AC",X"EC",X"DB",X"F6",
		X"4E",X"0B",X"2B",X"79",X"F7",X"49",X"4B",X"6F",X"FB",X"FB",X"FA",X"FA",X"7E",X"77",X"67",X"75",
		X"6F",X"2F",X"AB",X"A2",X"92",X"B2",X"16",X"77",X"5D",X"7D",X"ED",X"F7",X"B7",X"F6",X"F6",X"F6",
		X"51",X"54",X"54",X"44",X"40",X"44",X"54",X"50",X"20",X"01",X"25",X"25",X"A1",X"81",X"91",X"85",
		X"50",X"50",X"54",X"55",X"45",X"45",X"41",X"40",X"A4",X"84",X"14",X"15",X"51",X"10",X"21",X"08",
		X"00",X"00",X"33",X"00",X"00",X"33",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"33",X"00",X"00",
		X"33",X"00",X"00",X"33",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"33",X"00",X"00",X"00",X"00",
		X"00",X"00",X"33",X"00",X"00",X"33",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"33",X"00",X"00",
		X"33",X"00",X"00",X"33",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"33",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"F0",X"FE",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"66",X"00",X"99",X"00",X"E6",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C0",X"F9",X"F0",X"FE",X"FC",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"00",X"66",X"00",X"99",X"00",X"66",X"FF",X"FF",X"00",X"66",X"00",X"99",X"00",X"66",
		X"00",X"99",X"00",X"66",X"00",X"99",X"00",X"FF",X"00",X"99",X"00",X"66",X"00",X"99",X"00",X"FF",
		X"FF",X"FF",X"00",X"00",X"11",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"11",X"00",X"00",X"00",
		X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",
		X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",
		X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"AA",X"AA",X"55",X"55",X"AA",X"FF",X"55",X"55",X"AA",X"AA",X"55",X"55",X"AA",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"AA",X"AA",X"D5",X"D5",X"EA",X"FF",X"55",X"55",X"AA",X"AA",X"55",X"55",X"AA",X"FF",
		X"FF",X"FF",X"6D",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"B6",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"0A",X"04",X"1F",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"80",X"C0",X"E0",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FF",X"FF",X"AE",X"BF",X"AA",X"BF",X"BF",X"BF",
		X"AA",X"AA",X"AA",X"00",X"80",X"C0",X"E0",X"FF",X"BF",X"AA",X"BA",X"10",X"1F",X"10",X"10",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"FF",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"FF",X"FF",X"FF",X"C3",X"C3",X"C2",X"C3",X"C3",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"C3",X"C3",X"C3",X"C3",X"C3",X"C3",X"C3",X"C3",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"C2",X"C3",X"C3",X"FF",X"FF",X"FF",X"FF",X"FF",X"C0",X"C0",X"C0",X"C0",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"00",
		X"00",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"00",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"00",
		X"FF",X"80",X"C0",X"E0",X"F0",X"F8",X"FC",X"FE",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"80",X"C0",X"E0",X"F0",X"F8",X"FC",X"FF",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"31",X"33",X"33",X"73",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"30",X"30",X"30",X"30",X"37",X"30",X"30",X"30",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"30",X"30",X"30",X"30",X"37",X"30",X"30",X"30",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"30",X"30",X"30",X"30",X"37",X"30",X"30",X"30",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"01",X"DC",X"F8",X"F8",X"7E",X"78",X"3C",X"32",X"C0",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FA",X"F0",X"28",X"F2",X"53",X"E4",X"47",X"D7",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"48",X"A0",X"14",X"D2",X"8A",X"28",X"20",X"50",
		X"FF",X"FE",X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"D4",X"A0",X"84",X"58",X"D0",X"80",X"A4",X"58",
		X"FF",X"FF",X"BF",X"77",X"78",X"ED",X"73",X"F9",X"FF",X"FF",X"BF",X"9E",X"3F",X"9E",X"4E",X"A5",
		X"73",X"A1",X"53",X"0C",X"C6",X"17",X"4A",X"54",X"CC",X"C6",X"B7",X"E2",X"A5",X"42",X"37",X"16",
		X"0F",X"55",X"93",X"39",X"9C",X"11",X"38",X"74",X"69",X"C2",X"EC",X"8A",X"D4",X"78",X"F4",X"7E",
		X"B0",X"38",X"14",X"38",X"9E",X"1C",X"48",X"02",X"3D",X"5C",X"BA",X"1E",X"2D",X"87",X"0E",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FE",X"FC",X"FC",X"F8",X"F0",X"F0",X"E2",X"01",X"03",X"07",X"07",X"87",X"2F",X"2F",X"7F",
		X"CF",X"BF",X"BF",X"BF",X"BE",X"BE",X"BC",X"BC",X"6B",X"F5",X"E1",X"C1",X"00",X"00",X"00",X"00",
		X"DF",X"FF",X"BF",X"FF",X"BF",X"FF",X"BF",X"FF",X"DC",X"EE",X"FB",X"7D",X"EE",X"DF",X"FA",X"EE",
		X"FF",X"BF",X"BF",X"FF",X"BF",X"F7",X"BE",X"BF",X"7D",X"DA",X"E6",X"BD",X"F7",X"FE",X"39",X"9F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"2A",X"FF",X"FF",X"FF",X"FF",X"EF",X"AB",X"AB",X"AF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"0F",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",X"F0",X"F6",X"92",
		X"FF",X"FF",X"FE",X"FC",X"FB",X"F7",X"F6",X"FE",X"70",X"70",X"79",X"F4",X"78",X"78",X"78",X"78",
		X"FF",X"FF",X"FF",X"FF",X"BC",X"1C",X"05",X"0C",X"FF",X"FF",X"F9",X"FC",X"78",X"38",X"30",X"50",
		X"0C",X"1E",X"07",X"03",X"30",X"41",X"27",X"1F",X"FC",X"D4",X"34",X"67",X"4E",X"CC",X"E4",X"E0",
		X"BE",X"9E",X"1C",X"1C",X"0C",X"18",X"18",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"F8",X"FF",X"FE",X"F1",X"E1",X"81",X"01",X"01",X"01",
		X"F0",X"C3",X"84",X"00",X"00",X"FC",X"FA",X"FC",X"00",X"80",X"00",X"00",X"00",X"04",X"08",X"0C",
		X"2A",X"6A",X"6A",X"6A",X"2A",X"2A",X"2A",X"00",X"BF",X"BF",X"BF",X"FF",X"FF",X"FC",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"08",
		X"03",X"07",X"07",X"06",X"00",X"00",X"00",X"00",X"FF",X"FF",X"F8",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EC",X"E4",X"0E",X"05",X"02",X"00",X"00",X"00",X"1A",X"4D",X"9D",X"0C",X"10",X"38",X"1D",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"0E",X"02",X"00",X"00",X"00",X"00",X"00",
		X"CB",X"2E",X"17",X"AE",X"0C",X"05",X"06",X"39",X"F0",X"EA",X"64",X"F4",X"E0",X"60",X"A0",X"62",
		X"93",X"0A",X"89",X"08",X"1B",X"38",X"99",X"19",X"82",X"EA",X"A2",X"92",X"48",X"C0",X"C0",X"A2",
		X"00",X"00",X"07",X"0F",X"07",X"0F",X"2F",X"07",X"C0",X"D0",X"C8",X"E0",X"C8",X"C8",X"C0",X"E4",
		X"07",X"07",X"0E",X"0F",X"0F",X"01",X"00",X"00",X"C0",X"E0",X"F1",X"F9",X"FC",X"D2",X"01",X"19",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"F8",X"F2",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"F3",X"E0",X"C0",X"C0",X"80",X"80",X"0F",
		X"FF",X"FC",X"FC",X"FC",X"FD",X"FE",X"FE",X"FE",X"70",X"00",X"00",X"02",X"1C",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"0E",X"07",X"03",X"00",X"01",X"03",X"06",
		X"00",X"00",X"08",X"00",X"00",X"10",X"10",X"10",X"0D",X"8E",X"C6",X"37",X"0E",X"0F",X"0C",X"1E",
		X"00",X"20",X"98",X"E8",X"F1",X"19",X"CD",X"C9",X"00",X"00",X"00",X"00",X"00",X"30",X"31",X"21",
		X"91",X"31",X"39",X"38",X"9D",X"0D",X"14",X"04",X"41",X"79",X"71",X"F1",X"E0",X"E0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"0A",X"02",X"27",X"68",X"71",X"E4",
		X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"7F",X"FC",X"FA",X"10",X"22",X"10",X"10",X"60",X"F8",
		X"FC",X"FE",X"D1",X"B0",X"A0",X"E0",X"E0",X"D8",X"00",X"00",X"80",X"00",X"00",X"20",X"20",X"70",
		X"F8",X"DC",X"BC",X"AE",X"EE",X"A2",X"E0",X"A0",X"30",X"38",X"1C",X"18",X"00",X"00",X"00",X"00",
		X"BD",X"F7",X"FD",X"B3",X"FE",X"FE",X"40",X"00",X"DF",X"FA",X"FF",X"FD",X"EF",X"36",X"00",X"00",
		X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"40",X"44",X"65",X"63",X"A3",X"B7",X"BF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BE",X"BC",X"B8",X"F0",X"E0",X"E0",X"F0",X"F0",
		X"10",X"50",X"F8",X"FE",X"FE",X"CF",X"8F",X"07",X"0E",X"0C",X"0C",X"1C",X"38",X"38",X"78",X"79",
		X"01",X"03",X"07",X"03",X"00",X"04",X"06",X"06",X"D0",X"F0",X"E0",X"F0",X"F0",X"0F",X"03",X"01",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"80",X"83",X"87",
		X"81",X"87",X"1F",X"FE",X"C0",X"80",X"C0",X"00",X"FB",X"F1",X"80",X"00",X"00",X"00",X"01",X"01",
		X"00",X"00",X"00",X"00",X"04",X"0E",X"87",X"CF",X"01",X"0F",X"7F",X"1F",X"0B",X"02",X"30",X"A6",
		X"CF",X"8F",X"0F",X"13",X"1F",X"17",X"17",X"17",X"18",X"BB",X"F4",X"7C",X"96",X"FA",X"FE",X"FF",
		X"FE",X"EE",X"DC",X"FC",X"F0",X"49",X"02",X"CD",X"6C",X"26",X"FB",X"59",X"D8",X"D4",X"96",X"90",
		X"FF",X"3E",X"1E",X"1E",X"AE",X"AC",X"37",X"BF",X"90",X"12",X"04",X"1B",X"4D",X"41",X"00",X"00",
		X"A9",X"A9",X"A5",X"BC",X"9A",X"AB",X"BF",X"AF",X"20",X"20",X"90",X"08",X"C0",X"C0",X"E6",X"4C",
		X"BC",X"84",X"9C",X"D6",X"DE",X"DE",X"F6",X"F6",X"06",X"04",X"60",X"18",X"18",X"08",X"08",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"0F",X"0E",X"0F",X"3F",X"3D",X"3E",X"00",X"00",X"00",X"20",X"38",X"3C",X"7C",X"78",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"06",X"03",X"81",X"E0",X"F8",X"FE",X"FF",X"FF",X"61",X"04",X"FC",X"00",X"00",X"00",X"00",X"E0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"F8",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"00",X"00",X"00",X"E0",X"FC",X"FF",X"FF",X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"E1",X"FD",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"0F",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"07",X"07",X"03",X"02",X"05",X"02",X"2D",X"95",X"FF",X"EB",X"95",X"B5",X"EA",X"A5",X"52",X"25",
		X"DF",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C6",X"E4",X"C0",X"AA",X"E2",X"C4",X"A0",X"E2",
		X"FF",X"FF",X"BB",X"5C",X"D6",X"AB",X"92",X"6D",X"C1",X"C7",X"E7",X"4B",X"A1",X"CB",X"E2",X"7A",
		X"57",X"79",X"E9",X"68",X"6D",X"6A",X"6F",X"5F",X"B8",X"A8",X"D0",X"6C",X"DE",X"2C",X"1F",X"5F",
		X"6F",X"6D",X"4A",X"77",X"DE",X"C4",X"E1",X"F1",X"9E",X"3E",X"4F",X"AC",X"52",X"D7",X"71",X"3B",
		X"7E",X"6E",X"77",X"73",X"53",X"73",X"5B",X"71",X"0C",X"08",X"04",X"00",X"0C",X"02",X"02",X"84",
		X"68",X"18",X"0D",X"2D",X"01",X"7E",X"7E",X"7E",X"94",X"8C",X"8C",X"8B",X"9F",X"63",X"77",X"73",
		X"3F",X"7E",X"6E",X"7C",X"7C",X"FE",X"FE",X"FC",X"38",X"3C",X"32",X"78",X"70",X"68",X"42",X"E8",
		X"F8",X"FC",X"FD",X"FF",X"FF",X"FD",X"FE",X"FF",X"94",X"A4",X"48",X"B0",X"CA",X"F0",X"A8",X"52",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FD",X"FD",X"EB",X"FC",X"B5",
		X"FF",X"FE",X"FE",X"FC",X"F6",X"FF",X"FA",X"AF",X"DD",X"D7",X"DD",X"9B",X"DF",X"76",X"5D",X"35",
		X"7A",X"EF",X"BB",X"5A",X"F3",X"BB",X"6E",X"FF",X"F0",X"A0",X"F0",X"E0",X"B8",X"AC",X"9E",X"BE",
		X"DB",X"7B",X"7B",X"56",X"FB",X"5F",X"9D",X"DB",X"BD",X"EB",X"7B",X"FA",X"F7",X"BB",X"3B",X"96",
		X"F0",X"F8",X"F8",X"78",X"18",X"2C",X"20",X"FC",X"88",X"88",X"C0",X"40",X"C0",X"61",X"60",X"7C",
		X"F8",X"FD",X"7D",X"FF",X"5F",X"FF",X"BF",X"6F",X"FE",X"1C",X"88",X"88",X"C9",X"E1",X"E7",X"F7",
		X"7F",X"7F",X"7F",X"7F",X"78",X"91",X"40",X"53",X"CB",X"D3",X"EB",X"E3",X"09",X"7F",X"BF",X"FF",
		X"81",X"81",X"01",X"01",X"81",X"80",X"D0",X"C0",X"FF",X"F3",X"E1",X"F1",X"F8",X"7E",X"3F",X"1F",
		X"7E",X"FF",X"5F",X"7B",X"BE",X"5F",X"3F",X"FF",X"D0",X"A8",X"D4",X"68",X"D2",X"B0",X"24",X"D0",
		X"6F",X"BE",X"DF",X"7D",X"FF",X"FB",X"FF",X"7D",X"A8",X"D0",X"72",X"A8",X"52",X"F0",X"68",X"A4",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FE",X"FB",X"F9",X"EB",X"EA",
		X"FF",X"FF",X"FE",X"FA",X"FA",X"EA",X"E8",X"A9",X"A9",X"A1",X"E9",X"A9",X"8B",X"89",X"A2",X"AA",
		X"AD",X"7A",X"AD",X"DD",X"B4",X"3B",X"BF",X"AB",X"AF",X"ED",X"EA",X"7F",X"EA",X"67",X"DA",X"6D",
		X"DB",X"BE",X"BB",X"7D",X"AB",X"BB",X"BB",X"75",X"7F",X"F3",X"BA",X"6B",X"6F",X"6E",X"BB",X"7E",
		X"60",X"F8",X"9C",X"F8",X"EE",X"5F",X"D9",X"B9",X"79",X"39",X"3A",X"14",X"30",X"54",X"54",X"9E",
		X"B9",X"6F",X"DD",X"75",X"DC",X"DE",X"D2",X"BC",X"B9",X"98",X"B8",X"9A",X"93",X"B3",X"30",X"30",
		X"CD",X"99",X"48",X"43",X"A7",X"A0",X"B2",X"32",X"4F",X"1F",X"9C",X"1E",X"1C",X"98",X"A4",X"9C",
		X"93",X"03",X"58",X"4C",X"AC",X"AC",X"24",X"54",X"06",X"66",X"E1",X"C6",X"43",X"43",X"43",X"66",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"F2",X"E8",
		X"FF",X"FF",X"FE",X"F8",X"F0",X"E0",X"C0",X"F0",X"EE",X"92",X"0A",X"60",X"96",X"0A",X"0B",X"08",
		X"AE",X"A2",X"A2",X"8A",X"8A",X"A8",X"AA",X"6E",X"AA",X"CA",X"AA",X"A2",X"A8",X"AA",X"AB",X"A2",
		X"8A",X"BA",X"72",X"E2",X"AA",X"AE",X"A8",X"0A",X"AA",X"AE",X"4A",X"32",X"98",X"AA",X"AA",X"A2",
		X"F2",X"AE",X"FE",X"F6",X"7C",X"DE",X"D6",X"DF",X"C2",X"E1",X"E1",X"E9",X"49",X"45",X"54",X"75",
		X"BD",X"6D",X"F9",X"DB",X"FF",X"77",X"DF",X"5D",X"5A",X"B6",X"B7",X"F7",X"8B",X"5B",X"7A",X"FE",
		X"00",X"00",X"80",X"88",X"98",X"F8",X"F0",X"80",X"FA",X"FC",X"DE",X"FC",X"F8",X"E0",X"7C",X"7E",
		X"E1",X"69",X"7D",X"FD",X"D9",X"DF",X"DF",X"73",X"7E",X"7E",X"7E",X"3E",X"70",X"38",X"78",X"7C",
		X"FE",X"FF",X"FF",X"FB",X"FE",X"FF",X"FF",X"FF",X"D0",X"A8",X"D4",X"68",X"D2",X"B0",X"24",X"D0",
		X"FF",X"FE",X"FF",X"FD",X"FF",X"FB",X"FF",X"FD",X"A8",X"D0",X"72",X"A8",X"52",X"F0",X"68",X"A4",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"F8",X"F0",X"E0",X"C0",X"80",
		X"FF",X"FE",X"FC",X"F8",X"F0",X"E0",X"D2",X"83",X"12",X"15",X"12",X"45",X"67",X"33",X"3B",X"3B",
		X"02",X"03",X"03",X"02",X"02",X"00",X"10",X"68",X"19",X"0A",X"12",X"16",X"0B",X"1A",X"14",X"11",
		X"54",X"50",X"D8",X"F5",X"DB",X"9F",X"9B",X"13",X"3A",X"36",X"38",X"11",X"12",X"8A",X"CA",X"C6",
		X"F5",X"BE",X"AC",X"FD",X"DB",X"7D",X"FD",X"AD",X"D7",X"EB",X"EF",X"A7",X"FE",X"6B",X"DF",X"FD",
		X"BF",X"77",X"BD",X"9D",X"BF",X"F7",X"6F",X"BD",X"6F",X"CE",X"EF",X"6F",X"E9",X"FC",X"BD",X"ED",
		X"20",X"A8",X"AF",X"B0",X"03",X"09",X"05",X"10",X"7F",X"7E",X"7C",X"79",X"79",X"3B",X"B9",X"B9",
		X"0A",X"01",X"0A",X"05",X"02",X"01",X"0A",X"04",X"BB",X"79",X"FD",X"2B",X"B5",X"EF",X"57",X"BB",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"FA",X"F2",X"EA",X"C8",X"C0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"C1",X"C1",X"E3",X"F2",X"F8",X"FC",X"FE",
		X"01",X"03",X"85",X"BA",X"CE",X"9B",X"D3",X"0A",X"59",X"B0",X"12",X"A3",X"D1",X"B0",X"39",X"3A",
		X"40",X"B3",X"A5",X"D5",X"8A",X"E7",X"42",X"6C",X"AB",X"F1",X"B5",X"5C",X"5B",X"63",X"65",X"72",
		X"31",X"B9",X"21",X"3B",X"D5",X"4A",X"31",X"08",X"CA",X"4E",X"82",X"05",X"22",X"88",X"C6",X"A2",
		X"44",X"6C",X"11",X"45",X"13",X"55",X"16",X"93",X"52",X"61",X"21",X"40",X"49",X"80",X"82",X"C2",
		X"00",X"01",X"04",X"02",X"00",X"00",X"02",X"00",X"55",X"17",X"AB",X"5B",X"87",X"3D",X"D7",X"2B",
		X"01",X"04",X"00",X"02",X"00",X"00",X"04",X"01",X"4F",X"37",X"CD",X"9F",X"2B",X"97",X"2F",X"57",
		X"04",X"80",X"F0",X"F8",X"FC",X"FC",X"FF",X"FF",X"73",X"7B",X"D2",X"98",X"1B",X"13",X"03",X"82",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E0",X"E0",X"F8",X"FC",X"FC",X"FE",X"FF",X"FF",
		X"C3",X"9C",X"2C",X"60",X"00",X"88",X"88",X"08",X"A0",X"80",X"82",X"1E",X"19",X"0A",X"06",X"83",
		X"19",X"0B",X"1E",X"0B",X"1E",X"02",X"8A",X"E2",X"82",X"E0",X"A0",X"E8",X"88",X"1C",X"E8",X"AA",
		X"F2",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"2A",X"8B",X"E8",X"82",X"AA",X"FA",X"F9",X"FA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"E2",X"8A",X"08",X"A8",X"AA",X"AB",X"2A",X"9A",X"2C",X"EA",X"EC",X"A6",X"8E",X"AC",X"AC",
		X"BA",X"EA",X"EA",X"AA",X"AA",X"EB",X"F2",X"FE",X"B9",X"A2",X"A9",X"AA",X"44",X"A2",X"87",X"AD",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"47",X"AB",X"B6",X"A7",X"FA",X"F7",X"F9",X"FD",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"DB",X"7D",X"D5",X"FD",X"B6",X"65",X"DE",X"DD",X"DE",X"F7",X"77",X"E4",X"B7",X"B3",X"B6",X"D7",
		X"55",X"FD",X"DD",X"F7",X"FD",X"FB",X"FE",X"FF",X"BF",X"F7",X"4F",X"9D",X"D7",X"D7",X"77",X"D9",
		X"9A",X"BA",X"8F",X"97",X"25",X"AE",X"04",X"32",X"C5",X"D9",X"91",X"08",X"F1",X"A0",X"79",X"04",
		X"4D",X"BB",X"2A",X"84",X"39",X"D6",X"3D",X"95",X"1F",X"50",X"22",X"D7",X"63",X"E5",X"81",X"C1",
		X"3F",X"2E",X"3C",X"3F",X"0B",X"18",X"15",X"02",X"C4",X"E0",X"70",X"92",X"D1",X"63",X"AD",X"91",
		X"4C",X"5A",X"AF",X"A2",X"20",X"62",X"36",X"7D",X"1F",X"8F",X"FF",X"A7",X"5F",X"EB",X"7D",X"F3",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"E1",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FE",X"F0",X"00",X"0F",X"FF",X"FF",X"FF",X"FF",X"3F",X"3B",X"18",X"E1",X"F0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"E0",X"C0",X"C0",X"F7",X"01",X"FD",X"17",X"FF",X"7F",X"3F",X"38",X"FC",X"FD",X"FD",X"FC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FE",X"00",X"00",X"FF",X"FF",X"00",X"FF",X"87",X"C3",X"40",X"40",X"C0",X"C3",X"40",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F9",X"FF",X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",
		X"F0",X"E0",X"C3",X"07",X"0F",X"3F",X"FF",X"FF",X"0F",X"03",X"FC",X"FE",X"FE",X"FE",X"80",X"80",
		X"E0",X"80",X"3F",X"FF",X"00",X"C0",X"FC",X"F8",X"7F",X"00",X"1F",X"E0",X"20",X"07",X"04",X"07",
		X"F8",X"F8",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"07",X"07",X"07",X"07",X"07",X"07",X"8F",X"88",
		X"FF",X"00",X"FF",X"00",X"00",X"FF",X"00",X"00",X"FF",X"00",X"FF",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"F8",X"F0",X"F8",X"00",X"00",X"00",X"00",X"00",X"F8",X"F0",X"F8",X"00",X"00",X"00",
		X"FF",X"00",X"FF",X"00",X"00",X"FF",X"00",X"00",X"FF",X"00",X"FF",X"00",X"08",X"C4",X"04",X"0D",
		X"00",X"03",X"FF",X"F7",X"FB",X"01",X"00",X"00",X"7D",X"FD",X"E3",X"03",X"03",X"F0",X"FC",X"7C",
		X"1F",X"4F",X"FE",X"06",X"07",X"00",X"3F",X"C0",X"40",X"0F",X"7F",X"FF",X"FC",X"01",X"FF",X"00",
		X"C0",X"FF",X"FF",X"FF",X"C0",X"00",X"00",X"C0",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"03",X"27",X"EF",X"FE",X"0F",X"FF",X"9F",X"0F",X"56",X"C9",X"9A",X"E1",X"E8",X"92",X"68",X"C1",
		X"03",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"A8",X"CD",X"CE",X"EE",X"0C",X"0C",X"0C",X"0C",
		X"DF",X"00",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"9F",X"01",X"E0",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"07",X"C0",X"F8",X"FF",X"FF",X"FF",X"F0",X"F0",X"F1",X"61",X"1B",X"3B",X"CF",X"CF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"17",X"01",X"FD",X"F7",X"F0",X"FC",X"C0",X"C7",X"E0",X"E0",X"E0",X"E1",X"1D",X"1D",X"3B",X"CF",
		X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FE",X"43",X"41",X"7F",X"E7",X"FF",X"E7",X"F8",X"E2",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"82",X"FE",X"FD",X"FB",X"F7",X"EF",X"DC",X"BC",
		X"03",X"C0",X"F8",X"FF",X"FF",X"FF",X"0F",X"FF",X"80",X"00",X"00",X"FE",X"FD",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E0",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"87",X"03",X"81",
		X"00",X"00",X"FF",X"FF",X"FF",X"F8",X"F8",X"F8",X"F8",X"F8",X"00",X"00",X"00",X"FF",X"8F",X"8F",
		X"FC",X"86",X"87",X"FF",X"87",X"87",X"FF",X"FF",X"FC",X"F8",X"E0",X"E0",X"FF",X"FF",X"FF",X"FF",
		X"00",X"FF",X"F8",X"F0",X"F8",X"FF",X"FF",X"00",X"00",X"FF",X"F8",X"F0",X"F8",X"FF",X"FF",X"07",
		X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"07",X"06",X"04",X"04",X"04",X"05",X"05",X"05",
		X"00",X"FF",X"FF",X"F8",X"F0",X"F8",X"FF",X"FB",X"3F",X"FF",X"F0",X"F0",X"FC",X"FC",X"F0",X"F0",
		X"7B",X"7B",X"FB",X"FB",X"FB",X"FA",X"FA",X"FA",X"FC",X"F8",X"CF",X"CF",X"CF",X"7F",X"7F",X"7F",
		X"C0",X"03",X"46",X"03",X"40",X"03",X"46",X"03",X"01",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",
		X"40",X"00",X"C0",X"40",X"C0",X"40",X"C1",X"41",X"00",X"00",X"00",X"00",X"00",X"7C",X"FE",X"FC",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F1",X"F1",X"F3",X"F3",X"E3",X"E7",X"E7",X"E7",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C6",X"C6",X"CE",X"8E",X"8E",X"8E",X"8E",X"8E",
		X"9F",X"9F",X"9F",X"9D",X"1E",X"1F",X"1F",X"1F",X"8E",X"4B",X"1E",X"8F",X"0D",X"5E",X"9F",X"0E",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1E",X"1E",X"A7",X"F3",X"A1",X"E4",X"C8",X"EC",X"DC",X"7C",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"F8",X"F8",X"FF",X"FF",X"EF",X"9F",X"7F",X"3F",X"0F",X"03",
		X"F0",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"80",X"E0",X"F0",X"FC",X"FF",
		X"FF",X"FE",X"FD",X"FB",X"F3",X"F9",X"FC",X"FE",X"7F",X"F9",X"F9",X"FF",X"F3",X"F3",X"FF",X"79",
		X"FF",X"7F",X"3F",X"0F",X"03",X"01",X"00",X"00",X"39",X"9F",X"CC",X"E4",X"F3",X"F9",X"FC",X"7E",
		X"FF",X"F8",X"F8",X"FF",X"F0",X"F0",X"FF",X"F8",X"85",X"05",X"05",X"85",X"05",X"05",X"85",X"05",
		X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"05",X"85",X"83",X"87",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"87",X"87",X"FF",X"87",X"87",X"FF",X"FF",X"FF",X"C3",X"C3",X"FF",X"C3",X"C3",X"FF",
		X"FF",X"FF",X"FF",X"87",X"87",X"FF",X"87",X"87",X"FF",X"FF",X"FF",X"C3",X"C3",X"FF",X"C3",X"C3",
		X"FF",X"FF",X"E1",X"E1",X"FF",X"E1",X"E1",X"FF",X"E9",X"E9",X"E9",X"E9",X"EB",X"EB",X"EB",X"EB",
		X"FF",X"FF",X"FF",X"E1",X"E1",X"FF",X"E1",X"E1",X"EB",X"EB",X"EB",X"EB",X"E9",X"ED",X"ED",X"ED",
		X"F3",X"F3",X"E3",X"9F",X"9F",X"1F",X"FF",X"FF",X"FE",X"FC",X"F8",X"F0",X"E0",X"C0",X"80",X"00",
		X"FF",X"9F",X"9F",X"9F",X"F3",X"F3",X"F3",X"FE",X"80",X"C0",X"E0",X"F0",X"F8",X"FC",X"FE",X"7F",
		X"FF",X"FF",X"01",X"79",X"81",X"79",X"01",X"01",X"80",X"81",X"B3",X"A0",X"80",X"A0",X"A0",X"80",
		X"01",X"79",X"81",X"79",X"01",X"01",X"FF",X"FF",X"A0",X"A0",X"80",X"A0",X"B3",X"81",X"80",X"FC",
		X"00",X"FF",X"FE",X"00",X"00",X"00",X"00",X"00",X"8E",X"8E",X"8E",X"8E",X"8E",X"9E",X"9C",X"9C",
		X"00",X"00",X"00",X"00",X"FE",X"FF",X"00",X"00",X"9C",X"9C",X"9C",X"9C",X"9C",X"1C",X"1C",X"1C",
		X"1E",X"1E",X"1E",X"1E",X"1E",X"1E",X"1E",X"1E",X"7C",X"2A",X"04",X"09",X"14",X"1E",X"3C",X"39",
		X"1E",X"1E",X"1E",X"1E",X"1F",X"1F",X"1E",X"1E",X"36",X"7D",X"7C",X"F1",X"E4",X"EA",X"74",X"F9",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E0",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"F8",X"C7",X"FF",X"F8",X"FF",X"FF",X"F0",X"00",X"3E",X"FE",X"FE",X"00",X"80",X"FC",
		X"FF",X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FC",X"FF",X"FC",X"F3",X"3F",X"FC",X"FF",X"FF",
		X"F0",X"7B",X"00",X"7B",X"7B",X"00",X"00",X"7B",X"7E",X"FF",X"00",X"FF",X"FF",X"00",X"00",X"FF",
		X"F0",X"C7",X"3C",X"FF",X"FC",X"03",X"C3",X"FF",X"1F",X"E0",X"00",X"F7",X"00",X"F7",X"F7",X"FF",
		X"00",X"F1",X"06",X"8E",X"E6",X"03",X"00",X"FF",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"00",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"F8",X"01",X"E7",X"FF",X"E3",
		X"00",X"FF",X"00",X"00",X"00",X"F0",X"00",X"F0",X"00",X"00",X"1F",X"00",X"00",X"3F",X"7F",X"FF",
		X"F1",X"03",X"F3",X"07",X"77",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"3E",X"3C",
		X"00",X"00",X"FF",X"FF",X"E1",X"00",X"7F",X"7F",X"0F",X"00",X"FF",X"FF",X"C7",X"00",X"FF",X"FF",
		X"3F",X"BF",X"BF",X"BF",X"BF",X"00",X"00",X"F1",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"E3",
		X"FA",X"7A",X"7B",X"7B",X"7B",X"3B",X"BB",X"DB",X"7F",X"7F",X"CF",X"CF",X"CF",X"F8",X"F8",X"E0",
		X"DB",X"EB",X"EB",X"EB",X"EB",X"03",X"03",X"C3",X"E0",X"F8",X"F8",X"E0",X"E0",X"F8",X"C4",X"84",
		X"41",X"C0",X"40",X"C0",X"40",X"C0",X"00",X"43",X"8E",X"04",X"00",X"00",X"00",X"00",X"00",X"C0",
		X"06",X"43",X"00",X"43",X"06",X"43",X"00",X"7F",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"01",X"FF",
		X"00",X"00",X"F8",X"18",X"F8",X"00",X"FA",X"0D",X"1C",X"1C",X"1C",X"38",X"38",X"7A",X"FF",X"EF",
		X"0A",X"0F",X"FE",X"3F",X"1F",X"7D",X"FE",X"FF",X"1E",X"57",X"E9",X"E4",X"A1",X"F0",X"55",X"2A",
		X"1E",X"1E",X"18",X"3E",X"7F",X"BE",X"F6",X"EF",X"FA",X"78",X"75",X"3C",X"5A",X"91",X"2A",X"04",
		X"6F",X"F6",X"C7",X"AB",X"F2",X"6C",X"E8",X"C5",X"0A",X"9C",X"07",X"22",X"85",X"42",X"00",X"68",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"F8",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F0",X"F0",X"F0",X"70",X"70",X"F0",X"F8",X"FE",X"18",X"31",X"31",X"18",X"0C",X"06",X"3F",X"3F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"81",X"F3",X"F3",X"81",X"F1",X"00",X"00",X"FF",X"02",X"E7",X"E7",X"02",X"E3",X"00",X"00",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"07",X"C6",X"C5",X"07",X"C7",X"04",X"07",X"FF",X"0D",X"7F",X"FF",X"E3",X"01",X"00",X"E0",X"FE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"E0",X"E0",X"FF",X"FF",X"3F",X"00",X"02",X"02",X"00",X"09",X"FB",X"F7",X"D3",X"06",X"07",X"AB",
		X"CB",X"FF",X"FF",X"FF",X"FF",X"DF",X"AF",X"3D",X"C5",X"E1",X"C2",X"61",X"A9",X"C4",X"D0",X"B2",
		X"C5",X"F0",X"F8",X"D0",X"58",X"E9",X"F0",X"E3",X"FC",X"BA",X"1D",X"2C",X"2A",X"44",X"C6",X"E0",
		X"F1",X"B9",X"A8",X"D0",X"89",X"EC",X"BD",X"EF",X"92",X"E0",X"50",X"80",X"24",X"00",X"60",X"28",
		X"FD",X"F7",X"FF",X"FE",X"FB",X"FF",X"FE",X"FF",X"91",X"60",X"B4",X"C0",X"11",X"C8",X"F4",X"A2",
		X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"58",X"C4",X"B9",X"D0",X"EC",X"C9",X"BA",X"ED",
		X"FF",X"FC",X"FE",X"FE",X"FF",X"FE",X"FF",X"FF",X"EA",X"FC",X"E9",X"7A",X"1C",X"DA",X"1D",X"4C",
		X"FF",X"FE",X"FF",X"FD",X"FF",X"FB",X"FE",X"FD",X"89",X"86",X"EA",X"90",X"55",X"E2",X"B0",X"C9",
		X"FD",X"FE",X"FD",X"FA",X"FC",X"FE",X"FC",X"FB",X"6A",X"88",X"24",X"91",X"04",X"8A",X"C8",X"85",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"D0",X"45",X"D8",X"B5",X"EA",X"FE",X"FF",X"FF",
		X"B0",X"04",X"A0",X"68",X"80",X"20",X"A1",X"94",X"07",X"47",X"66",X"2F",X"65",X"EE",X"C7",X"B6",
		X"41",X"03",X"95",X"97",X"4F",X"9F",X"15",X"BE",X"C7",X"CB",X"C1",X"AD",X"D2",X"68",X"91",X"C8",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F5",X"FE",X"FB",X"FE",X"FF",X"FD",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C8",X"E2",X"94",X"F1",X"68",X"AA",X"D0",X"E5",X"8D",X"07",X"8F",X"5A",X"1C",X"39",X"0A",X"3E",
		X"40",X"D8",X"88",X"5D",X"BF",X"BF",X"FF",X"FF",X"74",X"BD",X"FE",X"FD",X"FE",X"FB",X"FF",X"FF",
		X"1F",X"1F",X"8B",X"57",X"03",X"03",X"85",X"16",X"54",X"88",X"C1",X"90",X"60",X"80",X"12",X"A0",
		X"8E",X"1E",X"BF",X"36",X"7F",X"5F",X"3E",X"2B",X"08",X"80",X"54",X"82",X"C8",X"94",X"E4",X"B0",
		X"C7",X"6F",X"CF",X"87",X"43",X"83",X"88",X"23",X"7A",X"DC",X"F5",X"EA",X"FD",X"78",X"D0",X"01",
		X"87",X"06",X"17",X"B7",X"3F",X"F7",X"F6",X"3F",X"54",X"A0",X"D4",X"A1",X"43",X"97",X"87",X"57",
		X"07",X"0B",X"17",X"8E",X"1F",X"0F",X"1F",X"2E",X"AA",X"40",X"94",X"A0",X"48",X"B0",X"04",X"A1",
		X"9F",X"1F",X"8E",X"1F",X"0F",X"07",X"0B",X"07",X"50",X"84",X"D0",X"84",X"40",X"A9",X"C0",X"70",
		X"4F",X"0F",X"8F",X"07",X"07",X"03",X"83",X"02",X"A8",X"58",X"D2",X"E0",X"B4",X"E0",X"48",X"B0",
		X"00",X"81",X"43",X"01",X"03",X"87",X"03",X"07",X"F9",X"C0",X"AA",X"A8",X"D2",X"48",X"E4",X"98",
		X"88",X"28",X"41",X"EA",X"30",X"7C",X"39",X"7C",X"0A",X"1D",X"0E",X"1E",X"3A",X"1C",X"3D",X"52",
		X"28",X"BC",X"1A",X"3C",X"9E",X"6E",X"14",X"88",X"1C",X"9F",X"3C",X"1E",X"3D",X"1E",X"8F",X"0E",
		X"87",X"8B",X"47",X"AF",X"27",X"4F",X"E3",X"45",X"A8",X"62",X"E4",X"56",X"CC",X"98",X"F4",X"F8",
		X"73",X"E9",X"74",X"30",X"70",X"1A",X"90",X"42",X"DA",X"ED",X"FA",X"D4",X"52",X"28",X"80",X"20",
		X"43",X"61",X"23",X"71",X"28",X"70",X"E4",X"38",X"F7",X"E2",X"F9",X"F0",X"F9",X"EB",X"B7",X"55",
		X"70",X"65",X"B4",X"7B",X"51",X"28",X"38",X"11",X"2E",X"1D",X"1D",X"4C",X"08",X"A0",X"00",X"00",
		X"DA",X"E3",X"C2",X"ED",X"D2",X"CB",X"90",X"FD",X"00",X"24",X"08",X"05",X"04",X"02",X"00",X"40",
		X"B8",X"FC",X"F3",X"7B",X"E7",X"7B",X"2F",X"0F",X"C0",X"A0",X"02",X"40",X"A0",X"50",X"94",X"EA",
		X"00",X"24",X"88",X"0D",X"1A",X"8C",X"5E",X"1D",X"8D",X"47",X"16",X"0D",X"06",X"0F",X"16",X"0C",
		X"0E",X"9D",X"0D",X"1E",X"88",X"2C",X"04",X"80",X"5E",X"36",X"3D",X"66",X"73",X"C1",X"A0",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
