library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity time_pilot_char_grphx is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of time_pilot_char_grphx is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"88",X"99",X"99",X"99",X"99",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"00",
		X"70",X"30",X"10",X"32",X"32",X"32",X"30",X"1E",X"00",X"80",X"C4",X"C4",X"C4",X"C4",X"80",X"0E",
		X"CC",X"EE",X"BB",X"99",X"88",X"CC",X"CC",X"00",X"00",X"00",X"00",X"EE",X"EE",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"4C",X"4C",X"0C",X"04",
		X"00",X"00",X"00",X"00",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"62",X"40",X"C0",X"00",
		X"00",X"00",X"67",X"23",X"03",X"03",X"01",X"77",X"00",X"00",X"68",X"68",X"68",X"2C",X"C0",X"F7",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"11",X"00",X"00",X"07",X"1F",
		X"00",X"00",X"01",X"CF",X"16",X"96",X"3C",X"8F",X"00",X"00",X"80",X"C4",X"00",X"00",X"80",X"08",
		X"0F",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"F1",X"70",X"00",X"00",X"11",X"00",X"00",
		X"CF",X"F8",X"E1",X"87",X"43",X"ED",X"10",X"00",X"0C",X"80",X"80",X"00",X"00",X"C4",X"80",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"00",X"CC",X"EE",X"22",X"22",X"22",X"EE",X"CC",X"00",
		X"FF",X"FF",X"11",X"00",X"11",X"FF",X"FF",X"00",X"00",X"88",X"CC",X"EE",X"CC",X"88",X"00",X"00",
		X"FF",X"FF",X"11",X"33",X"11",X"FF",X"FF",X"00",X"EE",X"EE",X"CC",X"88",X"CC",X"EE",X"EE",X"00",
		X"00",X"11",X"11",X"11",X"11",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"77",X"CC",X"88",X"88",X"77",X"33",X"00",X"88",X"CC",X"22",X"22",X"66",X"CC",X"88",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"99",X"99",X"99",X"99",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"00",
		X"00",X"66",X"99",X"99",X"BB",X"FF",X"66",X"00",X"CC",X"EE",X"AA",X"AA",X"22",X"22",X"CC",X"00",
		X"00",X"00",X"00",X"0F",X"FC",X"4B",X"FB",X"3C",X"00",X"00",X"00",X"0C",X"E6",X"4B",X"FB",X"87",
		X"00",X"00",X"00",X"00",X"00",X"10",X"A9",X"5A",X"00",X"00",X"00",X"00",X"00",X"80",X"48",X"A4",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"00",X"00",X"00",
		X"33",X"23",X"01",X"91",X"91",X"81",X"81",X"93",X"00",X"88",X"88",X"08",X"08",X"0C",X"5D",X"5D",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"EE",X"77",X"33",X"77",X"EE",X"CC",X"00",X"66",X"EE",X"CC",X"88",X"CC",X"EE",X"66",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"EE",X"22",X"22",X"22",X"66",X"44",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"11",X"33",X"33",X"33",X"33",X"33",X"00",X"FF",X"FF",X"F8",X"F7",X"F7",X"F8",X"FF",
		X"00",X"88",X"CC",X"E2",X"FD",X"FD",X"F3",X"FF",X"00",X"00",X"00",X"00",X"00",X"88",X"CC",X"CC",
		X"33",X"33",X"33",X"33",X"33",X"11",X"00",X"00",X"F9",X"F6",X"F6",X"F6",X"F6",X"FF",X"FF",X"00",
		X"F3",X"FD",X"FD",X"FD",X"EC",X"CC",X"88",X"00",X"CC",X"CC",X"88",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"FF",X"CC",X"66",X"33",X"11",X"00",X"88",X"EE",X"EE",X"88",X"88",X"88",X"88",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"88",X"88",X"FF",X"FF",X"00",X"00",X"00",X"66",X"22",X"22",X"EE",X"EE",X"00",X"66",X"66",
		X"00",X"00",X"CC",X"CC",X"22",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"00",X"00",X"00",
		X"1E",X"0F",X"0F",X"07",X"16",X"3C",X"07",X"03",X"F7",X"F6",X"F4",X"E5",X"E5",X"E5",X"E5",X"F0",
		X"F3",X"F3",X"79",X"79",X"79",X"3C",X"3C",X"16",X"E9",X"E9",X"C3",X"C3",X"C2",X"86",X"86",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"FF",X"88",X"88",X"88",X"FF",X"77",X"00",X"AA",X"CC",X"EE",X"AA",X"22",X"EE",X"CC",X"00",
		X"33",X"44",X"88",X"AA",X"AA",X"99",X"44",X"33",X"CC",X"22",X"11",X"55",X"55",X"99",X"22",X"CC",
		X"00",X"00",X"00",X"00",X"03",X"03",X"01",X"77",X"00",X"00",X"00",X"00",X"68",X"2C",X"C0",X"F7",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"07",X"5A",X"5A",X"78",X"07",X"00",
		X"00",X"11",X"0F",X"C3",X"5B",X"4B",X"0F",X"11",X"00",X"EE",X"0C",X"0C",X"EE",X"0C",X"0C",X"EE",
		X"88",X"99",X"99",X"99",X"FF",X"FF",X"00",X"00",X"22",X"22",X"22",X"22",X"EE",X"EE",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"01",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",
		X"67",X"67",X"67",X"23",X"03",X"03",X"01",X"77",X"68",X"68",X"68",X"68",X"68",X"2C",X"C0",X"F7",
		X"FF",X"FF",X"77",X"33",X"77",X"FF",X"FF",X"00",X"EE",X"EE",X"00",X"88",X"00",X"EE",X"EE",X"00",
		X"99",X"99",X"99",X"88",X"CC",X"77",X"33",X"00",X"EE",X"EE",X"22",X"22",X"66",X"CC",X"88",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"11",X"33",X"77",X"FF",X"FF",X"00",X"EE",X"EE",X"CC",X"88",X"00",X"EE",X"EE",X"00",
		X"33",X"44",X"88",X"AA",X"AA",X"99",X"44",X"33",X"CC",X"22",X"11",X"55",X"55",X"99",X"22",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"33",X"44",X"88",X"00",X"00",X"00",X"00",X"00",X"88",X"44",X"22",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"EE",
		X"00",X"99",X"99",X"99",X"DD",X"77",X"33",X"00",X"CC",X"EE",X"22",X"22",X"22",X"EE",X"CC",X"00",
		X"11",X"11",X"11",X"FF",X"11",X"11",X"11",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"00",X"CC",X"EE",X"22",X"22",X"22",X"EE",X"CC",X"00",
		X"0F",X"84",X"08",X"08",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"08",X"08",X"08",X"08",X"08",X"08",X"0C",X"86",
		X"00",X"00",X"01",X"91",X"91",X"81",X"81",X"93",X"00",X"00",X"88",X"08",X"08",X"0C",X"5D",X"5D",
		X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"84",X"0C",X"08",X"08",X"08",X"08",X"08",X"08",
		X"00",X"00",X"FF",X"FF",X"44",X"00",X"00",X"00",X"22",X"22",X"EE",X"EE",X"22",X"22",X"00",X"00",
		X"00",X"00",X"44",X"AA",X"99",X"AA",X"44",X"00",X"22",X"44",X"44",X"AA",X"22",X"AA",X"44",X"00",
		X"00",X"00",X"74",X"30",X"10",X"10",X"00",X"00",X"00",X"00",X"F3",X"62",X"62",X"40",X"C0",X"00",
		X"00",X"89",X"8B",X"9B",X"EF",X"8B",X"03",X"FE",X"5A",X"5A",X"7E",X"DA",X"5A",X"78",X"C0",X"EE",
		X"16",X"16",X"16",X"12",X"03",X"03",X"03",X"01",X"0C",X"0C",X"0C",X"08",X"08",X"08",X"08",X"00",
		X"00",X"33",X"44",X"55",X"55",X"44",X"33",X"00",X"00",X"CC",X"22",X"AA",X"AA",X"22",X"CC",X"00",
		X"00",X"00",X"16",X"16",X"03",X"01",X"01",X"01",X"00",X"88",X"88",X"C8",X"C0",X"2C",X"2C",X"3C",
		X"FF",X"FF",X"11",X"11",X"11",X"FF",X"FF",X"00",X"EE",X"EE",X"00",X"00",X"00",X"EE",X"EE",X"00",
		X"08",X"08",X"0C",X"86",X"E1",X"0F",X"0C",X"08",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"FF",X"88",X"88",X"88",X"FF",X"77",X"00",X"CC",X"EE",X"22",X"22",X"22",X"EE",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"22",X"22",X"22",X"22",X"EE",X"EE",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"EE",X"FF",X"BB",X"99",X"88",X"88",X"00",X"22",X"22",X"22",X"AA",X"EE",X"EE",X"66",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"61",X"00",X"00",X"00",X"00",X"00",X"00",X"2C",X"2C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"99",X"99",X"99",X"FF",X"FF",X"00",X"00",X"22",X"22",X"22",X"22",X"EE",X"EE",X"00",X"00",
		X"77",X"FF",X"99",X"99",X"99",X"FF",X"66",X"00",X"88",X"CC",X"66",X"22",X"22",X"22",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"FF",X"99",X"88",X"88",X"FF",X"FF",X"00",X"22",X"66",X"EE",X"CC",X"88",X"EE",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"16",X"3C",X"3C",X"79",X"79",X"79",X"F3",X"F3",X"0C",X"86",X"86",X"C2",X"C3",X"C3",X"E9",X"E9",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3C",X"3C",X"16",X"03",X"03",X"03",X"07",X"0F",X"CB",X"CA",X"C2",X"C2",X"C3",X"E1",X"87",X"87",
		X"88",X"DD",X"FF",X"BB",X"99",X"88",X"00",X"00",X"CC",X"EE",X"22",X"22",X"22",X"66",X"44",X"00",
		X"00",X"99",X"99",X"99",X"DD",X"77",X"33",X"00",X"CC",X"EE",X"22",X"22",X"22",X"EE",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"88",X"FF",X"FF",X"88",X"88",X"00",X"00",X"22",X"22",X"EE",X"EE",X"22",X"22",X"00",X"00",
		X"77",X"FF",X"88",X"88",X"88",X"FF",X"77",X"00",X"CC",X"EE",X"22",X"22",X"22",X"EE",X"CC",X"00",
		X"3C",X"79",X"3C",X"1E",X"16",X"70",X"35",X"1E",X"F8",X"FC",X"ED",X"EF",X"E5",X"E9",X"F8",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"88",X"FF",X"FF",X"88",X"88",X"00",X"00",X"00",X"00",X"EE",X"EE",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"01",X"01",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"EF",X"8B",X"03",X"FE",X"00",X"00",X"00",X"00",X"5A",X"78",X"C0",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"77",X"CC",X"88",X"CC",X"77",X"33",X"00",X"EE",X"EE",X"88",X"88",X"88",X"EE",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"16",X"03",X"03",X"61",X"00",X"00",X"00",X"00",X"48",X"48",X"2C",X"2C",
		X"00",X"00",X"EE",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"CC",X"88",X"88",X"CC",X"77",X"33",X"00",X"44",X"66",X"22",X"22",X"66",X"CC",X"88",X"00",
		X"00",X"FF",X"BF",X"17",X"13",X"03",X"21",X"30",X"00",X"00",X"BE",X"1F",X"1F",X"1F",X"3E",X"BE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"CC",X"66",X"33",X"11",X"FF",X"FF",X"00",X"22",X"66",X"EE",X"CC",X"88",X"EE",X"EE",X"00",
		X"30",X"10",X"01",X"01",X"00",X"00",X"00",X"00",X"BE",X"8C",X"4C",X"4C",X"4C",X"4C",X"0C",X"04",
		X"88",X"CC",X"66",X"33",X"11",X"FF",X"FF",X"00",X"22",X"66",X"EE",X"CC",X"88",X"EE",X"EE",X"00",
		X"99",X"99",X"99",X"88",X"CC",X"77",X"33",X"00",X"EE",X"EE",X"22",X"22",X"66",X"CC",X"88",X"00",
		X"00",X"33",X"77",X"CC",X"88",X"CC",X"77",X"33",X"00",X"EE",X"EE",X"88",X"88",X"88",X"EE",X"EE",
		X"11",X"BB",X"AA",X"AA",X"AA",X"EE",X"EE",X"00",X"CC",X"EE",X"22",X"22",X"22",X"66",X"44",X"00",
		X"77",X"FF",X"88",X"88",X"88",X"FF",X"FF",X"00",X"00",X"88",X"88",X"88",X"88",X"EE",X"EE",X"00",
		X"0C",X"08",X"08",X"08",X"0C",X"0C",X"0C",X"C3",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0E",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"FF",
		X"00",X"00",X"1E",X"1E",X"16",X"03",X"03",X"61",X"00",X"00",X"80",X"48",X"48",X"48",X"2C",X"2C",
		X"77",X"FF",X"99",X"99",X"99",X"FF",X"66",X"00",X"88",X"CC",X"66",X"22",X"22",X"22",X"00",X"00",
		X"33",X"77",X"CC",X"88",X"88",X"FF",X"FF",X"00",X"88",X"CC",X"66",X"22",X"22",X"EE",X"EE",X"00",
		X"77",X"FF",X"88",X"88",X"88",X"FF",X"FF",X"00",X"00",X"88",X"88",X"88",X"88",X"EE",X"EE",X"00",
		X"EE",X"FF",X"11",X"11",X"FF",X"EE",X"00",X"00",X"00",X"00",X"EE",X"EE",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"01",X"00",X"00",X"00",X"01",X"07",X"1E",X"0F",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"00",
		X"66",X"FF",X"99",X"99",X"99",X"FF",X"FF",X"00",X"CC",X"EE",X"22",X"22",X"22",X"EE",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"2C",X"3C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DA",X"29",X"10",X"00",X"00",X"00",X"00",X"00",X"A4",X"48",X"80",X"00",X"00",X"00",X"00",X"00",
		X"01",X"03",X"0B",X"0F",X"2D",X"34",X"16",X"16",X"86",X"86",X"87",X"C3",X"C3",X"E1",X"8F",X"CB",
		X"FC",X"74",X"74",X"30",X"10",X"10",X"00",X"00",X"73",X"73",X"F3",X"62",X"62",X"40",X"C0",X"00",
		X"88",X"44",X"22",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"44",X"22",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"44",X"00",X"00",X"00",X"22",X"22",X"EE",X"EE",X"22",X"22",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"01",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"88",X"44",X"33",X"00",X"00",X"00",X"00",X"00",X"22",X"44",X"88",X"00",X"00",X"00",
		X"66",X"FF",X"BB",X"99",X"99",X"CC",X"44",X"00",X"22",X"22",X"AA",X"AA",X"EE",X"EE",X"66",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"CC",X"22",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"EE",X"22",X"22",X"22",X"66",X"44",X"00",
		X"00",X"55",X"DD",X"99",X"99",X"FF",X"66",X"00",X"CC",X"EE",X"22",X"22",X"22",X"66",X"44",X"00",
		X"00",X"00",X"00",X"00",X"91",X"81",X"81",X"93",X"00",X"00",X"00",X"00",X"08",X"0C",X"5D",X"5D",
		X"01",X"01",X"03",X"07",X"1E",X"16",X"16",X"3C",X"87",X"87",X"87",X"C3",X"C3",X"CB",X"E9",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"77",X"CC",X"88",X"CC",X"77",X"33",X"00",X"EE",X"EE",X"88",X"88",X"88",X"EE",X"EE",X"00",
		X"00",X"00",X"8B",X"9B",X"EF",X"8B",X"03",X"FE",X"00",X"00",X"7E",X"DA",X"5A",X"78",X"C0",X"EE",
		X"00",X"61",X"1E",X"1E",X"12",X"03",X"03",X"61",X"00",X"00",X"80",X"48",X"48",X"48",X"2C",X"2C",
		X"66",X"FF",X"BB",X"99",X"99",X"CC",X"44",X"00",X"22",X"22",X"AA",X"AA",X"EE",X"EE",X"66",X"00",
		X"CC",X"EE",X"FF",X"BB",X"99",X"88",X"88",X"00",X"22",X"22",X"22",X"AA",X"EE",X"EE",X"66",X"00",
		X"08",X"00",X"00",X"08",X"0E",X"C3",X"E1",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"F7",
		X"00",X"01",X"01",X"12",X"34",X"34",X"7C",X"FC",X"0C",X"04",X"86",X"42",X"63",X"63",X"F3",X"73",
		X"77",X"FF",X"88",X"88",X"88",X"FF",X"77",X"00",X"AA",X"CC",X"EE",X"AA",X"22",X"EE",X"CC",X"00",
		X"11",X"BB",X"AA",X"AA",X"AA",X"EE",X"EE",X"00",X"CC",X"EE",X"22",X"22",X"22",X"66",X"44",X"00",
		X"00",X"55",X"55",X"FF",X"55",X"55",X"22",X"00",X"88",X"44",X"44",X"EE",X"44",X"44",X"00",X"00",
		X"CC",X"EE",X"BB",X"99",X"88",X"CC",X"CC",X"00",X"00",X"00",X"00",X"EE",X"EE",X"00",X"00",X"00",
		X"66",X"FF",X"99",X"99",X"99",X"FF",X"FF",X"00",X"CC",X"EE",X"22",X"22",X"22",X"EE",X"EE",X"00",
		X"01",X"03",X"03",X"03",X"12",X"16",X"16",X"16",X"00",X"08",X"08",X"08",X"08",X"0C",X"0C",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"81",X"93",X"00",X"00",X"00",X"00",X"00",X"00",X"5D",X"5D",
		X"3C",X"1E",X"1E",X"1E",X"3C",X"3C",X"F3",X"F1",X"E9",X"CB",X"CB",X"CB",X"E9",X"FE",X"F8",X"CB",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"11",X"00",X"11",X"FF",X"FF",X"00",X"00",X"88",X"CC",X"EE",X"CC",X"88",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"BF",X"17",X"13",X"03",X"21",X"30",X"00",X"00",X"BE",X"1F",X"1F",X"1F",X"3E",X"BE",
		X"08",X"00",X"00",X"00",X"08",X"0F",X"0E",X"84",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"EE",X"77",X"33",X"77",X"EE",X"CC",X"00",X"66",X"EE",X"CC",X"88",X"CC",X"EE",X"66",X"00",
		X"FF",X"FF",X"11",X"33",X"77",X"FF",X"FF",X"00",X"EE",X"EE",X"CC",X"88",X"00",X"EE",X"EE",X"00",
		X"EE",X"FF",X"11",X"11",X"FF",X"EE",X"00",X"00",X"00",X"00",X"EE",X"EE",X"00",X"00",X"00",X"00",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"88",
		X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"4C",X"4C",X"4C",X"4C",X"0C",X"04",
		X"03",X"03",X"03",X"16",X"16",X"1E",X"3C",X"3C",X"08",X"08",X"08",X"0C",X"0C",X"0E",X"86",X"86",
		X"FF",X"FF",X"11",X"11",X"11",X"FF",X"FF",X"00",X"EE",X"EE",X"00",X"00",X"00",X"EE",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"22",X"22",X"22",X"22",X"EE",X"EE",X"00",X"00",
		X"86",X"0C",X"08",X"08",X"08",X"0C",X"0C",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"44",X"22",X"11",X"77",X"11",X"22",X"44",X"00",X"44",X"88",X"00",X"CC",X"00",X"88",X"44",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"01",X"01",X"03",X"07",X"09",X"00",X"00",X"78",X"78",X"E1",X"C3",X"87",X"87",X"0C",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"CC",X"88",X"88",X"CC",X"77",X"33",X"00",X"44",X"66",X"22",X"22",X"66",X"CC",X"88",X"00",
		X"88",X"DD",X"FF",X"BB",X"99",X"88",X"00",X"00",X"CC",X"EE",X"22",X"22",X"22",X"66",X"44",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"54",X"54",
		X"00",X"00",X"70",X"10",X"70",X"F0",X"F0",X"F0",X"00",X"00",X"80",X"80",X"C4",X"A2",X"A2",X"E6",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"76",X"45",X"45",X"44",X"00",X"00",X"00",X"00",
		X"F0",X"3C",X"1E",X"1E",X"16",X"10",X"00",X"00",X"A2",X"A2",X"E6",X"A2",X"A2",X"C4",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"34",X"34",X"7C",X"FC",X"00",X"00",X"00",X"00",X"63",X"63",X"F3",X"73",
		X"00",X"00",X"01",X"12",X"34",X"34",X"7C",X"FC",X"00",X"00",X"86",X"42",X"63",X"63",X"F3",X"73",
		X"00",X"66",X"99",X"99",X"BB",X"FF",X"66",X"00",X"CC",X"EE",X"AA",X"AA",X"22",X"22",X"CC",X"00",
		X"00",X"11",X"11",X"11",X"11",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"FF",X"99",X"88",X"88",X"FF",X"FF",X"00",X"22",X"66",X"EE",X"CC",X"88",X"EE",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"93",X"57",X"93",X"A1",X"B0",X"90",X"90",X"80",X"FF",X"9D",X"1D",X"3F",X"1D",X"5D",X"CC",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"88",X"FF",X"FF",X"88",X"88",X"00",X"00",X"00",X"00",X"EE",X"EE",X"00",X"00",X"00",X"00",
		X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"21",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"BE",
		X"FD",X"5A",X"FA",X"5A",X"0F",X"00",X"00",X"00",X"F7",X"4B",X"FB",X"4A",X"0C",X"00",X"00",X"00",
		X"08",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"B0",X"90",X"90",X"80",X"00",X"00",X"00",X"00",X"1D",X"5D",X"CC",X"88",
		X"00",X"00",X"00",X"00",X"03",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"C0",X"2C",X"2C",X"3C",
		X"33",X"77",X"CC",X"88",X"88",X"77",X"33",X"00",X"88",X"CC",X"22",X"22",X"66",X"CC",X"88",X"00",
		X"88",X"44",X"22",X"11",X"44",X"AA",X"44",X"00",X"44",X"AA",X"44",X"00",X"88",X"44",X"22",X"00",
		X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"03",
		X"FF",X"FF",X"11",X"33",X"11",X"FF",X"FF",X"00",X"EE",X"EE",X"CC",X"88",X"CC",X"EE",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1E",X"3C",X"3C",X"3D",X"78",X"F2",X"F3",X"79",X"E9",X"E1",X"F4",X"FC",X"FE",X"FC",X"ED",X"E9",
		X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"00",X"00",X"08",X"08",X"0C",X"0C",X"86",X"87",
		X"33",X"77",X"CC",X"88",X"88",X"FF",X"FF",X"00",X"88",X"CC",X"66",X"22",X"22",X"EE",X"EE",X"00",
		X"00",X"55",X"DD",X"99",X"99",X"FF",X"66",X"00",X"CC",X"EE",X"22",X"22",X"22",X"66",X"44",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"7C",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"F3",X"73",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"FF",
		X"3C",X"3C",X"1E",X"16",X"16",X"03",X"03",X"03",X"86",X"86",X"0E",X"0C",X"0C",X"08",X"08",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"FF",X"CC",X"66",X"33",X"11",X"00",X"88",X"EE",X"EE",X"88",X"88",X"88",X"88",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"01",X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"3C",X"07",X"03",
		X"FF",X"FF",X"77",X"33",X"77",X"FF",X"FF",X"00",X"EE",X"EE",X"00",X"88",X"00",X"EE",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"77",X"00",X"00",X"00",X"66",X"66",X"00",X"88",X"CC",
		X"00",X"00",X"00",X"00",X"13",X"03",X"21",X"30",X"00",X"00",X"00",X"00",X"1F",X"1F",X"3E",X"BE",
		X"00",X"00",X"93",X"A1",X"B0",X"90",X"90",X"80",X"00",X"00",X"1D",X"3F",X"1D",X"5D",X"CC",X"88",
		X"00",X"00",X"16",X"16",X"03",X"01",X"01",X"01",X"00",X"00",X"88",X"C8",X"C0",X"2C",X"2C",X"3C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"88",X"FF",X"FF",X"88",X"88",X"00",X"00",X"22",X"22",X"EE",X"EE",X"22",X"22",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"88",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"11",X"11",X"11",X"11",X"11",X"33",X"33",X"33",X"88",X"88",X"88",X"88",X"88",X"CC",X"CC",X"CC",
		X"11",X"11",X"11",X"11",X"33",X"33",X"33",X"77",X"88",X"88",X"88",X"88",X"CC",X"CC",X"CC",X"EE",
		X"11",X"11",X"33",X"33",X"33",X"77",X"77",X"77",X"88",X"88",X"CC",X"CC",X"CC",X"EE",X"EE",X"EE",
		X"33",X"33",X"33",X"33",X"33",X"33",X"77",X"77",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"EE",X"EE",
		X"33",X"33",X"33",X"33",X"33",X"77",X"77",X"FF",X"CC",X"CC",X"CC",X"CC",X"CC",X"EE",X"EE",X"FF",
		X"33",X"33",X"33",X"33",X"77",X"77",X"FF",X"FF",X"CC",X"CC",X"CC",X"CC",X"EE",X"EE",X"FF",X"FF",
		X"77",X"77",X"77",X"FF",X"FF",X"FF",X"FF",X"FF",X"EE",X"EE",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"77",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"33",X"33",X"77",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"33",X"33",X"77",X"77",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"EF",X"FC",X"FC",X"FC",X"FC",X"FC",X"FF",X"FF",X"7F",X"33",X"33",X"33",X"33",X"33",X"FF",
		X"00",X"00",X"33",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"11",X"33",X"FF",X"FF",X"FF",X"CF",X"0F",X"FC",X"FC",X"FC",X"DA",X"AD",X"0E",X"0E",X"6C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"66",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"ED",X"FC",X"FC",X"FE",X"FF",X"77",X"77",X"0F",X"86",X"80",X"00",X"33",X"FF",X"FF",X"EF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"33",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"D1",X"FF",X"00",X"00",X"00",X"00",X"00",X"FC",X"FC",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"66",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"0F",X"00",X"00",X"00",X"00",X"80",X"FC",X"FC",X"FC",X"96",X"43",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"33",X"11",X"00",X"00",X"00",X"0C",X"FC",X"FC",X"FC",X"FC",X"EC",X"EC",X"44",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"FF",X"FF",X"FC",X"1E",X"0F",X"0F",X"0C",X"00",X"FC",X"FC",X"BC",X"1E",X"96",X"02",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",X"CF",X"3F",X"0F",X"FF",X"FF",X"FF",X"8F",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"EF",X"FC",X"0F",X"33",X"77",X"FF",X"FF",X"EF",X"0F",X"80",X"00",X"FC",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"0F",X"1E",X"DE",X"FF",X"FF",X"33",X"11",X"42",X"96",X"1E",X"BC",X"FC",X"FC",X"FC",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CF",X"FF",X"FF",X"FF",X"FF",X"0E",X"1E",X"FD",X"CF",X"1E",X"BC",X"FC",X"EC",X"1E",X"BC",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"01",X"00",X"00",X"00",X"00",X"44",X"EC",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"DF",X"CF",X"EF",X"77",X"11",X"00",X"8F",X"CF",X"FF",X"7F",X"7B",X"C0",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"77",X"FF",X"FF",X"FF",X"9F",X"0F",X"0E",X"00",X"00",X"88",X"CC",X"EC",X"EC",X"FC",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"EC",X"44",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EF",X"FF",X"FF",X"FF",X"FF",X"33",X"11",X"00",X"0F",X"CF",X"FF",X"FF",X"FF",X"CF",X"EF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"00",X"00",X"00",X"44",X"EC",X"EC",X"FC",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"66",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"FF",X"17",X"00",X"00",X"00",X"77",X"FF",X"EC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"EF",X"CF",X"DF",X"FF",X"FF",X"EF",X"ED",X"80",X"7B",X"7F",X"FF",X"CF",X"8F",X"0F",X"0F",
		X"00",X"00",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"33",X"11",X"0C",X"0F",X"1E",X"FC",X"FC",X"FC",X"FC",X"FC",X"ED",X"C7",X"1E",X"BC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"33",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"FF",X"FF",X"EF",X"9F",X"3F",X"77",X"77",X"0C",X"80",X"D1",X"F7",X"FF",X"FF",X"EF",X"8F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CF",X"FF",X"FF",X"FC",X"FC",X"FC",X"FC",X"FC",X"0C",X"C0",X"C0",X"00",X"CF",X"FF",X"77",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",
		X"47",X"8F",X"EF",X"FF",X"FF",X"FC",X"ED",X"FF",X"3F",X"E0",X"E0",X"C0",X"80",X"0C",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"1F",X"00",X"00",X"00",X"00",X"00",X"FC",X"FC",X"FC",X"FC",X"0F",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"EF",X"FC",X"0F",X"00",X"00",X"00",X"FF",X"FF",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"EF",X"FC",X"9E",X"07",X"EC",X"FF",X"FF",X"8F",X"0F",X"08",X"00",X"00",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"1E",X"BC",X"FF",X"FF",X"7F",X"1F",X"8F",X"07",X"1E",X"FC",X"FC",X"FC",X"FC",X"FC",X"EC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"FF",X"FF",X"FF",X"11",X"00",X"00",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"EC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"33",X"33",X"0F",X"FC",X"FC",X"E8",X"00",X"1E",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CF",X"FF",X"FF",X"FF",X"EC",X"07",X"9E",X"FC",X"3F",X"FF",X"FF",X"FF",X"11",X"00",X"00",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"8F",X"0F",X"08",X"00",X"00",X"11",X"FF",X"FC",X"FC",X"9E",X"03",X"EC",X"FC",X"FC",X"FC",
		X"07",X"9E",X"FC",X"EF",X"EF",X"FF",X"FF",X"FF",X"33",X"80",X"0C",X"0F",X"0F",X"8F",X"EF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
