library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity prog is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of prog is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"F3",X"C3",X"DF",X"0A",X"0F",X"C3",X"11",X"18",X"C3",X"09",X"14",X"23",X"22",
		X"C3",X"62",X"19",X"C3",X"06",X"04",X"00",X"23",X"C3",X"C5",X"0A",X"C9",X"C3",X"46",X"14",X"36",
		X"C3",X"E3",X"1B",X"C3",X"8A",X"18",X"73",X"59",X"C3",X"04",X"1C",X"C3",X"B4",X"07",X"34",X"3A",
		X"C3",X"1C",X"1A",X"C3",X"70",X"1E",X"21",X"FC",X"C3",X"92",X"14",X"91",X"07",X"01",X"1A",X"1A",
		X"A2",X"48",X"3E",X"06",X"32",X"FA",X"40",X"CD",X"5C",X"07",X"2A",X"FE",X"43",X"7D",X"E6",X"1F",
		X"FE",X"1A",X"38",X"02",X"D6",X"1A",X"6F",X"7C",X"E6",X"1F",X"FE",X"1A",X"38",X"02",X"D6",X"06",
		X"0F",X"0F",X"0F",X"67",X"E6",X"E0",X"B5",X"6F",X"7C",X"E6",X"03",X"67",X"11",X"A2",X"48",X"19",
		X"7D",X"E6",X"1F",X"FE",X"14",X"30",X"14",X"FE",X"0A",X"38",X"10",X"E5",X"29",X"29",X"29",X"7C",
		X"E1",X"E6",X"1F",X"FE",X"1B",X"30",X"04",X"FE",X"09",X"30",X"20",X"36",X"39",X"E5",X"CD",X"5C",
		X"07",X"E1",X"01",X"00",X"08",X"09",X"00",X"07",X"07",X"E6",X"07",X"28",X"0C",X"FE",X"03",X"38",
		X"04",X"36",X"F1",X"18",X"06",X"36",X"F5",X"18",X"02",X"36",X"F2",X"3A",X"FA",X"40",X"3D",X"32",
		X"FA",X"40",X"20",X"93",X"3E",X"01",X"F7",X"18",X"89",X"C9",X"00",X"CC",X"00",X"D0",X"00",X"D4",
		X"00",X"D8",X"00",X"DC",X"00",X"E0",X"00",X"E4",X"00",X"01",X"01",X"39",X"01",X"02",X"61",X"2E",
		X"01",X"02",X"3C",X"3D",X"01",X"02",X"3E",X"3F",X"01",X"02",X"40",X"41",X"01",X"02",X"42",X"43",
		X"01",X"02",X"44",X"45",X"01",X"02",X"46",X"47",X"CD",X"34",X"14",X"FD",X"BE",X"14",X"C0",X"FD",
		X"5E",X"15",X"FD",X"56",X"16",X"EB",X"E9",X"CD",X"34",X"14",X"2A",X"FE",X"40",X"01",X"17",X"00",
		X"09",X"06",X"05",X"BE",X"23",X"28",X"05",X"23",X"23",X"10",X"F8",X"C9",X"5E",X"23",X"56",X"EB",
		X"E9",X"21",X"29",X"01",X"18",X"08",X"21",X"2C",X"01",X"18",X"03",X"21",X"39",X"01",X"3E",X"2E",
		X"46",X"23",X"5E",X"23",X"56",X"12",X"10",X"F9",X"C9",X"01",X"92",X"4A",X"06",X"52",X"49",X"53",
		X"49",X"75",X"49",X"0C",X"4B",X"14",X"4B",X"51",X"49",X"06",X"C7",X"48",X"F6",X"48",X"49",X"49",
		X"4E",X"49",X"A4",X"49",X"03",X"4B",X"FD",X"21",X"09",X"18",X"3E",X"80",X"F7",X"C3",X"E5",X"12",
		X"3E",X"04",X"F7",X"2A",X"03",X"40",X"FD",X"21",X"89",X"01",X"7D",X"FE",X"A0",X"DA",X"0F",X"13",
		X"7C",X"FE",X"60",X"DA",X"E5",X"12",X"18",X"E8",X"C3",X"A9",X"23",X"C3",X"3D",X"27",X"C3",X"3D",
		X"27",X"CD",X"38",X"27",X"C3",X"A9",X"23",X"CD",X"38",X"27",X"C3",X"46",X"01",X"CD",X"42",X"27",
		X"C3",X"50",X"01",X"CD",X"3D",X"27",X"C3",X"46",X"01",X"4B",X"06",X"D9",X"15",X"68",X"10",X"5C",
		X"05",X"21",X"C3",X"49",X"11",X"9F",X"15",X"06",X"0B",X"40",X"0E",X"87",X"CD",X"19",X"00",X"21",
		X"C3",X"51",X"01",X"01",X"0D",X"3E",X"F5",X"CD",X"88",X"02",X"CD",X"B3",X"26",X"3A",X"15",X"40",
		X"FE",X"02",X"38",X"12",X"21",X"EC",X"49",X"11",X"0E",X"23",X"CD",X"87",X"0B",X"21",X"4A",X"49",
		X"11",X"15",X"23",X"CD",X"87",X"0B",X"3A",X"15",X"40",X"E6",X"0F",X"32",X"06",X"4B",X"3E",X"01",
		X"F7",X"01",X"08",X"00",X"E7",X"E7",X"DB",X"03",X"2F",X"E6",X"30",X"28",X"D0",X"E6",X"20",X"08",
		X"3A",X"15",X"40",X"47",X"08",X"28",X"09",X"05",X"05",X"FA",X"AD",X"01",X"3E",X"02",X"18",X"03",
		X"05",X"3E",X"01",X"32",X"C0",X"40",X"78",X"32",X"15",X"40",X"3E",X"01",X"32",X"CF",X"40",X"32",
		X"D0",X"40",X"CD",X"8C",X"22",X"CD",X"FA",X"1E",X"3E",X"00",X"32",X"C1",X"40",X"21",X"0D",X"41",
		X"01",X"18",X"00",X"CD",X"CE",X"15",X"21",X"C2",X"40",X"01",X"06",X"00",X"CD",X"CE",X"15",X"3A",
		X"27",X"43",X"6F",X"3A",X"21",X"43",X"67",X"C3",X"CB",X"42",X"DD",X"2A",X"28",X"02",X"CD",X"80",
		X"02",X"CD",X"02",X"21",X"CD",X"63",X"05",X"CD",X"5F",X"23",X"CD",X"C0",X"06",X"3E",X"20",X"F7",
		X"21",X"2E",X"06",X"11",X"02",X"40",X"01",X"03",X"00",X"ED",X"B0",X"21",X"ED",X"40",X"36",X"03",
		X"21",X"FC",X"40",X"7E",X"EE",X"01",X"77",X"CB",X"47",X"CA",X"5F",X"06",X"FD",X"21",X"83",X"1A",
		X"CD",X"32",X"04",X"3E",X"0F",X"D7",X"FD",X"21",X"D8",X"06",X"CD",X"F6",X"18",X"FD",X"7E",X"09",
		X"D7",X"CD",X"71",X"19",X"CD",X"7B",X"19",X"3E",X"20",X"F7",X"CD",X"10",X"1A",X"C3",X"94",X"12",
		X"21",X"80",X"48",X"01",X"20",X"1C",X"3E",X"2E",X"C5",X"E5",X"77",X"23",X"0D",X"20",X"FB",X"E1",
		X"01",X"20",X"00",X"09",X"C1",X"10",X"F1",X"C9",X"21",X"8A",X"73",X"71",X"23",X"70",X"2C",X"73",
		X"4E",X"0D",X"06",X"00",X"25",X"2E",X"7A",X"09",X"09",X"7E",X"23",X"46",X"21",X"8A",X"73",X"A6",
		X"2C",X"4F",X"78",X"A6",X"47",X"79",X"C9",X"21",X"8D",X"73",X"71",X"06",X"00",X"21",X"3C",X"71",
		X"09",X"7E",X"07",X"C9",X"21",X"8E",X"73",X"71",X"00",X"00",X"00",X"CD",X"25",X"24",X"CD",X"E3",
		X"06",X"CD",X"1B",X"04",X"CD",X"2E",X"25",X"FD",X"CB",X"00",X"56",X"28",X"05",X"11",X"C5",X"1B",
		X"18",X"03",X"11",X"D6",X"0B",X"FD",X"6E",X"02",X"FD",X"66",X"03",X"E5",X"CD",X"D0",X"14",X"E1",
		X"01",X"00",X"08",X"09",X"01",X"06",X"01",X"FD",X"7E",X"01",X"CD",X"88",X"02",X"3E",X"10",X"F7",
		X"FD",X"CB",X"00",X"66",X"28",X"32",X"3A",X"03",X"40",X"FD",X"BE",X"06",X"38",X"05",X"FD",X"BE",
		X"07",X"38",X"05",X"3E",X"02",X"F7",X"18",X"EE",X"FD",X"CB",X"00",X"F6",X"FD",X"CB",X"00",X"AE",
		X"CD",X"2E",X"25",X"FD",X"6E",X"02",X"FD",X"66",X"03",X"01",X"00",X"08",X"09",X"01",X"06",X"01",
		X"FD",X"7E",X"01",X"E6",X"F7",X"CD",X"88",X"02",X"FD",X"CB",X"00",X"56",X"28",X"05",X"11",X"CD",
		X"1B",X"18",X"03",X"11",X"DE",X"0B",X"FD",X"6E",X"02",X"FD",X"66",X"03",X"CD",X"D0",X"14",X"3E",
		X"04",X"F7",X"FD",X"6E",X"02",X"FD",X"66",X"03",X"FD",X"CB",X"00",X"56",X"28",X"0A",X"11",X"D5",
		X"1B",X"CD",X"D0",X"14",X"3E",X"7E",X"18",X"08",X"11",X"FC",X"0E",X"CD",X"D0",X"14",X"3E",X"93",
		X"FD",X"6E",X"04",X"FD",X"66",X"05",X"77",X"01",X"00",X"08",X"09",X"FD",X"7E",X"01",X"77",X"CD",
		X"1B",X"1B",X"3E",X"04",X"F7",X"FD",X"6E",X"04",X"FD",X"66",X"05",X"FD",X"CB",X"00",X"56",X"28",
		X"04",X"36",X"7F",X"18",X"02",X"36",X"94",X"3E",X"04",X"F7",X"FD",X"6E",X"04",X"FD",X"66",X"05",
		X"FD",X"CB",X"00",X"56",X"28",X"04",X"36",X"80",X"18",X"02",X"36",X"95",X"3E",X"04",X"F7",X"FD",
		X"6E",X"04",X"FD",X"66",X"05",X"FD",X"CB",X"00",X"56",X"28",X"0A",X"2B",X"11",X"DB",X"1B",X"E5",
		X"CD",X"D0",X"14",X"18",X"0B",X"01",X"DF",X"FF",X"09",X"11",X"02",X"0F",X"E5",X"CD",X"D0",X"14",
		X"E1",X"01",X"00",X"08",X"09",X"01",X"03",X"02",X"FD",X"7E",X"01",X"CD",X"88",X"02",X"3E",X"04",
		X"F7",X"FD",X"6E",X"04",X"FD",X"66",X"05",X"FD",X"CB",X"00",X"56",X"28",X"03",X"2B",X"18",X"04",
		X"01",X"DF",X"FF",X"09",X"01",X"03",X"02",X"CD",X"86",X"02",X"CD",X"C3",X"20",X"3E",X"20",X"F7",
		X"FD",X"CB",X"00",X"6E",X"CA",X"D7",X"02",X"FD",X"CB",X"00",X"AE",X"FD",X"CB",X"00",X"66",X"C2",
		X"D7",X"02",X"CD",X"95",X"18",X"FD",X"36",X"00",X"00",X"C9",X"CB",X"3A",X"03",X"40",X"FD",X"BE",
		X"06",X"38",X"0A",X"FD",X"BE",X"07",X"30",X"05",X"3E",X"02",X"F7",X"18",X"EE",X"FD",X"CB",X"00",
		X"EE",X"C9",X"FD",X"7E",X"00",X"A7",X"20",X"04",X"3E",X"0F",X"CF",X"C9",X"32",X"FD",X"40",X"FD",
		X"23",X"FD",X"7E",X"00",X"2A",X"03",X"40",X"CB",X"5F",X"C4",X"66",X"04",X"CB",X"57",X"C4",X"63",
		X"04",X"CB",X"4F",X"C4",X"60",X"04",X"CB",X"47",X"C4",X"5D",X"04",X"18",X"0E",X"2D",X"18",X"07",
		X"2C",X"18",X"04",X"24",X"18",X"01",X"25",X"22",X"03",X"40",X"C9",X"3A",X"FD",X"40",X"3D",X"32",
		X"FD",X"40",X"28",X"05",X"3E",X"01",X"F7",X"18",X"C8",X"FD",X"23",X"18",X"B5",X"81",X"09",X"E3",
		X"09",X"E6",X"12",X"E9",X"09",X"EC",X"09",X"EC",X"12",X"EC",X"09",X"EE",X"12",X"EC",X"12",X"E9",
		X"1B",X"E3",X"09",X"E6",X"12",X"E9",X"12",X"E9",X"12",X"E6",X"09",X"E6",X"09",X"E6",X"24",X"E3",
		X"00",X"3E",X"01",X"F7",X"01",X"08",X"00",X"E7",X"E7",X"DB",X"03",X"2F",X"E6",X"30",X"28",X"0A",
		X"CD",X"7B",X"19",X"3E",X"14",X"F7",X"3E",X"0A",X"CF",X"C9",X"21",X"7C",X"41",X"CD",X"02",X"1B",
		X"E6",X"02",X"BE",X"77",X"20",X"DB",X"23",X"BE",X"28",X"D7",X"77",X"A7",X"28",X"D3",X"3A",X"7B",
		X"41",X"FE",X"1C",X"28",X"3E",X"30",X"57",X"FE",X"1A",X"28",X"34",X"30",X"2E",X"4F",X"CB",X"21",
		X"06",X"00",X"21",X"F2",X"24",X"09",X"5E",X"23",X"56",X"13",X"1A",X"47",X"21",X"7E",X"41",X"7E",
		X"FE",X"0A",X"38",X"07",X"CD",X"7B",X"19",X"3E",X"0A",X"CF",X"C9",X"3C",X"77",X"5F",X"16",X"00",
		X"EB",X"19",X"70",X"21",X"07",X"4A",X"CD",X"87",X"0B",X"18",X"96",X"06",X"2E",X"18",X"DD",X"06",
		X"2D",X"18",X"D9",X"21",X"7E",X"41",X"7E",X"A7",X"CA",X"A1",X"04",X"E5",X"5F",X"16",X"00",X"EB",
		X"19",X"36",X"2E",X"21",X"07",X"4A",X"CD",X"87",X"0B",X"E1",X"35",X"C3",X"A1",X"04",X"CD",X"4C",
		X"26",X"3E",X"0B",X"D7",X"CD",X"7B",X"19",X"3E",X"0A",X"CF",X"C9",X"11",X"20",X"00",X"DD",X"7E",
		X"00",X"A7",X"C8",X"47",X"DD",X"23",X"DD",X"7E",X"00",X"FE",X"2E",X"28",X"08",X"77",X"19",X"10",
		X"FC",X"DD",X"23",X"18",X"E9",X"19",X"10",X"FD",X"DD",X"23",X"18",X"E2",X"82",X"FF",X"07",X"0B",
		X"08",X"2F",X"4B",X"21",X"7F",X"50",X"01",X"02",X"1D",X"3E",X"FF",X"CD",X"88",X"02",X"21",X"9D",
		X"50",X"01",X"02",X"1C",X"3E",X"F0",X"CD",X"88",X"02",X"21",X"9E",X"50",X"01",X"01",X"08",X"3E",
		X"F5",X"CD",X"88",X"02",X"21",X"FE",X"52",X"01",X"01",X"09",X"3E",X"F2",X"CD",X"88",X"02",X"21",
		X"81",X"50",X"01",X"1C",X"01",X"3E",X"F8",X"CD",X"88",X"02",X"21",X"A1",X"50",X"01",X"01",X"1A",
		X"CD",X"88",X"02",X"21",X"BC",X"50",X"01",X"01",X"1A",X"CD",X"88",X"02",X"21",X"E1",X"53",X"01",
		X"1C",X"01",X"CD",X"88",X"02",X"21",X"A2",X"50",X"01",X"1A",X"1A",X"3E",X"F1",X"CD",X"88",X"02",
		X"21",X"BE",X"48",X"11",X"8A",X"14",X"CD",X"87",X"0B",X"CD",X"70",X"26",X"CD",X"8C",X"24",X"CD",
		X"7D",X"24",X"3A",X"C0",X"40",X"CB",X"47",X"20",X"0C",X"21",X"1E",X"4B",X"11",X"C8",X"14",X"CD",
		X"87",X"0B",X"CD",X"94",X"24",X"DD",X"21",X"85",X"19",X"21",X"81",X"48",X"CD",X"B8",X"1F",X"DD",
		X"21",X"8C",X"19",X"21",X"A1",X"48",X"CD",X"3B",X"05",X"DD",X"21",X"8C",X"19",X"21",X"BC",X"48",
		X"CD",X"3B",X"05",X"DD",X"21",X"8F",X"19",X"21",X"E1",X"4B",X"CD",X"B8",X"1F",X"C9",X"94",X"F8",
		X"A9",X"48",X"CA",X"48",X"80",X"AC",X"98",X"F8",X"D6",X"4B",X"B7",X"4B",X"14",X"33",X"94",X"F8",
		X"89",X"49",X"AA",X"49",X"84",X"AC",X"98",X"F4",X"D6",X"4B",X"B7",X"4B",X"14",X"3C",X"64",X"D0",
		X"40",X"11",X"20",X"20",X"29",X"29",X"29",X"7C",X"07",X"07",X"07",X"E6",X"F0",X"B0",X"D6",X"20",
		X"ED",X"44",X"92",X"67",X"7D",X"B1",X"ED",X"44",X"93",X"6F",X"C9",X"92",X"EC",X"FF",X"0B",X"08",
		X"2F",X"4B",X"3A",X"BF",X"40",X"A7",X"C8",X"3A",X"15",X"40",X"A7",X"C8",X"C3",X"FB",X"0F",X"CD",
		X"38",X"27",X"FD",X"21",X"58",X"0B",X"CD",X"32",X"04",X"3E",X"0F",X"D7",X"21",X"26",X"06",X"11",
		X"39",X"41",X"CD",X"48",X"27",X"3E",X"01",X"D7",X"21",X"ED",X"40",X"36",X"00",X"CD",X"71",X"19",
		X"CD",X"7B",X"19",X"3E",X"F7",X"32",X"02",X"40",X"CD",X"80",X"02",X"3E",X"02",X"F7",X"CD",X"63",
		X"05",X"CD",X"5F",X"23",X"3E",X"07",X"32",X"02",X"40",X"3E",X"02",X"F7",X"CD",X"10",X"1A",X"FD",
		X"21",X"39",X"41",X"CD",X"75",X"1D",X"FD",X"21",X"59",X"41",X"CD",X"75",X"1D",X"3E",X"40",X"F7",
		X"CD",X"7B",X"19",X"CD",X"71",X"19",X"AF",X"32",X"39",X"41",X"32",X"59",X"41",X"C3",X"94",X"12",
		X"FD",X"21",X"CD",X"06",X"CD",X"F6",X"18",X"FD",X"7E",X"09",X"D7",X"18",X"F3",X"80",X"F9",X"40",
		X"0A",X"20",X"51",X"49",X"27",X"1C",X"10",X"08",X"80",X"F8",X"40",X"05",X"08",X"D6",X"48",X"D6",
		X"1F",X"11",X"66",X"01",X"06",X"20",X"E7",X"3E",X"30",X"F7",X"01",X"06",X"20",X"EF",X"C9",X"FD",
		X"20",X"68",X"18",X"05",X"20",X"3F",X"20",X"18",X"21",X"21",X"00",X"44",X"F9",X"EB",X"11",X"7C",
		X"01",X"E5",X"D5",X"3E",X"13",X"2A",X"FE",X"43",X"29",X"22",X"FE",X"43",X"01",X"15",X"83",X"09",
		X"30",X"03",X"22",X"FE",X"43",X"3D",X"20",X"ED",X"3A",X"FE",X"43",X"33",X"F5",X"1B",X"7A",X"B3",
		X"20",X"E1",X"0E",X"C8",X"06",X"15",X"CD",X"19",X"00",X"0E",X"80",X"06",X"02",X"CD",X"19",X"00",
		X"21",X"BF",X"14",X"4E",X"0C",X"11",X"7E",X"41",X"06",X"00",X"ED",X"B0",X"3E",X"FF",X"32",X"BF",
		X"40",X"06",X"07",X"0E",X"80",X"CD",X"19",X"00",X"01",X"06",X"01",X"E7",X"C3",X"4F",X"07",X"C3",
		X"4F",X"07",X"06",X"03",X"1A",X"BE",X"C0",X"1B",X"2B",X"10",X"F9",X"C9",X"2A",X"FE",X"43",X"29",
		X"17",X"17",X"AD",X"17",X"AD",X"1F",X"1F",X"2F",X"E6",X"01",X"B5",X"6F",X"22",X"FE",X"43",X"C9",
		X"84",X"06",X"01",X"01",X"00",X"88",X"49",X"B9",X"00",X"08",X"88",X"49",X"88",X"0C",X"01",X"01",
		X"AF",X"08",X"21",X"C4",X"40",X"11",X"18",X"40",X"CD",X"52",X"07",X"30",X"0A",X"08",X"3E",X"01",
		X"08",X"21",X"C2",X"40",X"CD",X"6F",X"08",X"21",X"C7",X"40",X"11",X"18",X"40",X"CD",X"52",X"07",
		X"30",X"0A",X"21",X"C5",X"40",X"CD",X"6F",X"08",X"08",X"3E",X"02",X"08",X"08",X"A7",X"CA",X"44",
		X"08",X"3D",X"32",X"C1",X"40",X"A7",X"28",X"05",X"CD",X"BE",X"15",X"18",X"03",X"CD",X"AD",X"15",
		X"21",X"7E",X"41",X"36",X"00",X"23",X"01",X"0A",X"00",X"3E",X"2E",X"CD",X"D0",X"15",X"CD",X"80",
		X"02",X"CD",X"63",X"05",X"21",X"37",X"49",X"0E",X"87",X"11",X"F7",X"23",X"06",X"0B",X"CD",X"19",
		X"00",X"21",X"46",X"49",X"11",X"0A",X"24",X"06",X"0B",X"0E",X"87",X"CD",X"19",X"00",X"21",X"C3",
		X"49",X"16",X"15",X"1E",X"9F",X"06",X"0B",X"0E",X"87",X"CD",X"19",X"00",X"3E",X"F5",X"01",X"01",
		X"0D",X"21",X"C3",X"51",X"CD",X"88",X"02",X"CD",X"B3",X"26",X"3E",X"0A",X"06",X"1A",X"21",X"F2",
		X"24",X"5E",X"23",X"56",X"23",X"13",X"12",X"3C",X"10",X"F7",X"5E",X"23",X"56",X"13",X"EB",X"11",
		X"1B",X"24",X"CD",X"87",X"0B",X"3E",X"01",X"F7",X"CD",X"52",X"0A",X"CD",X"CF",X"24",X"CD",X"A1",
		X"04",X"3E",X"0A",X"D7",X"21",X"7E",X"41",X"7E",X"A7",X"20",X"09",X"01",X"0B",X"00",X"11",X"BF",
		X"14",X"EB",X"ED",X"B0",X"CD",X"AD",X"15",X"01",X"06",X"02",X"EF",X"CD",X"71",X"19",X"CD",X"7B",
		X"19",X"3E",X"FF",X"32",X"BF",X"40",X"3A",X"15",X"40",X"A7",X"20",X"0F",X"3A",X"C6",X"42",X"6F",
		X"3A",X"A8",X"42",X"67",X"C3",X"CB",X"42",X"DD",X"2A",X"F0",X"42",X"C9",X"CD",X"78",X"08",X"11",
		X"16",X"40",X"01",X"03",X"00",X"ED",X"B0",X"C9",X"84",X"0B",X"01",X"02",X"00",X"15",X"4B",X"B9",
		X"00",X"09",X"15",X"4B",X"CD",X"4A",X"14",X"3A",X"06",X"40",X"E6",X"FE",X"D3",X"06",X"F6",X"01",
		X"D3",X"06",X"32",X"06",X"40",X"3A",X"ED",X"40",X"CB",X"47",X"28",X"0C",X"CD",X"6D",X"25",X"CD",
		X"94",X"1E",X"CD",X"9A",X"19",X"CD",X"C7",X"21",X"CD",X"84",X"15",X"CD",X"53",X"1F",X"CD",X"52",
		X"06",X"CD",X"AD",X"09",X"CD",X"A3",X"20",X"CD",X"3C",X"21",X"CD",X"62",X"20",X"CD",X"94",X"23",
		X"C9",X"40",X"49",X"88",X"18",X"02",X"01",X"3E",X"02",X"D7",X"CD",X"71",X"19",X"CD",X"7B",X"19",
		X"AF",X"32",X"04",X"41",X"01",X"05",X"FF",X"E7",X"01",X"06",X"78",X"EF",X"3A",X"C1",X"40",X"CB",
		X"47",X"20",X"05",X"3A",X"CF",X"40",X"18",X"03",X"3A",X"D0",X"40",X"FD",X"E5",X"FE",X"05",X"38",
		X"10",X"FE",X"09",X"38",X"06",X"FD",X"21",X"AD",X"10",X"18",X"0A",X"FD",X"21",X"38",X"13",X"18",
		X"04",X"FD",X"21",X"58",X"27",X"CD",X"0A",X"0F",X"FD",X"E1",X"FD",X"6E",X"12",X"FD",X"66",X"13",
		X"06",X"04",X"11",X"02",X"41",X"CD",X"9C",X"24",X"CD",X"E5",X"26",X"CD",X"92",X"09",X"3A",X"39",
		X"41",X"A7",X"28",X"2B",X"FD",X"21",X"39",X"41",X"E6",X"BF",X"32",X"39",X"41",X"AF",X"32",X"EF",
		X"40",X"32",X"EE",X"40",X"CD",X"95",X"18",X"CD",X"25",X"24",X"3A",X"39",X"41",X"E6",X"04",X"28",
		X"05",X"11",X"CD",X"1B",X"18",X"03",X"11",X"DE",X"0B",X"2A",X"3B",X"41",X"CD",X"D0",X"14",X"3E",
		X"0D",X"D7",X"3A",X"C1",X"40",X"CB",X"47",X"20",X"19",X"21",X"0D",X"41",X"01",X"12",X"00",X"CD",
		X"CE",X"15",X"3A",X"CF",X"40",X"3C",X"32",X"CF",X"40",X"3A",X"F0",X"40",X"3C",X"32",X"F0",X"40",
		X"18",X"1D",X"21",X"1F",X"41",X"01",X"12",X"00",X"CD",X"CE",X"15",X"3A",X"D0",X"40",X"3C",X"FE",
		X"11",X"38",X"02",X"3E",X"01",X"32",X"D0",X"40",X"3A",X"F1",X"40",X"3C",X"32",X"F1",X"40",X"C3",
		X"64",X"13",X"3E",X"20",X"F7",X"FD",X"2A",X"FE",X"40",X"FD",X"6E",X"08",X"FD",X"66",X"09",X"11",
		X"02",X"40",X"01",X"03",X"00",X"ED",X"B0",X"3E",X"03",X"32",X"ED",X"40",X"C9",X"01",X"08",X"02",
		X"3A",X"07",X"41",X"A7",X"20",X"0D",X"3A",X"15",X"40",X"FE",X"09",X"28",X"06",X"D2",X"00",X"00",
		X"E7",X"E7",X"C9",X"EF",X"EF",X"C9",X"01",X"F0",X"48",X"21",X"07",X"23",X"DF",X"C9",X"06",X"06",
		X"3A",X"C1",X"40",X"CB",X"47",X"20",X"06",X"DD",X"21",X"0D",X"41",X"18",X"04",X"DD",X"21",X"1F",
		X"41",X"DD",X"7E",X"00",X"CB",X"7F",X"C8",X"DD",X"5E",X"01",X"DD",X"56",X"02",X"DD",X"23",X"DD",
		X"23",X"DD",X"23",X"EB",X"FE",X"80",X"20",X"0A",X"7E",X"FE",X"39",X"20",X"02",X"36",X"2E",X"10",
		X"E0",X"C9",X"CB",X"5F",X"20",X"17",X"CB",X"57",X"20",X"0E",X"CB",X"4F",X"20",X"05",X"11",X"01",
		X"00",X"18",X"0D",X"11",X"FF",X"FF",X"18",X"08",X"11",X"E0",X"FF",X"18",X"03",X"11",X"20",X"00",
		X"7E",X"FE",X"39",X"28",X"07",X"FE",X"2E",X"20",X"B8",X"19",X"18",X"F4",X"36",X"2E",X"18",X"B1",
		X"AF",X"32",X"C1",X"40",X"3E",X"01",X"32",X"F0",X"40",X"32",X"CF",X"40",X"32",X"D0",X"40",X"3C",
		X"32",X"C0",X"40",X"CD",X"80",X"02",X"CD",X"02",X"21",X"CD",X"63",X"05",X"CD",X"5F",X"23",X"C3",
		X"94",X"12",X"3E",X"10",X"32",X"7B",X"41",X"CD",X"88",X"0A",X"3E",X"06",X"F7",X"CD",X"02",X"1B",
		X"E6",X"0C",X"28",X"F6",X"08",X"3E",X"2E",X"CD",X"9A",X"0A",X"CB",X"39",X"08",X"E6",X"04",X"20",
		X"08",X"79",X"FE",X"1D",X"30",X"08",X"3C",X"18",X"05",X"79",X"A7",X"28",X"01",X"3D",X"32",X"7B",
		X"41",X"3E",X"29",X"CD",X"9A",X"0A",X"18",X"D2",X"3E",X"29",X"CD",X"9A",X"0A",X"3E",X"04",X"F7",
		X"3E",X"2E",X"CD",X"9A",X"0A",X"3E",X"04",X"F7",X"18",X"EE",X"21",X"F2",X"24",X"ED",X"4B",X"7B",
		X"41",X"06",X"00",X"CB",X"21",X"09",X"5E",X"23",X"56",X"12",X"C9",X"82",X"FF",X"05",X"1A",X"1A",
		X"DB",X"4B",X"21",X"CE",X"48",X"01",X"03",X"17",X"CD",X"86",X"02",X"CD",X"F6",X"18",X"FD",X"7E",
		X"09",X"D7",X"3E",X"20",X"F7",X"3E",X"04",X"CF",X"C9",X"81",X"F8",X"40",X"05",X"0A",X"EF",X"48",
		X"25",X"23",X"06",X"08",X"81",X"F8",X"40",X"05",X"0A",X"EF",X"48",X"3B",X"23",X"06",X"08",X"ED",
		X"56",X"21",X"A8",X"1F",X"11",X"00",X"40",X"01",X"10",X"00",X"ED",X"B0",X"21",X"00",X"40",X"01",
		X"FF",X"10",X"0C",X"ED",X"A3",X"20",X"FB",X"DB",X"0E",X"C3",X"7B",X"0D",X"3E",X"80",X"D3",X"06",
		X"DB",X"0E",X"C3",X"82",X"0D",X"07",X"07",X"07",X"B3",X"5F",X"AF",X"D3",X"06",X"D3",X"0C",X"7B",
		X"EE",X"18",X"5F",X"08",X"0E",X"0B",X"21",X"9F",X"15",X"46",X"23",X"ED",X"B3",X"DB",X"03",X"E6",
		X"F0",X"0F",X"0F",X"0F",X"0F",X"57",X"3E",X"01",X"D3",X"0A",X"DB",X"03",X"E6",X"F0",X"B2",X"57",
		X"AF",X"D3",X"0A",X"7A",X"EE",X"02",X"57",X"FB",X"08",X"C2",X"F1",X"06",X"08",X"C2",X"5F",X"63",
		X"31",X"00",X"44",X"CD",X"C8",X"15",X"3E",X"01",X"D3",X"06",X"C3",X"4A",X"0B",X"81",X"F8",X"40",
		X"05",X"0A",X"6F",X"49",X"51",X"23",X"06",X"08",X"80",X"00",X"30",X"04",X"80",X"00",X"10",X"01",
		X"20",X"00",X"30",X"04",X"20",X"00",X"20",X"04",X"40",X"00",X"0C",X"05",X"C0",X"00",X"28",X"01",
		X"10",X"00",X"04",X"01",X"38",X"04",X"80",X"00",X"08",X"01",X"60",X"00",X"20",X"01",X"C0",X"00",
		X"30",X"01",X"FF",X"00",X"80",X"00",X"00",X"1A",X"A7",X"C8",X"47",X"13",X"1A",X"77",X"C5",X"01",
		X"20",X"00",X"09",X"C1",X"13",X"10",X"F5",X"C9",X"FD",X"2A",X"FE",X"40",X"FD",X"6E",X"0C",X"FD",
		X"66",X"0D",X"11",X"D9",X"40",X"06",X"00",X"4E",X"23",X"ED",X"B0",X"21",X"D9",X"40",X"22",X"D7",
		X"40",X"FD",X"6E",X"0E",X"FD",X"66",X"0F",X"22",X"D5",X"40",X"2A",X"03",X"40",X"7C",X"D6",X"08",
		X"E6",X"F8",X"67",X"7D",X"D6",X"08",X"E6",X"F8",X"6F",X"22",X"D2",X"40",X"AF",X"32",X"D4",X"40",
		X"3E",X"01",X"32",X"D1",X"40",X"C9",X"06",X"01",X"85",X"86",X"87",X"88",X"89",X"8A",X"06",X"01",
		X"8B",X"8C",X"8D",X"8E",X"89",X"8A",X"11",X"89",X"41",X"01",X"07",X"00",X"ED",X"B0",X"11",X"90",
		X"41",X"21",X"8C",X"41",X"01",X"04",X"00",X"ED",X"B0",X"2A",X"8E",X"41",X"22",X"94",X"41",X"3A",
		X"89",X"41",X"E6",X"06",X"3A",X"8B",X"41",X"20",X"1E",X"3D",X"E6",X"07",X"87",X"4F",X"87",X"81",
		X"4F",X"06",X"00",X"3A",X"89",X"41",X"E6",X"0C",X"20",X"08",X"21",X"1C",X"26",X"09",X"22",X"96",
		X"41",X"C9",X"21",X"E8",X"14",X"18",X"F6",X"E6",X"07",X"3C",X"87",X"4F",X"87",X"81",X"3D",X"18",
		X"DF",X"3A",X"89",X"41",X"CB",X"57",X"C2",X"55",X"0E",X"CB",X"5F",X"C2",X"AB",X"0D",X"CB",X"4F",
		X"C2",X"DF",X"0C",X"3E",X"01",X"F7",X"ED",X"5B",X"92",X"41",X"3A",X"8B",X"41",X"E6",X"07",X"FE",
		X"01",X"28",X"61",X"1A",X"FE",X"2E",X"28",X"0C",X"06",X"03",X"2A",X"96",X"41",X"BE",X"28",X"17",
		X"23",X"23",X"10",X"F9",X"01",X"20",X"00",X"EB",X"09",X"3A",X"91",X"41",X"3D",X"28",X"0D",X"32",
		X"91",X"41",X"22",X"92",X"41",X"18",X"CF",X"23",X"7E",X"12",X"18",X"E8",X"3A",X"90",X"41",X"3D",
		X"28",X"15",X"32",X"90",X"41",X"3A",X"8D",X"41",X"32",X"91",X"41",X"2A",X"94",X"41",X"23",X"22",
		X"94",X"41",X"22",X"92",X"41",X"18",X"AC",X"3A",X"8B",X"41",X"3C",X"47",X"3A",X"8A",X"41",X"B8",
		X"28",X"09",X"78",X"32",X"8B",X"41",X"CD",X"EE",X"0B",X"18",X"98",X"21",X"89",X"41",X"CB",X"BE",
		X"3E",X"05",X"CF",X"C9",X"1A",X"FE",X"39",X"28",X"18",X"FE",X"2E",X"20",X"A7",X"1B",X"1A",X"FE",
		X"6F",X"28",X"0A",X"FE",X"55",X"28",X"06",X"3E",X"2E",X"13",X"12",X"18",X"97",X"3E",X"54",X"18",
		X"F8",X"1B",X"1A",X"FE",X"2E",X"28",X"04",X"3E",X"6F",X"18",X"EE",X"3E",X"55",X"18",X"EA",X"3E",
		X"01",X"F7",X"ED",X"5B",X"92",X"41",X"3A",X"8B",X"41",X"E6",X"07",X"FE",X"06",X"28",X"61",X"1A",
		X"FE",X"2E",X"28",X"0C",X"06",X"03",X"2A",X"96",X"41",X"BE",X"28",X"17",X"2B",X"2B",X"10",X"F9",
		X"01",X"E0",X"FF",X"EB",X"09",X"3A",X"91",X"41",X"3D",X"28",X"0D",X"32",X"91",X"41",X"22",X"92",
		X"41",X"18",X"CF",X"2B",X"7E",X"12",X"18",X"E8",X"3A",X"90",X"41",X"3D",X"28",X"15",X"32",X"90",
		X"41",X"3A",X"8D",X"41",X"32",X"91",X"41",X"2A",X"94",X"41",X"2B",X"22",X"92",X"41",X"22",X"94",
		X"41",X"18",X"AC",X"3A",X"8B",X"41",X"3D",X"47",X"3A",X"8A",X"41",X"B8",X"28",X"09",X"78",X"32",
		X"8B",X"41",X"CD",X"EE",X"0B",X"18",X"98",X"21",X"89",X"41",X"CB",X"BE",X"3E",X"05",X"CF",X"C9",
		X"1A",X"FE",X"69",X"28",X"18",X"FE",X"2E",X"20",X"A7",X"13",X"1A",X"FE",X"6A",X"28",X"0A",X"FE",
		X"4A",X"28",X"06",X"3E",X"2E",X"1B",X"12",X"18",X"97",X"3E",X"4B",X"18",X"F8",X"13",X"1A",X"FE",
		X"2E",X"28",X"04",X"3E",X"6A",X"18",X"EE",X"3E",X"4A",X"18",X"EA",X"3C",X"E6",X"07",X"5F",X"C3",
		X"FC",X"0A",X"2F",X"E6",X"07",X"07",X"C3",X"05",X"0B",X"FD",X"73",X"4E",X"CD",X"C4",X"43",X"5F",
		X"21",X"DF",X"70",X"4E",X"06",X"00",X"CD",X"98",X"43",X"2E",X"ED",X"77",X"2E",X"FA",X"4E",X"2C",
		X"46",X"2E",X"EE",X"71",X"23",X"70",X"2E",X"FD",X"4E",X"06",X"C8",X"3E",X"01",X"F7",X"ED",X"5B",
		X"92",X"41",X"3A",X"8B",X"41",X"E6",X"07",X"FE",X"02",X"28",X"61",X"1A",X"FE",X"2E",X"28",X"0C",
		X"06",X"03",X"2A",X"96",X"41",X"BE",X"28",X"14",X"23",X"23",X"10",X"F9",X"13",X"3A",X"90",X"41",
		X"3D",X"28",X"0E",X"32",X"90",X"41",X"ED",X"53",X"92",X"41",X"18",X"D2",X"23",X"7E",X"12",X"18",
		X"EB",X"3A",X"91",X"41",X"3D",X"28",X"18",X"32",X"91",X"41",X"3A",X"8C",X"41",X"32",X"90",X"41",
		X"2A",X"94",X"41",X"01",X"20",X"00",X"09",X"22",X"94",X"41",X"22",X"92",X"41",X"18",X"AC",X"3A",
		X"8B",X"41",X"3C",X"47",X"3A",X"8A",X"41",X"B8",X"28",X"09",X"78",X"32",X"8B",X"41",X"CD",X"EE",
		X"0B",X"18",X"98",X"21",X"89",X"41",X"CB",X"BE",X"3E",X"05",X"CF",X"C9",X"1A",X"FE",X"61",X"28",
		X"22",X"FE",X"2E",X"20",X"A7",X"EB",X"01",X"E0",X"FF",X"01",X"E0",X"FF",X"09",X"7E",X"FE",X"62",
		X"28",X"0D",X"FE",X"3C",X"28",X"09",X"3E",X"2E",X"A7",X"ED",X"42",X"EB",X"12",X"18",X"8D",X"3E",
		X"3D",X"18",X"F5",X"EB",X"01",X"E0",X"FF",X"09",X"7E",X"FE",X"2E",X"28",X"04",X"3E",X"62",X"18",
		X"E7",X"3E",X"3C",X"18",X"E3",X"3E",X"01",X"F7",X"ED",X"5B",X"92",X"41",X"3A",X"8B",X"41",X"E6",
		X"07",X"FE",X"07",X"28",X"61",X"1A",X"FE",X"2E",X"28",X"0C",X"06",X"03",X"2A",X"96",X"41",X"BE",
		X"28",X"14",X"2B",X"2B",X"10",X"F9",X"1B",X"3A",X"90",X"41",X"3D",X"28",X"0E",X"32",X"90",X"41",
		X"ED",X"53",X"92",X"41",X"18",X"D2",X"2B",X"7E",X"12",X"18",X"EB",X"3A",X"91",X"41",X"3D",X"28",
		X"18",X"32",X"91",X"41",X"3A",X"8C",X"41",X"32",X"90",X"41",X"2A",X"94",X"41",X"01",X"E0",X"FF",
		X"09",X"22",X"92",X"41",X"22",X"94",X"41",X"18",X"AC",X"3A",X"8B",X"41",X"3D",X"47",X"3A",X"8A",
		X"41",X"B8",X"28",X"09",X"78",X"32",X"8B",X"41",X"CD",X"EE",X"0B",X"18",X"98",X"21",X"89",X"41",
		X"CB",X"BE",X"3E",X"05",X"CF",X"C9",X"1A",X"FE",X"39",X"28",X"1F",X"FE",X"2E",X"20",X"A7",X"EB",
		X"01",X"20",X"00",X"09",X"7E",X"FE",X"67",X"28",X"0D",X"FE",X"47",X"28",X"09",X"3E",X"2E",X"A7",
		X"ED",X"42",X"EB",X"12",X"18",X"90",X"3E",X"46",X"18",X"F5",X"EB",X"01",X"20",X"00",X"09",X"7E",
		X"FE",X"2E",X"28",X"04",X"3E",X"67",X"18",X"E7",X"3E",X"47",X"18",X"E3",X"04",X"01",X"8F",X"90",
		X"91",X"92",X"03",X"02",X"98",X"2E",X"99",X"2E",X"96",X"97",X"3A",X"04",X"41",X"E6",X"80",X"28",
		X"05",X"3E",X"0D",X"D7",X"18",X"F4",X"FD",X"7E",X"00",X"32",X"04",X"41",X"FD",X"23",X"FD",X"7E",
		X"01",X"D3",X"05",X"01",X"06",X"04",X"E7",X"3E",X"02",X"F7",X"3A",X"04",X"41",X"E6",X"01",X"28",
		X"04",X"01",X"06",X"04",X"EF",X"FD",X"7E",X"00",X"D6",X"02",X"F7",X"FD",X"23",X"FD",X"23",X"FD",
		X"7E",X"00",X"A7",X"20",X"D9",X"3E",X"FF",X"D3",X"05",X"01",X"06",X"04",X"EF",X"AF",X"32",X"04",
		X"41",X"3E",X"0D",X"CF",X"C9",X"CD",X"80",X"02",X"CD",X"02",X"21",X"CD",X"63",X"05",X"CD",X"5F",
		X"23",X"CD",X"E8",X"00",X"CD",X"CE",X"09",X"CD",X"98",X"0B",X"CD",X"E1",X"1F",X"3E",X"05",X"32",
		X"F8",X"40",X"FD",X"2A",X"FE",X"40",X"FD",X"6E",X"06",X"FD",X"66",X"07",X"01",X"01",X"05",X"CD",
		X"86",X"02",X"3E",X"08",X"F7",X"FD",X"2A",X"FE",X"40",X"FD",X"6E",X"06",X"FD",X"66",X"07",X"11",
		X"DB",X"1F",X"CD",X"87",X"0B",X"3E",X"08",X"F7",X"3A",X"F8",X"40",X"3D",X"32",X"F8",X"40",X"20",
		X"D1",X"3A",X"C1",X"40",X"CB",X"47",X"20",X"05",X"21",X"F0",X"40",X"18",X"03",X"21",X"F1",X"40",
		X"7E",X"D9",X"F5",X"CD",X"00",X"20",X"3E",X"2E",X"77",X"23",X"77",X"F1",X"3D",X"D9",X"77",X"FD",
		X"2A",X"FE",X"40",X"FD",X"6E",X"0A",X"FD",X"66",X"0B",X"11",X"02",X"40",X"01",X"03",X"00",X"ED",
		X"B0",X"3E",X"01",X"32",X"ED",X"40",X"21",X"00",X"02",X"22",X"F2",X"40",X"21",X"00",X"04",X"22",
		X"F4",X"40",X"2A",X"03",X"40",X"22",X"F6",X"40",X"3E",X"01",X"F7",X"01",X"C7",X"08",X"C5",X"CD",
		X"84",X"25",X"CD",X"F7",X"00",X"CD",X"11",X"1D",X"C3",X"1B",X"1F",X"AF",X"32",X"BF",X"40",X"CD",
		X"10",X"1A",X"CD",X"AD",X"15",X"CD",X"7B",X"19",X"CD",X"71",X"19",X"21",X"0D",X"41",X"01",X"24",
		X"00",X"CD",X"CE",X"15",X"CD",X"80",X"02",X"CD",X"63",X"05",X"21",X"37",X"49",X"11",X"41",X"1F",
		X"CD",X"87",X"0B",X"21",X"77",X"51",X"01",X"01",X"0D",X"3E",X"F4",X"CD",X"88",X"02",X"11",X"91",
		X"01",X"01",X"06",X"78",X"EF",X"01",X"05",X"FF",X"E7",X"01",X"06",X"02",X"E7",X"D5",X"AF",X"32",
		X"ED",X"40",X"32",X"EE",X"40",X"32",X"04",X"41",X"CD",X"DE",X"17",X"21",X"4E",X"49",X"11",X"8B",
		X"20",X"CD",X"87",X"0B",X"21",X"26",X"4A",X"11",X"9B",X"20",X"CD",X"87",X"0B",X"21",X"26",X"52",
		X"01",X"01",X"08",X"3E",X"F2",X"C3",X"88",X"02",X"91",X"09",X"01",X"0B",X"08",X"44",X"4A",X"06",
		X"08",X"0F",X"38",X"08",X"23",X"23",X"23",X"23",X"23",X"10",X"F6",X"C9",X"35",X"20",X"F5",X"C5",
		X"32",X"19",X"40",X"3E",X"FE",X"0F",X"10",X"FD",X"F3",X"DD",X"A6",X"00",X"DD",X"77",X"00",X"23",
		X"5E",X"23",X"56",X"23",X"4E",X"23",X"46",X"23",X"C5",X"FD",X"E1",X"EB",X"D5",X"DD",X"E5",X"11",
		X"A4",X"10",X"D5",X"E9",X"DD",X"E1",X"E1",X"3A",X"19",X"40",X"C1",X"18",X"CC",X"81",X"06",X"DD",
		X"06",X"D2",X"06",X"C9",X"06",X"E4",X"06",X"DD",X"06",X"D2",X"06",X"E1",X"06",X"DB",X"06",X"D2",
		X"06",X"E6",X"06",X"DB",X"06",X"D2",X"06",X"E4",X"06",X"DD",X"06",X"D2",X"06",X"EB",X"06",X"DD",
		X"06",X"D7",X"06",X"ED",X"06",X"E1",X"06",X"DB",X"06",X"EE",X"06",X"E4",X"06",X"DD",X"24",X"EE",
		X"00",X"AF",X"B1",X"5F",X"7E",X"D6",X"0A",X"D6",X"01",X"9F",X"B3",X"4F",X"7E",X"D6",X"06",X"D6",
		X"01",X"2A",X"03",X"40",X"7D",X"D6",X"08",X"A0",X"6F",X"7C",X"D6",X"08",X"A0",X"67",X"22",X"D2",
		X"40",X"DD",X"2A",X"D5",X"40",X"DD",X"CB",X"00",X"76",X"28",X"07",X"DD",X"E5",X"3E",X"02",X"CF",
		X"DD",X"E1",X"2A",X"D7",X"40",X"3A",X"D4",X"40",X"CB",X"47",X"C2",X"CD",X"11",X"CB",X"4F",X"C2",
		X"A9",X"11",X"CB",X"57",X"C2",X"7A",X"11",X"3A",X"D3",X"40",X"DD",X"BE",X"04",X"F5",X"DC",X"F1",
		X"11",X"F1",X"47",X"3A",X"D4",X"40",X"CB",X"9F",X"32",X"D4",X"40",X"DD",X"CB",X"00",X"5E",X"28",
		X"2C",X"78",X"BE",X"30",X"1F",X"70",X"DD",X"4E",X"01",X"06",X"00",X"21",X"3B",X"1B",X"09",X"5E",
		X"23",X"56",X"C5",X"FD",X"E5",X"D5",X"FD",X"E1",X"CD",X"0A",X"0F",X"FD",X"E1",X"C1",X"CD",X"B2",
		X"22",X"CD",X"85",X"24",X"3A",X"D4",X"40",X"E6",X"0F",X"C2",X"01",X"11",X"C9",X"DD",X"CB",X"00",
		X"56",X"28",X"F1",X"7E",X"B8",X"30",X"ED",X"70",X"18",X"EA",X"3A",X"D3",X"40",X"DD",X"BE",X"02",
		X"28",X"05",X"F5",X"D4",X"0D",X"12",X"F1",X"47",X"3A",X"D4",X"40",X"CB",X"97",X"32",X"D4",X"40",
		X"DD",X"CB",X"00",X"56",X"28",X"06",X"7E",X"B8",X"30",X"CA",X"18",X"A9",X"DD",X"CB",X"00",X"5E",
		X"28",X"C2",X"78",X"BE",X"30",X"BE",X"70",X"18",X"BB",X"3A",X"D2",X"40",X"DD",X"BE",X"06",X"28",
		X"05",X"F5",X"D4",X"17",X"12",X"F1",X"47",X"3A",X"D4",X"40",X"CB",X"8F",X"32",X"D4",X"40",X"DD",
		X"CB",X"00",X"4E",X"28",X"02",X"18",X"CF",X"DD",X"CB",X"00",X"46",X"18",X"D3",X"3A",X"D2",X"40",
		X"DD",X"BE",X"08",X"F5",X"DC",X"12",X"12",X"F1",X"47",X"3A",X"D4",X"40",X"CB",X"87",X"32",X"D4",
		X"40",X"DD",X"CB",X"00",X"46",X"28",X"03",X"C3",X"41",X"11",X"DD",X"CB",X"00",X"4E",X"C3",X"71",
		X"11",X"DD",X"7E",X"05",X"A7",X"F2",X"30",X"12",X"CB",X"BF",X"21",X"00",X"28",X"06",X"00",X"4F",
		X"09",X"3A",X"D2",X"40",X"BE",X"38",X"01",X"23",X"23",X"7E",X"7E",X"18",X"23",X"DD",X"7E",X"03",
		X"18",X"E2",X"DD",X"7E",X"09",X"18",X"03",X"DD",X"7E",X"07",X"A7",X"F2",X"30",X"12",X"CB",X"BF",
		X"21",X"00",X"28",X"06",X"00",X"4F",X"09",X"3A",X"D3",X"40",X"BE",X"38",X"01",X"23",X"23",X"7E",
		X"32",X"D1",X"40",X"FD",X"2A",X"FE",X"40",X"DD",X"21",X"00",X"00",X"FD",X"4E",X"0E",X"FD",X"46",
		X"0F",X"DD",X"09",X"A7",X"20",X"03",X"76",X"00",X"00",X"3D",X"87",X"4F",X"87",X"87",X"81",X"4F",
		X"06",X"00",X"DD",X"09",X"DD",X"22",X"D5",X"40",X"3A",X"D1",X"40",X"4F",X"21",X"D8",X"40",X"09",
		X"22",X"D7",X"40",X"C9",X"06",X"00",X"21",X"44",X"72",X"09",X"09",X"7E",X"23",X"46",X"21",X"22",
		X"74",X"77",X"23",X"70",X"2E",X"21",X"4E",X"CD",X"93",X"52",X"6F",X"26",X"00",X"C3",X"48",X"54",
		X"2A",X"22",X"74",X"36",X"FF",X"C3",X"5E",X"54",X"2A",X"22",X"74",X"36",X"00",X"C3",X"5E",X"54",
		X"01",X"24",X"74",X"CD",X"21",X"2A",X"49",X"01",X"0A",X"12",X"CD",X"86",X"02",X"3E",X"80",X"F7",
		X"21",X"51",X"49",X"11",X"27",X"1C",X"CD",X"87",X"0B",X"21",X"51",X"51",X"01",X"01",X"0F",X"3E",
		X"F0",X"CD",X"88",X"02",X"21",X"2E",X"49",X"11",X"41",X"1F",X"CD",X"87",X"0B",X"21",X"2E",X"51",
		X"01",X"01",X"11",X"3E",X"F4",X"CD",X"88",X"02",X"3E",X"40",X"F7",X"CD",X"42",X"00",X"FD",X"21",
		X"CD",X"06",X"CD",X"F6",X"18",X"FD",X"7E",X"09",X"D7",X"CD",X"71",X"19",X"CD",X"7B",X"19",X"3E",
		X"40",X"F7",X"C3",X"2E",X"02",X"FD",X"6E",X"00",X"FD",X"66",X"01",X"11",X"89",X"41",X"CD",X"E6",
		X"0B",X"CD",X"31",X"0C",X"3E",X"05",X"D7",X"3E",X"08",X"F7",X"FD",X"6E",X"02",X"FD",X"66",X"03",
		X"11",X"89",X"41",X"CD",X"E6",X"0B",X"CD",X"31",X"0C",X"3E",X"05",X"D7",X"3E",X"08",X"F7",X"FD",
		X"6E",X"04",X"FD",X"66",X"05",X"11",X"89",X"41",X"CD",X"E6",X"0B",X"CD",X"31",X"0C",X"3E",X"05",
		X"D7",X"FD",X"6E",X"06",X"FD",X"66",X"07",X"11",X"89",X"41",X"CD",X"E6",X"0B",X"CD",X"31",X"0C",
		X"3E",X"05",X"D7",X"3E",X"08",X"F7",X"18",X"AD",X"81",X"0A",X"E7",X"0A",X"E9",X"0A",X"EB",X"0A",
		X"E1",X"0A",X"E4",X"0A",X"E7",X"0A",X"E4",X"0A",X"E7",X"0A",X"E9",X"0A",X"DF",X"0A",X"E1",X"0A",
		X"E4",X"1E",X"E1",X"00",X"88",X"53",X"90",X"53",X"B2",X"53",X"D0",X"53",X"EB",X"53",X"21",X"21",
		X"74",X"7E",X"D6",X"10",X"CD",X"7B",X"19",X"CD",X"71",X"19",X"01",X"06",X"78",X"EF",X"AF",X"32",
		X"ED",X"40",X"AF",X"32",X"EE",X"40",X"32",X"EF",X"40",X"32",X"39",X"41",X"32",X"59",X"41",X"32",
		X"98",X"41",X"32",X"A4",X"41",X"32",X"89",X"41",X"32",X"04",X"41",X"32",X"06",X"41",X"CD",X"10",
		X"1A",X"CD",X"80",X"02",X"CD",X"63",X"05",X"C3",X"9A",X"13",X"21",X"72",X"49",X"11",X"E0",X"15",
		X"CD",X"87",X"0B",X"21",X"72",X"51",X"01",X"01",X"0E",X"3E",X"F4",X"CD",X"88",X"02",X"3A",X"C1",
		X"40",X"CB",X"47",X"20",X"05",X"11",X"EF",X"15",X"18",X"03",X"11",X"F8",X"15",X"21",X"CF",X"49",
		X"CD",X"87",X"0B",X"21",X"CC",X"49",X"11",X"01",X"16",X"CD",X"87",X"0B",X"21",X"CC",X"51",X"01",
		X"01",X"08",X"3E",X"F0",X"CD",X"88",X"02",X"3E",X"10",X"F7",X"3A",X"C1",X"40",X"CB",X"47",X"20",
		X"05",X"3A",X"CF",X"40",X"18",X"03",X"3A",X"D0",X"40",X"CD",X"8D",X"21",X"32",X"0A",X"41",X"0F",
		X"0F",X"0F",X"0F",X"E6",X"0F",X"20",X"02",X"3E",X"2E",X"32",X"8C",X"4A",X"3E",X"08",X"F7",X"3A",
		X"0A",X"41",X"E6",X"0F",X"32",X"AC",X"4A",X"3A",X"C1",X"40",X"CB",X"47",X"20",X"05",X"21",X"0D",
		X"41",X"18",X"03",X"21",X"1F",X"41",X"7E",X"E6",X"80",X"20",X"09",X"CD",X"42",X"00",X"FD",X"21",
		X"7D",X"04",X"18",X"04",X"FD",X"21",X"A1",X"21",X"CD",X"0A",X"0F",X"3E",X"0D",X"D7",X"CD",X"7B",
		X"19",X"C3",X"55",X"0F",X"3A",X"C1",X"40",X"CB",X"47",X"20",X"05",X"3A",X"CF",X"40",X"18",X"03",
		X"3A",X"D0",X"40",X"FE",X"11",X"D8",X"D6",X"10",X"18",X"F9",X"21",X"02",X"40",X"3A",X"05",X"41",
		X"A7",X"28",X"13",X"7E",X"C6",X"08",X"D3",X"02",X"23",X"7E",X"2F",X"D6",X"20",X"D3",X"03",X"23",
		X"7E",X"2F",X"D3",X"04",X"18",X"0B",X"7E",X"D3",X"02",X"23",X"7E",X"D3",X"03",X"23",X"7E",X"D3",
		X"04",X"DD",X"21",X"C8",X"40",X"DB",X"02",X"DD",X"77",X"00",X"DB",X"06",X"DD",X"77",X"01",X"DB",
		X"0A",X"DD",X"77",X"02",X"DB",X"0E",X"DD",X"77",X"03",X"C9",X"07",X"1C",X"0C",X"18",X"1B",X"0E",
		X"29",X"01",X"FD",X"E5",X"DD",X"E5",X"C5",X"D5",X"E5",X"F5",X"08",X"D9",X"C5",X"D5",X"E5",X"F5",
		X"3A",X"87",X"42",X"6F",X"3A",X"A1",X"42",X"67",X"CD",X"D8",X"43",X"AF",X"32",X"00",X"48",X"F1",
		X"E1",X"D1",X"C1",X"D9",X"08",X"F1",X"E1",X"D1",X"C1",X"DD",X"E1",X"FD",X"E1",X"FB",X"C9",X"08",
		X"11",X"12",X"29",X"1C",X"0C",X"18",X"1B",X"0E",X"07",X"1C",X"0C",X"18",X"1B",X"0E",X"29",X"02",
		X"1A",X"4F",X"13",X"1A",X"47",X"13",X"C5",X"E5",X"1A",X"77",X"23",X"13",X"0D",X"20",X"F9",X"E1",
		X"01",X"20",X"00",X"09",X"C1",X"10",X"EF",X"C9",X"39",X"61",X"39",X"61",X"39",X"61",X"61",X"62",
		X"61",X"3C",X"2E",X"3D",X"62",X"63",X"3C",X"3E",X"3D",X"3F",X"63",X"64",X"3E",X"40",X"3F",X"41",
		X"64",X"65",X"40",X"42",X"41",X"43",X"65",X"66",X"42",X"44",X"43",X"45",X"66",X"67",X"44",X"46",
		X"45",X"47",X"67",X"39",X"46",X"2E",X"47",X"39",X"3A",X"ED",X"40",X"E6",X"02",X"20",X"5B",X"2A",
		X"D5",X"40",X"FD",X"2A",X"FE",X"40",X"CB",X"7E",X"28",X"16",X"3A",X"06",X"41",X"A7",X"20",X"4A",
		X"FD",X"6E",X"0A",X"FD",X"66",X"0B",X"11",X"02",X"40",X"01",X"03",X"00",X"ED",X"B0",X"18",X"35",
		X"CB",X"76",X"28",X"36",X"7E",X"32",X"01",X"48",X"3A",X"33",X"43",X"6F",X"3A",X"6F",X"43",X"67",
		X"CD",X"D8",X"43",X"1A",X"FE",X"36",X"38",X"0C",X"FE",X"70",X"30",X"08",X"FE",X"56",X"38",X"1A",
		X"FE",X"60",X"30",X"16",X"FD",X"6E",X"08",X"FD",X"66",X"09",X"11",X"02",X"40",X"01",X"03",X"00",
		X"ED",X"B0",X"3E",X"02",X"CF",X"AF",X"32",X"CC",X"40",X"C9",X"DB",X"02",X"E6",X"10",X"28",X"F5",
		X"3E",X"01",X"CF",X"C9",X"DD",X"21",X"1A",X"40",X"21",X"1C",X"40",X"DD",X"7E",X"00",X"A7",X"C4",
		X"6F",X"10",X"DD",X"23",X"21",X"44",X"40",X"DD",X"7E",X"00",X"A7",X"C4",X"6F",X"10",X"C9",X"0D",
		X"B2",X"2E",X"1D",X"0A",X"12",X"1D",X"18",X"2E",X"0C",X"18",X"1B",X"19",X"2D",X"DB",X"00",X"CB",
		X"4F",X"20",X"0B",X"01",X"08",X"01",X"E7",X"E7",X"3E",X"FF",X"32",X"05",X"41",X"C9",X"01",X"08",
		X"01",X"EF",X"EF",X"AF",X"32",X"05",X"41",X"C9",X"21",X"10",X"40",X"01",X"F0",X"01",X"3E",X"00",
		X"57",X"72",X"23",X"0B",X"78",X"B1",X"20",X"F9",X"C9",X"81",X"01",X"EE",X"0B",X"08",X"44",X"4A",
		X"0E",X"15",X"0E",X"1D",X"B8",X"1C",X"2E",X"0A",X"1D",X"1D",X"0A",X"0C",X"14",X"2E",X"B3",X"08",
		X"19",X"15",X"0A",X"22",X"0E",X"1B",X"2E",X"01",X"08",X"19",X"15",X"0A",X"22",X"0E",X"1B",X"2E",
		X"02",X"06",X"15",X"0E",X"1F",X"0E",X"15",X"2C",X"06",X"00",X"21",X"C7",X"26",X"09",X"3A",X"C1",
		X"40",X"CB",X"47",X"20",X"05",X"11",X"C2",X"40",X"18",X"03",X"11",X"C5",X"40",X"06",X"03",X"AF",
		X"1A",X"8E",X"27",X"12",X"13",X"23",X"10",X"F8",X"C9",X"06",X"00",X"21",X"C7",X"26",X"09",X"3A",
		X"C1",X"40",X"CB",X"47",X"20",X"05",X"11",X"C2",X"40",X"18",X"03",X"11",X"C5",X"40",X"06",X"03",
		X"AF",X"1A",X"9E",X"27",X"12",X"13",X"23",X"10",X"F8",X"1B",X"20",X"01",X"C9",X"AF",X"12",X"1B",
		X"12",X"1B",X"12",X"37",X"C9",X"DD",X"FD",X"E5",X"D1",X"01",X"04",X"00",X"18",X"06",X"FD",X"E5",
		X"D1",X"01",X"0C",X"00",X"ED",X"B0",X"FD",X"6E",X"05",X"FD",X"66",X"06",X"7E",X"FE",X"39",X"20",
		X"07",X"FD",X"46",X"00",X"CB",X"78",X"20",X"0C",X"3E",X"01",X"F7",X"FD",X"CB",X"00",X"BE",X"FD",
		X"7E",X"09",X"CF",X"C9",X"FD",X"6E",X"05",X"FD",X"66",X"06",X"FD",X"7E",X"04",X"CB",X"58",X"C2",
		X"D2",X"16",X"CB",X"50",X"C2",X"5D",X"17",X"CB",X"48",X"C2",X"0D",X"17",X"FD",X"86",X"02",X"CB",
		X"5F",X"20",X"0C",X"FD",X"77",X"04",X"CD",X"C9",X"17",X"FD",X"7E",X"03",X"F7",X"18",X"C2",X"E6",
		X"07",X"FD",X"77",X"04",X"E5",X"23",X"CD",X"C3",X"17",X"CD",X"B5",X"17",X"11",X"20",X"00",X"E1",
		X"36",X"2E",X"19",X"10",X"FB",X"FD",X"7E",X"05",X"E6",X"1F",X"FD",X"BE",X"01",X"30",X"AC",X"C3",
		X"A9",X"16",X"FD",X"86",X"02",X"CB",X"5F",X"20",X"08",X"FD",X"77",X"04",X"CD",X"C9",X"17",X"18",
		X"C8",X"E6",X"07",X"FD",X"77",X"04",X"E5",X"11",X"20",X"00",X"19",X"CD",X"C3",X"17",X"CD",X"B5",
		X"17",X"E1",X"36",X"2E",X"23",X"0D",X"20",X"FA",X"FD",X"6E",X"05",X"FD",X"66",X"06",X"29",X"29",
		X"29",X"7C",X"E6",X"1F",X"FD",X"BE",X"01",X"D2",X"7B",X"16",X"C3",X"A9",X"16",X"FD",X"96",X"02",
		X"FA",X"1C",X"17",X"20",X"21",X"FD",X"BE",X"04",X"28",X"1C",X"18",X"25",X"08",X"7D",X"E6",X"1F",
		X"5F",X"FD",X"7E",X"01",X"BB",X"D2",X"7B",X"16",X"2B",X"08",X"E6",X"07",X"28",X"15",X"4F",X"FD",
		X"7E",X"04",X"A7",X"79",X"20",X"0D",X"E6",X"07",X"FD",X"77",X"04",X"CD",X"C3",X"17",X"C3",X"A9",
		X"16",X"E6",X"07",X"FD",X"77",X"04",X"E5",X"CD",X"C3",X"17",X"CD",X"B5",X"17",X"E1",X"11",X"20",
		X"00",X"23",X"0D",X"20",X"FC",X"36",X"2E",X"19",X"10",X"FB",X"C3",X"A9",X"16",X"FD",X"96",X"02",
		X"FA",X"6C",X"17",X"20",X"29",X"FD",X"BE",X"04",X"28",X"24",X"18",X"2D",X"08",X"5D",X"54",X"29",
		X"29",X"29",X"7C",X"E6",X"1F",X"6F",X"FD",X"7E",X"01",X"BD",X"D2",X"7B",X"16",X"21",X"E0",X"FF",
		X"19",X"08",X"E6",X"07",X"28",X"15",X"4F",X"FD",X"7E",X"04",X"A7",X"79",X"20",X"0D",X"E6",X"07",
		X"FD",X"77",X"04",X"CD",X"C3",X"17",X"C3",X"A9",X"16",X"E6",X"07",X"FD",X"77",X"04",X"E5",X"CD",
		X"C3",X"17",X"CD",X"B5",X"17",X"E1",X"11",X"20",X"00",X"19",X"10",X"FD",X"36",X"2E",X"23",X"0D",
		X"20",X"FA",X"C3",X"A9",X"16",X"FD",X"6E",X"07",X"FD",X"66",X"08",X"7E",X"23",X"66",X"6F",X"4E",
		X"23",X"46",X"C9",X"FD",X"75",X"05",X"FD",X"74",X"06",X"FD",X"5E",X"07",X"FD",X"56",X"08",X"87",
		X"4F",X"06",X"00",X"EB",X"09",X"7E",X"23",X"66",X"6F",X"EB",X"CD",X"D0",X"14",X"C9",X"FD",X"21",
		X"EB",X"17",X"CD",X"F6",X"18",X"FD",X"7E",X"09",X"D7",X"18",X"F3",X"81",X"F8",X"40",X"FF",X"0A",
		X"F2",X"48",X"82",X"20",X"07",X"08",X"7E",X"A7",X"C8",X"23",X"4E",X"23",X"46",X"23",X"5E",X"23",
		X"56",X"23",X"EB",X"CD",X"88",X"02",X"EB",X"18",X"ED",X"3B",X"00",X"AB",X"0A",X"09",X"1A",X"86",
		X"18",X"4F",X"ED",X"57",X"F3",X"F5",X"AF",X"08",X"FD",X"E5",X"DD",X"21",X"6D",X"40",X"21",X"6F",
		X"40",X"DD",X"7E",X"00",X"A7",X"C4",X"3D",X"18",X"DD",X"23",X"21",X"97",X"40",X"DD",X"7E",X"00",
		X"A7",X"C4",X"3D",X"18",X"FD",X"E1",X"08",X"47",X"F1",X"78",X"E0",X"FB",X"C9",X"06",X"08",X"0F",
		X"38",X"08",X"23",X"23",X"23",X"23",X"23",X"10",X"F6",X"C9",X"32",X"6C",X"40",X"79",X"BE",X"28",
		X"05",X"3A",X"6C",X"40",X"18",X"EC",X"C5",X"3E",X"FE",X"0F",X"10",X"FD",X"DD",X"A6",X"00",X"DD",
		X"77",X"00",X"08",X"F6",X"FF",X"F5",X"23",X"5E",X"23",X"56",X"23",X"4E",X"23",X"46",X"23",X"C5",
		X"FD",X"E1",X"EB",X"D5",X"DD",X"E5",X"11",X"7B",X"18",X"D5",X"E9",X"DD",X"E1",X"E1",X"F1",X"08",
		X"C1",X"3A",X"6C",X"40",X"18",X"C1",X"84",X"FF",X"06",X"1A",X"1A",X"DB",X"4B",X"07",X"B2",X"2E",
		X"01",X"09",X"08",X"00",X"2E",X"FD",X"E5",X"E1",X"01",X"08",X"00",X"09",X"FD",X"5E",X"02",X"FD",
		X"56",X"03",X"01",X"06",X"00",X"ED",X"B0",X"EB",X"FD",X"6E",X"04",X"FD",X"66",X"05",X"FD",X"CB",
		X"00",X"56",X"28",X"03",X"2B",X"18",X"04",X"01",X"DF",X"FF",X"09",X"E5",X"EB",X"01",X"03",X"00",
		X"ED",X"B0",X"01",X"1D",X"00",X"EB",X"09",X"EB",X"01",X"03",X"00",X"ED",X"B0",X"EB",X"FD",X"6E",
		X"02",X"FD",X"66",X"03",X"01",X"00",X"08",X"09",X"EB",X"01",X"06",X"00",X"ED",X"B0",X"EB",X"E1",
		X"01",X"00",X"08",X"09",X"EB",X"01",X"03",X"00",X"ED",X"B0",X"EB",X"01",X"1D",X"00",X"09",X"EB",
		X"01",X"03",X"00",X"ED",X"B0",X"C9",X"FD",X"6E",X"01",X"FD",X"66",X"02",X"FD",X"7E",X"03",X"77",
		X"FD",X"6E",X"07",X"FD",X"66",X"08",X"0E",X"01",X"46",X"FD",X"6E",X"05",X"FD",X"66",X"06",X"FD",
		X"CB",X"00",X"46",X"20",X"05",X"CD",X"86",X"02",X"18",X"0A",X"11",X"00",X"08",X"19",X"FD",X"7E",
		X"0A",X"CD",X"88",X"02",X"FD",X"7E",X"04",X"F7",X"FD",X"5E",X"07",X"FD",X"56",X"08",X"FD",X"6E",
		X"05",X"FD",X"66",X"06",X"E5",X"D5",X"CD",X"87",X"0B",X"E1",X"0E",X"01",X"46",X"E1",X"11",X"00",
		X"08",X"19",X"FD",X"7E",X"0A",X"0F",X"0F",X"0F",X"0F",X"CD",X"88",X"02",X"FD",X"7E",X"04",X"F7",
		X"FD",X"6E",X"01",X"FD",X"66",X"02",X"35",X"20",X"A7",X"00",X"00",X"00",X"00",X"FD",X"7E",X"09",
		X"CF",X"C9",X"E1",X"FD",X"E5",X"D1",X"DD",X"21",X"6D",X"40",X"FD",X"21",X"6F",X"40",X"C3",X"28",
		X"1A",X"AF",X"21",X"6C",X"40",X"77",X"23",X"77",X"23",X"77",X"C9",X"AF",X"21",X"19",X"40",X"77",
		X"23",X"77",X"23",X"77",X"C9",X"01",X"35",X"1A",X"31",X"01",X"34",X"00",X"1A",X"33",X"00",X"01",
		X"32",X"1A",X"31",X"01",X"30",X"00",X"02",X"01",X"57",X"56",X"06",X"F8",X"21",X"03",X"40",X"16",
		X"00",X"3A",X"EE",X"40",X"4F",X"3A",X"ED",X"40",X"E6",X"02",X"28",X"03",X"AF",X"18",X"03",X"CD",
		X"02",X"1B",X"B1",X"4F",X"3A",X"EF",X"40",X"2F",X"A1",X"4F",X"7E",X"5F",X"CB",X"19",X"30",X"01",
		X"3D",X"CB",X"19",X"30",X"01",X"3C",X"77",X"A0",X"08",X"7B",X"A0",X"5F",X"08",X"BB",X"28",X"08",
		X"38",X"04",X"CB",X"CA",X"18",X"02",X"CB",X"C2",X"23",X"7E",X"5F",X"CB",X"19",X"30",X"01",X"3C",
		X"CB",X"19",X"30",X"01",X"3D",X"77",X"A0",X"08",X"7B",X"A0",X"5F",X"08",X"BB",X"28",X"08",X"38",
		X"04",X"CB",X"D2",X"18",X"02",X"CB",X"DA",X"7A",X"E6",X"0F",X"28",X"0C",X"32",X"D4",X"40",X"21",
		X"ED",X"40",X"CB",X"4E",X"C0",X"CD",X"F1",X"10",X"C9",X"98",X"08",X"01",X"1A",X"1A",X"A2",X"48",
		X"21",X"AA",X"1F",X"11",X"02",X"40",X"01",X"03",X"00",X"ED",X"B0",X"C9",X"E1",X"FD",X"E5",X"D1",
		X"DD",X"21",X"1A",X"40",X"FD",X"21",X"1C",X"40",X"01",X"28",X"00",X"08",X"ED",X"57",X"F3",X"F5",
		X"D5",X"D9",X"01",X"00",X"08",X"DD",X"7E",X"00",X"FE",X"FF",X"20",X"10",X"DD",X"23",X"D9",X"FD",
		X"09",X"D9",X"DD",X"7E",X"00",X"FE",X"FF",X"20",X"03",X"C3",X"00",X"00",X"CB",X"3F",X"30",X"06",
		X"0C",X"10",X"F9",X"C3",X"00",X"00",X"F6",X"80",X"05",X"28",X"04",X"CB",X"3F",X"10",X"FC",X"DD",
		X"B6",X"00",X"DD",X"77",X"00",X"79",X"87",X"87",X"81",X"4F",X"FD",X"09",X"D9",X"08",X"FD",X"77",
		X"00",X"FD",X"75",X"01",X"FD",X"74",X"02",X"FD",X"73",X"03",X"FD",X"72",X"04",X"FD",X"E1",X"F1",
		X"E0",X"FB",X"C9",X"80",X"00",X"10",X"04",X"40",X"00",X"20",X"04",X"20",X"00",X"08",X"01",X"20",
		X"00",X"08",X"01",X"80",X"00",X"40",X"04",X"20",X"00",X"18",X"04",X"08",X"00",X"08",X"08",X"80",
		X"00",X"10",X"01",X"10",X"00",X"10",X"01",X"80",X"00",X"18",X"09",X"80",X"00",X"08",X"00",X"28",
		X"08",X"20",X"00",X"08",X"08",X"20",X"00",X"08",X"08",X"60",X"00",X"08",X"01",X"30",X"00",X"18",
		X"08",X"80",X"00",X"10",X"0A",X"40",X"00",X"08",X"08",X"C0",X"00",X"10",X"01",X"40",X"00",X"04",
		X"08",X"20",X"00",X"04",X"08",X"60",X"00",X"28",X"01",X"40",X"00",X"20",X"01",X"40",X"00",X"08",
		X"01",X"80",X"00",X"20",X"04",X"60",X"00",X"08",X"02",X"40",X"00",X"08",X"04",X"80",X"00",X"18",
		X"06",X"40",X"00",X"10",X"04",X"C0",X"00",X"20",X"05",X"80",X"00",X"08",X"01",X"40",X"00",X"20",
		X"04",X"00",X"DB",X"00",X"E6",X"02",X"20",X"07",X"3A",X"C1",X"40",X"CB",X"47",X"20",X"04",X"DB",
		X"01",X"2F",X"C9",X"DB",X"01",X"2F",X"0F",X"0F",X"0F",X"0F",X"C9",X"3E",X"08",X"F7",X"FD",X"CB",
		X"00",X"F6",X"01",X"06",X"10",X"E7",X"FD",X"7E",X"00",X"E6",X"0C",X"32",X"EF",X"40",X"07",X"CB",
		X"67",X"28",X"02",X"3E",X"04",X"32",X"EE",X"40",X"C3",X"2E",X"25",X"59",X"1B",X"00",X"5D",X"1B",
		X"00",X"61",X"1B",X"00",X"65",X"1B",X"00",X"69",X"1B",X"00",X"6D",X"1B",X"00",X"71",X"1B",X"00",
		X"21",X"F6",X"70",X"73",X"23",X"77",X"21",X"AB",X"72",X"81",X"03",X"FA",X"00",X"81",X"03",X"FA",
		X"00",X"81",X"03",X"FB",X"00",X"81",X"03",X"FC",X"00",X"81",X"03",X"FD",X"00",X"81",X"03",X"FE",
		X"00",X"81",X"03",X"FE",X"00",X"DF",X"70",X"4E",X"79",X"12",X"2E",X"F0",X"36",X"07",X"23",X"36",
		X"00",X"DD",X"21",X"B0",X"40",X"DD",X"7E",X"19",X"07",X"07",X"07",X"07",X"E6",X"F0",X"5F",X"DD",
		X"7E",X"18",X"E6",X"0F",X"B3",X"5F",X"DD",X"7E",X"1A",X"E6",X"4B",X"F6",X"48",X"57",X"3A",X"05",
		X"41",X"A7",X"28",X"02",X"13",X"FE",X"1B",X"C9",X"21",X"A2",X"50",X"18",X"03",X"21",X"A2",X"48",
		X"0E",X"1A",X"11",X"20",X"00",X"E5",X"DD",X"7E",X"00",X"A7",X"C4",X"BD",X"1F",X"DD",X"23",X"E1",
		X"19",X"0D",X"20",X"F1",X"C9",X"06",X"01",X"70",X"71",X"72",X"73",X"74",X"75",X"06",X"01",X"76",
		X"77",X"78",X"79",X"74",X"75",X"04",X"01",X"7A",X"7B",X"7C",X"7D",X"03",X"02",X"2E",X"81",X"82",
		X"83",X"2E",X"84",X"F5",X"E5",X"21",X"00",X"40",X"78",X"06",X"00",X"09",X"47",X"ED",X"57",X"EA",
		X"FA",X"1B",X"78",X"B6",X"77",X"ED",X"79",X"E1",X"F1",X"C9",X"78",X"F3",X"B6",X"77",X"ED",X"79",
		X"E1",X"FB",X"F1",X"C9",X"F5",X"E5",X"21",X"00",X"40",X"78",X"06",X"00",X"09",X"47",X"ED",X"57",
		X"EA",X"1C",X"1C",X"78",X"2F",X"A6",X"77",X"ED",X"79",X"E1",X"F1",X"C9",X"78",X"2F",X"F3",X"A6",
		X"77",X"ED",X"79",X"E1",X"FB",X"F1",X"C9",X"0F",X"2E",X"2E",X"12",X"17",X"1C",X"0E",X"1B",X"1D",
		X"2E",X"0C",X"18",X"12",X"17",X"2E",X"2E",X"ED",X"5B",X"E9",X"40",X"3A",X"33",X"43",X"6F",X"3A",
		X"6F",X"43",X"67",X"CD",X"D8",X"43",X"ED",X"53",X"0B",X"41",X"DD",X"21",X"98",X"41",X"0E",X"02",
		X"DD",X"7E",X"00",X"CB",X"7F",X"C4",X"DB",X"1C",X"EB",X"11",X"0C",X"00",X"DD",X"19",X"EB",X"0D",
		X"20",X"EE",X"21",X"89",X"41",X"CB",X"7E",X"28",X"1A",X"7E",X"4F",X"E6",X"0C",X"28",X"0A",X"CB",
		X"61",X"28",X"15",X"79",X"EE",X"1C",X"4F",X"18",X"0F",X"CB",X"61",X"28",X"0B",X"79",X"EE",X"13",
		X"4F",X"18",X"05",X"0E",X"80",X"18",X"01",X"4E",X"3A",X"C1",X"40",X"E6",X"01",X"20",X"05",X"21",
		X"0D",X"41",X"18",X"03",X"21",X"1F",X"41",X"06",X"06",X"CB",X"7E",X"28",X"08",X"23",X"23",X"23",
		X"10",X"F7",X"CD",X"00",X"00",X"71",X"23",X"73",X"23",X"72",X"C9",X"23",X"70",X"2C",X"73",X"CD",
		X"9B",X"5D",X"21",X"62",X"74",X"7E",X"2C",X"46",X"D3",X"F2",X"2C",X"7E",X"D6",X"31",X"C2",X"C7",
		X"5D",X"2C",X"36",X"20",X"C3",X"CA",X"5D",X"2C",X"36",X"00",X"2E",X"62",X"4E",X"2C",X"46",X"48",
		X"79",X"E6",X"0F",X"2E",X"65",X"B6",X"D3",X"F1",X"DB",X"F0",X"2C",X"DD",X"7E",X"00",X"E6",X"0C",
		X"20",X"0A",X"CD",X"FF",X"1C",X"C0",X"CD",X"84",X"1E",X"C0",X"18",X"08",X"CD",X"62",X"1E",X"C0",
		X"CD",X"6D",X"1E",X"C0",X"0E",X"80",X"DD",X"5E",X"0A",X"DD",X"56",X"0B",X"E1",X"18",X"89",X"D5",
		X"DD",X"6E",X"05",X"DD",X"66",X"06",X"29",X"29",X"29",X"EB",X"29",X"29",X"29",X"7A",X"D1",X"94",
		X"C9",X"3E",X"01",X"D7",X"CD",X"71",X"19",X"CD",X"7B",X"19",X"CD",X"6F",X"1D",X"AF",X"21",X"ED",
		X"40",X"36",X"00",X"CD",X"37",X"1C",X"3E",X"F7",X"32",X"02",X"40",X"CD",X"80",X"02",X"3E",X"02",
		X"F7",X"AF",X"32",X"04",X"41",X"3E",X"FF",X"D3",X"05",X"01",X"06",X"04",X"EF",X"CD",X"63",X"05",
		X"CD",X"5F",X"23",X"CD",X"E8",X"00",X"CD",X"CE",X"09",X"CD",X"E1",X"1F",X"3E",X"07",X"32",X"02",
		X"40",X"3E",X"02",X"F7",X"CD",X"10",X"1A",X"FD",X"21",X"39",X"41",X"FD",X"CB",X"00",X"7E",X"C4",
		X"75",X"1D",X"FD",X"21",X"59",X"41",X"FD",X"CB",X"00",X"7E",X"C4",X"75",X"1D",X"18",X"68",X"01",
		X"06",X"08",X"E7",X"EF",X"C9",X"FD",X"CB",X"00",X"B6",X"AF",X"32",X"EE",X"40",X"32",X"EF",X"40",
		X"CD",X"95",X"18",X"CD",X"25",X"24",X"FD",X"6E",X"02",X"FD",X"66",X"03",X"01",X"00",X"08",X"09",
		X"01",X"06",X"01",X"FD",X"7E",X"01",X"CD",X"88",X"02",X"FD",X"CB",X"00",X"56",X"28",X"05",X"11",
		X"1C",X"21",X"18",X"03",X"11",X"2C",X"21",X"FD",X"6E",X"02",X"FD",X"66",X"03",X"CD",X"D0",X"14",
		X"01",X"06",X"40",X"E7",X"3E",X"04",X"F7",X"FD",X"CB",X"00",X"56",X"28",X"05",X"11",X"24",X"21",
		X"18",X"03",X"11",X"34",X"21",X"FD",X"6E",X"02",X"FD",X"66",X"03",X"CD",X"D0",X"14",X"01",X"06",
		X"40",X"EF",X"3E",X"04",X"F7",X"18",X"C2",X"3E",X"60",X"F7",X"CD",X"7B",X"19",X"01",X"06",X"78",
		X"EF",X"CD",X"10",X"1A",X"3A",X"C0",X"40",X"CB",X"4F",X"20",X"14",X"3A",X"F0",X"40",X"A7",X"C2",
		X"5C",X"1E",X"FD",X"21",X"4D",X"0B",X"CD",X"B2",X"0A",X"3E",X"04",X"D7",X"C3",X"80",X"07",X"3A",
		X"C1",X"40",X"E6",X"01",X"20",X"2B",X"3A",X"F0",X"40",X"A7",X"28",X"12",X"3A",X"F1",X"40",X"A7",
		X"CA",X"5C",X"1E",X"3E",X"01",X"32",X"C1",X"40",X"CD",X"BE",X"15",X"C3",X"5C",X"1E",X"FD",X"21",
		X"C9",X"0A",X"CD",X"B2",X"0A",X"3E",X"04",X"D7",X"3A",X"F1",X"40",X"A7",X"20",X"E5",X"C3",X"80",
		X"07",X"3A",X"F1",X"40",X"A7",X"28",X"12",X"3A",X"F0",X"40",X"A7",X"CA",X"5C",X"1E",X"3E",X"00",
		X"32",X"C1",X"40",X"CD",X"AD",X"15",X"C3",X"5C",X"1E",X"FD",X"21",X"D4",X"0A",X"CD",X"B2",X"0A",
		X"3E",X"04",X"D7",X"3A",X"F0",X"40",X"A7",X"20",X"E5",X"C3",X"80",X"07",X"00",X"00",X"00",X"C3",
		X"64",X"13",X"DD",X"7E",X"05",X"E6",X"1F",X"6F",X"7B",X"E6",X"1F",X"95",X"C9",X"DD",X"6E",X"05",
		X"DD",X"66",X"06",X"29",X"29",X"29",X"D5",X"EB",X"29",X"29",X"29",X"7A",X"D1",X"94",X"C8",X"3C",
		X"C8",X"3D",X"3D",X"C9",X"DD",X"7E",X"05",X"E6",X"1F",X"6F",X"7B",X"E6",X"1F",X"95",X"C8",X"3C",
		X"C8",X"3D",X"3D",X"C9",X"3A",X"C1",X"40",X"CB",X"47",X"20",X"05",X"3A",X"CF",X"40",X"18",X"03",
		X"3A",X"D0",X"40",X"0E",X"08",X"FE",X"11",X"38",X"0A",X"FE",X"21",X"38",X"02",X"00",X"0D",X"0D",
		X"0D",X"0D",X"00",X"3A",X"CD",X"40",X"3C",X"32",X"CD",X"40",X"B9",X"38",X"3C",X"AF",X"32",X"CD",
		X"40",X"21",X"02",X"40",X"3A",X"CE",X"40",X"A7",X"20",X"17",X"7E",X"E6",X"07",X"FE",X"06",X"20",
		X"09",X"3E",X"FF",X"32",X"CE",X"40",X"06",X"06",X"18",X"1A",X"3C",X"47",X"18",X"16",X"00",X"00",
		X"00",X"7E",X"E6",X"07",X"20",X"09",X"3E",X"00",X"32",X"CE",X"40",X"06",X"00",X"18",X"05",X"3D",
		X"47",X"00",X"00",X"00",X"7E",X"E6",X"F8",X"B0",X"77",X"C9",X"21",X"17",X"1F",X"DB",X"00",X"E6",
		X"0C",X"0F",X"0F",X"4F",X"06",X"00",X"09",X"7E",X"32",X"F0",X"40",X"08",X"3A",X"C0",X"40",X"CB",
		X"4F",X"C8",X"08",X"32",X"F1",X"40",X"C9",X"02",X"03",X"04",X"05",X"3E",X"1E",X"32",X"09",X"41",
		X"3E",X"F0",X"F7",X"3A",X"09",X"41",X"3D",X"32",X"09",X"41",X"20",X"F4",X"3A",X"39",X"41",X"E6",
		X"80",X"20",X"09",X"CD",X"E3",X"06",X"3E",X"32",X"F7",X"CD",X"03",X"22",X"3E",X"20",X"F7",X"18",
		X"EB",X"11",X"2E",X"2E",X"0C",X"1B",X"0A",X"23",X"22",X"2E",X"0B",X"0A",X"15",X"15",X"18",X"18",
		X"17",X"2E",X"2E",X"21",X"12",X"40",X"01",X"07",X"04",X"E7",X"01",X"08",X"00",X"E7",X"E7",X"DB",
		X"03",X"2F",X"E6",X"40",X"BE",X"77",X"C0",X"23",X"BE",X"C8",X"77",X"A7",X"01",X"0D",X"01",X"28",
		X"02",X"E7",X"C9",X"EF",X"DB",X"00",X"E6",X"E0",X"C8",X"07",X"07",X"07",X"4F",X"06",X"00",X"21",
		X"A0",X"1F",X"09",X"7E",X"21",X"14",X"40",X"11",X"15",X"40",X"86",X"FE",X"0C",X"30",X"02",X"77",
		X"C9",X"D6",X"0C",X"08",X"1A",X"FE",X"09",X"28",X"05",X"D2",X"00",X"00",X"3C",X"12",X"08",X"18",
		X"EA",X"03",X"04",X"06",X"0C",X"18",X"24",X"30",X"00",X"00",X"F7",X"80",X"00",X"FF",X"00",X"14",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DD",X"7E",X"00",X"A7",X"C8",X"47",X"DD",X"23",
		X"DD",X"7E",X"00",X"FE",X"2E",X"28",X"08",X"77",X"23",X"10",X"FC",X"DD",X"23",X"18",X"E9",X"23",
		X"10",X"FD",X"DD",X"23",X"18",X"E2",X"04",X"10",X"18",X"0A",X"15",X"05",X"1C",X"1D",X"0A",X"1B",
		X"1D",X"3A",X"C1",X"40",X"CB",X"47",X"20",X"05",X"3A",X"F0",X"40",X"18",X"03",X"3A",X"F1",X"40",
		X"A7",X"C8",X"F5",X"CD",X"00",X"20",X"11",X"96",X"19",X"CD",X"D0",X"14",X"F1",X"3D",X"18",X"F0",
		X"07",X"4F",X"06",X"00",X"FD",X"2A",X"FE",X"40",X"FD",X"6E",X"10",X"FD",X"66",X"11",X"09",X"5E",
		X"23",X"56",X"EB",X"C9",X"21",X"03",X"00",X"4D",X"79",X"86",X"4F",X"23",X"7C",X"FE",X"28",X"20",
		X"F7",X"79",X"FE",X"6A",X"28",X"0A",X"2E",X"60",X"26",X"0A",X"2B",X"2B",X"D1",X"E3",X"E5",X"D5",
		X"CA",X"64",X"13",X"43",X"20",X"46",X"20",X"4A",X"20",X"4E",X"20",X"52",X"20",X"56",X"20",X"5A",
		X"20",X"5E",X"20",X"01",X"01",X"39",X"02",X"01",X"55",X"54",X"02",X"01",X"53",X"52",X"02",X"01",
		X"51",X"50",X"02",X"01",X"4F",X"4E",X"02",X"01",X"4D",X"4C",X"02",X"01",X"4B",X"4A",X"02",X"01",
		X"2E",X"69",X"21",X"10",X"40",X"DB",X"03",X"2F",X"E6",X"04",X"BE",X"77",X"C0",X"23",X"BE",X"C8",
		X"77",X"A7",X"C0",X"3A",X"15",X"40",X"FE",X"09",X"C8",X"D2",X"00",X"00",X"3C",X"32",X"15",X"40",
		X"C9",X"C9",X"08",X"5C",X"2E",X"19",X"1E",X"1C",X"11",X"2E",X"5C",X"0F",X"01",X"19",X"15",X"0A",
		X"22",X"0E",X"1B",X"2E",X"2E",X"0B",X"1E",X"1D",X"1D",X"18",X"17",X"07",X"0C",X"1B",X"0E",X"0D",
		X"12",X"1D",X"2C",X"DB",X"03",X"E6",X"02",X"C0",X"21",X"7E",X"41",X"7E",X"A7",X"C8",X"EB",X"21",
		X"BF",X"14",X"CD",X"B8",X"21",X"ED",X"B0",X"21",X"BE",X"49",X"01",X"01",X"0A",X"CD",X"86",X"02",
		X"C3",X"70",X"26",X"3E",X"20",X"F7",X"FD",X"CB",X"00",X"B6",X"AF",X"32",X"EF",X"40",X"32",X"EE",
		X"40",X"01",X"06",X"10",X"EF",X"C9",X"11",X"20",X"20",X"7C",X"D6",X"20",X"ED",X"44",X"92",X"67",
		X"E6",X"07",X"47",X"7D",X"ED",X"44",X"93",X"6F",X"E6",X"07",X"4F",X"7C",X"1F",X"1F",X"1F",X"1F",
		X"CB",X"1D",X"1F",X"CB",X"1D",X"1F",X"CB",X"1D",X"E6",X"4B",X"F6",X"48",X"67",X"C9",X"81",X"10",
		X"F0",X"00",X"CD",X"34",X"14",X"CB",X"27",X"4F",X"06",X"00",X"21",X"3E",X"28",X"09",X"5E",X"23",
		X"56",X"ED",X"53",X"FE",X"40",X"FD",X"21",X"00",X"00",X"FD",X"19",X"C9",X"06",X"01",X"9A",X"9B",
		X"9C",X"9D",X"9E",X"9F",X"06",X"01",X"A0",X"A1",X"A2",X"A3",X"A4",X"A5",X"06",X"01",X"A6",X"A7",
		X"A8",X"A9",X"AA",X"AB",X"06",X"01",X"AC",X"AD",X"AE",X"AF",X"B0",X"B1",X"DB",X"03",X"E6",X"08",
		X"C0",X"3A",X"BF",X"40",X"A7",X"C0",X"CD",X"C8",X"15",X"3E",X"FF",X"32",X"07",X"41",X"21",X"2A",
		X"49",X"01",X"0A",X"12",X"CD",X"86",X"02",X"21",X"CF",X"49",X"11",X"85",X"21",X"CD",X"87",X"0B",
		X"FD",X"21",X"7A",X"21",X"CD",X"F6",X"18",X"FD",X"7E",X"09",X"D7",X"CD",X"80",X"02",X"AF",X"32",
		X"07",X"41",X"3E",X"FF",X"32",X"BF",X"40",X"C3",X"DF",X"0A",X"81",X"F8",X"40",X"18",X"04",X"CF",
		X"49",X"85",X"21",X"12",X"F0",X"07",X"1D",X"2E",X"12",X"2E",X"15",X"2E",X"1D",X"08",X"AF",X"08",
		X"D6",X"0A",X"38",X"06",X"08",X"C6",X"10",X"27",X"18",X"F5",X"C6",X"0A",X"4F",X"08",X"81",X"27",
		X"C9",X"81",X"18",X"EB",X"12",X"ED",X"08",X"EB",X"18",X"E7",X"18",X"E7",X"12",X"E7",X"08",X"E4",
		X"12",X"E7",X"08",X"E8",X"18",X"E7",X"00",X"B3",X"4E",X"0C",X"06",X"00",X"C9",X"42",X"4F",X"21",
		X"C7",X"36",X"09",X"7E",X"07",X"C9",X"4E",X"3A",X"ED",X"40",X"E6",X"02",X"C0",X"3A",X"39",X"41",
		X"E6",X"80",X"C0",X"06",X"F8",X"2A",X"03",X"40",X"7D",X"A0",X"6F",X"3A",X"F6",X"40",X"A0",X"BD",
		X"20",X"0A",X"7C",X"A0",X"67",X"3A",X"F7",X"40",X"A0",X"BC",X"28",X"0A",X"22",X"F6",X"40",X"2A",
		X"F2",X"40",X"22",X"F4",X"40",X"C9",X"2A",X"F4",X"40",X"01",X"01",X"00",X"A7",X"ED",X"42",X"22",
		X"F4",X"40",X"C0",X"3A",X"03",X"40",X"E6",X"F8",X"47",X"21",X"3F",X"41",X"D6",X"14",X"77",X"23",
		X"78",X"C6",X"14",X"77",X"2A",X"03",X"40",X"CD",X"D6",X"20",X"ED",X"5B",X"D5",X"40",X"1A",X"E6",
		X"0C",X"20",X"09",X"3A",X"04",X"40",X"FE",X"80",X"38",X"06",X"18",X"21",X"E6",X"04",X"28",X"1D",
		X"3E",X"88",X"32",X"39",X"41",X"01",X"C0",X"00",X"09",X"E5",X"01",X"C0",X"4B",X"37",X"ED",X"42",
		X"38",X"28",X"E1",X"26",X"4B",X"7D",X"E6",X"DF",X"F6",X"C0",X"6F",X"18",X"1E",X"3E",X"84",X"32",
		X"39",X"41",X"01",X"80",X"FF",X"09",X"E5",X"01",X"A0",X"48",X"37",X"ED",X"42",X"30",X"0B",X"E1",
		X"26",X"48",X"7D",X"E6",X"BF",X"F6",X"A0",X"6F",X"18",X"01",X"E1",X"22",X"3B",X"41",X"3A",X"39",
		X"41",X"E6",X"04",X"28",X"05",X"01",X"21",X"00",X"18",X"03",X"01",X"E1",X"FF",X"09",X"22",X"3D",
		X"41",X"FD",X"21",X"39",X"41",X"FD",X"36",X"01",X"F4",X"C3",X"CB",X"02",X"DB",X"00",X"E6",X"10",
		X"20",X"05",X"21",X"AA",X"22",X"18",X"03",X"21",X"AE",X"22",X"E5",X"11",X"31",X"41",X"01",X"04",
		X"00",X"ED",X"B0",X"E1",X"01",X"04",X"00",X"ED",X"B0",X"C9",X"00",X"00",X"50",X"00",X"00",X"00",
		X"00",X"01",X"CD",X"08",X"16",X"3E",X"FF",X"32",X"06",X"41",X"3A",X"C1",X"40",X"CB",X"47",X"20",
		X"08",X"21",X"31",X"41",X"11",X"C4",X"40",X"18",X"06",X"21",X"35",X"41",X"11",X"C7",X"40",X"CB",
		X"7E",X"C0",X"23",X"23",X"23",X"CD",X"52",X"07",X"D8",X"3A",X"C1",X"40",X"CB",X"47",X"20",X"17",
		X"21",X"31",X"41",X"CB",X"FE",X"FD",X"E5",X"FD",X"21",X"FE",X"20",X"CD",X"0A",X"0F",X"FD",X"E1",
		X"21",X"F0",X"40",X"34",X"C3",X"E1",X"1F",X"21",X"35",X"41",X"CB",X"FE",X"FD",X"E5",X"FD",X"21",
		X"FE",X"20",X"CD",X"0A",X"0F",X"FD",X"E1",X"21",X"F1",X"40",X"34",X"C3",X"E1",X"1F",X"06",X"29",
		X"2E",X"18",X"1B",X"2E",X"29",X"0F",X"02",X"19",X"15",X"0A",X"22",X"0E",X"1B",X"2E",X"2E",X"0B",
		X"1E",X"1D",X"1D",X"18",X"17",X"15",X"5C",X"2E",X"01",X"19",X"15",X"0A",X"22",X"0E",X"1B",X"2E",
		X"10",X"0A",X"16",X"0E",X"2E",X"18",X"1F",X"0E",X"1B",X"2E",X"5C",X"15",X"5C",X"2E",X"02",X"19",
		X"15",X"0A",X"22",X"0E",X"1B",X"2E",X"10",X"0A",X"16",X"0E",X"2E",X"18",X"1F",X"0E",X"1B",X"2E",
		X"5C",X"0D",X"5C",X"2E",X"10",X"0A",X"16",X"0E",X"2E",X"18",X"1F",X"0E",X"1B",X"2E",X"5C",X"FD",
		X"2A",X"FE",X"40",X"FD",X"5E",X"00",X"FD",X"56",X"01",X"DD",X"21",X"00",X"00",X"DD",X"19",X"CD",
		X"AD",X"1B",X"FD",X"6E",X"02",X"FD",X"66",X"03",X"CD",X"F6",X"17",X"11",X"D6",X"1F",X"FD",X"6E",
		X"04",X"FD",X"66",X"05",X"CD",X"87",X"0B",X"11",X"DB",X"1F",X"FD",X"6E",X"06",X"FD",X"66",X"07",
		X"CD",X"87",X"0B",X"C9",X"3A",X"08",X"41",X"A7",X"28",X"05",X"3D",X"32",X"08",X"41",X"C9",X"3E",
		X"C0",X"32",X"08",X"41",X"01",X"01",X"00",X"E7",X"C9",X"3E",X"80",X"F7",X"CD",X"D0",X"23",X"21",
		X"70",X"07",X"FD",X"21",X"98",X"41",X"CD",X"5E",X"16",X"FD",X"7E",X"09",X"D7",X"3E",X"02",X"F7",
		X"21",X"7C",X"07",X"FD",X"21",X"98",X"41",X"CD",X"56",X"16",X"FD",X"7E",X"09",X"D7",X"18",X"DF",
		X"3E",X"80",X"F7",X"21",X"78",X"08",X"FD",X"21",X"A4",X"41",X"CD",X"5E",X"16",X"FD",X"7E",X"09",
		X"D7",X"3E",X"30",X"F7",X"21",X"C3",X"08",X"FD",X"21",X"A4",X"41",X"CD",X"56",X"16",X"FD",X"7E",
		X"09",X"D7",X"3E",X"20",X"F7",X"18",X"DC",X"12",X"17",X"0A",X"16",X"0E",X"2E",X"2E",X"1B",X"0E",
		X"10",X"12",X"1C",X"1D",X"1B",X"0A",X"1D",X"12",X"18",X"17",X"10",X"17",X"0A",X"16",X"0E",X"2E",
		X"2E",X"29",X"29",X"29",X"29",X"29",X"29",X"29",X"29",X"29",X"29",X"09",X"2D",X"2E",X"2E",X"2E",
		X"B4",X"B5",X"2E",X"B6",X"B7",X"FD",X"E5",X"E1",X"01",X"08",X"00",X"09",X"EB",X"FD",X"6E",X"02",
		X"FD",X"66",X"03",X"01",X"06",X"00",X"ED",X"B0",X"FD",X"6E",X"04",X"FD",X"66",X"05",X"FD",X"CB",
		X"00",X"56",X"28",X"03",X"2B",X"18",X"04",X"01",X"DF",X"FF",X"09",X"E5",X"01",X"03",X"00",X"ED",
		X"B0",X"01",X"1D",X"00",X"09",X"01",X"03",X"00",X"ED",X"B0",X"FD",X"6E",X"02",X"FD",X"66",X"03",
		X"01",X"00",X"08",X"09",X"01",X"06",X"00",X"ED",X"B0",X"E1",X"01",X"00",X"08",X"09",X"01",X"03",
		X"00",X"ED",X"B0",X"01",X"1D",X"00",X"09",X"01",X"03",X"00",X"ED",X"B0",X"C9",X"21",X"FD",X"49",
		X"11",X"18",X"40",X"18",X"15",X"3A",X"C1",X"40",X"CB",X"47",X"20",X"08",X"21",X"BD",X"48",X"11",
		X"C4",X"40",X"18",X"06",X"21",X"1D",X"4B",X"11",X"C7",X"40",X"06",X"06",X"0E",X"00",X"CB",X"40",
		X"20",X"09",X"1A",X"0F",X"0F",X"0F",X"0F",X"CD",X"B9",X"24",X"05",X"05",X"20",X"02",X"CB",X"C1",
		X"04",X"1A",X"CD",X"B9",X"24",X"1B",X"10",X"EA",X"C9",X"E6",X"0F",X"28",X"0A",X"CB",X"C1",X"77",
		X"C5",X"01",X"20",X"00",X"09",X"C1",X"C9",X"CB",X"41",X"20",X"F4",X"3E",X"2E",X"18",X"F0",X"3E",
		X"15",X"32",X"7A",X"41",X"3E",X"F0",X"F7",X"3A",X"7A",X"41",X"3D",X"32",X"7A",X"41",X"20",X"F4",
		X"FD",X"21",X"A8",X"26",X"CD",X"F6",X"18",X"FD",X"7E",X"09",X"D7",X"CD",X"7B",X"19",X"3E",X"0A",
		X"CF",X"C9",X"F2",X"48",X"32",X"49",X"72",X"49",X"B2",X"49",X"F2",X"49",X"32",X"4A",X"72",X"4A",
		X"B2",X"4A",X"F2",X"4A",X"32",X"4B",X"72",X"4B",X"F0",X"48",X"30",X"49",X"70",X"49",X"B0",X"49",
		X"F0",X"49",X"30",X"4A",X"70",X"4A",X"B0",X"4A",X"F0",X"4A",X"30",X"4B",X"70",X"4B",X"EE",X"48",
		X"2E",X"49",X"6E",X"49",X"AE",X"49",X"EE",X"49",X"2E",X"4A",X"6E",X"4A",X"CE",X"4A",X"3E",X"01",
		X"F7",X"21",X"CD",X"40",X"7E",X"FE",X"06",X"30",X"02",X"36",X"06",X"23",X"FD",X"7E",X"00",X"E6",
		X"04",X"28",X"19",X"CB",X"7E",X"28",X"0B",X"3A",X"02",X"40",X"E6",X"07",X"FE",X"04",X"30",X"02",
		X"36",X"00",X"FD",X"7E",X"00",X"E6",X"60",X"EE",X"40",X"28",X"D3",X"C9",X"CB",X"7E",X"20",X"F2",
		X"3A",X"02",X"40",X"E6",X"07",X"FE",X"03",X"38",X"E9",X"36",X"FF",X"18",X"E5",X"DD",X"21",X"B5",
		X"40",X"DD",X"7E",X"16",X"E6",X"08",X"C8",X"3A",X"CC",X"40",X"FE",X"02",X"D2",X"18",X"15",X"3C",
		X"32",X"CC",X"40",X"C9",X"FD",X"2A",X"FE",X"40",X"FD",X"6E",X"12",X"FD",X"66",X"13",X"E5",X"11",
		X"16",X"26",X"CD",X"87",X"0B",X"E1",X"11",X"00",X"08",X"19",X"01",X"01",X"05",X"3E",X"F4",X"CD",
		X"88",X"02",X"21",X"D9",X"26",X"11",X"01",X"41",X"01",X"03",X"00",X"ED",X"B0",X"3E",X"80",X"F7",
		X"FD",X"6E",X"12",X"FD",X"66",X"13",X"01",X"01",X"05",X"CD",X"86",X"02",X"3E",X"10",X"F7",X"FD",
		X"6E",X"12",X"FD",X"66",X"13",X"11",X"02",X"41",X"06",X"04",X"CD",X"9C",X"24",X"3E",X"05",X"32",
		X"00",X"41",X"3E",X"F0",X"F7",X"3A",X"00",X"41",X"3D",X"32",X"00",X"41",X"20",X"F4",X"FD",X"6E",
		X"12",X"FD",X"66",X"13",X"01",X"01",X"05",X"CD",X"86",X"02",X"3E",X"10",X"F7",X"21",X"CA",X"26",
		X"11",X"01",X"41",X"CD",X"3E",X"16",X"FD",X"6E",X"12",X"FD",X"66",X"13",X"11",X"02",X"41",X"06",
		X"04",X"CD",X"9C",X"24",X"3E",X"10",X"F7",X"21",X"03",X"41",X"11",X"15",X"26",X"CD",X"52",X"07",
		X"20",X"CC",X"C9",X"00",X"00",X"00",X"05",X"0B",X"18",X"17",X"1E",X"1C",X"39",X"55",X"39",X"6F",
		X"2E",X"54",X"54",X"52",X"6F",X"6E",X"55",X"53",X"52",X"50",X"6E",X"6D",X"53",X"51",X"50",X"4E",
		X"6D",X"6C",X"51",X"4F",X"4E",X"4C",X"6C",X"6B",X"4F",X"4D",X"4C",X"4A",X"6B",X"6A",X"4D",X"4B",
		X"4B",X"2E",X"6A",X"69",X"4A",X"69",X"69",X"39",X"69",X"39",X"69",X"39",X"3E",X"05",X"32",X"F8",
		X"40",X"21",X"BE",X"49",X"01",X"01",X"0A",X"CD",X"86",X"02",X"3E",X"05",X"F7",X"CD",X"70",X"26",
		X"3E",X"05",X"F7",X"3A",X"F8",X"40",X"3D",X"32",X"F8",X"40",X"20",X"E5",X"3E",X"0B",X"CF",X"C9",
		X"21",X"7E",X"41",X"7E",X"FE",X"02",X"38",X"29",X"FE",X"04",X"38",X"20",X"FE",X"06",X"38",X"17",
		X"FE",X"08",X"38",X"0E",X"FE",X"0A",X"38",X"05",X"11",X"BE",X"49",X"18",X"17",X"11",X"DE",X"49",
		X"18",X"12",X"11",X"FE",X"49",X"18",X"0D",X"11",X"1E",X"4A",X"18",X"08",X"11",X"3E",X"4A",X"18",
		X"03",X"11",X"5E",X"4A",X"EB",X"C3",X"87",X"0B",X"80",X"79",X"41",X"05",X"1E",X"46",X"49",X"0A",
		X"24",X"0C",X"00",X"21",X"03",X"49",X"11",X"8D",X"18",X"CD",X"87",X"0B",X"21",X"03",X"51",X"01",
		X"01",X"07",X"3E",X"F6",X"C3",X"88",X"02",X"10",X"00",X"00",X"20",X"00",X"00",X"00",X"01",X"00",
		X"00",X"02",X"00",X"00",X"03",X"00",X"00",X"05",X"00",X"00",X"10",X"00",X"C9",X"2A",X"B8",X"73",
		X"23",X"22",X"B8",X"73",X"21",X"3E",X"05",X"32",X"F8",X"40",X"FD",X"2A",X"FE",X"40",X"FD",X"6E",
		X"04",X"FD",X"66",X"05",X"01",X"01",X"04",X"CD",X"86",X"02",X"3E",X"08",X"F7",X"FD",X"2A",X"FE",
		X"40",X"FD",X"6E",X"04",X"FD",X"66",X"05",X"11",X"D6",X"1F",X"CD",X"87",X"0B",X"3E",X"08",X"F7",
		X"3A",X"F8",X"40",X"3D",X"32",X"F8",X"40",X"20",X"D1",X"21",X"01",X"41",X"CD",X"0E",X"16",X"CD",
		X"85",X"24",X"3E",X"04",X"F7",X"FD",X"6E",X"12",X"FD",X"66",X"13",X"01",X"01",X"05",X"CD",X"86",
		X"02",X"3E",X"40",X"F7",X"3E",X"03",X"CF",X"C9",X"21",X"0E",X"06",X"18",X"08",X"21",X"16",X"06",
		X"18",X"03",X"21",X"1E",X"06",X"11",X"59",X"41",X"FD",X"E5",X"D5",X"FD",X"E1",X"01",X"08",X"00",
		X"ED",X"B0",X"CD",X"C8",X"02",X"FD",X"E1",X"C9",X"81",X"08",X"DD",X"08",X"E1",X"08",X"E4",X"08",
		X"E6",X"08",X"E1",X"08",X"E4",X"08",X"E6",X"08",X"E9",X"08",X"E4",X"08",X"E6",X"08",X"E9",X"08",
		X"EB",X"08",X"E6",X"08",X"E9",X"08",X"EB",X"08",X"ED",X"08",X"E9",X"08",X"EB",X"08",X"ED",X"28",
		X"EE",X"00",X"3A",X"73",X"21",X"C0",X"73",X"4E",X"2E",X"3C",X"71",X"23",X"36",X"00",X"01",X"C2",
		X"73",X"11",X"E2",X"70",X"CD",X"1F",X"3A",X"21",X"E2",X"70",X"4E",X"06",X"00",X"CD",X"ED",X"42",
		X"21",X"F4",X"70",X"4E",X"2C",X"46",X"2A",X"C2",X"73",X"09",X"22",X"F4",X"70",X"3E",X"FF",X"21",
		X"F4",X"70",X"96",X"2C",X"4F",X"3E",X"00",X"9E",X"9F",X"2A",X"F4",X"70",X"2B",X"22",X"EE",X"70",
		X"EB",X"21",X"44",X"71",X"19",X"4F",X"7E",X"D6",X"0A",X"C6",X"FF",X"9F",X"A1",X"0F",X"D2",X"F4",
		X"48",X"21",X"38",X"73",X"36",X"01",X"23",X"36",X"00",X"01",X"44",X"71",X"2C",X"71",X"23",X"70",
		X"2C",X"36",X"FF",X"23",X"36",X"00",X"01",X"C2",X"73",X"11",X"E2",X"70",X"CD",X"1F",X"3A",X"0E",
		X"0F",X"CD",X"15",X"42",X"21",X"EE",X"70",X"4E",X"2C",X"46",X"24",X"2E",X"44",X"09",X"7E",X"D6",
		X"A8",X"04",X"02",X"70",X"08",X"04",X"38",X"0A",X"09",X"60",X"07",X"08",X"78",X"0D",X"0C",X"40",
		X"04",X"0E",X"40",X"07",X"06",X"58",X"0A",X"0B",X"78",X"0D",X"0C",X"88",X"05",X"04",X"30",X"04",
		X"05",X"A8",X"09",X"08",X"38",X"0C",X"0B",X"70",X"0F",X"10",X"78",X"11",X"0F",X"80",X"10",X"06",
		X"21",X"C8",X"73",X"77",X"D6",X"30",X"9F",X"2E",X"CB",X"4F",X"7E",X"2E",X"C8",X"96",X"9F",X"C5",
		X"60",X"28",X"60",X"28",X"5D",X"2A",X"60",X"28",X"5D",X"2A",X"A5",X"2C",X"5D",X"2A",X"A5",X"2C",
		X"60",X"28",X"60",X"28",X"5D",X"2A",X"60",X"28",X"5D",X"2A",X"A5",X"2C",X"5D",X"2A",X"A5",X"2C",
		X"86",X"28",X"B8",X"29",X"D6",X"48",X"27",X"4B",X"DC",X"29",X"DF",X"29",X"E2",X"29",X"ED",X"29",
		X"4F",X"2A",X"BB",X"48",X"02",X"11",X"01",X"02",X"68",X"01",X"04",X"46",X"01",X"0A",X"71",X"01",
		X"0C",X"77",X"01",X"00",X"00",X"00",X"14",X"39",X"01",X"33",X"00",X"04",X"39",X"08",X"2E",X"02",
		X"39",X"03",X"2E",X"03",X"39",X"00",X"03",X"39",X"0E",X"2E",X"03",X"39",X"00",X"03",X"39",X"0F",
		X"2E",X"02",X"39",X"00",X"02",X"39",X"10",X"2E",X"02",X"39",X"00",X"02",X"39",X"0B",X"2E",X"02",
		X"39",X"03",X"2E",X"02",X"39",X"01",X"32",X"05",X"2E",X"01",X"BA",X"00",X"02",X"39",X"0C",X"2E",
		X"01",X"39",X"05",X"2E",X"01",X"39",X"00",X"02",X"39",X"04",X"2E",X"02",X"39",X"07",X"2E",X"01",
		X"39",X"00",X"01",X"39",X"05",X"2E",X"02",X"39",X"07",X"2E",X"02",X"39",X"08",X"2E",X"01",X"39",
		X"00",X"01",X"39",X"06",X"2E",X"01",X"39",X"07",X"2E",X"03",X"39",X"07",X"2E",X"01",X"39",X"00",
		X"01",X"39",X"06",X"2E",X"02",X"39",X"06",X"2E",X"02",X"39",X"07",X"2E",X"02",X"39",X"00",X"01",
		X"39",X"06",X"2E",X"02",X"39",X"05",X"2E",X"02",X"39",X"06",X"2E",X"04",X"39",X"00",X"01",X"39",
		X"06",X"2E",X"02",X"39",X"04",X"2E",X"02",X"39",X"07",X"2E",X"04",X"39",X"00",X"01",X"39",X"06",
		X"2E",X"02",X"39",X"0C",X"2E",X"05",X"39",X"00",X"07",X"2E",X"02",X"39",X"0D",X"2E",X"04",X"39",
		X"00",X"07",X"2E",X"02",X"39",X"06",X"2E",X"02",X"39",X"07",X"2E",X"02",X"39",X"00",X"06",X"2E",
		X"04",X"39",X"05",X"2E",X"02",X"39",X"07",X"2E",X"02",X"39",X"00",X"06",X"2E",X"04",X"39",X"05",
		X"2E",X"03",X"39",X"06",X"2E",X"02",X"39",X"00",X"05",X"2E",X"04",X"39",X"06",X"2E",X"04",X"39",
		X"05",X"2E",X"02",X"39",X"00",X"05",X"2E",X"01",X"33",X"02",X"39",X"06",X"2E",X"01",X"39",X"04",
		X"2E",X"01",X"39",X"05",X"2E",X"01",X"39",X"00",X"06",X"2E",X"01",X"39",X"12",X"2E",X"01",X"39",
		X"00",X"06",X"2E",X"01",X"39",X"12",X"2E",X"01",X"39",X"00",X"06",X"2E",X"02",X"39",X"10",X"2E",
		X"02",X"39",X"00",X"06",X"2E",X"04",X"39",X"0E",X"2E",X"02",X"39",X"00",X"06",X"2E",X"05",X"39",
		X"04",X"2E",X"02",X"39",X"06",X"2E",X"03",X"39",X"00",X"05",X"2E",X"01",X"33",X"14",X"39",X"00",
		X"37",X"1E",X"03",X"CD",X"10",X"49",X"2F",X"0F",X"F2",X"05",X"02",X"AF",X"50",X"F2",X"07",X"04",
		X"EF",X"50",X"F2",X"04",X"03",X"6F",X"51",X"F6",X"06",X"06",X"B6",X"50",X"F5",X"04",X"06",X"10",
		X"52",X"F6",X"05",X"07",X"02",X"53",X"F5",X"01",X"07",X"07",X"53",X"00",X"64",X"28",X"D0",X"64",
		X"D0",X"40",X"0A",X"00",X"38",X"E8",X"A8",X"A8",X"60",X"38",X"70",X"70",X"00",X"80",X"00",X"38",
		X"02",X"08",X"01",X"E0",X"01",X"A8",X"05",X"04",X"00",X"A0",X"03",X"40",X"01",X"E0",X"02",X"A8",
		X"04",X"01",X"00",X"E0",X"03",X"A8",X"80",X"E0",X"03",X"70",X"09",X"08",X"00",X"A0",X"03",X"40",
		X"05",X"A0",X"02",X"70",X"08",X"01",X"00",X"38",X"83",X"08",X"05",X"A0",X"01",X"60",X"06",X"01",
		X"00",X"38",X"07",X"08",X"01",X"58",X"05",X"00",X"06",X"04",X"00",X"A0",X"86",X"40",X"06",X"58",
		X"08",X"00",X"07",X"01",X"09",X"A0",X"09",X"40",X"05",X"68",X"04",X"60",X"07",X"01",X"0C",X"E0",
		X"09",X"A8",X"89",X"68",X"03",X"38",X"0A",X"40",X"00",X"E0",X"0A",X"A8",X"07",X"30",X"09",X"00",
		X"0A",X"C2",X"4B",X"A2",X"4B",X"C4",X"4B",X"A4",X"4B",X"82",X"4B",X"84",X"4B",X"83",X"2A",X"C9",
		X"2B",X"C9",X"48",X"C7",X"48",X"ED",X"2B",X"F0",X"2B",X"F3",X"2B",X"03",X"2C",X"97",X"2C",X"CA",
		X"48",X"03",X"16",X"01",X"05",X"50",X"01",X"07",X"46",X"01",X"0B",X"6B",X"01",X"0D",X"7D",X"01",
		X"0F",X"83",X"01",X"05",X"2E",X"01",X"33",X"01",X"39",X"01",X"35",X"05",X"31",X"01",X"34",X"0C",
		X"39",X"00",X"06",X"2E",X"01",X"39",X"08",X"2E",X"02",X"39",X"05",X"2E",X"04",X"39",X"00",X"06",
		X"2E",X"01",X"39",X"11",X"2E",X"02",X"39",X"00",X"06",X"2E",X"01",X"39",X"11",X"2E",X"02",X"39",
		X"00",X"06",X"2E",X"01",X"39",X"11",X"2E",X"02",X"39",X"00",X"06",X"2E",X"01",X"39",X"01",X"33",
		X"07",X"2E",X"03",X"39",X"07",X"2E",X"01",X"39",X"00",X"05",X"2E",X"01",X"33",X"01",X"39",X"01",
		X"32",X"05",X"31",X"01",X"30",X"06",X"39",X"05",X"2E",X"01",X"39",X"00",X"05",X"2E",X"0E",X"39",
		X"06",X"2E",X"01",X"39",X"00",X"06",X"2E",X"03",X"39",X"04",X"2E",X"05",X"39",X"07",X"2E",X"01",
		X"39",X"00",X"06",X"2E",X"02",X"39",X"06",X"2E",X"03",X"39",X"07",X"2E",X"02",X"39",X"00",X"0E",
		X"2E",X"03",X"39",X"05",X"2E",X"04",X"39",X"00",X"01",X"39",X"0D",X"2E",X"02",X"39",X"05",X"2E",
		X"05",X"39",X"00",X"02",X"39",X"0B",X"2E",X"03",X"39",X"05",X"2E",X"05",X"39",X"00",X"02",X"39",
		X"06",X"2E",X"01",X"39",X"05",X"2E",X"01",X"39",X"05",X"2E",X"06",X"39",X"00",X"01",X"39",X"06",
		X"2E",X"03",X"39",X"04",X"2E",X"01",X"39",X"05",X"2E",X"06",X"39",X"00",X"01",X"39",X"05",X"2E",
		X"03",X"39",X"05",X"2E",X"01",X"39",X"06",X"2E",X"05",X"39",X"00",X"01",X"39",X"06",X"2E",X"01",
		X"39",X"06",X"2E",X"02",X"39",X"06",X"2E",X"04",X"39",X"00",X"01",X"39",X"06",X"2E",X"02",X"39",
		X"05",X"2E",X"03",X"39",X"07",X"2E",X"02",X"39",X"00",X"01",X"39",X"07",X"2E",X"02",X"39",X"05",
		X"2E",X"03",X"39",X"07",X"2E",X"01",X"39",X"00",X"01",X"39",X"07",X"2E",X"03",X"39",X"05",X"2E",
		X"03",X"39",X"06",X"2E",X"01",X"39",X"00",X"02",X"39",X"06",X"2E",X"02",X"39",X"08",X"2E",X"01",
		X"39",X"06",X"2E",X"01",X"39",X"00",X"02",X"39",X"16",X"2E",X"02",X"39",X"00",X"04",X"39",X"14",
		X"2E",X"02",X"39",X"00",X"04",X"39",X"0A",X"2E",X"01",X"39",X"08",X"2E",X"03",X"39",X"00",X"05",
		X"39",X"02",X"2E",X"02",X"39",X"04",X"2E",X"03",X"39",X"06",X"2E",X"04",X"39",X"00",X"1A",X"39",
		X"00",X"CD",X"AC",X"44",X"21",X"D7",X"70",X"77",X"C3",X"F2",X"05",X"07",X"A2",X"50",X"F5",X"01",
		X"07",X"A7",X"50",X"F6",X"07",X"07",X"A9",X"50",X"F2",X"02",X"07",X"B0",X"50",X"F5",X"07",X"02",
		X"4A",X"52",X"F5",X"03",X"07",X"12",X"53",X"F5",X"04",X"06",X"28",X"53",X"00",X"24",X"80",X"C8",
		X"24",X"D0",X"C0",X"0F",X"E8",X"A8",X"68",X"A8",X"88",X"68",X"00",X"38",X"60",X"08",X"50",X"A8",
		X"78",X"68",X"60",X"80",X"00",X"E0",X"01",X"A8",X"02",X"E0",X"01",X"A8",X"0F",X"08",X"00",X"A0",
		X"01",X"68",X"03",X"E0",X"02",X"A8",X"8C",X"08",X"00",X"60",X"02",X"08",X"03",X"E0",X"03",X"A8",
		X"8F",X"01",X"09",X"38",X"0E",X"08",X"04",X"A0",X"03",X"88",X"05",X"01",X"00",X"38",X"0E",X"08",
		X"05",X"80",X"04",X"68",X"06",X"01",X"09",X"38",X"08",X"08",X"06",X"60",X"05",X"40",X"07",X"04",
		X"00",X"38",X"08",X"08",X"07",X"38",X"06",X"00",X"07",X"04",X"00",X"60",X"09",X"40",X"92",X"60",
		X"0E",X"00",X"08",X"04",X"00",X"A0",X"95",X"68",X"08",X"60",X"98",X"00",X"09",X"02",X"00",X"E0",
		X"0A",X"A8",X"09",X"50",X"0B",X"00",X"0A",X"02",X"0C",X"E0",X"0B",X"A8",X"09",X"60",X"0F",X"58",
		X"0A",X"01",X"00",X"A0",X"0F",X"78",X"0D",X"A0",X"02",X"68",X"09",X"08",X"09",X"70",X"0C",X"68",
		X"0E",X"A0",X"02",X"68",X"09",X"08",X"00",X"60",X"0D",X"40",X"9B",X"A0",X"03",X"68",X"08",X"40",
		X"00",X"E0",X"0F",X"A8",X"0C",X"A0",X"01",X"68",X"0B",X"A2",X"48",X"C2",X"48",X"A4",X"48",X"C4",
		X"48",X"E2",X"48",X"E4",X"48",X"CB",X"2C",X"63",X"2E",X"53",X"4B",X"3B",X"4B",X"91",X"2E",X"94",
		X"2E",X"97",X"2E",X"AA",X"2E",X"5C",X"2F",X"52",X"4B",X"06",X"1B",X"01",X"0E",X"6E",X"01",X"10",
		X"46",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1A",X"39",X"00",X"03",X"39",
		X"02",X"2E",X"01",X"39",X"02",X"2E",X"08",X"39",X"03",X"2E",X"02",X"39",X"03",X"2E",X"02",X"39",
		X"00",X"02",X"39",X"08",X"2E",X"06",X"39",X"04",X"2E",X"01",X"39",X"04",X"2E",X"01",X"39",X"00",
		X"01",X"39",X"0A",X"2E",X"04",X"39",X"0A",X"2E",X"01",X"39",X"00",X"01",X"39",X"0A",X"2E",X"02",
		X"39",X"0C",X"2E",X"01",X"39",X"00",X"01",X"39",X"06",X"2E",X"01",X"39",X"04",X"2E",X"01",X"39",
		X"0C",X"2E",X"01",X"39",X"00",X"01",X"39",X"05",X"2E",X"03",X"39",X"08",X"2E",X"03",X"39",X"05",
		X"2E",X"01",X"39",X"00",X"02",X"39",X"05",X"2E",X"03",X"39",X"07",X"2E",X"02",X"39",X"06",X"2E",
		X"01",X"39",X"00",X"03",X"39",X"04",X"2E",X"03",X"39",X"06",X"2E",X"03",X"39",X"06",X"2E",X"01",
		X"39",X"00",X"02",X"39",X"05",X"2E",X"03",X"39",X"06",X"2E",X"02",X"39",X"06",X"2E",X"02",X"39",
		X"00",X"02",X"39",X"05",X"2E",X"03",X"39",X"03",X"2E",X"05",X"39",X"04",X"2E",X"04",X"39",X"00",
		X"01",X"39",X"05",X"2E",X"05",X"39",X"03",X"2E",X"04",X"39",X"04",X"2E",X"04",X"39",X"00",X"01",
		X"39",X"05",X"2E",X"06",X"39",X"03",X"2E",X"03",X"39",X"05",X"2E",X"03",X"39",X"00",X"01",X"39",
		X"04",X"2E",X"08",X"39",X"03",X"2E",X"02",X"39",X"06",X"2E",X"02",X"39",X"00",X"01",X"39",X"04",
		X"2E",X"02",X"39",X"03",X"2E",X"02",X"39",X"05",X"2E",X"02",X"39",X"06",X"2E",X"01",X"39",X"00",
		X"01",X"39",X"03",X"2E",X"03",X"39",X"0A",X"2E",X"02",X"39",X"06",X"2E",X"01",X"39",X"00",X"01",
		X"39",X"04",X"2E",X"01",X"39",X"0B",X"2E",X"03",X"39",X"05",X"2E",X"01",X"39",X"00",X"01",X"39",
		X"04",X"2E",X"01",X"39",X"0B",X"2E",X"03",X"39",X"05",X"2E",X"01",X"39",X"00",X"01",X"39",X"04",
		X"2E",X"01",X"39",X"04",X"2E",X"02",X"39",X"05",X"2E",X"03",X"39",X"05",X"2E",X"01",X"39",X"00",
		X"02",X"39",X"03",X"2E",X"01",X"39",X"04",X"2E",X"01",X"39",X"01",X"35",X"05",X"2E",X"01",X"34",
		X"01",X"39",X"01",X"35",X"05",X"2E",X"01",X"34",X"00",X"01",X"39",X"09",X"2E",X"01",X"39",X"01",
		X"33",X"05",X"2E",X"01",X"33",X"01",X"39",X"01",X"33",X"00",X"01",X"39",X"09",X"2E",X"01",X"39",
		X"01",X"33",X"06",X"2E",X"01",X"39",X"01",X"33",X"00",X"01",X"39",X"09",X"2E",X"01",X"39",X"01",
		X"33",X"06",X"2E",X"01",X"39",X"01",X"33",X"00",X"02",X"39",X"07",X"2E",X"02",X"39",X"01",X"33",
		X"06",X"2E",X"01",X"39",X"01",X"33",X"00",X"03",X"39",X"02",X"2E",X"01",X"39",X"02",X"2E",X"03",
		X"39",X"01",X"33",X"06",X"2E",X"01",X"39",X"01",X"33",X"00",X"0B",X"39",X"01",X"33",X"05",X"2E",
		X"01",X"33",X"01",X"39",X"01",X"33",X"05",X"2E",X"01",X"33",X"00",X"2A",X"0C",X"74",X"09",X"23",
		X"22",X"0C",X"74",X"F5",X"05",X"07",X"A7",X"50",X"F2",X"08",X"03",X"A2",X"51",X"F4",X"07",X"03",
		X"0C",X"52",X"F5",X"02",X"05",X"6C",X"52",X"F5",X"06",X"02",X"02",X"53",X"F6",X"07",X"07",X"0D",
		X"53",X"F5",X"01",X"07",X"15",X"53",X"F4",X"05",X"07",X"16",X"53",X"F5",X"01",X"07",X"1B",X"53",
		X"00",X"44",X"70",X"38",X"44",X"30",X"40",X"12",X"00",X"40",X"68",X"00",X"28",X"48",X"80",X"E8",
		X"A8",X"88",X"48",X"E8",X"B0",X"B0",X"88",X"88",X"78",X"48",X"80",X"00",X"40",X"02",X"08",X"01",
		X"48",X"12",X"00",X"01",X"04",X"00",X"68",X"03",X"48",X"01",X"48",X"11",X"00",X"02",X"04",X"00",
		X"98",X"9E",X"70",X"02",X"48",X"AD",X"00",X"03",X"04",X"00",X"E0",X"04",X"A0",X"03",X"28",X"05",
		X"00",X"04",X"02",X"00",X"E0",X"05",X"A0",X"03",X"48",X"06",X"30",X"04",X"02",X"00",X"E0",X"06",
		X"88",X"10",X"80",X"07",X"50",X"05",X"02",X"09",X"E0",X"07",X"88",X"0E",X"A8",X"A1",X"88",X"06",
		X"08",X"00",X"E0",X"08",X"A8",X"09",X"E0",X"08",X"B0",X"07",X"08",X"0C",X"A0",X"08",X"88",X"0A",
		X"E0",X"09",X"B0",X"07",X"08",X"00",X"80",X"09",X"48",X"0B",X"E0",X"0A",X"B0",X"0E",X"08",X"09",
		X"40",X"0A",X"38",X"0C",X"E0",X"0B",X"B0",X"0D",X"01",X"00",X"30",X"0B",X"08",X"0C",X"E0",X"0C",
		X"B0",X"0D",X"01",X"00",X"40",X"0E",X"08",X"0D",X"A8",X"A4",X"88",X"12",X"01",X"00",X"80",X"07",
		X"48",X"0D",X"A8",X"0A",X"88",X"A7",X"01",X"09",X"68",X"10",X"48",X"12",X"80",X"0E",X"78",X"11",
		X"08",X"0F",X"80",X"06",X"70",X"AA",X"80",X"0E",X"50",X"03",X"08",X"00",X"68",X"10",X"48",X"12",
		X"70",X"0F",X"50",X"02",X"40",X"00",X"40",X"AA",X"08",X"12",X"80",X"0D",X"50",X"01",X"D6",X"4B",
		X"D8",X"4B",X"B6",X"4B",X"B8",X"4B",X"96",X"4B",X"98",X"4B",X"2E",X"13",X"5E",X"CD",X"15",X"50",
		X"5F",X"21",X"13",X"74",X"4E",X"CD",X"E8",X"4E",X"21",X"13",X"74",X"34",X"C2",X"5A",X"50",X"C9",
		X"21",X"19",X"74",X"36",X"00",X"2D",X"36",X"00",X"0E",X"1B",X"0D",X"79",X"21",X"18",X"74",X"96",
		X"DA",X"B0",X"50",X"4E",X"CD",X"DB",X"4E",X"0F",X"D2",X"9F",X"50",X"21",X"19",X"74",X"34",X"21",
		X"19",X"74",X"7E",X"D6",X"02",X"DA",X"AB",X"50",X"3E",X"FF",X"C9",X"2D",X"34",X"C2",X"88",X"50",
		X"AF",X"C9",X"21",X"1A",X"74",X"36",X"00",X"0E",X"1B",X"0D",X"79",X"21",X"1A",X"74",X"96",X"DA",
		X"D3",X"50",X"4E",X"CD",X"DB",X"4E",X"0F",X"D2",X"CC",X"50",X"AF",X"C9",X"21",X"1A",X"74",X"34",
		X"C2",X"B7",X"50",X"3E",X"FF",X"C9",X"CD",X"12",X"50",X"CD",X"C3",X"46",X"CD",X"D2",X"43",X"21",
		X"07",X"74",X"77",X"2C",X"36",X"00",X"21",X"07",X"74",X"7E",X"D6",X"41",X"9F",X"2F",X"4F",X"3E",
		X"5A",X"96",X"9F",X"2F",X"A1",X"5F",X"7E",X"D6",X"30",X"9F",X"2F",X"D5",X"4F",X"3E",X"39",X"96",
		X"A8",X"04",X"02",X"70",X"08",X"04",X"38",X"0A",X"09",X"60",X"07",X"08",X"78",X"0D",X"0C",X"40",
		X"04",X"0E",X"40",X"07",X"06",X"58",X"0A",X"0B",X"78",X"0D",X"0C",X"88",X"05",X"04",X"30",X"04",
		X"05",X"A8",X"09",X"08",X"38",X"0C",X"0B",X"70",X"0F",X"10",X"78",X"11",X"0F",X"80",X"10",X"06",
		X"21",X"C8",X"73",X"77",X"D6",X"30",X"9F",X"2E",X"CB",X"4F",X"7E",X"2E",X"C8",X"96",X"9F",X"C5",
		X"60",X"28",X"60",X"28",X"5D",X"2A",X"60",X"28",X"5D",X"2A",X"A5",X"2C",X"5D",X"2A",X"A5",X"2C",
		X"60",X"28",X"60",X"28",X"5D",X"2A",X"60",X"28",X"5D",X"2A",X"A5",X"2C",X"5D",X"2A",X"A5",X"2C",
		X"86",X"28",X"B8",X"29",X"D6",X"48",X"27",X"4B",X"DC",X"29",X"DF",X"29",X"E2",X"29",X"ED",X"29",
		X"4F",X"2A",X"BB",X"48",X"02",X"11",X"01",X"02",X"68",X"01",X"04",X"46",X"01",X"0A",X"71",X"01",
		X"0C",X"77",X"01",X"00",X"00",X"00",X"14",X"39",X"01",X"33",X"00",X"04",X"39",X"08",X"2E",X"02",
		X"39",X"03",X"2E",X"03",X"39",X"00",X"03",X"39",X"0E",X"2E",X"03",X"39",X"00",X"03",X"39",X"0F",
		X"2E",X"02",X"39",X"00",X"02",X"39",X"10",X"2E",X"02",X"39",X"00",X"02",X"39",X"0B",X"2E",X"02",
		X"39",X"03",X"2E",X"02",X"39",X"01",X"32",X"05",X"2E",X"01",X"BA",X"00",X"02",X"39",X"0C",X"2E",
		X"01",X"39",X"05",X"2E",X"01",X"39",X"00",X"02",X"39",X"04",X"2E",X"02",X"39",X"07",X"2E",X"01",
		X"39",X"00",X"01",X"39",X"05",X"2E",X"02",X"39",X"07",X"2E",X"02",X"39",X"08",X"2E",X"01",X"39",
		X"00",X"01",X"39",X"06",X"2E",X"01",X"39",X"07",X"2E",X"03",X"39",X"07",X"2E",X"01",X"39",X"00",
		X"01",X"39",X"06",X"2E",X"02",X"39",X"06",X"2E",X"02",X"39",X"07",X"2E",X"02",X"39",X"00",X"01",
		X"39",X"06",X"2E",X"02",X"39",X"05",X"2E",X"02",X"39",X"06",X"2E",X"04",X"39",X"00",X"01",X"39",
		X"06",X"2E",X"02",X"39",X"04",X"2E",X"02",X"39",X"07",X"2E",X"04",X"39",X"00",X"01",X"39",X"06",
		X"2E",X"02",X"39",X"0C",X"2E",X"05",X"39",X"00",X"07",X"2E",X"02",X"39",X"0D",X"2E",X"04",X"39",
		X"00",X"07",X"2E",X"02",X"39",X"06",X"2E",X"02",X"39",X"07",X"2E",X"02",X"39",X"00",X"06",X"2E",
		X"04",X"39",X"05",X"2E",X"02",X"39",X"07",X"2E",X"02",X"39",X"00",X"06",X"2E",X"04",X"39",X"05",
		X"2E",X"03",X"39",X"06",X"2E",X"02",X"39",X"00",X"05",X"2E",X"04",X"39",X"06",X"2E",X"04",X"39",
		X"05",X"2E",X"02",X"39",X"00",X"05",X"2E",X"01",X"33",X"02",X"39",X"06",X"2E",X"01",X"39",X"04",
		X"2E",X"01",X"39",X"05",X"2E",X"01",X"39",X"00",X"06",X"2E",X"01",X"39",X"12",X"2E",X"01",X"39",
		X"00",X"06",X"2E",X"01",X"39",X"12",X"2E",X"01",X"39",X"00",X"06",X"2E",X"02",X"39",X"10",X"2E",
		X"02",X"39",X"00",X"06",X"2E",X"04",X"39",X"0E",X"2E",X"02",X"39",X"00",X"06",X"2E",X"05",X"39",
		X"04",X"2E",X"02",X"39",X"06",X"2E",X"03",X"39",X"00",X"05",X"2E",X"01",X"33",X"14",X"39",X"00",
		X"37",X"1E",X"03",X"CD",X"10",X"49",X"2F",X"0F",X"F2",X"05",X"02",X"AF",X"50",X"F2",X"07",X"04",
		X"EF",X"50",X"F2",X"04",X"03",X"6F",X"51",X"F6",X"06",X"06",X"B6",X"50",X"F5",X"04",X"06",X"10",
		X"52",X"F6",X"05",X"07",X"02",X"53",X"F5",X"01",X"07",X"07",X"53",X"00",X"64",X"28",X"D0",X"64",
		X"D0",X"40",X"0A",X"00",X"38",X"E8",X"A8",X"A8",X"60",X"38",X"70",X"70",X"00",X"80",X"00",X"38",
		X"02",X"08",X"01",X"E0",X"01",X"A8",X"05",X"04",X"00",X"A0",X"03",X"40",X"01",X"E0",X"02",X"A8",
		X"04",X"01",X"00",X"E0",X"03",X"A8",X"80",X"E0",X"03",X"70",X"09",X"08",X"00",X"A0",X"03",X"40",
		X"05",X"A0",X"02",X"70",X"08",X"01",X"00",X"38",X"83",X"08",X"05",X"A0",X"01",X"60",X"06",X"01",
		X"00",X"38",X"07",X"08",X"01",X"58",X"05",X"00",X"06",X"04",X"00",X"A0",X"86",X"40",X"06",X"58",
		X"08",X"00",X"07",X"01",X"09",X"A0",X"09",X"40",X"05",X"68",X"04",X"60",X"07",X"01",X"0C",X"E0",
		X"09",X"A8",X"89",X"68",X"03",X"38",X"0A",X"40",X"00",X"E0",X"0A",X"A8",X"07",X"30",X"09",X"00",
		X"0A",X"C2",X"4B",X"A2",X"4B",X"C4",X"4B",X"A4",X"4B",X"82",X"4B",X"84",X"4B",X"83",X"2A",X"C9",
		X"2B",X"C9",X"48",X"C7",X"48",X"ED",X"2B",X"F0",X"2B",X"F3",X"2B",X"03",X"2C",X"97",X"2C",X"CA",
		X"48",X"03",X"16",X"01",X"05",X"50",X"01",X"07",X"46",X"01",X"0B",X"6B",X"01",X"0D",X"7D",X"01",
		X"0F",X"83",X"01",X"05",X"2E",X"01",X"33",X"01",X"39",X"01",X"35",X"05",X"31",X"01",X"34",X"0C",
		X"39",X"00",X"06",X"2E",X"01",X"39",X"08",X"2E",X"02",X"39",X"05",X"2E",X"04",X"39",X"00",X"06",
		X"2E",X"01",X"39",X"11",X"2E",X"02",X"39",X"00",X"06",X"2E",X"01",X"39",X"11",X"2E",X"02",X"39",
		X"00",X"06",X"2E",X"01",X"39",X"11",X"2E",X"02",X"39",X"00",X"06",X"2E",X"01",X"39",X"01",X"33",
		X"07",X"2E",X"03",X"39",X"07",X"2E",X"01",X"39",X"00",X"05",X"2E",X"01",X"33",X"01",X"39",X"01",
		X"32",X"05",X"31",X"01",X"30",X"06",X"39",X"05",X"2E",X"01",X"39",X"00",X"05",X"2E",X"0E",X"39",
		X"06",X"2E",X"01",X"39",X"00",X"06",X"2E",X"03",X"39",X"04",X"2E",X"05",X"39",X"07",X"2E",X"01",
		X"39",X"00",X"06",X"2E",X"02",X"39",X"06",X"2E",X"03",X"39",X"07",X"2E",X"02",X"39",X"00",X"0E",
		X"2E",X"03",X"39",X"05",X"2E",X"04",X"39",X"00",X"01",X"39",X"0D",X"2E",X"02",X"39",X"05",X"2E",
		X"05",X"39",X"00",X"02",X"39",X"0B",X"2E",X"03",X"39",X"05",X"2E",X"05",X"39",X"00",X"02",X"39",
		X"06",X"2E",X"01",X"39",X"05",X"2E",X"01",X"39",X"05",X"2E",X"06",X"39",X"00",X"01",X"39",X"06",
		X"2E",X"03",X"39",X"04",X"2E",X"01",X"39",X"05",X"2E",X"06",X"39",X"00",X"01",X"39",X"05",X"2E",
		X"03",X"39",X"05",X"2E",X"01",X"39",X"06",X"2E",X"05",X"39",X"00",X"01",X"39",X"06",X"2E",X"01",
		X"39",X"06",X"2E",X"02",X"39",X"06",X"2E",X"04",X"39",X"00",X"01",X"39",X"06",X"2E",X"02",X"39",
		X"05",X"2E",X"03",X"39",X"07",X"2E",X"02",X"39",X"00",X"01",X"39",X"07",X"2E",X"02",X"39",X"05",
		X"2E",X"03",X"39",X"07",X"2E",X"01",X"39",X"00",X"01",X"39",X"07",X"2E",X"03",X"39",X"05",X"2E",
		X"03",X"39",X"06",X"2E",X"01",X"39",X"00",X"02",X"39",X"06",X"2E",X"02",X"39",X"08",X"2E",X"01",
		X"39",X"06",X"2E",X"01",X"39",X"00",X"02",X"39",X"16",X"2E",X"02",X"39",X"00",X"04",X"39",X"14",
		X"2E",X"02",X"39",X"00",X"04",X"39",X"0A",X"2E",X"01",X"39",X"08",X"2E",X"03",X"39",X"00",X"05",
		X"39",X"02",X"2E",X"02",X"39",X"04",X"2E",X"03",X"39",X"06",X"2E",X"04",X"39",X"00",X"1A",X"39",
		X"00",X"CD",X"AC",X"44",X"21",X"D7",X"70",X"77",X"C3",X"F2",X"05",X"07",X"A2",X"50",X"F5",X"01",
		X"07",X"A7",X"50",X"F6",X"07",X"07",X"A9",X"50",X"F2",X"02",X"07",X"B0",X"50",X"F5",X"07",X"02",
		X"4A",X"52",X"F5",X"03",X"07",X"12",X"53",X"F5",X"04",X"06",X"28",X"53",X"00",X"24",X"80",X"C8",
		X"24",X"D0",X"C0",X"0F",X"E8",X"A8",X"68",X"A8",X"88",X"68",X"00",X"38",X"60",X"08",X"50",X"A8",
		X"78",X"68",X"60",X"80",X"00",X"E0",X"01",X"A8",X"02",X"E0",X"01",X"A8",X"0F",X"08",X"00",X"A0",
		X"01",X"68",X"03",X"E0",X"02",X"A8",X"8C",X"08",X"00",X"60",X"02",X"08",X"03",X"E0",X"03",X"A8",
		X"8F",X"01",X"09",X"38",X"0E",X"08",X"04",X"A0",X"03",X"88",X"05",X"01",X"00",X"38",X"0E",X"08",
		X"05",X"80",X"04",X"68",X"06",X"01",X"09",X"38",X"08",X"08",X"06",X"60",X"05",X"40",X"07",X"04",
		X"00",X"38",X"08",X"08",X"07",X"38",X"06",X"00",X"07",X"04",X"00",X"60",X"09",X"40",X"92",X"60",
		X"0E",X"00",X"08",X"04",X"00",X"A0",X"95",X"68",X"08",X"60",X"98",X"00",X"09",X"02",X"00",X"E0",
		X"0A",X"A8",X"09",X"50",X"0B",X"00",X"0A",X"02",X"0C",X"E0",X"0B",X"A8",X"09",X"60",X"0F",X"58",
		X"0A",X"01",X"00",X"A0",X"0F",X"78",X"0D",X"A0",X"02",X"68",X"09",X"08",X"09",X"70",X"0C",X"68",
		X"0E",X"A0",X"02",X"68",X"09",X"08",X"00",X"60",X"0D",X"40",X"9B",X"A0",X"03",X"68",X"08",X"40",
		X"00",X"E0",X"0F",X"A8",X"0C",X"A0",X"01",X"68",X"0B",X"A2",X"48",X"C2",X"48",X"A4",X"48",X"C4",
		X"48",X"E2",X"48",X"E4",X"48",X"CB",X"2C",X"63",X"2E",X"53",X"4B",X"3B",X"4B",X"91",X"2E",X"94",
		X"2E",X"97",X"2E",X"AA",X"2E",X"5C",X"2F",X"52",X"4B",X"06",X"1B",X"01",X"0E",X"6E",X"01",X"10",
		X"46",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1A",X"39",X"00",X"03",X"39",
		X"02",X"2E",X"01",X"39",X"02",X"2E",X"08",X"39",X"03",X"2E",X"02",X"39",X"03",X"2E",X"02",X"39",
		X"00",X"02",X"39",X"08",X"2E",X"06",X"39",X"04",X"2E",X"01",X"39",X"04",X"2E",X"01",X"39",X"00",
		X"01",X"39",X"0A",X"2E",X"04",X"39",X"0A",X"2E",X"01",X"39",X"00",X"01",X"39",X"0A",X"2E",X"02",
		X"39",X"0C",X"2E",X"01",X"39",X"00",X"01",X"39",X"06",X"2E",X"01",X"39",X"04",X"2E",X"01",X"39",
		X"0C",X"2E",X"01",X"39",X"00",X"01",X"39",X"05",X"2E",X"03",X"39",X"08",X"2E",X"03",X"39",X"05",
		X"2E",X"01",X"39",X"00",X"02",X"39",X"05",X"2E",X"03",X"39",X"07",X"2E",X"02",X"39",X"06",X"2E",
		X"01",X"39",X"00",X"03",X"39",X"04",X"2E",X"03",X"39",X"06",X"2E",X"03",X"39",X"06",X"2E",X"01",
		X"39",X"00",X"02",X"39",X"05",X"2E",X"03",X"39",X"06",X"2E",X"02",X"39",X"06",X"2E",X"02",X"39",
		X"00",X"02",X"39",X"05",X"2E",X"03",X"39",X"03",X"2E",X"05",X"39",X"04",X"2E",X"04",X"39",X"00",
		X"01",X"39",X"05",X"2E",X"05",X"39",X"03",X"2E",X"04",X"39",X"04",X"2E",X"04",X"39",X"00",X"01",
		X"39",X"05",X"2E",X"06",X"39",X"03",X"2E",X"03",X"39",X"05",X"2E",X"03",X"39",X"00",X"01",X"39",
		X"04",X"2E",X"08",X"39",X"03",X"2E",X"02",X"39",X"06",X"2E",X"02",X"39",X"00",X"01",X"39",X"04",
		X"2E",X"02",X"39",X"03",X"2E",X"02",X"39",X"05",X"2E",X"02",X"39",X"06",X"2E",X"01",X"39",X"00",
		X"01",X"39",X"03",X"2E",X"03",X"39",X"0A",X"2E",X"02",X"39",X"06",X"2E",X"01",X"39",X"00",X"01",
		X"39",X"04",X"2E",X"01",X"39",X"0B",X"2E",X"03",X"39",X"05",X"2E",X"01",X"39",X"00",X"01",X"39",
		X"04",X"2E",X"01",X"39",X"0B",X"2E",X"03",X"39",X"05",X"2E",X"01",X"39",X"00",X"01",X"39",X"04",
		X"2E",X"01",X"39",X"04",X"2E",X"02",X"39",X"05",X"2E",X"03",X"39",X"05",X"2E",X"01",X"39",X"00",
		X"02",X"39",X"03",X"2E",X"01",X"39",X"04",X"2E",X"01",X"39",X"01",X"35",X"05",X"2E",X"01",X"34",
		X"01",X"39",X"01",X"35",X"05",X"2E",X"01",X"34",X"00",X"01",X"39",X"09",X"2E",X"01",X"39",X"01",
		X"33",X"05",X"2E",X"01",X"33",X"01",X"39",X"01",X"33",X"00",X"01",X"39",X"09",X"2E",X"01",X"39",
		X"01",X"33",X"06",X"2E",X"01",X"39",X"01",X"33",X"00",X"01",X"39",X"09",X"2E",X"01",X"39",X"01",
		X"33",X"06",X"2E",X"01",X"39",X"01",X"33",X"00",X"02",X"39",X"07",X"2E",X"02",X"39",X"01",X"33",
		X"06",X"2E",X"01",X"39",X"01",X"33",X"00",X"03",X"39",X"02",X"2E",X"01",X"39",X"02",X"2E",X"03",
		X"39",X"01",X"33",X"06",X"2E",X"01",X"39",X"01",X"33",X"00",X"0B",X"39",X"01",X"33",X"05",X"2E",
		X"01",X"33",X"01",X"39",X"01",X"33",X"05",X"2E",X"01",X"33",X"00",X"2A",X"0C",X"74",X"09",X"23",
		X"22",X"0C",X"74",X"F5",X"05",X"07",X"A7",X"50",X"F2",X"08",X"03",X"A2",X"51",X"F4",X"07",X"03",
		X"0C",X"52",X"F5",X"02",X"05",X"6C",X"52",X"F5",X"06",X"02",X"02",X"53",X"F6",X"07",X"07",X"0D",
		X"53",X"F5",X"01",X"07",X"15",X"53",X"F4",X"05",X"07",X"16",X"53",X"F5",X"01",X"07",X"1B",X"53",
		X"00",X"44",X"70",X"38",X"44",X"30",X"40",X"12",X"00",X"40",X"68",X"00",X"28",X"48",X"80",X"E8",
		X"A8",X"88",X"48",X"E8",X"B0",X"B0",X"88",X"88",X"78",X"48",X"80",X"00",X"40",X"02",X"08",X"01",
		X"48",X"12",X"00",X"01",X"04",X"00",X"68",X"03",X"48",X"01",X"48",X"11",X"00",X"02",X"04",X"00",
		X"98",X"9E",X"70",X"02",X"48",X"AD",X"00",X"03",X"04",X"00",X"E0",X"04",X"A0",X"03",X"28",X"05",
		X"00",X"04",X"02",X"00",X"E0",X"05",X"A0",X"03",X"48",X"06",X"30",X"04",X"02",X"00",X"E0",X"06",
		X"88",X"10",X"80",X"07",X"50",X"05",X"02",X"09",X"E0",X"07",X"88",X"0E",X"A8",X"A1",X"88",X"06",
		X"08",X"00",X"E0",X"08",X"A8",X"09",X"E0",X"08",X"B0",X"07",X"08",X"0C",X"A0",X"08",X"88",X"0A",
		X"E0",X"09",X"B0",X"07",X"08",X"00",X"80",X"09",X"48",X"0B",X"E0",X"0A",X"B0",X"0E",X"08",X"09",
		X"40",X"0A",X"38",X"0C",X"E0",X"0B",X"B0",X"0D",X"01",X"00",X"30",X"0B",X"08",X"0C",X"E0",X"0C",
		X"B0",X"0D",X"01",X"00",X"40",X"0E",X"08",X"0D",X"A8",X"A4",X"88",X"12",X"01",X"00",X"80",X"07",
		X"48",X"0D",X"A8",X"0A",X"88",X"A7",X"01",X"09",X"68",X"10",X"48",X"12",X"80",X"0E",X"78",X"11",
		X"08",X"0F",X"80",X"06",X"70",X"AA",X"80",X"0E",X"50",X"03",X"08",X"00",X"68",X"10",X"48",X"12",
		X"70",X"0F",X"50",X"02",X"40",X"00",X"40",X"AA",X"08",X"12",X"80",X"0D",X"50",X"01",X"D6",X"4B",
		X"D8",X"4B",X"B6",X"4B",X"B8",X"4B",X"96",X"4B",X"98",X"4B",X"2E",X"13",X"5E",X"CD",X"15",X"50",
		X"5F",X"21",X"13",X"74",X"4E",X"CD",X"E8",X"4E",X"21",X"13",X"74",X"34",X"C2",X"5A",X"50",X"C9",
		X"21",X"19",X"74",X"36",X"00",X"2D",X"36",X"00",X"0E",X"1B",X"0D",X"79",X"21",X"18",X"74",X"96",
		X"DA",X"B0",X"50",X"4E",X"CD",X"DB",X"4E",X"0F",X"D2",X"9F",X"50",X"21",X"19",X"74",X"34",X"21",
		X"19",X"74",X"7E",X"D6",X"02",X"DA",X"AB",X"50",X"3E",X"FF",X"C9",X"2D",X"34",X"C2",X"88",X"50",
		X"AF",X"C9",X"21",X"1A",X"74",X"36",X"00",X"0E",X"1B",X"0D",X"79",X"21",X"1A",X"74",X"96",X"DA",
		X"D3",X"50",X"4E",X"CD",X"DB",X"4E",X"0F",X"D2",X"CC",X"50",X"AF",X"C9",X"21",X"1A",X"74",X"34",
		X"C2",X"B7",X"50",X"3E",X"FF",X"C9",X"CD",X"12",X"50",X"CD",X"C3",X"46",X"CD",X"D2",X"43",X"21",
		X"07",X"74",X"77",X"2C",X"36",X"00",X"21",X"07",X"74",X"7E",X"D6",X"41",X"9F",X"2F",X"4F",X"3E",
		X"5A",X"96",X"9F",X"2F",X"A1",X"5F",X"7E",X"D6",X"30",X"9F",X"2F",X"D5",X"4F",X"3E",X"39",X"96",
		X"A8",X"04",X"02",X"70",X"08",X"04",X"38",X"0A",X"09",X"60",X"07",X"08",X"78",X"0D",X"0C",X"40",
		X"04",X"0E",X"40",X"07",X"06",X"58",X"0A",X"0B",X"78",X"0D",X"0C",X"88",X"05",X"04",X"30",X"04",
		X"05",X"A8",X"09",X"08",X"38",X"0C",X"0B",X"70",X"0F",X"10",X"78",X"11",X"0F",X"80",X"10",X"06",
		X"21",X"C8",X"73",X"77",X"D6",X"30",X"9F",X"2E",X"CB",X"4F",X"7E",X"2E",X"C8",X"96",X"9F",X"C5",
		X"60",X"28",X"60",X"28",X"5D",X"2A",X"60",X"28",X"5D",X"2A",X"A5",X"2C",X"5D",X"2A",X"A5",X"2C",
		X"60",X"28",X"60",X"28",X"5D",X"2A",X"60",X"28",X"5D",X"2A",X"A5",X"2C",X"5D",X"2A",X"A5",X"2C",
		X"86",X"28",X"B8",X"29",X"D6",X"48",X"27",X"4B",X"DC",X"29",X"DF",X"29",X"E2",X"29",X"ED",X"29",
		X"4F",X"2A",X"BB",X"48",X"02",X"11",X"01",X"02",X"68",X"01",X"04",X"46",X"01",X"0A",X"71",X"01",
		X"0C",X"77",X"01",X"00",X"00",X"00",X"14",X"39",X"01",X"33",X"00",X"04",X"39",X"08",X"2E",X"02",
		X"39",X"03",X"2E",X"03",X"39",X"00",X"03",X"39",X"0E",X"2E",X"03",X"39",X"00",X"03",X"39",X"0F",
		X"2E",X"02",X"39",X"00",X"02",X"39",X"10",X"2E",X"02",X"39",X"00",X"02",X"39",X"0B",X"2E",X"02",
		X"39",X"03",X"2E",X"02",X"39",X"01",X"32",X"05",X"2E",X"01",X"BA",X"00",X"02",X"39",X"0C",X"2E",
		X"01",X"39",X"05",X"2E",X"01",X"39",X"00",X"02",X"39",X"04",X"2E",X"02",X"39",X"07",X"2E",X"01",
		X"39",X"00",X"01",X"39",X"05",X"2E",X"02",X"39",X"07",X"2E",X"02",X"39",X"08",X"2E",X"01",X"39",
		X"00",X"01",X"39",X"06",X"2E",X"01",X"39",X"07",X"2E",X"03",X"39",X"07",X"2E",X"01",X"39",X"00",
		X"01",X"39",X"06",X"2E",X"02",X"39",X"06",X"2E",X"02",X"39",X"07",X"2E",X"02",X"39",X"00",X"01",
		X"39",X"06",X"2E",X"02",X"39",X"05",X"2E",X"02",X"39",X"06",X"2E",X"04",X"39",X"00",X"01",X"39",
		X"06",X"2E",X"02",X"39",X"04",X"2E",X"02",X"39",X"07",X"2E",X"04",X"39",X"00",X"01",X"39",X"06",
		X"2E",X"02",X"39",X"0C",X"2E",X"05",X"39",X"00",X"07",X"2E",X"02",X"39",X"0D",X"2E",X"04",X"39",
		X"00",X"07",X"2E",X"02",X"39",X"06",X"2E",X"02",X"39",X"07",X"2E",X"02",X"39",X"00",X"06",X"2E",
		X"04",X"39",X"05",X"2E",X"02",X"39",X"07",X"2E",X"02",X"39",X"00",X"06",X"2E",X"04",X"39",X"05",
		X"2E",X"03",X"39",X"06",X"2E",X"02",X"39",X"00",X"05",X"2E",X"04",X"39",X"06",X"2E",X"04",X"39",
		X"05",X"2E",X"02",X"39",X"00",X"05",X"2E",X"01",X"33",X"02",X"39",X"06",X"2E",X"01",X"39",X"04",
		X"2E",X"01",X"39",X"05",X"2E",X"01",X"39",X"00",X"06",X"2E",X"01",X"39",X"12",X"2E",X"01",X"39",
		X"00",X"06",X"2E",X"01",X"39",X"12",X"2E",X"01",X"39",X"00",X"06",X"2E",X"02",X"39",X"10",X"2E",
		X"02",X"39",X"00",X"06",X"2E",X"04",X"39",X"0E",X"2E",X"02",X"39",X"00",X"06",X"2E",X"05",X"39",
		X"04",X"2E",X"02",X"39",X"06",X"2E",X"03",X"39",X"00",X"05",X"2E",X"01",X"33",X"14",X"39",X"00",
		X"37",X"1E",X"03",X"CD",X"10",X"49",X"2F",X"0F",X"F2",X"05",X"02",X"AF",X"50",X"F2",X"07",X"04",
		X"EF",X"50",X"F2",X"04",X"03",X"6F",X"51",X"F6",X"06",X"06",X"B6",X"50",X"F5",X"04",X"06",X"10",
		X"52",X"F6",X"05",X"07",X"02",X"53",X"F5",X"01",X"07",X"07",X"53",X"00",X"64",X"28",X"D0",X"64",
		X"D0",X"40",X"0A",X"00",X"38",X"E8",X"A8",X"A8",X"60",X"38",X"70",X"70",X"00",X"80",X"00",X"38",
		X"02",X"08",X"01",X"E0",X"01",X"A8",X"05",X"04",X"00",X"A0",X"03",X"40",X"01",X"E0",X"02",X"A8",
		X"04",X"01",X"00",X"E0",X"03",X"A8",X"80",X"E0",X"03",X"70",X"09",X"08",X"00",X"A0",X"03",X"40",
		X"05",X"A0",X"02",X"70",X"08",X"01",X"00",X"38",X"83",X"08",X"05",X"A0",X"01",X"60",X"06",X"01",
		X"00",X"38",X"07",X"08",X"01",X"58",X"05",X"00",X"06",X"04",X"00",X"A0",X"86",X"40",X"06",X"58",
		X"08",X"00",X"07",X"01",X"09",X"A0",X"09",X"40",X"05",X"68",X"04",X"60",X"07",X"01",X"0C",X"E0",
		X"09",X"A8",X"89",X"68",X"03",X"38",X"0A",X"40",X"00",X"E0",X"0A",X"A8",X"07",X"30",X"09",X"00",
		X"0A",X"C2",X"4B",X"A2",X"4B",X"C4",X"4B",X"A4",X"4B",X"82",X"4B",X"84",X"4B",X"83",X"2A",X"C9",
		X"2B",X"C9",X"48",X"C7",X"48",X"ED",X"2B",X"F0",X"2B",X"F3",X"2B",X"03",X"2C",X"97",X"2C",X"CA",
		X"48",X"03",X"16",X"01",X"05",X"50",X"01",X"07",X"46",X"01",X"0B",X"6B",X"01",X"0D",X"7D",X"01",
		X"0F",X"83",X"01",X"05",X"2E",X"01",X"33",X"01",X"39",X"01",X"35",X"05",X"31",X"01",X"34",X"0C",
		X"39",X"00",X"06",X"2E",X"01",X"39",X"08",X"2E",X"02",X"39",X"05",X"2E",X"04",X"39",X"00",X"06",
		X"2E",X"01",X"39",X"11",X"2E",X"02",X"39",X"00",X"06",X"2E",X"01",X"39",X"11",X"2E",X"02",X"39",
		X"00",X"06",X"2E",X"01",X"39",X"11",X"2E",X"02",X"39",X"00",X"06",X"2E",X"01",X"39",X"01",X"33",
		X"07",X"2E",X"03",X"39",X"07",X"2E",X"01",X"39",X"00",X"05",X"2E",X"01",X"33",X"01",X"39",X"01",
		X"32",X"05",X"31",X"01",X"30",X"06",X"39",X"05",X"2E",X"01",X"39",X"00",X"05",X"2E",X"0E",X"39",
		X"06",X"2E",X"01",X"39",X"00",X"06",X"2E",X"03",X"39",X"04",X"2E",X"05",X"39",X"07",X"2E",X"01",
		X"39",X"00",X"06",X"2E",X"02",X"39",X"06",X"2E",X"03",X"39",X"07",X"2E",X"02",X"39",X"00",X"0E",
		X"2E",X"03",X"39",X"05",X"2E",X"04",X"39",X"00",X"01",X"39",X"0D",X"2E",X"02",X"39",X"05",X"2E",
		X"05",X"39",X"00",X"02",X"39",X"0B",X"2E",X"03",X"39",X"05",X"2E",X"05",X"39",X"00",X"02",X"39",
		X"06",X"2E",X"01",X"39",X"05",X"2E",X"01",X"39",X"05",X"2E",X"06",X"39",X"00",X"01",X"39",X"06",
		X"2E",X"03",X"39",X"04",X"2E",X"01",X"39",X"05",X"2E",X"06",X"39",X"00",X"01",X"39",X"05",X"2E",
		X"03",X"39",X"05",X"2E",X"01",X"39",X"06",X"2E",X"05",X"39",X"00",X"01",X"39",X"06",X"2E",X"01",
		X"39",X"06",X"2E",X"02",X"39",X"06",X"2E",X"04",X"39",X"00",X"01",X"39",X"06",X"2E",X"02",X"39",
		X"05",X"2E",X"03",X"39",X"07",X"2E",X"02",X"39",X"00",X"01",X"39",X"07",X"2E",X"02",X"39",X"05",
		X"2E",X"03",X"39",X"07",X"2E",X"01",X"39",X"00",X"01",X"39",X"07",X"2E",X"03",X"39",X"05",X"2E",
		X"03",X"39",X"06",X"2E",X"01",X"39",X"00",X"02",X"39",X"06",X"2E",X"02",X"39",X"08",X"2E",X"01",
		X"39",X"06",X"2E",X"01",X"39",X"00",X"02",X"39",X"16",X"2E",X"02",X"39",X"00",X"04",X"39",X"14",
		X"2E",X"02",X"39",X"00",X"04",X"39",X"0A",X"2E",X"01",X"39",X"08",X"2E",X"03",X"39",X"00",X"05",
		X"39",X"02",X"2E",X"02",X"39",X"04",X"2E",X"03",X"39",X"06",X"2E",X"04",X"39",X"00",X"1A",X"39",
		X"00",X"CD",X"AC",X"44",X"21",X"D7",X"70",X"77",X"C3",X"F2",X"05",X"07",X"A2",X"50",X"F5",X"01",
		X"07",X"A7",X"50",X"F6",X"07",X"07",X"A9",X"50",X"F2",X"02",X"07",X"B0",X"50",X"F5",X"07",X"02",
		X"4A",X"52",X"F5",X"03",X"07",X"12",X"53",X"F5",X"04",X"06",X"28",X"53",X"00",X"24",X"80",X"C8",
		X"24",X"D0",X"C0",X"0F",X"E8",X"A8",X"68",X"A8",X"88",X"68",X"00",X"38",X"60",X"08",X"50",X"A8",
		X"78",X"68",X"60",X"80",X"00",X"E0",X"01",X"A8",X"02",X"E0",X"01",X"A8",X"0F",X"08",X"00",X"A0",
		X"01",X"68",X"03",X"E0",X"02",X"A8",X"8C",X"08",X"00",X"60",X"02",X"08",X"03",X"E0",X"03",X"A8",
		X"8F",X"01",X"09",X"38",X"0E",X"08",X"04",X"A0",X"03",X"88",X"05",X"01",X"00",X"38",X"0E",X"08",
		X"05",X"80",X"04",X"68",X"06",X"01",X"09",X"38",X"08",X"08",X"06",X"60",X"05",X"40",X"07",X"04",
		X"00",X"38",X"08",X"08",X"07",X"38",X"06",X"00",X"07",X"04",X"00",X"60",X"09",X"40",X"92",X"60",
		X"0E",X"00",X"08",X"04",X"00",X"A0",X"95",X"68",X"08",X"60",X"98",X"00",X"09",X"02",X"00",X"E0",
		X"0A",X"A8",X"09",X"50",X"0B",X"00",X"0A",X"02",X"0C",X"E0",X"0B",X"A8",X"09",X"60",X"0F",X"58",
		X"0A",X"01",X"00",X"A0",X"0F",X"78",X"0D",X"A0",X"02",X"68",X"09",X"08",X"09",X"70",X"0C",X"68",
		X"0E",X"A0",X"02",X"68",X"09",X"08",X"00",X"60",X"0D",X"40",X"9B",X"A0",X"03",X"68",X"08",X"40",
		X"00",X"E0",X"0F",X"A8",X"0C",X"A0",X"01",X"68",X"0B",X"A2",X"48",X"C2",X"48",X"A4",X"48",X"C4",
		X"48",X"E2",X"48",X"E4",X"48",X"CB",X"2C",X"63",X"2E",X"53",X"4B",X"3B",X"4B",X"91",X"2E",X"94",
		X"2E",X"97",X"2E",X"AA",X"2E",X"5C",X"2F",X"52",X"4B",X"06",X"1B",X"01",X"0E",X"6E",X"01",X"10",
		X"46",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1A",X"39",X"00",X"03",X"39",
		X"02",X"2E",X"01",X"39",X"02",X"2E",X"08",X"39",X"03",X"2E",X"02",X"39",X"03",X"2E",X"02",X"39",
		X"00",X"02",X"39",X"08",X"2E",X"06",X"39",X"04",X"2E",X"01",X"39",X"04",X"2E",X"01",X"39",X"00",
		X"01",X"39",X"0A",X"2E",X"04",X"39",X"0A",X"2E",X"01",X"39",X"00",X"01",X"39",X"0A",X"2E",X"02",
		X"39",X"0C",X"2E",X"01",X"39",X"00",X"01",X"39",X"06",X"2E",X"01",X"39",X"04",X"2E",X"01",X"39",
		X"0C",X"2E",X"01",X"39",X"00",X"01",X"39",X"05",X"2E",X"03",X"39",X"08",X"2E",X"03",X"39",X"05",
		X"2E",X"01",X"39",X"00",X"02",X"39",X"05",X"2E",X"03",X"39",X"07",X"2E",X"02",X"39",X"06",X"2E",
		X"01",X"39",X"00",X"03",X"39",X"04",X"2E",X"03",X"39",X"06",X"2E",X"03",X"39",X"06",X"2E",X"01",
		X"39",X"00",X"02",X"39",X"05",X"2E",X"03",X"39",X"06",X"2E",X"02",X"39",X"06",X"2E",X"02",X"39",
		X"00",X"02",X"39",X"05",X"2E",X"03",X"39",X"03",X"2E",X"05",X"39",X"04",X"2E",X"04",X"39",X"00",
		X"01",X"39",X"05",X"2E",X"05",X"39",X"03",X"2E",X"04",X"39",X"04",X"2E",X"04",X"39",X"00",X"01",
		X"39",X"05",X"2E",X"06",X"39",X"03",X"2E",X"03",X"39",X"05",X"2E",X"03",X"39",X"00",X"01",X"39",
		X"04",X"2E",X"08",X"39",X"03",X"2E",X"02",X"39",X"06",X"2E",X"02",X"39",X"00",X"01",X"39",X"04",
		X"2E",X"02",X"39",X"03",X"2E",X"02",X"39",X"05",X"2E",X"02",X"39",X"06",X"2E",X"01",X"39",X"00",
		X"01",X"39",X"03",X"2E",X"03",X"39",X"0A",X"2E",X"02",X"39",X"06",X"2E",X"01",X"39",X"00",X"01",
		X"39",X"04",X"2E",X"01",X"39",X"0B",X"2E",X"03",X"39",X"05",X"2E",X"01",X"39",X"00",X"01",X"39",
		X"04",X"2E",X"01",X"39",X"0B",X"2E",X"03",X"39",X"05",X"2E",X"01",X"39",X"00",X"01",X"39",X"04",
		X"2E",X"01",X"39",X"04",X"2E",X"02",X"39",X"05",X"2E",X"03",X"39",X"05",X"2E",X"01",X"39",X"00",
		X"02",X"39",X"03",X"2E",X"01",X"39",X"04",X"2E",X"01",X"39",X"01",X"35",X"05",X"2E",X"01",X"34",
		X"01",X"39",X"01",X"35",X"05",X"2E",X"01",X"34",X"00",X"01",X"39",X"09",X"2E",X"01",X"39",X"01",
		X"33",X"05",X"2E",X"01",X"33",X"01",X"39",X"01",X"33",X"00",X"01",X"39",X"09",X"2E",X"01",X"39",
		X"01",X"33",X"06",X"2E",X"01",X"39",X"01",X"33",X"00",X"01",X"39",X"09",X"2E",X"01",X"39",X"01",
		X"33",X"06",X"2E",X"01",X"39",X"01",X"33",X"00",X"02",X"39",X"07",X"2E",X"02",X"39",X"01",X"33",
		X"06",X"2E",X"01",X"39",X"01",X"33",X"00",X"03",X"39",X"02",X"2E",X"01",X"39",X"02",X"2E",X"03",
		X"39",X"01",X"33",X"06",X"2E",X"01",X"39",X"01",X"33",X"00",X"0B",X"39",X"01",X"33",X"05",X"2E",
		X"01",X"33",X"01",X"39",X"01",X"33",X"05",X"2E",X"01",X"33",X"00",X"2A",X"0C",X"74",X"09",X"23",
		X"22",X"0C",X"74",X"F5",X"05",X"07",X"A7",X"50",X"F2",X"08",X"03",X"A2",X"51",X"F4",X"07",X"03",
		X"0C",X"52",X"F5",X"02",X"05",X"6C",X"52",X"F5",X"06",X"02",X"02",X"53",X"F6",X"07",X"07",X"0D",
		X"53",X"F5",X"01",X"07",X"15",X"53",X"F4",X"05",X"07",X"16",X"53",X"F5",X"01",X"07",X"1B",X"53",
		X"00",X"44",X"70",X"38",X"44",X"30",X"40",X"12",X"00",X"40",X"68",X"00",X"28",X"48",X"80",X"E8",
		X"A8",X"88",X"48",X"E8",X"B0",X"B0",X"88",X"88",X"78",X"48",X"80",X"00",X"40",X"02",X"08",X"01",
		X"48",X"12",X"00",X"01",X"04",X"00",X"68",X"03",X"48",X"01",X"48",X"11",X"00",X"02",X"04",X"00",
		X"98",X"9E",X"70",X"02",X"48",X"AD",X"00",X"03",X"04",X"00",X"E0",X"04",X"A0",X"03",X"28",X"05",
		X"00",X"04",X"02",X"00",X"E0",X"05",X"A0",X"03",X"48",X"06",X"30",X"04",X"02",X"00",X"E0",X"06",
		X"88",X"10",X"80",X"07",X"50",X"05",X"02",X"09",X"E0",X"07",X"88",X"0E",X"A8",X"A1",X"88",X"06",
		X"08",X"00",X"E0",X"08",X"A8",X"09",X"E0",X"08",X"B0",X"07",X"08",X"0C",X"A0",X"08",X"88",X"0A",
		X"E0",X"09",X"B0",X"07",X"08",X"00",X"80",X"09",X"48",X"0B",X"E0",X"0A",X"B0",X"0E",X"08",X"09",
		X"40",X"0A",X"38",X"0C",X"E0",X"0B",X"B0",X"0D",X"01",X"00",X"30",X"0B",X"08",X"0C",X"E0",X"0C",
		X"B0",X"0D",X"01",X"00",X"40",X"0E",X"08",X"0D",X"A8",X"A4",X"88",X"12",X"01",X"00",X"80",X"07",
		X"48",X"0D",X"A8",X"0A",X"88",X"A7",X"01",X"09",X"68",X"10",X"48",X"12",X"80",X"0E",X"78",X"11",
		X"08",X"0F",X"80",X"06",X"70",X"AA",X"80",X"0E",X"50",X"03",X"08",X"00",X"68",X"10",X"48",X"12",
		X"70",X"0F",X"50",X"02",X"40",X"00",X"40",X"AA",X"08",X"12",X"80",X"0D",X"50",X"01",X"D6",X"4B",
		X"D8",X"4B",X"B6",X"4B",X"B8",X"4B",X"96",X"4B",X"98",X"4B",X"2E",X"13",X"5E",X"CD",X"15",X"50",
		X"5F",X"21",X"13",X"74",X"4E",X"CD",X"E8",X"4E",X"21",X"13",X"74",X"34",X"C2",X"5A",X"50",X"C9",
		X"21",X"19",X"74",X"36",X"00",X"2D",X"36",X"00",X"0E",X"1B",X"0D",X"79",X"21",X"18",X"74",X"96",
		X"DA",X"B0",X"50",X"4E",X"CD",X"DB",X"4E",X"0F",X"D2",X"9F",X"50",X"21",X"19",X"74",X"34",X"21",
		X"19",X"74",X"7E",X"D6",X"02",X"DA",X"AB",X"50",X"3E",X"FF",X"C9",X"2D",X"34",X"C2",X"88",X"50",
		X"AF",X"C9",X"21",X"1A",X"74",X"36",X"00",X"0E",X"1B",X"0D",X"79",X"21",X"1A",X"74",X"96",X"DA",
		X"D3",X"50",X"4E",X"CD",X"DB",X"4E",X"0F",X"D2",X"CC",X"50",X"AF",X"C9",X"21",X"1A",X"74",X"34",
		X"C2",X"B7",X"50",X"3E",X"FF",X"C9",X"CD",X"12",X"50",X"CD",X"C3",X"46",X"CD",X"D2",X"43",X"21",
		X"07",X"74",X"77",X"2C",X"36",X"00",X"21",X"07",X"74",X"7E",X"D6",X"41",X"9F",X"2F",X"4F",X"3E",
		X"5A",X"96",X"9F",X"2F",X"A1",X"5F",X"7E",X"D6",X"30",X"9F",X"2F",X"D5",X"4F",X"3E",X"39",X"96");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
