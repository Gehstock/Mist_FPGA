library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity gfx1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of gfx1 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"7C",X"82",X"82",X"82",X"7C",X"00",X"00",X"00",X"00",X"42",X"FE",X"02",X"00",X"00",X"00",
		X"00",X"46",X"8A",X"92",X"92",X"62",X"00",X"00",X"00",X"84",X"82",X"92",X"B2",X"CC",X"00",X"00",
		X"00",X"18",X"28",X"48",X"FE",X"08",X"00",X"00",X"00",X"E4",X"A2",X"A2",X"A2",X"9C",X"00",X"00",
		X"00",X"3C",X"52",X"92",X"92",X"8C",X"00",X"00",X"00",X"80",X"80",X"9E",X"A0",X"C0",X"00",X"00",
		X"00",X"6C",X"92",X"92",X"92",X"6C",X"00",X"00",X"00",X"62",X"92",X"92",X"94",X"78",X"00",X"00",
		X"00",X"7E",X"90",X"90",X"90",X"7E",X"00",X"00",X"00",X"FE",X"92",X"92",X"92",X"6C",X"00",X"00",
		X"00",X"7C",X"82",X"82",X"82",X"44",X"00",X"00",X"00",X"FE",X"82",X"82",X"82",X"7C",X"00",X"00",
		X"00",X"FE",X"92",X"92",X"92",X"82",X"00",X"00",X"00",X"FE",X"90",X"90",X"90",X"80",X"00",X"00",
		X"00",X"7C",X"82",X"82",X"92",X"9E",X"00",X"00",X"00",X"FE",X"10",X"10",X"10",X"FE",X"00",X"00",
		X"00",X"00",X"82",X"FE",X"82",X"00",X"00",X"00",X"00",X"04",X"02",X"02",X"02",X"FC",X"00",X"00",
		X"00",X"FE",X"10",X"38",X"44",X"82",X"00",X"00",X"00",X"FE",X"02",X"02",X"02",X"02",X"00",X"00",
		X"00",X"FE",X"40",X"30",X"40",X"FE",X"00",X"00",X"00",X"FE",X"20",X"10",X"08",X"FE",X"00",X"00",
		X"00",X"7C",X"82",X"82",X"82",X"7C",X"00",X"00",X"00",X"FE",X"90",X"90",X"90",X"60",X"00",X"00",
		X"00",X"7C",X"82",X"8A",X"84",X"7A",X"00",X"00",X"00",X"FE",X"90",X"98",X"94",X"62",X"00",X"00",
		X"00",X"64",X"92",X"92",X"92",X"4C",X"00",X"00",X"00",X"80",X"80",X"FE",X"80",X"80",X"00",X"00",
		X"00",X"FC",X"02",X"02",X"02",X"FC",X"00",X"00",X"00",X"F8",X"04",X"02",X"04",X"F8",X"00",X"00",
		X"00",X"FE",X"04",X"18",X"04",X"FE",X"00",X"00",X"00",X"C6",X"28",X"10",X"28",X"C6",X"00",X"00",
		X"00",X"C0",X"20",X"1E",X"20",X"C0",X"00",X"00",X"00",X"86",X"8A",X"92",X"A2",X"C2",X"00",X"00",
		X"00",X"7C",X"82",X"BA",X"8A",X"7A",X"00",X"00",X"00",X"38",X"44",X"82",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"82",X"44",X"38",X"00",X"00",X"00",X"40",X"80",X"9A",X"A0",X"40",X"00",X"00",
		X"00",X"10",X"10",X"7C",X"10",X"10",X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"00",X"00",
		X"00",X"44",X"28",X"FE",X"28",X"44",X"00",X"00",X"00",X"04",X"08",X"10",X"20",X"40",X"00",X"00",
		X"00",X"28",X"28",X"28",X"28",X"28",X"00",X"00",X"00",X"00",X"06",X"06",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3C",X"3C",X"3F",X"3F",X"3F",X"3F",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"3C",X"3C",X"FC",X"FC",X"FC",X"FC",X"00",X"00",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",
		X"00",X"00",X"3F",X"3F",X"3F",X"3F",X"3C",X"3C",X"00",X"00",X"FC",X"FC",X"FC",X"FC",X"3C",X"3C",
		X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"28",X"10",X"00",X"00",X"00",
		X"00",X"10",X"38",X"6C",X"38",X"10",X"00",X"00",X"10",X"54",X"38",X"EE",X"38",X"54",X"10",X"00",
		X"00",X"10",X"54",X"38",X"EE",X"38",X"54",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"54",X"38",X"EE",X"38",X"54",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"54",X"38",X"EE",X"38",X"54",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"54",X"38",X"EE",X"38",X"54",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"54",X"38",X"EE",X"38",X"54",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"54",X"38",X"EE",X"38",X"54",X"10",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"54",X"38",X"EE",X"38",X"54",X"10",X"00",X"00",
		X"08",X"2A",X"1C",X"77",X"1C",X"2A",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"15",X"0E",X"3B",X"0E",X"15",X"04",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",
		X"02",X"0A",X"07",X"1D",X"07",X"0A",X"02",X"00",X"00",X"80",X"00",X"C0",X"00",X"80",X"00",X"00",
		X"01",X"05",X"03",X"0E",X"03",X"05",X"01",X"00",X"00",X"40",X"80",X"E0",X"80",X"40",X"00",X"00",
		X"00",X"02",X"01",X"07",X"01",X"02",X"00",X"00",X"80",X"A0",X"C0",X"70",X"C0",X"A0",X"80",X"00",
		X"00",X"01",X"00",X"03",X"00",X"01",X"00",X"00",X"40",X"50",X"E0",X"B8",X"E0",X"50",X"40",X"00",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"20",X"A8",X"70",X"DC",X"70",X"A8",X"20",X"00",
		X"1C",X"3E",X"7F",X"7F",X"7F",X"3E",X"1C",X"00",X"01",X"06",X"18",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"20",X"28",X"30",X"3C",X"00",X"00",X"00",X"00",X"04",X"14",X"0C",X"3C",X"00",X"00",
		X"00",X"00",X"3C",X"30",X"28",X"20",X"00",X"00",X"00",X"00",X"3C",X"0C",X"14",X"04",X"00",X"00",
		X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"10",X"54",X"38",X"EE",X"38",X"54",X"10",X"00",X"00",X"10",X"54",X"38",X"EE",X"38",X"54",X"10",
		X"10",X"00",X"10",X"54",X"38",X"EE",X"38",X"54",X"54",X"10",X"00",X"10",X"54",X"38",X"EE",X"38",
		X"38",X"54",X"10",X"00",X"10",X"54",X"38",X"EE",X"EE",X"38",X"54",X"10",X"00",X"10",X"54",X"38",
		X"38",X"EE",X"38",X"54",X"10",X"00",X"10",X"54",X"54",X"38",X"EE",X"38",X"54",X"10",X"00",X"10",
		X"10",X"54",X"38",X"EE",X"38",X"54",X"10",X"00",X"08",X"2A",X"1C",X"77",X"1C",X"2A",X"08",X"00",
		X"04",X"15",X"0E",X"BB",X"0E",X"15",X"04",X"00",X"02",X"8A",X"07",X"DD",X"07",X"8A",X"02",X"00",
		X"01",X"45",X"83",X"EE",X"83",X"45",X"01",X"00",X"80",X"A2",X"C1",X"77",X"C1",X"A2",X"80",X"00",
		X"40",X"51",X"E0",X"BB",X"E0",X"51",X"40",X"00",X"20",X"A8",X"70",X"DD",X"70",X"A8",X"20",X"00",
		X"FF",X"FF",X"C6",X"C0",X"C0",X"80",X"00",X"00",X"FF",X"FF",X"EF",X"EF",X"EF",X"EF",X"00",X"00",
		X"FF",X"FF",X"FF",X"7F",X"7F",X"FF",X"0F",X"03",X"FF",X"FF",X"80",X"00",X"1C",X"FF",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"A0",X"00",X"0F",X"1F",X"0F",X"1F",X"07",X"0B",X"02",X"00",
		X"FF",X"FF",X"E3",X"E0",X"E0",X"C0",X"00",X"00",X"FF",X"83",X"83",X"83",X"83",X"83",X"83",X"00",
		X"FF",X"FF",X"FF",X"7F",X"7F",X"FF",X"1E",X"06",X"FF",X"FF",X"80",X"00",X"38",X"FF",X"00",X"00",
		X"FF",X"FF",X"D8",X"C0",X"C0",X"80",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7E",X"28",
		X"FF",X"FF",X"FF",X"7F",X"7F",X"FF",X"0F",X"03",X"FF",X"FF",X"80",X"00",X"0E",X"FF",X"00",X"00",
		X"00",X"10",X"28",X"28",X"10",X"00",X"00",X"00",X"00",X"10",X"28",X"44",X"44",X"44",X"28",X"00",
		X"00",X"00",X"10",X"00",X"44",X"44",X"00",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"C6",X"FF",X"FF",
		X"00",X"00",X"EF",X"EF",X"EF",X"EF",X"FF",X"FF",X"03",X"0F",X"FF",X"7F",X"7F",X"FF",X"FF",X"FF",
		X"00",X"00",X"FF",X"1C",X"00",X"80",X"FF",X"FF",X"00",X"A0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"02",X"0B",X"07",X"1F",X"0F",X"1F",X"0F",X"00",X"00",X"C0",X"E0",X"E0",X"E3",X"FF",X"FF",
		X"00",X"83",X"83",X"83",X"83",X"83",X"83",X"FF",X"06",X"1E",X"FF",X"7F",X"7F",X"FF",X"FF",X"FF",
		X"00",X"00",X"FF",X"38",X"00",X"80",X"FF",X"FF",X"00",X"00",X"80",X"C0",X"C0",X"D8",X"FF",X"FF",
		X"28",X"7E",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"03",X"0F",X"FF",X"7F",X"7F",X"FF",X"FF",X"FF",
		X"00",X"00",X"FF",X"0E",X"00",X"80",X"FF",X"FF",X"00",X"00",X"00",X"10",X"28",X"28",X"10",X"00",
		X"00",X"28",X"44",X"44",X"44",X"28",X"10",X"00",X"82",X"00",X"44",X"44",X"00",X"10",X"00",X"00",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",
		X"FF",X"FF",X"C6",X"C0",X"C0",X"80",X"00",X"00",X"FF",X"DF",X"EF",X"EF",X"EF",X"EF",X"00",X"00",
		X"FF",X"FF",X"FF",X"7F",X"7F",X"FF",X"0F",X"03",X"FF",X"80",X"0C",X"18",X"8C",X"FF",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"A0",X"00",X"0F",X"1F",X"0F",X"1F",X"07",X"0B",X"02",X"00",
		X"FF",X"FF",X"E3",X"E0",X"E0",X"C0",X"00",X"00",X"FF",X"C7",X"E7",X"E3",X"E3",X"E3",X"E3",X"00",
		X"FF",X"FF",X"FF",X"7F",X"7F",X"FF",X"1E",X"06",X"FF",X"80",X"18",X"30",X"98",X"FF",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"A0",X"00",X"0F",X"1F",X"0F",X"1F",X"07",X"0B",X"02",X"00",
		X"00",X"00",X"80",X"C0",X"C0",X"C6",X"FF",X"FF",X"00",X"00",X"EF",X"EF",X"EF",X"EF",X"DF",X"FF",
		X"03",X"0F",X"FF",X"7F",X"7F",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"8C",X"18",X"0C",X"80",X"FF",
		X"00",X"A0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"02",X"0B",X"07",X"1F",X"0F",X"1F",X"0F",
		X"00",X"00",X"C0",X"E0",X"E0",X"E3",X"FF",X"FF",X"00",X"E3",X"E3",X"E3",X"E3",X"E7",X"C7",X"FF",
		X"06",X"1E",X"FF",X"7F",X"7F",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"98",X"30",X"18",X"80",X"FF",
		X"00",X"A0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"02",X"0B",X"07",X"1F",X"0F",X"1F",X"0F",
		X"3C",X"42",X"99",X"A5",X"A5",X"A5",X"42",X"3C",X"00",X"00",X"00",X"FA",X"00",X"00",X"00",X"00",
		X"FE",X"90",X"98",X"94",X"62",X"00",X"FC",X"02",X"02",X"FC",X"00",X"FE",X"92",X"92",X"92",X"6C",
		X"FE",X"92",X"92",X"82",X"00",X"FE",X"20",X"10",X"08",X"FE",X"00",X"FE",X"82",X"82",X"82",X"7C",
		X"00",X"00",X"D0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"00",X"00",
		X"3C",X"3C",X"3F",X"3F",X"3F",X"3F",X"3C",X"3C",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"84",X"82",X"92",X"B2",X"CC",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"18",X"28",X"48",X"FE",X"08",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
