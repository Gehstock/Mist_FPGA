library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity mw04 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of mw04 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"01",X"B8",X"03",X"5C",X"07",X"EE",X"0E",X"F3",X"19",X"FF",X"1F",X"F8",X"03",X"FF",X"1F",X"F3",
		X"19",X"EE",X"0E",X"5C",X"07",X"B8",X"03",X"B0",X"01",X"00",X"00",X"3B",X"18",X"00",X"00",X"80",
		X"07",X"80",X"0F",X"C0",X"1D",X"E0",X"3B",X"F8",X"67",X"5E",X"7C",X"C7",X"08",X"5E",X"7C",X"F8",
		X"67",X"E0",X"3B",X"C0",X"1D",X"80",X"0F",X"80",X"07",X"00",X"00",X"1B",X"18",X"00",X"00",X"80",
		X"07",X"80",X"0F",X"C0",X"1D",X"E0",X"3B",X"F8",X"7F",X"5E",X"7C",X"FF",X"08",X"5E",X"7C",X"F8",
		X"7F",X"E0",X"3B",X"C0",X"1D",X"80",X"0F",X"80",X"07",X"00",X"00",X"7B",X"18",X"00",X"00",X"F0",
		X"0F",X"80",X"1F",X"80",X"34",X"E0",X"6F",X"38",X"79",X"9E",X"30",X"BF",X"1F",X"9E",X"30",X"38",
		X"79",X"E0",X"6F",X"80",X"34",X"80",X"1F",X"F0",X"0F",X"00",X"00",X"5B",X"18",X"00",X"00",X"F0",
		X"0F",X"80",X"1F",X"80",X"34",X"E0",X"6F",X"38",X"7F",X"9E",X"36",X"B1",X"1F",X"9E",X"36",X"38",
		X"7F",X"E0",X"6F",X"80",X"34",X"80",X"1F",X"F0",X"0F",X"00",X"00",X"BB",X"18",X"00",X"00",X"F0",
		X"0F",X"C8",X"13",X"40",X"02",X"E0",X"07",X"70",X"5F",X"BF",X"7B",X"58",X"70",X"BF",X"7B",X"70",
		X"5F",X"E0",X"07",X"40",X"02",X"C8",X"13",X"F0",X"0F",X"00",X"00",X"9B",X"18",X"00",X"00",X"F0",
		X"0F",X"C8",X"13",X"40",X"02",X"E0",X"07",X"70",X"5F",X"BF",X"7B",X"5E",X"7C",X"BF",X"7B",X"70",
		X"5F",X"E0",X"07",X"40",X"02",X"C8",X"13",X"F0",X"0F",X"00",X"00",X"FB",X"18",X"00",X"00",X"F0",
		X"01",X"F8",X"03",X"0C",X"06",X"06",X"0C",X"E3",X"18",X"BF",X"1F",X"1F",X"1F",X"BF",X"1F",X"E3",
		X"18",X"06",X"0C",X"0C",X"06",X"F8",X"03",X"F0",X"01",X"00",X"00",X"1B",X"19",X"00",X"00",X"F0",
		X"01",X"F8",X"03",X"0C",X"07",X"06",X"0F",X"E3",X"1F",X"B3",X"19",X"13",X"19",X"B3",X"19",X"FF",
		X"18",X"1E",X"0C",X"1C",X"06",X"F8",X"03",X"F0",X"01",X"00",X"00",X"3B",X"19",X"00",X"00",X"F0",
		X"01",X"F8",X"03",X"EC",X"06",X"E6",X"0C",X"E3",X"18",X"B3",X"19",X"13",X"19",X"B3",X"19",X"E3",
		X"18",X"E6",X"0C",X"EC",X"06",X"F8",X"03",X"F0",X"01",X"00",X"00",X"DB",X"18",X"00",X"00",X"F0",
		X"01",X"F8",X"03",X"1C",X"06",X"1E",X"0C",X"FF",X"18",X"B3",X"19",X"13",X"19",X"B3",X"19",X"E3",
		X"1F",X"06",X"0F",X"0C",X"07",X"F8",X"03",X"F0",X"01",X"00",X"00",X"68",X"19",X"00",X"1C",X"2A",
		X"75",X"6B",X"75",X"3D",X"2F",X"1E",X"0C",X"00",X"75",X"19",X"00",X"0C",X"1E",X"2F",X"3B",X"65",
		X"7B",X"7D",X"32",X"1C",X"00",X"82",X"19",X"00",X"18",X"3C",X"7E",X"5A",X"5F",X"6B",X"57",X"2A",
		X"1C",X"00",X"5B",X"19",X"00",X"1C",X"26",X"5B",X"6F",X"5D",X"72",X"7E",X"3C",X"18",X"00",X"59",
		X"1A",X"03",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"1F",X"00",X"00",X"00",X"00",
		X"3E",X"00",X"00",X"00",X"00",X"7C",X"00",X"00",X"00",X"00",X"F8",X"00",X"00",X"00",X"00",X"F0",
		X"01",X"00",X"00",X"00",X"E0",X"03",X"00",X"00",X"00",X"C0",X"0F",X"00",X"00",X"00",X"80",X"1F",
		X"00",X"00",X"00",X"00",X"2F",X"00",X"00",X"10",X"00",X"7E",X"00",X"00",X"00",X"00",X"7E",X"00",
		X"00",X"00",X"00",X"FC",X"00",X"00",X"00",X"00",X"E8",X"03",X"00",X"00",X"00",X"D0",X"0B",X"00",
		X"00",X"00",X"F0",X"15",X"00",X"00",X"00",X"A0",X"2B",X"00",X"00",X"00",X"40",X"55",X"00",X"00",
		X"00",X"80",X"EA",X"00",X"00",X"00",X"00",X"DD",X"03",X"00",X"00",X"00",X"36",X"05",X"00",X"00",
		X"00",X"AA",X"08",X"00",X"00",X"00",X"1C",X"1B",X"00",X"00",X"00",X"58",X"36",X"00",X"00",X"00",
		X"A0",X"59",X"00",X"00",X"00",X"40",X"67",X"00",X"00",X"00",X"C0",X"CC",X"01",X"00",X"00",X"80",
		X"45",X"01",X"00",X"00",X"00",X"AB",X"03",X"00",X"00",X"00",X"50",X"06",X"00",X"00",X"00",X"A4",
		X"0C",X"00",X"00",X"00",X"8C",X"05",X"00",X"00",X"00",X"18",X"09",X"00",X"00",X"00",X"30",X"11",
		X"00",X"00",X"00",X"40",X"02",X"00",X"00",X"00",X"80",X"04",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"8F",X"19",X"03",X"00",X"00",X"00",X"00",
		X"0F",X"00",X"00",X"00",X"00",X"1F",X"00",X"00",X"00",X"00",X"3E",X"00",X"00",X"00",X"00",X"7C",
		X"00",X"00",X"00",X"00",X"F8",X"00",X"00",X"00",X"00",X"F0",X"01",X"00",X"00",X"00",X"E0",X"07",
		X"00",X"00",X"00",X"C0",X"0F",X"00",X"00",X"00",X"80",X"1F",X"00",X"00",X"00",X"00",X"2F",X"00",
		X"00",X"00",X"00",X"6E",X"00",X"00",X"00",X"00",X"DA",X"00",X"00",X"00",X"00",X"EC",X"01",X"00",
		X"00",X"00",X"A8",X"03",X"00",X"00",X"00",X"5C",X"0B",X"00",X"00",X"00",X"E0",X"16",X"00",X"00",
		X"00",X"A0",X"2D",X"00",X"00",X"00",X"C0",X"71",X"00",X"00",X"00",X"80",X"E5",X"00",X"00",X"00",
		X"00",X"CB",X"01",X"00",X"00",X"00",X"36",X"05",X"00",X"00",X"00",X"68",X"02",X"00",X"00",X"00",
		X"94",X"0C",X"00",X"00",X"00",X"48",X"39",X"00",X"00",X"00",X"90",X"52",X"00",X"00",X"00",X"20",
		X"A5",X"00",X"00",X"00",X"C0",X"48",X"01",X"00",X"00",X"80",X"05",X"02",X"00",X"00",X"00",X"2B",
		X"05",X"00",X"00",X"00",X"54",X"0A",X"00",X"00",X"00",X"A8",X"14",X"00",X"00",X"00",X"94",X"01",
		X"00",X"00",X"00",X"08",X"01",X"00",X"00",X"00",X"10",X"02",X"00",X"00",X"00",X"20",X"04",X"00",
		X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"23",X"1B",X"00",X"00",X"20",X"00",X"30",X"00",X"30",X"00",X"30",X"00",X"34",
		X"00",X"3C",X"00",X"2C",X"00",X"7C",X"00",X"7C",X"00",X"3C",X"00",X"3C",X"00",X"3C",X"00",X"3C",
		X"00",X"3C",X"00",X"BC",X"00",X"7C",X"00",X"7C",X"00",X"7C",X"01",X"FE",X"00",X"7E",X"00",X"FE",
		X"00",X"FE",X"01",X"7E",X"03",X"FE",X"0F",X"7E",X"0F",X"FC",X"01",X"FC",X"03",X"FC",X"00",X"7C",
		X"01",X"7C",X"02",X"7C",X"04",X"3C",X"00",X"38",X"00",X"3C",X"00",X"7A",X"00",X"B8",X"00",X"38",
		X"00",X"10",X"00",X"00",X"00",X"75",X"1B",X"40",X"A0",X"00",X"60",X"FF",X"F0",X"FF",X"60",X"00",
		X"A0",X"40",X"82",X"1B",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"00",X"6C",X"00",X"FE",X"03",X"6C",X"00",X"38",X"00",X"F7",X"01",X"7F",X"1F",X"1E",X"FE",X"7F",
		X"1F",X"F7",X"01",X"38",X"00",X"6C",X"00",X"FE",X"03",X"6C",X"00",X"00",X"00",X"B9",X"1B",X"00",
		X"00",X"1C",X"0E",X"3B",X"3B",X"0E",X"1C",X"00",X"00",X"AD",X"1B",X"00",X"00",X"1C",X"0E",X"3F",
		X"3F",X"0E",X"1C",X"00",X"00",X"E3",X"1B",X"3E",X"7C",X"63",X"C6",X"DD",X"BB",X"DD",X"BB",X"63",
		X"C6",X"3E",X"7C",X"00",X"00",X"00",X"00",X"3E",X"7C",X"63",X"C6",X"DD",X"BB",X"DD",X"BB",X"63",
		X"C6",X"3E",X"7C",X"C5",X"1B",X"3E",X"7C",X"6B",X"B6",X"D5",X"AB",X"D5",X"AB",X"6B",X"D6",X"BE",
		X"7D",X"C0",X"03",X"C0",X"03",X"BE",X"7D",X"6B",X"D6",X"D5",X"AB",X"D5",X"AB",X"6B",X"D6",X"3E",
		X"7C",X"0D",X"1C",X"00",X"00",X"3C",X"05",X"FF",X"1F",X"3C",X"05",X"00",X"00",X"01",X"1C",X"00",
		X"00",X"3C",X"05",X"F7",X"1F",X"3C",X"05",X"00",X"00",X"80",X"00",X"80",X"02",X"50",X"48",X"54",
		X"21",X"2A",X"04",X"40",X"0B",X"A8",X"24",X"D2",X"0D",X"E0",X"0A",X"F8",X"C7",X"F0",X"24",X"61",
		X"04",X"D8",X"1A",X"54",X"25",X"00",X"02",X"88",X"15",X"A4",X"22",X"00",X"00",X"80",X"00",X"54",
		X"2A",X"BB",X"56",X"30",X"E8",X"30",X"56",X"B3",X"2A",X"94",X"80",X"B4",X"28",X"1D",X"80",X"43",
		X"52",X"24",X"80",X"5C",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"10",X"20",X"00",X"40",X"20",
		X"39",X"12",X"2A",X"80",X"C8",X"46",X"09",X"04",X"10",X"95",X"8F",X"A7",X"02",X"00",X"88",X"F1",
		X"5E",X"04",X"00",X"55",X"34",X"29",X"22",X"90",X"B2",X"D2",X"76",X"11",X"24",X"F5",X"6F",X"4B",
		X"08",X"40",X"FF",X"FF",X"BB",X"02",X"C0",X"FF",X"FF",X"7F",X"02",X"BB",X"FF",X"FF",X"FF",X"DD",
		X"C0",X"FF",X"FF",X"7F",X"00",X"20",X"DF",X"FF",X"1F",X"03",X"00",X"F5",X"EF",X"C9",X"20",X"92",
		X"EC",X"52",X"76",X"49",X"48",X"CA",X"7C",X"77",X"10",X"04",X"A5",X"97",X"0D",X"00",X"10",X"52",
		X"6A",X"55",X"09",X"08",X"28",X"D5",X"22",X"13",X"00",X"94",X"38",X"05",X"00",X"00",X"04",X"10",
		X"08",X"00",X"00",X"20",X"10",X"00",X"00",X"1A",X"2C",X"0C",X"03",X"0D",X"18",X"0C",X"14",X"12",
		X"17",X"10",X"2E",X"1D",X"12",X"16",X"0E",X"00",X"18",X"28",X"05",X"03",X"1B",X"0E",X"0A",X"0D",
		X"22",X"00",X"10",X"29",X"12",X"00",X"10",X"0A",X"16",X"0E",X"2E",X"18",X"1F",X"0E",X"1B",X"2E",
		X"19",X"15",X"0A",X"22",X"0E",X"1B",X"2E",X"01",X"00",X"10",X"29",X"12",X"00",X"10",X"0A",X"16",
		X"0E",X"2E",X"18",X"1F",X"0E",X"1B",X"2E",X"19",X"15",X"0A",X"22",X"0E",X"1B",X"2E",X"02",X"00",
		X"10",X"2B",X"0D",X"00",X"1D",X"1B",X"22",X"2E",X"19",X"15",X"0A",X"22",X"0E",X"1B",X"24",X"01",
		X"25",X"00",X"10",X"2B",X"0D",X"00",X"1D",X"1B",X"22",X"2E",X"19",X"15",X"0A",X"22",X"0E",X"1B",
		X"24",X"02",X"25",X"00",X"1E",X"25",X"1A",X"00",X"1C",X"0C",X"18",X"1B",X"0E",X"24",X"01",X"25",
		X"2E",X"11",X"12",X"2B",X"1C",X"0C",X"18",X"1B",X"0E",X"2E",X"1C",X"0C",X"18",X"1B",X"0E",X"24",
		X"02",X"25",X"00",X"1C",X"2D",X"05",X"00",X"19",X"18",X"12",X"17",X"1D",X"00",X"01",X"36",X"06",
		X"00",X"0C",X"1B",X"0E",X"0D",X"12",X"1D",X"00",X"01",X"25",X"06",X"00",X"0E",X"17",X"0E",X"1B",
		X"10",X"22",X"00",X"14",X"30",X"04",X"0F",X"19",X"1E",X"1C",X"11",X"01",X"12",X"2A",X"0F",X"0F",
		X"01",X"2E",X"19",X"15",X"0A",X"22",X"0E",X"1B",X"2E",X"0B",X"1E",X"1D",X"1D",X"18",X"17",X"00",
		X"10",X"2A",X"10",X"0F",X"02",X"2E",X"19",X"15",X"0A",X"22",X"0E",X"1B",X"1C",X"2E",X"0B",X"1E",
		X"1D",X"1D",X"18",X"17",X"00",X"03",X"27",X"15",X"00",X"27",X"2E",X"1C",X"11",X"12",X"17",X"2E",
		X"17",X"12",X"11",X"18",X"17",X"2E",X"14",X"12",X"14",X"0A",X"14",X"1E",X"2E",X"27",X"00",X"1A",
		X"2C",X"0A",X"1F",X"18",X"23",X"16",X"0A",X"2E",X"2E",X"20",X"0A",X"1B",X"1C",X"01",X"18",X"2F",
		X"05",X"1F",X"15",X"0E",X"1D",X"2F",X"1C",X"01",X"16",X"2B",X"0C",X"1F",X"1D",X"1B",X"0A",X"1F",
		X"0E",X"15",X"29",X"0F",X"12",X"10",X"11",X"1D",X"01",X"14",X"2B",X"0B",X"1F",X"1C",X"19",X"0A",
		X"0C",X"0E",X"2E",X"20",X"18",X"1B",X"15",X"0D",X"00",X"10",X"2E",X"07",X"00",X"27",X"1C",X"0C",
		X"18",X"1B",X"0E",X"27",X"01",X"0E",X"2B",X"0E",X"00",X"1E",X"0F",X"18",X"2E",X"2E",X"2E",X"2E",
		X"01",X"00",X"00",X"2C",X"05",X"00",X"00",X"01",X"0C",X"2B",X"0C",X"00",X"16",X"0E",X"1D",X"0E",
		X"18",X"2E",X"2E",X"05",X"00",X"2C",X"07",X"00",X"01",X"0A",X"2B",X"0A",X"00",X"0C",X"18",X"16",
		X"0E",X"1D",X"2E",X"2E",X"08",X"00",X"00",X"00",X"12",X"2A",X"0F",X"00",X"27",X"0C",X"11",X"0A",
		X"1B",X"10",X"0E",X"2E",X"0E",X"17",X"0E",X"1B",X"10",X"22",X"27",X"01",X"10",X"2B",X"0F",X"00",
		X"0D",X"18",X"0C",X"14",X"12",X"17",X"10",X"2E",X"2E",X"2A",X"01",X"05",X"00",X"00",X"00",X"01",
		X"0E",X"29",X"13",X"00",X"27",X"0C",X"1B",X"0A",X"1C",X"11",X"2E",X"15",X"18",X"1C",X"1D",X"2E",
		X"0E",X"17",X"0E",X"1B",X"10",X"22",X"27",X"01",X"0C",X"2B",X"0F",X"00",X"1E",X"0F",X"18",X"2E",
		X"2E",X"2E",X"2E",X"2E",X"2E",X"2B",X"01",X"05",X"00",X"00",X"00",X"01",X"0A",X"2B",X"0E",X"00",
		X"16",X"0E",X"1D",X"0E",X"18",X"2E",X"2E",X"2E",X"2E",X"2B",X"08",X"00",X"00",X"00",X"01",X"08",
		X"2B",X"0F",X"00",X"0C",X"18",X"16",X"0E",X"1D",X"2E",X"2E",X"2E",X"2E",X"2B",X"02",X"00",X"00",
		X"00",X"00",X"01",X"06",X"2B",X"0F",X"00",X"16",X"12",X"1C",X"1C",X"12",X"15",X"0E",X"2E",X"2E",
		X"2B",X"01",X"00",X"00",X"00",X"00",X"00",X"14",X"2D",X"0B",X"00",X"12",X"17",X"1C",X"0E",X"1B",
		X"1D",X"2E",X"0C",X"18",X"12",X"17",X"01",X"12",X"2B",X"0E",X"00",X"01",X"2E",X"18",X"1B",X"2E",
		X"02",X"2E",X"19",X"15",X"0A",X"22",X"0E",X"1B",X"1C",X"01",X"10",X"2B",X"0F",X"00",X"01",X"2E",
		X"19",X"15",X"0A",X"22",X"0E",X"1B",X"2E",X"01",X"2E",X"0C",X"18",X"12",X"17",X"01",X"0E",X"2A",
		X"11",X"00",X"02",X"2E",X"19",X"15",X"0A",X"22",X"0E",X"1B",X"1C",X"2E",X"02",X"2E",X"0C",X"18",
		X"12",X"17",X"1C",X"00",X"DE",X"88",X"D0",X"B8",X"C2",X"26",X"B6",X"CC",X"B0",X"60",X"A8",X"44",
		X"A6",X"9C",X"9A",X"FC",X"8B",X"C8",X"7C",X"90",X"76",X"24",X"7C",X"90",X"68",X"C0",X"60",X"60",
		X"4C",X"DC",X"48",X"84",X"3E",X"30",X"34",X"F8",X"2C",X"48",X"18",X"30",X"07",X"07",X"07",X"07",
		X"45",X"1F",X"0A",X"15",X"0A",X"40",X"1F",X"15",X"0A",X"15",X"51",X"1F",X"00",X"0A",X"07",X"0A",
		X"00",X"58",X"1F",X"00",X"05",X"0E",X"05",X"00",X"5F",X"1F",X"00",X"0A",X"0D",X"0A",X"00",X"4A",
		X"1F",X"00",X"05",X"0B",X"05",X"00",X"66",X"1F",X"FF",X"0F",X"6A",X"1F",X"00",X"00",X"80",X"07",
		X"E0",X"1B",X"F8",X"77",X"47",X"5C",X"FC",X"77",X"F0",X"3B",X"E0",X"1D",X"C0",X"0F",X"80",X"07",
		X"00",X"00",X"A6",X"1F",X"00",X"00",X"00",X"00",X"D8",X"00",X"DC",X"01",X"FE",X"03",X"73",X"06",
		X"FD",X"05",X"FF",X"07",X"FF",X"07",X"FF",X"07",X"FD",X"05",X"73",X"06",X"FE",X"03",X"DC",X"01",
		X"D8",X"00",X"00",X"00",X"00",X"00",X"CA",X"1F",X"00",X"00",X"00",X"00",X"F8",X"00",X"DC",X"01",
		X"DE",X"03",X"53",X"06",X"DD",X"05",X"DF",X"07",X"DF",X"07",X"DF",X"07",X"FD",X"05",X"73",X"06",
		X"FE",X"03",X"FC",X"01",X"F8",X"00",X"00",X"00",X"00",X"00",X"82",X"1F",X"00",X"00",X"00",X"00",
		X"F8",X"00",X"FC",X"01",X"FE",X"03",X"73",X"06",X"FD",X"05",X"DF",X"07",X"DF",X"07",X"DF",X"07",
		X"DD",X"05",X"53",X"06",X"DE",X"03",X"DC",X"01",X"F8",X"00",X"00",X"00",X"00",X"00",X"3A",X"2A",
		X"21",X"FE",X"10",X"E2",X"EE",X"1F",X"C3",X"4A",X"07",X"FF",X"85",X"78",X"E9",X"01",X"6C",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
