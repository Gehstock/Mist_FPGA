library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity f1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of f1 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"1C",X"00",X"1C",X"00",X"1C",X"00",
		X"1C",X"00",X"1C",X"00",X"1C",X"00",X"2A",X"00",X"55",X"00",X"55",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"20",X"00",X"20",X"00",X"20",X"00",X"70",X"00",X"70",X"00",X"70",X"00",
		X"70",X"00",X"70",X"00",X"70",X"00",X"A8",X"00",X"54",X"01",X"54",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"C0",X"01",X"C0",X"01",X"C0",X"01",
		X"C0",X"01",X"C0",X"01",X"C0",X"01",X"A0",X"02",X"50",X"05",X"50",X"05",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"07",X"00",X"07",X"00",X"07",
		X"00",X"07",X"00",X"07",X"00",X"07",X"80",X"0A",X"40",X"15",X"40",X"15",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"00",X"1C",X"00",X"3E",X"00",X"1C",X"00",X"08",X"00",X"08",X"00",
		X"08",X"00",X"5D",X"00",X"7F",X"00",X"7F",X"00",X"7F",X"00",X"49",X"00",X"41",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"20",X"00",X"70",X"00",X"F8",X"00",X"70",X"00",X"20",X"00",X"20",X"00",
		X"20",X"00",X"74",X"01",X"FC",X"01",X"FC",X"01",X"FC",X"01",X"24",X"01",X"04",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"00",X"C0",X"01",X"E0",X"03",X"C0",X"01",X"80",X"00",X"80",X"00",
		X"80",X"00",X"D0",X"05",X"F0",X"07",X"F0",X"07",X"F0",X"07",X"90",X"04",X"10",X"04",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"07",X"80",X"0F",X"00",X"07",X"00",X"02",X"00",X"02",
		X"00",X"02",X"40",X"17",X"C0",X"1F",X"C0",X"1F",X"C0",X"1F",X"40",X"12",X"40",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"00",X"1C",X"00",X"3E",X"00",X"2A",X"00",X"2A",X"00",X"2A",X"00",
		X"3E",X"00",X"3E",X"00",X"2A",X"00",X"14",X"00",X"14",X"00",X"22",X"00",X"55",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"20",X"00",X"70",X"00",X"F8",X"00",X"A8",X"00",X"A8",X"00",X"A8",X"00",
		X"F8",X"00",X"F8",X"00",X"A8",X"00",X"50",X"00",X"50",X"00",X"88",X"00",X"54",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"00",X"C0",X"01",X"E0",X"03",X"A0",X"02",X"A0",X"02",X"A0",X"02",
		X"E0",X"03",X"E0",X"03",X"A0",X"02",X"40",X"01",X"40",X"01",X"20",X"02",X"50",X"05",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"07",X"80",X"0F",X"80",X"0A",X"80",X"0A",X"80",X"0A",
		X"80",X"0F",X"80",X"0F",X"80",X"0A",X"00",X"05",X"00",X"05",X"80",X"08",X"40",X"15",X"00",X"00",
		X"03",X"C0",X"00",X"07",X"E0",X"00",X"0D",X"B0",X"00",X"19",X"98",X"00",X"11",X"88",X"00",X"91",
		X"89",X"00",X"D5",X"AB",X"00",X"FD",X"BF",X"00",X"FD",X"BF",X"00",X"D5",X"AB",X"00",X"91",X"89",
		X"00",X"11",X"88",X"00",X"19",X"98",X"00",X"0D",X"B0",X"00",X"07",X"E0",X"00",X"03",X"C0",X"00",
		X"0C",X"00",X"03",X"1C",X"80",X"03",X"34",X"C0",X"02",X"64",X"60",X"02",X"44",X"20",X"02",X"44",
		X"26",X"02",X"54",X"AF",X"02",X"F4",X"FF",X"02",X"F4",X"FF",X"02",X"54",X"AF",X"02",X"44",X"26",
		X"02",X"44",X"20",X"02",X"64",X"60",X"02",X"34",X"C0",X"02",X"1C",X"80",X"03",X"0C",X"00",X"03",
		X"30",X"00",X"0C",X"70",X"00",X"0E",X"D0",X"00",X"0B",X"90",X"81",X"09",X"10",X"81",X"08",X"10",
		X"99",X"08",X"50",X"BD",X"0A",X"D0",X"FF",X"0B",X"D0",X"FF",X"0B",X"50",X"BD",X"0A",X"10",X"99",
		X"08",X"10",X"81",X"08",X"90",X"81",X"09",X"D0",X"00",X"0B",X"70",X"00",X"0E",X"30",X"00",X"0C",
		X"C0",X"00",X"30",X"C0",X"01",X"38",X"40",X"03",X"2C",X"40",X"06",X"26",X"40",X"04",X"22",X"40",
		X"64",X"22",X"40",X"F5",X"2A",X"40",X"FF",X"2F",X"40",X"FF",X"2F",X"40",X"F5",X"2A",X"40",X"64",
		X"22",X"40",X"04",X"22",X"40",X"06",X"26",X"40",X"03",X"2C",X"C0",X"01",X"38",X"C0",X"00",X"30",
		X"00",X"00",X"00",X"72",X"02",X"00",X"15",X"05",X"00",X"34",X"05",X"00",X"42",X"05",X"00",X"41",
		X"05",X"00",X"37",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C8",X"09",X"00",X"54",X"14",
		X"00",X"D0",X"14",X"00",X"08",X"15",X"00",X"04",X"15",X"00",X"DC",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"20",X"27",X"00",X"50",X"51",X"00",X"40",X"53",X"00",X"20",X"54",X"00",X"10",
		X"54",X"00",X"70",X"23",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"9C",X"00",X"40",X"45",
		X"01",X"00",X"4D",X"01",X"80",X"50",X"01",X"40",X"50",X"01",X"C0",X"8D",X"00",X"00",X"00",X"00",
		X"F0",X"0F",X"00",X"FE",X"7F",X"00",X"9F",X"F9",X"00",X"FE",X"7F",X"00",X"F8",X"1F",X"00",X"E0",
		X"07",X"00",X"30",X"0C",X"00",X"18",X"18",X"00",X"C0",X"3F",X"00",X"F8",X"FF",X"01",X"7C",X"E6",
		X"03",X"F8",X"FF",X"01",X"E0",X"7F",X"00",X"80",X"1F",X"00",X"C0",X"30",X"00",X"60",X"60",X"00",
		X"00",X"FF",X"00",X"E0",X"FF",X"07",X"F0",X"99",X"0F",X"E0",X"FF",X"07",X"80",X"FF",X"01",X"00",
		X"7E",X"00",X"00",X"C3",X"00",X"80",X"81",X"01",X"00",X"FC",X"03",X"80",X"FF",X"1F",X"C0",X"67",
		X"3E",X"80",X"FF",X"1F",X"00",X"FE",X"07",X"00",X"F8",X"01",X"00",X"0C",X"03",X"00",X"06",X"06",
		X"02",X"00",X"07",X"00",X"02",X"00",X"07",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"00",X"0E",X"00",X"04",X"00",X"0E",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"00",X"1C",X"00",X"08",X"00",X"1C",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"00",X"38",X"00",X"10",X"00",X"38",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"00",X"70",X"00",X"20",X"00",X"70",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"00",X"E0",X"00",X"40",X"00",X"E0",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"C0",X"01",X"80",X"00",X"C0",X"01",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"80",X"03",X"00",X"01",X"80",X"03",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"00",X"08",X"00",X"1C",X"00",X"1C",X"00",X"1C",X"00",X"14",X"00",
		X"3E",X"00",X"3E",X"00",X"2A",X"00",X"7F",X"00",X"6B",X"00",X"49",X"00",X"55",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"20",X"00",X"20",X"00",X"70",X"00",X"70",X"00",X"70",X"00",X"50",X"00",
		X"F8",X"00",X"F8",X"00",X"A8",X"00",X"FC",X"01",X"AC",X"01",X"24",X"01",X"54",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"00",X"80",X"00",X"C0",X"01",X"C0",X"01",X"C0",X"01",X"40",X"01",
		X"E0",X"03",X"E0",X"03",X"A0",X"02",X"F0",X"07",X"B0",X"06",X"90",X"04",X"50",X"05",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"02",X"00",X"07",X"00",X"07",X"00",X"07",X"00",X"05",
		X"80",X"0F",X"80",X"0F",X"80",X"0A",X"C0",X"1F",X"C0",X"1A",X"40",X"12",X"40",X"15",X"00",X"00",
		X"CD",X"FB",X"15",X"2A",X"74",X"20",X"44",X"4D",X"21",X"68",X"20",X"CD",X"76",X"14",X"C9",X"3A",
		X"12",X"20",X"E6",X"03",X"CA",X"B4",X"16",X"3D",X"CA",X"DE",X"16",X"3D",X"CA",X"08",X"17",X"C3",
		X"32",X"17",X"CD",X"6F",X"18",X"3A",X"12",X"20",X"E6",X"01",X"CA",X"9C",X"18",X"C3",X"C7",X"18",
		X"00",X"00",X"00",X"00",X"00",X"00",X"CD",X"D0",X"14",X"1E",X"10",X"CD",X"2A",X"15",X"C9",X"CD",
		X"D0",X"14",X"1E",X"10",X"CD",X"B7",X"15",X"C9",X"3A",X"12",X"20",X"E6",X"03",X"CA",X"BD",X"19",
		X"3D",X"CA",X"E7",X"19",X"C9",X"C3",X"5E",X"14",X"C3",X"6C",X"14",X"C3",X"93",X"1A",X"3A",X"6B",
		X"20",X"FE",X"50",X"D8",X"3E",X"FF",X"32",X"C9",X"21",X"C3",X"00",X"14",X"AF",X"21",X"C9",X"21",
		X"BE",X"77",X"C0",X"C3",X"00",X"14",X"C5",X"E5",X"E5",X"7D",X"C6",X"13",X"6F",X"7E",X"B7",X"CA",
		X"88",X"14",X"36",X"00",X"23",X"4E",X"23",X"46",X"E1",X"CD",X"F1",X"14",X"1E",X"10",X"CD",X"42",
		X"15",X"E1",X"C1",X"23",X"23",X"E5",X"CD",X"F1",X"14",X"1E",X"10",X"CD",X"CD",X"15",X"E1",X"CD",
		X"F2",X"15",X"C9",X"C5",X"E5",X"E5",X"7D",X"C6",X"13",X"6F",X"7E",X"B7",X"CA",X"B5",X"14",X"36",
		X"00",X"23",X"4E",X"23",X"46",X"E1",X"CD",X"D0",X"14",X"1E",X"10",X"CD",X"2A",X"15",X"E1",X"C1",
		X"23",X"23",X"E5",X"CD",X"D0",X"14",X"1E",X"10",X"CD",X"B7",X"15",X"E1",X"CD",X"F2",X"15",X"C9",
		X"7E",X"07",X"07",X"07",X"07",X"E6",X"60",X"81",X"D2",X"DC",X"14",X"04",X"4F",X"7E",X"0F",X"0F",
		X"0F",X"E6",X"1F",X"5F",X"23",X"6E",X"26",X"00",X"29",X"29",X"29",X"29",X"29",X"16",X"24",X"19",
		X"C9",X"7E",X"E6",X"01",X"32",X"F0",X"21",X"7E",X"0F",X"E6",X"03",X"07",X"07",X"07",X"07",X"5F",
		X"07",X"81",X"D2",X"06",X"15",X"04",X"4F",X"7B",X"81",X"D2",X"0D",X"15",X"04",X"4F",X"C3",X"DD",
		X"14",X"7E",X"E6",X"01",X"32",X"F0",X"21",X"7E",X"0F",X"E6",X"03",X"07",X"07",X"07",X"5F",X"07",
		X"83",X"81",X"D2",X"26",X"15",X"04",X"4F",X"C3",X"DD",X"14",X"0A",X"2F",X"A6",X"77",X"03",X"23",
		X"0A",X"2F",X"A6",X"77",X"03",X"7D",X"C6",X"1F",X"D2",X"3C",X"15",X"24",X"6F",X"1D",X"C2",X"2A",
		X"15",X"C9",X"7B",X"B7",X"C8",X"3A",X"F0",X"21",X"B7",X"C2",X"8F",X"15",X"0A",X"2F",X"A6",X"77",
		X"03",X"23",X"0A",X"2F",X"A6",X"77",X"03",X"23",X"0A",X"2F",X"A6",X"77",X"03",X"7D",X"C6",X"1E",
		X"D2",X"64",X"15",X"24",X"6F",X"1D",X"C2",X"4C",X"15",X"C9",X"0A",X"57",X"B7",X"17",X"B6",X"77",
		X"7A",X"17",X"03",X"23",X"0A",X"57",X"17",X"B6",X"77",X"7A",X"17",X"03",X"23",X"0A",X"17",X"B6",
		X"77",X"03",X"7D",X"C6",X"1E",X"D2",X"89",X"15",X"24",X"6F",X"1D",X"C2",X"6A",X"15",X"C9",X"0A",
		X"2F",X"57",X"37",X"17",X"A6",X"77",X"7A",X"17",X"03",X"23",X"0A",X"2F",X"57",X"17",X"A6",X"77",
		X"7A",X"17",X"03",X"23",X"0A",X"2F",X"17",X"A6",X"77",X"03",X"7D",X"C6",X"1E",X"D2",X"B1",X"15",
		X"24",X"6F",X"1D",X"C2",X"8F",X"15",X"C9",X"0A",X"B6",X"77",X"03",X"23",X"0A",X"B6",X"77",X"03",
		X"7D",X"C6",X"1F",X"D2",X"C7",X"15",X"24",X"6F",X"1D",X"C2",X"B7",X"15",X"C9",X"7B",X"B7",X"C8",
		X"3A",X"F0",X"21",X"B7",X"C2",X"6A",X"15",X"0A",X"B6",X"77",X"03",X"23",X"0A",X"B6",X"77",X"03",
		X"23",X"0A",X"B6",X"77",X"03",X"7D",X"C6",X"1E",X"D2",X"EC",X"15",X"24",X"6F",X"1D",X"C2",X"D7",
		X"15",X"C9",X"5E",X"23",X"56",X"2B",X"2B",X"72",X"2B",X"73",X"C9",X"21",X"6B",X"20",X"3A",X"22",
		X"20",X"B7",X"CA",X"5B",X"14",X"3A",X"90",X"21",X"B7",X"C2",X"13",X"16",X"3A",X"50",X"23",X"B7",
		X"CA",X"19",X"16",X"36",X"C0",X"2B",X"36",X"78",X"C9",X"3A",X"21",X"20",X"96",X"DA",X"61",X"16",
		X"C6",X"0E",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"86",X"77",X"3A",X"72",X"20",X"BE",X"D2",X"32",
		X"16",X"77",X"CD",X"A1",X"16",X"21",X"6A",X"20",X"3A",X"20",X"20",X"96",X"DA",X"57",X"16",X"0F",
		X"0F",X"0F",X"E6",X"1F",X"86",X"77",X"79",X"BE",X"D2",X"4F",X"16",X"CD",X"6C",X"16",X"77",X"78",
		X"BE",X"D8",X"CD",X"6C",X"16",X"77",X"C9",X"0F",X"0F",X"0F",X"F6",X"E0",X"86",X"77",X"C3",X"46",
		X"16",X"0F",X"0F",X"0F",X"0F",X"F6",X"F0",X"86",X"77",X"C3",X"32",X"16",X"F5",X"E5",X"D5",X"21",
		X"A9",X"21",X"36",X"02",X"3A",X"29",X"20",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"FE",X"07",X"DA",
		X"84",X"16",X"3E",X"07",X"11",X"99",X"16",X"83",X"D2",X"8C",X"16",X"14",X"5F",X"23",X"7E",X"B7",
		X"C2",X"95",X"16",X"1A",X"77",X"D1",X"E1",X"F1",X"C9",X"2D",X"2D",X"1E",X"1E",X"0F",X"0F",X"08",
		X"08",X"7E",X"0F",X"0F",X"0F",X"E6",X"1E",X"21",X"9D",X"19",X"85",X"D2",X"AF",X"16",X"24",X"6F",
		X"46",X"23",X"4E",X"C9",X"3A",X"10",X"22",X"B7",X"C8",X"2A",X"0A",X"22",X"44",X"4D",X"21",X"03",
		X"22",X"11",X"09",X"22",X"CD",X"80",X"17",X"EB",X"2B",X"2B",X"CD",X"53",X"18",X"23",X"13",X"CD",
		X"53",X"18",X"2A",X"0C",X"22",X"44",X"4D",X"21",X"00",X"22",X"CD",X"A3",X"14",X"C9",X"3A",X"30",
		X"22",X"B7",X"C8",X"2A",X"2A",X"22",X"44",X"4D",X"21",X"23",X"22",X"11",X"29",X"22",X"CD",X"80",
		X"17",X"EB",X"2B",X"2B",X"CD",X"53",X"18",X"23",X"13",X"CD",X"53",X"18",X"2A",X"2C",X"22",X"44",
		X"4D",X"21",X"20",X"22",X"CD",X"A3",X"14",X"C9",X"3A",X"50",X"22",X"B7",X"C8",X"2A",X"4A",X"22",
		X"44",X"4D",X"21",X"43",X"22",X"11",X"49",X"22",X"CD",X"80",X"17",X"EB",X"2B",X"2B",X"CD",X"53",
		X"18",X"23",X"13",X"CD",X"53",X"18",X"2A",X"4C",X"22",X"44",X"4D",X"21",X"40",X"22",X"CD",X"A3",
		X"14",X"C9",X"3A",X"70",X"22",X"B7",X"C8",X"2A",X"6A",X"22",X"44",X"4D",X"21",X"63",X"22",X"11",
		X"69",X"22",X"CD",X"80",X"17",X"EB",X"2B",X"2B",X"CD",X"53",X"18",X"23",X"13",X"CD",X"53",X"18",
		X"2A",X"6C",X"22",X"44",X"4D",X"21",X"60",X"22",X"CD",X"A3",X"14",X"C9",X"C5",X"7E",X"B8",X"DC",
		X"AD",X"17",X"7E",X"91",X"47",X"DA",X"7E",X"17",X"CD",X"B5",X"17",X"3A",X"D7",X"20",X"B7",X"C2",
		X"7E",X"17",X"78",X"0F",X"0F",X"0F",X"E6",X"1F",X"47",X"7E",X"90",X"77",X"C1",X"C9",X"C1",X"C9",
		X"E5",X"7D",X"C6",X"0E",X"6F",X"7E",X"B7",X"E1",X"C2",X"BD",X"17",X"3A",X"04",X"20",X"B7",X"C2",
		X"BD",X"17",X"CD",X"5C",X"17",X"E5",X"CD",X"A1",X"16",X"E1",X"2B",X"1B",X"1B",X"1B",X"CD",X"A2",
		X"17",X"C9",X"7E",X"B8",X"DC",X"AD",X"17",X"7E",X"B9",X"D4",X"B5",X"17",X"C9",X"1A",X"FE",X"80",
		X"D8",X"2F",X"3C",X"12",X"C9",X"1A",X"FE",X"80",X"D0",X"2F",X"3C",X"12",X"C9",X"CD",X"C3",X"17",
		X"C3",X"95",X"17",X"7E",X"B8",X"DC",X"AD",X"17",X"3A",X"6B",X"20",X"C6",X"18",X"BE",X"D0",X"06",
		X"00",X"70",X"2B",X"70",X"7D",X"C6",X"0E",X"6F",X"70",X"23",X"70",X"2B",X"2B",X"2B",X"2B",X"46",
		X"2B",X"4E",X"E5",X"CD",X"F1",X"17",X"E1",X"7D",X"D6",X"0C",X"6F",X"CD",X"36",X"14",X"C1",X"C1",
		X"C9",X"7D",X"C6",X"07",X"6F",X"AF",X"BE",X"C8",X"77",X"23",X"4E",X"23",X"46",X"C9",X"CD",X"04");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
