library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity satans_hollow_sp_bits_4 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of satans_hollow_sp_bits_4 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"DD",X"00",
		X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"E0",X"7D",X"00",
		X"00",X"D7",X"76",X"00",X"00",X"77",X"76",X"00",X"00",X"E0",X"7D",X"00",X"00",X"E0",X"6D",X"00",
		X"00",X"E0",X"66",X"00",X"00",X"60",X"76",X"00",X"00",X"DD",X"76",X"00",X"DD",X"66",X"76",X"00",
		X"77",X"66",X"76",X"00",X"00",X"77",X"76",X"00",X"00",X"E0",X"76",X"00",X"00",X"E0",X"6D",X"00",
		X"00",X"E0",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"77",X"DD",X"00",X"00",X"77",X"DD",X"00",
		X"00",X"E0",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"DD",X"00",
		X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"E0",X"7D",X"00",
		X"00",X"D7",X"76",X"00",X"06",X"77",X"76",X"00",X"00",X"E0",X"7D",X"00",X"00",X"E0",X"6D",X"00",
		X"00",X"E0",X"66",X"00",X"00",X"60",X"76",X"00",X"DD",X"DD",X"76",X"00",X"00",X"66",X"76",X"00",
		X"00",X"66",X"76",X"00",X"77",X"77",X"76",X"00",X"00",X"E0",X"76",X"00",X"00",X"E0",X"6D",X"00",
		X"00",X"E0",X"DD",X"00",X"00",X"60",X"DD",X"00",X"00",X"77",X"DD",X"00",X"00",X"77",X"DD",X"00",
		X"00",X"E0",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"DD",X"00",
		X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"07",X"E0",X"7D",X"00",
		X"06",X"D7",X"76",X"00",X"06",X"77",X"76",X"00",X"07",X"E0",X"7D",X"00",X"00",X"E0",X"0D",X"00",
		X"00",X"E0",X"66",X"00",X"00",X"60",X"76",X"00",X"00",X"DD",X"76",X"00",X"DD",X"66",X"76",X"00",
		X"77",X"66",X"76",X"00",X"00",X"77",X"76",X"00",X"00",X"E0",X"76",X"00",X"00",X"E0",X"6D",X"00",
		X"00",X"E0",X"DD",X"00",X"00",X"60",X"DD",X"00",X"00",X"77",X"DD",X"00",X"00",X"77",X"DD",X"00",
		X"00",X"E0",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"DD",X"00",
		X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"E0",X"7D",X"00",
		X"DD",X"D7",X"76",X"00",X"77",X"77",X"76",X"00",X"00",X"E0",X"7D",X"00",X"00",X"E0",X"0D",X"00",
		X"00",X"E0",X"66",X"00",X"00",X"60",X"76",X"00",X"0D",X"DD",X"76",X"00",X"00",X"66",X"76",X"00",
		X"00",X"66",X"76",X"00",X"07",X"77",X"76",X"00",X"00",X"E0",X"76",X"00",X"00",X"E0",X"6D",X"00",
		X"00",X"E0",X"DD",X"00",X"00",X"60",X"DD",X"00",X"00",X"77",X"DD",X"00",X"00",X"77",X"DD",X"00",
		X"00",X"E0",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"DD",X"00",
		X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"07",X"E0",X"7D",X"00",
		X"06",X"D7",X"76",X"00",X"06",X"77",X"76",X"00",X"07",X"E0",X"7D",X"00",X"00",X"E0",X"6D",X"00",
		X"00",X"E0",X"66",X"00",X"00",X"60",X"76",X"00",X"00",X"DD",X"76",X"00",X"DD",X"66",X"76",X"00",
		X"77",X"66",X"76",X"00",X"00",X"77",X"76",X"00",X"00",X"E0",X"76",X"00",X"00",X"E0",X"6D",X"00",
		X"00",X"E0",X"DD",X"00",X"07",X"60",X"DD",X"00",X"06",X"77",X"DD",X"00",X"06",X"77",X"DD",X"00",
		X"07",X"E0",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"DD",X"00",
		X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"E0",X"7D",X"00",
		X"DD",X"D7",X"76",X"00",X"77",X"77",X"76",X"00",X"00",X"E0",X"7D",X"00",X"00",X"E0",X"6D",X"00",
		X"00",X"E0",X"66",X"00",X"00",X"60",X"76",X"00",X"0D",X"DD",X"76",X"00",X"00",X"66",X"76",X"00",
		X"00",X"66",X"76",X"00",X"07",X"77",X"76",X"00",X"00",X"E0",X"76",X"00",X"00",X"E0",X"6D",X"00",
		X"00",X"E0",X"DD",X"00",X"00",X"60",X"DD",X"00",X"DD",X"77",X"DD",X"00",X"77",X"77",X"DD",X"00",
		X"00",X"E0",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"31",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"10",
		X"10",X"10",X"11",X"31",X"F1",X"21",X"44",X"11",X"5F",X"22",X"34",X"23",X"51",X"42",X"22",X"11",
		X"1C",X"44",X"11",X"31",X"16",X"22",X"31",X"10",X"33",X"22",X"41",X"00",X"16",X"22",X"41",X"00",
		X"1C",X"22",X"31",X"00",X"51",X"44",X"11",X"00",X"5F",X"42",X"22",X"00",X"F1",X"22",X"24",X"00",
		X"11",X"21",X"33",X"10",X"00",X"10",X"11",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"14",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"23",X"00",X"00",X"00",
		X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"9F",X"00",X"00",X"00",X"99",X"00",
		X"00",X"99",X"90",X"00",X"00",X"CC",X"09",X"F0",X"00",X"99",X"09",X"F0",X"00",X"00",X"09",X"F0",
		X"00",X"0F",X"00",X"F0",X"00",X"FC",X"90",X"F0",X"00",X"CC",X"90",X"F0",X"00",X"CC",X"C9",X"F0",
		X"00",X"C9",X"09",X"F0",X"00",X"C9",X"99",X"F0",X"00",X"FC",X"99",X"F0",X"00",X"CC",X"FF",X"F0",
		X"00",X"CF",X"F9",X"F0",X"00",X"0F",X"99",X"F0",X"00",X"0F",X"9C",X"F0",X"00",X"00",X"09",X"F0",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"90",X"F0",X"00",X"FF",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"00",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"CC",X"FF",X"00",X"00",X"99",X"F0",X"00",
		X"00",X"00",X"F0",X"00",X"09",X"FF",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"90",X"90",X"00",X"00",X"00",X"90",X"00",
		X"00",X"90",X"00",X"90",X"00",X"00",X"00",X"90",X"99",X"00",X"00",X"90",X"99",X"99",X"90",X"90",
		X"69",X"99",X"90",X"90",X"69",X"99",X"99",X"00",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"00",
		X"69",X"99",X"99",X"00",X"69",X"99",X"99",X"90",X"99",X"99",X"99",X"00",X"99",X"99",X"90",X"99",
		X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"09",X"00",X"09",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"0C",X"CC",X"00",
		X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",
		X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",
		X"00",X"CC",X"CC",X"00",X"00",X"CC",X"C0",X"00",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"99",X"90",X"00",
		X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"F9",X"66",X"00",
		X"90",X"F9",X"C6",X"00",X"59",X"F9",X"CC",X"00",X"50",X"59",X"CC",X"00",X"55",X"55",X"CC",X"00",
		X"55",X"66",X"CC",X"00",X"95",X"66",X"CC",X"00",X"00",X"CC",X"6C",X"00",X"00",X"CC",X"CC",X"00",
		X"09",X"CC",X"CC",X"00",X"09",X"C6",X"CC",X"00",X"00",X"C6",X"CC",X"00",X"00",X"6C",X"CC",X"00",
		X"00",X"CC",X"CC",X"00",X"00",X"CC",X"66",X"00",X"00",X"CC",X"00",X"00",X"00",X"6C",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",
		X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",
		X"BB",X"BB",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"90",X"00",X"00",X"DD",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"90",X"00",X"00",X"DD",X"00",X"00",X"00",
		X"00",X"90",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"02",X"00",X"00",
		X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"29",X"00",
		X"00",X"00",X"22",X"00",X"90",X"00",X"22",X"40",X"49",X"00",X"99",X"00",X"90",X"99",X"99",X"00",
		X"00",X"22",X"99",X"00",X"00",X"02",X"99",X"00",X"00",X"00",X"22",X"40",X"00",X"00",X"22",X"00",
		X"00",X"00",X"22",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",
		X"00",X"02",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"20",X"00",X"00",
		X"99",X"B0",X"00",X"00",X"BB",X"BB",X"00",X"00",X"B1",X"11",X"00",X"00",X"9A",X"91",X"00",X"00",
		X"1B",X"9B",X"00",X"00",X"B1",X"B9",X"B0",X"00",X"B1",X"BB",X"1B",X"00",X"91",X"B9",X"B1",X"00",
		X"91",X"BB",X"11",X"00",X"B1",X"B9",X"BB",X"00",X"B9",X"BB",X"B9",X"00",X"BB",X"BB",X"B9",X"00",
		X"BB",X"11",X"B9",X"00",X"BB",X"11",X"B9",X"B0",X"BB",X"99",X"19",X"BB",X"BB",X"BB",X"19",X"BB",
		X"BB",X"BB",X"B9",X"B0",X"BB",X"BB",X"B9",X"00",X"BB",X"BB",X"B9",X"00",X"BB",X"BB",X"B9",X"00",
		X"B9",X"BB",X"BB",X"00",X"B9",X"BB",X"BB",X"00",X"91",X"BB",X"BB",X"00",X"91",X"BB",X"BB",X"00",
		X"91",X"B9",X"B0",X"00",X"B1",X"91",X"00",X"00",X"A1",X"91",X"00",X"00",X"1B",X"1B",X"00",X"00",
		X"BB",X"BB",X"00",X"00",X"BB",X"00",X"00",X"00",X"B9",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"B0",
		X"00",X"00",X"0B",X"B0",X"00",X"00",X"BB",X"B0",X"00",X"00",X"BB",X"00",X"F0",X"00",X"B9",X"00",
		X"7F",X"00",X"BB",X"00",X"0F",X"00",X"BB",X"00",X"0F",X"00",X"1B",X"00",X"0F",X"00",X"90",X"00",
		X"07",X"09",X"99",X"00",X"97",X"77",X"99",X"00",X"FF",X"FF",X"99",X"00",X"07",X"00",X"90",X"00",
		X"07",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"7F",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"BB",X"99",X"00",X"99",X"BB",X"11",X"00",X"99",X"B9",X"11",X"00",X"99",X"99",X"BB",
		X"00",X"09",X"91",X"BB",X"00",X"09",X"91",X"BB",X"00",X"00",X"91",X"BB",X"00",X"00",X"91",X"BB",
		X"00",X"00",X"91",X"BB",X"00",X"0A",X"11",X"B9",X"00",X"C0",X"11",X"B9",X"00",X"00",X"B1",X"91",
		X"00",X"00",X"B9",X"9B",X"00",X"00",X"BB",X"90",X"00",X"09",X"90",X"00",X"00",X"91",X"99",X"00",
		X"00",X"11",X"09",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"19",X"BB",X"00",X"00",X"B9",X"BB",X"00",X"00",X"B9",X"B0",X"00",X"00",X"B9",X"00",X"00",X"00",
		X"19",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",
		X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"8F",X"C8",X"88",X"88",X"F9",X"9C",
		X"88",X"88",X"99",X"C8",X"88",X"88",X"89",X"98",X"88",X"88",X"F8",X"C8",X"88",X"88",X"9F",X"98",
		X"88",X"88",X"99",X"C8",X"88",X"88",X"99",X"C8",X"88",X"88",X"97",X"C1",X"88",X"88",X"77",X"18",
		X"88",X"88",X"79",X"C8",X"88",X"88",X"79",X"C8",X"88",X"9F",X"99",X"CC",X"88",X"F9",X"99",X"CC",
		X"88",X"8F",X"89",X"C8",X"88",X"88",X"89",X"98",X"88",X"88",X"99",X"98",X"88",X"88",X"97",X"C8",
		X"88",X"88",X"99",X"C8",X"88",X"88",X"F9",X"98",X"88",X"88",X"89",X"98",X"88",X"88",X"99",X"98",
		X"88",X"88",X"99",X"98",X"88",X"88",X"79",X"98",X"88",X"88",X"99",X"94",X"88",X"88",X"FF",X"98",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"00",X"BB",X"BB",X"99",X"00",X"BB",X"9B",X"11",X"00",X"BB",X"B9",X"11",X"00",X"BB",X"99",X"BB",
		X"00",X"BB",X"99",X"BB",X"00",X"BB",X"91",X"BB",X"00",X"BB",X"91",X"BB",X"00",X"BA",X"1A",X"BB",
		X"00",X"AA",X"1C",X"BB",X"00",X"AA",X"1C",X"BB",X"00",X"AA",X"CC",X"B9",X"00",X"AB",X"CC",X"99",
		X"00",X"BB",X"C9",X"9B",X"00",X"BB",X"BB",X"99",X"00",X"BB",X"BB",X"91",X"00",X"9B",X"99",X"11",
		X"00",X"1B",X"09",X"11",X"00",X"9B",X"00",X"11",X"00",X"B1",X"00",X"19",X"00",X"11",X"00",X"90",
		X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"91",X"BB",X"B0",X"00",X"1B",X"BB",X"B0",X"00",X"1B",X"B1",X"00",X"00",X"BB",X"B1",X"00",X"00",
		X"1B",X"11",X"00",X"00",X"BB",X"11",X"00",X"00",X"1B",X"11",X"00",X"00",X"B1",X"19",X"00",X"00",
		X"11",X"11",X"00",X"00",X"91",X"00",X"00",X"00",X"1B",X"00",X"00",X"00",X"B1",X"00",X"00",X"00",
		X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"FD",X"00",X"00",X"00",X"FD",X"00",X"00",
		X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"E0",X"00",
		X"00",X"DD",X"E0",X"00",X"00",X"DD",X"E0",X"00",X"00",X"DE",X"E0",X"00",X"00",X"DD",X"E0",X"00",
		X"00",X"DD",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",
		X"00",X"00",X"23",X"00",X"00",X"00",X"32",X"00",X"00",X"33",X"32",X"00",X"00",X"39",X"33",X"00",
		X"00",X"33",X"23",X"00",X"00",X"00",X"22",X"40",X"00",X"00",X"33",X"00",X"00",X"33",X"33",X"00",
		X"00",X"33",X"33",X"00",X"00",X"22",X"32",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"33",X"00",
		X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"30",X"00",X"00",X"02",X"00",X"00",
		X"00",X"02",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"23",X"00",X"00",X"00",X"23",X"00",X"00",
		X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"55",X"00",X"00",X"CC",X"55",X"00",
		X"99",X"CC",X"00",X"00",X"99",X"CC",X"00",X"00",X"99",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"C5",X"00",X"00",
		X"00",X"C5",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"CC",X"C5",X"00",X"00",X"CC",X"C5",X"00",
		X"99",X"CC",X"05",X"00",X"99",X"CC",X"00",X"00",X"00",X"5C",X"00",X"00",X"00",X"55",X"50",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"CC",X"00",X"00",X"99",X"CC",X"00",X"99",X"99",X"55",X"00",X"99",X"99",X"55",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"CC",X"99",X"CC",X"00",X"CC",X"99",X"CC",X"00",
		X"55",X"CC",X"55",X"00",X"55",X"CC",X"55",X"00",X"99",X"9C",X"99",X"00",X"99",X"CC",X"99",X"00",
		X"00",X"CC",X"CC",X"99",X"00",X"99",X"CC",X"99",X"00",X"99",X"55",X"00",X"00",X"99",X"55",X"00",
		X"CC",X"99",X"99",X"00",X"CC",X"99",X"99",X"00",X"CC",X"99",X"CC",X"00",X"CC",X"99",X"CC",X"00",
		X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"55",X"00",X"00",X"CC",X"55",X"00",X"00",X"CC",
		X"99",X"CC",X"00",X"CC",X"99",X"CC",X"00",X"CC",X"55",X"55",X"CC",X"00",X"55",X"55",X"CC",X"00",
		X"CC",X"99",X"55",X"00",X"CC",X"99",X"55",X"00",X"CC",X"99",X"99",X"00",X"CC",X"99",X"59",X"00",
		X"55",X"FF",X"99",X"00",X"55",X"F9",X"99",X"00",X"55",X"FF",X"99",X"00",X"55",X"FF",X"99",X"00",
		X"99",X"FF",X"55",X"CC",X"99",X"9F",X"55",X"CC",X"99",X"99",X"55",X"00",X"99",X"99",X"55",X"00",
		X"55",X"99",X"55",X"00",X"55",X"99",X"55",X"00",X"CC",X"99",X"99",X"00",X"CC",X"99",X"99",X"00",
		X"CC",X"55",X"99",X"CC",X"CC",X"55",X"99",X"CC",X"55",X"CC",X"55",X"00",X"55",X"CC",X"55",X"00",
		X"55",X"00",X"CC",X"00",X"55",X"00",X"CC",X"00",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"90",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"99",X"00",X"00",X"99",X"99",
		X"99",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",X"99",X"00",X"99",X"99",X"C9",X"99",X"99",X"99",
		X"C9",X"99",X"F9",X"00",X"CC",X"FF",X"CC",X"00",X"CC",X"99",X"9C",X"CC",X"CC",X"9C",X"99",X"9C",
		X"CC",X"99",X"99",X"99",X"99",X"C9",X"FF",X"99",X"FC",X"CC",X"99",X"99",X"FF",X"FF",X"C9",X"00",
		X"9F",X"CC",X"99",X"00",X"9F",X"CC",X"99",X"00",X"9F",X"FF",X"99",X"00",X"99",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"90",X"00",X"90",
		X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"99",X"00",X"09",
		X"00",X"90",X"00",X"99",X"09",X"00",X"00",X"09",X"09",X"00",X"00",X"09",X"99",X"99",X"00",X"99",
		X"99",X"99",X"00",X"00",X"9F",X"FF",X"99",X"00",X"9F",X"CC",X"99",X"00",X"9F",X"99",X"99",X"00",
		X"FF",X"9F",X"C9",X"00",X"FC",X"9C",X"99",X"99",X"99",X"C9",X"FF",X"99",X"9C",X"99",X"99",X"99",
		X"9C",X"9C",X"99",X"9C",X"CC",X"99",X"9C",X"CC",X"CC",X"F9",X"CC",X"00",X"C9",X"99",X"F9",X"00",
		X"99",X"99",X"99",X"99",X"99",X"00",X"99",X"99",X"F9",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"99",X"00",X"90",X"00",X"99",
		X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",
		X"99",X"99",X"90",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"00",X"99",X"99",X"00",
		X"90",X"00",X"C9",X"90",X"99",X"00",X"C9",X"90",X"00",X"C0",X"CC",X"00",X"00",X"9C",X"99",X"00",
		X"90",X"99",X"99",X"00",X"90",X"99",X"99",X"00",X"90",X"CC",X"09",X"00",X"90",X"0C",X"09",X"00",
		X"90",X"00",X"09",X"00",X"90",X"00",X"09",X"FF",X"90",X"00",X"09",X"0F",X"00",X"00",X"00",X"0F",
		X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",X"90",X"F0",
		X"00",X"00",X"90",X"F0",X"00",X"00",X"99",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",X"CF",X"00",
		X"00",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"30",X"00",X"00",X"00",X"23",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"02",X"00",X"00",
		X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",
		X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"23",X"00",
		X"00",X"00",X"22",X"00",X"30",X"00",X"22",X"40",X"43",X"00",X"33",X"00",X"20",X"33",X"33",X"00",
		X"00",X"22",X"33",X"00",X"00",X"02",X"33",X"00",X"00",X"00",X"22",X"40",X"00",X"00",X"22",X"00",
		X"00",X"00",X"22",X"00",X"00",X"00",X"23",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",
		X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",
		X"00",X"02",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"23",X"00",X"00",X"00",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"99",X"30",X"00",
		X"00",X"30",X"30",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"23",X"00",X"00",X"00",X"23",X"00",
		X"00",X"00",X"23",X"00",X"00",X"22",X"23",X"00",X"00",X"33",X"23",X"00",X"00",X"33",X"33",X"00",
		X"00",X"03",X"33",X"00",X"00",X"00",X"23",X"00",X"00",X"02",X"22",X"00",X"00",X"22",X"32",X"00",
		X"00",X"33",X"32",X"00",X"22",X"33",X"33",X"00",X"23",X"22",X"00",X"00",X"33",X"33",X"00",X"00",
		X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",
		X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"40",X"20",X"00",X"00",X"93",X"20",X"00",
		X"00",X"13",X"30",X"00",X"00",X"93",X"33",X"00",X"00",X"40",X"33",X"00",X"00",X"00",X"33",X"00",
		X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",
		X"00",X"20",X"23",X"00",X"00",X"32",X"23",X"00",X"00",X"33",X"23",X"00",X"22",X"03",X"23",X"00",
		X"32",X"00",X"33",X"00",X"33",X"00",X"23",X"00",X"03",X"22",X"23",X"00",X"00",X"33",X"23",X"00",
		X"00",X"33",X"23",X"00",X"00",X"23",X"32",X"00",X"00",X"32",X"33",X"00",X"00",X"33",X"03",X"00",
		X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"03",X"34",X"00",
		X"00",X"03",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"03",X"00",X"00",
		X"00",X"03",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"23",X"00",X"00",X"00",X"23",X"00",X"00",
		X"00",X"23",X"00",X"00",X"00",X"23",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"32",X"00",X"00",
		X"00",X"32",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"03",X"30",X"00",
		X"00",X"60",X"30",X"00",X"00",X"60",X"30",X"00",X"00",X"66",X"30",X"00",X"00",X"66",X"30",X"00",
		X"00",X"60",X"30",X"00",X"00",X"60",X"30",X"00",X"00",X"60",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"99",X"00",X"00",X"03",X"30",X"00",
		X"00",X"33",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",
		X"00",X"30",X"00",X"00",X"00",X"32",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"03",X"00",X"00",
		X"00",X"03",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"33",X"00",X"00",
		X"00",X"23",X"00",X"00",X"00",X"23",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"32",X"00",X"00",
		X"00",X"32",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",
		X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"23",X"00",X"00",X"00",X"03",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"93",X"00",X"00",X"00",X"13",X"00",
		X"00",X"00",X"93",X"00",X"00",X"00",X"40",X"00",X"00",X"03",X"00",X"00",X"00",X"03",X"00",X"00",
		X"00",X"03",X"02",X"00",X"00",X"03",X"23",X"00",X"00",X"03",X"30",X"00",X"00",X"03",X"30",X"00",
		X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",
		X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"60",X"00",X"00",X"33",X"60",X"00",
		X"00",X"32",X"60",X"00",X"00",X"32",X"60",X"00",X"00",X"22",X"60",X"00",X"00",X"23",X"00",X"00",
		X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"36",X"00",X"00",X"00",X"30",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"03",X"00",X"00",X"00",
		X"03",X"03",X"00",X"00",X"03",X"33",X"00",X"00",X"03",X"32",X"00",X"00",X"33",X"32",X"00",X"00",
		X"33",X"22",X"22",X"00",X"33",X"20",X"33",X"00",X"33",X"22",X"33",X"00",X"33",X"22",X"33",X"00",
		X"33",X"33",X"30",X"00",X"33",X"23",X"00",X"00",X"33",X"22",X"00",X"00",X"33",X"22",X"00",X"00",
		X"30",X"23",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",
		X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"34",X"00",
		X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",
		X"03",X"00",X"00",X"00",X"33",X"03",X"00",X"00",X"33",X"33",X"00",X"00",X"33",X"33",X"00",X"00",
		X"33",X"32",X"00",X"00",X"33",X"32",X"00",X"00",X"33",X"22",X"00",X"00",X"33",X"23",X"00",X"00",
		X"22",X"33",X"20",X"00",X"33",X"22",X"22",X"00",X"00",X"22",X"33",X"00",X"00",X"23",X"33",X"00",
		X"00",X"33",X"33",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",
		X"00",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"D0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"0D",X"D0",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"00",X"00",X"0D",X"D0",X"00",X"00",X"D0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"0D",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"CF",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"F0",
		X"00",X"00",X"90",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"9F",
		X"00",X"00",X"00",X"0F",X"90",X"00",X"09",X"0F",X"90",X"00",X"09",X"FF",X"90",X"00",X"09",X"00",
		X"90",X"09",X"09",X"00",X"90",X"99",X"09",X"00",X"90",X"99",X"99",X"00",X"90",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"90",X"C9",X"00",X"99",X"00",X"C9",X"90",X"90",X"00",X"99",X"90",
		X"00",X"99",X"99",X"00",X"99",X"F0",X"90",X"00",X"9F",X"00",X"00",X"00",X"09",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",
		X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",
		X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"88",X"00",X"00",X"88",X"88",X"00",X"00",
		X"88",X"88",X"00",X"00",X"88",X"88",X"00",X"00",X"88",X"88",X"00",X"00",X"88",X"88",X"80",X"00",
		X"88",X"88",X"88",X"00",X"88",X"88",X"88",X"00",X"88",X"88",X"88",X"00",X"88",X"88",X"88",X"00",
		X"88",X"89",X"88",X"00",X"88",X"C8",X"88",X"00",X"8C",X"5C",X"88",X"00",X"99",X"99",X"88",X"88",
		X"CC",X"C9",X"88",X"88",X"89",X"55",X"98",X"00",X"88",X"88",X"88",X"00",X"8C",X"88",X"88",X"00",
		X"88",X"88",X"88",X"00",X"88",X"88",X"88",X"00",X"88",X"C8",X"88",X"00",X"88",X"88",X"88",X"00",
		X"88",X"88",X"80",X"00",X"88",X"88",X"00",X"00",X"88",X"88",X"00",X"00",X"88",X"88",X"00",X"00",
		X"88",X"88",X"00",X"00",X"08",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"90",X"90",X"00",X"00",X"00",X"90",X"00",
		X"00",X"90",X"00",X"90",X"00",X"00",X"00",X"90",X"99",X"00",X"00",X"90",X"99",X"99",X"90",X"90",
		X"69",X"99",X"90",X"90",X"69",X"99",X"99",X"00",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"00",
		X"69",X"99",X"99",X"00",X"69",X"99",X"99",X"90",X"99",X"99",X"99",X"00",X"99",X"99",X"90",X"99",
		X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"09",X"00",X"90",X"0D",X"00",
		X"00",X"90",X"D0",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"00",X"D0",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"00",X"00",X"00",X"D0",X"00",X"00",X"0D",X"00",
		X"00",X"00",X"D0",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"C9",X"00",X"00",X"00",X"CC",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"F9",X"00",X"00",
		X"00",X"9C",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"9C",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"C0",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"99",X"C0",X"00",
		X"00",X"99",X"90",X"00",X"00",X"99",X"C0",X"00",X"00",X"99",X"90",X"00",X"00",X"F9",X"00",X"00",
		X"00",X"9C",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"C9",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"9C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",
		X"55",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"50",X"00",X"00",
		X"FF",X"55",X"00",X"00",X"5F",X"F5",X"00",X"00",X"5F",X"FF",X"00",X"00",X"5F",X"FF",X"00",X"00",
		X"5F",X"5F",X"00",X"00",X"55",X"55",X"00",X"00",X"05",X"05",X"00",X"00",X"05",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"99",X"90",X"00",
		X"00",X"30",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",
		X"00",X"00",X"29",X"00",X"00",X"22",X"29",X"00",X"00",X"99",X"29",X"00",X"00",X"99",X"99",X"00",
		X"00",X"09",X"99",X"00",X"00",X"00",X"29",X"00",X"00",X"02",X"22",X"00",X"00",X"22",X"92",X"00",
		X"00",X"99",X"92",X"00",X"22",X"99",X"99",X"00",X"29",X"22",X"00",X"00",X"99",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"FF",X"00",X"00",X"EE",X"FF",
		X"00",X"00",X"E0",X"FF",X"00",X"00",X"E0",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"0F",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"FE",X"FF",X"00",X"00",X"EE",X"FF",X"99",X"99",X"0E",X"FF",X"00",X"00",X"EE",X"FF",
		X"00",X"00",X"EE",X"FF",X"00",X"00",X"F0",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"0F",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"E0",X"FF",X"00",X"00",X"EE",X"FF",X"00",X"00",X"0E",X"FF",
		X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"40",X"20",X"00",X"00",X"93",X"20",X"00",
		X"00",X"13",X"90",X"00",X"00",X"93",X"99",X"00",X"00",X"40",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"20",X"29",X"00",X"00",X"92",X"29",X"00",X"00",X"99",X"29",X"00",X"22",X"09",X"29",X"00",
		X"92",X"00",X"99",X"00",X"99",X"00",X"29",X"00",X"09",X"22",X"29",X"00",X"00",X"99",X"29",X"00",
		X"00",X"99",X"29",X"00",X"00",X"29",X"92",X"00",X"00",X"92",X"99",X"00",X"00",X"99",X"09",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"09",X"94",X"00",
		X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",
		X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"92",X"00",X"00",
		X"00",X"92",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"90",X"00",
		X"00",X"60",X"90",X"00",X"00",X"60",X"90",X"00",X"00",X"66",X"90",X"00",X"00",X"66",X"90",X"00",
		X"00",X"60",X"90",X"00",X"00",X"60",X"90",X"00",X"00",X"60",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"30",X"00",
		X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",
		X"00",X"90",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"92",X"00",X"00",
		X"00",X"92",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"93",X"00",X"00",X"00",X"13",X"00",
		X"00",X"00",X"93",X"00",X"00",X"00",X"40",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"09",X"02",X"00",X"00",X"09",X"29",X"00",X"00",X"09",X"90",X"00",X"00",X"09",X"90",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"60",X"00",X"00",X"99",X"60",X"00",
		X"00",X"92",X"60",X"00",X"00",X"92",X"60",X"00",X"00",X"22",X"60",X"00",X"00",X"29",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"96",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",
		X"09",X"09",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"92",X"00",X"00",X"99",X"92",X"00",X"00",
		X"99",X"22",X"22",X"00",X"99",X"20",X"99",X"00",X"99",X"22",X"99",X"00",X"99",X"22",X"99",X"00",
		X"99",X"99",X"90",X"00",X"99",X"29",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"22",X"00",X"00",
		X"90",X"29",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"94",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",
		X"09",X"00",X"00",X"00",X"99",X"09",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"92",X"00",X"00",X"99",X"92",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"29",X"00",X"00",
		X"22",X"99",X"20",X"00",X"99",X"22",X"22",X"00",X"00",X"22",X"99",X"00",X"00",X"29",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
