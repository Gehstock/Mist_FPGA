library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity cclimber_tile_bit1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of cclimber_tile_bit1 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"1C",X"26",X"63",X"63",X"63",X"32",X"1C",X"00",X"0C",X"1C",X"0C",X"0C",X"0C",X"0C",X"3F",X"00",
		X"3E",X"63",X"07",X"1E",X"3C",X"70",X"7F",X"00",X"3F",X"06",X"0C",X"1E",X"03",X"63",X"3E",X"00",
		X"0E",X"1E",X"36",X"66",X"7F",X"06",X"06",X"00",X"3E",X"30",X"3E",X"03",X"03",X"33",X"1E",X"00",
		X"1E",X"30",X"60",X"7E",X"63",X"63",X"3E",X"00",X"3F",X"23",X"06",X"0C",X"18",X"18",X"18",X"00",
		X"3C",X"62",X"72",X"3C",X"4F",X"43",X"3E",X"00",X"3E",X"63",X"63",X"3F",X"03",X"06",X"3C",X"00",
		X"1C",X"36",X"63",X"63",X"7F",X"63",X"63",X"00",X"7E",X"63",X"63",X"7E",X"63",X"63",X"7E",X"00",
		X"1E",X"33",X"60",X"60",X"60",X"33",X"1E",X"00",X"7C",X"66",X"63",X"63",X"63",X"66",X"7C",X"00",
		X"3F",X"30",X"30",X"3E",X"30",X"30",X"3F",X"00",X"7F",X"60",X"60",X"7E",X"60",X"60",X"60",X"00",
		X"1F",X"30",X"60",X"67",X"63",X"33",X"1F",X"00",X"63",X"63",X"63",X"7F",X"63",X"63",X"63",X"00",
		X"3F",X"0C",X"0C",X"0C",X"0C",X"0C",X"3F",X"00",X"03",X"03",X"03",X"03",X"03",X"63",X"3E",X"00",
		X"63",X"66",X"6C",X"78",X"7C",X"6E",X"67",X"00",X"30",X"30",X"30",X"30",X"30",X"30",X"3F",X"00",
		X"63",X"77",X"7F",X"7F",X"6B",X"63",X"63",X"00",X"63",X"73",X"7B",X"7F",X"6F",X"67",X"63",X"00",
		X"3E",X"63",X"63",X"63",X"63",X"63",X"3E",X"00",X"7E",X"63",X"63",X"63",X"7E",X"60",X"60",X"00",
		X"3E",X"63",X"63",X"63",X"6F",X"66",X"3D",X"00",X"7E",X"63",X"63",X"67",X"7C",X"6E",X"67",X"00",
		X"3C",X"66",X"60",X"3E",X"03",X"63",X"3E",X"00",X"3F",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"00",
		X"63",X"63",X"63",X"63",X"63",X"63",X"3E",X"00",X"63",X"63",X"63",X"77",X"3E",X"1C",X"08",X"00",
		X"63",X"63",X"6B",X"7F",X"7F",X"36",X"22",X"00",X"63",X"77",X"3E",X"1C",X"3E",X"77",X"63",X"00",
		X"33",X"33",X"12",X"1E",X"0C",X"0C",X"0C",X"00",X"7F",X"07",X"0E",X"1C",X"38",X"70",X"7F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"06",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",
		X"00",X"00",X"00",X"18",X"1C",X"04",X"08",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"07",X"07",X"07",X"07",X"03",X"03",X"07",X"01",X"80",X"80",X"80",X"80",X"80",X"C0",X"C0",X"E0",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"A0",X"D0",X"C8",X"00",X"00",X"00",X"00",
		X"04",X"02",X"03",X"01",X"01",X"01",X"01",X"03",X"00",X"00",X"00",X"80",X"C0",X"C0",X"C0",X"C0",
		X"03",X"03",X"0B",X"0D",X"07",X"03",X"03",X"03",X"80",X"00",X"00",X"00",X"C0",X"C0",X"E0",X"A0",
		X"0F",X"0F",X"0B",X"03",X"03",X"01",X"01",X"00",X"00",X"80",X"80",X"D0",X"D0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"7C",X"6E",X"2C",X"20",X"10",X"00",X"00",
		X"20",X"60",X"60",X"C0",X"E0",X"E0",X"E0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"80",X"80",X"90",X"50",X"78",X"38",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"09",X"07",X"1E",X"11",X"07",X"14",X"23",X"60",X"C0",X"20",X"70",X"90",X"70",X"C8",X"F8",
		X"04",X"03",X"C0",X"01",X"00",X"01",X"00",X"00",X"24",X"E4",X"02",X"A0",X"00",X"40",X"00",X"00",
		X"00",X"00",X"10",X"18",X"06",X"0A",X"24",X"0B",X"00",X"00",X"00",X"00",X"40",X"68",X"B8",X"C4",
		X"04",X"03",X"24",X"23",X"04",X"03",X"4C",X"43",X"68",X"84",X"60",X"80",X"40",X"80",X"40",X"80",
		X"01",X"22",X"21",X"07",X"04",X"83",X"81",X"00",X"10",X"E0",X"90",X"70",X"C0",X"BA",X"65",X"DA",
		X"01",X"05",X"05",X"02",X"04",X"02",X"00",X"00",X"B0",X"74",X"68",X"88",X"34",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"C4",X"B2",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",
		X"18",X"B7",X"8C",X"1B",X"06",X"4D",X"43",X"06",X"40",X"10",X"20",X"80",X"00",X"C0",X"00",X"E0",
		X"17",X"17",X"07",X"03",X"03",X"07",X"07",X"0F",X"E0",X"E0",X"E0",X"C0",X"C0",X"F8",X"F0",X"E0",
		X"0F",X"0A",X"09",X"00",X"00",X"00",X"00",X"00",X"F0",X"A0",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"01",X"03",X"03",X"01",X"01",X"03",X"03",X"03",X"00",X"80",X"80",X"C0",X"C0",X"C0",X"80",X"80",
		X"03",X"03",X"03",X"03",X"07",X"0F",X"1F",X"1F",X"80",X"00",X"00",X"D0",X"F0",X"E0",X"C0",X"C0",
		X"1F",X"0F",X"07",X"07",X"03",X"03",X"01",X"05",X"E0",X"C0",X"E0",X"F0",X"F0",X"FC",X"FF",X"F9",
		X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7C",X"FE",X"54",X"38",X"00",X"00",X"00",X"00",
		X"20",X"60",X"C0",X"E0",X"F0",X"F0",X"E0",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"60",X"70",X"30",X"36",X"3F",X"BE",X"FF",X"FF",X"00",X"00",X"00",X"00",X"80",X"40",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"7F",X"3F",X"5F",X"1F",X"0F",X"87",X"11",
		X"FC",X"F8",X"F1",X"E3",X"C7",X"CF",X"FF",X"FF",X"FC",X"FE",X"FF",X"F7",X"EE",X"FC",X"F1",X"88",
		X"F1",X"E3",X"C7",X"CF",X"7F",X"7F",X"3F",X"07",X"FF",X"FE",X"FE",X"F8",X"F8",X"E0",X"E3",X"E3",
		X"8F",X"0F",X"3F",X"3F",X"FE",X"FF",X"FF",X"FF",X"FE",X"DF",X"BF",X"7F",X"FE",X"FE",X"FC",X"FC",
		X"1C",X"3F",X"3F",X"7F",X"7F",X"FE",X"FC",X"F8",X"00",X"87",X"FF",X"FF",X"3B",X"3D",X"7F",X"FF",
		X"FC",X"FF",X"FF",X"F8",X"F8",X"E0",X"E3",X"83",X"01",X"88",X"E0",X"FC",X"FE",X"FC",X"F8",X"FC",
		X"0E",X"1F",X"7B",X"77",X"EF",X"DE",X"7C",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"7F",X"3F",X"5F",X"1F",X"0F",X"87",X"11",
		X"FC",X"F8",X"F1",X"E3",X"C7",X"CF",X"FF",X"FF",X"FC",X"FE",X"FF",X"F7",X"EE",X"FC",X"F1",X"88",
		X"F1",X"E3",X"C7",X"CF",X"7F",X"7F",X"3F",X"07",X"FF",X"FE",X"FE",X"F8",X"F8",X"E0",X"E3",X"E3",
		X"8F",X"0F",X"3F",X"3F",X"FE",X"FF",X"FF",X"FF",X"FE",X"DF",X"BF",X"7F",X"FE",X"FE",X"FC",X"FC",
		X"1C",X"3F",X"3F",X"7F",X"7F",X"FE",X"FC",X"F8",X"00",X"87",X"FF",X"FF",X"3B",X"3D",X"7F",X"FF",
		X"FC",X"FF",X"FF",X"F8",X"F8",X"E0",X"E3",X"83",X"01",X"88",X"E0",X"FC",X"FE",X"FC",X"F8",X"FC",
		X"0E",X"1F",X"7B",X"77",X"EF",X"DE",X"7C",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"7F",X"3F",X"5F",X"1F",X"0F",X"87",X"11",
		X"FC",X"F8",X"F1",X"E3",X"C7",X"CF",X"FF",X"FF",X"FC",X"FE",X"FF",X"F7",X"EE",X"FC",X"F1",X"88",
		X"F1",X"E3",X"C7",X"CF",X"7F",X"7F",X"3F",X"07",X"FF",X"FE",X"FE",X"F8",X"F8",X"E0",X"E3",X"E3",
		X"8F",X"0F",X"3F",X"3F",X"FE",X"FF",X"FF",X"FF",X"FE",X"DF",X"BF",X"7F",X"FE",X"FE",X"FC",X"FC",
		X"1C",X"3F",X"3F",X"7F",X"7F",X"FE",X"FC",X"F8",X"00",X"87",X"FF",X"FF",X"3B",X"3D",X"7F",X"FF",
		X"FC",X"FF",X"FF",X"F8",X"F8",X"E0",X"E3",X"83",X"01",X"88",X"E0",X"FC",X"FE",X"FC",X"F8",X"FC",
		X"0E",X"1F",X"7B",X"77",X"EF",X"DE",X"7C",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"7F",X"3F",X"5F",X"1F",X"0F",X"87",X"11",
		X"FC",X"F8",X"F1",X"E3",X"C7",X"CF",X"FF",X"FF",X"FC",X"FE",X"FF",X"F7",X"EE",X"FC",X"F1",X"88",
		X"F1",X"E3",X"C7",X"CF",X"7F",X"7F",X"3F",X"07",X"FF",X"FE",X"FE",X"F8",X"F8",X"E0",X"E3",X"E3",
		X"8F",X"0F",X"3F",X"3F",X"FE",X"FF",X"FF",X"FF",X"FE",X"DF",X"BF",X"7F",X"FE",X"FE",X"FC",X"FC",
		X"1C",X"3F",X"3F",X"7F",X"7F",X"FE",X"FC",X"F8",X"00",X"87",X"FF",X"FF",X"3B",X"3D",X"7F",X"FF",
		X"FC",X"FF",X"FF",X"F8",X"F8",X"E0",X"E3",X"83",X"01",X"88",X"E0",X"FC",X"FE",X"FC",X"F8",X"FC",
		X"0E",X"1F",X"7B",X"77",X"EF",X"DE",X"7C",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"1F",X"01",X"07",X"1F",X"0F",X"07",X"07",X"FC",X"FC",X"C8",X"E0",X"F0",X"FC",X"F8",X"F8",
		X"06",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"B0",X"80",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",
		X"07",X"07",X"07",X"0F",X"0F",X"1F",X"1F",X"1F",X"F0",X"F0",X"F8",X"FC",X"FE",X"FE",X"FE",X"FE",
		X"09",X"01",X"03",X"01",X"00",X"00",X"00",X"00",X"FE",X"FE",X"F8",X"FC",X"EE",X"26",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"07",X"0F",X"1F",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",
		X"1F",X"1F",X"1F",X"1F",X"3F",X"3F",X"1F",X"1E",X"C0",X"E0",X"F0",X"F0",X"C0",X"A0",X"F8",X"FC",
		X"3F",X"3F",X"13",X"07",X"0F",X"3F",X"1F",X"1F",X"F8",X"F8",X"80",X"E0",X"F8",X"F0",X"E0",X"E0",
		X"0D",X"01",X"03",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",
		X"0F",X"0F",X"1F",X"3F",X"7F",X"7F",X"7F",X"7F",X"E0",X"E0",X"E0",X"F0",X"F0",X"F8",X"F8",X"F8",
		X"7F",X"7F",X"1F",X"3F",X"77",X"64",X"00",X"00",X"90",X"80",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"00",X"00",X"00",X"00",X"40",X"E0",X"F0",X"F8",
		X"03",X"07",X"0F",X"0F",X"03",X"05",X"1F",X"3F",X"F8",X"F8",X"F8",X"F8",X"FC",X"FC",X"F8",X"78",
		X"47",X"E6",X"E0",X"4F",X"2A",X"57",X"39",X"3E",X"60",X"08",X"DD",X"7E",X"01",X"BC",X"20",X"06",
		X"DD",X"7E",X"00",X"BD",X"28",X"0C",X"5E",X"23",X"7E",X"57",X"E6",X"E0",X"23",X"B9",X"30",X"19",
		X"2B",X"2B",X"78",X"A7",X"28",X"87",X"2B",X"77",X"E5",X"2A",X"2D",X"39",X"AF",X"CD",X"11",X"21",
		X"E1",X"2B",X"77",X"22",X"57",X"39",X"AF",X"3C",X"C9",X"C5",X"E5",X"DD",X"73",X"52",X"7A",X"E6",
		X"1F",X"87",X"87",X"5F",X"16",X"00",X"21",X"62",X"23",X"19",X"E5",X"FD",X"E3",X"FD",X"CB",X"FE",
		X"7E",X"28",X"0C",X"2A",X"59",X"39",X"36",X"00",X"23",X"36",X"00",X"23",X"22",X"59",X"39",X"CD",
		X"C6",X"20",X"2B",X"46",X"E5",X"2B",X"CB",X"7B",X"28",X"02",X"CB",X"FE",X"4E",X"78",X"07",X"AA",
		X"E6",X"01",X"AA",X"07",X"E6",X"03",X"67",X"FD",X"7E",X"FF",X"24",X"25",X"28",X"04",X"0F",X"0F",
		X"18",X"F9",X"E6",X"03",X"28",X"14",X"FE",X"02",X"38",X"0A",X"28",X"0C",X"D5",X"DD",X"5E",X"52",
		X"CD",X"FC",X"20",X"D1",X"CB",X"B8",X"18",X"02",X"CB",X"F8",X"E1",X"70",X"FD",X"46",X"FE",X"CB",
		X"68",X"20",X"10",X"DD",X"CB",X"08",X"4E",X"28",X"08",X"CB",X"76",X"28",X"04",X"CB",X"72",X"20",
		X"02",X"CB",X"E8",X"21",X"BC",X"21",X"FD",X"5E",X"00",X"16",X"00",X"FD",X"19",X"FD",X"E3",X"E3",
		X"E5",X"CD",X"C6",X"20",X"22",X"59",X"39",X"CB",X"79",X"C2",X"B7",X"21",X"CB",X"68",X"28",X"3C",
		X"CD",X"DA",X"20",X"CB",X"60",X"28",X"0F",X"AF",X"BA",X"20",X"05",X"7B",X"FE",X"11",X"38",X"06",
		X"CD",X"1E",X"24",X"11",X"11",X"00",X"D5",X"CD",X"C6",X"20",X"CD",X"DA",X"20",X"21",X"00",X"00",
		X"78",X"C1",X"CB",X"77",X"20",X"0E",X"CB",X"5F",X"20",X"03",X"79",X"B0",X"C9",X"CB",X"FC",X"19",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"4C",X"A9",X"C2",X"20",X"FC",X"E4",X"C2",X"20",
		X"FC",X"BB",X"62",X"20",X"FC",X"A2",X"62",X"20",X"FC",X"AC",X"81",X"08",X"50",X"48",X"81",X"08",
		X"50",X"3C",X"81",X"08",X"50",X"31",X"81",X"60",X"50",X"34",X"81",X"60",X"50",X"29",X"62",X"20",
		X"FC",X"3E",X"62",X"30",X"FC",X"4B",X"62",X"30",X"FC",X"51",X"62",X"20",X"FC",X"81",X"81",X"08",
		X"50",X"27",X"81",X"08",X"50",X"15",X"81",X"08",X"50",X"17",X"63",X"30",X"FC",X"33",X"05",X"00",
		X"00",X"00",X"06",X"00",X"00",X"00",X"C8",X"D8",X"2B",X"C9",X"D8",X"2B",X"C9",X"D0",X"2B",X"C9",
		X"28",X"FC",X"D0",X"2B",X"C9",X"C0",X"2B",X"C9",X"C8",X"2B",X"C9",X"2B",X"ED",X"52",X"C9",X"C8",
		X"D5",X"C5",X"CD",X"3F",X"24",X"C1",X"EB",X"CD",X"59",X"24",X"EB",X"E1",X"A7",X"ED",X"52",X"C9",
		X"41",X"EB",X"C8",X"CB",X"3C",X"CB",X"1D",X"10",X"FA",X"C9",X"41",X"EB",X"C8",X"CB",X"25",X"CB",
		X"14",X"DC",X"1E",X"24",X"10",X"F7",X"C9",X"2E",X"01",X"C8",X"EB",X"4D",X"44",X"3D",X"C8",X"F5",
		X"C5",X"EB",X"CD",X"59",X"24",X"C1",X"F1",X"18",X"F4",X"EB",X"ED",X"4A",X"E0",X"08",X"F6",X"0D",
		X"08",X"C9",X"EB",X"ED",X"42",X"18",X"F5",X"7B",X"B1",X"6F",X"7A",X"B0",X"67",X"C9",X"7B",X"A9",
		X"6F",X"7A",X"A8",X"67",X"C9",X"7B",X"A1",X"6F",X"7A",X"A0",X"67",X"C9",X"28",X"DF",X"21",X"00",
		X"00",X"3E",X"10",X"CB",X"23",X"CB",X"12",X"CB",X"15",X"CB",X"14",X"13",X"A7",X"ED",X"42",X"30",
		X"01",X"07",X"0F",X"1B",X"07",X"1B",X"03",X"0F",X"C0",X"F0",X"F8",X"E0",X"F0",X"F8",X"FC",X"E4",
		X"3F",X"17",X"0F",X"1F",X"F7",X"62",X"04",X"00",X"F0",X"F8",X"FE",X"EA",X"F0",X"7E",X"1A",X"00",
		X"01",X"07",X"0F",X"1B",X"07",X"1B",X"03",X"0F",X"C0",X"F0",X"F8",X"E0",X"F0",X"F8",X"FC",X"E4",
		X"3F",X"17",X"0F",X"1F",X"F7",X"62",X"04",X"00",X"F0",X"F8",X"FE",X"EA",X"F0",X"7E",X"1A",X"00",
		X"01",X"07",X"0F",X"1B",X"07",X"1B",X"03",X"0F",X"C0",X"F0",X"F8",X"E0",X"F0",X"F8",X"FC",X"E4",
		X"3F",X"17",X"0F",X"1F",X"F7",X"62",X"04",X"00",X"F0",X"F8",X"FE",X"EA",X"F0",X"7E",X"1A",X"00",
		X"00",X"01",X"06",X"39",X"42",X"82",X"A1",X"80",X"38",X"C4",X"0C",X"F0",X"00",X"F0",X"0C",X"02",
		X"60",X"10",X"10",X"10",X"13",X"0A",X"0A",X"1E",X"01",X"01",X"01",X"01",X"C2",X"21",X"41",X"7F",
		X"1C",X"25",X"7A",X"40",X"81",X"A5",X"81",X"42",X"78",X"84",X"04",X"78",X"80",X"00",X"F0",X"0C",
		X"3C",X"10",X"10",X"10",X"13",X"0A",X"0A",X"1E",X"02",X"01",X"01",X"01",X"C2",X"21",X"41",X"3F",
		X"F3",X"8C",X"F0",X"08",X"0A",X"74",X"83",X"78",X"CF",X"31",X"0F",X"10",X"50",X"2E",X"C1",X"1E",
		X"04",X"04",X"08",X"30",X"40",X"9E",X"E2",X"01",X"20",X"20",X"10",X"0C",X"02",X"79",X"47",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"FC",X"F8",X"F8",X"F8",X"F8",X"F0",X"F0",X"FC",X"FC",X"F8",X"F0",X"F0",X"F8",X"F8",X"FC",
		X"FF",X"FE",X"FC",X"FC",X"FE",X"FE",X"FE",X"FC",X"FF",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",
		X"FC",X"FC",X"F8",X"F8",X"F8",X"FE",X"FE",X"FF",X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",X"FC",X"FC",
		X"F0",X"F0",X"F0",X"F0",X"E0",X"E0",X"E0",X"F0",X"FE",X"FE",X"FC",X"FC",X"F8",X"F8",X"F0",X"F0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"39",X"22",X"2B",X"39",X"CD",X"49",X"1F",X"38",X"56",X"DD",X"CB",X"54",X"5E",X"28",X"45",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"07",
		X"00",X"00",X"80",X"F0",X"FE",X"FF",X"FF",X"FF",X"FF",X"1F",X"03",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"7F",X"3F",X"1F",X"0F",X"07",X"03",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"C0",X"F0",X"FC",X"FF",
		X"C0",X"F0",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"02",X"04",X"08",X"10",X"08",X"04",X"03",
		X"80",X"40",X"20",X"10",X"08",X"04",X"02",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"E0",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"0F",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"F8",X"FF",X"24",X"03",X"02",X"26",X"37",X"00",X"DF",X"0E",
		X"2C",X"18",X"27",X"3E",X"01",X"CF",X"18",X"10",X"AF",X"CF",X"0E",X"0C",X"18",X"1C",X"3E",X"81",
		X"CF",X"0E",X"2D",X"18",X"15",X"3E",X"81",X"CF",X"0E",X"0D",X"18",X"0E",X"3E",X"40",X"CF",X"18",
		X"E9",X"3E",X"41",X"CF",X"18",X"F2",X"AF",X"FE",X"01",X"C9",X"79",X"08",X"79",X"CB",X"71",X"28",
		X"1D",X"21",X"A8",X"17",X"CD",X"30",X"00",X"D8",X"08",X"47",X"08",X"78",X"E6",X"20",X"B1",X"DD",
		X"77",X"06",X"0E",X"01",X"FE",X"06",X"30",X"06",X"DD",X"CB",X"54",X"76",X"20",X"0F",X"2A",X"77",
		X"39",X"11",X"06",X"39",X"E6",X"3F",X"12",X"D7",X"20",X"CC",X"22",X"77",X"39",X"DD",X"71",X"51",
		X"CB",X"71",X"20",X"20",X"CB",X"69",X"28",X"1C",X"DD",X"CB",X"51",X"FE",X"3E",X"20",X"B9",X"20",
		X"13",X"0E",X"C0",X"21",X"FC",X"0F",X"18",X"E2",X"CB",X"71",X"C2",X"1D",X"16",X"DD",X"7E",X"51",
		X"E6",X"1F",X"3D",X"E7",X"08",X"CB",X"77",X"28",X"EF",X"DD",X"7E",X"06",X"FE",X"38",X"38",X"08",
		X"FE",X"3B",X"30",X"04",X"DD",X"36",X"06",X"06",X"E6",X"1F",X"FE",X"19",X"20",X"0A",X"DD",X"CB",
		X"0E",X"6E",X"DD",X"CB",X"0E",X"EE",X"18",X"0C",X"FE",X"1A",X"20",X"0B",X"DD",X"CB",X"0E",X"76",
		X"DD",X"CB",X"0E",X"F6",X"CC",X"49",X"18",X"DD",X"7E",X"06",X"CB",X"67",X"28",X"07",X"07",X"07",
		X"E6",X"30",X"DD",X"77",X"06",X"BF",X"C9",X"AB",X"41",X"42",X"43",X"44",X"45",X"48",X"4C",X"46",
		X"49",X"52",X"53",X"CB",X"CE",X"01",X"D0",X"03",X"D2",X"05",X"06",X"D3",X"09",X"D7",X"81",X"46",
		X"1D",X"07",X"81",X"43",X"10",X"00",X"81",X"45",X"14",X"02",X"81",X"4C",X"18",X"04",X"82",X"58",
		X"59",X"19",X"1A",X"08",X"A1",X"50",X"1C",X"DD",X"CB",X"08",X"86",X"DD",X"CB",X"09",X"AE",X"21",
		X"00",X"00",X"22",X"37",X"39",X"21",X"3F",X"3B",X"22",X"59",X"39",X"C9",X"2A",X"25",X"39",X"E5",
		X"11",X"7F",X"3A",X"A7",X"ED",X"52",X"ED",X"5B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"24",X"24",X"24",X"24",X"24",X"00",X"24",X"24",
		X"77",X"55",X"55",X"55",X"55",X"55",X"77",X"00",X"06",X"02",X"02",X"02",X"02",X"02",X"07",X"00",
		X"06",X"09",X"01",X"01",X"06",X"08",X"0F",X"00",X"06",X"09",X"01",X"06",X"01",X"09",X"06",X"00",
		X"02",X"06",X"0A",X"12",X"12",X"1F",X"02",X"00",X"0F",X"08",X"08",X"07",X"01",X"09",X"0F",X"00",
		X"06",X"09",X"08",X"0E",X"09",X"09",X"06",X"00",X"0F",X"01",X"02",X"04",X"08",X"08",X"08",X"00",
		X"06",X"09",X"09",X"06",X"09",X"09",X"06",X"00",X"06",X"09",X"09",X"07",X"01",X"09",X"06",X"00",
		X"67",X"25",X"25",X"25",X"25",X"25",X"77",X"00",X"00",X"03",X"0C",X"13",X"24",X"44",X"88",X"88",
		X"FF",X"00",X"7F",X"80",X"00",X"00",X"00",X"00",X"80",X"60",X"18",X"C6",X"21",X"11",X"09",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"04",X"0A",X"15",X"09",X"09",X"30",
		X"00",X"00",X"80",X"40",X"40",X"20",X"20",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"0B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"07",X"1B",X"24",X"48",X"50",X"90",X"90",X"20",X"80",X"40",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"B1",X"BB",X"3F",X"3F",X"1F",X"00",X"00",X"00",X"FF",X"80",X"FF",X"00",X"FC",
		X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"0A",X"0A",X"12",X"12",
		X"88",X"84",X"44",X"42",X"21",X"18",X"07",X"00",X"00",X"00",X"00",X"00",X"C0",X"38",X"07",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"0E",X"0A",X"0E",X"00",X"00",X"00",X"00",
		X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"A0",X"90",X"50",X"50",X"50",X"50",X"50",X"50",
		X"1D",X"08",X"09",X"1D",X"09",X"00",X"00",X"00",X"00",X"40",X"C0",X"C0",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"24",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"02",X"02",X"02",X"04",X"04",X"04",X"20",X"40",X"40",X"40",X"80",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"0F",X"0F",X"07",X"05",X"00",X"00",X"00",
		X"00",X"F0",X"58",X"B7",X"D4",X"EB",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"30",X"00",X"00",
		X"12",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"50",
		X"06",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"08",X"84",X"42",X"21",X"11",X"11",X"11",
		X"00",X"00",X"00",X"0C",X"0A",X"0A",X"0A",X"0A",X"30",X"30",X"30",X"28",X"28",X"18",X"18",X"15",
		X"50",X"50",X"60",X"A0",X"A0",X"A1",X"A1",X"42",X"00",X"00",X"00",X"00",X"F0",X"68",X"98",X"98",
		X"00",X"00",X"00",X"00",X"60",X"50",X"50",X"31",X"00",X"00",X"00",X"00",X"38",X"7C",X"C6",X"86",
		X"3C",X"00",X"00",X"30",X"2C",X"13",X"16",X"29",X"00",X"00",X"00",X"00",X"00",X"C0",X"40",X"40",
		X"00",X"00",X"00",X"1E",X"21",X"5C",X"62",X"61",X"09",X"09",X"09",X"09",X"91",X"52",X"22",X"82",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"36",X"49",
		X"00",X"00",X"00",X"00",X"00",X"80",X"81",X"82",X"00",X"00",X"00",X"00",X"00",X"EF",X"1C",X"12",
		X"00",X"00",X"00",X"00",X"03",X"04",X"89",X"92",X"14",X"14",X"14",X"14",X"D8",X"E8",X"28",X"18",
		X"88",X"84",X"42",X"21",X"18",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"FF",X"00",
		X"11",X"21",X"22",X"44",X"88",X"07",X"FF",X"00",X"12",X"11",X"29",X"55",X"A2",X"C2",X"03",X"00",
		X"15",X"0A",X"08",X"05",X"88",X"76",X"F9",X"00",X"43",X"83",X"83",X"05",X"86",X"FA",X"FC",X"00",
		X"28",X"30",X"30",X"30",X"2C",X"23",X"1F",X"00",X"29",X"55",X"6A",X"A4",X"A3",X"C0",X"00",X"00",
		X"8A",X"8C",X"94",X"68",X"10",X"8F",X"7F",X"00",X"31",X"31",X"52",X"52",X"A2",X"21",X"C0",X"00",
		X"40",X"80",X"80",X"80",X"4C",X"34",X"F8",X"00",X"A0",X"C0",X"A0",X"50",X"49",X"26",X"1F",X"00",
		X"42",X"24",X"23",X"CC",X"13",X"20",X"C0",X"00",X"00",X"00",X"01",X"81",X"61",X"DF",X"3E",X"00",
		X"92",X"A3",X"43",X"43",X"22",X"1F",X"FC",X"00",X"83",X"06",X"06",X"0C",X"94",X"68",X"F1",X"00",
		X"A2",X"A3",X"A5",X"A5",X"C4",X"C2",X"C1",X"00",X"54",X"14",X"14",X"18",X"A8",X"57",X"EF",X"00",
		X"18",X"18",X"18",X"24",X"54",X"AB",X"C7",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"01",X"01",X"03",X"03",X"03",X"07",
		X"00",X"FA",X"8B",X"A5",X"E9",X"4F",X"11",X"BB",X"00",X"3C",X"18",X"31",X"31",X"61",X"63",X"FE",
		X"00",X"70",X"C9",X"83",X"83",X"86",X"8B",X"F1",X"00",X"E7",X"93",X"1B",X"1A",X"1C",X"34",X"EE",
		X"00",X"1C",X"88",X"90",X"D0",X"70",X"60",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"18",X"01",X"B6",X"77",X"3C",X"C9",X"1E",X"08",X"DD",X"36",X"0C",X"06",X"DD",X"CB",X"50",X"DE",
		X"53",X"CD",X"83",X"1C",X"21",X"12",X"10",X"ED",X"7B",X"4B",X"39",X"DD",X"21",X"FF",X"38",X"E9",
		X"21",X"6E",X"10",X"30",X"F2",X"C2",X"69",X"1B",X"EB",X"E5",X"2B",X"36",X"0D",X"22",X"0F",X"39",
		X"16",X"10",X"CD",X"83",X"1C",X"D1",X"C3",X"8E",X"2B",X"21",X"FA",X"10",X"18",X"E5",X"21",X"52",
		X"45",X"3E",X"4C",X"DD",X"CB",X"0F",X"76",X"28",X"05",X"21",X"41",X"42",X"3E",X"53",X"22",X"E3",
		X"38",X"32",X"E5",X"38",X"3E",X"32",X"32",X"CC",X"38",X"AF",X"32",X"09",X"39",X"21",X"00",X"00",
		X"22",X"65",X"39",X"22",X"75",X"39",X"22",X"5F",X"39",X"22",X"67",X"39",X"22",X"1D",X"39",X"22",
		X"3B",X"39",X"22",X"3D",X"39",X"22",X"1F",X"39",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
