library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity dotron_bg_bits_1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of dotron_bg_bits_1 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"FF",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"54",X"00",X"55",X"50",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"54",X"00",X"55",X"00",X"55",X"40",
		X"55",X"40",X"55",X"50",X"55",X"50",X"55",X"50",X"55",X"50",X"55",X"50",X"55",X"40",X"55",X"40",
		X"55",X"00",X"55",X"00",X"54",X"00",X"50",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"54",X"55",X"40",X"40",X"00",
		X"54",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"54",X"00",X"55",X"40",X"55",X"54",X"55",X"55",
		X"50",X"00",X"54",X"00",X"55",X"00",X"55",X"40",X"55",X"50",X"55",X"54",X"55",X"55",X"55",X"55",
		X"40",X"00",X"50",X"00",X"50",X"00",X"54",X"00",X"54",X"00",X"55",X"00",X"55",X"00",X"55",X"00",
		X"00",X"00",X"55",X"00",X"55",X"54",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"54",X"00",
		X"01",X"55",X"05",X"55",X"05",X"55",X"05",X"55",X"05",X"55",X"05",X"55",X"01",X"55",X"01",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"15",X"00",X"55",X"01",X"55",
		X"00",X"00",X"00",X"15",X"05",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"7F",X"FD",X"7D",X"5D",X"7D",X"5D",X"75",X"5D",X"75",X"5D",X"75",X"5D",X"7F",X"FD",
		X"55",X"55",X"57",X"55",X"57",X"55",X"57",X"55",X"57",X"D5",X"57",X"D5",X"57",X"D5",X"57",X"D5",
		X"55",X"55",X"7F",X"FD",X"75",X"5D",X"75",X"55",X"7F",X"FD",X"55",X"7D",X"55",X"7D",X"7F",X"FD",
		X"55",X"55",X"5F",X"FD",X"5D",X"55",X"7F",X"55",X"7D",X"55",X"7D",X"55",X"7D",X"5D",X"7F",X"FD",
		X"55",X"55",X"5D",X"55",X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",X"7F",X"FD",X"5F",X"55",X"5F",X"55",
		X"55",X"55",X"7F",X"FD",X"55",X"5D",X"55",X"5D",X"7F",X"FD",X"7D",X"55",X"7D",X"5D",X"7F",X"FD",
		X"55",X"55",X"7F",X"FD",X"55",X"5D",X"55",X"5D",X"7F",X"FD",X"7D",X"5D",X"7D",X"5D",X"7F",X"FD",
		X"55",X"55",X"7F",X"FD",X"75",X"55",X"75",X"55",X"7D",X"55",X"7D",X"55",X"7D",X"55",X"7D",X"55",
		X"55",X"55",X"5F",X"F5",X"5D",X"75",X"5D",X"75",X"7F",X"FD",X"7D",X"5D",X"7D",X"5D",X"7F",X"FD",
		X"55",X"55",X"7F",X"FD",X"75",X"5D",X"75",X"5D",X"7F",X"FD",X"7D",X"55",X"7D",X"55",X"7F",X"FD",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"FF",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"15",X"55",X"01",X"55",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"01",X"00",X"05",X"00",X"05",X"00",X"15",X"00",X"15",X"00",X"55",X"00",X"55",X"00",X"55",
		X"00",X"05",X"00",X"15",X"00",X"55",X"01",X"55",X"05",X"55",X"15",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"15",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"15",X"01",X"55",X"15",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"55",X"15",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"55",X"00",X"55",X"00",X"15",X"00",X"05",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"FF",X"08",X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"08",X"44",X"09",X"55",X"09",X"55",
		X"09",X"55",X"09",X"55",X"09",X"55",X"0A",X"66",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"FA",X"AA",
		X"FB",X"BB",X"0B",X"FF",X"0B",X"FF",X"0B",X"FF",X"0B",X"FF",X"0B",X"77",X"09",X"55",X"09",X"55",
		X"C0",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"03",X"80",X"0D",X"80",X"09",X"80",X"35",
		X"80",X"25",X"80",X"D5",X"80",X"95",X"80",X"A6",X"83",X"AA",X"82",X"AA",X"82",X"AA",X"BE",X"AA",
		X"BE",X"AA",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",
		X"80",X"03",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",
		X"09",X"55",X"09",X"55",X"09",X"55",X"09",X"55",X"09",X"55",X"09",X"55",X"09",X"55",X"0A",X"AA",
		X"EE",X"EE",X"2F",X"FE",X"3F",X"FE",X"2F",X"FE",X"FF",X"FE",X"B7",X"78",X"55",X"58",X"55",X"58",
		X"55",X"60",X"55",X"5C",X"55",X"58",X"A6",X"68",X"AA",X"AB",X"2A",X"AA",X"2A",X"AA",X"EA",X"AA",
		X"00",X"A5",X"00",X"09",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FC",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"55",X"55",X"AA",X"55",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"55",X"55",X"AA",X"AA",
		X"00",X"FF",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"91",X"00",X"95",X"00",X"AA",
		X"55",X"60",X"55",X"80",X"55",X"80",X"56",X"00",X"58",X"00",X"60",X"00",X"80",X"00",X"00",X"00",
		X"FF",X"F5",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"AA",X"A8",
		X"FF",X"FF",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"AA",X"AA",
		X"00",X"BF",X"00",X"95",X"00",X"95",X"00",X"95",X"00",X"95",X"00",X"95",X"00",X"95",X"00",X"AA",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"3D",
		X"00",X"00",X"C0",X"00",X"30",X"00",X"0C",X"00",X"03",X"00",X"11",X"C0",X"55",X"80",X"55",X"70",
		X"00",X"FF",X"0F",X"00",X"30",X"00",X"C0",X"00",X"00",X"00",X"11",X"11",X"55",X"55",X"55",X"56",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"55",X"55",X"AA",X"AA",
		X"FF",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"12",X"00",X"56",X"00",X"AA",X"00",
		X"55",X"68",X"55",X"80",X"56",X"00",X"68",X"00",X"A8",X"00",X"A0",X"00",X"A0",X"00",X"AF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"AF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"AA",X"AA",
		X"FF",X"F5",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"AA",X"A8",
		X"55",X"60",X"55",X"80",X"55",X"80",X"56",X"00",X"58",X"00",X"60",X"00",X"80",X"00",X"00",X"00",
		X"FF",X"FF",X"2F",X"FE",X"2F",X"FE",X"2F",X"FE",X"FF",X"F8",X"9D",X"D8",X"55",X"58",X"55",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"CC",X"F3",X"CC",X"CC",X"CC",X"C0",X"CC",
		X"FF",X"FF",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"FF",X"FF",
		X"FB",X"BB",X"0B",X"FF",X"0B",X"FF",X"0B",X"FF",X"02",X"FF",X"02",X"DD",X"02",X"55",X"00",X"95",
		X"00",X"95",X"03",X"55",X"02",X"55",X"02",X"99",X"0E",X"AA",X"0A",X"AA",X"0A",X"AA",X"FA",X"AA",
		X"55",X"A3",X"56",X"03",X"58",X"03",X"A0",X"03",X"A0",X"03",X"80",X"03",X"80",X"03",X"BF",X"FF",
		X"03",X"FF",X"3C",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"44",X"44",X"55",X"55",X"55",X"5A",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"3D",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"95",X"00",X"25",X"00",X"25",X"00",X"09",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"5F",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"95",X"55",X"29",X"55",X"02",X"AA",
		X"FF",X"FF",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"AA",X"AA",
		X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"FF",X"FF",
		X"BF",X"FF",X"C0",X"03",X"80",X"03",X"F0",X"03",X"E0",X"03",X"DC",X"03",X"57",X"03",X"55",X"F3",
		X"FF",X"FF",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"0C",X"00",X"34",X"00",X"25",X"00",X"D5",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"44",X"55",X"55",X"AA",X"AA",
		X"C0",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",
		X"C0",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",
		X"00",X"0A",X"00",X"2A",X"00",X"AA",X"02",X"AA",X"02",X"AA",X"0A",X"AB",X"0A",X"A3",X"0A",X"A3",
		X"0A",X"A3",X"0A",X"A3",X"0A",X"AB",X"02",X"AA",X"02",X"AA",X"00",X"AA",X"00",X"2A",X"00",X"0A",
		X"CA",X"A0",X"CA",X"A0",X"EA",X"A0",X"AA",X"80",X"AA",X"80",X"AA",X"00",X"A8",X"00",X"A0",X"00",
		X"A0",X"00",X"A8",X"00",X"AA",X"00",X"AA",X"80",X"AA",X"80",X"EA",X"A0",X"CA",X"A0",X"CA",X"A0",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"80",X"AA",X"80",X"AA",X"80",X"AA",X"80",X"AA",X"80",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"80",X"AA",X"AA",X"AA",X"AA",
		X"A8",X"00",X"A8",X"00",X"A8",X"00",X"A8",X"00",X"A8",X"00",X"00",X"00",X"A8",X"00",X"A8",X"00",
		X"A8",X"00",X"A8",X"00",X"A8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"2A",X"AA",X"2A",X"AA",
		X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"AA",X"00",X"00",X"00",X"00",
		X"AA",X"80",X"AA",X"80",X"AA",X"80",X"AA",X"80",X"AA",X"80",X"AA",X"80",X"00",X"00",X"00",X"00",
		X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"EA",X"AA",X"EA",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",
		X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"00",
		X"00",X"00",X"A0",X"00",X"A8",X"00",X"AA",X"00",X"AA",X"80",X"AA",X"80",X"AA",X"A0",X"2A",X"A0",
		X"2A",X"A0",X"2A",X"A8",X"0A",X"A8",X"FA",X"AB",X"FF",X"FF",X"80",X"00",X"A0",X"00",X"A8",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",X"A8",X"AA",X"A8",X"2A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FA",X"00",X"0A",X"00",X"0A",X"00",X"0A",
		X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"0A",X"00",X"00",X"00",X"00",
		X"A8",X"0A",X"A8",X"02",X"A8",X"00",X"A8",X"00",X"A8",X"00",X"A8",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"00",X"AA",X"80",X"AA",X"A0",X"2A",X"A8",X"0A",X"AA",X"02",X"AA",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"2A",X"AB",X"0A",X"AA",X"0A",X"AA",X"02",X"AA",X"00",X"AA",X"80",X"0A",X"00",X"03",X"00",X"03",
		X"EA",X"A8",X"AA",X"A0",X"AA",X"A0",X"AA",X"80",X"AA",X"00",X"A0",X"00",X"C0",X"00",X"C0",X"00",
		X"AA",X"83",X"AA",X"83",X"AA",X"03",X"AA",X"FF",X"AA",X"FF",X"AA",X"83",X"AA",X"83",X"2A",X"A3",
		X"00",X"0A",X"00",X"AA",X"02",X"AA",X"0A",X"AA",X"0A",X"AA",X"2A",X"AA",X"2A",X"AB",X"2A",X"A3",
		X"A0",X"00",X"AA",X"00",X"AA",X"80",X"AA",X"A0",X"AA",X"A0",X"AA",X"A8",X"EA",X"A8",X"CA",X"A8",
		X"C2",X"AA",X"C2",X"AA",X"C0",X"AA",X"FF",X"AA",X"FF",X"AA",X"C2",X"AA",X"C2",X"AA",X"CA",X"A8",
		X"2A",X"A0",X"2A",X"A0",X"2A",X"A0",X"2A",X"A0",X"2A",X"A0",X"2A",X"A0",X"00",X"00",X"00",X"00",
		X"2A",X"AA",X"2A",X"AA",X"2A",X"AA",X"EA",X"AA",X"EA",X"AF",X"2A",X"A0",X"2A",X"A0",X"2A",X"A0",
		X"20",X"00",X"28",X"00",X"2A",X"00",X"2A",X"80",X"2A",X"A0",X"2A",X"A8",X"2A",X"AA",X"2A",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"30",X"30",X"C0",X"30",X"C0",X"3C",X"C0",
		X"A0",X"00",X"A8",X"00",X"AA",X"00",X"AA",X"BF",X"FF",X"EA",X"00",X"0A",X"00",X"02",X"00",X"00",
		X"0A",X"A8",X"0A",X"A8",X"0A",X"A8",X"FA",X"AB",X"AA",X"AB",X"AA",X"A8",X"AA",X"A8",X"AA",X"A8",
		X"2A",X"A8",X"0A",X"A8",X"02",X"A8",X"00",X"A8",X"00",X"28",X"00",X"08",X"00",X"00",X"00",X"00",
		X"0A",X"A8",X"0A",X"A8",X"0A",X"A8",X"0A",X"A8",X"0A",X"A8",X"0A",X"A8",X"0A",X"A8",X"0A",X"A8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"0C",X"0C",X"CC",X"CF",X"CC",X"CC",X"CF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"00",X"33",X"00",X"3C",X"00",X"3F",
		X"0F",X"C0",X"30",X"30",X"C3",X"0C",X"CC",X"0C",X"CC",X"0C",X"C3",X"0C",X"30",X"30",X"0F",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"00",X"03",X"00",X"03",X"FF",X"FF",X"FF",X"FF",X"00",X"03",X"00",X"03",X"00",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"F0",X"FF",X"FC",X"00",X"3F",X"00",X"0F",X"00",X"03",
		X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",
		X"00",X"00",X"33",X"F3",X"33",X"33",X"33",X"33",X"33",X"F3",X"30",X"33",X"30",X"33",X"00",X"00",
		X"00",X"00",X"F3",X"F0",X"30",X"30",X"F3",X"F0",X"30",X"30",X"30",X"30",X"F3",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"30",X"00",X"F0",X"00",X"30",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"00",X"33",X"00",X"33",X"00",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"0C",X"33",X"CC",X"33",X"3C",X"33",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C3",X"3C",X"F3",X"3C",X"CF",X"30",X"C3",X"3C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"C0",X"CC",X"F3",X"F0",X"CC",X"CC",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C3",X"0C",X"CC",X"CF",X"CF",X"CC",X"CC",X"CC",
		X"0F",X"C0",X"30",X"30",X"C3",X"0C",X"CC",X"CC",X"CF",X"CC",X"CC",X"CC",X"30",X"30",X"0F",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"3C",X"3F",X"33",X"30",X"3F",X"3C",X"33",X"30",X"33",X"30",X"3F",X"30",X"00",X"00",
		X"00",X"00",X"0F",X"00",X"30",X"C0",X"30",X"00",X"30",X"00",X"30",X"C0",X"0F",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"C0",X"CC",X"CC",X"CC",X"33",X"F0",X"33",
		X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"FF",X"3F",X"C0",X"FC",X"00",X"F0",X"00",X"F0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C3",X"0C",X"CC",X"C3",X"0F",X"C3",X"0C",X"C3",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"F0",X"3F",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"FF",X"D7",
		X"FF",X"57",X"3F",X"57",X"0F",X"55",X"01",X"55",X"01",X"55",X"01",X"55",X"11",X"55",X"01",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"44",X"50",X"44",X"54",X"44",X"54",X"44",X"54",X"44",X"54",X"44",
		X"00",X"00",X"00",X"00",X"01",X"10",X"01",X"00",X"00",X"00",X"01",X"10",X"11",X"00",X"51",X"54",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"54",X"54",X"55",X"04",X"55",X"45",X"55",X"45",X"55",X"45",X"55",X"45",X"55",X"50",X"55",X"14",
		X"50",X"54",X"50",X"54",X"00",X"55",X"50",X"55",X"51",X"55",X"10",X"55",X"41",X"55",X"51",X"55",
		X"00",X"00",X"00",X"00",X"10",X"04",X"01",X"04",X"00",X"15",X"01",X"15",X"40",X"05",X"00",X"45",
		X"00",X"00",X"01",X"00",X"41",X"50",X"05",X"50",X"15",X"54",X"10",X"50",X"15",X"50",X"17",X"50",
		X"00",X"00",X"40",X"00",X"54",X"00",X"44",X"50",X"50",X"44",X"44",X"44",X"44",X"44",X"41",X"50",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",
		X"55",X"54",X"51",X"54",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"5D",X"55",X"55",
		X"54",X"55",X"5D",X"55",X"55",X"55",X"55",X"55",X"57",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"50",X"45",X"10",X"55",X"14",X"55",X"44",X"55",X"50",X"55",X"54",X"55",X"55",X"15",X"51",X"55",
		X"15",X"54",X"11",X"55",X"51",X"54",X"11",X"50",X"45",X"50",X"55",X"54",X"15",X"54",X"11",X"54",
		X"15",X"4C",X"15",X"55",X"15",X"55",X"15",X"55",X"15",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"04",X"04",X"55",X"14",X"45",X"14",X"55",X"11",X"55",X"11",X"55",X"55",X"55",X"11",X"55",X"45",
		X"00",X"00",X"57",X"50",X"01",X"01",X"11",X"15",X"01",X"15",X"11",X"15",X"11",X"15",X"07",X"41",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"10",X"11",X"10",X"44",X"10",X"04",X"00",X"44",X"14",
		X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"10",X"01",X"10",X"00",X"10",X"01",X"50",X"15",X"54",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"D4",X"55",X"55",X"55",X"54",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"5C",X"55",X"D4",X"55",X"55",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"54",
		X"57",X"55",X"55",X"75",X"55",X"5D",X"55",X"55",X"55",X"75",X"55",X"55",X"55",X"55",X"55",X"55",
		X"45",X"05",X"45",X"41",X"45",X"55",X"45",X"D4",X"44",X"54",X"01",X"05",X"51",X"50",X"51",X"55",
		X"10",X"00",X"00",X"14",X"50",X"10",X"10",X"10",X"10",X"15",X"10",X"54",X"00",X"51",X"10",X"14",
		X"01",X"00",X"01",X"50",X"11",X"04",X"01",X"01",X"41",X"45",X"41",X"15",X"41",X"55",X"41",X"54",
		X"00",X"00",X"00",X"40",X"00",X"55",X"45",X"41",X"45",X"55",X"55",X"04",X"55",X"05",X"5D",X"15",
		X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"05",X"50",X"05",X"50",X"05",X"54",X"45",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"04",X"05",
		X"00",X"00",X"10",X"00",X"10",X"10",X"54",X"04",X"55",X"00",X"55",X"00",X"55",X"55",X"75",X"55",
		X"00",X"40",X"00",X"40",X"00",X"54",X"00",X"50",X"51",X"45",X"01",X"45",X"41",X"45",X"45",X"45",
		X"00",X"00",X"00",X"01",X"05",X"51",X"45",X"51",X"45",X"45",X"55",X"55",X"55",X"15",X"55",X"55",
		X"15",X"54",X"57",X"54",X"55",X"54",X"55",X"54",X"55",X"54",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"01",X"00",X"01",X"00",X"11",X"15",X"11",X"15",X"05",X"55",X"51",X"55",X"41",X"55",X"41",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"54",X"5D",X"D5",X"55",X"55",X"55",X"55",X"55",X"D5",
		X"14",X"10",X"14",X"14",X"05",X"05",X"45",X"45",X"05",X"45",X"45",X"54",X"51",X"55",X"45",X"55",
		X"41",X"55",X"05",X"55",X"55",X"55",X"15",X"55",X"15",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"15",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"45",X"54",X"45",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"45",X"44",X"45",X"40",X"45",X"55",X"05",X"55",X"45",X"51",X"15",X"55",X"55",X"55",X"55",
		X"45",X"45",X"51",X"45",X"54",X"15",X"54",X"45",X"55",X"55",X"55",X"15",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"D5",X"5D",X"55",X"55",X"55",X"55",X"D5",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"57",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"5F",X"FF",X"F5",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"FF",X"FF",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"57",X"55",X"5D",X"55",X"F5",
		X"55",X"5D",X"55",X"F5",X"57",X"55",X"5D",X"55",X"F5",X"55",X"55",X"56",X"55",X"59",X"55",X"65",
		X"55",X"55",X"55",X"55",X"56",X"AA",X"59",X"55",X"A5",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"AA",X"AA",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"57",X"55",X"5D",X"55",X"F5",X"57",X"55",X"5D",X"55",
		X"57",X"55",X"5D",X"55",X"F5",X"55",X"55",X"55",X"55",X"5A",X"55",X"65",X"55",X"95",X"56",X"55",
		X"56",X"95",X"59",X"55",X"65",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"54",X"00",X"51",X"55",X"45",X"55",X"15",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"57",
		X"55",X"55",X"55",X"57",X"55",X"5D",X"55",X"F5",X"57",X"55",X"5D",X"55",X"F5",X"55",X"55",X"55",
		X"F5",X"55",X"55",X"55",X"55",X"56",X"55",X"59",X"55",X"A5",X"56",X"55",X"59",X"55",X"65",X"55",
		X"69",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"54",X"55",X"51",X"55",X"45",X"55",X"15",X"54",X"55",X"51",X"57",X"45",X"5D",X"15",X"5D",
		X"55",X"55",X"57",X"FF",X"5D",X"55",X"75",X"55",X"D5",X"55",X"55",X"55",X"56",X"AA",X"59",X"55",
		X"55",X"55",X"FF",X"FF",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"AA",X"AA",X"55",X"55",
		X"14",X"00",X"15",X"50",X"15",X"55",X"15",X"55",X"95",X"55",X"95",X"55",X"95",X"55",X"95",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"57",X"55",X"5D",X"55",X"F5",
		X"55",X"5D",X"55",X"F5",X"57",X"55",X"5D",X"55",X"F5",X"55",X"55",X"55",X"55",X"55",X"55",X"56",
		X"55",X"56",X"55",X"59",X"55",X"65",X"55",X"95",X"5A",X"55",X"65",X"55",X"95",X"55",X"55",X"55",
		X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"54",X"55",X"51",X"55",X"45",X"55",X"15",X"54",X"55",X"51",X"55",X"45",X"55",X"15",X"57",
		X"55",X"75",X"55",X"D5",X"57",X"55",X"5D",X"56",X"75",X"59",X"D5",X"65",X"D5",X"95",X"55",X"95",
		X"65",X"55",X"65",X"55",X"95",X"55",X"54",X"00",X"51",X"55",X"45",X"55",X"45",X"55",X"15",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"95",X"55",X"95",X"55",X"95",X"55",X"95",X"55",X"15",X"55",X"15",X"55",X"15",X"55",X"15",X"55",
		X"94",X"00",X"95",X"50",X"95",X"55",X"95",X"55",X"15",X"55",X"15",X"55",X"15",X"55",X"15",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"57",X"55",X"5D",X"55",X"F5",X"57",X"55",X"5D",X"55",
		X"57",X"55",X"5D",X"55",X"F5",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"59",X"55",X"65",
		X"55",X"69",X"55",X"95",X"56",X"55",X"59",X"55",X"A5",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"54",X"55",X"51",X"55",X"45",X"55",X"15",X"54",X"55",X"51",X"55",X"45",X"55",X"15",X"57",
		X"55",X"5D",X"55",X"75",X"55",X"D5",X"57",X"55",X"5D",X"56",X"75",X"56",X"D5",X"59",X"55",X"65",
		X"56",X"54",X"59",X"51",X"65",X"51",X"95",X"45",X"55",X"15",X"54",X"55",X"54",X"57",X"51",X"5D",
		X"57",X"FF",X"5D",X"55",X"5D",X"55",X"75",X"55",X"D5",X"55",X"D6",X"AA",X"59",X"55",X"59",X"55",
		X"FF",X"FF",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"AA",X"AA",X"55",X"55",X"55",X"55",
		X"95",X"55",X"95",X"55",X"95",X"55",X"15",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"54",X"00",X"55",X"50",X"55",X"55",X"55",X"55",X"55",X"55",X"95",X"55",X"95",X"55",X"95",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"57",
		X"55",X"55",X"55",X"57",X"55",X"5D",X"55",X"F5",X"57",X"55",X"5D",X"55",X"F5",X"55",X"55",X"55",
		X"F5",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"5A",X"55",X"65",X"55",X"95",X"56",X"55",
		X"56",X"95",X"59",X"55",X"65",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"54",X"55",X"51",X"55",X"45",X"55",X"15",X"54",X"55",X"51",X"55",X"45",X"55",X"15",X"55",
		X"55",X"5D",X"55",X"5D",X"55",X"75",X"55",X"D5",X"57",X"55",X"5D",X"55",X"75",X"56",X"D5",X"59",
		X"55",X"95",X"56",X"55",X"59",X"55",X"59",X"54",X"65",X"51",X"95",X"45",X"55",X"45",X"55",X"15",
		X"45",X"5D",X"15",X"75",X"15",X"D5",X"55",X"D6",X"57",X"56",X"5D",X"59",X"75",X"65",X"75",X"65",
		X"65",X"55",X"65",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"95",X"00",X"95",X"55",X"95",X"55",X"95",X"55",X"15",X"55",X"15",X"55",X"15",X"55",X"15",X"55",
		X"94",X"00",X"95",X"50",X"95",X"55",X"95",X"55",X"95",X"55",X"95",X"55",X"95",X"55",X"95",X"55",
		X"55",X"5D",X"55",X"F5",X"57",X"55",X"5D",X"55",X"F5",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"59",X"55",X"A5",X"56",X"55",X"59",X"55",X"65",X"55",
		X"69",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"54",X"55",X"51",X"55",X"45",X"55",X"15",X"54",X"55",X"51",X"55",X"45",X"55",X"15",X"55",
		X"55",X"57",X"55",X"5D",X"55",X"75",X"55",X"D5",X"55",X"D5",X"57",X"55",X"5D",X"55",X"75",X"55",
		X"55",X"65",X"55",X"65",X"55",X"95",X"56",X"55",X"59",X"55",X"65",X"54",X"95",X"54",X"95",X"51",
		X"54",X"55",X"51",X"57",X"51",X"57",X"45",X"5D",X"15",X"75",X"55",X"75",X"55",X"D5",X"57",X"55",
		X"D5",X"95",X"56",X"55",X"56",X"55",X"59",X"55",X"65",X"55",X"65",X"55",X"95",X"55",X"95",X"55",
		X"95",X"55",X"95",X"55",X"95",X"55",X"95",X"55",X"95",X"55",X"95",X"55",X"95",X"55",X"95",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"95",X"55",X"95",X"55",X"95",X"55",X"95",X"55",
		X"15",X"55",X"15",X"55",X"15",X"55",X"95",X"55",X"95",X"55",X"95",X"55",X"95",X"55",X"95",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"56",X"55",X"59",X"55",X"65",X"55",X"95",X"5A",X"55",X"65",X"55",X"95",X"55",X"55",X"55",
		X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"54",X"55",X"51",X"55",X"45",X"55",X"15",X"54",X"55",X"51",X"55",X"45",X"55",X"15",X"55",
		X"55",X"55",X"55",X"57",X"55",X"5D",X"55",X"75",X"55",X"D5",X"57",X"55",X"5D",X"55",X"5D",X"55",
		X"D5",X"56",X"55",X"59",X"55",X"65",X"55",X"95",X"56",X"55",X"56",X"55",X"59",X"55",X"65",X"55",
		X"55",X"45",X"55",X"15",X"55",X"15",X"54",X"55",X"51",X"55",X"45",X"57",X"45",X"5D",X"15",X"5D",
		X"57",X"56",X"5D",X"59",X"75",X"59",X"D5",X"65",X"D5",X"95",X"55",X"95",X"56",X"55",X"59",X"55",
		X"95",X"55",X"95",X"55",X"95",X"55",X"95",X"55",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"80",X"01",X"80",X"00",X"80",X"00",X"80",X"00",
		X"15",X"55",X"15",X"55",X"15",X"55",X"15",X"55",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"55",X"00",X"15",X"00",X"15",X"00",X"05",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"54",X"55",X"51",X"55",X"45",X"55",X"15",X"54",X"55",X"51",X"55",X"45",X"55",X"15",X"55",
		X"55",X"55",X"55",X"55",X"55",X"57",X"55",X"5D",X"55",X"75",X"55",X"D5",X"57",X"55",X"5D",X"55",
		X"75",X"55",X"D5",X"56",X"55",X"59",X"55",X"59",X"55",X"65",X"55",X"95",X"56",X"55",X"59",X"55",
		X"95",X"54",X"55",X"51",X"55",X"51",X"55",X"45",X"55",X"15",X"54",X"55",X"54",X"55",X"51",X"55",
		X"55",X"75",X"55",X"D5",X"55",X"D5",X"57",X"55",X"5D",X"56",X"5D",X"56",X"75",X"59",X"D5",X"65",
		X"59",X"55",X"65",X"55",X"95",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"05",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"15",X"55",X"15",X"55",X"05",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"54",X"55",X"51",X"55",X"45",X"55",X"15",X"54",X"55",X"51",X"55",X"45",X"55",X"15",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"57",X"55",X"5D",X"55",X"75",X"55",X"D5",X"57",X"55",
		X"75",X"55",X"D5",X"55",X"D5",X"55",X"55",X"56",X"55",X"59",X"55",X"65",X"55",X"95",X"55",X"95",
		X"65",X"55",X"65",X"55",X"95",X"55",X"55",X"54",X"55",X"51",X"55",X"45",X"55",X"45",X"55",X"15",
		X"45",X"57",X"15",X"57",X"15",X"5D",X"55",X"75",X"55",X"75",X"55",X"D5",X"57",X"55",X"57",X"55",
		X"55",X"65",X"55",X"95",X"56",X"55",X"56",X"55",X"59",X"55",X"65",X"55",X"65",X"55",X"95",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"15",X"01",X"55",X"15",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"95",X"00",X"95",X"55",X"95",X"55",X"95",X"55",X"95",X"55",X"95",X"55",X"95",X"55",X"95",X"55",
		X"55",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"95",X"55",X"95",X"55",X"95",X"55",
		X"15",X"00",X"15",X"55",X"15",X"55",X"15",X"55",X"15",X"55",X"95",X"55",X"95",X"55",X"95",X"55",
		X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"55",X"05",X"55",X"15",X"55",X"55",X"55",X"55",X"55",
		X"01",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"54",X"00",X"55",X"50",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"40",X"00",X"54",X"00",X"55",X"40",X"55",X"50",X"55",X"54",X"55",X"55",
		X"05",X"55",X"01",X"55",X"01",X"55",X"00",X"55",X"00",X"55",X"00",X"15",X"00",X"15",X"00",X"05",
		X"55",X"54",X"55",X"51",X"55",X"45",X"55",X"15",X"54",X"55",X"51",X"55",X"45",X"55",X"15",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"57",X"55",X"5D",X"55",X"5D",X"55",X"75",X"55",X"D5",
		X"5D",X"55",X"75",X"55",X"D5",X"55",X"55",X"55",X"55",X"56",X"55",X"56",X"55",X"59",X"55",X"65",
		X"56",X"55",X"59",X"55",X"65",X"55",X"95",X"55",X"55",X"55",X"55",X"54",X"55",X"54",X"55",X"51",
		X"54",X"55",X"51",X"55",X"51",X"55",X"45",X"55",X"15",X"57",X"55",X"57",X"55",X"5D",X"55",X"75",
		X"5D",X"56",X"75",X"56",X"75",X"59",X"D5",X"59",X"55",X"65",X"55",X"95",X"55",X"95",X"56",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"15",X"55",X"01",X"55",X"00",X"15",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"55",
		X"55",X"55",X"15",X"55",X"05",X"55",X"01",X"55",X"00",X"15",X"00",X"01",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"05",X"55",X"00",X"15",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"40",
		X"55",X"55",X"55",X"55",X"55",X"54",X"55",X"50",X"55",X"00",X"50",X"00",X"00",X"00",X"00",X"00",
		X"00",X"05",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"15",X"55",X"15",X"55",X"05",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"57",X"55",X"5D",X"55",X"75",X"55",X"D5",
		X"57",X"55",X"5D",X"55",X"75",X"55",X"D5",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"55",X"59",
		X"55",X"95",X"56",X"55",X"59",X"55",X"59",X"55",X"65",X"55",X"95",X"55",X"55",X"55",X"55",X"55",
		X"55",X"45",X"55",X"15",X"55",X"15",X"54",X"55",X"51",X"55",X"45",X"55",X"45",X"55",X"15",X"55",
		X"55",X"D5",X"55",X"D5",X"57",X"55",X"5D",X"55",X"5D",X"55",X"75",X"56",X"D5",X"59",X"D5",X"59",
		X"59",X"55",X"59",X"55",X"65",X"55",X"95",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"05",X"55",X"01",X"55",X"01",X"55",X"00",X"55",X"00",X"55",X"00",X"15",X"00",X"15",X"00",X"05",
		X"55",X"D5",X"57",X"55",X"5D",X"55",X"75",X"55",X"D5",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"65",X"55",X"65",X"55",X"95",X"56",X"55",X"59",X"55",X"65",X"55",X"95",X"55",X"95",X"55",
		X"55",X"54",X"55",X"51",X"55",X"51",X"55",X"45",X"55",X"15",X"54",X"55",X"54",X"55",X"51",X"55",
		X"55",X"57",X"55",X"5D",X"55",X"5D",X"55",X"75",X"55",X"D5",X"57",X"55",X"57",X"55",X"5D",X"55",
		X"55",X"65",X"55",X"65",X"55",X"95",X"56",X"55",X"56",X"55",X"59",X"55",X"65",X"55",X"65",X"55",
		X"55",X"56",X"55",X"59",X"55",X"65",X"55",X"95",X"56",X"55",X"56",X"55",X"59",X"55",X"65",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"54",X"55",X"54",X"55",X"51",X"55",X"45",X"55",X"15",
		X"51",X"55",X"45",X"55",X"15",X"55",X"55",X"57",X"55",X"57",X"55",X"5D",X"55",X"75",X"55",X"75",
		X"75",X"55",X"75",X"56",X"D5",X"56",X"55",X"59",X"55",X"65",X"55",X"65",X"55",X"95",X"55",X"95",
		X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"54",X"55",X"51",
		X"55",X"15",X"54",X"55",X"51",X"55",X"45",X"55",X"45",X"55",X"15",X"55",X"55",X"55",X"55",X"57",
		X"55",X"D5",X"57",X"55",X"5D",X"55",X"5D",X"55",X"75",X"55",X"D5",X"55",X"D5",X"56",X"55",X"59",
		X"56",X"55",X"59",X"55",X"59",X"55",X"65",X"55",X"95",X"55",X"95",X"55",X"55",X"55",X"55",X"55",
		X"55",X"51",X"55",X"45",X"55",X"15",X"54",X"55",X"54",X"55",X"51",X"55",X"45",X"55",X"15",X"55",
		X"55",X"5D",X"55",X"5D",X"55",X"75",X"55",X"D5",X"55",X"D5",X"57",X"55",X"5D",X"55",X"75",X"55",
		X"55",X"59",X"55",X"65",X"55",X"95",X"55",X"95",X"56",X"55",X"56",X"55",X"59",X"55",X"65",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",
		X"55",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"15",X"55",X"55",X"55",X"55",X"57",X"55",X"57",X"55",X"5D",X"55",X"75",X"55",X"75",X"55",X"D5",
		X"75",X"55",X"D5",X"55",X"55",X"56",X"55",X"56",X"55",X"59",X"55",X"65",X"55",X"65",X"55",X"95",
		X"65",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"57",X"55",X"57",X"55",X"5D",X"55",X"75",X"55",X"D5",X"55",X"55",X"55",X"55",X"55",X"55",X"56",
		X"56",X"55",X"56",X"55",X"59",X"55",X"59",X"55",X"65",X"55",X"95",X"55",X"95",X"55",X"55",X"55",
		X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A5",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"40",
		X"55",X"59",X"55",X"59",X"55",X"65",X"55",X"95",X"55",X"95",X"56",X"55",X"59",X"55",X"59",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"55",
		X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"A5",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"40",
		X"65",X"55",X"65",X"55",X"95",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"55",X"01",X"55",X"05",X"55",
		X"00",X"01",X"00",X"55",X"05",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"A5",X"55",X"A5",X"55",X"A5",X"55",X"A5",X"55",X"A5",X"55",X"A5",X"55",X"A5",X"55",X"A5",X"55",
		X"05",X"55",X"05",X"55",X"05",X"55",X"05",X"55",X"05",X"55",X"05",X"55",X"05",X"55",X"05",X"55",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"05",X"00",X"05",X"00",X"15",X"00",X"15",X"00",X"55",
		X"15",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"A5",X"55",X"A5",X"55",X"A5",X"55",X"A5",X"55",X"A5",X"55",X"A5",X"55",X"A5",X"55",X"A5",X"55",
		X"05",X"55",X"05",X"55",X"05",X"55",X"05",X"55",X"05",X"55",X"05",X"55",X"05",X"55",X"05",X"55",
		X"50",X"00",X"40",X"00",X"40",X"01",X"00",X"05",X"00",X"05",X"00",X"15",X"00",X"15",X"00",X"55",
		X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"00",
		X"BF",X"FF",X"95",X"55",X"95",X"55",X"95",X"55",X"95",X"55",X"AA",X"AA",X"95",X"55",X"95",X"55",
		X"95",X"55",X"95",X"55",X"95",X"55",X"80",X"00",X"95",X"55",X"95",X"55",X"95",X"55",X"95",X"55",
		X"BF",X"FF",X"95",X"55",X"15",X"55",X"15",X"55",X"15",X"55",X"2A",X"AA",X"95",X"55",X"95",X"55",
		X"95",X"55",X"95",X"55",X"15",X"55",X"00",X"00",X"15",X"55",X"15",X"55",X"95",X"55",X"95",X"55",
		X"00",X"00",X"00",X"00",X"40",X"00",X"50",X"00",X"50",X"00",X"54",X"00",X"54",X"00",X"55",X"00",
		X"55",X"54",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"55",X"00",X"55",X"40",X"55",X"50",
		X"40",X"00",X"55",X"00",X"55",X"50",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"50",X"00",X"40",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"57",X"55",X"7F",X"D5",X"57",X"75",X"57",X"55",X"57",X"55",X"5D",X"D5",X"5D",X"D5",X"5D",X"75");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
