library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity popeye_sp_bits_1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of popeye_sp_bits_1 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"C0",X"00",X"E1",X"00",X"F1",X"00",X"F8",X"00",X"FC",X"00",X"F8",X"00",X"F0",
		X"0F",X"00",X"07",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"1F",X"00",X"1E",
		X"00",X"18",X"00",X"30",X"00",X"19",X"00",X"1B",X"00",X"3E",X"00",X"10",X"00",X"00",X"00",X"00",
		X"F0",X"E0",X"E0",X"3F",X"7F",X"7F",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"C0",X"80",X"80",X"00",X"00",
		X"00",X"00",X"00",X"01",X"03",X"03",X"07",X"07",X"07",X"87",X"C7",X"C7",X"E2",X"E0",X"E0",X"E0",
		X"E0",X"C0",X"F0",X"38",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"14",X"1E",X"3F",X"1F",X"0F",X"0F",X"0F",X"0E",
		X"0C",X"1C",X"18",X"38",X"30",X"70",X"60",X"60",X"E0",X"E0",X"70",X"70",X"20",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"17",X"3B",X"0F",X"0F",X"01",X"00",X"19",X"3E",X"3F",X"1F",X"0C",X"00",
		X"01",X"01",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"33",X"37",X"3F",X"3F",X"3F",X"FB",X"F1",X"F0",
		X"B0",X"B0",X"B0",X"A0",X"E0",X"E0",X"F0",X"F8",X"FE",X"FE",X"5E",X"5E",X"DF",X"7F",X"FF",X"FF",
		X"BF",X"7F",X"6E",X"DC",X"C0",X"00",X"00",X"FF",X"FF",X"1F",X"1F",X"3F",X"3F",X"7F",X"3F",X"1F",
		X"0F",X"0F",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"0E",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"07",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"80",X"C0",X"00",X"20",X"70",X"78",X"FC",X"FF",X"FF",X"F8",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"01",
		X"0D",X"0C",X"86",X"81",X"C0",X"40",X"00",X"07",X"23",X"1F",X"02",X"04",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"07",X"07",
		X"03",X"01",X"00",X"00",X"00",X"00",X"04",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"7C",X"FF",X"FF",X"F9",X"E0",X"00",X"00",X"00",X"40",X"40",X"40",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"BF",X"9F",X"8F",X"DE",
		X"BE",X"7F",X"7F",X"1F",X"7F",X"FF",X"FF",X"9F",X"7B",X"FB",X"E7",X"FF",X"7E",X"00",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"03",X"01",X"01",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"03",X"03",X"01",X"0F",X"1F",X"3F",X"3F",X"7F",X"7F",X"7F",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"38",X"70",X"FE",X"F1",X"FC",X"60",X"78",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"1F",X"DF",X"8F",X"CF",X"EF",
		X"FF",X"FF",X"87",X"03",X"01",X"01",X"01",X"01",X"C1",X"39",X"7D",X"FF",X"D4",X"34",X"38",X"1C",
		X"03",X"03",X"01",X"01",X"01",X"00",X"00",X"00",X"03",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"07",X"07",X"07",X"0F",X"1E",X"1F",X"1E",X"1F",X"0D",X"0E",X"03",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"60",X"20",X"80",X"E0",X"F0",X"F8",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"F0",X"C0",X"80",X"00",X"00",
		X"FF",X"0F",X"7F",X"FF",X"FF",X"FF",X"F8",X"F0",X"E1",X"E3",X"E3",X"E3",X"E3",X"E3",X"E3",X"E3",
		X"80",X"00",X"23",X"63",X"E3",X"E3",X"E1",X"71",X"11",X"01",X"F1",X"F0",X"F0",X"F8",X"F0",X"E0",
		X"C6",X"8F",X"9F",X"1F",X"3F",X"3F",X"3E",X"3E",X"1C",X"80",X"C1",X"FF",X"FF",X"FF",X"3F",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"07",X"07",X"07",
		X"0F",X"0F",X"0F",X"0F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"0F",X"0F",
		X"0F",X"07",X"07",X"07",X"03",X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"04",X"00",X"10",X"00",X"00",X"20",X"00",X"00",X"20",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"50",X"04",
		X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"20",X"00",X"08",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"04",X"04",X"04",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"08",X"08",X"00",X"00",X"10",X"20",X"40",X"40",X"80",X"80",X"80",X"80",X"00",X"00",
		X"00",X"00",X"30",X"30",X"30",X"30",X"30",X"F0",X"F0",X"30",X"30",X"30",X"F0",X"F0",X"00",X"00",
		X"00",X"01",X"03",X"07",X"07",X"07",X"07",X"06",X"06",X"06",X"FE",X"FE",X"06",X"06",X"FE",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"03",X"07",X"0F",X"1F",X"3F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"7C",X"38",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"7F",X"60",X"60",X"60",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"7F",X"7F",X"3F",X"1F",X"7F",X"7F",X"7F",X"3F",X"1F",X"7F",X"7F",X"7F",X"3F",X"1F",X"00",
		X"78",X"7C",X"60",X"60",X"60",X"61",X"61",X"60",X"60",X"60",X"60",X"60",X"60",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"1F",X"3F",X"7F",X"7F",X"7F",X"7C",X"3C",X"1E",X"0F",X"07",X"00",
		X"00",X"00",X"0C",X"0C",X"00",X"00",X"18",X"31",X"73",X"63",X"E3",X"E3",X"C3",X"C1",X"00",X"00",
		X"00",X"00",X"0F",X"0F",X"03",X"03",X"03",X"0F",X"0F",X"03",X"03",X"03",X"0F",X"0F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E3",X"E3",X"F3",X"FF",X"FF",X"FE",
		X"FF",X"FF",X"FF",X"E3",X"C0",X"E0",X"60",X"70",X"78",X"3C",X"3E",X"1F",X"07",X"01",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FC",X"F8",X"F0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"78",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CC",X"CC",X"CF",X"CF",X"0F",X"0F",
		X"CF",X"CF",X"0C",X"1C",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7E",X"7E",X"7E",X"7E",X"70",X"60",X"66",X"66",X"60",X"70",X"FF",X"FF",X"FF",X"FF",X"FE",X"F0",
		X"00",X"C0",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"0F",X"CF",X"CF",X"CF",X"CF",
		X"CF",X"CF",X"0C",X"1C",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3F",X"3F",X"3F",X"3F",X"38",X"30",X"33",X"33",X"30",X"38",X"FF",X"FF",X"BF",X"0F",X"01",X"00",
		X"00",X"F0",X"F8",X"7D",X"DE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"0F",X"CF",X"CF",X"0C",X"0C",X"CC",X"CC",X"0C",X"0C",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",
		X"FF",X"07",X"00",X"00",X"00",X"01",X"03",X"07",X"0F",X"1F",X"3F",X"7F",X"7F",X"7E",X"BC",X"F8",
		X"F8",X"F8",X"F8",X"F8",X"FC",X"FE",X"FF",X"FF",X"7F",X"7F",X"7F",X"3F",X"1F",X"1F",X"0F",X"17",
		X"1E",X"3E",X"3F",X"3F",X"1E",X"1E",X"1E",X"1E",X"1E",X"0E",X"0F",X"0F",X"07",X"00",X"00",X"00",
		X"FF",X"07",X"00",X"00",X"00",X"01",X"03",X"07",X"0F",X"1F",X"3F",X"7F",X"7E",X"7C",X"BC",X"FC",
		X"FC",X"FC",X"FC",X"FC",X"E0",X"E0",X"FC",X"FC",X"60",X"60",X"7F",X"3F",X"1F",X"1F",X"0F",X"17",
		X"00",X"E0",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"00",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"1F",X"1F",X"0F",X"01",X"00",
		X"20",X"99",X"83",X"C5",X"C1",X"6C",X"62",X"62",X"61",X"01",X"00",X"05",X"4D",X"26",X"16",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"0F",X"07",X"0F",X"07",X"00",
		X"00",X"01",X"03",X"05",X"0E",X"03",X"01",X"00",X"00",X"00",X"00",X"05",X"4D",X"26",X"16",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"A0",X"A0",X"A8",X"48",X"50",X"10",X"00",X"08",
		X"10",X"10",X"20",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"40",X"40",X"40",X"40",X"48",X"09",X"29",X"20",X"04",X"04",X"01",X"E3",X"E7",X"37",
		X"1D",X"1D",X"0F",X"0F",X"06",X"00",X"04",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"81",X"01",X"51",X"42",X"92",X"22",X"44",X"05",
		X"09",X"08",X"90",X"50",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"01",X"03",X"07",X"E7",X"FD",X"3D",X"0F",X"4F",
		X"06",X"22",X"04",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",
		X"00",X"C0",X"00",X"80",X"78",X"00",X"30",X"0F",X"00",X"80",X"7F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"01",X"03",X"07",X"E7",X"FD",X"3D",X"0F",X"0F",
		X"06",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"1C",X"20",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"47",X"C0",X"F8",X"77",X"3F",X"01",X"02",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"C0",X"60",X"60",X"70",X"30",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",
		X"10",X"08",X"00",X"04",X"84",X"89",X"92",X"84",X"80",X"88",X"82",X"80",X"80",X"80",X"80",X"40",
		X"30",X"78",X"F8",X"F8",X"F1",X"69",X"03",X"07",X"1F",X"FF",X"EB",X"D7",X"0B",X"1F",X"1D",X"09",
		X"01",X"01",X"81",X"01",X"81",X"81",X"81",X"81",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"3F",X"3F",X"1C",X"E0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"38",X"F8",X"D8",X"D9",X"DC",X"8C",X"8F",X"1F",X"3F",
		X"1E",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"E0",X"E0",X"E0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"03",X"03",X"01",X"00",
		X"00",X"00",X"00",X"00",X"17",X"3B",X"0F",X"0F",X"01",X"00",X"19",X"3E",X"3F",X"1F",X"0C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"3C",X"18",X"18",X"3C",X"FF",X"FF",X"FF",X"FF",
		X"01",X"01",X"01",X"03",X"02",X"02",X"02",X"01",X"06",X"04",X"08",X"00",X"00",X"01",X"1D",X"1C",
		X"1F",X"4F",X"76",X"7C",X"7E",X"63",X"07",X"1F",X"1F",X"1F",X"1E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"3C",X"18",X"18",X"3C",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C4",X"F0",X"F8",X"98",X"98",X"30",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"F0",X"F8",X"FC",X"FC",X"F8",X"78",X"90",X"E1",X"7B",X"BD",X"DC",X"EE",X"F2",X"FD",X"FE",
		X"F8",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"BF",X"DF",
		X"FF",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"38",X"60",X"7E",X"1F",X"03",X"00",X"40",X"60",X"10",X"0E",X"01",X"40",X"40",X"20",X"10",
		X"0E",X"01",X"40",X"40",X"60",X"38",X"1F",X"07",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EF",X"F7",X"FB",X"FB",X"FD",X"7D",X"DE",X"3E",X"2C",X"1C",X"08",X"18",X"58",X"68",X"EC",X"AC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"20",X"F0",X"F0",X"E0",X"80",X"80",
		X"00",X"78",X"7D",X"5E",X"5F",X"6F",X"EF",X"EF",X"E7",X"F3",X"F3",X"F3",X"F3",X"F9",X"F9",X"F9",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"23",X"47",X"47",X"13",X"21",X"41",
		X"1F",X"0F",X"0F",X"0F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"0F",X"1F",
		X"1F",X"1F",X"1F",X"FF",X"FF",X"FF",X"FF",X"EF",X"77",X"F7",X"77",X"17",X"37",X"77",X"37",X"3B",
		X"00",X"00",X"80",X"CF",X"DF",X"EF",X"EF",X"EF",X"E7",X"F3",X"F3",X"F3",X"F3",X"F9",X"F9",X"F9",
		X"F9",X"F9",X"F9",X"F9",X"F3",X"F3",X"F7",X"E7",X"EF",X"DF",X"DF",X"BF",X"3F",X"7E",X"F8",X"C0",
		X"00",X"00",X"F0",X"FC",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"6F",X"17",X"37",X"77",X"37",X"3B",
		X"7B",X"7B",X"F7",X"B7",X"6F",X"EF",X"9F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"0F",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"1F",X"1F",X"3F",X"7F",X"FF",X"E7",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"F8",X"FF",X"7F",X"3F",
		X"3E",X"3E",X"1D",X"1F",X"17",X"09",X"00",X"00",X"02",X"03",X"01",X"01",X"00",X"00",X"00",X"00",
		X"07",X"83",X"86",X"06",X"05",X"07",X"87",X"C5",X"43",X"41",X"00",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C7",X"8F",X"7F",X"FF",X"FF",X"FF",X"FC",X"BE",X"7D",X"7F",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"F0",
		X"98",X"CC",X"EC",X"F6",X"FA",X"FD",X"7E",X"BE",X"DF",X"DF",X"DF",X"FF",X"FF",X"FB",X"FD",X"FD",
		X"FE",X"FE",X"FE",X"FE",X"FC",X"F8",X"C0",X"80",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"E0",
		X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",X"F0",X"F0",X"E0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"C0",X"F0",X"1C",X"E7",X"F9",X"FE",X"FF",X"FF",
		X"1F",X"CF",X"E7",X"EF",X"FD",X"FE",X"FF",X"7F",X"FF",X"DF",X"EF",X"F7",X"FB",X"FD",X"FE",X"FE",
		X"FF",X"FF",X"BF",X"BF",X"5F",X"5F",X"DF",X"BF",X"7E",X"7C",X"F2",X"F3",X"EB",X"D7",X"F7",X"CF",
		X"BF",X"FF",X"FF",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"00",X"00",X"00",
		X"00",X"04",X"04",X"04",X"04",X"84",X"70",X"00",X"FF",X"FF",X"00",X"7F",X"FF",X"FF",X"FF",X"9F",
		X"7C",X"FF",X"FF",X"FF",X"FF",X"FF",X"E0",X"DE",X"FF",X"FF",X"FF",X"7F",X"3F",X"FF",X"02",X"FE",
		X"FD",X"FD",X"FD",X"FD",X"FC",X"BC",X"7C",X"7D",X"3F",X"AF",X"9E",X"9E",X"9D",X"1B",X"0F",X"0F",
		X"07",X"01",X"00",X"00",X"30",X"39",X"3F",X"1F",X"FF",X"FF",X"3F",X"FF",X"FF",X"EE",X"9C",X"0C",
		X"98",X"B8",X"B0",X"F0",X"FE",X"FE",X"FC",X"F8",X"F0",X"F8",X"F8",X"F9",X"FB",X"FB",X"F9",X"F9",
		X"F8",X"F3",X"F7",X"FB",X"FB",X"FB",X"FB",X"F7",X"EE",X"DE",X"BC",X"FC",X"FC",X"FF",X"FF",X"FE",
		X"FF",X"FF",X"7F",X"B6",X"01",X"39",X"4C",X"46",X"63",X"11",X"08",X"04",X"63",X"F3",X"70",X"A0",
		X"7D",X"5A",X"36",X"EC",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"01",X"01",X"00",X"00",
		X"01",X"05",X"05",X"07",X"07",X"07",X"03",X"03",X"03",X"03",X"07",X"07",X"07",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"1F",X"1F",X"1F",X"1F",X"1F",X"0F",X"07",X"07",X"07",X"03",X"03",X"01",X"01",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"0D",X"0B",X"07",X"05",X"04",
		X"04",X"06",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"F8",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"FF",X"DF",X"BF",X"FB",X"ED",X"0F",
		X"CF",X"EF",X"EF",X"FF",X"7F",X"BF",X"FF",X"FF",X"F3",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"04",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"03",X"03",X"03",
		X"3F",X"3F",X"1F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"07",X"4F",X"FF",X"FF",X"7F",X"3B",
		X"CB",X"FD",X"76",X"0F",X"3F",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"C0",X"F0",X"FC",X"FE",X"FC",X"F0",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"CF",
		X"00",X"00",X"00",X"01",X"07",X"0C",X"08",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"1F",X"1F",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"00",X"80",X"80",X"00",X"00",X"00",X"80",X"C0",X"40",X"40",X"00",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"02",X"02",X"02",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FE",X"FF",X"07",X"F1",X"FC",X"FE",X"FE",X"FE",X"0F",X"01",X"00",X"00",X"00",X"F8",X"07",
		X"00",X"00",X"00",X"00",X"F8",X"07",X"00",X"00",X"00",X"00",X"FC",X"FF",X"07",X"00",X"01",X"FF",
		X"7B",X"7B",X"FC",X"FF",X"EC",X"E9",X"DB",X"BC",X"7E",X"FF",X"F3",X"06",X"04",X"04",X"00",X"00",
		X"01",X"02",X"04",X"04",X"00",X"00",X"01",X"06",X"04",X"00",X"00",X"01",X"07",X"06",X"03",X"00",
		X"00",X"02",X"03",X"00",X"00",X"1F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"81",X"7E",
		X"F3",X"F8",X"FD",X"FE",X"FF",X"FF",X"1F",X"EF",X"F7",X"F7",X"F7",X"F7",X"F3",X"E5",X"ED",X"DD",
		X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"B7",X"9A",X"00",X"C0",
		X"B0",X"CC",X"7C",X"00",X"C4",X"EE",X"FE",X"D4",X"A8",X"00",X"90",X"F0",X"70",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"7F",X"FE",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"1D",
		X"81",X"7B",X"FF",X"FB",X"F7",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"F7",X"7B",X"7D",
		X"7B",X"7B",X"FC",X"FF",X"EF",X"EF",X"DF",X"BE",X"7E",X"FE",X"FE",X"70",X"00",X"0F",X"07",X"07",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"0B",X"0B",
		X"0B",X"0D",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3E",X"DE",X"EE",X"72",X"BC",X"FE",X"FF",X"FF",X"FE",X"FE",X"FC",X"1C",X"F0",X"EE",X"DF",X"BF",
		X"FF",X"FF",X"FF",X"FF",X"FE",X"FD",X"FD",X"FB",X"7B",X"7F",X"BF",X"BF",X"D7",X"C7",X"CF",X"87",
		X"37",X"6F",X"5F",X"7F",X"7F",X"5F",X"3F",X"17",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"BB",X"77",X"F7",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"EF",X"F7",X"FB",X"FD",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"DD",X"E4",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"03",X"03",X"07",X"07",X"07",X"07",X"07",X"07",
		X"07",X"07",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"1D",X"1A",X"17",X"1E",X"1D",X"0B",X"07",X"02",
		X"00",X"00",X"00",X"07",X"0F",X"1F",X"7F",X"FF",X"FF",X"FF",X"7F",X"8F",X"73",X"F5",X"EA",X"FD",
		X"DF",X"EF",X"FD",X"F9",X"F9",X"FF",X"FF",X"FF",X"F7",X"F3",X"F3",X"F3",X"67",X"67",X"67",X"4F",
		X"CF",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"F8",
		X"00",X"00",X"00",X"3E",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"7C",X"33",X"1F",X"3A",X"65",
		X"DE",X"DF",X"BF",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"FF",X"DF",X"DE",X"E9",X"E3",X"F7",X"FF",
		X"FF",X"FF",X"FF",X"BF",X"7F",X"3F",X"8E",X"9E",X"BE",X"1D",X"1D",X"3D",X"3D",X"7B",X"F7",X"E7",
		X"36",X"35",X"6D",X"7F",X"7F",X"7F",X"7F",X"7F",X"3F",X"3F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"3E",X"1F",X"1F",X"0F",X"0F",X"07",X"07",
		X"07",X"07",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"60",X"70",X"70",X"B8",X"AF",X"6F",X"6F",X"6F",X"EF",X"CF",X"DF",X"DF",X"9F",X"BF",X"BE",
		X"7D",X"63",X"0F",X"1F",X"03",X"09",X"09",X"04",X"04",X"04",X"04",X"04",X"04",X"08",X"08",X"30",
		X"00",X"00",X"00",X"01",X"1F",X"3F",X"7F",X"7F",X"00",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C7",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"CF",X"F1",X"FF",X"F5",X"F8",X"A3",X"C5",X"88",
		X"08",X"1E",X"23",X"20",X"00",X"11",X"3B",X"3F",X"13",X"0A",X"04",X"06",X"03",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"19",
		X"1F",X"1F",X"0F",X"1F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"1F",X"0F",X"FF",X"FF",X"3F",X"0F",
		X"1F",X"3B",X"73",X"63",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"7F",X"FF",X"FE",X"FC",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",
		X"00",X"00",X"08",X"0C",X"00",X"00",X"0F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"7F",X"0F",X"7D",
		X"00",X"00",X"00",X"00",X"00",X"08",X"01",X"07",X"0F",X"0F",X"3F",X"3F",X"3F",X"3F",X"0F",X"7D",
		X"00",X"00",X"00",X"80",X"E0",X"F0",X"F0",X"F0",X"E0",X"F8",X"FE",X"FF",X"FF",X"FF",X"FF",X"0F",
		X"1E",X"E6",X"F8",X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F3",X"E3",X"DB",X"FF",X"FF",X"FF",X"7F",X"3F",X"BF",X"DF",X"DE",X"EC",X"E0",X"E0",X"E0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"09",X"1C",X"1E",X"3F",X"3F",X"3F",X"3F",X"0F",X"7D",
		X"BB",X"77",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"02",X"0A",X"02",X"00",X"08",X"1D",X"1F",X"02",X"05",X"00",X"02",X"03",X"01",X"00",X"00",X"00",
		X"00",X"00",X"01",X"01",X"03",X"07",X"09",X"1E",X"16",X"1D",X"1B",X"06",X"05",X"03",X"00",X"00",
		X"00",X"00",X"00",X"08",X"0C",X"00",X"C0",X"E0",X"F0",X"FC",X"FC",X"FC",X"FF",X"FF",X"FF",X"0F",
		X"00",X"00",X"00",X"20",X"31",X"07",X"07",X"0F",X"3F",X"7F",X"7F",X"7F",X"3F",X"3F",X"0F",X"7D",
		X"00",X"80",X"C0",X"00",X"1E",X"7F",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"0F",
		X"1E",X"E6",X"F8",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"3E",X"BE",X"DC",X"DC",X"E8",X"E0",X"E0",X"E0",X"C0",
		X"00",X"00",X"10",X"38",X"78",X"FC",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"7D",
		X"BB",X"77",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"EF",X"F7",X"7B",X"7D",X"7E",X"BF",X"BF",X"FF",X"FF",X"3F",X"0D",X"00",X"00",X"00",
		X"00",X"01",X"0F",X"00",X"08",X"1D",X"1F",X"0A",X"05",X"00",X"02",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"E0",X"F0",X"F0",
		X"F0",X"F8",X"FA",X"FA",X"FA",X"F6",X"77",X"77",X"76",X"7E",X"7E",X"7C",X"3C",X"38",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"04",X"F0",X"FE",X"FF",X"FF",X"1F",X"EF",X"77",X"FB",
		X"FB",X"FD",X"FD",X"FE",X"FE",X"FE",X"FF",X"FD",X"FC",X"78",X"38",X"30",X"20",X"40",X"D0",X"D8",
		X"D8",X"3C",X"FE",X"CF",X"3F",X"7F",X"FF",X"FF",X"FE",X"FE",X"FC",X"F8",X"E0",X"C0",X"C0",X"80",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"07",X"00",X"03",X"03",X"03",X"01",X"00",X"00",X"00",X"00",
		X"01",X"03",X"07",X"0F",X"31",X"F1",X"F9",X"FC",X"00",X"00",X"F9",X"F1",X"F3",X"F3",X"C6",X"C7",
		X"C7",X"C0",X"E0",X"E0",X"E0",X"E0",X"DC",X"1F",X"0F",X"07",X"3F",X"7F",X"67",X"0F",X"1D",X"19",
		X"18",X"B8",X"F6",X"FE",X"FC",X"F8",X"FE",X"FF",X"FF",X"38",X"98",X"58",X"70",X"70",X"70",X"E0",
		X"E0",X"E0",X"F8",X"7C",X"78",X"7B",X"37",X"0F",X"00",X"00",X"00",X"3C",X"66",X"67",X"6F",X"77",
		X"C3",X"DB",X"FB",X"DB",X"9B",X"79",X"EF",X"BE",X"BF",X"9F",X"FA",X"60",X"A0",X"10",X"00",X"00",
		X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"01",X"01",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"03",X"01",X"01",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"03",X"01",X"03",X"03",X"05",X"2C",X"1F",X"07",X"0B",X"0B",X"05",X"02",X"01",X"00",X"00",X"00",
		X"07",X"0F",X"0C",X"0C",X"0F",X"07",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"79",X"F9",X"FF",X"FE",X"FD",X"FD",X"FB",
		X"FF",X"FF",X"FF",X"FF",X"7F",X"BE",X"41",X"7F",X"FF",X"FD",X"F4",X"E0",X"03",X"03",X"07",X"07",
		X"0C",X"37",X"7F",X"3F",X"3F",X"3F",X"3F",X"3B",X"1B",X"1F",X"0D",X"0F",X"07",X"00",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"3E",X"7F",X"FF",X"BF",X"9B",X"01",
		X"01",X"03",X"03",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"08",X"04",X"03",X"01",
		X"03",X"07",X"0F",X"0F",X"13",X"04",X"04",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"04",X"0C",X"18",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C7",X"CC",X"18",X"10",X"00",X"00",X"00",X"00",X"18",X"1C",X"0C",X"07",X"00",X"00",X"00",X"00",
		X"9E",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"1C",X"BC",X"EE",X"C8",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"20",X"31",X"33",X"06",X"04",X"00",X"00",X"07",X"06",X"06",X"03",X"01",X"00",
		X"E3",X"F3",X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"FC",X"38",X"30",X"20",X"20",
		X"1F",X"31",X"61",X"40",X"00",X"00",X"00",X"00",X"60",X"71",X"33",X"1E",X"00",X"00",X"00",X"00",
		X"EF",X"FF",X"71",X"60",X"60",X"60",X"60",X"60",X"60",X"71",X"7F",X"6F",X"60",X"60",X"70",X"40",
		X"00",X"00",X"00",X"00",X"78",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"70",X"F1",X"B9",X"23",
		X"3F",X"78",X"E0",X"E0",X"F0",X"F0",X"7C",X"3F",X"0F",X"03",X"00",X"00",X"40",X"60",X"71",X"3F",
		X"0F",X"18",X"18",X"18",X"1C",X"1F",X"0F",X"03",X"10",X"18",X"1C",X"0F",X"00",X"00",X"00",X"00",
		X"E0",X"30",X"38",X"18",X"18",X"18",X"F8",X"18",X"18",X"32",X"67",X"C7",X"00",X"00",X"00",X"00",
		X"BC",X"BC",X"EE",X"C6",X"86",X"86",X"86",X"86",X"86",X"86",X"C7",X"04",X"00",X"00",X"00",X"00",
		X"EF",X"F9",X"60",X"60",X"61",X"67",X"6F",X"78",X"60",X"61",X"73",X"3F",X"00",X"00",X"00",X"00",
		X"C0",X"60",X"70",X"30",X"30",X"30",X"F2",X"33",X"33",X"63",X"C2",X"90",X"18",X"18",X"0C",X"0F",
		X"01",X"03",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"05",X"07",X"06",
		X"F3",X"61",X"61",X"61",X"61",X"61",X"61",X"61",X"63",X"77",X"7D",X"39",X"00",X"00",X"00",X"00",
		X"FC",X"70",X"38",X"38",X"1C",X"0E",X"0E",X"07",X"07",X"03",X"06",X"06",X"0C",X"18",X"30",X"7C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7B",X"7F",X"7D",X"78",X"78",X"78",X"78",X"78",X"78",X"7D",X"7F",X"7B",X"78",X"78",X"78",X"78",
		X"CF",X"CF",X"CF",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"F0",X"F0",X"C0",X"C0",X"00",X"00",
		X"00",X"00",X"40",X"80",X"D8",X"D9",X"03",X"07",X"07",X"07",X"07",X"07",X"07",X"03",X"01",X"00",
		X"01",X"07",X"0F",X"1E",X"1E",X"3E",X"3E",X"00",X"00",X"3E",X"3E",X"1E",X"1E",X"0F",X"07",X"01",
		X"06",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"83",X"C3",X"E3",X"F3",X"F3",X"F3",X"F3",X"F3",X"F3",X"E3",X"C1",X"80",X"00",X"00",X"00",X"00",
		X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"1E",X"1E",X"1E",X"1E",
		X"EF",X"FF",X"F7",X"E3",X"E3",X"E3",X"E3",X"E3",X"E3",X"F7",X"FF",X"EF",X"00",X"00",X"00",X"00",
		X"F0",X"B8",X"1C",X"1E",X"1E",X"1E",X"1E",X"1E",X"1E",X"1C",X"B8",X"F0",X"00",X"00",X"00",X"00",
		X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"7C",X"FC",X"FC",X"BC",X"3C",X"00",X"00",X"00",X"00",
		X"07",X"87",X"C7",X"E7",X"E7",X"E7",X"E7",X"E7",X"E7",X"C7",X"87",X"03",X"00",X"00",X"00",X"00",
		X"7B",X"7B",X"79",X"79",X"78",X"78",X"78",X"78",X"F8",X"F8",X"78",X"78",X"00",X"00",X"00",X"00",
		X"3E",X"3E",X"3C",X"FC",X"F8",X"78",X"78",X"F0",X"F0",X"E0",X"E0",X"E0",X"C0",X"C0",X"80",X"80",
		X"E0",X"E1",X"E3",X"E7",X"E7",X"E7",X"E7",X"E7",X"E7",X"E3",X"F9",X"F8",X"E0",X"E0",X"C0",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"87",X"C7",X"E7",X"E7",X"E7",X"E7",X"E7",X"E7",X"C7",X"87",X"07",X"07",X"07",X"07",X"07",
		X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3E",X"3F",X"1F",X"0E",X"00",X"00",X"00",X"00",
		X"3E",X"77",X"E3",X"E3",X"E3",X"03",X"FF",X"FF",X"E3",X"E3",X"77",X"3E",X"00",X"00",X"00",X"00",
		X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3E",X"1F",X"DF",X"CE",X"00",X"00",X"00",X"00",
		X"E7",X"E7",X"E7",X"E7",X"E7",X"E7",X"E7",X"E7",X"E7",X"E7",X"E7",X"07",X"07",X"E7",X"E7",X"E7",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"06",X"0E",X"0E",X"1E",
		X"0E",X"86",X"C0",X"E0",X"F0",X"F0",X"E0",X"C0",X"C0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"03",X"0F",X"3F",X"63",X"9B",X"7F",X"FF",X"F3",X"C3",X"83",X"03",X"03",X"03",X"03",X"83",
		X"03",X"03",X"03",X"0F",X"0F",X"03",X"03",X"07",X"0E",X"0C",X"0C",X"0C",X"0C",X"06",X"02",X"00",
		X"00",X"02",X"06",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"06",X"02",X"00",X"00",X"02",X"06",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"0D",X"08",X"0D",X"0F",X"1E",X"3E",X"33",X"31",X"31",X"39",X"3F",X"1F",X"1F",X"0F",X"07",
		X"F1",X"F3",X"67",X"6D",X"DC",X"F8",X"71",X"3B",X"1E",X"4C",X"8C",X"18",X"00",X"21",X"61",X"00",
		X"00",X"00",X"C0",X"F0",X"F8",X"F8",X"F7",X"FF",X"FF",X"EF",X"E0",X"E0",X"C0",X"C4",X"8C",X"8C",
		X"44",X"44",X"8B",X"8A",X"17",X"17",X"20",X"20",X"40",X"A0",X"F0",X"E0",X"F0",X"F0",X"E0",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"DC",X"7C",X"3C",X"18",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"F0",X"F8",X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",X"F8",X"FC",X"FC",X"FC",X"FC",
		X"00",X"00",X"03",X"02",X"07",X"07",X"00",X"00",X"00",X"A0",X"F0",X"E0",X"F0",X"F0",X"E0",X"80",
		X"00",X"00",X"80",X"DC",X"DE",X"CE",X"C4",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"01",X"07",
		X"00",X"00",X"03",X"03",X"01",X"01",X"03",X"01",X"01",X"03",X"03",X"01",X"00",X"00",X"00",X"00",
		X"07",X"0E",X"0C",X"1C",X"18",X"18",X"18",X"10",X"10",X"D0",X"F0",X"F0",X"6A",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"C7",X"EE",X"FC",X"3C",X"0E",X"07",
		X"C2",X"F0",X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"40",X"40",X"00",X"20",X"20",X"20",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"01",X"01",X"01",X"01",X"01",X"03",X"03",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"0F",X"FF",X"FD",X"1C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"F0",X"F0",X"F8",X"F8",X"F8",
		X"C0",X"F9",X"F8",X"F8",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"F8",X"F0",X"60",X"60",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"06",X"1C",X"78",X"F0",X"E0",X"C0",
		X"00",X"40",X"02",X"0C",X"00",X"02",X"06",X"0C",X"1C",X"19",X"3B",X"37",X"3F",X"7F",X"7B",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"F8",X"3C",X"7C",X"FE",X"DF",X"B3",X"30",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"78",X"7C",X"30",X"30",
		X"C0",X"F1",X"FB",X"FB",X"FD",X"FC",X"FC",X"FE",X"FE",X"FE",X"FE",X"FE",X"FC",X"F8",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"03",X"03",X"07",X"06",X"07",X"06",X"05",X"04",X"34",X"3C",X"3C",X"1A",X"00",X"00",X"00",
		X"7C",X"FE",X"D4",X"00",X"30",X"38",X"0D",X"01",X"09",X"10",X"12",X"77",X"E6",X"E1",X"60",X"00",
		X"07",X"0F",X"0E",X"0C",X"00",X"18",X"78",X"FF",X"FE",X"FE",X"FE",X"EE",X"47",X"6F",X"3F",X"1F",
		X"00",X"00",X"01",X"03",X"03",X"1B",X"78",X"FF",X"FE",X"FE",X"FE",X"EE",X"47",X"6F",X"3F",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"40",X"20",X"00",X"00",X"B0",X"FC",X"84",X"7A",X"7D",X"B2",X"30",
		X"C0",X"F0",X"FB",X"FB",X"FD",X"FC",X"FC",X"FC",X"FC",X"FC",X"F8",X"F0",X"E0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"00",X"00",X"60",X"60",X"FC",X"F8",X"F8",X"08",X"00",
		X"00",X"F8",X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"61",X"00",X"00",X"00",
		X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"0C",X"18",X"F8",X"FC",X"1E",
		X"00",X"00",X"C0",X"F0",X"F8",X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"18",X"3C",X"06",X"7B",X"7E",X"30",
		X"C0",X"F0",X"FB",X"FB",X"F9",X"FC",X"FC",X"FC",X"FC",X"FC",X"F8",X"F0",X"E0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"FC",X"C4",X"BA",X"7D",X"FA",X"30",
		X"C0",X"F0",X"FA",X"FB",X"F9",X"FC",X"FC",X"FC",X"FC",X"FC",X"F8",X"F0",X"E0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"F8",X"7C",X"3C",X"18",X"18",X"10",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"F8",X"1F",X"0F",X"07",
		X"C3",X"E3",X"F1",X"F8",X"F8",X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"FF",
		X"60",X"19",X"00",X"00",X"00",X"20",X"00",X"00",X"08",X"00",X"00",X"03",X"03",X"06",X"03",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"03",X"06",X"06",X"07",X"07",X"06",X"06",X"06",X"07",X"07",X"06",X"06",X"07",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"03",X"06",X"06",X"07",X"07",X"06",X"06",X"06",X"FE",X"FE",X"06",X"06",X"FE",X"FE",
		X"FF",X"FF",X"FF",X"FF",X"FC",X"F1",X"63",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",
		X"FF",X"FE",X"00",X"83",X"83",X"81",X"89",X"8D",X"8D",X"89",X"81",X"C3",X"E7",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",
		X"0F",X"07",X"07",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"07",X"C0",X"FE",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"E0",X"01",X"0F",X"FF",X"FF",
		X"F8",X"C0",X"00",X"00",X"01",X"01",X"03",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"1C",X"EC",X"F4",X"F8",X"FC",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"81",X"E3",X"FB",X"FC",X"FF",X"FF",X"FF",X"FE",X"7E",X"3D",X"3B",X"7F",X"7F",X"7F",X"7F",X"FF",
		X"07",X"1F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FD",X"FC",X"0C",X"F0",X"FE",X"FF",X"FF",X"FF",X"FF",
		X"FB",X"C7",X"DF",X"DF",X"BE",X"7E",X"DE",X"EC",X"F0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"80",X"C0",X"40",X"C0",X"00",X"80",X"80",X"C0",X"F0",X"E0",X"80",X"40",X"C0",X"80",X"00",X"00",
		X"FF",X"FF",X"FF",X"1F",X"E3",X"FD",X"FE",X"FF",X"FF",X"FE",X"FE",X"FC",X"FC",X"FC",X"FC",X"F8",
		X"88",X"20",X"7C",X"4C",X"4B",X"9B",X"97",X"97",X"37",X"2F",X"27",X"C1",X"C1",X"E0",X"F0",X"F8",
		X"F8",X"F8",X"F8",X"80",X"7C",X"FE",X"E0",X"DC",X"B8",X"70",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"40",X"61",X"01",X"03",X"07",X"0F",X"0F",X"1F",X"1F",X"1F",X"1F",X"0F",X"00",X"00",
		X"00",X"00",X"40",X"81",X"CD",X"FD",X"FB",X"FB",X"3B",X"1B",X"0B",X"00",X"00",X"00",X"01",X"07",
		X"07",X"0B",X"1B",X"3F",X"3F",X"3C",X"3B",X"17",X"07",X"03",X"00",X"00",X"04",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"17",X"3B",X"7B",X"63",X"FB",X"F1",X"47",X"EF",X"EF",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"06",X"06",
		X"17",X"73",X"FB",X"FB",X"FB",X"F9",X"F9",X"FC",X"FC",X"FC",X"FD",X"F9",X"E9",X"C3",X"83",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"C0",X"80",X"84",X"88",X"80",X"C0",X"00",X"00",X"00",X"80",X"C0",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"7C",X"FC",X"FC",X"F4",
		X"E4",X"40",X"03",X"07",X"06",X"0C",X"38",X"3F",X"0F",X"0F",X"0F",X"1F",X"3F",X"3F",X"0F",X"03",
		X"10",X"18",X"80",X"00",X"80",X"00",X"00",X"00",X"10",X"48",X"E8",X"E0",X"E0",X"60",X"60",X"70",
		X"30",X"B8",X"BD",X"9D",X"DD",X"D8",X"D8",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"E0",
		X"C0",X"C0",X"42",X"04",X"00",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1C",X"0E",X"07",X"3F",X"7E",X"F0",X"60",X"00",X"00",X"0C",X"0F",X"07",X"07",X"07",X"0F",X"0F",
		X"0F",X"1F",X"3F",X"1F",X"1F",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"03",X"1F",X"3E",X"7C",X"F8",X"E3",X"DF",X"BE",X"3A",X"13",X"01",X"00",X"00",X"81",X"00",
		X"F0",X"F0",X"F9",X"FB",X"EF",X"DF",X"FB",X"7D",X"9C",X"E8",X"20",X"D0",X"50",X"70",X"6C",X"F4",
		X"F8",X"70",X"F0",X"F0",X"52",X"BE",X"F4",X"E8",X"D8",X"B0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"61",X"03",X"03",X"01",X"01",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",
		X"00",X"02",X"03",X"03",X"03",X"03",X"01",X"01",X"03",X"03",X"07",X"07",X"17",X"19",X"1F",X"1E",
		X"3C",X"78",X"78",X"F8",X"7C",X"7E",X"7F",X"7F",X"3F",X"3F",X"1F",X"1F",X"0F",X"07",X"01",X"00",
		X"00",X"00",X"00",X"3E",X"7C",X"FC",X"F8",X"FE",X"FF",X"FC",X"F3",X"6F",X"1B",X"0F",X"3F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"3F",X"FD",X"F0",X"E0",X"C0",X"00",X"00",X"C0",X"A0",X"E0",
		X"80",X"C0",X"C0",X"C0",X"F4",X"DC",X"9C",X"38",X"30",X"68",X"D8",X"B0",X"60",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"78",X"A0",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"02",X"03",X"03",X"07",X"07",
		X"07",X"03",X"03",X"01",X"01",X"01",X"00",X"81",X"FF",X"FF",X"FF",X"81",X"03",X"07",X"0F",X"0F",
		X"17",X"3C",X"3B",X"17",X"07",X"06",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"7F",X"7F",X"7F",X"FF",X"FF",X"CF",X"5B",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"7C",X"5E",X"FF",X"FF",X"FF",X"FE",X"1C",X"E8",X"F0",
		X"D8",X"E8",X"F0",X"F8",X"F8",X"FC",X"FC",X"FC",X"FF",X"DF",X"EB",X"F3",X"67",X"7F",X"7F",X"F2",
		X"F2",X"64",X"CC",X"8C",X"1C",X"FC",X"FC",X"EC",X"70",X"79",X"F9",X"B9",X"7B",X"F3",X"FF",X"F7",
		X"EF",X"E7",X"66",X"E3",X"E3",X"E1",X"E0",X"70",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"04",X"05",X"09",X"0B",
		X"13",X"17",X"E7",X"07",X"0F",X"0E",X"1E",X"1E",X"1C",X"08",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"20",X"10",X"08",X"08",X"08",X"C8",X"E8",X"E8",X"EE",X"F3",X"8F",
		X"FF",X"FF",X"0F",X"F3",X"FD",X"FE",X"FF",X"FF",X"FE",X"FE",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"0C",X"00",X"70",X"4D",X"4B",X"8B",X"95",X"96",X"16",X"2C",X"28",X"C0",X"C0",X"E0",X"F0",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"0F",X"1F",X"1F",X"37",X"2F",X"6F",X"5E",X"1E",X"4E",X"7C",X"FC",X"F8",X"FC",X"71",X"3B",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"01",X"00",X"02",X"0F",X"1F",X"3F",X"E7",X"FB",X"FD",X"FF",
		X"FF",X"0F",X"F3",X"FD",X"FE",X"BF",X"FF",X"FF",X"7F",X"BE",X"FE",X"7C",X"7C",X"FC",X"FC",X"F8",
		X"C8",X"C0",X"30",X"4C",X"48",X"88",X"90",X"90",X"10",X"28",X"20",X"C0",X"C0",X"E0",X"F0",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"06",X"0E",X"0E",X"0D",X"05",X"06",X"03",X"01",X"00",X"00",X"00",X"01",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"8F",X"1F",X"1F",X"3E",X"3E",X"E7",X"FB",X"FB",X"FF",X"FF",
		X"FF",X"3F",X"C7",X"F9",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F9",X"F8",
		X"09",X"01",X"70",X"4D",X"4B",X"8A",X"94",X"94",X"10",X"28",X"20",X"C0",X"C0",X"E0",X"F0",X"F8",
		X"F8",X"F8",X"F8",X"80",X"7D",X"FE",X"E0",X"DC",X"B0",X"70",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"07",X"07",X"0F",X"0B",X"0D",X"07",X"02",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",
		X"03",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"F0",X"E0",X"E1",X"00",X"F0",X"FC",X"FC",X"FE",X"08",
		X"F2",X"FD",X"FE",X"FF",X"FF",X"FF",X"FE",X"FE",X"FC",X"FC",X"F8",X"F8",X"78",X"B8",X"D8",X"D8",
		X"D8",X"AC",X"76",X"F7",X"FF",X"7C",X"18",X"80",X"C0",X"80",X"80",X"F0",X"F8",X"7C",X"7B",X"2D",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"07",X"07",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"07",X"0F",
		X"0E",X"1A",X"19",X"1C",X"3F",X"3F",X"3F",X"3F",X"1D",X"0E",X"06",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FC",X"38",X"C0",X"E0",X"D8",X"E8",X"F0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"9F",X"BF",X"7F",X"FF",X"FF",X"FF",
		X"0E",X"F3",X"FD",X"FE",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"FF",X"7F",X"FF",X"FF",X"FF",X"F7",
		X"F7",X"F4",X"2F",X"9B",X"BC",X"FC",X"78",X"18",X"80",X"C0",X"80",X"80",X"F0",X"B8",X"DC",X"5B",
		X"00",X"00",X"00",X"00",X"00",X"40",X"61",X"07",X"1E",X"1E",X"1E",X"BF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"06",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"1F",X"E3",X"FD",X"FE",X"FF",X"FF",X"EF",X"FE",X"CE",X"9E",X"AF",X"F7",X"FF",X"FF",X"EF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"BE",X"EF",X"F7",X"FB",X"FD",X"FE",X"0F",
		X"F3",X"FD",X"FE",X"FF",X"FF",X"FF",X"FE",X"FE",X"FC",X"FC",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"D8",X"E8",X"F7",X"FE",X"FF",X"7B",X"1D",X"80",X"C0",X"80",X"80",X"F0",X"F8",X"7C",X"7B",X"2D",
		X"AF",X"EC",X"DE",X"FE",X"FE",X"DC",X"5E",X"BE",X"FF",X"F1",X"CE",X"7C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"38",X"7C",X"7E",
		X"FA",X"FE",X"FD",X"FD",X"FC",X"FC",X"7C",X"7C",X"78",X"2C",X"D6",X"DE",X"64",X"7C",X"18",X"00",
		X"01",X"03",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"CF",X"F3",X"FD",X"FD",X"FE",X"FE",
		X"0F",X"F3",X"FD",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FD",X"F8",X"F8",X"F8",X"F8",X"F9",
		X"FB",X"F7",X"EF",X"DB",X"FD",X"FC",X"78",X"18",X"80",X"C0",X"80",X"80",X"F0",X"B8",X"DC",X"5B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"18",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"0F",X"1F",X"1F",
		X"3F",X"0E",X"72",X"6E",X"6E",X"72",X"3E",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"1E",X"37",X"29",X"36",
		X"00",X"00",X"00",X"00",X"00",X"40",X"60",X"00",X"04",X"0E",X"1F",X"3F",X"47",X"3B",X"FD",X"FF",
		X"FF",X"0F",X"F3",X"FD",X"FE",X"FF",X"FF",X"EF",X"FE",X"CE",X"9E",X"AF",X"F7",X"FF",X"FF",X"EF",
		X"DE",X"D6",X"D9",X"DF",X"AE",X"B0",X"F8",X"78",X"18",X"80",X"C0",X"80",X"80",X"F8",X"BC",X"5B",
		X"DD",X"BF",X"FC",X"FE",X"7E",X"7E",X"DC",X"5E",X"BE",X"FF",X"F1",X"CE",X"7C",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"1E",X"37",X"29",X"36",
		X"37",X"0B",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"03",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
