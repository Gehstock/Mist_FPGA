library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity tron_bg_bits_2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of tron_bg_bits_2 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"00",X"07",X"00",X"05",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",
		X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"07",X"00",X"07",X"00",X"0D",
		X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",
		X"00",X"0D",X"00",X"0C",X"00",X"07",X"00",X"0F",X"00",X"0F",X"00",X"0D",X"00",X"07",X"00",X"0F",
		X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0D",X"00",X"07",
		X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"05",X"00",X"0F",X"00",X"0F",X"00",X"0F",
		X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"05",X"00",X"0F",X"00",X"05",X"00",X"0F",X"00",X"0F",
		X"00",X"0F",X"00",X"0F",X"00",X"07",X"00",X"0D",X"00",X"0F",X"00",X"07",X"00",X"0D",X"00",X"07",
		X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"07",X"00",X"0F",
		X"7F",X"FF",X"DF",X"55",X"7F",X"7F",X"7F",X"7D",X"DF",X"7D",X"DF",X"7D",X"DF",X"7D",X"F7",X"DD",
		X"FD",X"F7",X"FD",X"F7",X"FD",X"F5",X"F5",X"F7",X"DD",X"F7",X"7D",X"F7",X"7D",X"DF",X"7D",X"DF",
		X"FF",X"FF",X"55",X"5F",X"FF",X"DF",X"55",X"5F",X"FF",X"FF",X"FF",X"FF",X"D5",X"7F",X"DF",X"7F",
		X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"AA",X"AA",
		X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",
		X"7F",X"5D",X"7D",X"DD",X"77",X"DD",X"77",X"DD",X"5F",X"DD",X"7F",X"DD",X"7F",X"DD",X"7F",X"DD",
		X"75",X"55",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"55",X"57",X"7F",X"F7",X"7F",X"F7",X"7F",X"F7",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",
		X"F5",X"55",X"F7",X"FF",X"F7",X"FF",X"F7",X"FF",X"F7",X"FF",X"F7",X"FF",X"F7",X"FF",X"F7",X"FF",
		X"FD",X"FD",X"FD",X"F7",X"FF",X"5F",X"FF",X"FD",X"57",X"F7",X"F7",X"FD",X"F7",X"FF",X"FD",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"DF",X"FF",X"F7",X"FF",X"F7",X"FF",
		X"FF",X"FF",X"FF",X"FD",X"FF",X"F7",X"FF",X"DF",X"FF",X"DF",X"FF",X"DD",X"F7",X"F7",X"F7",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"55",X"FF",X"7F",X"FF",X"7F",X"FF",X"75",X"FF",X"57",X"FF",X"FF",
		X"FD",X"F7",X"F7",X"FD",X"F3",X"FF",X"DF",X"FF",X"DF",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F7",X"FF",X"F7",X"FF",X"DF",X"FF",X"DF",X"FF",X"DF",X"FF",X"DF",X"FF",X"F5",X"55",X"FF",X"FF",
		X"FF",X"FF",X"D5",X"55",X"DF",X"FF",X"DF",X"F5",X"DF",X"DF",X"DF",X"F7",X"DF",X"FD",X"F7",X"FF",
		X"D5",X"77",X"FF",X"77",X"FF",X"77",X"FF",X"77",X"FF",X"77",X"FF",X"77",X"55",X"7D",X"FF",X"FF",
		X"FF",X"77",X"FF",X"77",X"FF",X"77",X"D5",X"77",X"DF",X"F7",X"DF",X"F7",X"DF",X"F7",X"DF",X"F7",
		X"F7",X"DF",X"FD",X"F7",X"7D",X"F7",X"DF",X"7D",X"F7",X"DF",X"FD",X"F7",X"FF",X"77",X"FF",X"77",
		X"F7",X"FD",X"DF",X"F7",X"7F",X"DF",X"FF",X"DF",X"FF",X"F7",X"D7",X"FD",X"7D",X"FF",X"DF",X"7F",
		X"F7",X"FF",X"F7",X"FF",X"F7",X"FF",X"F5",X"FF",X"DD",X"FF",X"7D",X"F5",X"FD",X"DF",X"FD",X"7F",
		X"FF",X"77",X"FF",X"7D",X"FF",X"5F",X"FF",X"77",X"FF",X"7D",X"D5",X"7F",X"DF",X"FF",X"DF",X"FF",
		X"55",X"55",X"FF",X"FF",X"FF",X"FF",X"FD",X"55",X"5F",X"7F",X"77",X"DF",X"7D",X"F7",X"7F",X"7D",
		X"55",X"55",X"FF",X"FF",X"55",X"55",X"FF",X"FF",X"55",X"55",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"F5",X"FF",X"5F",X"D5",X"FF",X"7F",X"FF",X"FF",X"55",X"FD",X"FF",
		X"55",X"55",X"FF",X"FF",X"55",X"55",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"55",
		X"55",X"F7",X"FF",X"DF",X"55",X"7D",X"FF",X"F7",X"55",X"5F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"57",X"FF",X"FF",X"FF",X"55",X"FF",X"FF",X"7F",X"FF",X"DF",X"FF",X"7F",X"FD",X"FF",X"57",X"FF",
		X"FF",X"F7",X"FF",X"FD",X"55",X"57",X"FF",X"FF",X"FF",X"FF",X"FD",X"55",X"FD",X"FD",X"FD",X"F7",
		X"F7",X"7F",X"F7",X"7F",X"77",X"7F",X"D7",X"DF",X"FF",X"DF",X"FF",X"DF",X"57",X"F7",X"F7",X"F7",
		X"FF",X"F7",X"FF",X"DF",X"55",X"7F",X"FF",X"FD",X"55",X"7D",X"FF",X"77",X"FD",X"F7",X"F7",X"DF",
		X"7F",X"DD",X"DF",X"DD",X"F7",X"DD",X"3D",X"DD",X"CF",X"5D",X"F3",X"FD",X"F3",X"FD",X"FC",X"FD",
		X"55",X"55",X"FF",X"FD",X"55",X"5D",X"FF",X"DD",X"FF",X"DD",X"FF",X"DD",X"FF",X"DD",X"FF",X"DD",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"55",X"55",X"FF",X"FF",X"55",X"55",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"F7",X"FD",X"57",X"FD",X"FF",X"FD",X"55",X"FF",X"FF",X"55",X"55",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"DF",X"FF",X"F7",X"FF",X"F7",X"FF",X"F7",X"FF",X"FD",X"FF",X"FD",X"FF",X"F7",X"FF",X"F7",
		X"DF",X"FD",X"DF",X"FD",X"DF",X"FD",X"DD",X"55",X"DD",X"FF",X"DD",X"55",X"DF",X"FF",X"DF",X"FF",
		X"DF",X"F7",X"FF",X"DF",X"FF",X"7F",X"FF",X"7F",X"FD",X"FD",X"F7",X"F7",X"5F",X"F7",X"FF",X"F7",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DD",X"DF",X"DD",X"DF",X"DD",X"F7",X"DF",X"77",X"F7",X"77",X"77",X"7D",X"F7",X"DD",X"FD",X"DF",
		X"DF",X"F7",X"DF",X"F7",X"DF",X"F7",X"DF",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",X"FD",X"FD",
		X"DF",X"FD",X"7F",X"F7",X"7F",X"F7",X"FF",X"DF",X"FF",X"DF",X"FF",X"7F",X"FF",X"7F",X"FF",X"7F",
		X"DF",X"DF",X"DF",X"DF",X"DF",X"DF",X"DF",X"DF",X"DF",X"DF",X"DF",X"DF",X"DF",X"DF",X"DF",X"F7",
		X"DF",X"DF",X"DF",X"DF",X"DF",X"DF",X"DF",X"DF",X"D7",X"DF",X"DD",X"DF",X"DF",X"5F",X"DF",X"DF",
		X"DF",X"FF",X"F7",X"FF",X"FD",X"FF",X"57",X"FF",X"FF",X"FF",X"5F",X"D5",X"DF",X"DF",X"DF",X"DF",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"5D",X"DD",X"FD",X"D7",X"55",X"DF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DF",X"FF",X"DD",X"55",X"DD",X"FF",X"DD",X"D5",X"DD",X"DF",X"DD",X"DF",X"DD",X"DF",X"DD",X"DD",
		X"DD",X"F7",X"DD",X"F7",X"DD",X"F7",X"DD",X"F7",X"DD",X"F7",X"5D",X"F7",X"FD",X"F7",X"FD",X"F7",
		X"F7",X"7D",X"F7",X"7F",X"F7",X"7F",X"F7",X"55",X"F7",X"FF",X"F7",X"55",X"77",X"7F",X"D7",X"7F",
		X"FF",X"7F",X"FF",X"DF",X"FF",X"F7",X"FF",X"DF",X"FF",X"7F",X"FF",X"7D",X"FD",X"FD",X"FD",X"F7",
		X"FF",X"F7",X"55",X"57",X"FF",X"FF",X"57",X"FF",X"F7",X"FF",X"DF",X"FF",X"7F",X"FF",X"FF",X"FF",
		X"55",X"7D",X"FF",X"77",X"FF",X"77",X"57",X"77",X"F7",X"77",X"77",X"77",X"77",X"77",X"77",X"77",
		X"DF",X"D7",X"F5",X"FD",X"FF",X"5F",X"FF",X"F5",X"5F",X"FF",X"F7",X"FF",X"FD",X"7F",X"FF",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",
		X"FD",X"DD",X"FD",X"DD",X"F7",X"DF",X"DF",X"DF",X"DF",X"7F",X"DD",X"FF",X"DD",X"FF",X"DD",X"FF",
		X"F7",X"77",X"F7",X"77",X"F7",X"77",X"F7",X"77",X"F7",X"77",X"F7",X"77",X"DF",X"77",X"7F",X"77",
		X"FF",X"FF",X"7F",X"FF",X"D7",X"FF",X"FD",X"7F",X"7F",X"DF",X"D7",X"F5",X"FD",X"7F",X"FF",X"D7",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"3D",X"75",X"CD",X"75",X"F3",X"DF",X"5C",X"35",X"5C",X"35",X"F7",X"CF",X"DD",X"73",X"7D",X"7C",
		X"FD",X"FF",X"FD",X"7D",X"F7",X"DD",X"DF",X"F7",X"7F",X"DD",X"FF",X"7D",X"FD",X"F7",X"F7",X"DF",
		X"7F",X"7F",X"DF",X"DF",X"F7",X"F7",X"F7",X"F7",X"7D",X"FD",X"DF",X"77",X"F7",X"DF",X"FD",X"5F",
		X"FD",X"7F",X"F5",X"DF",X"DF",X"77",X"7F",X"DD",X"DF",X"DF",X"F7",X"F7",X"F7",X"FD",X"FD",X"FF",
		X"DD",X"F7",X"DD",X"DD",X"7D",X"DD",X"7D",X"DD",X"55",X"DD",X"FF",X"DD",X"FD",X"5D",X"FD",X"FD",
		X"FF",X"7D",X"FF",X"7D",X"FF",X"D7",X"F7",X"FF",X"DD",X"FF",X"DD",X"FF",X"DD",X"FF",X"DD",X"FF",
		X"FD",X"FD",X"FD",X"FD",X"D7",X"FD",X"DF",X"FD",X"DF",X"FD",X"DF",X"FD",X"DF",X"FD",X"D5",X"7D",
		X"F7",X"F7",X"DF",X"DF",X"7F",X"7F",X"FF",X"7F",X"FD",X"F7",X"F7",X"DD",X"F7",X"DD",X"DF",X"7D",
		X"F7",X"5F",X"F7",X"7D",X"F7",X"F7",X"F7",X"DF",X"F7",X"DF",X"F7",X"7F",X"D7",X"7F",X"7F",X"7F",
		X"FD",X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",X"55",X"FF",X"FD",X"FD",X"55",X"FD",X"F7",X"FD",X"F7",
		X"77",X"FD",X"77",X"FF",X"77",X"FF",X"77",X"FF",X"77",X"FF",X"77",X"D5",X"77",X"DF",X"77",X"DF",
		X"F7",X"F7",X"F7",X"FD",X"F7",X"FF",X"F7",X"FF",X"F7",X"FD",X"F5",X"F7",X"F7",X"77",X"F7",X"DF",
		X"FF",X"CF",X"7F",X"CF",X"7F",X"F3",X"7F",X"FC",X"7F",X"FC",X"7F",X"FC",X"7F",X"FC",X"FF",X"FC",
		X"FF",X"77",X"FF",X"D7",X"5F",X"F7",X"F7",X"FF",X"FD",X"FF",X"7F",X"7F",X"DF",X"DF",X"F7",X"F7",
		X"FF",X"7F",X"FF",X"7F",X"FF",X"7F",X"FF",X"7F",X"FF",X"7F",X"FD",X"5F",X"F7",X"FF",X"FD",X"FF",
		X"55",X"57",X"FF",X"FF",X"FF",X"FD",X"55",X"57",X"FF",X"FF",X"FF",X"FF",X"55",X"55",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"F5",X"55",X"DF",X"FF",X"7F",X"FF",X"FF",X"55",X"FD",X"FF",X"F7",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"55",X"57",X"FF",X"FF",X"FF",X"FF",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FD",X"5F",X"FF",X"F5",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"D5",X"FF",X"FF",X"57",X"FF",X"FD",
		X"FD",X"FD",X"FD",X"F7",X"7D",X"F7",X"D5",X"DF",X"FF",X"F5",X"55",X"FF",X"FF",X"57",X"FF",X"FD",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"5D",X"DF",X"FD",X"DF",X"FD",X"DF",X"FD",
		X"FF",X"7F",X"FF",X"7F",X"03",X"7F",X"F3",X"77",X"F3",X"75",X"F3",X"77",X"F3",X"77",X"F3",X"77",
		X"DF",X"FD",X"DF",X"F7",X"DF",X"F7",X"DF",X"DF",X"DF",X"7F",X"DF",X"7D",X"DD",X"F7",X"D7",X"F7",
		X"77",X"7D",X"DF",X"7D",X"FF",X"7D",X"FF",X"77",X"5F",X"77",X"77",X"77",X"77",X"5F",X"77",X"7F",
		X"DD",X"FF",X"DD",X"FF",X"DD",X"FF",X"DD",X"FF",X"DD",X"FF",X"DD",X"FF",X"DD",X"FF",X"DD",X"FF",
		X"FF",X"DD",X"FF",X"77",X"FD",X"DF",X"F5",X"DF",X"DF",X"7F",X"7D",X"FF",X"55",X"55",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"55",X"55",X"FF",X"FF",X"FF",X"FF",X"55",X"55",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FD",X"DC",X"FD",X"DC",X"FD",X"DC",X"FD",X"DC",X"FD",X"DC",X"5D",X"DC",X"F5",X"DF",X"FF",X"D7",
		X"7F",X"37",X"DF",X"37",X"F7",X"3D",X"F7",X"3F",X"F7",X"00",X"F7",X"FC",X"F7",X"FC",X"FD",X"FC",
		X"FF",X"7F",X"FF",X"7F",X"FF",X"55",X"FF",X"FF",X"FF",X"FF",X"FD",X"55",X"F7",X"FF",X"DF",X"55",
		X"DF",X"77",X"DF",X"77",X"DF",X"77",X"DF",X"77",X"DF",X"77",X"DF",X"77",X"DF",X"77",X"DF",X"77",
		X"73",X"7D",X"73",X"7D",X"73",X"7D",X"73",X"7D",X"73",X"7D",X"73",X"7D",X"73",X"75",X"F3",X"5D",
		X"CD",X"F7",X"F1",X"DD",X"F3",X"7D",X"FC",X"7D",X"FF",X"DF",X"FF",X"DF",X"FF",X"F7",X"FF",X"F7",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FD",X"DF",X"FD",X"DF",X"FD",X"DF",X"FD",X"DF",X"FD",X"D5",X"FD",X"FF",X"3D",X"FF",X"3D",X"FF",
		X"FF",X"FF",X"FF",X"DF",X"7F",X"77",X"DF",X"77",X"F7",X"77",X"F7",X"77",X"F7",X"77",X"F7",X"77",
		X"FF",X"FF",X"FF",X"FF",X"55",X"55",X"FF",X"FF",X"FF",X"FF",X"55",X"55",X"FF",X"FF",X"57",X"FD",
		X"77",X"7F",X"77",X"7F",X"77",X"7F",X"77",X"7F",X"77",X"7F",X"77",X"DF",X"77",X"F7",X"77",X"FD",
		X"FF",X"7F",X"FF",X"DF",X"FF",X"F7",X"FF",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"7F",X"FF",X"DF",X"FF",X"DF",X"FF",
		X"FD",X"FF",X"F7",X"7F",X"F7",X"DF",X"DF",X"F7",X"7F",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DF",X"DF",X"DF",X"DF",X"7F",X"7F",X"7F",X"7F",X"FD",X"FF",X"FD",X"FF",X"F7",X"FF",X"F7",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"55",X"FD",X"FD",X"F7",X"F7",X"F7",X"F7",X"DF",
		X"D7",X"F7",X"FD",X"77",X"FF",X"D7",X"FF",X"FF",X"F5",X"7F",X"DF",X"DF",X"77",X"F7",X"75",X"FD",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DF",X"F7",X"DF",X"DF",X"5F",X"DF",X"FF",X"7F",X"FF",X"7F",X"55",X"FF",X"FD",X"FF",X"57",X"FF",
		X"FF",X"7F",X"FF",X"7F",X"7F",X"7F",X"DF",X"7F",X"F7",X"75",X"F7",X"77",X"F7",X"77",X"F7",X"77",
		X"F7",X"7F",X"F7",X"75",X"F7",X"77",X"F7",X"77",X"57",X"77",X"FF",X"7D",X"FF",X"7F",X"FF",X"7F",
		X"DF",X"FF",X"DF",X"FF",X"DF",X"F5",X"DF",X"F7",X"DF",X"57",X"F7",X"7F",X"F7",X"7F",X"F7",X"7F",
		X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",X"DF",X"F7",X"DF",X"F7",X"DF",X"F7",X"DF",X"F7",X"DF",X"F5",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"75",X"55",X"77",X"FF",X"77",X"FF",X"77",X"FF",
		X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",X"FF",X"FD",X"5D",X"5D",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"FF",X"F7",X"FF",X"F7",X"FD",X"F5",X"D7",X"7F",X"DF",X"7F",X"DF",X"55",X"DF",X"FF",X"DF",X"FF",
		X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",X"FD",X"F7",X"FD",X"F7",X"FF",X"77",X"FF",X"77",X"FF",X"77",
		X"FF",X"77",X"FF",X"77",X"FF",X"77",X"55",X"77",X"FF",X"F7",X"FF",X"F7",X"55",X"57",X"FF",X"FF",
		X"FD",X"F7",X"FD",X"F7",X"FD",X"F7",X"FD",X"F7",X"FD",X"F7",X"FD",X"F7",X"F7",X"77",X"DF",X"77",
		X"DD",X"F7",X"DD",X"F7",X"DD",X"F7",X"DD",X"F7",X"7D",X"F7",X"7D",X"F7",X"FD",X"F7",X"FD",X"F7",
		X"7F",X"F7",X"7F",X"F7",X"7F",X"F5",X"7F",X"F7",X"7F",X"DF",X"7F",X"7F",X"75",X"FF",X"5F",X"FF",
		X"FF",X"7F",X"FF",X"7F",X"FF",X"7F",X"FF",X"DF",X"FF",X"DF",X"FF",X"DF",X"FF",X"F7",X"FF",X"F7",
		X"FF",X"F7",X"FF",X"F7",X"FF",X"D7",X"FF",X"77",X"F5",X"F7",X"DF",X"F7",X"7F",X"F7",X"7F",X"F7",
		X"FF",X"77",X"FF",X"77",X"FF",X"77",X"FF",X"77",X"FD",X"57",X"F7",X"7F",X"DF",X"75",X"7D",X"F7",
		X"5F",X"77",X"DF",X"77",X"DF",X"77",X"7F",X"77",X"FF",X"77",X"FF",X"77",X"FF",X"77",X"FF",X"77",
		X"FF",X"7D",X"FF",X"7D",X"FF",X"7F",X"FF",X"7F",X"FF",X"7F",X"FF",X"75",X"FF",X"75",X"FF",X"77",
		X"FF",X"F7",X"FF",X"77",X"FD",X"77",X"F7",X"77",X"DF",X"77",X"DF",X"77",X"7F",X"77",X"FF",X"77",
		X"F7",X"FF",X"FD",X"FF",X"7F",X"7F",X"DF",X"DF",X"F7",X"F7",X"FD",X"FD",X"FF",X"7F",X"FF",X"D5",
		X"5F",X"FF",X"DF",X"FF",X"D5",X"55",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"55",X"55",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"F5",X"FF",X"5F",X"F5",X"FF",X"5F",X"FF",X"D7",X"FF",X"FD",X"FF",
		X"FF",X"FF",X"FD",X"55",X"57",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"55",X"55",
		X"FF",X"F7",X"FF",X"5F",X"FD",X"FF",X"57",X"FD",X"FF",X"F7",X"FF",X"DF",X"FF",X"7F",X"55",X"FF",
		X"D7",X"DD",X"DD",X"F7",X"DD",X"FF",X"DF",X"7F",X"DF",X"7F",X"DF",X"DF",X"DF",X"F7",X"5F",X"FD",
		X"FD",X"FF",X"55",X"FF",X"FF",X"FF",X"FF",X"FF",X"55",X"55",X"FF",X"FF",X"55",X"55",X"F7",X"FF",
		X"FD",X"7F",X"FD",X"FF",X"FF",X"7F",X"FF",X"7F",X"5F",X"DF",X"DF",X"F7",X"F7",X"F5",X"FD",X"FD",
		X"DF",X"FD",X"7F",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"55",X"55",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"00",X"F0",X"00",X"FC",X"00",X"FF",X"00",X"FF",X"C0",X"FF",X"F0",X"FF",X"FC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"00",X"FF",X"C0",X"FF",X"C0",X"FF",X"F0",X"FF",X"F0",X"FF",X"FC",X"FF",X"FC",X"FF",X"FF",
		X"00",X"00",X"C0",X"00",X"C0",X"00",X"F0",X"00",X"F0",X"00",X"FC",X"00",X"FC",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"FF",X"00",X"FF",X"F0",
		X"00",X"00",X"00",X"00",X"C0",X"00",X"FF",X"00",X"FF",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FC",X"00",X"FF",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",
		X"FE",X"BF",X"FE",X"BF",X"FE",X"BF",X"FE",X"BF",X"FE",X"BF",X"FE",X"BF",X"FE",X"BF",X"FE",X"BF",
		X"FE",X"BF",X"FE",X"BF",X"FE",X"BF",X"AA",X"BF",X"AA",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FC",X"3F",X"FC",X"3F",X"FC",X"3F",X"FC",X"3F",X"FC",X"3F",X"FC",X"3F",X"FC",X"3F",X"FC",X"3F",
		X"FC",X"3F",X"FC",X"3F",X"FC",X"3F",X"00",X"3F",X"00",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"15",X"55",X"00",X"00",
		X"15",X"55",X"15",X"55",X"15",X"55",X"15",X"55",X"15",X"55",X"15",X"55",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"FF",X"57",X"FF",X"57",X"FF",X"5F",X"FF",X"5F",X"FF",X"7F",X"FF",X"7F",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"55",X"00",X"55",X"00",
		X"00",X"15",X"00",X"55",X"00",X"55",X"01",X"55",X"01",X"55",X"05",X"55",X"05",X"55",X"15",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"15",X"00",X"15",X"00",X"15",
		X"00",X"00",X"00",X"03",X"00",X"0F",X"00",X"3F",X"00",X"FF",X"03",X"FF",X"0F",X"FF",X"3F",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"00",X"0F",X"00",X"3F",X"00",X"FF",X"03",X"FF",X"0F",X"FF",X"3F",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"54",X"00",X"54",X"00",X"50",X"00",X"40",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"40",X"55",X"40",X"55",X"40",X"55",X"40",X"55",X"40",X"55",X"00",X"55",X"00",X"55",X"00",
		X"00",X"00",X"00",X"03",X"00",X"0F",X"00",X"3F",X"00",X"FF",X"03",X"FF",X"0F",X"FF",X"3F",X"FF",
		X"FF",X"FB",X"FF",X"FB",X"FF",X"FB",X"FF",X"FB",X"FF",X"FB",X"FF",X"FB",X"FF",X"FB",X"AA",X"AB",
		X"FF",X"FB",X"FF",X"FB",X"FF",X"FB",X"FF",X"FB",X"FF",X"FB",X"FF",X"FB",X"FF",X"FB",X"FF",X"FB",
		X"FF",X"FF",X"FF",X"FF",X"AA",X"AB",X"FF",X"FB",X"FF",X"FB",X"FF",X"FB",X"FF",X"FB",X"FF",X"FB",
		X"FF",X"FF",X"FF",X"FF",X"AA",X"BF",X"FF",X"BF",X"FF",X"EF",X"FF",X"EF",X"FF",X"FB",X"FF",X"FE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",X"EF",X"FF",X"BF",X"BF",X"BF",X"EA",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"AA",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"AF",X"FF",X"FA",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"EA",X"FF",X"EF",X"FF",X"EF",X"FF",X"EF",X"FF",X"AF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"AA",X"EB",X"FF",X"BF",X"FF",X"FF",X"FF",
		X"FE",X"AF",X"FB",X"FF",X"EF",X"FF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FB",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"FF",X"EF",X"FF",X"FA",X"AF",
		X"FB",X"FF",X"EF",X"FF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",X"EF",X"FF",X"BF",X"FE",X"FF",
		X"FF",X"EF",X"FF",X"FB",X"FF",X"FB",X"FF",X"FE",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"EF",X"FF",X"EF",X"FF",X"FB",X"FF",X"FB",X"FF",X"FE",X"FF",X"FE",X"FF",X"FF",X"BF",X"FF",X"BF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FA",X"AF",X"EF",X"FF",X"BF",X"FF",X"BF",X"FF",
		X"FF",X"FA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"BF",X"FF",X"BF",X"FF",X"BF",X"FF",X"BF",X"FF",X"BF",X"FF",X"BF",X"FF",X"BF",X"FF",X"BF",X"FF",
		X"FF",X"FA",X"FE",X"A0",X"F8",X"0F",X"E3",X"FF",X"8F",X"FF",X"BF",X"FF",X"BF",X"FF",X"BF",X"FF",
		X"FF",X"FA",X"FE",X"A0",X"F8",X"00",X"E0",X"00",X"80",X"00",X"80",X"03",X"BF",X"FF",X"BF",X"FF",
		X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",
		X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",
		X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"05",X"55",X"05",X"55",X"05",X"55",X"05",X"55",X"05",X"55",X"05",X"55",X"05",X"55",X"05",X"55",
		X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",
		X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"05",X"55",X"05",X"55",X"05",X"55",X"05",X"55",X"05",X"55",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"C0",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",
		X"C5",X"55",X"C5",X"55",X"C5",X"55",X"C5",X"55",X"C5",X"55",X"C5",X"55",X"C5",X"55",X"00",X"00",
		X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"FF",X"FC",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FC",X"FF",X"FC",
		X"C5",X"00",X"C4",X"00",X"C0",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"05",X"55",X"05",X"55",
		X"C5",X"55",X"C5",X"55",X"C5",X"55",X"C5",X"54",X"C5",X"50",X"C5",X"50",X"C5",X"40",X"C5",X"00",
		X"C0",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FC",X"FF",X"FC",X"FF",X"F0",X"FF",X"C0",X"FF",X"00",X"FC",X"00",X"FC",X"00",X"F0",X"00",
		X"00",X"3C",X"00",X"3C",X"00",X"FC",X"03",X"FC",X"0F",X"FC",X"0F",X"FC",X"FF",X"FC",X"FF",X"FC",
		X"FF",X"00",X"FC",X"00",X"F0",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"00",X"00",X"C0",X"00",X"30",X"00",X"0C",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"05",X"55",X"05",X"55",X"05",X"55",X"05",X"55",X"05",X"55",X"05",X"50",X"05",X"00",X"00",X"00",
		X"05",X"55",X"05",X"55",X"FD",X"55",X"03",X"D5",X"00",X"F5",X"00",X"35",X"00",X"0D",X"00",X"0D",
		X"00",X"0D",X"00",X"0D",X"00",X"35",X"00",X"F5",X"00",X"D5",X"01",X"55",X"05",X"55",X"05",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"F0",X"00",X"FC",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"C0",X"FF",X"C0",X"FF",X"F0",X"FF",X"F0",X"FF",X"F0",X"FF",X"FC",X"FF",X"FC",
		X"05",X"55",X"05",X"55",X"05",X"55",X"05",X"55",X"05",X"55",X"05",X"55",X"05",X"55",X"00",X"00",
		X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",
		X"C0",X"00",X"C0",X"00",X"30",X"00",X"30",X"00",X"30",X"00",X"0C",X"00",X"0C",X"00",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"00",X"00",X"C0",X"00",X"30",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"30",X"00",X"30",X"00",X"C0",X"03",X"00",X"0C",X"00",X"30",X"00",X"F0",X"00",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"0C",
		X"C0",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"05",X"55",X"05",X"55",X"05",X"55",X"05",X"55",X"05",X"55",X"05",X"55",X"05",X"55",
		X"05",X"55",X"05",X"55",X"05",X"54",X"C5",X"50",X"C5",X"50",X"C5",X"40",X"C5",X"00",X"C4",X"00",
		X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"0C",X"00",X"30",X"00",X"30",
		X"00",X"C0",X"03",X"00",X"0C",X"00",X"30",X"00",X"30",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"55",X"05",X"55",
		X"00",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"F0",X"FF",X"F0",X"FF",X"C0",X"FF",X"00",X"FC",X"00",X"F0",X"00",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"AA",X"AA",
		X"80",X"00",X"20",X"00",X"08",X"00",X"02",X"00",X"00",X"80",X"00",X"20",X"00",X"08",X"00",X"02",
		X"80",X"02",X"20",X"08",X"08",X"20",X"02",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",
		X"AA",X"00",X"82",X"00",X"82",X"00",X"82",X"00",X"82",X"00",X"82",X"00",X"82",X"00",X"82",X"00",
		X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"20",X"00",X"08",X"00",X"02",X"AA",
		X"82",X"AA",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"AA",X"AA",
		X"00",X"80",X"00",X"80",X"00",X"80",X"02",X"00",X"02",X"00",X"02",X"00",X"08",X"00",X"08",X"00",
		X"80",X"00",X"20",X"00",X"08",X"00",X"02",X"00",X"00",X"80",X"00",X"20",X"00",X"08",X"00",X"02",
		X"00",X"02",X"00",X"0A",X"00",X"22",X"00",X"82",X"02",X"02",X"08",X"02",X"20",X"02",X"80",X"02",
		X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",
		X"AA",X"AA",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",
		X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",
		X"80",X"00",X"20",X"00",X"08",X"00",X"02",X"00",X"00",X"80",X"00",X"20",X"00",X"08",X"00",X"02",
		X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",X"80",X"02",
		X"08",X"00",X"20",X"00",X"80",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"28",X"02",X"80",X"A8",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"00",X"05",X"00",X"15",X"00",X"55",X"00",X"55",X"01",X"55",X"05",X"55",X"05",X"55",
		X"00",X"03",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"55",X"05",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"BF",X"FE",X"BF",X"FE",X"BF",X"FE",X"AA",X"FE",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FC",X"3F",X"FC",X"3F",X"FC",X"3F",X"FC",X"00",X"FC",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"AA",X"AA",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"BF",X"FE",X"BF",X"FE",X"BF",X"FE",X"BF",X"FE",X"BF",X"FE",X"BF",X"FE",X"BF",X"FE",X"BF",
		X"FC",X"3F",X"FC",X"3F",X"FC",X"3F",X"FC",X"3F",X"FC",X"3F",X"FC",X"3F",X"FC",X"3F",X"FC",X"3F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"AA",X"FE",X"AA",X"FE",X"BF",X"FE",X"BF",X"FE",X"BF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"00",X"FC",X"00",X"FC",X"3F",X"FC",X"3F",X"FC",X"3F",
		X"FE",X"BF",X"FE",X"BF",X"FE",X"BF",X"AA",X"BF",X"AA",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FC",X"3F",X"FC",X"3F",X"FC",X"3F",X"00",X"3F",X"00",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"03",X"03",X"0C",X"3F",X"FF",X"F0",X"FF",X"F0",X"0C",X"3F",X"03",X"03",X"00",X"00",
		X"00",X"EA",X"00",X"EA",X"00",X"EA",X"00",X"EA",X"00",X"EA",X"00",X"EA",X"00",X"E8",X"00",X"00",
		X"00",X"30",X"00",X"30",X"00",X"30",X"00",X"FF",X"00",X"FA",X"00",X"3A",X"00",X"0E",X"00",X"03",
		X"EA",X"AA",X"3A",X"A9",X"0E",X"A5",X"03",X"95",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"AA",X"3A",X"AA",X"EA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"0E",X"00",X"3A",X"00",X"EA",X"03",X"AA",
		X"AA",X"A8",X"AA",X"A4",X"AA",X"94",X"AA",X"94",X"AA",X"54",X"A9",X"54",X"A5",X"54",X"95",X"54",
		X"3A",X"AA",X"EA",X"AA",X"EA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"3A",X"00",X"EA",X"00",X"EA",X"FF",X"AA",X"03",X"AA",X"FF",X"AA",X"0E",X"AA",X"0E",X"AA",
		X"00",X"03",X"00",X"03",X"00",X"0E",X"FF",X"FE",X"00",X"0E",X"FF",X"FE",X"00",X"3A",X"00",X"3A",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"03",
		X"EF",X"FE",X"EB",X"FA",X"EA",X"EA",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A9",X"55",X"A9",X"55",X"A5",X"55",X"A5",X"55",X"95",X"55",X"95",X"55",X"55",X"55",X"55",X"55",
		X"AA",X"A4",X"AA",X"A4",X"AA",X"A4",X"AA",X"94",X"AA",X"94",X"AA",X"94",X"AA",X"54",X"AA",X"54",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A9",X"AA",X"A9",X"AA",X"A9",X"AA",X"A9",X"AA",X"A5",
		X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"EA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",
		X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"FF",X"C0",X"00",X"C0",
		X"30",X"03",X"0C",X"03",X"03",X"0C",X"C0",X"CC",X"B0",X"30",X"AC",X"00",X"AB",X"00",X"AA",X"C0",
		X"03",X"00",X"03",X"00",X"0C",X"00",X"0F",X"FF",X"30",X"00",X"3F",X"FF",X"C0",X"00",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"30",X"00",X"30",X"00",X"30",X"FF",X"FF",X"00",X"30",X"FF",X"FF",X"00",X"30",X"00",X"30",
		X"AC",X"30",X"AB",X"0C",X"AB",X"0C",X"AA",X"C3",X"AA",X"C3",X"AA",X"C0",X"AA",X"B0",X"AA",X"B0",
		X"C3",X"00",X"C3",X"00",X"B3",X"00",X"B0",X"C0",X"B0",X"C0",X"B0",X"C0",X"AC",X"30",X"AC",X"30",
		X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"03",X"00",X"C3",X"00",X"C3",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",
		X"00",X"30",X"00",X"30",X"00",X"30",X"00",X"30",X"00",X"30",X"00",X"30",X"00",X"30",X"00",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"30",X"00",X"30",X"00",X"30",X"00",X"30",X"00",X"30",X"00",X"30",X"00",X"30",X"00",X"30",
		X"00",X"30",X"00",X"30",X"00",X"30",X"FF",X"FF",X"00",X"30",X"FF",X"FF",X"00",X"30",X"00",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"C0",X"00",X"30",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"2A",X"AA",X"2A",X"AA",X"0A",X"AA",X"0A",X"AA",X"0A",X"AA",X"02",X"AA",X"00",X"AA",X"00",X"2A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"54",X"55",X"54",X"55",X"50",X"55",X"40",X"55",X"00",X"54",X"00",X"50",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"05",X"55",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"15",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"05",X"55",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"05",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"55",X"55",X"55",X"55",X"55",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"05",X"55",X"05",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",
		X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"50",X"05",X"50",X"00",X"00",X"00",X"00",
		X"50",X"05",X"50",X"05",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"05",X"55",X"05",X"55",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",
		X"00",X"00",X"00",X"00",X"50",X"05",X"50",X"05",X"50",X"05",X"50",X"05",X"50",X"05",X"50",X"05",
		X"05",X"05",X"05",X"05",X"05",X"00",X"05",X"00",X"05",X"50",X"05",X"50",X"00",X"00",X"00",X"00",
		X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"55",X"00",X"55",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"55",X"05",X"55",X"05",X"05",X"05",X"05",
		X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"05",X"00",X"05",
		X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"55",X"05",X"55",X"00",X"00",X"00",X"00",
		X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"55",X"00",X"55",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"55",X"05",X"55",X"05",X"00",X"05",X"00",
		X"00",X"00",X"00",X"00",X"05",X"00",X"05",X"00",X"55",X"55",X"55",X"55",X"05",X"55",X"05",X"55",
		X"50",X"05",X"50",X"05",X"50",X"05",X"50",X"05",X"50",X"55",X"50",X"55",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",
		X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"50",X"05",X"50",X"05",
		X"50",X"05",X"50",X"05",X"50",X"05",X"50",X"05",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",
		X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",
		X"05",X"00",X"05",X"00",X"05",X"55",X"05",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"50",X"05",X"50",X"05",X"50",X"05",X"50",X"05",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"55",X"05",X"55",X"05",X"00",X"05",X"00",
		X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"00",X"50",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"05",X"55",X"05",X"55",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"00",
		X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"50",X"00",X"50",X"00",
		X"00",X"05",X"00",X"05",X"00",X"05",X"00",X"05",X"55",X"55",X"55",X"55",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",X"05",X"55",X"05",X"55",X"00",X"05",X"00",X"05",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"FF",X"00",X"FF",X"F0",
		X"00",X"00",X"00",X"00",X"C0",X"00",X"FF",X"00",X"FF",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FC",X"00",X"FF",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"00",
		X"FE",X"BF",X"FE",X"BF",X"FE",X"BF",X"FE",X"BF",X"FE",X"BF",X"FE",X"BF",X"FE",X"BF",X"FE",X"BF",
		X"FE",X"BF",X"FE",X"BF",X"FE",X"BF",X"AA",X"BF",X"AA",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FC",X"3F",X"FC",X"3F",X"FC",X"3F",X"FC",X"3F",X"FC",X"3F",X"FC",X"3F",X"FC",X"3F",X"FC",X"3F",
		X"FC",X"3F",X"FC",X"3F",X"FC",X"3F",X"00",X"3F",X"00",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"15",X"55",X"00",X"00",
		X"15",X"55",X"15",X"55",X"15",X"55",X"15",X"55",X"15",X"55",X"15",X"55",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"FF",X"57",X"FF",X"57",X"FF",X"5F",X"FF",X"5F",X"FF",X"7F",X"FF",X"7F",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"55",X"00",X"55",X"00",
		X"00",X"15",X"00",X"55",X"00",X"55",X"01",X"55",X"01",X"55",X"05",X"55",X"05",X"55",X"15",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"15",X"00",X"15",X"00",X"15",
		X"00",X"00",X"00",X"03",X"00",X"0F",X"00",X"3F",X"00",X"FF",X"03",X"FF",X"0F",X"FF",X"3F",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"00",X"0F",X"00",X"3F",X"00",X"FF",X"03",X"FF",X"0F",X"FF",X"3F",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"54",X"00",X"54",X"00",X"50",X"00",X"40",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"40",X"55",X"40",X"55",X"40",X"55",X"40",X"55",X"40",X"55",X"00",X"55",X"00",X"55",X"00",
		X"00",X"00",X"00",X"03",X"00",X"0F",X"00",X"3F",X"00",X"FF",X"03",X"FF",X"0F",X"FF",X"3F",X"FF",
		X"FF",X"FB",X"FF",X"FB",X"FF",X"FB",X"FF",X"FB",X"FF",X"FB",X"FF",X"FB",X"FF",X"FB",X"AA",X"AB",
		X"FF",X"FB",X"FF",X"FB",X"FF",X"FB",X"FF",X"FB",X"FF",X"FB",X"FF",X"FB",X"FF",X"FB",X"FF",X"FB",
		X"FF",X"FF",X"FF",X"FF",X"AA",X"AB",X"FF",X"FB",X"FF",X"FB",X"FF",X"FB",X"FF",X"FB",X"FF",X"FB",
		X"FF",X"FF",X"FF",X"FF",X"AA",X"BF",X"FF",X"BF",X"FF",X"EF",X"FF",X"EF",X"FF",X"FB",X"FF",X"FE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",X"EF",X"FF",X"BF",X"BF",X"BF",X"EA",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"AA",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"AF",X"FF",X"FA",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"EA",X"FF",X"EF",X"FF",X"EF",X"FF",X"EF",X"FF",X"AF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"AA",X"EB",X"FF",X"BF",X"FF",X"FF",X"FF",
		X"FE",X"AF",X"FB",X"FF",X"EF",X"FF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FB",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"FF",X"EF",X"FF",X"FA",X"AF",
		X"FB",X"FF",X"EF",X"FF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",X"EF",X"FF",X"BF",X"FE",X"FF",
		X"FF",X"EF",X"FF",X"FB",X"FF",X"FB",X"FF",X"FE",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"EF",X"FF",X"EF",X"FF",X"FB",X"FF",X"FB",X"FF",X"FE",X"FF",X"FE",X"FF",X"FF",X"BF",X"FF",X"BF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FA",X"AF",X"EF",X"FF",X"BF",X"FF",X"BF",X"FF",
		X"FF",X"FA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"BF",X"FF",X"BF",X"FF",X"BF",X"FF",X"BF",X"FF",X"BF",X"FF",X"BF",X"FF",X"BF",X"FF",X"BF",X"FF",
		X"FF",X"FA",X"FE",X"A0",X"F8",X"0F",X"E3",X"FF",X"8F",X"FF",X"BF",X"FF",X"BF",X"FF",X"BF",X"FF",
		X"FF",X"FA",X"FE",X"A0",X"F8",X"00",X"E0",X"00",X"80",X"00",X"80",X"03",X"BF",X"FF",X"BF",X"FF",
		X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00",X"C0",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
