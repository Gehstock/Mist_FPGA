library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity spy_hunter_sound_cpu is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of spy_hunter_sound_cpu is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"F3",X"00",X"00",X"00",X"31",X"FF",X"83",X"ED",X"56",X"18",X"55",X"06",X"06",X"11",X"09",X"00",
		X"DD",X"21",X"BC",X"82",X"DD",X"7E",X"01",X"FE",X"FF",X"28",X"13",X"DD",X"4E",X"02",X"21",X"27",
		X"00",X"E5",X"DD",X"6E",X"00",X"67",X"E9",X"11",X"09",X"00",X"DD",X"36",X"02",X"00",X"DD",X"19",
		X"10",X"E2",X"C9",X"85",X"6F",X"D0",X"24",X"C9",X"F5",X"3A",X"00",X"E0",X"3A",X"75",X"83",X"3D",
		X"28",X"06",X"32",X"75",X"83",X"F1",X"FB",X"C9",X"3C",X"32",X"74",X"83",X"3E",X"06",X"32",X"75",
		X"83",X"F1",X"FB",X"C9",X"C5",X"42",X"21",X"00",X"00",X"54",X"78",X"B7",X"C3",X"E7",X"00",X"FF",
		X"21",X"00",X"B0",X"36",X"0F",X"21",X"02",X"B0",X"36",X"F0",X"3A",X"00",X"F0",X"CB",X"47",X"20",
		X"4F",X"CB",X"4F",X"20",X"2E",X"AF",X"32",X"77",X"83",X"CD",X"29",X"05",X"CD",X"E1",X"05",X"3A",
		X"77",X"83",X"FE",X"00",X"28",X"1D",X"CB",X"67",X"20",X"05",X"01",X"00",X"10",X"18",X"03",X"01",
		X"00",X"80",X"11",X"01",X"00",X"60",X"69",X"32",X"00",X"D0",X"37",X"3F",X"ED",X"52",X"20",X"FC",
		X"2F",X"18",X"F2",X"3E",X"FF",X"32",X"00",X"D0",X"3A",X"00",X"F0",X"CB",X"57",X"20",X"08",X"CD",
		X"55",X"06",X"18",X"EF",X"3A",X"00",X"F0",X"CB",X"5F",X"20",X"F9",X"CD",X"7C",X"06",X"18",X"F4",
		X"06",X"00",X"CD",X"38",X"06",X"06",X"FF",X"CD",X"38",X"06",X"06",X"55",X"CD",X"38",X"06",X"06",
		X"AA",X"CD",X"38",X"06",X"AF",X"32",X"77",X"83",X"CD",X"29",X"05",X"CD",X"E1",X"05",X"3A",X"77",
		X"83",X"32",X"00",X"C0",X"CD",X"EE",X"00",X"28",X"03",X"19",X"10",X"FD",X"C1",X"C9",X"31",X"FF",
		X"83",X"F3",X"ED",X"56",X"CD",X"13",X"01",X"CD",X"AD",X"07",X"FB",X"AF",X"32",X"74",X"83",X"CD",
		X"82",X"01",X"CD",X"0B",X"00",X"CD",X"AD",X"07",X"00",X"00",X"00",X"3A",X"74",X"83",X"B7",X"28",
		X"FA",X"18",X"E8",X"21",X"3C",X"1E",X"06",X"20",X"11",X"20",X"80",X"DD",X"21",X"00",X"80",X"7E",
		X"DD",X"77",X"00",X"2F",X"12",X"13",X"23",X"DD",X"23",X"10",X"F4",X"06",X"06",X"11",X"09",X"00",
		X"DD",X"21",X"BC",X"82",X"DD",X"36",X"00",X"FF",X"DD",X"36",X"01",X"FF",X"DD",X"36",X"02",X"00",
		X"DD",X"36",X"03",X"00",X"DD",X"36",X"04",X"00",X"DD",X"36",X"05",X"00",X"DD",X"36",X"06",X"00",
		X"DD",X"19",X"10",X"E0",X"06",X"03",X"21",X"6B",X"83",X"36",X"00",X"23",X"10",X"FB",X"3E",X"01",
		X"32",X"0C",X"83",X"32",X"20",X"83",X"3D",X"32",X"1F",X"83",X"3A",X"00",X"90",X"E6",X"80",X"32",
		X"6E",X"83",X"3E",X"55",X"32",X"71",X"83",X"3E",X"06",X"32",X"75",X"83",X"3E",X"52",X"32",X"76",
		X"83",X"C9",X"3A",X"6E",X"83",X"47",X"3A",X"00",X"90",X"A8",X"CB",X"7F",X"20",X"31",X"CB",X"40",
		X"28",X"1E",X"CB",X"80",X"78",X"32",X"6E",X"83",X"CD",X"E0",X"01",X"3A",X"70",X"83",X"CB",X"47",
		X"28",X"0E",X"CD",X"95",X"02",X"CD",X"A3",X"03",X"CD",X"06",X"04",X"CD",X"02",X"19",X"18",X"23",
		X"CD",X"A3",X"03",X"3A",X"6F",X"83",X"CB",X"47",X"28",X"19",X"CD",X"02",X"19",X"18",X"14",X"78",
		X"2F",X"CB",X"C7",X"32",X"6E",X"83",X"CD",X"A3",X"03",X"3A",X"6F",X"83",X"CB",X"47",X"28",X"03",
		X"CD",X"02",X"19",X"3E",X"01",X"32",X"20",X"83",X"32",X"0C",X"83",X"3D",X"32",X"1F",X"83",X"C9",
		X"3E",X"01",X"32",X"70",X"83",X"DD",X"21",X"00",X"90",X"DD",X"46",X"00",X"CB",X"70",X"28",X"23",
		X"FD",X"21",X"00",X"80",X"FD",X"7E",X"0F",X"E6",X"8F",X"4F",X"78",X"17",X"E6",X"70",X"B1",X"FD",
		X"77",X"0F",X"FD",X"7E",X"1F",X"E6",X"8F",X"4F",X"78",X"17",X"17",X"17",X"17",X"E6",X"70",X"B1",
		X"FD",X"77",X"1F",X"DD",X"7E",X"01",X"4F",X"FE",X"00",X"28",X"23",X"CB",X"7F",X"28",X"6E",X"DD",
		X"7E",X"02",X"CB",X"7F",X"20",X"67",X"79",X"E6",X"7F",X"4F",X"06",X"06",X"FD",X"21",X"BC",X"82",
		X"11",X"09",X"00",X"FD",X"7E",X"06",X"B9",X"CC",X"61",X"02",X"FD",X"19",X"10",X"F5",X"FD",X"21",
		X"6B",X"83",X"DD",X"46",X"02",X"78",X"E6",X"7F",X"28",X"24",X"CB",X"77",X"20",X"20",X"FD",X"77",
		X"01",X"DD",X"7E",X"01",X"CB",X"7F",X"C0",X"DD",X"7E",X"03",X"FE",X"00",X"C8",X"FD",X"77",X"02",
		X"C9",X"DD",X"7E",X"03",X"E5",X"FD",X"6E",X"07",X"FD",X"66",X"08",X"77",X"E1",X"C9",X"DD",X"4E",
		X"01",X"79",X"FE",X"00",X"20",X"09",X"DD",X"7E",X"03",X"FE",X"00",X"20",X"D4",X"18",X"09",X"CB",
		X"79",X"28",X"CE",X"CB",X"78",X"20",X"CA",X"AF",X"32",X"70",X"83",X"18",X"C4",X"79",X"E6",X"7F",
		X"32",X"6B",X"83",X"18",X"A9",X"06",X"03",X"21",X"6B",X"83",X"C5",X"7E",X"4F",X"FE",X"00",X"CA",
		X"66",X"03",X"3A",X"76",X"83",X"91",X"DA",X"66",X"03",X"79",X"FE",X"06",X"20",X"04",X"F3",X"C3",
		X"00",X"00",X"79",X"FE",X"01",X"20",X"0C",X"DD",X"21",X"00",X"80",X"DD",X"7E",X"1F",X"F6",X"80",
		X"DD",X"77",X"1F",X"79",X"FE",X"02",X"20",X"0F",X"DD",X"21",X"00",X"80",X"DD",X"7E",X"1F",X"E6",
		X"7F",X"DD",X"77",X"1F",X"CD",X"6D",X"03",X"79",X"FE",X"03",X"20",X"03",X"CD",X"6D",X"03",X"79",
		X"FE",X"04",X"20",X"07",X"3E",X"52",X"32",X"76",X"83",X"18",X"0A",X"79",X"FE",X"05",X"20",X"05",
		X"3E",X"52",X"32",X"76",X"83",X"79",X"D9",X"6F",X"26",X"00",X"54",X"5D",X"29",X"29",X"19",X"19",
		X"19",X"11",X"01",X"08",X"19",X"EB",X"1A",X"FE",X"00",X"20",X"1F",X"01",X"0C",X"83",X"60",X"69",
		X"3E",X"06",X"08",X"13",X"1A",X"FE",X"00",X"28",X"4A",X"7E",X"CD",X"33",X"00",X"1A",X"77",X"60",
		X"69",X"34",X"08",X"3D",X"FE",X"00",X"20",X"EA",X"18",X"39",X"3E",X"06",X"21",X"20",X"83",X"08",
		X"13",X"1A",X"FE",X"00",X"28",X"2D",X"7E",X"CD",X"33",X"00",X"1A",X"77",X"26",X"00",X"6F",X"29",
		X"01",X"46",X"0A",X"09",X"01",X"20",X"83",X"0A",X"CB",X"27",X"E5",X"21",X"33",X"83",X"CD",X"33",
		X"00",X"EB",X"E3",X"7E",X"12",X"23",X"13",X"7E",X"12",X"0A",X"3C",X"02",X"D1",X"60",X"69",X"08",
		X"3D",X"20",X"CC",X"D9",X"AF",X"77",X"23",X"C1",X"05",X"C2",X"9A",X"02",X"C9",X"D9",X"DD",X"21",
		X"BC",X"82",X"01",X"09",X"00",X"11",X"0C",X"83",X"3E",X"01",X"12",X"62",X"6B",X"3E",X"06",X"08",
		X"DD",X"7E",X"03",X"FE",X"00",X"28",X"0B",X"1A",X"CD",X"33",X"00",X"DD",X"7E",X"03",X"77",X"62",
		X"6B",X"34",X"DD",X"09",X"08",X"3D",X"20",X"E7",X"3E",X"00",X"32",X"1F",X"83",X"3C",X"32",X"20",
		X"83",X"D9",X"C9",X"AF",X"32",X"6F",X"83",X"21",X"0C",X"83",X"7E",X"D6",X"01",X"28",X"2A",X"11",
		X"09",X"00",X"4F",X"DD",X"21",X"BC",X"82",X"06",X"06",X"23",X"7E",X"DD",X"BE",X"04",X"20",X"13",
		X"AF",X"DD",X"77",X"06",X"DD",X"77",X"04",X"DD",X"77",X"05",X"3C",X"32",X"6F",X"83",X"0D",X"20",
		X"E2",X"18",X"06",X"DD",X"19",X"10",X"E4",X"18",X"F5",X"21",X"1F",X"83",X"7E",X"4F",X"FE",X"00",
		X"C8",X"3E",X"01",X"32",X"6F",X"83",X"06",X"06",X"21",X"5C",X"1E",X"DD",X"21",X"BC",X"82",X"11",
		X"09",X"00",X"79",X"A6",X"28",X"0A",X"AF",X"DD",X"77",X"06",X"DD",X"77",X"04",X"DD",X"77",X"05",
		X"DD",X"19",X"23",X"10",X"ED",X"C9",X"3A",X"20",X"83",X"D6",X"01",X"C8",X"08",X"CD",X"38",X"04",
		X"CD",X"54",X"04",X"79",X"CB",X"27",X"21",X"33",X"83",X"CD",X"33",X"00",X"7A",X"FE",X"00",X"20",
		X"11",X"CB",X"7E",X"20",X"0A",X"E5",X"CD",X"95",X"04",X"E1",X"7A",X"FE",X"00",X"20",X"03",X"CD",
		X"CE",X"04",X"23",X"36",X"00",X"08",X"18",X"D1",X"06",X"00",X"0E",X"01",X"16",X"01",X"3A",X"20",
		X"83",X"5F",X"21",X"33",X"83",X"23",X"7A",X"BB",X"C8",X"23",X"23",X"78",X"BE",X"30",X"02",X"46",
		X"4A",X"14",X"18",X"F2",X"79",X"CB",X"27",X"21",X"33",X"83",X"CD",X"33",X"00",X"C5",X"06",X"06",
		X"4E",X"11",X"09",X"00",X"21",X"5C",X"1E",X"DD",X"21",X"BC",X"82",X"7E",X"A1",X"28",X"1D",X"DD",
		X"7E",X"04",X"FE",X"00",X"20",X"16",X"21",X"20",X"83",X"C1",X"79",X"CD",X"33",X"00",X"7E",X"DD",
		X"77",X"04",X"DD",X"70",X"05",X"AF",X"DD",X"77",X"03",X"16",X"01",X"C9",X"DD",X"19",X"23",X"10",
		X"DA",X"16",X"00",X"C1",X"C9",X"26",X"06",X"11",X"09",X"00",X"DD",X"21",X"BC",X"82",X"DD",X"7E",
		X"04",X"FE",X"00",X"20",X"15",X"79",X"21",X"20",X"83",X"CD",X"33",X"00",X"7E",X"DD",X"77",X"04",
		X"DD",X"70",X"05",X"AF",X"DD",X"77",X"03",X"16",X"01",X"C9",X"DD",X"19",X"25",X"20",X"DF",X"16",
		X"00",X"21",X"33",X"83",X"79",X"CB",X"27",X"CD",X"33",X"00",X"F6",X"3F",X"77",X"C9",X"16",X"FF",
		X"1E",X"00",X"E5",X"C5",X"4E",X"06",X"00",X"DD",X"21",X"BC",X"82",X"21",X"5C",X"1E",X"7E",X"A1",
		X"28",X"08",X"DD",X"7E",X"05",X"BA",X"30",X"02",X"57",X"58",X"D5",X"11",X"09",X"00",X"DD",X"19",
		X"D1",X"23",X"04",X"78",X"FE",X"06",X"20",X"E6",X"C1",X"7A",X"B8",X"30",X"24",X"21",X"20",X"83",
		X"79",X"CD",X"33",X"00",X"4E",X"6B",X"26",X"00",X"54",X"5D",X"29",X"29",X"29",X"19",X"EB",X"DD",
		X"21",X"BC",X"82",X"DD",X"19",X"DD",X"71",X"04",X"DD",X"70",X"05",X"AF",X"DD",X"77",X"03",X"E1",
		X"C9",X"E1",X"C0",X"CB",X"76",X"C8",X"E5",X"18",X"D4",X"DD",X"21",X"D1",X"05",X"AF",X"F5",X"DD",
		X"6E",X"00",X"DD",X"66",X"01",X"7C",X"B5",X"20",X"0A",X"F1",X"47",X"3A",X"77",X"83",X"B0",X"32",
		X"77",X"83",X"C9",X"DD",X"5E",X"04",X"DD",X"56",X"05",X"DD",X"4E",X"02",X"DD",X"46",X"03",X"ED",
		X"B0",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"DD",X"5E",X"02",X"DD",X"56",X"03",X"7A",X"B3",X"28",
		X"11",X"06",X"02",X"3E",X"00",X"77",X"BE",X"C2",X"CC",X"05",X"F6",X"FF",X"10",X"F7",X"23",X"1B",
		X"18",X"EB",X"DD",X"66",X"01",X"DD",X"6E",X"00",X"DD",X"5E",X"02",X"DD",X"56",X"03",X"7A",X"B3",
		X"28",X"06",X"36",X"00",X"23",X"1B",X"18",X"F6",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"DD",X"5E",
		X"02",X"DD",X"56",X"03",X"7A",X"B3",X"28",X"14",X"7E",X"FE",X"00",X"20",X"2F",X"3E",X"01",X"77",
		X"BE",X"C2",X"CC",X"05",X"CB",X"27",X"30",X"F7",X"23",X"1B",X"18",X"E8",X"AF",X"DD",X"66",X"05",
		X"DD",X"6E",X"04",X"DD",X"56",X"01",X"DD",X"5E",X"00",X"DD",X"4E",X"02",X"DD",X"46",X"03",X"ED",
		X"B0",X"47",X"F1",X"B0",X"11",X"07",X"00",X"DD",X"19",X"C3",X"2E",X"05",X"DD",X"7E",X"06",X"18",
		X"DC",X"00",X"80",X"00",X"02",X"00",X"80",X"10",X"00",X"82",X"00",X"02",X"00",X"80",X"10",X"00",
		X"00",X"DD",X"21",X"1D",X"06",X"16",X"00",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"DD",X"4E",X"00",
		X"DD",X"46",X"01",X"78",X"B1",X"28",X"1A",X"AF",X"86",X"23",X"0D",X"20",X"FB",X"05",X"20",X"F8",
		X"DD",X"BE",X"04",X"28",X"05",X"7A",X"DD",X"B6",X"05",X"57",X"01",X"06",X"00",X"DD",X"09",X"18",
		X"D6",X"7A",X"B7",X"C8",X"47",X"3A",X"77",X"83",X"B0",X"32",X"77",X"83",X"C9",X"00",X"10",X"00",
		X"00",X"D7",X"01",X"00",X"10",X"00",X"10",X"BD",X"02",X"00",X"00",X"00",X"20",X"00",X"04",X"00",
		X"00",X"00",X"30",X"00",X"08",X"00",X"00",X"29",X"3A",X"00",X"90",X"B8",X"20",X"FA",X"3A",X"01",
		X"90",X"B8",X"20",X"F4",X"3A",X"02",X"90",X"B8",X"20",X"EE",X"3A",X"03",X"90",X"B8",X"20",X"E8",
		X"78",X"32",X"00",X"C0",X"C9",X"06",X"00",X"CD",X"B5",X"06",X"0E",X"00",X"3E",X"AD",X"CD",X"F5",
		X"06",X"0E",X"01",X"3E",X"07",X"CD",X"F5",X"06",X"06",X"01",X"CD",X"B5",X"06",X"0E",X"00",X"3E",
		X"AD",X"CD",X"F5",X"06",X"0E",X"01",X"3E",X"77",X"CD",X"F5",X"06",X"C9",X"CD",X"55",X"06",X"16",
		X"10",X"3E",X"00",X"1E",X"FF",X"06",X"00",X"0E",X"00",X"CD",X"F5",X"06",X"2F",X"0E",X"01",X"CD",
		X"F5",X"06",X"06",X"01",X"32",X"78",X"83",X"E6",X"7F",X"CD",X"F5",X"06",X"3A",X"78",X"83",X"2F",
		X"0E",X"00",X"CD",X"F5",X"06",X"3C",X"E6",X"0F",X"47",X"07",X"07",X"07",X"07",X"B0",X"1D",X"20",
		X"FD",X"15",X"20",X"CF",X"C9",X"CD",X"0C",X"07",X"36",X"00",X"DD",X"36",X"00",X"F4",X"36",X"01",
		X"DD",X"36",X"00",X"01",X"36",X"02",X"DD",X"36",X"00",X"FA",X"36",X"03",X"DD",X"36",X"00",X"00",
		X"36",X"04",X"DD",X"36",X"00",X"7D",X"36",X"05",X"DD",X"36",X"00",X"00",X"36",X"08",X"DD",X"36",
		X"00",X"0B",X"36",X"09",X"DD",X"36",X"00",X"0B",X"36",X"0A",X"DD",X"36",X"00",X"0B",X"36",X"07",
		X"DD",X"36",X"00",X"F8",X"C9",X"CD",X"0C",X"07",X"32",X"72",X"83",X"AF",X"A9",X"28",X"09",X"36",
		X"0F",X"3A",X"72",X"83",X"DD",X"77",X"00",X"C9",X"36",X"0E",X"18",X"F5",X"32",X"72",X"83",X"AF",
		X"A8",X"3A",X"72",X"83",X"20",X"08",X"21",X"00",X"A0",X"DD",X"21",X"02",X"A0",X"C9",X"21",X"00",
		X"B0",X"DD",X"21",X"02",X"B0",X"C9",X"21",X"F4",X"07",X"16",X"00",X"19",X"56",X"21",X"E8",X"07",
		X"79",X"CB",X"27",X"5F",X"7A",X"16",X"00",X"19",X"5E",X"23",X"56",X"6F",X"26",X"00",X"19",X"11",
		X"40",X"80",X"19",X"C9",X"21",X"62",X"1E",X"CB",X"27",X"D2",X"53",X"07",X"24",X"CD",X"33",X"00",
		X"C3",X"56",X"07",X"CD",X"33",X"00",X"E5",X"1E",X"38",X"51",X"CD",X"54",X"00",X"11",X"EC",X"1C",
		X"19",X"C5",X"4E",X"23",X"46",X"60",X"69",X"C1",X"D1",X"1A",X"77",X"23",X"13",X"1A",X"77",X"C9",
		X"C5",X"3E",X"06",X"90",X"47",X"57",X"1E",X"38",X"CD",X"54",X"00",X"EB",X"FD",X"21",X"EC",X"1C",
		X"FD",X"19",X"16",X"00",X"58",X"21",X"3E",X"82",X"19",X"FD",X"7E",X"14",X"4F",X"FE",X"0F",X"7E",
		X"20",X"17",X"CB",X"27",X"CB",X"27",X"CB",X"27",X"CB",X"27",X"E6",X"F0",X"47",X"FD",X"6E",X"12",
		X"FD",X"66",X"13",X"7E",X"A1",X"B0",X"77",X"C1",X"C9",X"E6",X"0F",X"18",X"EF",X"01",X"1F",X"00",
		X"21",X"00",X"80",X"11",X"20",X"80",X"09",X"EB",X"09",X"06",X"0F",X"DD",X"21",X"00",X"B0",X"1A",
		X"BE",X"28",X"07",X"77",X"DD",X"70",X"00",X"32",X"02",X"B0",X"1B",X"2B",X"05",X"F2",X"BF",X"07",
		X"06",X"0F",X"DD",X"21",X"00",X"A0",X"1A",X"BE",X"28",X"07",X"77",X"DD",X"70",X"00",X"32",X"02",
		X"A0",X"1B",X"2B",X"05",X"F2",X"D6",X"07",X"C9",X"00",X"00",X"55",X"00",X"AA",X"00",X"FF",X"00",
		X"54",X"01",X"A9",X"01",X"00",X"11",X"22",X"33",X"44",X"4D",X"49",X"44",X"57",X"41",X"59",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"01",X"02",X"03",X"04",X"05",X"06",X"00",X"01",X"02",X"03",X"04",X"05",X"06",
		X"01",X"07",X"07",X"07",X"07",X"07",X"07",X"00",X"07",X"07",X"07",X"07",X"07",X"07",X"01",X"08",
		X"00",X"00",X"00",X"00",X"00",X"01",X"09",X"0A",X"0B",X"0C",X"00",X"00",X"01",X"47",X"00",X"00",
		X"00",X"00",X"00",X"00",X"47",X"00",X"00",X"00",X"00",X"00",X"01",X"40",X"00",X"00",X"00",X"00",
		X"00",X"00",X"26",X"00",X"00",X"00",X"00",X"00",X"01",X"10",X"00",X"00",X"00",X"00",X"00",X"01",
		X"11",X"00",X"00",X"00",X"00",X"00",X"01",X"12",X"13",X"14",X"15",X"16",X"17",X"00",X"12",X"13",
		X"14",X"15",X"16",X"17",X"01",X"18",X"19",X"1A",X"1B",X"1C",X"00",X"00",X"18",X"19",X"1A",X"1B",
		X"1C",X"00",X"01",X"1D",X"1E",X"1F",X"20",X"00",X"00",X"00",X"1D",X"1E",X"1F",X"20",X"00",X"00",
		X"01",X"21",X"22",X"23",X"00",X"00",X"00",X"00",X"21",X"22",X"23",X"00",X"00",X"00",X"01",X"24",
		X"25",X"00",X"00",X"00",X"00",X"00",X"24",X"25",X"00",X"00",X"00",X"00",X"01",X"26",X"00",X"00",
		X"00",X"00",X"00",X"00",X"2B",X"00",X"00",X"00",X"00",X"00",X"01",X"27",X"00",X"00",X"00",X"00",
		X"00",X"00",X"27",X"00",X"00",X"00",X"00",X"00",X"00",X"2A",X"00",X"00",X"00",X"00",X"00",X"01",
		X"29",X"00",X"00",X"00",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"00",X"00",X"01",X"2A",X"00",
		X"00",X"00",X"00",X"00",X"01",X"2B",X"00",X"00",X"00",X"00",X"00",X"01",X"2C",X"00",X"00",X"00",
		X"00",X"00",X"01",X"2D",X"00",X"00",X"00",X"00",X"00",X"00",X"2D",X"00",X"00",X"00",X"00",X"00",
		X"01",X"2E",X"2F",X"00",X"00",X"00",X"00",X"00",X"2E",X"2F",X"35",X"36",X"41",X"42",X"01",X"35",
		X"36",X"00",X"00",X"00",X"00",X"01",X"41",X"42",X"00",X"00",X"00",X"00",X"01",X"30",X"00",X"00",
		X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"01",X"31",X"00",X"00",X"00",X"00",
		X"00",X"01",X"32",X"00",X"00",X"00",X"00",X"00",X"01",X"33",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"00",X"00",X"00",X"00",X"00",X"01",X"34",X"00",X"00",X"00",X"00",X"00",X"00",X"34",X"00",
		X"00",X"00",X"00",X"00",X"01",X"37",X"28",X"3F",X"00",X"00",X"00",X"00",X"37",X"28",X"3F",X"00",
		X"00",X"00",X"01",X"38",X"00",X"00",X"00",X"00",X"00",X"01",X"39",X"00",X"00",X"00",X"00",X"00",
		X"00",X"39",X"00",X"00",X"00",X"00",X"00",X"01",X"3A",X"00",X"00",X"00",X"00",X"00",X"00",X"3A",
		X"00",X"00",X"00",X"00",X"00",X"01",X"3B",X"00",X"00",X"00",X"00",X"00",X"00",X"3B",X"00",X"00",
		X"00",X"00",X"00",X"01",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"00",X"00",X"00",X"00",
		X"00",X"01",X"3D",X"00",X"00",X"00",X"00",X"00",X"00",X"3D",X"00",X"00",X"00",X"00",X"00",X"01",
		X"3E",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"3D",X"3C",X"3B",X"00",X"00",X"01",X"0F",X"00",
		X"00",X"00",X"00",X"00",X"01",X"0D",X"00",X"00",X"00",X"00",X"00",X"01",X"43",X"00",X"00",X"00",
		X"00",X"00",X"01",X"44",X"00",X"00",X"00",X"00",X"00",X"01",X"45",X"00",X"00",X"00",X"00",X"00",
		X"01",X"46",X"00",X"00",X"00",X"00",X"00",X"00",X"43",X"44",X"45",X"46",X"00",X"00",X"01",X"48",
		X"49",X"4A",X"48",X"49",X"4A",X"00",X"31",X"00",X"00",X"00",X"00",X"00",X"01",X"4B",X"00",X"00",
		X"00",X"00",X"00",X"00",X"4B",X"00",X"00",X"00",X"00",X"00",X"01",X"4C",X"4D",X"00",X"00",X"00",
		X"00",X"00",X"4C",X"4D",X"00",X"00",X"00",X"00",X"01",X"4E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"4E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"02",X"02",X"04",X"03",X"08",X"04",
		X"10",X"05",X"20",X"06",X"FF",X"90",X"82",X"81",X"C2",X"77",X"C4",X"77",X"C8",X"77",X"D0",X"77",
		X"82",X"0D",X"C2",X"1E",X"82",X"0F",X"82",X"29",X"82",X"32",X"81",X"80",X"82",X"80",X"84",X"64",
		X"88",X"80",X"90",X"7F",X"A0",X"80",X"81",X"7C",X"82",X"62",X"84",X"80",X"88",X"71",X"90",X"82",
		X"81",X"7C",X"82",X"51",X"88",X"50",X"90",X"71",X"81",X"80",X"88",X"80",X"90",X"81",X"82",X"2C",
		X"88",X"4D",X"C8",X"2C",X"E0",X"50",X"81",X"7E",X"C1",X"7D",X"88",X"70",X"88",X"70",X"C2",X"31",
		X"84",X"66",X"90",X"80",X"84",X"65",X"81",X"7F",X"88",X"57",X"81",X"7E",X"84",X"67",X"C8",X"2C",
		X"90",X"81",X"84",X"66",X"A0",X"60",X"C2",X"3F",X"E0",X"50",X"E0",X"50",X"E0",X"50",X"E0",X"50",
		X"E0",X"50",X"E0",X"50",X"82",X"70",X"C8",X"2C",X"90",X"82",X"84",X"67",X"E0",X"50",X"E0",X"50",
		X"E0",X"50",X"E0",X"50",X"82",X"50",X"89",X"51",X"92",X"51",X"A4",X"51",X"88",X"56",X"E0",X"50",
		X"C1",X"50",X"81",X"7C",X"BE",X"0C",X"FF",X"FF",X"FF",X"FF",X"CC",X"0C",X"DA",X"0C",X"6D",X"18",
		X"EC",X"0C",X"FA",X"0C",X"6D",X"18",X"0F",X"0D",X"1D",X"0D",X"6D",X"18",X"32",X"0D",X"40",X"0D",
		X"6D",X"18",X"55",X"0D",X"63",X"0D",X"6D",X"18",X"78",X"0D",X"86",X"0D",X"6D",X"18",X"9E",X"0D",
		X"AC",X"0D",X"7B",X"18",X"BE",X"0D",X"CC",X"0D",X"6D",X"18",X"E1",X"0D",X"ED",X"0D",X"04",X"16",
		X"1E",X"0E",X"2A",X"0E",X"04",X"16",X"3C",X"0E",X"48",X"0E",X"04",X"16",X"5D",X"0E",X"69",X"0E",
		X"04",X"16",X"BA",X"0E",X"C8",X"0E",X"74",X"18",X"DD",X"0E",X"EB",X"0E",X"88",X"18",X"15",X"0F",
		X"21",X"0F",X"6D",X"18",X"2D",X"0F",X"39",X"0F",X"6D",X"18",X"4B",X"0F",X"59",X"0F",X"95",X"18",
		X"7D",X"0F",X"D1",X"0F",X"88",X"18",X"8B",X"0F",X"D1",X"0F",X"88",X"18",X"99",X"0F",X"D1",X"0F",
		X"88",X"18",X"A7",X"0F",X"D1",X"0F",X"88",X"18",X"B5",X"0F",X"D1",X"0F",X"88",X"18",X"C3",X"0F",
		X"D1",X"0F",X"88",X"18",X"FA",X"0F",X"40",X"10",X"88",X"18",X"08",X"10",X"40",X"10",X"88",X"18",
		X"16",X"10",X"40",X"10",X"88",X"18",X"24",X"10",X"40",X"10",X"88",X"18",X"32",X"10",X"40",X"10",
		X"88",X"18",X"5D",X"10",X"8D",X"10",X"88",X"18",X"69",X"10",X"8D",X"10",X"88",X"18",X"75",X"10",
		X"8D",X"10",X"88",X"18",X"81",X"10",X"8D",X"10",X"88",X"18",X"AA",X"10",X"CE",X"10",X"88",X"18",
		X"B6",X"10",X"CE",X"10",X"88",X"18",X"C2",X"10",X"CE",X"10",X"88",X"18",X"EB",X"10",X"03",X"11",
		X"88",X"18",X"F7",X"10",X"03",X"11",X"88",X"18",X"20",X"11",X"2C",X"11",X"A2",X"18",X"F6",X"15",
		X"1C",X"17",X"17",X"16",X"41",X"14",X"88",X"14",X"AF",X"18",X"BA",X"11",X"C8",X"11",X"6D",X"18",
		X"D7",X"11",X"E5",X"11",X"74",X"18",X"F4",X"11",X"02",X"12",X"74",X"18",X"11",X"12",X"1D",X"12",
		X"88",X"18",X"37",X"12",X"45",X"12",X"88",X"18",X"61",X"12",X"9B",X"12",X"DC",X"18",X"AA",X"12",
		X"BA",X"12",X"DC",X"18",X"E7",X"12",X"F5",X"12",X"88",X"18",X"12",X"13",X"20",X"13",X"C9",X"18",
		X"4D",X"13",X"70",X"13",X"95",X"18",X"7F",X"13",X"8B",X"13",X"88",X"18",X"96",X"13",X"B1",X"13",
		X"A4",X"13",X"61",X"12",X"D5",X"13",X"DC",X"18",X"AA",X"12",X"F3",X"13",X"DC",X"18",X"23",X"14",
		X"4F",X"14",X"AF",X"18",X"18",X"15",X"24",X"15",X"88",X"18",X"4D",X"15",X"A8",X"15",X"EF",X"18",
		X"5B",X"15",X"A8",X"15",X"EF",X"18",X"C6",X"15",X"46",X"16",X"17",X"16",X"D2",X"15",X"24",X"16",
		X"17",X"16",X"DE",X"15",X"46",X"16",X"17",X"16",X"EA",X"15",X"35",X"16",X"17",X"16",X"31",X"14",
		X"4F",X"14",X"AF",X"18",X"69",X"15",X"77",X"15",X"BC",X"18",X"61",X"12",X"6D",X"17",X"DC",X"18",
		X"AA",X"12",X"7C",X"17",X"DC",X"18",X"57",X"16",X"75",X"16",X"EF",X"18",X"61",X"16",X"86",X"16",
		X"EF",X"18",X"61",X"16",X"97",X"16",X"EF",X"18",X"6B",X"16",X"A8",X"16",X"EF",X"18",X"7E",X"0E",
		X"8E",X"0E",X"DC",X"18",X"41",X"14",X"D0",X"14",X"AF",X"18",X"23",X"14",X"D0",X"14",X"AF",X"18",
		X"31",X"14",X"D0",X"14",X"AF",X"18",X"8B",X"17",X"A5",X"17",X"95",X"18",X"B4",X"17",X"D8",X"17",
		X"DC",X"18",X"C6",X"17",X"D8",X"17",X"DC",X"18",X"25",X"18",X"33",X"18",X"C9",X"18",X"CD",X"65",
		X"19",X"00",X"00",X"FF",X"0A",X"00",X"FF",X"C9",X"CD",X"70",X"07",X"C9",X"CD",X"65",X"19",X"01",
		X"02",X"FF",X"0A",X"01",X"00",X"DE",X"02",X"01",X"FF",X"C9",X"CD",X"6A",X"1A",X"C7",X"0C",X"00",
		X"01",X"00",X"04",X"01",X"03",X"01",X"34",X"00",X"04",X"01",X"FD",X"00",X"CD",X"65",X"19",X"01",
		X"02",X"FF",X"0A",X"01",X"00",X"AA",X"02",X"01",X"FF",X"C9",X"CD",X"6A",X"1A",X"C7",X"0C",X"00",
		X"01",X"00",X"01",X"3C",X"00",X"04",X"01",X"03",X"01",X"34",X"00",X"04",X"01",X"FD",X"00",X"CD",
		X"65",X"19",X"01",X"02",X"FF",X"0A",X"01",X"00",X"7B",X"02",X"01",X"FF",X"C9",X"CD",X"6A",X"1A",
		X"C7",X"0C",X"00",X"01",X"00",X"01",X"78",X"00",X"04",X"01",X"03",X"01",X"34",X"00",X"04",X"01",
		X"FD",X"00",X"CD",X"65",X"19",X"01",X"02",X"FF",X"0A",X"01",X"00",X"52",X"02",X"01",X"FF",X"C9",
		X"CD",X"6A",X"1A",X"C7",X"0C",X"00",X"01",X"00",X"01",X"B4",X"00",X"04",X"01",X"03",X"01",X"34",
		X"00",X"04",X"01",X"FD",X"00",X"CD",X"65",X"19",X"01",X"02",X"FF",X"0A",X"01",X"00",X"2D",X"02",
		X"01",X"FF",X"C9",X"CD",X"6A",X"1A",X"C7",X"0C",X"00",X"01",X"00",X"01",X"F0",X"00",X"04",X"01",
		X"03",X"01",X"34",X"00",X"04",X"01",X"FD",X"00",X"CD",X"65",X"19",X"01",X"02",X"FF",X"0A",X"01",
		X"00",X"0C",X"02",X"01",X"FF",X"C9",X"CD",X"6A",X"1A",X"C7",X"0C",X"00",X"01",X"00",X"01",X"C8",
		X"00",X"01",X"64",X"00",X"04",X"01",X"03",X"01",X"34",X"00",X"04",X"01",X"FD",X"00",X"CD",X"65",
		X"19",X"01",X"05",X"FF",X"0A",X"0E",X"00",X"50",X"02",X"00",X"FF",X"C9",X"CD",X"6A",X"1A",X"C7",
		X"0C",X"00",X"01",X"FF",X"02",X"01",X"07",X"01",X"07",X"00",X"07",X"01",X"FE",X"00",X"CD",X"65",
		X"19",X"01",X"01",X"FF",X"0A",X"03",X"00",X"A9",X"02",X"00",X"FF",X"C9",X"CD",X"6A",X"1A",X"C7",
		X"0C",X"00",X"01",X"04",X"04",X"01",X"03",X"02",X"02",X"FF",X"01",X"05",X"00",X"05",X"01",X"FE",
		X"00",X"CD",X"65",X"19",X"01",X"08",X"FF",X"0A",X"07",X"18",X"1E",X"FF",X"C9",X"CD",X"6A",X"1A",
		X"FF",X"0D",X"00",X"01",X"00",X"07",X"02",X"01",X"01",X"14",X"00",X"0E",X"03",X"FF",X"00",X"CD",
		X"7B",X"1B",X"0D",X"0E",X"01",X"FF",X"01",X"02",X"01",X"01",X"03",X"FF",X"00",X"CD",X"6A",X"1A",
		X"C7",X"0C",X"02",X"02",X"FF",X"05",X"01",X"F0",X"FF",X"05",X"02",X"10",X"00",X"00",X"CD",X"65",
		X"19",X"01",X"08",X"FF",X"0A",X"07",X"18",X"19",X"FF",X"C9",X"CD",X"6A",X"1A",X"FF",X"0D",X"00",
		X"01",X"00",X"07",X"02",X"01",X"01",X"12",X"00",X"0E",X"03",X"FF",X"00",X"CD",X"65",X"19",X"01",
		X"07",X"FF",X"0A",X"00",X"18",X"16",X"FF",X"C9",X"CD",X"6A",X"1A",X"FF",X"0D",X"00",X"01",X"00",
		X"01",X"0F",X"00",X"05",X"02",X"03",X"01",X"0A",X"00",X"0F",X"05",X"FF",X"00",X"CD",X"65",X"19",
		X"01",X"07",X"FF",X"0A",X"00",X"18",X"11",X"FF",X"C9",X"CD",X"6A",X"1A",X"FF",X"0D",X"00",X"01",
		X"00",X"01",X"0F",X"00",X"05",X"02",X"03",X"01",X"08",X"00",X"0F",X"05",X"FF",X"00",X"CD",X"65",
		X"19",X"01",X"01",X"FF",X"0A",X"00",X"00",X"81",X"02",X"00",X"2A",X"01",X"FF",X"C9",X"CD",X"6A",
		X"1A",X"9A",X"0E",X"01",X"01",X"00",X"07",X"C0",X"01",X"00",X"CD",X"6A",X"1A",X"A9",X"0E",X"00",
		X"01",X"00",X"05",X"01",X"02",X"08",X"50",X"FF",X"00",X"CD",X"6A",X"1A",X"C7",X"0C",X"02",X"02",
		X"00",X"90",X"04",X"02",X"00",X"FF",X"03",X"02",X"00",X"00",X"CD",X"65",X"19",X"10",X"07",X"FF",
		X"0A",X"0E",X"04",X"10",X"2A",X"0B",X"FF",X"C9",X"CD",X"6A",X"1A",X"C8",X"0C",X"00",X"01",X"00",
		X"04",X"06",X"FF",X"02",X"02",X"FF",X"03",X"14",X"01",X"07",X"0B",X"01",X"00",X"CD",X"65",X"19",
		X"01",X"04",X"FF",X"0A",X"0C",X"18",X"A8",X"04",X"1F",X"FF",X"C9",X"CD",X"7B",X"1B",X"06",X"0F",
		X"01",X"1C",X"01",X"01",X"EA",X"01",X"01",X"13",X"00",X"01",X"01",X"F7",X"01",X"01",X"08",X"01",
		X"01",X"F7",X"01",X"01",X"09",X"00",X"CD",X"6A",X"1A",X"C7",X"0C",X"00",X"01",X"FF",X"03",X"02",
		X"01",X"01",X"01",X"FD",X"00",X"CD",X"65",X"19",X"10",X"00",X"FF",X"0A",X"0F",X"04",X"0B",X"FF",
		X"C9",X"CD",X"6A",X"1A",X"C7",X"0C",X"00",X"01",X"00",X"0F",X"01",X"FF",X"00",X"CD",X"65",X"19",
		X"10",X"04",X"FF",X"0A",X"0D",X"04",X"04",X"FF",X"C9",X"CD",X"6A",X"1A",X"C7",X"0C",X"00",X"01",
		X"00",X"01",X"07",X"F3",X"01",X"0D",X"0D",X"01",X"08",X"F3",X"00",X"CD",X"65",X"19",X"10",X"0B",
		X"FF",X"2A",X"0B",X"0A",X"0F",X"04",X"1F",X"FF",X"C9",X"CD",X"6A",X"1A",X"6B",X"0F",X"00",X"01",
		X"00",X"04",X"04",X"FF",X"01",X"01",X"04",X"0F",X"06",X"FF",X"00",X"CD",X"6A",X"1A",X"C8",X"0C",
		X"01",X"01",X"00",X"03",X"05",X"00",X"01",X"02",X"FB",X"1E",X"03",X"00",X"00",X"CD",X"65",X"19",
		X"01",X"04",X"FF",X"0A",X"0F",X"18",X"00",X"2A",X"04",X"FF",X"C9",X"CD",X"65",X"19",X"01",X"04",
		X"FF",X"0A",X"0F",X"18",X"04",X"2A",X"04",X"FF",X"C9",X"CD",X"65",X"19",X"01",X"04",X"FF",X"0A",
		X"0F",X"18",X"08",X"2A",X"04",X"FF",X"C9",X"CD",X"65",X"19",X"01",X"04",X"FF",X"0A",X"0F",X"18",
		X"0C",X"2A",X"04",X"FF",X"C9",X"CD",X"65",X"19",X"01",X"04",X"FF",X"0A",X"0F",X"18",X"10",X"2A",
		X"04",X"FF",X"C9",X"CD",X"65",X"19",X"01",X"04",X"FF",X"0A",X"0F",X"18",X"14",X"2A",X"04",X"FF",
		X"C9",X"CD",X"7B",X"1B",X"DF",X"0F",X"01",X"FF",X"05",X"01",X"02",X"05",X"01",X"FE",X"00",X"CD",
		X"6A",X"1A",X"C7",X"0C",X"00",X"01",X"00",X"01",X"08",X"00",X"03",X"01",X"FB",X"01",X"03",X"00",
		X"03",X"01",X"05",X"01",X"20",X"00",X"0F",X"0A",X"FF",X"00",X"CD",X"65",X"19",X"01",X"04",X"FF",
		X"0A",X"0F",X"18",X"00",X"2A",X"04",X"FF",X"C9",X"CD",X"65",X"19",X"01",X"04",X"FF",X"0A",X"0F",
		X"18",X"04",X"2A",X"04",X"FF",X"C9",X"CD",X"65",X"19",X"01",X"04",X"FF",X"0A",X"0F",X"18",X"08",
		X"2A",X"04",X"FF",X"C9",X"CD",X"65",X"19",X"01",X"04",X"FF",X"0A",X"0F",X"18",X"0C",X"2A",X"04",
		X"FF",X"C9",X"CD",X"65",X"19",X"01",X"04",X"FF",X"0A",X"0F",X"18",X"10",X"2A",X"04",X"FF",X"C9",
		X"CD",X"7B",X"1B",X"4E",X"10",X"01",X"FF",X"06",X"01",X"02",X"06",X"01",X"FE",X"00",X"CD",X"6A",
		X"1A",X"C7",X"0C",X"00",X"01",X"00",X"01",X"10",X"00",X"0F",X"09",X"FF",X"00",X"CD",X"65",X"19",
		X"01",X"04",X"FF",X"18",X"00",X"0A",X"0F",X"FF",X"C9",X"CD",X"65",X"19",X"01",X"04",X"FF",X"18",
		X"02",X"0A",X"0F",X"FF",X"C9",X"CD",X"65",X"19",X"01",X"04",X"FF",X"18",X"04",X"0A",X"0F",X"FF",
		X"C9",X"CD",X"65",X"19",X"01",X"04",X"FF",X"18",X"06",X"0A",X"0F",X"FF",X"C9",X"CD",X"7B",X"1B",
		X"9B",X"10",X"01",X"FF",X"04",X"01",X"04",X"04",X"01",X"FC",X"00",X"CD",X"6A",X"1A",X"C7",X"0C",
		X"00",X"01",X"00",X"01",X"0C",X"00",X"0F",X"08",X"FF",X"00",X"CD",X"65",X"19",X"01",X"02",X"FF",
		X"0A",X"0F",X"18",X"10",X"FF",X"C9",X"CD",X"65",X"19",X"01",X"02",X"FF",X"0A",X"0F",X"18",X"15",
		X"FF",X"C9",X"CD",X"65",X"19",X"01",X"02",X"FF",X"0A",X"0F",X"18",X"18",X"FF",X"C9",X"CD",X"7B",
		X"1B",X"DC",X"10",X"01",X"FF",X"04",X"01",X"02",X"04",X"01",X"FE",X"00",X"CD",X"6A",X"1A",X"C7",
		X"0C",X"00",X"01",X"00",X"01",X"18",X"00",X"0F",X"0E",X"FF",X"00",X"CD",X"65",X"19",X"01",X"07",
		X"FF",X"0A",X"0F",X"18",X"00",X"FF",X"C9",X"CD",X"65",X"19",X"01",X"07",X"FF",X"0A",X"0F",X"18",
		X"02",X"FF",X"C9",X"CD",X"7B",X"1B",X"11",X"11",X"01",X"FF",X"07",X"01",X"02",X"07",X"01",X"FE",
		X"00",X"CD",X"6A",X"1A",X"C7",X"0C",X"00",X"01",X"00",X"01",X"0A",X"00",X"0F",X"07",X"FF",X"00",
		X"CD",X"65",X"19",X"10",X"06",X"FF",X"0A",X"0C",X"04",X"1E",X"FF",X"C9",X"CD",X"6A",X"1A",X"3E",
		X"11",X"00",X"01",X"01",X"03",X"03",X"01",X"01",X"04",X"F1",X"01",X"09",X"0C",X"00",X"CD",X"6A",
		X"1A",X"C7",X"0C",X"01",X"01",X"FF",X"01",X"09",X"F1",X"01",X"07",X"F1",X"01",X"05",X"0F",X"01",
		X"03",X"0F",X"00",X"CD",X"65",X"19",X"10",X"08",X"FF",X"0A",X"0E",X"04",X"18",X"2C",X"23",X"2A",
		X"08",X"FF",X"C9",X"CD",X"33",X"1A",X"00",X"0A",X"0A",X"CD",X"33",X"1A",X"01",X"2C",X"2C",X"CD",
		X"C9",X"1C",X"20",X"CD",X"33",X"1A",X"02",X"2A",X"2A",X"C9",X"CD",X"6A",X"1A",X"89",X"11",X"00",
		X"01",X"FF",X"07",X"01",X"FE",X"01",X"30",X"0E",X"00",X"CD",X"70",X"07",X"CD",X"6A",X"1A",X"9B",
		X"11",X"02",X"01",X"FF",X"04",X"21",X"FF",X"04",X"17",X"01",X"00",X"CD",X"6A",X"1A",X"B6",X"11",
		X"01",X"01",X"FF",X"06",X"20",X"01",X"07",X"18",X"FF",X"04",X"20",X"02",X"03",X"20",X"FE",X"07",
		X"18",X"01",X"08",X"20",X"FF",X"00",X"CD",X"A9",X"1C",X"C9",X"CD",X"65",X"19",X"10",X"03",X"FF",
		X"0A",X"0F",X"04",X"1E",X"2A",X"03",X"FF",X"C9",X"CD",X"6A",X"1A",X"C7",X"0C",X"00",X"01",X"FF",
		X"01",X"04",X"F1",X"01",X"08",X"0F",X"00",X"CD",X"65",X"19",X"10",X"0F",X"FF",X"0A",X"0F",X"04",
		X"00",X"2A",X"0F",X"FF",X"C9",X"CD",X"6A",X"1A",X"C8",X"0C",X"00",X"01",X"07",X"08",X"03",X"FF",
		X"07",X"02",X"01",X"00",X"CD",X"65",X"19",X"10",X"0F",X"FF",X"0A",X"0F",X"2A",X"0F",X"04",X"1F",
		X"FF",X"C9",X"CD",X"6A",X"1A",X"C8",X"0C",X"00",X"01",X"00",X"0F",X"0F",X"FF",X"0F",X"0F",X"01",
		X"00",X"CD",X"65",X"19",X"01",X"03",X"FF",X"0A",X"05",X"18",X"85",X"FF",X"C9",X"CD",X"7B",X"1B",
		X"2B",X"12",X"01",X"05",X"03",X"01",X"FD",X"02",X"01",X"02",X"00",X"CD",X"6A",X"1A",X"C7",X"0C",
		X"00",X"01",X"00",X"0A",X"03",X"01",X"00",X"CD",X"65",X"19",X"01",X"08",X"FF",X"0A",X"0C",X"18",
		X"00",X"04",X"08",X"FF",X"C9",X"CD",X"7B",X"1B",X"52",X"12",X"01",X"00",X"50",X"01",X"02",X"FF",
		X"FE",X"00",X"CD",X"6A",X"1A",X"C7",X"0C",X"00",X"01",X"FF",X"01",X"04",X"F4",X"03",X"01",X"04",
		X"00",X"CD",X"65",X"19",X"01",X"0F",X"FF",X"0A",X"0F",X"02",X"0F",X"2A",X"0F",X"00",X"FF",X"FF",
		X"C9",X"CD",X"6A",X"1A",X"C7",X"0C",X"00",X"01",X"FF",X"01",X"03",X"F1",X"01",X"06",X"0F",X"00",
		X"CD",X"70",X"07",X"CD",X"6A",X"1A",X"71",X"12",X"01",X"01",X"00",X"03",X"60",X"FF",X"02",X"50",
		X"FF",X"02",X"40",X"FF",X"01",X"40",X"FF",X"FF",X"FF",X"00",X"00",X"CD",X"6A",X"1A",X"80",X"12",
		X"02",X"01",X"FF",X"04",X"08",X"F0",X"04",X"08",X"10",X"00",X"CD",X"65",X"19",X"01",X"0F",X"FF",
		X"0A",X"0F",X"02",X"00",X"00",X"10",X"2A",X"0F",X"FF",X"C9",X"CD",X"6A",X"1A",X"80",X"12",X"02",
		X"01",X"FF",X"03",X"01",X"FF",X"01",X"06",X"03",X"00",X"CD",X"6A",X"1A",X"D8",X"12",X"00",X"01",
		X"FF",X"05",X"01",X"01",X"05",X"02",X"FF",X"00",X"CD",X"6A",X"1A",X"C8",X"0C",X"01",X"01",X"FF",
		X"05",X"01",X"FF",X"05",X"02",X"01",X"00",X"CD",X"65",X"19",X"11",X"06",X"FF",X"18",X"A0",X"0A",
		X"0F",X"04",X"0C",X"FF",X"C9",X"CD",X"7B",X"1B",X"03",X"13",X"01",X"00",X"50",X"01",X"FE",X"FF",
		X"FF",X"00",X"00",X"CD",X"6A",X"1A",X"C7",X"0C",X"00",X"01",X"FF",X"01",X"03",X"F1",X"01",X"06",
		X"0F",X"00",X"CD",X"65",X"19",X"10",X"04",X"FF",X"0A",X"09",X"2A",X"04",X"04",X"04",X"FF",X"C9",
		X"CD",X"6A",X"1A",X"2F",X"13",X"02",X"01",X"FF",X"03",X"0A",X"FF",X"03",X"0F",X"01",X"00",X"CD",
		X"6A",X"1A",X"3E",X"13",X"00",X"01",X"FF",X"03",X"0A",X"01",X"03",X"0F",X"FF",X"00",X"CD",X"6A",
		X"1A",X"C8",X"0C",X"01",X"01",X"FF",X"03",X"0A",X"FF",X"03",X"0F",X"01",X"00",X"CD",X"65",X"19",
		X"10",X"0B",X"FF",X"0A",X"0F",X"04",X"1F",X"2A",X"0B",X"FF",X"C9",X"CD",X"6A",X"1A",X"C8",X"0C",
		X"01",X"01",X"00",X"01",X"2C",X"00",X"01",X"01",X"04",X"0F",X"02",X"FF",X"0F",X"06",X"01",X"00",
		X"CD",X"6A",X"1A",X"5B",X"13",X"00",X"01",X"00",X"01",X"4B",X"00",X"0F",X"06",X"FF",X"00",X"CD",
		X"65",X"19",X"01",X"08",X"FF",X"18",X"A0",X"0A",X"0C",X"FF",X"C9",X"CD",X"7B",X"1B",X"52",X"12",
		X"01",X"00",X"FF",X"FF",X"00",X"00",X"CD",X"65",X"19",X"10",X"0F",X"FF",X"04",X"06",X"2A",X"0F",
		X"0A",X"04",X"FF",X"C9",X"CD",X"33",X"1A",X"00",X"0A",X"0A",X"CD",X"33",X"1A",X"01",X"2A",X"2A",
		X"C9",X"CD",X"6A",X"1A",X"C3",X"13",X"00",X"01",X"00",X"0A",X"01",X"01",X"01",X"1C",X"00",X"09",
		X"0A",X"FF",X"00",X"CD",X"6A",X"1A",X"C8",X"0C",X"01",X"01",X"00",X"07",X"03",X"FF",X"03",X"09",
		X"FF",X"02",X"28",X"01",X"00",X"CD",X"70",X"07",X"CD",X"6A",X"1A",X"05",X"14",X"01",X"01",X"FF",
		X"01",X"01",X"F8",X"04",X"B0",X"01",X"03",X"B0",X"FF",X"02",X"B0",X"01",X"03",X"B0",X"FF",X"01",
		X"01",X"08",X"00",X"CD",X"70",X"07",X"CD",X"6A",X"1A",X"14",X"14",X"01",X"01",X"00",X"01",X"01",
		X"F8",X"FF",X"FF",X"00",X"00",X"CD",X"6A",X"1A",X"71",X"12",X"02",X"01",X"FF",X"04",X"08",X"F0",
		X"04",X"08",X"10",X"00",X"CD",X"6A",X"1A",X"71",X"12",X"02",X"01",X"FF",X"03",X"01",X"FF",X"01",
		X"06",X"03",X"00",X"CD",X"65",X"19",X"01",X"01",X"FF",X"0A",X"0A",X"02",X"00",X"00",X"59",X"FF",
		X"C9",X"CD",X"65",X"19",X"11",X"04",X"FF",X"0A",X"0A",X"02",X"00",X"00",X"6B",X"04",X"1A",X"FF",
		X"C9",X"CD",X"65",X"19",X"01",X"01",X"FF",X"0A",X"0A",X"02",X"00",X"00",X"62",X"FF",X"C9",X"CD",
		X"6A",X"1A",X"C1",X"14",X"01",X"02",X"02",X"05",X"01",X"03",X"00",X"02",X"02",X"FA",X"FF",X"05",
		X"01",X"04",X"00",X"02",X"02",X"F9",X"FF",X"05",X"01",X"05",X"00",X"02",X"02",X"F8",X"FF",X"05",
		X"01",X"06",X"00",X"02",X"02",X"F7",X"FF",X"05",X"01",X"07",X"00",X"02",X"02",X"F6",X"FF",X"05",
		X"01",X"08",X"00",X"02",X"02",X"F5",X"FF",X"00",X"CD",X"6A",X"1A",X"C1",X"14",X"01",X"02",X"02",
		X"02",X"02",X"FA",X"FF",X"05",X"01",X"03",X"00",X"02",X"02",X"F9",X"FF",X"05",X"01",X"04",X"00",
		X"02",X"02",X"F8",X"FF",X"05",X"01",X"05",X"00",X"02",X"02",X"F7",X"FF",X"05",X"01",X"07",X"00",
		X"02",X"02",X"F6",X"FF",X"05",X"01",X"06",X"00",X"02",X"02",X"F5",X"FF",X"05",X"01",X"08",X"00",
		X"00",X"CD",X"6A",X"1A",X"C7",X"0C",X"00",X"01",X"FF",X"04",X"05",X"01",X"02",X"02",X"FE",X"00",
		X"CD",X"6A",X"1A",X"09",X"15",X"01",X"02",X"00",X"06",X"01",X"03",X"00",X"02",X"01",X"FA",X"FF",
		X"06",X"01",X"04",X"00",X"02",X"01",X"F9",X"FF",X"06",X"01",X"05",X"00",X"02",X"01",X"F8",X"FF",
		X"06",X"01",X"06",X"00",X"02",X"01",X"F7",X"FF",X"06",X"01",X"07",X"00",X"02",X"01",X"F6",X"FF",
		X"06",X"01",X"08",X"00",X"02",X"01",X"F5",X"FF",X"00",X"CD",X"6A",X"1A",X"C7",X"0C",X"00",X"01",
		X"00",X"05",X"0C",X"01",X"0C",X"01",X"FF",X"00",X"CD",X"65",X"19",X"01",X"02",X"FF",X"0A",X"0C",
		X"18",X"8C",X"FF",X"C9",X"CD",X"7B",X"1B",X"35",X"15",X"01",X"09",X"03",X"01",X"FE",X"02",X"01",
		X"0A",X"01",X"01",X"EA",X"00",X"CD",X"6A",X"1A",X"C7",X"0C",X"00",X"01",X"00",X"01",X"04",X"F4",
		X"01",X"06",X"0F",X"05",X"06",X"FF",X"05",X"03",X"FF",X"05",X"01",X"FF",X"00",X"CD",X"65",X"19",
		X"01",X"09",X"FF",X"0A",X"07",X"02",X"0C",X"00",X"00",X"FF",X"C9",X"CD",X"65",X"19",X"01",X"08",
		X"FF",X"0A",X"09",X"02",X"0A",X"00",X"00",X"FF",X"C9",X"CD",X"65",X"19",X"01",X"09",X"FF",X"0A",
		X"00",X"00",X"FF",X"02",X"0F",X"FF",X"C9",X"CD",X"6A",X"1A",X"86",X"15",X"00",X"01",X"01",X"01",
		X"01",X"0F",X"05",X"05",X"FD",X"00",X"CD",X"6A",X"1A",X"C7",X"0C",X"01",X"01",X"01",X"01",X"01",
		X"F6",X"05",X"05",X"02",X"00",X"CD",X"33",X"1A",X"00",X"0A",X"0A",X"CD",X"33",X"1A",X"01",X"00",
		X"00",X"CD",X"33",X"1A",X"02",X"00",X"00",X"C9",X"CD",X"6A",X"1A",X"B7",X"15",X"02",X"01",X"FF",
		X"02",X"01",X"01",X"01",X"01",X"FE",X"00",X"CD",X"6A",X"1A",X"C7",X"0C",X"00",X"01",X"FF",X"04",
		X"10",X"01",X"FF",X"FF",X"00",X"00",X"CD",X"65",X"19",X"01",X"0B",X"00",X"0A",X"0D",X"2A",X"0B",
		X"FF",X"C9",X"CD",X"65",X"19",X"01",X"0B",X"00",X"0A",X"0D",X"2A",X"0B",X"FF",X"C9",X"CD",X"65",
		X"19",X"01",X"09",X"00",X"0A",X"0D",X"2A",X"09",X"FF",X"C9",X"CD",X"65",X"19",X"01",X"09",X"00",
		X"0A",X"0D",X"2A",X"09",X"FF",X"C9",X"CD",X"65",X"19",X"01",X"09",X"FF",X"0A",X"0D",X"02",X"0F",
		X"00",X"FF",X"FF",X"C9",X"CD",X"33",X"1A",X"00",X"0A",X"0A",X"CD",X"33",X"1A",X"01",X"18",X"18",
		X"CD",X"33",X"1A",X"02",X"00",X"00",X"C9",X"CD",X"33",X"1A",X"00",X"02",X"02",X"CD",X"33",X"1A",
		X"01",X"0A",X"0A",X"C9",X"CD",X"6A",X"1A",X"C7",X"0C",X"00",X"02",X"FF",X"02",X"01",X"00",X"FF",
		X"01",X"01",X"00",X"02",X"00",X"CD",X"6A",X"1A",X"C7",X"0C",X"00",X"02",X"FF",X"03",X"01",X"00",
		X"FF",X"01",X"01",X"00",X"03",X"00",X"CD",X"6A",X"1A",X"C7",X"0C",X"00",X"02",X"FF",X"01",X"01",
		X"00",X"03",X"03",X"01",X"00",X"FF",X"00",X"CD",X"65",X"19",X"01",X"0B",X"00",X"0A",X"0F",X"FF",
		X"C9",X"CD",X"65",X"19",X"01",X"0A",X"00",X"0A",X"0F",X"FF",X"C9",X"CD",X"65",X"19",X"01",X"09",
		X"00",X"0A",X"0F",X"FF",X"C9",X"CD",X"6A",X"1A",X"B9",X"16",X"01",X"02",X"FF",X"03",X"04",X"9D",
		X"FF",X"03",X"02",X"63",X"00",X"00",X"CD",X"6A",X"1A",X"C8",X"16",X"01",X"02",X"FF",X"03",X"04",
		X"B1",X"FF",X"03",X"02",X"4F",X"00",X"00",X"CD",X"6A",X"1A",X"C8",X"16",X"01",X"02",X"FF",X"03",
		X"02",X"C5",X"FF",X"03",X"01",X"3B",X"00",X"00",X"CD",X"6A",X"1A",X"D7",X"16",X"01",X"02",X"FF",
		X"03",X"02",X"CF",X"FF",X"03",X"01",X"31",X"00",X"00",X"CD",X"6A",X"1A",X"E6",X"16",X"02",X"01",
		X"FF",X"01",X"0C",X"FF",X"01",X"04",X"01",X"00",X"CD",X"6A",X"1A",X"F8",X"16",X"02",X"01",X"FF",
		X"01",X"06",X"FF",X"01",X"02",X"01",X"00",X"CD",X"6A",X"1A",X"0A",X"17",X"02",X"01",X"FF",X"01",
		X"03",X"FF",X"01",X"01",X"01",X"00",X"CD",X"6A",X"1A",X"C7",X"0C",X"00",X"01",X"FF",X"01",X"0C",
		X"00",X"03",X"04",X"FF",X"03",X"02",X"01",X"00",X"CD",X"6A",X"1A",X"C7",X"0C",X"00",X"01",X"FF",
		X"01",X"06",X"00",X"03",X"02",X"FF",X"03",X"01",X"01",X"00",X"CD",X"6A",X"1A",X"C7",X"0C",X"00",
		X"01",X"FF",X"01",X"03",X"00",X"01",X"03",X"FD",X"01",X"01",X"03",X"00",X"CD",X"6A",X"1A",X"2B",
		X"17",X"00",X"01",X"FF",X"05",X"01",X"FF",X"01",X"01",X"05",X"00",X"CD",X"6A",X"1A",X"C7",X"0C",
		X"01",X"01",X"FF",X"01",X"28",X"FC",X"01",X"07",X"04",X"01",X"1E",X"FA",X"01",X"05",X"06",X"01",
		X"32",X"FD",X"01",X"08",X"03",X"01",X"28",X"FB",X"01",X"0A",X"05",X"01",X"1E",X"FD",X"01",X"0C",
		X"03",X"00",X"CD",X"70",X"07",X"CD",X"6A",X"1A",X"71",X"12",X"01",X"01",X"00",X"01",X"01",X"F8",
		X"01",X"30",X"01",X"02",X"40",X"01",X"02",X"50",X"01",X"03",X"50",X"01",X"00",X"CD",X"6A",X"1A",
		X"52",X"17",X"02",X"01",X"FF",X"04",X"08",X"F0",X"04",X"08",X"10",X"00",X"CD",X"6A",X"1A",X"52",
		X"17",X"02",X"01",X"FF",X"03",X"01",X"FF",X"01",X"06",X"03",X"00",X"CD",X"65",X"19",X"10",X"06",
		X"FF",X"0A",X"0F",X"04",X"0F",X"2A",X"06",X"FF",X"C9",X"CD",X"6A",X"1A",X"C8",X"0C",X"01",X"01",
		X"00",X"06",X"0F",X"FF",X"00",X"CD",X"6A",X"1A",X"99",X"17",X"00",X"01",X"00",X"02",X"09",X"00",
		X"08",X"09",X"FF",X"00",X"CD",X"65",X"19",X"11",X"0B",X"FF",X"0A",X"0A",X"2A",X"0B",X"04",X"01",
		X"00",X"B8",X"02",X"00",X"FF",X"C9",X"CD",X"65",X"19",X"11",X"0B",X"FF",X"0A",X"0A",X"2A",X"0B",
		X"04",X"01",X"00",X"30",X"02",X"02",X"FF",X"C9",X"CD",X"6A",X"1A",X"0F",X"18",X"00",X"01",X"00",
		X"05",X"01",X"01",X"01",X"0A",X"00",X"05",X"01",X"FD",X"01",X"0F",X"00",X"05",X"01",X"03",X"01",
		X"0F",X"00",X"08",X"0A",X"FF",X"07",X"05",X"FF",X"00",X"CD",X"6A",X"1A",X"0F",X"18",X"02",X"01",
		X"00",X"0F",X"02",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"63",X"00",X"08",X"13",X"01",X"00",X"CD",
		X"6A",X"1A",X"C8",X"0C",X"01",X"01",X"00",X"05",X"01",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"63",
		X"00",X"08",X"13",X"01",X"00",X"CD",X"65",X"19",X"10",X"00",X"FF",X"0A",X"0C",X"04",X"12",X"2A",
		X"00",X"FF",X"C9",X"CD",X"6A",X"1A",X"42",X"18",X"00",X"01",X"FF",X"05",X"07",X"FF",X"05",X"0A",
		X"01",X"00",X"CD",X"6A",X"1A",X"5A",X"18",X"02",X"01",X"FF",X"01",X"10",X"F8",X"01",X"14",X"04",
		X"01",X"20",X"05",X"01",X"15",X"F7",X"01",X"1F",X"08",X"00",X"CD",X"6A",X"1A",X"C8",X"0C",X"01",
		X"01",X"FF",X"05",X"01",X"01",X"05",X"03",X"FF",X"00",X"00",X"00",X"00",X"00",X"CD",X"33",X"1A",
		X"00",X"0A",X"0A",X"C9",X"CD",X"33",X"1A",X"00",X"2A",X"2A",X"C9",X"CD",X"33",X"1A",X"00",X"0A",
		X"0A",X"CD",X"33",X"1A",X"01",X"0A",X"0A",X"C9",X"CD",X"33",X"1A",X"00",X"0A",X"0A",X"CD",X"33",
		X"1A",X"01",X"18",X"18",X"C9",X"CD",X"33",X"1A",X"00",X"0A",X"0A",X"CD",X"33",X"1A",X"01",X"2A",
		X"2A",X"C9",X"CD",X"33",X"1A",X"00",X"0A",X"0A",X"CD",X"33",X"1A",X"01",X"04",X"04",X"C9",X"CD",
		X"33",X"1A",X"00",X"0A",X"0A",X"CD",X"33",X"1A",X"01",X"00",X"00",X"C9",X"CD",X"33",X"1A",X"00",
		X"0A",X"0A",X"CD",X"33",X"1A",X"01",X"02",X"02",X"C9",X"CD",X"33",X"1A",X"00",X"0A",X"0A",X"CD",
		X"33",X"1A",X"01",X"2A",X"2A",X"CD",X"33",X"1A",X"02",X"04",X"04",X"C9",X"CD",X"33",X"1A",X"00",
		X"0A",X"0A",X"CD",X"33",X"1A",X"01",X"2A",X"2A",X"CD",X"33",X"1A",X"02",X"00",X"00",X"C9",X"CD",
		X"33",X"1A",X"00",X"0A",X"0A",X"CD",X"33",X"1A",X"01",X"00",X"00",X"CD",X"33",X"1A",X"02",X"02",
		X"02",X"C9",X"DD",X"21",X"BC",X"82",X"06",X"00",X"DD",X"7E",X"04",X"DD",X"BE",X"03",X"28",X"49",
		X"DD",X"77",X"03",X"DD",X"36",X"02",X"01",X"26",X"00",X"DD",X"6E",X"04",X"29",X"54",X"5D",X"19",
		X"19",X"11",X"E4",X"0A",X"19",X"5E",X"23",X"56",X"DD",X"E5",X"E5",X"EB",X"11",X"31",X"19",X"D5",
		X"E9",X"E1",X"DD",X"E1",X"23",X"7E",X"DD",X"77",X"00",X"23",X"7E",X"DD",X"77",X"01",X"DD",X"7E",
		X"04",X"FE",X"00",X"28",X"14",X"23",X"23",X"7E",X"FE",X"FF",X"28",X"0D",X"DD",X"E5",X"57",X"2B",
		X"5E",X"EB",X"11",X"57",X"19",X"D5",X"E9",X"DD",X"E1",X"11",X"09",X"00",X"DD",X"19",X"04",X"78",
		X"FE",X"06",X"20",X"A4",X"C9",X"50",X"1E",X"38",X"CD",X"54",X"00",X"11",X"EC",X"1C",X"19",X"E5",
		X"FD",X"E1",X"DD",X"E3",X"DD",X"CB",X"00",X"46",X"20",X"10",X"FD",X"7E",X"09",X"2F",X"4F",X"FD",
		X"5E",X"06",X"FD",X"56",X"07",X"1A",X"B1",X"12",X"18",X"0B",X"FD",X"5E",X"06",X"FD",X"56",X"07",
		X"1A",X"FD",X"A6",X"09",X"12",X"DD",X"CB",X"00",X"66",X"20",X"0A",X"FD",X"7E",X"08",X"2F",X"4F",
		X"1A",X"B1",X"12",X"18",X"05",X"1A",X"FD",X"A6",X"08",X"12",X"DD",X"4E",X"01",X"FD",X"7E",X"14",
		X"FE",X"0F",X"20",X"0A",X"79",X"CB",X"27",X"CB",X"27",X"CB",X"27",X"CB",X"27",X"4F",X"FD",X"5E",
		X"12",X"FD",X"56",X"13",X"1A",X"FD",X"A6",X"14",X"B1",X"12",X"DD",X"7E",X"02",X"4F",X"FE",X"FF",
		X"28",X"39",X"26",X"00",X"68",X"5D",X"54",X"29",X"29",X"29",X"19",X"11",X"BC",X"82",X"19",X"11",
		X"01",X"90",X"3E",X"06",X"CD",X"33",X"00",X"1A",X"E6",X"7F",X"77",X"23",X"FD",X"E5",X"D1",X"EB",
		X"79",X"CD",X"33",X"00",X"7E",X"12",X"23",X"13",X"66",X"6F",X"EB",X"72",X"21",X"03",X"90",X"7E",
		X"12",X"2B",X"7E",X"CB",X"77",X"28",X"04",X"E6",X"0F",X"13",X"12",X"DD",X"E5",X"E1",X"1E",X"03",
		X"16",X"00",X"19",X"D9",X"FD",X"E5",X"D1",X"D9",X"7E",X"FE",X"FF",X"28",X"12",X"D9",X"62",X"6B",
		X"CD",X"33",X"00",X"4E",X"23",X"46",X"D9",X"23",X"7E",X"D9",X"02",X"D9",X"23",X"18",X"E9",X"23",
		X"D1",X"E5",X"C9",X"DD",X"E1",X"48",X"DD",X"5E",X"00",X"CD",X"26",X"07",X"DD",X"5E",X"01",X"FD",
		X"E5",X"16",X"00",X"FD",X"19",X"FD",X"7E",X"00",X"77",X"23",X"FD",X"7E",X"01",X"77",X"FD",X"E1",
		X"DD",X"5E",X"02",X"FD",X"E5",X"FD",X"19",X"FD",X"7E",X"00",X"23",X"77",X"23",X"FD",X"7E",X"01",
		X"77",X"1E",X"03",X"DD",X"19",X"FD",X"E1",X"DD",X"E5",X"C9",X"FD",X"E1",X"C5",X"3E",X"06",X"90",
		X"4F",X"FD",X"5E",X"02",X"CD",X"26",X"07",X"C1",X"C5",X"E5",X"DD",X"E3",X"79",X"FE",X"00",X"28",
		X"33",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"DD",X"5E",X"02",X"DD",X"56",X"03",X"7E",X"12",X"FD",
		X"CB",X"03",X"4E",X"28",X"04",X"23",X"13",X"7E",X"12",X"FD",X"7E",X"06",X"DD",X"77",X"04",X"FD",
		X"7E",X"05",X"DD",X"77",X"05",X"AF",X"DD",X"77",X"06",X"FD",X"7E",X"04",X"DD",X"77",X"07",X"DD",
		X"E1",X"C3",X"72",X"1B",X"DD",X"35",X"04",X"28",X"05",X"DD",X"E1",X"C3",X"72",X"1B",X"FD",X"46",
		X"03",X"CB",X"48",X"26",X"00",X"DD",X"6E",X"06",X"54",X"5D",X"20",X"04",X"0E",X"03",X"18",X"03",
		X"0E",X"04",X"29",X"19",X"19",X"16",X"00",X"1E",X"05",X"19",X"EB",X"FD",X"E5",X"FD",X"19",X"DD",
		X"6E",X"00",X"DD",X"66",X"01",X"DD",X"5E",X"02",X"DD",X"56",X"03",X"CB",X"48",X"20",X"07",X"FD",
		X"7E",X"02",X"86",X"12",X"18",X"10",X"C5",X"4E",X"23",X"46",X"FD",X"6E",X"02",X"FD",X"66",X"03",
		X"09",X"C1",X"EB",X"73",X"23",X"72",X"DD",X"35",X"05",X"20",X"5D",X"DD",X"34",X"06",X"16",X"00",
		X"59",X"FD",X"19",X"FD",X"7E",X"00",X"FE",X"00",X"20",X"3C",X"DD",X"7E",X"07",X"FE",X"00",X"28",
		X"1D",X"FE",X"FF",X"28",X"03",X"DD",X"35",X"07",X"AF",X"DD",X"77",X"06",X"FD",X"E1",X"FD",X"7E",
		X"05",X"DD",X"77",X"05",X"FD",X"7E",X"06",X"DD",X"77",X"04",X"DD",X"E1",X"18",X"34",X"FD",X"E1",
		X"DD",X"E1",X"C1",X"3E",X"06",X"90",X"21",X"5C",X"1E",X"16",X"00",X"5F",X"19",X"3A",X"1F",X"83",
		X"B6",X"32",X"1F",X"83",X"18",X"1D",X"FD",X"7E",X"01",X"DD",X"77",X"04",X"FD",X"7E",X"00",X"DD",
		X"77",X"05",X"FD",X"E1",X"DD",X"E1",X"18",X"0A",X"FD",X"7E",X"01",X"DD",X"77",X"04",X"FD",X"E1",
		X"DD",X"E1",X"C1",X"FD",X"6E",X"00",X"FD",X"66",X"01",X"E5",X"C9",X"FD",X"E1",X"C5",X"3E",X"06",
		X"90",X"4F",X"FD",X"5E",X"02",X"CD",X"26",X"07",X"59",X"C1",X"C5",X"E5",X"DD",X"E3",X"79",X"FE",
		X"00",X"28",X"48",X"C5",X"4B",X"16",X"00",X"1E",X"09",X"19",X"71",X"C1",X"2B",X"DD",X"75",X"00",
		X"DD",X"74",X"01",X"DD",X"75",X"02",X"DD",X"74",X"03",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"DD",
		X"5E",X"02",X"DD",X"56",X"03",X"7E",X"12",X"FD",X"7E",X"05",X"DD",X"77",X"04",X"FD",X"7E",X"04",
		X"DD",X"77",X"05",X"AF",X"DD",X"77",X"06",X"FD",X"7E",X"03",X"DD",X"77",X"07",X"DD",X"7E",X"08",
		X"DD",X"4E",X"09",X"CD",X"44",X"07",X"DD",X"E1",X"C3",X"A0",X"1C",X"DD",X"35",X"04",X"28",X"05",
		X"DD",X"E1",X"C3",X"A0",X"1C",X"26",X"00",X"DD",X"6E",X"06",X"54",X"5D",X"0E",X"03",X"19",X"19",
		X"16",X"00",X"1E",X"04",X"19",X"EB",X"FD",X"E5",X"FD",X"19",X"DD",X"6E",X"00",X"DD",X"66",X"01",
		X"DD",X"5E",X"02",X"DD",X"56",X"03",X"FD",X"7E",X"02",X"CB",X"7F",X"CA",X"1E",X"1C",X"86",X"CB",
		X"7F",X"CA",X"2B",X"1C",X"CB",X"77",X"CA",X"2B",X"1C",X"C6",X"C0",X"C3",X"2B",X"1C",X"86",X"CB",
		X"7F",X"CA",X"2B",X"1C",X"CB",X"77",X"CA",X"2B",X"1C",X"C6",X"40",X"12",X"C5",X"DD",X"4E",X"09",
		X"CD",X"44",X"07",X"C1",X"DD",X"35",X"05",X"20",X"5D",X"DD",X"34",X"06",X"16",X"00",X"59",X"FD",
		X"19",X"FD",X"7E",X"00",X"FE",X"00",X"20",X"3C",X"DD",X"7E",X"07",X"FE",X"00",X"28",X"1D",X"FE",
		X"FF",X"28",X"03",X"DD",X"35",X"07",X"AF",X"DD",X"77",X"06",X"FD",X"E1",X"FD",X"7E",X"04",X"DD",
		X"77",X"05",X"FD",X"7E",X"05",X"DD",X"77",X"04",X"DD",X"E1",X"18",X"34",X"FD",X"E1",X"DD",X"E1",
		X"C1",X"3E",X"06",X"90",X"21",X"5C",X"1E",X"16",X"00",X"5F",X"19",X"3A",X"1F",X"83",X"B6",X"32",
		X"1F",X"83",X"18",X"1D",X"FD",X"7E",X"01",X"DD",X"77",X"04",X"FD",X"7E",X"00",X"DD",X"77",X"05",
		X"FD",X"E1",X"DD",X"E1",X"18",X"0A",X"FD",X"7E",X"01",X"DD",X"77",X"04",X"FD",X"E1",X"DD",X"E1",
		X"C1",X"FD",X"6E",X"00",X"FD",X"66",X"01",X"E5",X"C9",X"3E",X"06",X"90",X"6F",X"26",X"00",X"54",
		X"5D",X"29",X"19",X"FD",X"21",X"F2",X"82",X"EB",X"FD",X"19",X"FD",X"6E",X"00",X"FD",X"66",X"01",
		X"FD",X"7E",X"02",X"96",X"D8",X"3E",X"01",X"77",X"C9",X"DD",X"E1",X"FD",X"E5",X"E1",X"DD",X"5E",
		X"00",X"16",X"00",X"19",X"E5",X"68",X"26",X"00",X"54",X"5D",X"29",X"19",X"11",X"F2",X"82",X"19",
		X"D1",X"1A",X"77",X"13",X"23",X"1A",X"77",X"DD",X"23",X"DD",X"E5",X"C9",X"00",X"80",X"01",X"80",
		X"06",X"80",X"07",X"80",X"F7",X"FE",X"08",X"80",X"0B",X"80",X"0C",X"80",X"0D",X"80",X"0E",X"80",
		X"F0",X"00",X"48",X"80",X"59",X"80",X"6A",X"80",X"7B",X"80",X"8C",X"80",X"44",X"80",X"55",X"80",
		X"66",X"80",X"77",X"80",X"88",X"80",X"3E",X"82",X"F4",X"82",X"49",X"80",X"5A",X"80",X"6B",X"80",
		X"7C",X"80",X"8D",X"80",X"02",X"80",X"03",X"80",X"06",X"80",X"07",X"80",X"EF",X"FD",X"09",X"80",
		X"0B",X"80",X"0C",X"80",X"0D",X"80",X"0E",X"80",X"0F",X"00",X"9D",X"80",X"AE",X"80",X"BF",X"80",
		X"D0",X"80",X"E1",X"80",X"99",X"80",X"AA",X"80",X"BB",X"80",X"CC",X"80",X"DD",X"80",X"3F",X"82",
		X"F7",X"82",X"9E",X"80",X"AF",X"80",X"C0",X"80",X"D1",X"80",X"E2",X"80",X"04",X"80",X"05",X"80",
		X"06",X"80",X"07",X"80",X"DF",X"FB",X"0A",X"80",X"0B",X"80",X"0C",X"80",X"0D",X"80",X"0F",X"80",
		X"F0",X"00",X"F2",X"80",X"03",X"81",X"14",X"81",X"25",X"81",X"36",X"81",X"EE",X"80",X"FF",X"80",
		X"10",X"81",X"21",X"81",X"32",X"81",X"40",X"82",X"FA",X"82",X"F3",X"80",X"04",X"81",X"15",X"81",
		X"26",X"81",X"37",X"81",X"10",X"80",X"11",X"80",X"16",X"80",X"17",X"80",X"F7",X"FE",X"18",X"80",
		X"1B",X"80",X"1C",X"80",X"1D",X"80",X"1E",X"80",X"F0",X"00",X"47",X"81",X"58",X"81",X"69",X"81",
		X"7A",X"81",X"8B",X"81",X"43",X"81",X"54",X"81",X"65",X"81",X"76",X"81",X"87",X"81",X"41",X"82",
		X"FD",X"82",X"48",X"81",X"59",X"81",X"6A",X"81",X"7B",X"81",X"8C",X"81",X"12",X"80",X"13",X"80",
		X"16",X"80",X"17",X"80",X"EF",X"FD",X"19",X"80",X"1B",X"80",X"1C",X"80",X"1D",X"80",X"1E",X"80",
		X"0F",X"00",X"9C",X"81",X"AD",X"81",X"BE",X"81",X"CF",X"81",X"E0",X"81",X"98",X"81",X"A9",X"81",
		X"BA",X"81",X"CB",X"81",X"DC",X"81",X"42",X"82",X"00",X"83",X"9D",X"81",X"AE",X"81",X"BF",X"81",
		X"D0",X"81",X"E1",X"81",X"14",X"80",X"15",X"80",X"16",X"80",X"17",X"80",X"DF",X"FB",X"1A",X"80",
		X"1B",X"80",X"1C",X"80",X"1D",X"80",X"1F",X"80",X"F0",X"00",X"F1",X"81",X"02",X"82",X"13",X"82",
		X"24",X"82",X"35",X"82",X"ED",X"81",X"FE",X"81",X"0F",X"82",X"20",X"82",X"31",X"82",X"43",X"82",
		X"03",X"83",X"F2",X"81",X"03",X"82",X"14",X"82",X"25",X"82",X"36",X"82",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"01",X"02",X"04",X"08",
		X"10",X"20",X"D1",X"0F",X"60",X"0F",X"EE",X"0E",X"83",X"0E",X"18",X"0E",X"B2",X"0D",X"4D",X"0D",
		X"EE",X"0C",X"8E",X"0C",X"34",X"0C",X"DA",X"0B",X"84",X"0B",X"2F",X"0B",X"DF",X"0A",X"8F",X"0A",
		X"43",X"0A",X"F7",X"09",X"B0",X"09",X"68",X"09",X"24",X"09",X"E1",X"08",X"A1",X"08",X"61",X"08",
		X"25",X"08",X"E9",X"07",X"B0",X"07",X"77",X"07",X"42",X"07",X"0C",X"07",X"D9",X"06",X"A7",X"06",
		X"77",X"06",X"47",X"06",X"15",X"06",X"ED",X"05",X"C3",X"05",X"98",X"05",X"6F",X"05",X"47",X"05",
		X"21",X"05",X"FB",X"04",X"D8",X"04",X"B4",X"04",X"92",X"04",X"70",X"04",X"50",X"04",X"31",X"04",
		X"13",X"04",X"F4",X"03",X"D8",X"03",X"BC",X"03",X"9F",X"03",X"86",X"03",X"6D",X"03",X"53",X"03",
		X"3B",X"03",X"24",X"03",X"0D",X"03",X"F6",X"02",X"E1",X"02",X"CC",X"02",X"B8",X"02",X"A4",X"02",
		X"91",X"02",X"7E",X"02",X"6C",X"02",X"5A",X"02",X"49",X"02",X"38",X"02",X"28",X"02",X"18",X"02",
		X"09",X"02",X"FA",X"01",X"EC",X"01",X"DE",X"01",X"D1",X"01",X"C3",X"01",X"B7",X"01",X"AA",X"01",
		X"9E",X"01",X"92",X"01",X"86",X"01",X"7B",X"01",X"71",X"01",X"66",X"01",X"5C",X"01",X"52",X"01",
		X"48",X"01",X"3F",X"01",X"36",X"01",X"2D",X"01",X"25",X"01",X"1C",X"01",X"14",X"01",X"0C",X"01",
		X"04",X"01",X"FD",X"00",X"F6",X"00",X"EF",X"00",X"E8",X"00",X"E1",X"00",X"DB",X"00",X"D5",X"00",
		X"CF",X"00",X"C9",X"00",X"C4",X"00",X"BE",X"00",X"B8",X"00",X"B3",X"00",X"AE",X"00",X"A9",X"00",
		X"A4",X"00",X"9F",X"00",X"9B",X"00",X"96",X"00",X"92",X"00",X"8E",X"00",X"8A",X"00",X"86",X"00",
		X"82",X"00",X"7F",X"00",X"7B",X"00",X"77",X"00",X"74",X"00",X"71",X"00",X"6D",X"00",X"6A",X"00",
		X"67",X"00",X"64",X"00",X"62",X"00",X"5F",X"00",X"5C",X"00",X"59",X"00",X"56",X"00",X"54",X"00",
		X"52",X"00",X"50",X"00",X"4E",X"00",X"4B",X"00",X"49",X"00",X"47",X"00",X"45",X"00",X"43",X"00",
		X"41",X"00",X"3F",X"00",X"3D",X"00",X"3B",X"00",X"39",X"00",X"38",X"00",X"37",X"00",X"35",X"00",
		X"33",X"00",X"32",X"00",X"31",X"00",X"2F",X"00",X"2D",X"00",X"2C",X"00",X"2B",X"00",X"2A",X"00",
		X"29",X"00",X"27",X"00",X"26",X"00",X"26",X"00",X"25",X"00",X"24",X"00",X"23",X"00",X"22",X"00",
		X"21",X"00",X"20",X"00",X"1F",X"00",X"1E",X"00",X"1D",X"00",X"1C",X"00",X"1B",X"00",X"1B",X"00",
		X"1A",X"00",X"19",X"00",X"18",X"00",X"18",X"00",X"17",X"00",X"16",X"00",X"15",X"00",X"15",X"00",
		X"14",X"00",X"14",X"00",X"13",X"00",X"13",X"00",X"12",X"00",X"12",X"00",X"11",X"00",X"11",X"00",
		X"10",X"00",X"52",X"6F",X"62",X"65",X"72",X"74",X"20",X"4D",X"20",X"4C",X"69",X"62",X"62",X"65",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
