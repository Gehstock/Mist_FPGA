library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity sbagman_program is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of sbagman_program is
	type rom is array(0 to  24575) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"C3",X"A8",X"EC",X"9B",X"AE",X"7B",X"04",X"80",X"E4",X"0E",X"00",X"11",X"4F",X"92",X"60",X"A3",
		X"C4",X"F7",X"04",X"02",X"F7",X"FE",X"03",X"19",X"06",X"13",X"80",X"00",X"6D",X"9F",X"42",X"02",
		X"E2",X"16",X"00",X"08",X"97",X"73",X"58",X"00",X"B6",X"1F",X"00",X"08",X"85",X"57",X"00",X"01",
		X"F2",X"5B",X"01",X"00",X"A2",X"5C",X"00",X"10",X"F3",X"F5",X"C5",X"D5",X"E5",X"DD",X"E5",X"FD",
		X"E5",X"D9",X"C5",X"D5",X"E5",X"08",X"F5",X"CD",X"2E",X"D3",X"AF",X"32",X"00",X"A0",X"CD",X"91",
		X"CA",X"CD",X"65",X"15",X"3A",X"8C",X"62",X"FE",X"01",X"CC",X"89",X"16",X"3A",X"42",X"61",X"3C",
		X"32",X"42",X"61",X"3A",X"32",X"63",X"FE",X"01",X"CC",X"9E",X"11",X"3A",X"32",X"63",X"FE",X"01",
		X"CA",X"12",X"05",X"3A",X"74",X"62",X"FE",X"01",X"28",X"05",X"3A",X"ED",X"61",X"FE",X"00",X"CC",
		X"E8",X"0F",X"3A",X"6F",X"62",X"FE",X"01",X"CA",X"15",X"05",X"3A",X"10",X"62",X"FE",X"01",X"20",
		X"22",X"3A",X"54",X"60",X"FE",X"00",X"28",X"1B",X"3A",X"F2",X"61",X"FE",X"01",X"28",X"14",X"3A",
		X"ED",X"61",X"FE",X"01",X"28",X"0D",X"3A",X"82",X"65",X"FE",X"E9",X"D2",X"15",X"05",X"FE",X"0F",
		X"DA",X"15",X"05",X"3A",X"00",X"B8",X"21",X"A0",X"65",X"11",X"00",X"98",X"01",X"20",X"00",X"ED",
		X"B0",X"CD",X"09",X"CF",X"3A",X"C1",X"62",X"FE",X"00",X"28",X"04",X"3D",X"32",X"C1",X"62",X"CD",
		X"A7",X"CF",X"3A",X"51",X"63",X"FE",X"01",X"CC",X"E7",X"DB",X"3A",X"43",X"61",X"3C",X"32",X"43",
		X"61",X"CD",X"92",X"11",X"3A",X"6D",X"62",X"3C",X"32",X"6D",X"62",X"FD",X"21",X"B8",X"65",X"3A",
		X"0D",X"60",X"47",X"3A",X"99",X"60",X"B8",X"28",X"05",X"CD",X"8C",X"11",X"18",X"0B",X"DD",X"21",
		X"94",X"65",X"FD",X"21",X"B8",X"65",X"CD",X"D7",X"D6",X"FD",X"21",X"BC",X"65",X"3A",X"0D",X"60",
		X"47",X"3A",X"9A",X"60",X"B8",X"28",X"05",X"CD",X"8C",X"11",X"18",X"0B",X"DD",X"21",X"98",X"65",
		X"FD",X"21",X"BC",X"65",X"CD",X"D7",X"D6",X"3A",X"43",X"63",X"FE",X"01",X"28",X"0B",X"3A",X"53",
		X"60",X"FE",X"01",X"CA",X"EA",X"04",X"CD",X"80",X"05",X"3A",X"51",X"61",X"FE",X"01",X"CA",X"EA",
		X"04",X"CD",X"31",X"17",X"3A",X"00",X"B8",X"3A",X"AC",X"62",X"3C",X"32",X"AC",X"62",X"CD",X"AE",
		X"FE",X"CD",X"D3",X"E9",X"CD",X"6F",X"E7",X"CD",X"16",X"E6",X"CD",X"38",X"05",X"CD",X"37",X"C6",
		X"CD",X"B3",X"CE",X"CD",X"C4",X"D3",X"3A",X"00",X"B8",X"3A",X"71",X"62",X"32",X"72",X"62",X"3A",
		X"0C",X"57",X"32",X"71",X"62",X"FD",X"21",X"56",X"61",X"DD",X"21",X"94",X"65",X"11",X"48",X"61",
		X"CD",X"4C",X"05",X"FD",X"21",X"57",X"61",X"DD",X"21",X"98",X"65",X"11",X"49",X"61",X"CD",X"4C",
		X"05",X"2A",X"38",X"60",X"DD",X"21",X"EB",X"61",X"FD",X"21",X"3A",X"60",X"DD",X"7E",X"00",X"DD",
		X"A6",X"01",X"08",X"11",X"97",X"65",X"3A",X"99",X"60",X"47",X"3A",X"EB",X"61",X"FE",X"00",X"C4",
		X"77",X"CF",X"2A",X"78",X"60",X"DD",X"21",X"EC",X"61",X"FD",X"21",X"7A",X"60",X"11",X"9B",X"65",
		X"3E",X"00",X"08",X"3A",X"9A",X"60",X"47",X"3A",X"EC",X"61",X"FE",X"00",X"C4",X"77",X"CF",X"3A",
		X"ED",X"61",X"FE",X"00",X"CC",X"99",X"F1",X"CD",X"5E",X"11",X"CD",X"E8",X"08",X"3A",X"2C",X"60",
		X"FE",X"01",X"28",X"06",X"CD",X"84",X"08",X"3A",X"00",X"B8",X"CD",X"C2",X"08",X"AF",X"32",X"2C",
		X"60",X"3A",X"00",X"B8",X"CD",X"3E",X"F8",X"CD",X"92",X"07",X"CD",X"C6",X"CB",X"CD",X"D5",X"07",
		X"CD",X"82",X"09",X"CD",X"10",X"09",X"3A",X"00",X"B8",X"CD",X"9F",X"D5",X"CD",X"D6",X"D5",X"3A",
		X"ED",X"61",X"FE",X"00",X"CC",X"A6",X"09",X"3A",X"00",X"B8",X"CD",X"8A",X"DA",X"3A",X"26",X"60",
		X"E6",X"60",X"FE",X"00",X"28",X"17",X"3A",X"83",X"65",X"F5",X"3D",X"32",X"83",X"65",X"CD",X"A7",
		X"EA",X"F1",X"32",X"83",X"65",X"3A",X"C7",X"61",X"FE",X"00",X"CC",X"14",X"0E",X"CD",X"A7",X"EA",
		X"3A",X"4E",X"60",X"FE",X"00",X"20",X"57",X"CD",X"64",X"D4",X"3A",X"14",X"60",X"FE",X"01",X"28",
		X"0E",X"3A",X"E5",X"62",X"FE",X"01",X"28",X"07",X"3A",X"08",X"60",X"FE",X"01",X"28",X"3F",X"3A",
		X"BD",X"62",X"FE",X"00",X"20",X"38",X"3A",X"D2",X"62",X"FE",X"01",X"28",X"31",X"3A",X"95",X"62",
		X"FE",X"00",X"20",X"2A",X"3A",X"B0",X"62",X"FE",X"01",X"28",X"07",X"3A",X"AF",X"62",X"FE",X"01",
		X"28",X"1C",X"3A",X"14",X"60",X"FE",X"01",X"20",X"07",X"3A",X"12",X"60",X"FE",X"01",X"20",X"0E",
		X"FD",X"21",X"47",X"60",X"DD",X"21",X"80",X"65",X"CD",X"C6",X"0B",X"3A",X"00",X"B8",X"CD",X"C6",
		X"10",X"CD",X"0C",X"11",X"3E",X"01",X"32",X"8A",X"62",X"3A",X"0D",X"60",X"32",X"98",X"60",X"21",
		X"14",X"60",X"DD",X"21",X"80",X"65",X"CD",X"B1",X"0A",X"3A",X"00",X"B8",X"3A",X"F2",X"61",X"FE",
		X"00",X"20",X"60",X"3A",X"D2",X"62",X"FE",X"01",X"28",X"59",X"3A",X"E5",X"62",X"FE",X"01",X"28",
		X"52",X"3A",X"BD",X"62",X"FE",X"01",X"28",X"4B",X"3A",X"AF",X"62",X"FE",X"01",X"28",X"44",X"3A",
		X"0D",X"60",X"32",X"98",X"60",X"21",X"08",X"60",X"7E",X"FE",X"00",X"28",X"1F",X"3A",X"0D",X"60",
		X"FE",X"04",X"20",X"18",X"3A",X"13",X"60",X"FE",X"01",X"28",X"11",X"3A",X"14",X"60",X"FE",X"01",
		X"28",X"0A",X"3A",X"C7",X"61",X"FE",X"01",X"E5",X"CC",X"4B",X"D6",X"E1",X"FD",X"21",X"4D",X"60",
		X"DD",X"21",X"80",X"65",X"3A",X"14",X"60",X"4F",X"3A",X"13",X"60",X"06",X"19",X"CD",X"82",X"0B",
		X"3A",X"00",X"B8",X"3A",X"0D",X"60",X"32",X"98",X"60",X"DD",X"21",X"80",X"65",X"FD",X"21",X"14",
		X"60",X"CD",X"DB",X"0A",X"DD",X"21",X"80",X"65",X"21",X"14",X"60",X"CD",X"40",X"0A",X"3A",X"56",
		X"61",X"FE",X"00",X"20",X"63",X"3A",X"D6",X"62",X"FE",X"01",X"28",X"3B",X"3A",X"11",X"62",X"FE",
		X"00",X"20",X"34",X"3A",X"C4",X"62",X"FE",X"00",X"20",X"2D",X"3A",X"9D",X"62",X"FE",X"00",X"20",
		X"26",X"3A",X"B6",X"62",X"FE",X"01",X"28",X"0E",X"3A",X"B5",X"62",X"FE",X"01",X"28",X"18",X"3A",
		X"48",X"61",X"FE",X"01",X"28",X"11",X"3A",X"3B",X"60",X"FE",X"01",X"20",X"07",X"3A",X"12",X"60",
		X"FE",X"01",X"20",X"03",X"CD",X"C0",X"11",X"FD",X"21",X"57",X"60",X"FD",X"22",X"93",X"60",X"2A",
		X"38",X"60",X"22",X"44",X"60",X"21",X"35",X"60",X"FD",X"21",X"27",X"60",X"DD",X"21",X"94",X"65",
		X"3A",X"37",X"60",X"FE",X"01",X"C4",X"BB",X"05",X"3A",X"57",X"61",X"FE",X"00",X"20",X"69",X"3A",
		X"12",X"62",X"FE",X"00",X"20",X"3B",X"3A",X"DA",X"62",X"FE",X"01",X"28",X"34",X"3A",X"CB",X"62",
		X"FE",X"00",X"20",X"2D",X"3A",X"A5",X"62",X"FE",X"00",X"20",X"26",X"3A",X"BA",X"62",X"FE",X"01",
		X"28",X"0E",X"3A",X"B9",X"62",X"FE",X"01",X"28",X"18",X"3A",X"49",X"61",X"FE",X"01",X"28",X"11",
		X"3A",X"7B",X"60",X"FE",X"01",X"20",X"07",X"3A",X"12",X"60",X"FE",X"01",X"20",X"03",X"CD",X"EC",
		X"11",X"2A",X"78",X"60",X"22",X"44",X"60",X"FD",X"21",X"97",X"60",X"FD",X"22",X"93",X"60",X"2A",
		X"78",X"60",X"22",X"44",X"60",X"21",X"75",X"60",X"FD",X"21",X"67",X"60",X"DD",X"21",X"98",X"65",
		X"3A",X"77",X"60",X"FE",X"01",X"C4",X"BB",X"05",X"3A",X"9A",X"60",X"32",X"98",X"60",X"21",X"7B",
		X"60",X"DD",X"21",X"98",X"65",X"CD",X"B1",X"0A",X"3A",X"00",X"B8",X"3A",X"97",X"60",X"3C",X"32",
		X"97",X"60",X"FD",X"21",X"8F",X"60",X"21",X"77",X"60",X"DD",X"21",X"98",X"65",X"3A",X"EC",X"61",
		X"FE",X"01",X"28",X"27",X"3A",X"DA",X"62",X"FE",X"01",X"28",X"20",X"3A",X"CB",X"62",X"FE",X"00",
		X"20",X"19",X"3A",X"ED",X"62",X"FE",X"01",X"28",X"12",X"3A",X"9A",X"60",X"32",X"98",X"60",X"3A",
		X"7B",X"60",X"4F",X"3A",X"7A",X"60",X"06",X"26",X"CD",X"82",X"0B",X"3A",X"99",X"60",X"32",X"98",
		X"60",X"21",X"3B",X"60",X"DD",X"21",X"94",X"65",X"CD",X"B1",X"0A",X"3A",X"57",X"60",X"3C",X"32",
		X"57",X"60",X"FD",X"21",X"4F",X"60",X"21",X"37",X"60",X"DD",X"21",X"94",X"65",X"3A",X"EB",X"61",
		X"FE",X"01",X"28",X"27",X"3A",X"D6",X"62",X"FE",X"01",X"28",X"20",X"3A",X"C4",X"62",X"FE",X"00",
		X"20",X"19",X"3A",X"E9",X"62",X"FE",X"01",X"28",X"12",X"3A",X"99",X"60",X"32",X"98",X"60",X"3A",
		X"3B",X"60",X"4F",X"3A",X"3A",X"60",X"06",X"26",X"CD",X"82",X"0B",X"CD",X"E0",X"E3",X"CD",X"6D",
		X"E3",X"CD",X"89",X"E3",X"CD",X"30",X"E6",X"CD",X"B4",X"E1",X"CD",X"C0",X"E1",X"CD",X"CC",X"E1",
		X"CD",X"69",X"E8",X"CD",X"3C",X"E0",X"CD",X"42",X"DF",X"CD",X"13",X"DD",X"CD",X"0C",X"D6",X"3E",
		X"01",X"32",X"7F",X"62",X"CD",X"ED",X"F3",X"3A",X"00",X"B8",X"CD",X"11",X"D5",X"3A",X"F1",X"61",
		X"FE",X"00",X"CC",X"15",X"0F",X"3A",X"ED",X"61",X"FE",X"01",X"CD",X"61",X"E8",X"3A",X"5B",X"63",
		X"3C",X"32",X"5B",X"63",X"FE",X"0A",X"38",X"0A",X"AF",X"32",X"5B",X"63",X"CD",X"2E",X"16",X"CD",
		X"0F",X"56",X"CD",X"89",X"16",X"CD",X"4D",X"D3",X"3A",X"56",X"63",X"FE",X"00",X"C0",X"3A",X"00",
		X"B8",X"3E",X"01",X"32",X"00",X"A0",X"ED",X"56",X"F1",X"08",X"E1",X"D1",X"C1",X"D9",X"FD",X"E1",
		X"DD",X"E1",X"E1",X"D1",X"C1",X"F1",X"FB",X"C9",X"3A",X"59",X"61",X"47",X"3A",X"34",X"63",X"B0",
		X"FE",X"00",X"C8",X"3A",X"9F",X"65",X"3C",X"3C",X"32",X"9F",X"65",X"C9",X"FD",X"7E",X"00",X"FE",
		X"00",X"C8",X"2A",X"54",X"61",X"3A",X"53",X"61",X"FE",X"07",X"20",X"11",X"7E",X"FE",X"FF",X"28",
		X"14",X"DD",X"77",X"00",X"23",X"22",X"54",X"61",X"AF",X"32",X"53",X"61",X"C9",X"3A",X"53",X"61",
		X"3C",X"32",X"53",X"61",X"C9",X"3E",X"31",X"DD",X"77",X"00",X"AF",X"FD",X"77",X"00",X"12",X"C9",
		X"FD",X"21",X"51",X"61",X"DD",X"21",X"80",X"65",X"2A",X"54",X"61",X"FD",X"7E",X"00",X"FE",X"00",
		X"C8",X"3A",X"53",X"61",X"FE",X"07",X"20",X"11",X"7E",X"FE",X"FF",X"28",X"14",X"DD",X"77",X"00",
		X"23",X"22",X"54",X"61",X"AF",X"32",X"53",X"61",X"C9",X"3A",X"53",X"61",X"3C",X"32",X"53",X"61",
		X"C9",X"3E",X"01",X"32",X"52",X"61",X"C9",X"94",X"65",X"98",X"65",X"FD",X"7E",X"00",X"E6",X"10",
		X"FE",X"10",X"28",X"15",X"FD",X"7E",X"00",X"E6",X"20",X"FE",X"20",X"C0",X"E5",X"2A",X"44",X"60",
		X"7E",X"FE",X"FF",X"E1",X"C0",X"06",X"00",X"18",X"0C",X"E5",X"2A",X"44",X"60",X"2B",X"7E",X"FE",
		X"FF",X"E1",X"C0",X"06",X"80",X"7E",X"FE",X"0B",X"20",X"05",X"3E",X"01",X"77",X"18",X"02",X"3C",
		X"77",X"7E",X"FE",X"01",X"C8",X"FE",X"03",X"C8",X"FE",X"05",X"C8",X"FE",X"08",X"C8",X"FE",X"0A",
		X"CC",X"31",X"06",X"FE",X"02",X"CC",X"31",X"06",X"FE",X"04",X"CC",X"31",X"06",X"FE",X"07",X"CC",
		X"31",X"06",X"FE",X"09",X"CC",X"31",X"06",X"FE",X"06",X"20",X"09",X"3E",X"27",X"DD",X"77",X"00",
		X"CD",X"31",X"06",X"C9",X"FE",X"0B",X"20",X"08",X"3E",X"A7",X"DD",X"77",X"00",X"CD",X"31",X"06",
		X"C9",X"F5",X"C5",X"3A",X"F5",X"61",X"FE",X"00",X"20",X"14",X"3A",X"CF",X"61",X"FE",X"00",X"20",
		X"0D",X"3A",X"F3",X"61",X"FE",X"00",X"20",X"06",X"21",X"7B",X"D9",X"CD",X"84",X"EC",X"C1",X"F1",
		X"F5",X"78",X"FE",X"80",X"20",X"14",X"DD",X"7E",X"03",X"3D",X"DD",X"77",X"03",X"AF",X"FD",X"2A",
		X"93",X"60",X"FD",X"77",X"00",X"CD",X"C9",X"0F",X"F1",X"C9",X"DD",X"7E",X"03",X"3C",X"DD",X"77",
		X"03",X"AF",X"FD",X"2A",X"93",X"60",X"FD",X"77",X"00",X"CD",X"C9",X"0F",X"F1",X"C9",X"FD",X"7E",
		X"00",X"E6",X"80",X"FE",X"80",X"20",X"0F",X"E5",X"2A",X"44",X"60",X"CD",X"71",X"0D",X"E1",X"3A",
		X"0B",X"60",X"FE",X"02",X"28",X"1A",X"FD",X"7E",X"00",X"E6",X"40",X"FE",X"40",X"C0",X"E5",X"2A",
		X"44",X"60",X"CD",X"CC",X"0D",X"E1",X"3A",X"0B",X"60",X"FE",X"02",X"C0",X"06",X"80",X"28",X"02",
		X"06",X"00",X"7E",X"FE",X"0B",X"20",X"05",X"3E",X"01",X"77",X"18",X"02",X"3C",X"77",X"7E",X"FE",
		X"02",X"28",X"2B",X"FE",X"05",X"28",X"27",X"FE",X"09",X"28",X"23",X"FE",X"FF",X"28",X"1F",X"FE",
		X"04",X"CA",X"EE",X"06",X"FE",X"06",X"CC",X"22",X"07",X"FE",X"08",X"CC",X"22",X"07",X"FE",X"0A",
		X"CC",X"22",X"07",X"FE",X"01",X"20",X"19",X"3E",X"31",X"B0",X"DD",X"77",X"00",X"C9",X"F5",X"C5",
		X"47",X"3A",X"64",X"61",X"B8",X"30",X"03",X"C1",X"F1",X"C9",X"C1",X"F1",X"CD",X"22",X"07",X"C9",
		X"FE",X"03",X"20",X"07",X"3E",X"30",X"B0",X"DD",X"77",X"00",X"C9",X"FE",X"07",X"20",X"07",X"3E",
		X"2E",X"B0",X"DD",X"77",X"00",X"C9",X"FE",X"FF",X"20",X"07",X"3E",X"30",X"B0",X"DD",X"77",X"00",
		X"C9",X"C9",X"F5",X"C5",X"3A",X"F5",X"61",X"FE",X"00",X"20",X"14",X"3A",X"CF",X"61",X"FE",X"00",
		X"20",X"0D",X"3A",X"F3",X"61",X"FE",X"00",X"20",X"06",X"21",X"9F",X"D9",X"CD",X"84",X"EC",X"C1",
		X"AF",X"FD",X"2A",X"93",X"60",X"FD",X"77",X"00",X"78",X"FE",X"80",X"28",X"19",X"DD",X"7E",X"02",
		X"3C",X"DD",X"77",X"02",X"FE",X"F0",X"20",X"0C",X"3E",X"01",X"DD",X"77",X"02",X"3A",X"98",X"60",
		X"3C",X"32",X"98",X"60",X"F1",X"C9",X"DD",X"7E",X"02",X"3D",X"DD",X"77",X"02",X"FE",X"01",X"20",
		X"0C",X"3E",X"F0",X"DD",X"77",X"02",X"3A",X"98",X"60",X"3D",X"32",X"98",X"60",X"AF",X"FD",X"2A",
		X"93",X"60",X"FD",X"77",X"00",X"F1",X"C9",X"AF",X"32",X"1C",X"60",X"32",X"1D",X"60",X"32",X"1E",
		X"60",X"C9",X"21",X"1C",X"60",X"DD",X"21",X"8A",X"65",X"FD",X"21",X"82",X"65",X"11",X"04",X"00",
		X"7E",X"FE",X"01",X"28",X"01",X"C9",X"3E",X"01",X"32",X"30",X"60",X"3A",X"26",X"60",X"E6",X"08",
		X"FE",X"08",X"CC",X"C9",X"07",X"3A",X"26",X"60",X"E6",X"10",X"FE",X"10",X"CC",X"CF",X"07",X"3E",
		X"01",X"32",X"29",X"60",X"3D",X"32",X"2F",X"60",X"C9",X"3E",X"01",X"32",X"2D",X"60",X"C9",X"3E",
		X"01",X"32",X"2E",X"60",X"C9",X"3A",X"30",X"60",X"FE",X"01",X"C0",X"3A",X"2D",X"60",X"FE",X"01",
		X"CC",X"10",X"08",X"3A",X"2E",X"60",X"FE",X"01",X"CC",X"20",X"08",X"3A",X"2F",X"60",X"3C",X"FE",
		X"04",X"28",X"04",X"32",X"2F",X"60",X"C9",X"AF",X"32",X"2D",X"60",X"32",X"2E",X"60",X"32",X"30",
		X"60",X"32",X"29",X"60",X"32",X"25",X"60",X"CD",X"87",X"07",X"3E",X"20",X"32",X"80",X"65",X"C9",
		X"CD",X"30",X"08",X"CD",X"70",X"08",X"FD",X"7E",X"00",X"3D",X"3D",X"3D",X"FD",X"77",X"00",X"C9",
		X"CD",X"30",X"08",X"CD",X"53",X"08",X"FD",X"7E",X"00",X"3C",X"3C",X"3C",X"FD",X"77",X"00",X"C9",
		X"11",X"4F",X"08",X"3A",X"2F",X"60",X"FE",X"04",X"C8",X"83",X"5F",X"7A",X"CE",X"00",X"57",X"1A",
		X"47",X"3A",X"80",X"65",X"E6",X"08",X"B0",X"32",X"80",X"65",X"AF",X"32",X"25",X"60",X"C9",X"1D",
		X"1D",X"1D",X"1D",X"06",X"20",X"C5",X"2A",X"09",X"60",X"CD",X"71",X"0D",X"3A",X"0B",X"60",X"FE",
		X"02",X"20",X"02",X"C1",X"C9",X"3E",X"01",X"32",X"25",X"60",X"3D",X"32",X"29",X"60",X"C1",X"C9",
		X"06",X"20",X"C5",X"2A",X"09",X"60",X"CD",X"CC",X"0D",X"3A",X"0B",X"60",X"FE",X"02",X"20",X"E5",
		X"C1",X"10",X"EF",X"C9",X"2A",X"09",X"60",X"2B",X"2B",X"2B",X"7E",X"FE",X"DC",X"28",X"03",X"FE",
		X"0B",X"C0",X"3A",X"2A",X"60",X"FE",X"01",X"C8",X"3E",X"01",X"21",X"1E",X"60",X"01",X"03",X"00",
		X"ED",X"B9",X"C8",X"CD",X"E3",X"F4",X"78",X"FE",X"01",X"C0",X"3E",X"01",X"32",X"28",X"60",X"32",
		X"2A",X"60",X"3D",X"32",X"2B",X"60",X"3E",X"01",X"32",X"75",X"62",X"21",X"63",X"D9",X"CD",X"84",
		X"EC",X"C9",X"3A",X"2A",X"60",X"FE",X"01",X"C0",X"11",X"E3",X"08",X"3A",X"2B",X"60",X"FE",X"05",
		X"C8",X"83",X"5F",X"7A",X"CE",X"00",X"57",X"1A",X"32",X"80",X"65",X"3A",X"2B",X"60",X"3C",X"32",
		X"2B",X"60",X"C9",X"1C",X"1C",X"1C",X"1C",X"1B",X"3A",X"2A",X"60",X"FE",X"01",X"C0",X"CD",X"E3",
		X"F4",X"78",X"FE",X"00",X"C8",X"AF",X"32",X"2A",X"60",X"32",X"28",X"60",X"32",X"29",X"60",X"32",
		X"2B",X"60",X"32",X"60",X"61",X"3E",X"19",X"32",X"80",X"65",X"3E",X"01",X"32",X"2C",X"60",X"C9",
		X"3A",X"2A",X"60",X"FE",X"01",X"C8",X"3A",X"25",X"60",X"FE",X"01",X"C8",X"3A",X"83",X"65",X"3C",
		X"DD",X"21",X"8A",X"65",X"FD",X"21",X"1C",X"60",X"11",X"04",X"00",X"CD",X"2F",X"09",X"C9",X"DD",
		X"BE",X"01",X"20",X"47",X"F5",X"06",X"08",X"3A",X"82",X"65",X"D6",X"05",X"3C",X"F5",X"DD",X"BE",
		X"00",X"28",X"2F",X"F1",X"10",X"F6",X"18",X"2D",X"FD",X"7E",X"00",X"FE",X"00",X"20",X"17",X"E5",
		X"DD",X"E5",X"21",X"00",X"01",X"CD",X"90",X"5C",X"21",X"69",X"D9",X"CD",X"84",X"EC",X"3E",X"01",
		X"32",X"75",X"62",X"DD",X"E1",X"E1",X"3E",X"01",X"FD",X"77",X"00",X"3E",X"1A",X"32",X"80",X"65",
		X"F1",X"C9",X"F1",X"18",X"D3",X"AF",X"FD",X"77",X"00",X"F1",X"C9",X"F5",X"AF",X"FD",X"77",X"00",
		X"F1",X"C9",X"DD",X"21",X"19",X"60",X"FD",X"21",X"8B",X"65",X"3E",X"C1",X"08",X"CD",X"91",X"09",
		X"C9",X"3A",X"0D",X"60",X"3D",X"DD",X"BE",X"00",X"C2",X"A0",X"09",X"08",X"FD",X"77",X"00",X"C9",
		X"3E",X"FF",X"FD",X"77",X"00",X"C9",X"DD",X"21",X"16",X"60",X"FD",X"21",X"3C",X"0A",X"21",X"8A",
		X"65",X"CD",X"B5",X"09",X"C9",X"DD",X"7E",X"00",X"FE",X"00",X"C2",X"FD",X"09",X"7E",X"3D",X"77",
		X"F5",X"DD",X"7E",X"06",X"FE",X"00",X"28",X"13",X"3A",X"82",X"65",X"3D",X"32",X"82",X"65",X"3A",
		X"95",X"62",X"FE",X"00",X"20",X"05",X"3E",X"1A",X"32",X"80",X"65",X"F1",X"FD",X"BE",X"02",X"CA",
		X"E8",X"09",X"FE",X"00",X"CA",X"F5",X"09",X"C9",X"DD",X"7E",X"03",X"FD",X"BE",X"03",X"C0",X"3E",
		X"01",X"DD",X"77",X"00",X"C9",X"DD",X"7E",X"03",X"3D",X"DD",X"77",X"03",X"C9",X"7E",X"3C",X"77",
		X"F5",X"DD",X"7E",X"06",X"FE",X"00",X"28",X"13",X"3A",X"82",X"65",X"3C",X"32",X"82",X"65",X"3A",
		X"95",X"62",X"FE",X"00",X"20",X"05",X"3E",X"1A",X"32",X"80",X"65",X"F1",X"FD",X"BE",X"00",X"CA",
		X"27",X"0A",X"FE",X"FF",X"28",X"0E",X"C9",X"DD",X"7E",X"03",X"FD",X"BE",X"01",X"C0",X"3E",X"00",
		X"DD",X"77",X"00",X"C9",X"DD",X"7E",X"03",X"3C",X"DD",X"77",X"03",X"C9",X"B0",X"03",X"20",X"02",
		X"3A",X"12",X"60",X"FE",X"00",X"C8",X"3A",X"11",X"60",X"3C",X"32",X"11",X"60",X"FE",X"5F",X"C0",
		X"AF",X"32",X"11",X"60",X"32",X"12",X"60",X"3C",X"32",X"15",X"60",X"FD",X"21",X"72",X"0A",X"06",
		X"09",X"DD",X"7E",X"02",X"FD",X"BE",X"00",X"28",X"12",X"FD",X"23",X"10",X"F4",X"AF",X"77",X"2B",
		X"77",X"C9",X"C4",X"C5",X"C6",X"C7",X"C8",X"C9",X"CA",X"CB",X"CC",X"3A",X"87",X"65",X"D6",X"00",
		X"DD",X"BE",X"03",X"28",X"0E",X"D6",X"01",X"DD",X"BE",X"03",X"28",X"07",X"C6",X"02",X"DD",X"BE",
		X"03",X"20",X"DA",X"3A",X"98",X"60",X"FE",X"04",X"20",X"D3",X"3A",X"4E",X"60",X"FE",X"00",X"28",
		X"0A",X"7D",X"FE",X"14",X"20",X"05",X"3E",X"01",X"32",X"25",X"60",X"3E",X"01",X"77",X"2B",X"77",
		X"C9",X"3A",X"98",X"60",X"FE",X"04",X"20",X"0E",X"FD",X"21",X"C9",X"0A",X"06",X"12",X"7E",X"F5",
		X"CD",X"61",X"0A",X"F1",X"77",X"C9",X"AF",X"77",X"C9",X"B8",X"B9",X"BA",X"BB",X"BC",X"BD",X"BE",
		X"BF",X"C0",X"C1",X"C2",X"C3",X"C4",X"C5",X"C6",X"C7",X"C8",X"C9",X"3A",X"12",X"60",X"FE",X"00",
		X"C0",X"21",X"87",X"65",X"3A",X"10",X"60",X"FE",X"01",X"20",X"59",X"7E",X"FE",X"1A",X"38",X"4A",
		X"3A",X"15",X"60",X"FE",X"01",X"CA",X"03",X"0B",X"7E",X"FE",X"72",X"CA",X"7C",X"0B",X"FE",X"C2",
		X"CA",X"7C",X"0B",X"35",X"AF",X"32",X"15",X"60",X"FD",X"7E",X"00",X"FE",X"01",X"20",X"0F",X"DD",
		X"7E",X"03",X"3D",X"DD",X"77",X"03",X"3A",X"C7",X"61",X"FE",X"01",X"CC",X"9E",X"EB",X"FD",X"7E",
		X"27",X"FE",X"01",X"20",X"07",X"DD",X"7E",X"17",X"3D",X"DD",X"77",X"17",X"FD",X"7E",X"67",X"FE",
		X"01",X"C0",X"DD",X"7E",X"1B",X"3D",X"DD",X"77",X"1B",X"C9",X"3E",X"00",X"32",X"10",X"60",X"3C",
		X"32",X"12",X"60",X"C9",X"7E",X"FE",X"E1",X"30",X"2E",X"34",X"FD",X"7E",X"00",X"FE",X"01",X"20",
		X"0A",X"DD",X"7E",X"03",X"3C",X"DD",X"77",X"03",X"CD",X"9E",X"EB",X"FD",X"7E",X"27",X"FE",X"01",
		X"20",X"07",X"DD",X"7E",X"17",X"3C",X"DD",X"77",X"17",X"FD",X"7E",X"67",X"FE",X"01",X"C0",X"DD",
		X"7E",X"1B",X"3C",X"DD",X"77",X"1B",X"C9",X"3E",X"01",X"32",X"10",X"60",X"3E",X"01",X"32",X"12",
		X"60",X"C9",X"FE",X"01",X"28",X"32",X"7E",X"FE",X"00",X"28",X"2D",X"79",X"FE",X"00",X"C0",X"DD",
		X"7E",X"00",X"E6",X"80",X"B0",X"DD",X"77",X"00",X"DD",X"34",X"03",X"FD",X"34",X"00",X"3A",X"F5",
		X"61",X"FE",X"00",X"C0",X"3E",X"0D",X"47",X"3A",X"98",X"60",X"B8",X"C0",X"3E",X"01",X"32",X"F5",
		X"61",X"21",X"AB",X"D9",X"CD",X"84",X"EC",X"C9",X"AF",X"FD",X"77",X"00",X"C9",X"F1",X"AF",X"32",
		X"9B",X"60",X"FD",X"77",X"00",X"C9",X"3A",X"25",X"60",X"FE",X"01",X"C8",X"3A",X"28",X"60",X"FE",
		X"01",X"CA",X"BE",X"0B",X"3A",X"D3",X"62",X"FE",X"00",X"28",X"06",X"3D",X"32",X"D3",X"62",X"18",
		X"09",X"3A",X"26",X"60",X"E6",X"10",X"FE",X"10",X"20",X"12",X"2A",X"09",X"60",X"CD",X"1C",X"D1",
		X"28",X"0A",X"CD",X"71",X"0D",X"3A",X"0B",X"60",X"FE",X"02",X"28",X"1C",X"3A",X"26",X"60",X"E6",
		X"08",X"FE",X"08",X"C2",X"BE",X"0B",X"2A",X"09",X"60",X"CD",X"CC",X"0D",X"3A",X"0B",X"60",X"FE",
		X"02",X"C2",X"BE",X"0B",X"06",X"80",X"28",X"02",X"06",X"00",X"3A",X"C1",X"62",X"FE",X"16",X"30",
		X"05",X"3C",X"3C",X"32",X"C1",X"62",X"3A",X"06",X"60",X"FE",X"0B",X"20",X"1A",X"3E",X"01",X"32",
		X"06",X"60",X"C5",X"CD",X"C2",X"10",X"E5",X"DD",X"E5",X"D5",X"21",X"10",X"00",X"CD",X"90",X"5C",
		X"D1",X"DD",X"E1",X"E1",X"C1",X"18",X"14",X"3C",X"F5",X"3A",X"58",X"61",X"FE",X"00",X"28",X"07",
		X"CD",X"50",X"0D",X"FE",X"00",X"28",X"39",X"F1",X"32",X"06",X"60",X"3A",X"06",X"60",X"21",X"80",
		X"65",X"FE",X"02",X"CC",X"AD",X"0C",X"FE",X"05",X"CC",X"AD",X"0C",X"FE",X"09",X"CC",X"AD",X"0C",
		X"FE",X"FF",X"C8",X"FE",X"04",X"CC",X"AD",X"0C",X"FE",X"06",X"CC",X"AD",X"0C",X"FE",X"08",X"CC",
		X"AD",X"0C",X"FE",X"0A",X"CC",X"AD",X"0C",X"FE",X"01",X"20",X"07",X"3E",X"20",X"B0",X"77",X"C9",
		X"F1",X"C9",X"FE",X"03",X"20",X"05",X"3E",X"1F",X"B0",X"77",X"C9",X"FE",X"07",X"20",X"05",X"3E",
		X"1E",X"B0",X"77",X"C9",X"FE",X"FF",X"20",X"04",X"3E",X"80",X"77",X"C9",X"C9",X"F5",X"78",X"FE",
		X"80",X"28",X"5A",X"2A",X"09",X"60",X"CD",X"71",X"0D",X"3A",X"0B",X"60",X"FE",X"02",X"C2",X"BD",
		X"0B",X"3A",X"82",X"65",X"3C",X"32",X"82",X"65",X"3A",X"F3",X"61",X"FE",X"00",X"20",X"1A",X"CD",
		X"F3",X"0C",X"3A",X"F3",X"61",X"FE",X"00",X"20",X"10",X"CD",X"00",X"0D",X"3A",X"F3",X"61",X"FE",
		X"00",X"20",X"06",X"21",X"99",X"D9",X"CD",X"84",X"EC",X"3E",X"01",X"FD",X"77",X"00",X"32",X"9B",
		X"60",X"F1",X"C9",X"3A",X"CF",X"61",X"FE",X"00",X"C8",X"21",X"93",X"D9",X"CD",X"84",X"EC",X"C9",
		X"3A",X"C7",X"61",X"FE",X"00",X"C9",X"21",X"A5",X"D9",X"CD",X"84",X"EC",X"C9",X"2A",X"09",X"60",
		X"CD",X"CC",X"0D",X"3A",X"0B",X"60",X"FE",X"02",X"C2",X"BD",X"0B",X"3A",X"82",X"65",X"3D",X"32",
		X"82",X"65",X"CD",X"55",X"EA",X"3A",X"F3",X"61",X"FE",X"00",X"20",X"1A",X"CD",X"F3",X"0C",X"3A",
		X"F3",X"61",X"FE",X"00",X"20",X"10",X"CD",X"00",X"0D",X"3A",X"F3",X"61",X"FE",X"00",X"20",X"06",
		X"21",X"99",X"D9",X"CD",X"84",X"EC",X"3E",X"01",X"FD",X"77",X"00",X"32",X"9B",X"60",X"F1",X"C9",
		X"C5",X"06",X"02",X"3A",X"7C",X"62",X"FE",X"00",X"28",X"02",X"06",X"01",X"3A",X"5F",X"61",X"B8",
		X"C1",X"38",X"07",X"AF",X"32",X"5F",X"61",X"3E",X"00",X"C9",X"3C",X"32",X"5F",X"61",X"3E",X"01",
		X"C9",X"3A",X"ED",X"61",X"FE",X"01",X"20",X"06",X"3E",X"02",X"32",X"0B",X"60",X"C9",X"3A",X"F2",
		X"61",X"FE",X"01",X"28",X"F3",X"CD",X"C0",X"C0",X"3A",X"0B",X"60",X"FE",X"02",X"C8",X"7D",X"D6",
		X"21",X"6F",X"7C",X"DE",X"00",X"67",X"7E",X"CD",X"05",X"0E",X"3A",X"0B",X"60",X"FE",X"02",X"C0",
		X"2B",X"7E",X"CD",X"05",X"0E",X"23",X"23",X"CD",X"AB",X"0D",X"C9",X"7E",X"FE",X"FB",X"28",X"05",
		X"FE",X"FA",X"28",X"01",X"C9",X"DD",X"E5",X"CD",X"6D",X"C1",X"DD",X"E1",X"78",X"FE",X"05",X"D8",
		X"3E",X"01",X"32",X"0B",X"60",X"C9",X"3E",X"01",X"32",X"0B",X"60",X"C9",X"3A",X"ED",X"61",X"FE",
		X"01",X"20",X"06",X"3E",X"02",X"32",X"0B",X"60",X"C9",X"CD",X"A4",X"C0",X"3A",X"0B",X"60",X"FE",
		X"02",X"C8",X"7D",X"C6",X"1F",X"6F",X"7C",X"CE",X"00",X"67",X"7E",X"CD",X"05",X"0E",X"3A",X"0B",
		X"60",X"FE",X"02",X"C0",X"2B",X"7E",X"CD",X"05",X"0E",X"23",X"23",X"CD",X"AB",X"0D",X"C9",X"3E",
		X"02",X"32",X"0B",X"60",X"C9",X"4F",X"11",X"A7",X"1B",X"06",X"23",X"1A",X"B9",X"28",X"F0",X"13",
		X"10",X"F9",X"18",X"B2",X"3A",X"9B",X"60",X"FE",X"01",X"C8",X"3A",X"26",X"60",X"E6",X"20",X"FE",
		X"20",X"28",X"13",X"3A",X"26",X"60",X"E6",X"40",X"FE",X"40",X"C0",X"2A",X"09",X"60",X"7E",X"FE",
		X"FF",X"C0",X"06",X"00",X"18",X"0A",X"2A",X"09",X"60",X"2B",X"7E",X"FE",X"FF",X"C0",X"06",X"80",
		X"3A",X"07",X"60",X"FE",X"0B",X"20",X"07",X"3E",X"01",X"32",X"07",X"60",X"18",X"15",X"3C",X"F5",
		X"3A",X"58",X"61",X"FE",X"00",X"28",X"08",X"CD",X"50",X"0D",X"FE",X"00",X"CA",X"90",X"0C",X"F1",
		X"32",X"07",X"60",X"3A",X"07",X"60",X"FE",X"01",X"C8",X"FE",X"03",X"CC",X"DF",X"0E",X"FE",X"05",
		X"C8",X"FE",X"08",X"CC",X"DF",X"0E",X"FE",X"0A",X"C8",X"FE",X"02",X"CC",X"DF",X"0E",X"FE",X"04",
		X"CC",X"DF",X"0E",X"FE",X"07",X"CC",X"DF",X"0E",X"FE",X"09",X"CC",X"DF",X"0E",X"FE",X"06",X"20",
		X"0C",X"3E",X"12",X"32",X"80",X"65",X"CD",X"DF",X"0E",X"CD",X"AD",X"0E",X"C9",X"FE",X"0B",X"20",
		X"0B",X"3E",X"92",X"32",X"80",X"65",X"CD",X"DF",X"0E",X"CD",X"AD",X"0E",X"C9",X"3A",X"F3",X"61",
		X"FE",X"00",X"20",X"06",X"21",X"8D",X"D9",X"CD",X"84",X"EC",X"3A",X"58",X"61",X"FE",X"00",X"C8",
		X"3A",X"41",X"63",X"FE",X"01",X"28",X"0C",X"3E",X"3F",X"32",X"9C",X"65",X"3A",X"82",X"65",X"32",
		X"9E",X"65",X"C9",X"3E",X"31",X"32",X"9C",X"65",X"3A",X"82",X"65",X"32",X"9E",X"65",X"C9",X"F5",
		X"AF",X"32",X"1C",X"60",X"32",X"1D",X"60",X"32",X"1E",X"60",X"78",X"FE",X"80",X"20",X"13",X"3A",
		X"83",X"65",X"3D",X"32",X"83",X"65",X"DD",X"21",X"80",X"65",X"CD",X"C9",X"0F",X"CD",X"AD",X"0E",
		X"F1",X"C9",X"3A",X"83",X"65",X"3C",X"32",X"83",X"65",X"DD",X"21",X"80",X"65",X"CD",X"C9",X"0F",
		X"CD",X"AD",X"0E",X"F1",X"C9",X"3A",X"0F",X"91",X"FE",X"1E",X"28",X"06",X"3A",X"2F",X"91",X"FE",
		X"1E",X"C0",X"3A",X"00",X"60",X"FE",X"00",X"C8",X"3A",X"54",X"60",X"FE",X"01",X"C8",X"3A",X"26",
		X"60",X"E6",X"04",X"FE",X"04",X"28",X"1D",X"3A",X"00",X"60",X"FE",X"02",X"D8",X"3A",X"51",X"60",
		X"E6",X"04",X"FE",X"04",X"C0",X"3A",X"00",X"60",X"3D",X"27",X"32",X"00",X"60",X"3E",X"02",X"32",
		X"7D",X"61",X"18",X"05",X"3E",X"01",X"32",X"7D",X"61",X"AF",X"32",X"7C",X"61",X"3A",X"00",X"60",
		X"3D",X"27",X"32",X"00",X"60",X"3E",X"0A",X"32",X"7D",X"62",X"32",X"90",X"62",X"CD",X"17",X"D0",
		X"3E",X"01",X"32",X"10",X"62",X"CD",X"51",X"F9",X"CD",X"14",X"C3",X"3E",X"01",X"32",X"9A",X"60",
		X"AF",X"32",X"53",X"60",X"32",X"55",X"60",X"3C",X"32",X"54",X"60",X"AF",X"21",X"76",X"61",X"06",
		X"06",X"77",X"23",X"10",X"FC",X"3A",X"63",X"61",X"E6",X"03",X"C6",X"01",X"32",X"56",X"60",X"3C",
		X"32",X"7E",X"61",X"21",X"C3",X"91",X"22",X"C4",X"61",X"22",X"FA",X"61",X"3E",X"01",X"32",X"C6",
		X"61",X"32",X"FC",X"61",X"CD",X"C9",X"D7",X"CD",X"DB",X"CF",X"CD",X"E7",X"CF",X"AF",X"32",X"53",
		X"63",X"CD",X"F7",X"D0",X"AF",X"32",X"48",X"63",X"C9",X"DD",X"7E",X"02",X"D6",X"01",X"E6",X"F8",
		X"C6",X"04",X"DD",X"77",X"02",X"C9",X"E1",X"3A",X"51",X"61",X"FE",X"01",X"28",X"04",X"AF",X"32",
		X"48",X"63",X"3E",X"38",X"32",X"4D",X"63",X"C9",X"3A",X"4D",X"63",X"FE",X"38",X"28",X"05",X"2A",
		X"4E",X"63",X"18",X"03",X"2A",X"40",X"61",X"11",X"03",X"00",X"E5",X"19",X"7E",X"FE",X"FF",X"28",
		X"D5",X"7E",X"E1",X"47",X"3A",X"42",X"61",X"B8",X"C0",X"AF",X"32",X"42",X"61",X"11",X"B5",X"23",
		X"3A",X"48",X"63",X"FE",X"00",X"28",X"14",X"11",X"BF",X"23",X"3A",X"48",X"63",X"FE",X"01",X"28",
		X"0A",X"11",X"C9",X"23",X"FE",X"02",X"28",X"03",X"11",X"D3",X"23",X"CD",X"58",X"10",X"3E",X"0F",
		X"D3",X"08",X"3E",X"01",X"32",X"07",X"A0",X"2A",X"40",X"61",X"11",X"03",X"00",X"19",X"7E",X"FE",
		X"FF",X"28",X"0A",X"2A",X"40",X"61",X"11",X"04",X"00",X"19",X"22",X"40",X"61",X"2A",X"4E",X"63",
		X"11",X"04",X"00",X"19",X"22",X"4E",X"63",X"C9",X"7E",X"FE",X"FE",X"C8",X"AF",X"32",X"07",X"A0",
		X"3E",X"07",X"D3",X"08",X"C5",X"06",X"38",X"3A",X"48",X"63",X"FE",X"02",X"38",X"08",X"06",X"01",
		X"FE",X"02",X"28",X"02",X"06",X"07",X"78",X"C1",X"D3",X"09",X"0E",X"00",X"D5",X"CD",X"88",X"10",
		X"D1",X"EB",X"0E",X"08",X"CD",X"B5",X"10",X"C9",X"06",X"03",X"79",X"D3",X"08",X"7E",X"CD",X"9F",
		X"10",X"23",X"0C",X"10",X"F5",X"3E",X"06",X"D3",X"08",X"3A",X"4C",X"63",X"D3",X"09",X"C9",X"E5",
		X"87",X"26",X"00",X"6F",X"11",X"F5",X"D8",X"19",X"7E",X"D3",X"09",X"0C",X"79",X"D3",X"08",X"23",
		X"7E",X"D3",X"09",X"E1",X"C9",X"06",X"06",X"79",X"D3",X"08",X"0C",X"7E",X"D3",X"09",X"23",X"10",
		X"F6",X"C9",X"3A",X"43",X"61",X"C9",X"3A",X"58",X"61",X"FE",X"00",X"C8",X"3A",X"41",X"63",X"FE",
		X"01",X"20",X"04",X"CD",X"37",X"EC",X"C9",X"3A",X"83",X"65",X"D6",X"02",X"32",X"9F",X"65",X"3A",
		X"80",X"65",X"E6",X"7F",X"FE",X"12",X"C8",X"3A",X"80",X"65",X"E6",X"80",X"FE",X"80",X"20",X"0E",
		X"3A",X"82",X"65",X"C6",X"08",X"32",X"9E",X"65",X"3E",X"BF",X"32",X"9C",X"65",X"C9",X"3A",X"82",
		X"65",X"D6",X"08",X"32",X"9E",X"65",X"3E",X"3F",X"32",X"9C",X"65",X"C9",X"3A",X"CF",X"61",X"FE",
		X"00",X"C8",X"3A",X"80",X"65",X"E6",X"7F",X"FE",X"1F",X"06",X"37",X"28",X"0D",X"3A",X"80",X"65",
		X"E6",X"7F",X"FE",X"12",X"06",X"37",X"28",X"02",X"06",X"38",X"3A",X"83",X"65",X"32",X"9F",X"65",
		X"3A",X"80",X"65",X"E6",X"7F",X"FE",X"12",X"28",X"16",X"3A",X"80",X"65",X"E6",X"80",X"FE",X"80",
		X"28",X"0D",X"3A",X"82",X"65",X"C6",X"0C",X"32",X"9E",X"65",X"78",X"32",X"9C",X"65",X"C9",X"3A",
		X"82",X"65",X"D6",X"0C",X"32",X"9E",X"65",X"78",X"F6",X"80",X"32",X"9C",X"65",X"C9",X"3A",X"54",
		X"60",X"FE",X"01",X"28",X"0A",X"3A",X"50",X"60",X"E6",X"80",X"FE",X"80",X"28",X"12",X"C9",X"3A",
		X"26",X"60",X"E6",X"80",X"FE",X"80",X"20",X"0E",X"3A",X"50",X"60",X"E6",X"80",X"FE",X"80",X"C8",
		X"3E",X"01",X"32",X"60",X"61",X"C9",X"3E",X"00",X"32",X"60",X"61",X"C9",X"3E",X"FF",X"FD",X"77",
		X"03",X"C9",X"3A",X"10",X"62",X"FE",X"01",X"C0",X"3A",X"ED",X"61",X"FE",X"01",X"C8",X"3A",X"C0",
		X"61",X"FE",X"01",X"28",X"15",X"21",X"BD",X"61",X"11",X"00",X"A8",X"01",X"06",X"00",X"ED",X"B0",
		X"AF",X"32",X"03",X"A8",X"3E",X"01",X"32",X"C0",X"61",X"C9",X"3E",X"01",X"32",X"03",X"A8",X"C9",
		X"3A",X"99",X"60",X"32",X"98",X"60",X"2A",X"38",X"60",X"22",X"44",X"60",X"FD",X"21",X"57",X"60",
		X"FD",X"22",X"93",X"60",X"DD",X"2A",X"B7",X"05",X"21",X"34",X"60",X"FD",X"21",X"27",X"60",X"CD",
		X"7E",X"06",X"3A",X"00",X"B8",X"3A",X"98",X"60",X"32",X"99",X"60",X"C9",X"3A",X"9A",X"60",X"32",
		X"98",X"60",X"2A",X"78",X"60",X"22",X"44",X"60",X"FD",X"21",X"97",X"60",X"FD",X"22",X"93",X"60",
		X"DD",X"2A",X"B9",X"05",X"21",X"74",X"60",X"FD",X"21",X"67",X"60",X"CD",X"7E",X"06",X"3A",X"00",
		X"B8",X"3A",X"98",X"60",X"32",X"9A",X"60",X"C9",X"F3",X"3E",X"00",X"32",X"03",X"A0",X"CD",X"B7",
		X"C3",X"3E",X"3F",X"CD",X"A3",X"C3",X"CD",X"A4",X"F8",X"3E",X"01",X"32",X"0D",X"60",X"32",X"03",
		X"A0",X"32",X"98",X"60",X"32",X"99",X"60",X"32",X"9A",X"60",X"AF",X"32",X"08",X"60",X"32",X"37",
		X"60",X"32",X"4E",X"60",X"32",X"77",X"60",X"32",X"87",X"65",X"32",X"9A",X"65",X"32",X"9B",X"65",
		X"32",X"59",X"61",X"32",X"CF",X"61",X"32",X"E0",X"61",X"32",X"E1",X"61",X"3E",X"01",X"32",X"ED",
		X"61",X"CD",X"EE",X"C5",X"21",X"1D",X"90",X"11",X"20",X"00",X"3E",X"F0",X"06",X"20",X"77",X"E5",
		X"F5",X"7C",X"C6",X"08",X"67",X"3E",X"04",X"77",X"F1",X"E1",X"19",X"10",X"F1",X"21",X"00",X"00",
		X"22",X"F6",X"61",X"CD",X"42",X"15",X"3E",X"01",X"32",X"54",X"60",X"11",X"80",X"65",X"21",X"59",
		X"15",X"01",X"04",X"00",X"ED",X"B0",X"11",X"94",X"65",X"21",X"61",X"15",X"01",X"04",X"00",X"ED",
		X"B0",X"3A",X"74",X"62",X"FE",X"01",X"C8",X"11",X"00",X"4C",X"21",X"A5",X"91",X"3E",X"16",X"08",
		X"CD",X"F0",X"55",X"11",X"0B",X"4C",X"21",X"A6",X"91",X"3E",X"16",X"08",X"CD",X"F0",X"55",X"11",
		X"16",X"4C",X"21",X"A7",X"91",X"3E",X"16",X"08",X"CD",X"F0",X"55",X"11",X"21",X"4C",X"21",X"AA",
		X"91",X"3E",X"13",X"08",X"CD",X"F0",X"55",X"3A",X"00",X"B0",X"E6",X"20",X"FE",X"20",X"20",X"0A",
		X"3E",X"E1",X"32",X"CA",X"90",X"3E",X"13",X"32",X"CA",X"98",X"21",X"6B",X"93",X"0E",X"1A",X"CD",
		X"DD",X"23",X"FB",X"ED",X"56",X"FF",X"06",X"02",X"11",X"00",X"40",X"CD",X"42",X"15",X"1B",X"7A",
		X"FE",X"00",X"20",X"F7",X"3A",X"00",X"B0",X"E6",X"40",X"FE",X"40",X"20",X"11",X"E5",X"21",X"00",
		X"38",X"22",X"40",X"61",X"AF",X"32",X"42",X"61",X"3E",X"01",X"32",X"4A",X"63",X"E1",X"10",X"D8",
		X"06",X"05",X"DD",X"21",X"5B",X"92",X"DD",X"36",X"00",X"18",X"DD",X"36",X"01",X"17",X"DD",X"36",
		X"20",X"19",X"DD",X"36",X"21",X"16",X"DD",X"36",X"40",X"1A",X"DD",X"36",X"41",X"15",X"11",X"00",
		X"06",X"CD",X"42",X"15",X"1B",X"7A",X"FE",X"00",X"20",X"F7",X"DD",X"36",X"00",X"B7",X"DD",X"36",
		X"01",X"1C",X"DD",X"36",X"20",X"B6",X"DD",X"36",X"21",X"1B",X"DD",X"36",X"40",X"B2",X"DD",X"36",
		X"41",X"B5",X"11",X"00",X"06",X"CD",X"42",X"15",X"1B",X"7A",X"FE",X"00",X"20",X"F7",X"10",X"B2",
		X"11",X"00",X"40",X"CD",X"42",X"15",X"1B",X"7A",X"FE",X"00",X"20",X"F7",X"DD",X"21",X"6E",X"92",
		X"DD",X"36",X"00",X"16",X"DD",X"36",X"01",X"21",X"DD",X"36",X"1F",X"0E",X"DD",X"36",X"20",X"15",
		X"DD",X"36",X"21",X"20",X"DD",X"36",X"40",X"14",X"DD",X"36",X"41",X"1F",X"DD",X"36",X"61",X"1E",
		X"11",X"00",X"14",X"CD",X"42",X"15",X"1B",X"7A",X"FE",X"00",X"20",X"F7",X"DD",X"21",X"6E",X"92",
		X"DD",X"36",X"00",X"00",X"DD",X"36",X"01",X"B2",X"DD",X"36",X"1F",X"6A",X"DD",X"36",X"20",X"6B",
		X"DD",X"36",X"21",X"AD",X"DD",X"36",X"40",X"6C",X"DD",X"36",X"41",X"9B",X"DD",X"36",X"61",X"72",
		X"11",X"00",X"40",X"CD",X"42",X"15",X"1B",X"7A",X"FE",X"00",X"20",X"F7",X"DD",X"21",X"6E",X"92",
		X"DD",X"36",X"00",X"16",X"DD",X"36",X"01",X"21",X"DD",X"36",X"1F",X"0E",X"DD",X"36",X"20",X"15",
		X"DD",X"36",X"21",X"20",X"DD",X"36",X"40",X"14",X"DD",X"36",X"41",X"1F",X"DD",X"36",X"61",X"1E",
		X"DD",X"21",X"4D",X"92",X"DD",X"36",X"00",X"10",X"06",X"08",X"DD",X"21",X"91",X"91",X"DD",X"36",
		X"40",X"B8",X"11",X"00",X"07",X"CD",X"42",X"15",X"1B",X"7A",X"FE",X"00",X"20",X"F7",X"DD",X"36",
		X"00",X"BD",X"DD",X"36",X"20",X"BA",X"11",X"00",X"07",X"CD",X"42",X"15",X"1B",X"7A",X"FE",X"00",
		X"20",X"F7",X"DD",X"36",X"40",X"43",X"11",X"00",X"07",X"CD",X"42",X"15",X"1B",X"7A",X"FE",X"00",
		X"20",X"F7",X"DD",X"36",X"00",X"45",X"DD",X"36",X"20",X"44",X"DD",X"36",X"40",X"43",X"11",X"00",
		X"07",X"CD",X"42",X"15",X"1B",X"7A",X"FE",X"00",X"20",X"F7",X"10",X"B2",X"11",X"00",X"20",X"CD",
		X"42",X"15",X"1B",X"7A",X"FE",X"00",X"20",X"F7",X"DD",X"21",X"6E",X"92",X"DD",X"36",X"00",X"00",
		X"DD",X"36",X"01",X"B2",X"DD",X"36",X"1F",X"6A",X"DD",X"36",X"20",X"6B",X"DD",X"36",X"21",X"AD",
		X"DD",X"36",X"40",X"6C",X"DD",X"36",X"41",X"9B",X"DD",X"36",X"61",X"72",X"DD",X"21",X"4D",X"92",
		X"DD",X"36",X"00",X"62",X"21",X"6B",X"93",X"0E",X"1A",X"CD",X"DD",X"23",X"3E",X"30",X"32",X"94",
		X"65",X"3E",X"0C",X"32",X"95",X"65",X"3E",X"00",X"32",X"96",X"65",X"3E",X"D8",X"32",X"97",X"65",
		X"3E",X"80",X"32",X"27",X"60",X"11",X"00",X"20",X"CD",X"42",X"15",X"1B",X"7A",X"FE",X"00",X"20",
		X"F7",X"21",X"6B",X"93",X"0E",X"19",X"F3",X"E5",X"C5",X"CD",X"DD",X"23",X"C1",X"E1",X"FB",X"ED",
		X"56",X"FF",X"11",X"00",X"08",X"CD",X"42",X"15",X"1B",X"7A",X"FE",X"00",X"20",X"F7",X"11",X"E0",
		X"FF",X"19",X"0D",X"79",X"FE",X"FF",X"20",X"DE",X"AF",X"32",X"27",X"60",X"3E",X"2C",X"32",X"94",
		X"65",X"11",X"00",X"40",X"CD",X"42",X"15",X"1B",X"7A",X"FE",X"00",X"20",X"F7",X"3E",X"00",X"32",
		X"ED",X"61",X"06",X"01",X"21",X"80",X"65",X"3E",X"00",X"32",X"54",X"60",X"3A",X"00",X"60",X"FE",
		X"00",X"C0",X"3E",X"00",X"CD",X"A8",X"C3",X"3E",X"01",X"32",X"32",X"63",X"3E",X"00",X"32",X"03",
		X"A0",X"CD",X"B7",X"C3",X"3E",X"04",X"CD",X"A3",X"C3",X"DD",X"21",X"A1",X"1F",X"3A",X"00",X"B0",
		X"E6",X"20",X"FE",X"20",X"20",X"04",X"DD",X"21",X"A5",X"1D",X"CD",X"2A",X"D8",X"AF",X"32",X"32",
		X"63",X"C9",X"3A",X"00",X"60",X"FE",X"00",X"C8",X"3A",X"74",X"62",X"FE",X"01",X"C8",X"3E",X"00",
		X"32",X"ED",X"61",X"3A",X"00",X"B8",X"E1",X"18",X"A4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"CD",X"72",X"15",X"CD",X"8F",X"15",X"CD",X"AC",X"15",X"CD",X"C9",
		X"15",X"C9",X"3A",X"26",X"60",X"E6",X"01",X"47",X"3A",X"50",X"60",X"E6",X"01",X"B8",X"C8",X"3A",
		X"50",X"60",X"E6",X"01",X"FE",X"01",X"C0",X"3E",X"01",X"0E",X"01",X"CD",X"E6",X"15",X"C9",X"3A",
		X"26",X"60",X"E6",X"02",X"47",X"3A",X"50",X"60",X"E6",X"02",X"B8",X"C8",X"3A",X"50",X"60",X"E6",
		X"02",X"FE",X"02",X"C0",X"3E",X"02",X"0E",X"02",X"CD",X"E6",X"15",X"C9",X"3A",X"51",X"60",X"E6",
		X"01",X"47",X"3A",X"52",X"60",X"E6",X"01",X"B8",X"C8",X"3A",X"52",X"60",X"E6",X"01",X"FE",X"01",
		X"C0",X"3E",X"06",X"0E",X"05",X"CD",X"E6",X"15",X"C9",X"3A",X"51",X"60",X"E6",X"02",X"47",X"3A",
		X"52",X"60",X"E6",X"02",X"B8",X"C8",X"3A",X"52",X"60",X"E6",X"02",X"FE",X"02",X"C0",X"3E",X"0E",
		X"0E",X"0A",X"CD",X"E6",X"15",X"C9",X"F5",X"CD",X"82",X"16",X"F1",X"47",X"3A",X"63",X"61",X"E6",
		X"04",X"FE",X"04",X"78",X"28",X"01",X"87",X"21",X"E4",X"61",X"86",X"77",X"FE",X"02",X"D4",X"02",
		X"16",X"C9",X"21",X"E4",X"61",X"7E",X"FE",X"02",X"D8",X"3A",X"00",X"60",X"FE",X"90",X"C8",X"C6",
		X"01",X"27",X"32",X"00",X"60",X"21",X"E4",X"61",X"35",X"35",X"CD",X"D9",X"D4",X"20",X"0A",X"21",
		X"68",X"5B",X"22",X"40",X"61",X"AF",X"32",X"42",X"61",X"CD",X"2E",X"16",X"18",X"D4",X"3A",X"00",
		X"60",X"E6",X"0F",X"32",X"9F",X"90",X"3A",X"00",X"60",X"CB",X"0F",X"CB",X"0F",X"CB",X"0F",X"CB",
		X"0F",X"E6",X"0F",X"32",X"BF",X"90",X"3E",X"E0",X"06",X"06",X"21",X"BF",X"93",X"CD",X"73",X"C3",
		X"3A",X"56",X"60",X"FE",X"00",X"28",X"09",X"21",X"BF",X"93",X"47",X"3E",X"CA",X"CD",X"73",X"C3",
		X"3A",X"10",X"62",X"FE",X"01",X"C0",X"3E",X"11",X"32",X"DF",X"92",X"3E",X"13",X"32",X"BF",X"92",
		X"3E",X"24",X"32",X"9F",X"92",X"3A",X"D3",X"60",X"32",X"5F",X"92",X"C9",X"01",X"01",X"01",X"00",
		X"01",X"00",X"79",X"21",X"E5",X"61",X"86",X"77",X"C9",X"3A",X"26",X"60",X"32",X"50",X"60",X"AF",
		X"32",X"07",X"A0",X"CD",X"D9",X"16",X"47",X"CD",X"D9",X"16",X"B8",X"28",X"05",X"32",X"60",X"63",
		X"18",X"F1",X"2F",X"CD",X"F0",X"16",X"CD",X"05",X"17",X"32",X"26",X"60",X"3A",X"51",X"60",X"32",
		X"52",X"60",X"CD",X"E9",X"16",X"47",X"CD",X"E9",X"16",X"B8",X"28",X"05",X"32",X"60",X"63",X"18",
		X"F1",X"2F",X"CD",X"F0",X"16",X"32",X"51",X"60",X"3A",X"00",X"B0",X"2F",X"32",X"63",X"61",X"3E",
		X"01",X"32",X"07",X"A0",X"3E",X"63",X"D3",X"56",X"C9",X"3E",X"07",X"D3",X"08",X"3A",X"4D",X"63",
		X"D3",X"09",X"3E",X"0E",X"D3",X"08",X"DB",X"0C",X"C9",X"3E",X"0F",X"D3",X"08",X"DB",X"0C",X"C9",
		X"F5",X"3A",X"ED",X"61",X"FE",X"01",X"28",X"09",X"3A",X"F2",X"61",X"FE",X"01",X"28",X"02",X"F1",
		X"C9",X"F1",X"E6",X"03",X"C9",X"47",X"3A",X"00",X"B0",X"2F",X"CB",X"07",X"E6",X"01",X"4F",X"3A",
		X"7C",X"61",X"A1",X"32",X"FD",X"61",X"FE",X"01",X"28",X"02",X"78",X"C9",X"3A",X"51",X"60",X"E6",
		X"F8",X"4F",X"78",X"E6",X"07",X"B1",X"C9",X"3A",X"54",X"60",X"FE",X"00",X"C8",X"CD",X"00",X"55",
		X"C9",X"3A",X"54",X"60",X"FE",X"01",X"C8",X"3A",X"26",X"60",X"E6",X"03",X"32",X"26",X"60",X"DD",
		X"21",X"20",X"18",X"3A",X"41",X"63",X"FE",X"01",X"28",X"04",X"DD",X"21",X"48",X"18",X"FD",X"21",
		X"80",X"65",X"11",X"04",X"00",X"3A",X"88",X"62",X"FE",X"00",X"CC",X"F1",X"17",X"3A",X"88",X"62",
		X"FE",X"00",X"28",X"05",X"DD",X"19",X"3D",X"18",X"F7",X"3A",X"5D",X"63",X"FE",X"01",X"28",X"53",
		X"DD",X"7E",X"03",X"FE",X"FF",X"28",X"52",X"FE",X"FE",X"CA",X"E3",X"17",X"E6",X"80",X"FE",X"80",
		X"CC",X"BD",X"17",X"DD",X"7E",X"03",X"47",X"3A",X"26",X"60",X"E6",X"07",X"B0",X"32",X"26",X"60",
		X"FD",X"7E",X"02",X"DD",X"BE",X"00",X"C0",X"FD",X"7E",X"03",X"DD",X"BE",X"01",X"C0",X"3A",X"0D",
		X"60",X"DD",X"BE",X"02",X"C0",X"3A",X"88",X"62",X"3C",X"32",X"88",X"62",X"3A",X"26",X"60",X"E6",
		X"80",X"FE",X"80",X"C8",X"3A",X"26",X"60",X"E6",X"07",X"32",X"26",X"60",X"C9",X"3E",X"01",X"32",
		X"5D",X"63",X"C9",X"AF",X"32",X"5D",X"63",X"18",X"DC",X"3E",X"10",X"32",X"97",X"65",X"32",X"9B",
		X"65",X"3E",X"D0",X"32",X"96",X"65",X"3E",X"E0",X"32",X"9A",X"65",X"3A",X"87",X"65",X"FE",X"11",
		X"C0",X"18",X"C2",X"3A",X"8A",X"65",X"FE",X"60",X"C0",X"3A",X"19",X"60",X"FE",X"02",X"C0",X"18",
		X"B4",X"21",X"C3",X"91",X"22",X"C4",X"61",X"22",X"FA",X"61",X"3E",X"01",X"32",X"C6",X"61",X"32",
		X"FC",X"61",X"3E",X"05",X"32",X"99",X"60",X"32",X"9A",X"60",X"3E",X"20",X"32",X"96",X"65",X"32",
		X"9A",X"65",X"3E",X"A0",X"32",X"97",X"65",X"32",X"9B",X"65",X"3E",X"0C",X"32",X"7D",X"62",X"C9",
		X"61",X"70",X"02",X"10",X"64",X"A0",X"02",X"40",X"30",X"A0",X"02",X"08",X"2C",X"90",X"02",X"20",
		X"A4",X"90",X"01",X"08",X"A4",X"D8",X"01",X"40",X"2B",X"D8",X"01",X"08",X"2C",X"18",X"01",X"20",
		X"10",X"18",X"01",X"08",X"FF",X"FF",X"FF",X"08",X"2C",X"D8",X"01",X"10",X"2C",X"70",X"01",X"20",
		X"8B",X"68",X"02",X"10",X"8B",X"68",X"02",X"90",X"B9",X"68",X"02",X"10",X"B9",X"68",X"02",X"10",
		X"BC",X"50",X"02",X"20",X"29",X"50",X"03",X"10",X"2C",X"A0",X"03",X"40",X"60",X"A0",X"03",X"10",
		X"30",X"A0",X"03",X"08",X"2C",X"50",X"03",X"20",X"C0",X"50",X"02",X"08",X"BC",X"18",X"02",X"20",
		X"98",X"18",X"02",X"0C",X"70",X"18",X"02",X"08",X"60",X"18",X"02",X"0C",X"18",X"18",X"02",X"08",
		X"18",X"18",X"02",X"80",X"82",X"18",X"01",X"08",X"78",X"18",X"01",X"08",X"78",X"18",X"01",X"80",
		X"60",X"18",X"01",X"08",X"5A",X"18",X"01",X"08",X"59",X"18",X"01",X"80",X"56",X"18",X"01",X"08",
		X"76",X"18",X"02",X"10",X"70",X"18",X"02",X"08",X"70",X"18",X"02",X"80",X"88",X"18",X"02",X"10",
		X"8C",X"18",X"03",X"10",X"8C",X"50",X"03",X"40",X"6C",X"50",X"03",X"08",X"6C",X"50",X"03",X"80",
		X"8A",X"50",X"03",X"10",X"8C",X"50",X"03",X"10",X"8C",X"18",X"03",X"20",X"BC",X"18",X"02",X"08",
		X"BC",X"50",X"02",X"40",X"2C",X"50",X"03",X"10",X"2C",X"C0",X"03",X"40",X"60",X"C0",X"03",X"10",
		X"60",X"C0",X"03",X"80",X"60",X"C0",X"03",X"00",X"00",X"00",X"03",X"FE",X"60",X"C0",X"03",X"80",
		X"CB",X"C0",X"03",X"00",X"CC",X"C0",X"03",X"00",X"CC",X"80",X"03",X"20",X"80",X"80",X"03",X"08",
		X"C0",X"18",X"05",X"10",X"FF",X"FF",X"FF",X"10",X"7A",X"FD",X"21",X"4E",X"22",X"FE",X"34",X"D8",
		X"FD",X"21",X"5D",X"22",X"FE",X"38",X"D8",X"FD",X"21",X"E8",X"21",X"FE",X"44",X"D8",X"FD",X"21",
		X"09",X"22",X"FE",X"48",X"D8",X"FD",X"21",X"30",X"22",X"C9",X"DD",X"E5",X"FD",X"E5",X"E5",X"C5",
		X"D5",X"78",X"FE",X"01",X"20",X"06",X"FD",X"21",X"75",X"22",X"18",X"49",X"FE",X"02",X"20",X"13",
		X"47",X"3A",X"0D",X"60",X"B8",X"30",X"06",X"FD",X"21",X"93",X"22",X"18",X"38",X"FD",X"21",X"BA",
		X"22",X"18",X"32",X"FE",X"03",X"20",X"13",X"47",X"3A",X"0D",X"60",X"B8",X"30",X"06",X"FD",X"21",
		X"E1",X"22",X"18",X"21",X"FD",X"21",X"FF",X"22",X"18",X"1B",X"FE",X"04",X"20",X"13",X"47",X"3A",
		X"0D",X"60",X"B8",X"30",X"06",X"FD",X"21",X"1D",X"23",X"18",X"0A",X"FD",X"21",X"2C",X"23",X"18",
		X"04",X"FD",X"21",X"3B",X"23",X"D1",X"FD",X"7E",X"00",X"67",X"FD",X"7E",X"01",X"6F",X"AF",X"ED",
		X"52",X"28",X"10",X"FD",X"23",X"FD",X"23",X"FD",X"23",X"FD",X"7E",X"02",X"FE",X"FF",X"20",X"E6",
		X"C3",X"D1",X"19",X"FD",X"7E",X"02",X"FE",X"80",X"20",X"06",X"CD",X"A2",X"F6",X"C3",X"D1",X"19",
		X"FE",X"40",X"20",X"06",X"CD",X"C0",X"F6",X"C3",X"D1",X"19",X"DD",X"2A",X"95",X"60",X"DD",X"77",
		X"00",X"C1",X"E1",X"FD",X"E1",X"DD",X"E1",X"E1",X"C3",X"44",X"F6",X"0A",X"08",X"06",X"04",X"02",
		X"C7",X"C6",X"C5",X"C4",X"C3",X"C2",X"C1",X"C0",X"FF",X"F7",X"F5",X"F3",X"F2",X"DA",X"D9",X"D8",
		X"D7",X"D6",X"D5",X"D4",X"D3",X"D2",X"D1",X"D0",X"CF",X"CE",X"CD",X"CC",X"CB",X"CA",X"C9",X"C8",
		X"E9",X"C0",X"C1",X"C2",X"C3",X"C7",X"C6",X"C5",X"C4",X"B0",X"B1",X"B2",X"B3",X"4C",X"4D",X"4E",
		X"4F",X"E8",X"19",X"1B",X"1D",X"1F",X"21",X"23",X"25",X"28",X"41",X"35",X"04",X"5F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"0C",X"D0",X"18",X"20",X"0C",X"D0",X"18",X"26",
		X"11",X"1C",X"11",X"14",X"1F",X"1E",X"10",X"11",X"25",X"24",X"1F",X"1D",X"11",X"24",X"19",X"1F",
		X"1E",X"3F",X"8A",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"8F",X"3F",X"8C",X"90",X"90",
		X"90",X"90",X"90",X"90",X"90",X"90",X"8D",X"3F",X"13",X"15",X"10",X"1A",X"15",X"25",X"10",X"1C",
		X"15",X"10",X"12",X"11",X"17",X"1E",X"11",X"22",X"14",X"10",X"11",X"10",X"15",X"24",X"15",X"10",
		X"13",X"22",X"15",X"15",X"3F",X"20",X"11",X"22",X"10",X"26",X"11",X"1C",X"11",X"14",X"1F",X"1E",
		X"10",X"11",X"25",X"24",X"1F",X"1D",X"11",X"24",X"19",X"1F",X"1E",X"3F",X"00",X"42",X"01",X"1A",
		X"10",X"12",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"00",X"51",X"01",X"1A",
		X"1F",X"1A",X"1F",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"00",X"60",X"01",X"20",
		X"19",X"15",X"22",X"22",X"1F",X"24",X"10",X"10",X"10",X"10",X"10",X"10",X"00",X"79",X"01",X"17",
		X"11",X"23",X"24",X"1F",X"25",X"1E",X"15",X"24",X"10",X"10",X"10",X"10",X"00",X"89",X"01",X"16",
		X"11",X"1E",X"13",X"18",X"1F",X"19",X"23",X"10",X"10",X"10",X"10",X"10",X"54",X"93",X"05",X"67",
		X"93",X"01",X"B7",X"91",X"01",X"2F",X"91",X"01",X"67",X"93",X"02",X"63",X"93",X"02",X"38",X"92",
		X"02",X"78",X"91",X"02",X"8A",X"93",X"03",X"78",X"93",X"03",X"70",X"91",X"03",X"38",X"91",X"03",
		X"6A",X"93",X"04",X"0E",X"93",X"04",X"98",X"91",X"04",X"0E",X"92",X"05",X"6E",X"90",X"04",X"1C",
		X"92",X"05",X"FF",X"FF",X"FF",X"54",X"93",X"05",X"7B",X"92",X"01",X"6F",X"91",X"01",X"0F",X"91",
		X"01",X"67",X"93",X"02",X"8E",X"92",X"02",X"38",X"92",X"02",X"D8",X"92",X"02",X"8A",X"93",X"03",
		X"78",X"93",X"03",X"70",X"91",X"03",X"D8",X"91",X"03",X"8A",X"93",X"04",X"0E",X"93",X"04",X"78",
		X"90",X"04",X"E9",X"91",X"05",X"6E",X"90",X"04",X"1C",X"92",X"05",X"FF",X"FF",X"FF",X"54",X"93",
		X"05",X"94",X"92",X"01",X"6F",X"91",X"01",X"9B",X"90",X"01",X"94",X"92",X"02",X"8E",X"92",X"02",
		X"F8",X"91",X"02",X"58",X"92",X"02",X"23",X"92",X"03",X"1C",X"93",X"03",X"70",X"91",X"03",X"D8",
		X"91",X"03",X"38",X"93",X"04",X"0E",X"93",X"04",X"23",X"92",X"04",X"0E",X"93",X"05",X"6E",X"90",
		X"04",X"1C",X"92",X"05",X"FF",X"FF",X"FF",X"D9",X"D8",X"E9",X"E9",X"D7",X"D6",X"D5",X"E9",X"D2",
		X"D1",X"D4",X"D3",X"CE",X"CD",X"D0",X"CF",X"CB",X"CA",X"E9",X"CC",X"66",X"65",X"E9",X"C9",X"63",
		X"62",X"E9",X"64",X"60",X"5F",X"E9",X"61",X"E0",X"FF",X"F2",X"F3",X"F5",X"4C",X"4D",X"4E",X"4F",
		X"F7",X"4B",X"DF",X"DE",X"51",X"52",X"57",X"4A",X"49",X"C7",X"C6",X"C5",X"C4",X"C3",X"C2",X"C1",
		X"C0",X"E9",X"B3",X"B2",X"B1",X"B0",X"8F",X"8E",X"8D",X"E8",X"F1",X"F2",X"F3",X"F4",X"F5",X"F6",
		X"F7",X"30",X"A5",X"40",X"30",X"B0",X"40",X"30",X"BA",X"40",X"30",X"BE",X"40",X"31",X"05",X"80",
		X"31",X"10",X"80",X"31",X"1A",X"80",X"31",X"1D",X"80",X"35",X"47",X"80",X"35",X"4B",X"80",X"35",
		X"50",X"80",X"35",X"55",X"80",X"35",X"5E",X"80",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"2E",X"92",X"04",X"00",X"00",X"00",X"00",X"1B",X"92",X"01",X"0A",X"92",X"03",X"07",X"93",X"05",
		X"A3",X"91",X"02",X"54",X"52",X"4F",X"55",X"56",X"45",X"5A",X"3A",X"4C",X"41",X"3A",X"43",X"4C",
		X"45",X"46",X"FE",X"45",X"54",X"3A",X"44",X"45",X"4C",X"49",X"56",X"52",X"45",X"5A",X"3A",X"56",
		X"4F",X"54",X"52",X"45",X"FE",X"43",X"4F",X"4D",X"50",X"41",X"47",X"4E",X"4F",X"4E",X"3A",X"44",
		X"45",X"3A",X"43",X"45",X"4C",X"4C",X"55",X"4C",X"45",X"FE",X"3A",X"3A",X"3A",X"3A",X"3A",X"42",
		X"4F",X"4E",X"4E",X"45",X"3A",X"43",X"48",X"41",X"4E",X"43",X"45",X"3A",X"66",X"FE",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"46",X"4F",X"55",X"4E",X"44",X"3A",
		X"54",X"48",X"45",X"3A",X"4B",X"45",X"59",X"FE",X"41",X"4E",X"44",X"3A",X"52",X"45",X"4C",X"45",
		X"41",X"53",X"45",X"3A",X"59",X"4F",X"55",X"52",X"3A",X"46",X"52",X"49",X"45",X"4E",X"44",X"3A",
		X"FE",X"3A",X"3A",X"3A",X"3A",X"3A",X"47",X"4F",X"4F",X"44",X"3A",X"4C",X"55",X"43",X"4B",X"3A",
		X"66",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"42",X"52",
		X"41",X"56",X"4F",X"3A",X"FE",X"3A",X"FE",X"3A",X"FE",X"42",X"4F",X"4E",X"4E",X"45",X"3A",X"43",
		X"48",X"41",X"4E",X"43",X"45",X"3A",X"50",X"4F",X"55",X"52",X"3A",X"4C",X"45",X"FE",X"50",X"52",
		X"4F",X"43",X"48",X"41",X"49",X"4E",X"3A",X"44",X"45",X"46",X"49",X"FE",X"4D",X"41",X"49",X"53",
		X"3A",X"41",X"54",X"54",X"45",X"4E",X"54",X"49",X"4F",X"4E",X"3A",X"66",X"FE",X"47",X"45",X"4E",
		X"44",X"41",X"52",X"4D",X"45",X"53",X"3A",X"4F",X"4E",X"54",X"3A",X"52",X"45",X"43",X"55",X"FE",
		X"4F",X"52",X"44",X"52",X"45",X"3A",X"44",X"45",X"3A",X"54",X"49",X"52",X"45",X"52",X"3A",X"41",
		X"3A",X"56",X"55",X"45",X"FE",X"3A",X"FE",X"3A",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"43",X"4F",X"4E",X"47",X"52",X"41",X"54",X"55",X"4C",X"41",X"54",
		X"49",X"4F",X"4E",X"53",X"3A",X"FE",X"3A",X"FE",X"47",X"4F",X"4F",X"44",X"3A",X"4C",X"55",X"43",
		X"4B",X"3A",X"46",X"4F",X"52",X"3A",X"54",X"48",X"45",X"3A",X"4E",X"45",X"58",X"54",X"FE",X"43",
		X"48",X"41",X"4C",X"4C",X"45",X"4E",X"47",X"45",X"FE",X"42",X"55",X"54",X"3A",X"57",X"41",X"52",
		X"4E",X"49",X"4E",X"47",X"3A",X"66",X"FE",X"50",X"4F",X"4C",X"49",X"43",X"45",X"3A",X"48",X"41",
		X"56",X"45",X"3A",X"42",X"45",X"45",X"4E",X"3A",X"49",X"4E",X"53",X"54",X"52",X"55",X"43",X"54",
		X"45",X"44",X"FE",X"54",X"4F",X"3A",X"53",X"48",X"4F",X"4F",X"54",X"3A",X"4F",X"4E",X"3A",X"53",
		X"49",X"47",X"48",X"54",X"FE",X"3A",X"FE",X"3A",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"41",X"4C",X"43",X"41",X"54",X"52",X"41",X"5A",X"3A",X"50",X"52",
		X"49",X"53",X"4F",X"4E",X"3A",X"54",X"4F",X"3A",X"49",X"4E",X"54",X"45",X"52",X"50",X"4F",X"4C",
		X"FE",X"3A",X"65",X"53",X"54",X"4F",X"50",X"65",X"FE",X"5B",X"5B",X"5B",X"5B",X"5B",X"FE",X"3A",
		X"FE",X"3A",X"FE",X"42",X"41",X"47",X"4D",X"41",X"4E",X"3A",X"48",X"41",X"53",X"3A",X"45",X"53",
		X"43",X"41",X"50",X"45",X"44",X"3A",X"65",X"53",X"54",X"4F",X"50",X"65",X"FE",X"3A",X"FE",X"50",
		X"4F",X"4C",X"49",X"43",X"45",X"3A",X"41",X"52",X"45",X"3A",X"4F",X"4E",X"3A",X"48",X"49",X"53",
		X"3A",X"48",X"45",X"45",X"4C",X"53",X"FE",X"3A",X"65",X"53",X"54",X"4F",X"50",X"65",X"FE",X"48",
		X"45",X"3A",X"57",X"49",X"4C",X"4C",X"3A",X"50",X"52",X"4F",X"42",X"41",X"42",X"4C",X"59",X"3A",
		X"54",X"52",X"59",X"3A",X"54",X"4F",X"FE",X"52",X"45",X"43",X"4F",X"56",X"45",X"52",X"3A",X"54",
		X"48",X"45",X"3A",X"47",X"4F",X"4C",X"44",X"3A",X"42",X"41",X"47",X"53",X"3A",X"FE",X"3A",X"FE",
		X"57",X"48",X"45",X"4E",X"3A",X"48",X"45",X"3A",X"48",X"41",X"53",X"3A",X"54",X"48",X"45",X"4D",
		X"3A",X"41",X"4E",X"44",X"3A",X"54",X"48",X"45",X"FE",X"4B",X"45",X"59",X"3A",X"46",X"4F",X"55",
		X"4E",X"44",X"3A",X"49",X"4E",X"3A",X"54",X"48",X"45",X"3A",X"4D",X"49",X"4E",X"45",X"FE",X"48",
		X"45",X"3A",X"57",X"49",X"4C",X"4C",X"3A",X"54",X"52",X"59",X"3A",X"54",X"4F",X"3A",X"52",X"45",
		X"4C",X"45",X"41",X"53",X"45",X"FE",X"48",X"49",X"53",X"3A",X"46",X"52",X"49",X"45",X"4E",X"44",
		X"3A",X"4C",X"4F",X"43",X"4B",X"45",X"44",X"3A",X"49",X"4E",X"3A",X"54",X"48",X"45",X"FE",X"44",
		X"55",X"4E",X"47",X"45",X"4F",X"4E",X"3A",X"65",X"53",X"54",X"4F",X"50",X"65",X"FE",X"3A",X"FE",
		X"48",X"45",X"3A",X"57",X"49",X"4C",X"4C",X"3A",X"48",X"41",X"56",X"45",X"3A",X"53",X"49",X"58",
		X"3A",X"53",X"48",X"4F",X"54",X"53",X"FE",X"49",X"4E",X"3A",X"45",X"41",X"43",X"48",X"3A",X"52",
		X"45",X"56",X"4F",X"4C",X"56",X"45",X"52",X"3A",X"43",X"4F",X"4C",X"4C",X"45",X"43",X"54",X"45",
		X"44",X"FE",X"46",X"52",X"4F",X"4D",X"3A",X"54",X"48",X"45",X"3A",X"47",X"55",X"4E",X"53",X"4D",
		X"49",X"54",X"48",X"6A",X"53",X"3A",X"52",X"4F",X"4F",X"4D",X"FE",X"3A",X"FE",X"50",X"4F",X"4C",
		X"49",X"43",X"45",X"3A",X"48",X"41",X"56",X"45",X"3A",X"42",X"45",X"45",X"4E",X"3A",X"49",X"4E",
		X"53",X"54",X"52",X"55",X"43",X"54",X"45",X"44",X"FE",X"4E",X"4F",X"54",X"3A",X"54",X"4F",X"3A",
		X"53",X"48",X"4F",X"4F",X"54",X"3A",X"46",X"49",X"52",X"53",X"54",X"3A",X"65",X"53",X"54",X"4F",
		X"50",X"65",X"FE",X"3A",X"FE",X"3A",X"FE",X"3A",X"3A",X"3A",X"3A",X"47",X"4F",X"4F",X"44",X"3A",
		X"4C",X"55",X"43",X"4B",X"3A",X"66",X"FE",X"3A",X"5B",X"5B",X"5B",X"5B",X"3A",X"FE",X"3A",X"FE",
		X"3A",X"FE",X"65",X"4E",X"5B",X"42",X"FE",X"3A",X"FE",X"41",X"4E",X"59",X"3A",X"4C",X"49",X"4B",
		X"45",X"4E",X"45",X"53",X"53",X"3A",X"54",X"4F",X"3A",X"50",X"45",X"52",X"53",X"4F",X"4E",X"53",
		X"FE",X"41",X"4C",X"49",X"56",X"45",X"3A",X"4F",X"52",X"3A",X"44",X"45",X"41",X"44",X"3A",X"49",
		X"53",X"FE",X"43",X"4F",X"49",X"4E",X"43",X"49",X"44",X"45",X"4E",X"54",X"41",X"4C",X"FE",X"3A",
		X"FE",X"3A",X"FE",X"3A",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"50",X"45",X"4E",X"49",X"54",X"45",X"4E",X"54",X"49",X"45",X"52",X"3A",X"44",X"45",X"3A",
		X"43",X"41",X"59",X"45",X"4E",X"4E",X"45",X"3A",X"41",X"FE",X"49",X"4E",X"54",X"45",X"52",X"50",
		X"4F",X"4C",X"FE",X"5B",X"5B",X"5B",X"5B",X"5B",X"FE",X"3A",X"FE",X"3A",X"FE",X"4A",X"4F",X"45",
		X"3A",X"4C",X"45",X"3A",X"42",X"41",X"47",X"4E",X"41",X"52",X"44",X"3A",X"45",X"56",X"41",X"44",
		X"45",X"3A",X"65",X"53",X"54",X"4F",X"50",X"65",X"FE",X"3A",X"FE",X"47",X"41",X"53",X"54",X"4F",
		X"55",X"4E",X"45",X"54",X"3A",X"45",X"54",X"3A",X"50",X"49",X"45",X"52",X"52",X"4F",X"54",X"3A",
		X"41",X"3A",X"53",X"45",X"53",X"FE",X"54",X"52",X"4F",X"55",X"53",X"53",X"45",X"53",X"3A",X"65",
		X"53",X"54",X"4F",X"50",X"65",X"FE",X"3A",X"FE",X"3A",X"FE",X"43",X"48",X"45",X"52",X"43",X"48",
		X"45",X"52",X"41",X"3A",X"50",X"52",X"4F",X"42",X"41",X"42",X"4C",X"45",X"4D",X"45",X"4E",X"54",
		X"3A",X"41",X"FE",X"52",X"45",X"43",X"55",X"50",X"45",X"52",X"45",X"52",X"3A",X"53",X"41",X"43",
		X"53",X"3A",X"44",X"6A",X"4F",X"52",X"3A",X"65",X"53",X"54",X"4F",X"50",X"65",X"FE",X"45",X"54",
		X"3A",X"54",X"45",X"4E",X"54",X"45",X"52",X"41",X"3A",X"44",X"45",X"3A",X"44",X"45",X"4C",X"49",
		X"56",X"52",X"45",X"52",X"FE",X"43",X"4F",X"4D",X"50",X"41",X"52",X"53",X"45",X"3A",X"45",X"4E",
		X"46",X"45",X"52",X"4D",X"45",X"3A",X"41",X"55",X"3A",X"43",X"41",X"43",X"48",X"4F",X"54",X"FE",
		X"3A",X"FE",X"4A",X"4F",X"45",X"3A",X"50",X"41",X"53",X"3A",X"41",X"52",X"4D",X"45",X"3A",X"65",
		X"53",X"54",X"4F",X"50",X"65",X"FE",X"3A",X"FE",X"45",X"53",X"53",X"41",X"49",X"45",X"52",X"41",
		X"3A",X"53",X"55",X"52",X"45",X"4D",X"45",X"4E",X"54",X"3A",X"44",X"45",X"FE",X"50",X"45",X"4E",
		X"45",X"54",X"52",X"45",X"52",X"3A",X"44",X"41",X"4E",X"53",X"3A",X"4C",X"6A",X"41",X"52",X"4D",
		X"55",X"52",X"45",X"52",X"49",X"45",X"FE",X"50",X"4F",X"55",X"52",X"3A",X"53",X"6A",X"45",X"4D",
		X"50",X"41",X"52",X"45",X"52",X"3A",X"44",X"45",X"53",X"FE",X"52",X"45",X"56",X"4F",X"4C",X"56",
		X"45",X"52",X"53",X"3A",X"41",X"3A",X"53",X"49",X"58",X"3A",X"43",X"4F",X"55",X"50",X"53",X"FE",
		X"3A",X"FE",X"47",X"45",X"4E",X"44",X"41",X"52",X"4D",X"45",X"53",X"3A",X"4F",X"4E",X"54",X"3A",
		X"52",X"45",X"43",X"55",X"3A",X"4F",X"52",X"44",X"52",X"45",X"3A",X"44",X"45",X"FE",X"4E",X"45",
		X"3A",X"50",X"41",X"53",X"3A",X"54",X"49",X"52",X"45",X"52",X"3A",X"4C",X"45",X"53",X"3A",X"50",
		X"52",X"45",X"4D",X"49",X"45",X"52",X"53",X"FE",X"3A",X"FE",X"3A",X"FE",X"3A",X"3A",X"3A",X"3A",
		X"3A",X"42",X"4F",X"4E",X"4E",X"45",X"3A",X"43",X"48",X"41",X"4E",X"43",X"45",X"3A",X"66",X"FE",
		X"3A",X"5B",X"5B",X"5B",X"5B",X"3A",X"FE",X"3A",X"FE",X"3A",X"FE",X"65",X"4E",X"5B",X"42",X"FE",
		X"3A",X"FE",X"54",X"4F",X"55",X"54",X"45",X"3A",X"52",X"45",X"53",X"53",X"45",X"4D",X"42",X"4C",
		X"41",X"4E",X"43",X"45",X"3A",X"41",X"56",X"45",X"43",X"3A",X"44",X"45",X"53",X"FE",X"50",X"45",
		X"52",X"53",X"4F",X"4E",X"4E",X"41",X"47",X"45",X"53",X"3A",X"45",X"58",X"49",X"53",X"54",X"41",
		X"4E",X"54",X"53",X"3A",X"4F",X"55",X"FE",X"41",X"59",X"41",X"4E",X"54",X"3A",X"45",X"58",X"49",
		X"53",X"54",X"45",X"53",X"3A",X"4E",X"45",X"3A",X"53",X"41",X"55",X"52",X"41",X"49",X"54",X"3A",
		X"FE",X"45",X"54",X"52",X"45",X"3A",X"51",X"55",X"45",X"3A",X"50",X"55",X"52",X"45",X"3A",X"43",
		X"4F",X"49",X"4E",X"43",X"49",X"44",X"45",X"4E",X"43",X"45",X"FE",X"3A",X"FE",X"3A",X"FE",X"3A",
		X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"4B",X"B0",X"B1",
		X"B2",X"B3",X"4E",X"4F",X"4C",X"4D",X"E0",X"FF",X"DF",X"E5",X"E0",X"FD",X"FA",X"FC",X"49",X"4A",
		X"51",X"52",X"57",X"DE",X"A2",X"C2",X"A2",X"E2",X"40",X"A5",X"E0",X"40",X"A9",X"90",X"43",X"25",
		X"A0",X"43",X"30",X"B0",X"43",X"35",X"B0",X"43",X"3D",X"D0",X"40",X"B4",X"D0",X"41",X"54",X"E0",
		X"41",X"5D",X"D0",X"41",X"D4",X"90",X"FF",X"FF",X"FF",X"44",X"E5",X"A0",X"44",X"EC",X"B0",X"44",
		X"FA",X"D0",X"44",X"9A",X"60",X"44",X"9E",X"D0",X"47",X"05",X"E0",X"47",X"09",X"D0",X"47",X"26",
		X"B0",X"47",X"7E",X"90",X"47",X"7D",X"60",X"46",X"50",X"60",X"46",X"56",X"50",X"FF",X"FF",X"FF",
		X"48",X"A5",X"E0",X"48",X"AC",X"F0",X"49",X"A5",X"E0",X"49",X"AC",X"D0",X"4B",X"2C",X"E0",X"48",
		X"B2",X"70",X"48",X"BA",X"F0",X"48",X"BE",X"D0",X"4B",X"3A",X"D0",X"FF",X"FF",X"FF",X"31",X"A5",
		X"E0",X"31",X"F0",X"E0",X"31",X"FA",X"D0",X"31",X"AC",X"50",X"FF",X"FF",X"FF",X"36",X"D0",X"D0",
		X"37",X"70",X"D0",X"36",X"F9",X"90",X"36",X"79",X"50",X"36",X"CB",X"B0",X"37",X"69",X"A0",X"36",
		X"75",X"A0",X"FF",X"FF",X"FF",X"40",X"A5",X"80",X"40",X"A9",X"80",X"43",X"25",X"80",X"43",X"30",
		X"10",X"43",X"35",X"10",X"43",X"3D",X"80",X"40",X"B4",X"80",X"41",X"54",X"80",X"41",X"5D",X"80",
		X"FF",X"FF",X"FF",X"44",X"E5",X"40",X"44",X"EC",X"10",X"44",X"FA",X"80",X"44",X"9A",X"20",X"44",
		X"9E",X"40",X"47",X"05",X"40",X"47",X"09",X"40",X"47",X"26",X"10",X"47",X"7E",X"10",X"47",X"7D",
		X"40",X"46",X"50",X"20",X"46",X"56",X"40",X"FF",X"FF",X"FF",X"44",X"E5",X"80",X"44",X"EC",X"10",
		X"44",X"FA",X"80",X"44",X"9A",X"20",X"44",X"9E",X"80",X"47",X"05",X"80",X"47",X"09",X"10",X"47",
		X"26",X"20",X"47",X"7E",X"80",X"47",X"7D",X"20",X"46",X"50",X"20",X"46",X"56",X"40",X"FF",X"FF",
		X"FF",X"48",X"A5",X"40",X"48",X"AC",X"10",X"49",X"A5",X"40",X"49",X"AC",X"10",X"4B",X"2C",X"40",
		X"48",X"B2",X"10",X"48",X"BA",X"20",X"48",X"BE",X"40",X"4B",X"3A",X"10",X"FF",X"FF",X"FF",X"48",
		X"A5",X"80",X"48",X"AC",X"10",X"49",X"A5",X"80",X"49",X"AC",X"80",X"4B",X"2C",X"20",X"48",X"B2",
		X"20",X"48",X"BA",X"80",X"48",X"BE",X"80",X"4B",X"3A",X"80",X"FF",X"FF",X"FF",X"31",X"A5",X"40",
		X"31",X"F0",X"20",X"31",X"FA",X"40",X"31",X"AC",X"10",X"FF",X"FF",X"FF",X"31",X"A5",X"80",X"31",
		X"F0",X"20",X"31",X"FA",X"80",X"31",X"AC",X"10",X"FF",X"FF",X"FF",X"36",X"D0",X"40",X"37",X"70",
		X"40",X"36",X"F9",X"80",X"36",X"79",X"10",X"36",X"CB",X"20",X"37",X"69",X"20",X"36",X"75",X"80",
		X"FF",X"FF",X"FF",X"0E",X"10",X"42",X"59",X"10",X"56",X"41",X"4C",X"41",X"44",X"4F",X"4E",X"10",
		X"41",X"55",X"54",X"4F",X"4D",X"41",X"54",X"49",X"4F",X"4E",X"10",X"31",X"39",X"38",X"34",X"3F",
		X"BF",X"BE",X"FF",X"DF",X"DE",X"B0",X"B1",X"B2",X"B3",X"49",X"4A",X"4B",X"51",X"52",X"57",X"53",
		X"4E",X"4F",X"4C",X"4D",X"E0",X"08",X"04",X"02",X"01",X"E0",X"FF",X"DF",X"E9",X"DE",X"49",X"4A",
		X"4B",X"51",X"52",X"57",X"B3",X"B2",X"B1",X"B0",X"8F",X"8E",X"4E",X"4F",X"4D",X"4C",X"FB",X"B3",
		X"B2",X"B1",X"B0",X"4E",X"4F",X"4C",X"4D",X"E0",X"35",X"47",X"35",X"4B",X"35",X"50",X"35",X"55",
		X"35",X"5E",X"FF",X"FF",X"FF",X"1F",X"1F",X"1F",X"FF",X"09",X"00",X"1F",X"1F",X"1F",X"FF",X"1F",
		X"1F",X"1F",X"FF",X"20",X"00",X"1F",X"1F",X"1F",X"FF",X"1F",X"1F",X"1F",X"FF",X"20",X"00",X"1F",
		X"1F",X"1F",X"FF",X"1F",X"1F",X"1F",X"FF",X"30",X"00",X"1F",X"1F",X"1F",X"FF",X"3E",X"01",X"CD",
		X"E2",X"D8",X"06",X"12",X"E5",X"D1",X"7A",X"C6",X"08",X"57",X"3E",X"2C",X"E5",X"12",X"36",X"E0",
		X"13",X"23",X"10",X"F9",X"E1",X"DD",X"21",X"4E",X"25",X"11",X"E0",X"FF",X"19",X"3E",X"2C",X"08",
		X"CD",X"0F",X"25",X"DD",X"21",X"57",X"25",X"CD",X"0F",X"25",X"DD",X"21",X"61",X"25",X"CD",X"0F",
		X"25",X"DD",X"21",X"6B",X"25",X"CD",X"0F",X"25",X"DD",X"21",X"77",X"25",X"CD",X"0F",X"25",X"DD",
		X"21",X"86",X"25",X"CD",X"0F",X"25",X"DD",X"21",X"97",X"25",X"CD",X"0F",X"25",X"3E",X"28",X"08",
		X"DD",X"21",X"A8",X"25",X"CD",X"0F",X"25",X"DD",X"21",X"B9",X"25",X"CD",X"0F",X"25",X"DD",X"21",
		X"CA",X"25",X"CD",X"0F",X"25",X"DD",X"21",X"DB",X"25",X"CD",X"0F",X"25",X"DD",X"21",X"F0",X"25",
		X"CD",X"0F",X"25",X"DD",X"21",X"05",X"26",X"CD",X"0F",X"25",X"DD",X"21",X"1A",X"26",X"CD",X"0F",
		X"25",X"3E",X"18",X"08",X"DD",X"21",X"2F",X"26",X"CD",X"0F",X"25",X"3E",X"1C",X"08",X"FD",X"21",
		X"33",X"25",X"06",X"00",X"FD",X"09",X"FD",X"7E",X"00",X"FE",X"00",X"28",X"1A",X"FE",X"01",X"28",
		X"2C",X"FE",X"02",X"28",X"3E",X"FE",X"03",X"28",X"50",X"FE",X"10",X"28",X"62",X"FE",X"11",X"28",
		X"66",X"FE",X"12",X"28",X"6A",X"18",X"70",X"DD",X"21",X"44",X"26",X"CD",X"0F",X"25",X"DD",X"21",
		X"59",X"26",X"CD",X"0F",X"25",X"DD",X"21",X"63",X"26",X"CD",X"0F",X"25",X"C9",X"DD",X"21",X"82",
		X"26",X"CD",X"0F",X"25",X"DD",X"21",X"97",X"26",X"CD",X"0F",X"25",X"DD",X"21",X"A3",X"26",X"CD",
		X"0F",X"25",X"C9",X"DD",X"21",X"C2",X"26",X"CD",X"0F",X"25",X"DD",X"21",X"D7",X"26",X"CD",X"0F",
		X"25",X"DD",X"21",X"E2",X"26",X"CD",X"0F",X"25",X"C9",X"DD",X"21",X"02",X"27",X"CD",X"0F",X"25",
		X"DD",X"21",X"17",X"27",X"CD",X"0F",X"25",X"DD",X"21",X"21",X"27",X"CD",X"0F",X"25",X"C9",X"DD",
		X"21",X"6D",X"26",X"CD",X"0F",X"25",X"C9",X"DD",X"21",X"AD",X"26",X"CD",X"0F",X"25",X"C9",X"DD",
		X"21",X"ED",X"26",X"CD",X"0F",X"25",X"C9",X"DD",X"21",X"2B",X"27",X"CD",X"0F",X"25",X"C9",X"E5",
		X"DD",X"7E",X"00",X"DD",X"23",X"B9",X"41",X"30",X"01",X"47",X"78",X"FE",X"00",X"C8",X"DD",X"7E",
		X"00",X"77",X"E5",X"7C",X"C6",X"08",X"67",X"08",X"77",X"08",X"E1",X"19",X"DD",X"23",X"10",X"EA",
		X"E1",X"23",X"C9",X"13",X"03",X"12",X"02",X"11",X"01",X"13",X"03",X"12",X"02",X"11",X"01",X"13",
		X"03",X"12",X"02",X"11",X"01",X"13",X"03",X"12",X"02",X"11",X"01",X"13",X"03",X"00",X"08",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"01",X"02",X"09",X"E0",X"E0",X"03",X"04",X"05",X"06",X"07",X"08",
		X"09",X"09",X"E0",X"E0",X"0A",X"0B",X"0C",X"0D",X"6A",X"0F",X"62",X"0B",X"E0",X"E0",X"11",X"12",
		X"13",X"6C",X"6B",X"00",X"17",X"18",X"19",X"0E",X"1A",X"1B",X"1C",X"1D",X"72",X"9B",X"AD",X"B2",
		X"22",X"23",X"24",X"25",X"26",X"27",X"10",X"28",X"29",X"2A",X"2B",X"2C",X"2D",X"2E",X"2F",X"30",
		X"31",X"32",X"33",X"34",X"35",X"36",X"4D",X"10",X"37",X"38",X"39",X"3A",X"3B",X"3C",X"3D",X"3E",
		X"3F",X"40",X"41",X"42",X"43",X"44",X"45",X"50",X"10",X"46",X"47",X"48",X"49",X"4A",X"4B",X"4C",
		X"47",X"4E",X"4F",X"47",X"51",X"52",X"47",X"54",X"55",X"10",X"56",X"57",X"58",X"59",X"5A",X"5B",
		X"5C",X"5D",X"5E",X"5F",X"60",X"61",X"A2",X"63",X"64",X"65",X"10",X"66",X"67",X"68",X"69",X"5A",
		X"5B",X"5C",X"6D",X"6E",X"6F",X"70",X"71",X"A2",X"73",X"74",X"75",X"14",X"76",X"77",X"78",X"79",
		X"7A",X"7B",X"7C",X"7D",X"7E",X"7F",X"80",X"81",X"82",X"83",X"84",X"85",X"86",X"87",X"88",X"89",
		X"14",X"8A",X"8B",X"8C",X"8D",X"8E",X"8F",X"90",X"91",X"92",X"93",X"94",X"95",X"96",X"97",X"98",
		X"99",X"9A",X"99",X"9C",X"9D",X"14",X"9E",X"9F",X"A0",X"A1",X"A2",X"A3",X"A4",X"A5",X"A6",X"A7",
		X"A8",X"A9",X"AA",X"AB",X"AC",X"A2",X"AE",X"AF",X"B0",X"B1",X"14",X"9E",X"B3",X"B4",X"B5",X"B6",
		X"B7",X"A4",X"B9",X"A2",X"BB",X"BC",X"A2",X"BE",X"AB",X"C0",X"C1",X"C2",X"C3",X"53",X"B1",X"14",
		X"92",X"93",X"94",X"95",X"96",X"97",X"98",X"99",X"9A",X"9B",X"9C",X"9D",X"9E",X"9F",X"A0",X"A1",
		X"A2",X"A3",X"A4",X"A5",X"14",X"BD",X"BC",X"1F",X"20",X"B8",X"BB",X"AD",X"BC",X"BC",X"BC",X"BF",
		X"BC",X"C0",X"BC",X"BC",X"C1",X"BC",X"C2",X"BD",X"C3",X"09",X"91",X"91",X"25",X"26",X"B9",X"B1",
		X"B2",X"B6",X"B7",X"09",X"91",X"91",X"2D",X"2E",X"BA",X"B4",X"B5",X"1B",X"1C",X"14",X"BD",X"1F",
		X"20",X"B8",X"BB",X"AD",X"BC",X"BC",X"BC",X"BC",X"BF",X"BC",X"C0",X"BC",X"BC",X"C1",X"BC",X"C2",
		X"BD",X"C3",X"14",X"BD",X"BC",X"BC",X"00",X"01",X"02",X"03",X"04",X"05",X"06",X"07",X"BC",X"C0",
		X"BC",X"BC",X"C1",X"BC",X"C2",X"BD",X"C3",X"0B",X"91",X"91",X"08",X"09",X"0A",X"0B",X"0C",X"0D",
		X"0E",X"0F",X"10",X"09",X"91",X"91",X"11",X"12",X"13",X"1B",X"1C",X"1D",X"1E",X"14",X"BD",X"BC",
		X"00",X"01",X"02",X"03",X"04",X"05",X"06",X"07",X"BC",X"BC",X"C0",X"BC",X"BC",X"C1",X"BC",X"C2",
		X"BD",X"C3",X"14",X"BD",X"BC",X"1F",X"20",X"21",X"22",X"23",X"24",X"BC",X"BC",X"BF",X"BC",X"C0",
		X"BC",X"BC",X"C1",X"BC",X"C2",X"BD",X"C3",X"0A",X"91",X"91",X"25",X"26",X"27",X"28",X"29",X"2A",
		X"2B",X"2C",X"0A",X"91",X"91",X"2D",X"2E",X"2F",X"91",X"30",X"A6",X"A7",X"A8",X"14",X"BD",X"1F",
		X"20",X"21",X"22",X"23",X"24",X"BC",X"BC",X"BC",X"BF",X"BC",X"C0",X"BC",X"BC",X"C1",X"BC",X"C2",
		X"BD",X"C3",X"14",X"BD",X"BC",X"A9",X"AA",X"AB",X"AC",X"AD",X"BC",X"BC",X"BC",X"BF",X"BC",X"C0",
		X"BC",X"BC",X"C1",X"BC",X"C2",X"BD",X"C3",X"09",X"91",X"91",X"AE",X"AF",X"B0",X"B1",X"B2",X"B6",
		X"B7",X"09",X"91",X"91",X"91",X"91",X"B3",X"B4",X"B5",X"1B",X"1C",X"14",X"BD",X"A9",X"AA",X"AB",
		X"AC",X"AD",X"BC",X"BC",X"BC",X"BC",X"BF",X"BC",X"C0",X"BC",X"BC",X"C1",X"BC",X"C2",X"BD",X"C3",
		X"DA",X"D9",X"D8",X"D7",X"D6",X"D5",X"D4",X"D3",X"D2",X"D1",X"D0",X"CF",X"CE",X"CD",X"CC",X"CB",
		X"C9",X"C8",X"23",X"22",X"21",X"22",X"23",X"21",X"22",X"23",X"22",X"21",X"23",X"21",X"22",X"23",
		X"21",X"22",X"23",X"21",X"22",X"23",X"22",X"21",X"22",X"23",X"21",X"22",X"23",X"22",X"21",X"23",
		X"21",X"22",X"23",X"21",X"22",X"23",X"21",X"22",X"FF",X"18",X"17",X"16",X"15",X"14",X"15",X"14",
		X"16",X"15",X"16",X"14",X"15",X"14",X"16",X"15",X"14",X"16",X"15",X"14",X"FF",X"FF",X"70",X"F7",
		X"DF",X"FF",X"B9",X"C0",X"FC",X"FF",X"18",X"A0",X"99",X"F7",X"48",X"04",X"FF",X"DF",X"70",X"F2",
		X"F1",X"EF",X"10",X"30",X"A9",X"FB",X"08",X"0D",X"39",X"F3",X"20",X"3C",X"FD",X"F5",X"A9",X"51",
		X"F1",X"FF",X"08",X"34",X"FB",X"FF",X"B8",X"04",X"F1",X"FA",X"00",X"04",X"9D",X"2B",X"00",X"04",
		X"BF",X"BF",X"2D",X"75",X"E9",X"DF",X"C0",X"46",X"79",X"BE",X"28",X"94",X"FB",X"FF",X"F7",X"E7",
		X"FD",X"FF",X"09",X"7A",X"CB",X"FF",X"09",X"B0",X"DC",X"7F",X"B4",X"62",X"7D",X"F9",X"0C",X"8C",
		X"CA",X"D2",X"40",X"C5",X"DC",X"EB",X"48",X"21",X"EC",X"7E",X"84",X"14",X"F5",X"FD",X"59",X"F4",
		X"E8",X"6D",X"30",X"AD",X"EC",X"F6",X"20",X"D6",X"B8",X"FB",X"40",X"24",X"BC",X"2A",X"00",X"01",
		X"7F",X"FF",X"EB",X"EB",X"6D",X"AF",X"2A",X"27",X"FF",X"F7",X"9F",X"E5",X"BE",X"F7",X"9C",X"7C",
		X"FF",X"FF",X"54",X"DB",X"FE",X"FF",X"ED",X"76",X"9B",X"FF",X"9D",X"B6",X"23",X"F7",X"0B",X"05",
		X"14",X"FF",X"0B",X"88",X"E2",X"A3",X"00",X"60",X"EF",X"DF",X"9A",X"F6",X"FD",X"EF",X"1E",X"A6",
		X"BF",X"EA",X"2E",X"02",X"8D",X"AE",X"02",X"E6",X"D7",X"FF",X"8C",X"08",X"3D",X"AF",X"04",X"A8",
		X"DF",X"EF",X"AC",X"B6",X"AF",X"A7",X"A1",X"04",X"FD",X"FF",X"65",X"6D",X"FF",X"EF",X"3F",X"6E",
		X"BF",X"7F",X"CB",X"C2",X"FF",X"E3",X"8F",X"A5",X"FF",X"BF",X"9F",X"A7",X"BF",X"FF",X"20",X"88",
		X"7F",X"F6",X"00",X"14",X"99",X"27",X"12",X"A0",X"BF",X"FF",X"9B",X"F3",X"BF",X"EF",X"D3",X"80",
		X"0F",X"57",X"0F",X"62",X"F5",X"A6",X"44",X"A8",X"BF",X"FB",X"A4",X"20",X"25",X"A4",X"08",X"84",
		X"B7",X"CB",X"34",X"44",X"F7",X"FD",X"87",X"64",X"EF",X"FF",X"95",X"66",X"F7",X"FF",X"03",X"C9",
		X"EF",X"FD",X"97",X"B5",X"FF",X"EF",X"BF",X"69",X"57",X"6F",X"47",X"01",X"EF",X"EF",X"87",X"09",
		X"97",X"6F",X"04",X"40",X"55",X"CB",X"07",X"09",X"B7",X"8A",X"34",X"00",X"C7",X"EF",X"45",X"04",
		X"5F",X"AD",X"47",X"01",X"FF",X"FF",X"27",X"01",X"37",X"47",X"07",X"40",X"AD",X"CF",X"45",X"85",
		X"E7",X"ED",X"C2",X"55",X"B7",X"DD",X"1C",X"01",X"C7",X"F5",X"EB",X"4E",X"97",X"FF",X"1E",X"8C",
		X"FF",X"DF",X"1E",X"8F",X"EF",X"FD",X"0F",X"08",X"BF",X"0F",X"97",X"60",X"A7",X"BF",X"87",X"0E",
		X"87",X"14",X"00",X"00",X"0F",X"DF",X"00",X"08",X"2E",X"CE",X"51",X"48",X"D7",X"CF",X"02",X"00",
		X"9F",X"CD",X"87",X"08",X"E7",X"8F",X"3F",X"50",X"95",X"6D",X"01",X"08",X"6F",X"BD",X"05",X"C0",
		X"FD",X"A7",X"64",X"2E",X"BF",X"FF",X"1D",X"FB",X"BF",X"FF",X"17",X"B6",X"FF",X"FE",X"CA",X"0E",
		X"DF",X"FF",X"81",X"63",X"BC",X"BE",X"AB",X"86",X"FF",X"FF",X"8F",X"DF",X"9F",X"EF",X"07",X"A6",
		X"1B",X"6F",X"02",X"40",X"ED",X"D7",X"02",X"02",X"FF",X"B7",X"4C",X"13",X"F9",X"EF",X"06",X"AF",
		X"8D",X"36",X"28",X"81",X"9D",X"EF",X"06",X"24",X"FF",X"DF",X"9F",X"1A",X"2F",X"8F",X"02",X"35",
		X"3F",X"FF",X"26",X"A2",X"BF",X"E7",X"A8",X"00",X"EF",X"FF",X"67",X"A2",X"AE",X"8F",X"9B",X"25",
		X"0D",X"F7",X"84",X"19",X"FF",X"F5",X"9F",X"0C",X"BD",X"FF",X"2E",X"B6",X"FF",X"AF",X"4A",X"87",
		X"6F",X"BC",X"00",X"85",X"3F",X"AD",X"A2",X"E0",X"BF",X"AF",X"0E",X"BB",X"DB",X"FF",X"1C",X"2E",
		X"5E",X"A6",X"03",X"40",X"CC",X"FE",X"89",X"80",X"BD",X"F9",X"86",X"E5",X"9F",X"EF",X"2E",X"86",
		X"9F",X"FB",X"8D",X"88",X"BF",X"2F",X"C7",X"81",X"FF",X"FF",X"AF",X"C3",X"F7",X"EF",X"85",X"C9",
		X"AF",X"3F",X"87",X"B6",X"9F",X"DF",X"0F",X"48",X"FF",X"E9",X"B7",X"80",X"FF",X"EF",X"FF",X"CF",
		X"87",X"D7",X"87",X"09",X"6F",X"57",X"44",X"01",X"D7",X"A7",X"0F",X"48",X"FF",X"FB",X"08",X"54",
		X"FF",X"4B",X"04",X"01",X"DF",X"D7",X"05",X"00",X"A7",X"C5",X"17",X"43",X"A7",X"CF",X"C6",X"48",
		X"FF",X"DD",X"8F",X"63",X"AF",X"BF",X"97",X"2E",X"BF",X"5D",X"A1",X"87",X"D7",X"E9",X"27",X"61",
		X"BF",X"4F",X"87",X"C5",X"FF",X"57",X"C7",X"8D",X"27",X"E3",X"2D",X"CC",X"FF",X"FF",X"8F",X"E9",
		X"37",X"AF",X"03",X"45",X"CF",X"5F",X"04",X"14",X"F7",X"6D",X"2D",X"42",X"AF",X"11",X"84",X"C4",
		X"3F",X"CD",X"4F",X"08",X"55",X"4F",X"8D",X"01",X"C7",X"0B",X"04",X"0C",X"AF",X"DF",X"94",X"47",
		X"BF",X"FF",X"45",X"56",X"FF",X"F7",X"AF",X"56",X"9F",X"FF",X"AE",X"5F",X"FF",X"BF",X"88",X"CF",
		X"BB",X"67",X"ED",X"A5",X"FF",X"BF",X"2D",X"A5",X"FF",X"EB",X"0C",X"05",X"5F",X"F7",X"97",X"A6",
		X"EF",X"FF",X"00",X"A5",X"AF",X"FB",X"3C",X"C2",X"9F",X"BF",X"CC",X"EE",X"34",X"F6",X"06",X"08",
		X"33",X"A7",X"A4",X"AA",X"DD",X"FF",X"86",X"A6",X"CF",X"56",X"00",X"00",X"5D",X"F7",X"27",X"BC",
		X"FB",X"EF",X"32",X"6E",X"FF",X"DE",X"23",X"E4",X"FF",X"E7",X"DF",X"CE",X"B7",X"E7",X"64",X"FE",
		X"8F",X"BE",X"0D",X"B6",X"BF",X"FF",X"B6",X"36",X"1F",X"BC",X"8C",X"CE",X"FF",X"BF",X"0F",X"E7",
		X"AF",X"F7",X"84",X"0A",X"6D",X"ED",X"20",X"4A",X"FF",X"AF",X"AF",X"04",X"97",X"9E",X"87",X"00",
		X"7D",X"77",X"00",X"10",X"1F",X"A6",X"08",X"23",X"2C",X"07",X"04",X"80",X"FF",X"FF",X"20",X"84",
		X"FF",X"FD",X"0F",X"36",X"BF",X"DF",X"97",X"C0",X"FF",X"FF",X"F7",X"C9",X"F7",X"FF",X"EF",X"CF",
		X"A7",X"8D",X"46",X"39",X"FF",X"EF",X"A7",X"8D",X"EF",X"F7",X"25",X"19",X"BF",X"FF",X"CF",X"0D",
		X"DF",X"77",X"2C",X"89",X"3D",X"5D",X"06",X"08",X"6E",X"BF",X"9D",X"8B",X"5F",X"4D",X"85",X"01",
		X"C7",X"C9",X"00",X"00",X"DF",X"E5",X"93",X"15",X"77",X"4F",X"05",X"01",X"EF",X"7F",X"9E",X"11",
		X"FF",X"DF",X"57",X"11",X"FF",X"4F",X"07",X"11",X"B7",X"EF",X"1E",X"5D",X"C7",X"DF",X"9D",X"D5",
		X"77",X"AF",X"00",X"40",X"9F",X"FF",X"BE",X"8A",X"9F",X"87",X"97",X"43",X"FF",X"FD",X"3E",X"DE",
		X"8F",X"A9",X"45",X"40",X"87",X"85",X"01",X"88",X"AE",X"6F",X"00",X"77",X"1F",X"1F",X"87",X"05",
		X"0F",X"5A",X"04",X"08",X"D7",X"8D",X"47",X"50",X"2F",X"85",X"01",X"8C",X"97",X"97",X"8F",X"03",
		X"FD",X"BD",X"0B",X"06",X"AF",X"FF",X"DE",X"A4",X"FF",X"EF",X"3F",X"7F",X"DF",X"BF",X"2E",X"0E",
		X"3F",X"FE",X"2F",X"29",X"BF",X"F7",X"2B",X"22",X"BF",X"FF",X"9E",X"E4",X"BF",X"F7",X"B6",X"9F",
		X"EC",X"92",X"0C",X"21",X"3F",X"FF",X"0A",X"E4",X"B7",X"FF",X"98",X"BD",X"89",X"F7",X"3D",X"84",
		X"3F",X"CF",X"0D",X"C1",X"EF",X"4F",X"08",X"26",X"DF",X"B7",X"1D",X"84",X"BF",X"BF",X"4C",X"2E",
		X"4E",X"EC",X"21",X"26",X"AF",X"FF",X"0F",X"05",X"A7",X"FF",X"A5",X"6E",X"EF",X"F7",X"2E",X"A6",
		X"BF",X"AF",X"05",X"DF",X"28",X"FE",X"27",X"0F",X"BF",X"FF",X"A6",X"F7",X"EF",X"BF",X"E7",X"A6",
		X"0E",X"B3",X"82",X"24",X"BC",X"AA",X"07",X"14",X"7F",X"C7",X"1C",X"21",X"85",X"35",X"02",X"06",
		X"9F",X"F7",X"08",X"A0",X"36",X"F5",X"82",X"06",X"BE",X"E6",X"CC",X"01",X"0F",X"3F",X"02",X"65",
		X"D7",X"E5",X"04",X"09",X"FF",X"BF",X"94",X"49",X"FF",X"FF",X"07",X"0B",X"FF",X"FF",X"97",X"55",
		X"BF",X"5F",X"25",X"33",X"F7",X"EF",X"A7",X"C1",X"FF",X"FD",X"4F",X"4E",X"FF",X"FF",X"9D",X"C1",
		X"37",X"65",X"87",X"40",X"5F",X"D7",X"0E",X"07",X"9F",X"ED",X"05",X"44",X"CF",X"77",X"0F",X"00",
		X"A7",X"59",X"07",X"02",X"BD",X"BF",X"06",X"16",X"F7",X"ED",X"84",X"54",X"D7",X"FD",X"87",X"8C",
		X"C7",X"45",X"03",X"E1",X"FF",X"4E",X"5F",X"4C",X"5F",X"BF",X"85",X"16",X"FF",X"CF",X"F1",X"95",
		X"CB",X"9F",X"8F",X"02",X"EF",X"DF",X"47",X"C3",X"CF",X"5F",X"A1",X"CF",X"F7",X"FF",X"9D",X"49",
		X"0F",X"CD",X"01",X"08",X"D7",X"49",X"07",X"20",X"FF",X"EF",X"04",X"41",X"A7",X"8B",X"86",X"05",
		X"CF",X"ED",X"0F",X"45",X"CF",X"DF",X"A5",X"42",X"9F",X"EC",X"07",X"00",X"DF",X"8D",X"40",X"25",
		X"FF",X"FF",X"40",X"76",X"AF",X"B6",X"08",X"08",X"FF",X"EF",X"05",X"25",X"BE",X"FF",X"2E",X"C6",
		X"EF",X"A7",X"03",X"82",X"AF",X"B7",X"0C",X"14",X"FF",X"FF",X"B6",X"BF",X"3F",X"E7",X"40",X"A8",
		X"0F",X"BE",X"0F",X"04",X"01",X"16",X"00",X"00",X"3F",X"AB",X"86",X"66",X"EF",X"DF",X"04",X"20",
		X"1D",X"EF",X"29",X"40",X"E9",X"E5",X"0D",X"00",X"FF",X"FF",X"91",X"A2",X"0C",X"EE",X"16",X"04",
		X"BD",X"BF",X"6A",X"A6",X"26",X"8B",X"09",X"04",X"BD",X"EF",X"0F",X"E6",X"FF",X"EF",X"0D",X"FF",
		X"37",X"B3",X"9A",X"0E",X"EF",X"BD",X"82",X"B5",X"FF",X"FF",X"CD",X"22",X"F7",X"A5",X"A4",X"8A",
		X"5F",X"4F",X"07",X"82",X"65",X"06",X"04",X"04",X"FF",X"EA",X"94",X"61",X"AF",X"AE",X"4C",X"C2",
		X"9B",X"86",X"04",X"C0",X"DD",X"C6",X"84",X"80",X"6D",X"EF",X"06",X"A6",X"0F",X"EE",X"00",X"24",
		X"E3",X"D5",X"0F",X"C8",X"CF",X"D7",X"B5",X"01",X"FF",X"CF",X"03",X"0D",X"BF",X"89",X"86",X"04",
		X"DF",X"DF",X"D7",X"32",X"DF",X"1D",X"BF",X"51",X"A4",X"87",X"C5",X"40",X"ED",X"8F",X"C6",X"C1",
		X"9F",X"E3",X"10",X"00",X"87",X"89",X"05",X"40",X"17",X"3B",X"00",X"01",X"AF",X"49",X"84",X"00",
		X"FF",X"ED",X"47",X"61",X"77",X"FF",X"07",X"25",X"0F",X"75",X"05",X"04",X"97",X"F9",X"C0",X"50",
		X"EF",X"4C",X"05",X"49",X"27",X"0B",X"07",X"70",X"3F",X"59",X"03",X"85",X"FF",X"CD",X"27",X"04",
		X"CF",X"FF",X"8F",X"C9",X"7F",X"BD",X"C6",X"4B",X"FF",X"DF",X"04",X"85",X"87",X"DF",X"07",X"15",
		X"A7",X"41",X"04",X"0D",X"9F",X"44",X"03",X"08",X"F7",X"8D",X"01",X"41",X"87",X"0B",X"04",X"10",
		X"CD",X"4F",X"44",X"29",X"9F",X"85",X"05",X"46",X"0A",X"1C",X"04",X"08",X"B6",X"4D",X"8A",X"40",
		X"3F",X"BE",X"00",X"12",X"AF",X"3F",X"00",X"02",X"BF",X"EF",X"3B",X"AA",X"77",X"EE",X"94",X"14",
		X"DB",X"C7",X"84",X"24",X"8D",X"F7",X"2D",X"28",X"ED",X"FF",X"9F",X"AA",X"DF",X"F7",X"18",X"46",
		X"9C",X"64",X"10",X"00",X"DD",X"15",X"00",X"20",X"7B",X"2F",X"38",X"A4",X"2F",X"7E",X"12",X"54",
		X"9C",X"7E",X"04",X"20",X"AE",X"A5",X"08",X"50",X"17",X"F7",X"0B",X"E6",X"1E",X"F6",X"0C",X"84",
		X"BC",X"43",X"09",X"00",X"6F",X"CF",X"04",X"28",X"7F",X"B7",X"24",X"20",X"3F",X"FF",X"1B",X"8E",
		X"1B",X"D5",X"0C",X"26",X"1F",X"FB",X"25",X"64",X"FF",X"A7",X"A5",X"C2",X"2E",X"BF",X"0F",X"06",
		X"C7",X"E6",X"11",X"30",X"2C",X"A9",X"8C",X"80",X"96",X"9C",X"22",X"26",X"3D",X"A7",X"01",X"24",
		X"1F",X"23",X"04",X"21",X"1C",X"FE",X"86",X"24",X"8F",X"AF",X"02",X"06",X"8B",X"66",X"0A",X"30",
		X"97",X"67",X"87",X"17",X"BF",X"CF",X"0F",X"A2",X"FF",X"FF",X"0F",X"AB",X"FF",X"DD",X"FE",X"41",
		X"3F",X"F7",X"0C",X"10",X"9F",X"7F",X"03",X"09",X"9F",X"7D",X"02",X"40",X"F7",X"FD",X"CF",X"7D",
		X"C7",X"4B",X"05",X"D5",X"CF",X"45",X"05",X"40",X"1F",X"6F",X"17",X"88",X"8F",X"E3",X"95",X"00",
		X"1D",X"95",X"04",X"00",X"07",X"44",X"00",X"04",X"2F",X"B0",X"00",X"00",X"FF",X"E5",X"C6",X"09",
		X"DF",X"4F",X"0F",X"19",X"C7",X"F5",X"3E",X"04",X"9F",X"FF",X"67",X"20",X"DF",X"CF",X"9D",X"45",
		X"9D",X"7B",X"47",X"05",X"37",X"E9",X"CE",X"45",X"35",X"57",X"81",X"90",X"F7",X"FF",X"03",X"5D",
		X"54",X"CB",X"AF",X"2D",X"AF",X"28",X"26",X"00",X"9D",X"DF",X"07",X"80",X"EF",X"A7",X"05",X"08",
		X"6D",X"0D",X"04",X"00",X"97",X"45",X"04",X"04",X"C1",X"86",X"00",X"14",X"F7",X"5D",X"86",X"00",
		X"FF",X"FF",X"08",X"9F",X"AF",X"BF",X"A5",X"B4",X"BF",X"CF",X"9F",X"DB",X"BF",X"BF",X"27",X"EE",
		X"7D",X"37",X"1F",X"A6",X"BF",X"F7",X"80",X"8E",X"ED",X"6C",X"00",X"D4",X"BA",X"FF",X"57",X"E3",
		X"E7",X"E2",X"08",X"82",X"5B",X"3F",X"60",X"20",X"AF",X"F6",X"0E",X"01",X"23",X"AF",X"84",X"96",
		X"AF",X"BF",X"06",X"A2",X"2F",X"A4",X"84",X"02",X"B8",X"92",X"01",X"A0",X"BF",X"AF",X"04",X"90",
		X"BF",X"FE",X"8F",X"6C",X"FD",X"BA",X"FD",X"B2",X"BF",X"FF",X"8F",X"A5",X"FF",X"D7",X"06",X"90",
		X"B7",X"F7",X"8D",X"32",X"AD",X"AF",X"08",X"94",X"BF",X"AF",X"01",X"A4",X"BF",X"FE",X"BD",X"BB",
		X"A7",X"E6",X"9D",X"03",X"8E",X"EF",X"AC",X"21",X"77",X"FF",X"85",X"A7",X"37",X"9C",X"04",X"60",
		X"C9",X"EF",X"A6",X"7C",X"DE",X"EE",X"2A",X"0F",X"01",X"36",X"06",X"20",X"4C",X"F5",X"25",X"06",
		X"BF",X"C7",X"E3",X"0C",X"DF",X"BF",X"05",X"4B",X"FF",X"FF",X"AF",X"07",X"DF",X"DF",X"DE",X"04",
		X"A5",X"1D",X"01",X"19",X"BF",X"CF",X"B7",X"51",X"95",X"89",X"0D",X"80",X"FF",X"DF",X"C7",X"79",
		X"AF",X"57",X"2F",X"09",X"67",X"DF",X"0A",X"08",X"BF",X"C4",X"81",X"41",X"EF",X"16",X"05",X"02",
		X"A5",X"87",X"04",X"00",X"EF",X"0F",X"0C",X"4C",X"D7",X"C9",X"C7",X"25",X"F7",X"ED",X"87",X"89",
		X"F7",X"EF",X"E5",X"95",X"67",X"BF",X"4F",X"24",X"9F",X"3F",X"1F",X"CB",X"AF",X"DF",X"9C",X"01",
		X"47",X"49",X"10",X"00",X"57",X"FF",X"45",X"C2",X"57",X"1D",X"07",X"01",X"BF",X"EF",X"A5",X"90",
		X"B5",X"27",X"83",X"41",X"55",X"8F",X"57",X"01",X"1F",X"7D",X"04",X"44",X"8F",X"C5",X"04",X"05",
		X"91",X"80",X"01",X"00",X"CF",X"88",X"80",X"60",X"EC",X"69",X"05",X"00",X"C5",X"CF",X"97",X"01",
		X"8F",X"FF",X"2D",X"06",X"BF",X"EF",X"44",X"A1",X"ED",X"B7",X"8B",X"05",X"2D",X"F7",X"2A",X"AE",
		X"B7",X"EF",X"05",X"04",X"A5",X"24",X"E6",X"29",X"FF",X"FF",X"13",X"4F",X"3F",X"FF",X"6A",X"A6",
		X"7B",X"A3",X"00",X"80",X"CE",X"A7",X"04",X"04",X"3D",X"CF",X"84",X"80",X"9B",X"FD",X"00",X"06",
		X"AF",X"E6",X"0B",X"76",X"04",X"A6",X"00",X"04",X"FD",X"B2",X"28",X"27",X"2D",X"86",X"A1",X"04",
		X"4F",X"A7",X"20",X"A1",X"3F",X"FF",X"0D",X"62",X"AF",X"A6",X"B4",X"47",X"E7",X"EF",X"29",X"A0",
		X"DB",X"CF",X"0C",X"8A",X"AD",X"07",X"04",X"04",X"BF",X"F7",X"C8",X"3B",X"DF",X"F7",X"0E",X"24",
		X"34",X"A4",X"0A",X"02",X"B4",X"BD",X"08",X"A2",X"9F",X"E2",X"80",X"C0",X"34",X"F7",X"8C",X"05",
		X"BF",X"BD",X"81",X"6A",X"09",X"AE",X"00",X"00",X"7F",X"36",X"23",X"0B",X"3F",X"F9",X"88",X"26",
		X"8F",X"81",X"67",X"00",X"F7",X"D5",X"05",X"05",X"EF",X"AF",X"87",X"85",X"CF",X"8F",X"BC",X"84",
		X"BF",X"7B",X"0A",X"01",X"FF",X"AF",X"17",X"47",X"FF",X"17",X"41",X"98",X"EF",X"CF",X"97",X"4F",
		X"82",X"05",X"24",X"00",X"9F",X"69",X"86",X"04",X"8F",X"9B",X"17",X"94",X"C7",X"6F",X"42",X"09",
		X"AD",X"AF",X"44",X"0D",X"BF",X"2B",X"83",X"84",X"DD",X"0B",X"01",X"41",X"DF",X"F7",X"17",X"45",
		X"85",X"2F",X"07",X"44",X"F7",X"AD",X"06",X"81",X"E7",X"9D",X"FF",X"45",X"FD",X"BF",X"81",X"0D",
		X"FF",X"E9",X"97",X"01",X"AF",X"ED",X"96",X"25",X"B7",X"2E",X"07",X"A6",X"ED",X"FF",X"A7",X"A4",
		X"17",X"C9",X"20",X"01",X"44",X"4D",X"06",X"42",X"BB",X"5D",X"0D",X"08",X"2E",X"C9",X"07",X"04",
		X"DF",X"87",X"00",X"40",X"47",X"DD",X"04",X"00",X"25",X"8E",X"06",X"CE",X"5C",X"A7",X"97",X"58",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"46",X"E0",X"E0",
		X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"46",X"E0",X"E0",X"DB",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"46",X"E0",X"E0",
		X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"46",X"E0",X"E0",X"DB",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"46",X"E0",X"E0",
		X"50",X"13",X"DB",X"DB",X"DB",X"DB",X"DB",X"46",X"DB",X"DB",X"0F",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"81",X"4A",X"E0",X"50",X"DB",X"12",X"DB",X"DB",X"DB",X"0E",X"DB",X"46",X"4A",X"E0",
		X"50",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"46",X"E0",X"E0",X"50",X"46",X"4A",X"E0",X"50",X"E0",
		X"E0",X"E0",X"82",X"4B",X"49",X"5A",X"DB",X"5A",X"DB",X"5A",X"0F",X"5A",X"5A",X"46",X"4B",X"49",
		X"50",X"5A",X"DB",X"5A",X"DB",X"5A",X"DB",X"46",X"4A",X"E0",X"5A",X"46",X"4B",X"49",X"50",X"E0",
		X"E0",X"E0",X"82",X"E0",X"E0",X"5B",X"5A",X"5B",X"5A",X"5B",X"5A",X"5B",X"5B",X"46",X"E0",X"E0",
		X"5A",X"5B",X"5A",X"5B",X"5A",X"5B",X"5A",X"46",X"4B",X"49",X"5B",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"82",X"4C",X"4E",X"4C",X"4E",X"4C",X"4E",X"4C",X"4E",X"4C",X"4E",X"4C",X"4E",X"4C",
		X"4E",X"4C",X"4E",X"4C",X"4E",X"4C",X"4E",X"4C",X"4E",X"4C",X"4E",X"4C",X"4E",X"4C",X"50",X"E0",
		X"E0",X"E0",X"82",X"4D",X"4F",X"4D",X"4F",X"4D",X"4F",X"4D",X"4F",X"4D",X"4F",X"4D",X"4F",X"4D",
		X"4F",X"4D",X"4F",X"4D",X"4F",X"4D",X"4F",X"4D",X"4F",X"4D",X"4F",X"4D",X"4F",X"4D",X"50",X"E0",
		X"E0",X"E0",X"82",X"E0",X"E0",X"5A",X"5B",X"5A",X"5B",X"5A",X"5B",X"5A",X"5B",X"46",X"E0",X"E0",
		X"5A",X"5B",X"5A",X"5B",X"5A",X"5B",X"5A",X"46",X"4A",X"E0",X"BF",X"46",X"4A",X"E0",X"50",X"E0",
		X"E0",X"E0",X"82",X"E0",X"E0",X"5B",X"5A",X"5B",X"0F",X"5B",X"DB",X"5B",X"DB",X"46",X"E0",X"E0",
		X"5B",X"DB",X"5B",X"0C",X"5B",X"DB",X"5B",X"46",X"4B",X"49",X"BF",X"46",X"4B",X"49",X"50",X"E0",
		X"E0",X"E0",X"82",X"E0",X"E0",X"50",X"5B",X"5A",X"DB",X"12",X"DB",X"DB",X"DB",X"46",X"E0",X"E0",
		X"50",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"46",X"E0",X"E0",X"BF",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"82",X"E0",X"E0",X"50",X"0D",X"5B",X"DB",X"DB",X"DB",X"0C",X"DB",X"46",X"E0",X"E0",
		X"50",X"DB",X"0E",X"DB",X"DB",X"DB",X"DB",X"46",X"E0",X"E0",X"BF",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"82",X"E0",X"DF",X"FB",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"DB",X"46",X"4A",X"E0",
		X"50",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"46",X"E0",X"E0",X"BF",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"82",X"E0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"50",X"46",X"4B",X"49",
		X"50",X"DB",X"DB",X"DB",X"13",X"DB",X"DB",X"46",X"E0",X"E0",X"BF",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"82",X"E0",X"DE",X"FA",X"FD",X"FD",X"FD",X"FC",X"DE",X"DE",X"50",X"46",X"E0",X"DF",
		X"FB",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"F9",X"DF",X"DF",X"BF",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"82",X"4A",X"E0",X"50",X"DB",X"DB",X"DB",X"46",X"E0",X"E0",X"50",X"46",X"E0",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"83",X"4B",X"49",X"50",X"DB",X"0F",X"DB",X"46",X"E0",X"E0",X"50",X"46",X"E0",X"DE",
		X"FA",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FC",X"DE",X"DE",X"BF",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"DB",X"DB",X"DB",X"46",X"4A",X"E0",X"50",X"46",X"E0",X"E0",
		X"50",X"DB",X"DB",X"DB",X"DB",X"44",X"DB",X"46",X"4A",X"E0",X"BF",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"13",X"DB",X"DB",X"46",X"4B",X"49",X"50",X"46",X"E0",X"E0",
		X"50",X"DB",X"DB",X"0D",X"DB",X"45",X"DB",X"46",X"4B",X"49",X"BF",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"DB",X"DB",X"DB",X"46",X"E0",X"E0",X"50",X"46",X"4A",X"E0",
		X"50",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"46",X"E0",X"E0",X"BF",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"DB",X"DB",X"DB",X"46",X"E0",X"E0",X"50",X"46",X"4B",X"49",
		X"50",X"0E",X"DB",X"DB",X"DB",X"DB",X"DB",X"46",X"4A",X"E0",X"BF",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"DB",X"12",X"DB",X"46",X"E0",X"E0",X"50",X"46",X"E0",X"E0",
		X"50",X"DB",X"DB",X"DB",X"0C",X"DB",X"DB",X"46",X"4B",X"49",X"BF",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"DB",X"DB",X"DB",X"46",X"E0",X"E0",X"50",X"46",X"E0",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"BF",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"DB",X"DB",X"12",X"46",X"E0",X"E0",X"50",X"46",X"E0",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"BF",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"55",X"51",X"57",X"50",X"DB",X"DB",X"DB",X"46",X"E0",X"E0",X"50",X"46",X"E0",X"E0",
		X"50",X"0D",X"DB",X"DB",X"DB",X"DB",X"DB",X"46",X"E0",X"E0",X"BF",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"56",X"52",X"E0",X"50",X"44",X"DB",X"DB",X"46",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"50",X"DB",X"DB",X"DB",X"DB",X"0F",X"DB",X"46",X"4A",X"E0",X"BF",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"45",X"DB",X"DB",X"46",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"50",X"40",X"DB",X"DB",X"DB",X"DB",X"DB",X"DC",X"4B",X"49",X"BF",X"46",X"4A",X"E0",X"50",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"DB",X"DB",X"DB",X"46",X"E0",X"E0",X"50",X"12",X"DB",X"DB",
		X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"0E",X"46",X"E0",X"E0",X"BF",X"46",X"4B",X"49",X"50",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"DB",X"0D",X"DB",X"46",X"E0",X"E0",X"50",X"DB",X"DB",X"13",
		X"DB",X"DB",X"DB",X"12",X"DB",X"DB",X"DB",X"46",X"E0",X"E0",X"BF",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"DB",X"DB",X"DB",X"46",X"E0",X"E0",X"50",X"DB",X"DB",X"DB",
		X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"46",X"E0",X"E0",X"BF",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"DB",X"DB",X"DB",X"DB",X"46",X"E0",X"E0",X"DB",X"DB",X"DB",X"DB",
		X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"46",X"E0",X"E0",X"DB",X"46",X"E0",X"E0",X"DB",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"DB",X"DB",X"DB",X"DB",X"46",X"E0",X"E0",X"DB",X"DB",X"DB",X"DB",
		X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"46",X"E0",X"E0",X"DB",X"46",X"E0",X"E0",X"DB",X"E0",
		X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",
		X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",
		X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",
		X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"89",X"DB",X"DB",X"DB",X"45",X"DB",X"DB",X"DB",X"DB",X"DB",
		X"DB",X"13",X"DB",X"DB",X"DB",X"DB",X"DB",X"48",X"DB",X"DB",X"DB",X"DB",X"12",X"DB",X"DB",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"88",X"8A",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"0D",X"DB",X"DB",
		X"DB",X"DB",X"DB",X"DB",X"0E",X"DB",X"DB",X"DB",X"13",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"E0",
		X"E0",X"E0",X"81",X"E0",X"88",X"8A",X"E0",X"DB",X"5A",X"DB",X"5A",X"DB",X"5A",X"DB",X"5A",X"DB",
		X"5A",X"DB",X"5A",X"DB",X"5A",X"DB",X"5A",X"DB",X"5A",X"DB",X"5A",X"DB",X"5A",X"DB",X"DB",X"E0",
		X"E0",X"E0",X"82",X"88",X"87",X"8B",X"8C",X"5A",X"5B",X"5A",X"5B",X"5A",X"5B",X"5A",X"5B",X"5A",
		X"5B",X"5A",X"5B",X"5A",X"5B",X"5A",X"5B",X"5A",X"5B",X"5A",X"5B",X"5A",X"5B",X"5A",X"DB",X"E0",
		X"E0",X"E0",X"82",X"86",X"E0",X"8D",X"B2",X"B0",X"B2",X"B0",X"B2",X"B0",X"B2",X"B0",X"B2",X"B0",
		X"B2",X"B0",X"B2",X"B0",X"B2",X"B0",X"B2",X"B0",X"B2",X"B0",X"B2",X"B0",X"B2",X"B0",X"50",X"E0",
		X"E0",X"E0",X"82",X"85",X"E0",X"8F",X"B3",X"B1",X"B3",X"B1",X"B3",X"B1",X"B3",X"B1",X"B3",X"B1",
		X"B3",X"B1",X"B3",X"B1",X"B3",X"B1",X"B3",X"B1",X"B3",X"B1",X"B3",X"B1",X"B3",X"B1",X"50",X"E0",
		X"E0",X"E0",X"82",X"84",X"84",X"8E",X"B2",X"B0",X"B2",X"B0",X"B2",X"B0",X"B2",X"B0",X"B2",X"B0",
		X"B2",X"B0",X"B2",X"B0",X"B2",X"B0",X"B2",X"B0",X"B2",X"B0",X"B2",X"B0",X"B2",X"B0",X"50",X"E0",
		X"E0",X"E0",X"83",X"E0",X"E0",X"8F",X"B3",X"B1",X"B3",X"B1",X"B3",X"B1",X"B3",X"B1",X"B3",X"B1",
		X"B3",X"B1",X"B3",X"B1",X"B3",X"B1",X"B3",X"B1",X"B3",X"B1",X"B3",X"B1",X"B3",X"B1",X"50",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"5B",X"46",X"E0",X"E0",X"5A",X"5B",X"46",X"E0",X"E0",
		X"5A",X"5B",X"46",X"E0",X"E0",X"5A",X"5B",X"5A",X"5B",X"5A",X"5B",X"46",X"4A",X"E0",X"50",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"46",X"4A",X"E0",X"5B",X"DB",X"46",X"E0",X"E0",
		X"5B",X"DB",X"46",X"4A",X"E0",X"5B",X"DB",X"5B",X"DB",X"5B",X"DB",X"46",X"4B",X"49",X"50",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"46",X"4B",X"49",X"50",X"DB",X"46",X"4A",X"E0",
		X"50",X"12",X"46",X"4B",X"49",X"50",X"40",X"DB",X"DB",X"DB",X"DB",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"46",X"E0",X"E0",X"50",X"DB",X"46",X"4B",X"49",
		X"50",X"DB",X"46",X"E0",X"E0",X"50",X"DB",X"DB",X"DB",X"DB",X"DB",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"C0",X"DB",X"46",X"E0",X"E0",X"50",X"0C",X"46",X"E0",X"E0",
		X"50",X"DB",X"46",X"E0",X"E0",X"50",X"0F",X"DB",X"DB",X"DB",X"DB",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"C1",X"DB",X"46",X"E0",X"E0",X"50",X"DB",X"46",X"E0",X"E0",
		X"50",X"DB",X"46",X"DB",X"DB",X"50",X"DB",X"DB",X"DB",X"44",X"DB",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"C2",X"44",X"46",X"E0",X"E0",X"50",X"0D",X"46",X"E0",X"E0",
		X"50",X"DB",X"46",X"E0",X"E0",X"50",X"DB",X"DB",X"DB",X"45",X"DB",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"C3",X"45",X"46",X"E0",X"E0",X"50",X"DB",X"46",X"E0",X"E0",
		X"50",X"0D",X"46",X"E0",X"E0",X"50",X"DB",X"DB",X"13",X"DB",X"DB",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"C4",X"F8",X"DB",X"46",X"4A",X"E0",X"50",X"40",X"46",X"E0",X"E0",
		X"50",X"DB",X"46",X"E0",X"DF",X"FB",X"FE",X"FE",X"FE",X"DB",X"DB",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"C5",X"DB",X"DB",X"46",X"4B",X"49",X"50",X"DB",X"46",X"4A",X"E0",
		X"50",X"DB",X"46",X"E0",X"FF",X"FF",X"FF",X"FF",X"FF",X"DB",X"DB",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"C6",X"DB",X"12",X"46",X"E0",X"E0",X"50",X"12",X"46",X"4B",X"49",
		X"50",X"DB",X"46",X"E5",X"FD",X"FD",X"FC",X"DE",X"DE",X"DB",X"DB",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"C7",X"46",X"E4",X"F9",X"DF",X"DF",X"FB",X"FE",X"F9",X"DF",X"DF",
		X"50",X"DB",X"DB",X"0F",X"DB",X"DB",X"46",X"E0",X"E0",X"DB",X"0E",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"46",X"E0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"50",X"DB",X"DB",X"46",X"E4",X"FE",X"F9",X"DF",X"DF",X"DB",X"DB",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"46",X"E0",X"DE",X"FA",X"FD",X"FD",X"FD",X"FC",X"DE",X"DE",
		X"50",X"12",X"DB",X"46",X"E0",X"FF",X"FF",X"FF",X"FF",X"DB",X"DB",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"46",X"E0",X"E0",X"DB",X"DB",X"DB",X"13",X"46",X"4A",X"E0",
		X"50",X"46",X"DB",X"46",X"E0",X"DE",X"FA",X"FD",X"FD",X"DB",X"DB",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"46",X"E0",X"E0",X"DB",X"12",X"DB",X"DB",X"46",X"4B",X"49",
		X"50",X"46",X"E0",X"E0",X"E0",X"E0",X"DB",X"5A",X"DB",X"0D",X"DB",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"46",X"E0",X"DF",X"FB",X"FE",X"FE",X"FE",X"F9",X"DF",X"DF",
		X"50",X"46",X"E0",X"E0",X"E0",X"E0",X"5A",X"5B",X"DB",X"DB",X"DB",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"46",X"E0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"50",X"46",X"E0",X"E0",X"E0",X"E0",X"5B",X"5A",X"DB",X"DB",X"13",X"46",X"4A",X"E0",X"50",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"46",X"E5",X"FD",X"FD",X"FD",X"FD",X"FD",X"FC",X"DE",X"DE",
		X"50",X"46",X"E0",X"E0",X"E0",X"E0",X"5A",X"5B",X"DB",X"DB",X"DB",X"46",X"4B",X"49",X"50",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"DB",X"DB",X"44",X"DB",X"DB",X"DB",X"DB",X"46",X"E0",X"E0",
		X"50",X"46",X"5B",X"5A",X"5B",X"5A",X"5B",X"DB",X"DB",X"44",X"DB",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"E0",X"E0",
		X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"E0",X"E0",X"E0",X"DB",X"DB",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"E0",X"E0",
		X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"E0",X"E0",X"DB",X"DB",
		X"0A",X"00",X"00",X"0A",X"0A",X"00",X"00",X"0A",X"0E",X"00",X"00",X"0A",X"0F",X"00",X"00",X"0A",
		X"10",X"00",X"00",X"0A",X"11",X"00",X"00",X"0A",X"10",X"00",X"00",X"0A",X"11",X"00",X"00",X"0A",
		X"0A",X"00",X"00",X"0A",X"0A",X"00",X"00",X"0A",X"0E",X"00",X"00",X"0A",X"0F",X"00",X"00",X"0A",
		X"10",X"00",X"00",X"0A",X"11",X"00",X"00",X"0A",X"10",X"00",X"00",X"0A",X"11",X"00",X"00",X"0A",
		X"0A",X"1D",X"1A",X"0A",X"0A",X"1D",X"1A",X"0A",X"0E",X"22",X"1D",X"0A",X"0F",X"00",X"00",X"0A",
		X"10",X"22",X"1D",X"0A",X"11",X"00",X"00",X"0A",X"10",X"22",X"1D",X"0A",X"11",X"22",X"1D",X"0A",
		X"05",X"21",X"1D",X"0A",X"05",X"24",X"21",X"0A",X"09",X"00",X"00",X"0A",X"0A",X"24",X"21",X"0A",
		X"0B",X"00",X"00",X"0A",X"0C",X"00",X"00",X"0A",X"0B",X"00",X"00",X"0A",X"0C",X"00",X"00",X"0A",
		X"05",X"1D",X"18",X"0A",X"05",X"1D",X"18",X"0A",X"09",X"24",X"21",X"0A",X"0A",X"00",X"00",X"0A",
		X"0B",X"24",X"21",X"0A",X"0C",X"00",X"00",X"0A",X"0B",X"24",X"21",X"0A",X"0C",X"00",X"00",X"0A",
		X"0A",X"22",X"1D",X"0A",X"0A",X"26",X"22",X"0A",X"0E",X"00",X"00",X"0A",X"0F",X"26",X"22",X"0A",
		X"10",X"00",X"00",X"0A",X"11",X"00",X"00",X"0A",X"10",X"00",X"00",X"0A",X"11",X"00",X"00",X"0A",
		X"0A",X"22",X"1D",X"0A",X"0A",X"22",X"1D",X"0A",X"0E",X"26",X"22",X"0A",X"0F",X"00",X"00",X"0A",
		X"10",X"26",X"22",X"0A",X"11",X"00",X"00",X"0A",X"10",X"26",X"22",X"0A",X"11",X"26",X"22",X"0A",
		X"03",X"27",X"22",X"0A",X"03",X"2B",X"27",X"0A",X"07",X"00",X"00",X"0A",X"08",X"2B",X"27",X"0A",
		X"09",X"00",X"00",X"0A",X"0A",X"00",X"00",X"0A",X"09",X"00",X"00",X"0A",X"0A",X"2B",X"27",X"0A",
		X"05",X"29",X"24",X"0A",X"05",X"00",X"00",X"0A",X"09",X"29",X"24",X"0A",X"0A",X"29",X"24",X"0A",
		X"0B",X"27",X"21",X"0A",X"0C",X"21",X"1D",X"0A",X"0B",X"00",X"00",X"0A",X"0C",X"22",X"1D",X"0A",
		X"0A",X"00",X"00",X"0A",X"0A",X"00",X"00",X"0A",X"0E",X"00",X"00",X"0A",X"0F",X"00",X"00",X"0A",
		X"10",X"00",X"00",X"0A",X"11",X"00",X"00",X"0A",X"10",X"00",X"00",X"0A",X"11",X"00",X"00",X"0A",
		X"0A",X"00",X"00",X"0A",X"0A",X"00",X"00",X"0A",X"0E",X"00",X"00",X"0A",X"0F",X"00",X"00",X"0A",
		X"10",X"00",X"00",X"0A",X"11",X"00",X"00",X"0A",X"10",X"00",X"00",X"0A",X"11",X"00",X"00",X"0A",
		X"0A",X"1D",X"05",X"0A",X"0A",X"1D",X"05",X"0A",X"0E",X"22",X"0A",X"0A",X"0F",X"00",X"0A",X"0A",
		X"10",X"22",X"0A",X"0A",X"11",X"00",X"0A",X"0A",X"10",X"22",X"0A",X"0A",X"11",X"22",X"0A",X"0A",
		X"05",X"21",X"0C",X"0A",X"05",X"24",X"0C",X"0A",X"09",X"00",X"05",X"0A",X"0A",X"24",X"05",X"0A",
		X"0B",X"00",X"05",X"0A",X"0C",X"00",X"05",X"0A",X"0B",X"00",X"05",X"0A",X"0C",X"00",X"05",X"0A",
		X"05",X"1D",X"0C",X"0A",X"05",X"1D",X"0C",X"0A",X"09",X"24",X"05",X"0A",X"0A",X"00",X"05",X"0A",
		X"0B",X"24",X"05",X"0A",X"0C",X"00",X"05",X"0A",X"0B",X"24",X"05",X"0A",X"0C",X"00",X"05",X"0A",
		X"0A",X"22",X"05",X"0A",X"0A",X"26",X"05",X"0A",X"0E",X"00",X"0A",X"0A",X"0F",X"26",X"0A",X"0A",
		X"10",X"00",X"0A",X"0A",X"11",X"00",X"0A",X"0A",X"10",X"00",X"0A",X"0A",X"11",X"00",X"0A",X"0A",
		X"0A",X"22",X"05",X"0A",X"0A",X"22",X"05",X"0A",X"0E",X"26",X"0A",X"0A",X"0F",X"00",X"0A",X"0A",
		X"10",X"26",X"0A",X"0A",X"11",X"00",X"0A",X"0A",X"10",X"26",X"0A",X"0A",X"11",X"26",X"0A",X"0A",
		X"03",X"27",X"0A",X"0A",X"03",X"2B",X"0A",X"0A",X"07",X"00",X"03",X"0A",X"08",X"2B",X"03",X"0A",
		X"09",X"00",X"03",X"0A",X"0A",X"00",X"03",X"0A",X"09",X"00",X"03",X"0A",X"0A",X"2B",X"03",X"0A",
		X"05",X"29",X"0C",X"0A",X"05",X"00",X"0C",X"0A",X"09",X"29",X"05",X"0A",X"0A",X"29",X"05",X"0A",
		X"0B",X"27",X"05",X"0A",X"0C",X"21",X"05",X"0A",X"0B",X"00",X"05",X"0A",X"0C",X"22",X"05",X"0A",
		X"0A",X"00",X"00",X"0A",X"0A",X"00",X"00",X"0A",X"0E",X"00",X"00",X"0A",X"0F",X"00",X"00",X"0A",
		X"10",X"00",X"00",X"0A",X"11",X"00",X"00",X"0A",X"10",X"00",X"00",X"0A",X"11",X"00",X"00",X"0A",
		X"0A",X"00",X"00",X"0A",X"0A",X"00",X"00",X"0A",X"0E",X"00",X"00",X"0A",X"0F",X"00",X"00",X"0A",
		X"10",X"00",X"00",X"0A",X"11",X"00",X"00",X"0A",X"10",X"00",X"00",X"0A",X"11",X"00",X"00",X"0A",
		X"0A",X"1D",X"05",X"0A",X"0A",X"1D",X"05",X"0A",X"0E",X"22",X"0A",X"0A",X"0F",X"00",X"0A",X"0A",
		X"10",X"22",X"0A",X"0A",X"11",X"00",X"0A",X"0A",X"10",X"22",X"0A",X"0A",X"11",X"22",X"0A",X"0A",
		X"05",X"21",X"0C",X"0A",X"05",X"24",X"0C",X"0A",X"09",X"00",X"05",X"0A",X"0A",X"24",X"05",X"0A",
		X"0B",X"00",X"05",X"0A",X"0C",X"00",X"05",X"0A",X"0B",X"00",X"05",X"0A",X"0C",X"00",X"05",X"0A",
		X"05",X"1D",X"0C",X"0A",X"05",X"1D",X"0C",X"0A",X"09",X"24",X"05",X"0A",X"0A",X"00",X"05",X"0A",
		X"0B",X"24",X"05",X"0A",X"0C",X"00",X"05",X"0A",X"0B",X"24",X"05",X"0A",X"0C",X"00",X"05",X"0A",
		X"0A",X"22",X"05",X"0A",X"0A",X"26",X"05",X"0A",X"0E",X"00",X"0A",X"0A",X"0F",X"26",X"0A",X"0A",
		X"10",X"00",X"0A",X"0A",X"11",X"00",X"0A",X"0A",X"10",X"00",X"0A",X"0A",X"11",X"00",X"0A",X"0A",
		X"0A",X"22",X"05",X"0A",X"0A",X"22",X"05",X"0A",X"0E",X"26",X"0A",X"0A",X"0F",X"00",X"0A",X"0A",
		X"10",X"26",X"0A",X"0A",X"11",X"00",X"0A",X"0A",X"10",X"26",X"0A",X"0A",X"11",X"26",X"0A",X"0A",
		X"03",X"27",X"0A",X"0A",X"03",X"2B",X"0A",X"0A",X"07",X"00",X"03",X"0A",X"08",X"2B",X"03",X"0A",
		X"09",X"00",X"03",X"0A",X"0A",X"00",X"03",X"0A",X"09",X"00",X"03",X"0A",X"0A",X"2B",X"03",X"0A",
		X"05",X"29",X"0C",X"0A",X"05",X"00",X"0C",X"0A",X"09",X"29",X"05",X"0A",X"0A",X"29",X"05",X"0A",
		X"0B",X"27",X"05",X"0A",X"0C",X"21",X"05",X"0A",X"0B",X"00",X"05",X"0A",X"0C",X"22",X"05",X"0A",
		X"0A",X"00",X"05",X"0A",X"00",X"00",X"00",X"FF",X"00",X"00",X"1D",X"0A",X"00",X"00",X"00",X"0A",
		X"00",X"00",X"22",X"0A",X"00",X"00",X"00",X"0A",X"0A",X"05",X"26",X"0A",X"11",X"0A",X"00",X"0A",
		X"13",X"0A",X"00",X"0A",X"11",X"0A",X"00",X"0A",X"0A",X"05",X"26",X"0A",X"11",X"0A",X"00",X"0A",
		X"13",X"0A",X"00",X"0A",X"11",X"0A",X"00",X"0A",X"0A",X"05",X"26",X"0A",X"11",X"0A",X"00",X"0A",
		X"13",X"0A",X"00",X"0A",X"11",X"01",X"24",X"0A",X"0A",X"05",X"00",X"0A",X"11",X"0A",X"26",X"0A",
		X"13",X"0A",X"24",X"0A",X"11",X"0A",X"26",X"0A",X"0A",X"05",X"24",X"0A",X"11",X"0A",X"22",X"0A",
		X"13",X"0A",X"00",X"0A",X"11",X"0A",X"00",X"0A",X"0A",X"05",X"00",X"0A",X"11",X"0A",X"00",X"0A",
		X"13",X"0A",X"00",X"0A",X"11",X"0A",X"00",X"0A",X"0A",X"05",X"00",X"0A",X"11",X"0A",X"00",X"0A",
		X"13",X"0A",X"00",X"0A",X"11",X"0A",X"00",X"0A",X"0A",X"05",X"1D",X"0A",X"11",X"0A",X"00",X"0A",
		X"13",X"0A",X"22",X"0A",X"11",X"0A",X"00",X"0A",X"0A",X"05",X"26",X"0A",X"11",X"0A",X"00",X"0A",
		X"13",X"0A",X"00",X"0A",X"11",X"0A",X"00",X"0A",X"0A",X"05",X"22",X"0A",X"11",X"0A",X"00",X"0A",
		X"13",X"0A",X"26",X"0A",X"11",X"0A",X"00",X"0A",X"0A",X"05",X"29",X"0A",X"11",X"0A",X"00",X"0A",
		X"13",X"0A",X"00",X"0A",X"11",X"0A",X"2B",X"0A",X"0A",X"05",X"00",X"0A",X"11",X"0A",X"29",X"0A",
		X"13",X"0A",X"27",X"0A",X"11",X"0A",X"26",X"0A",X"05",X"0C",X"24",X"0A",X"0C",X"05",X"00",X"0A",
		X"0E",X"05",X"00",X"0A",X"0C",X"05",X"00",X"0A",X"05",X"0C",X"00",X"0A",X"0C",X"05",X"00",X"0A",
		X"0E",X"05",X"00",X"0A",X"0C",X"05",X"00",X"0A",X"0C",X"05",X"00",X"0A",X"0C",X"05",X"00",X"0A",
		X"0E",X"05",X"00",X"0A",X"0C",X"05",X"00",X"0A",X"05",X"0C",X"29",X"0A",X"0C",X"05",X"00",X"0A",
		X"0E",X"05",X"27",X"0A",X"0C",X"05",X"00",X"0A",X"0A",X"05",X"26",X"0A",X"11",X"0A",X"00",X"0A",
		X"13",X"0A",X"00",X"0A",X"11",X"0A",X"00",X"0A",X"0A",X"05",X"26",X"0A",X"11",X"0A",X"00",X"0A",
		X"13",X"0A",X"24",X"0A",X"11",X"0A",X"00",X"0A",X"0A",X"05",X"22",X"0A",X"11",X"0A",X"00",X"0A",
		X"13",X"0A",X"00",X"0A",X"11",X"0A",X"24",X"0A",X"0A",X"05",X"00",X"0A",X"11",X"0A",X"26",X"0A",
		X"13",X"0A",X"00",X"0A",X"11",X"0A",X"29",X"0A",X"03",X"0A",X"00",X"0A",X"0A",X"03",X"27",X"0A",
		X"0C",X"03",X"00",X"0A",X"0A",X"03",X"00",X"0A",X"03",X"0A",X"00",X"0A",X"0A",X"03",X"00",X"0A",
		X"0C",X"03",X"00",X"0A",X"0A",X"03",X"00",X"0A",X"03",X"0A",X"00",X"0A",X"0A",X"03",X"00",X"0A",
		X"0C",X"03",X"00",X"0A",X"0A",X"03",X"00",X"0A",X"03",X"0A",X"21",X"0A",X"0A",X"03",X"00",X"0A",
		X"0C",X"03",X"1F",X"0A",X"0A",X"03",X"00",X"0A",X"0A",X"05",X"1D",X"0A",X"11",X"0A",X"00",X"0A",
		X"13",X"0A",X"00",X"0A",X"11",X"0A",X"00",X"0A",X"0A",X"05",X"22",X"0A",X"11",X"0A",X"00",X"0A",
		X"13",X"0A",X"26",X"0A",X"11",X"0A",X"00",X"0A",X"05",X"0C",X"24",X"0A",X"0C",X"05",X"00",X"0A",
		X"0E",X"05",X"00",X"0A",X"0C",X"05",X"00",X"0A",X"05",X"0C",X"26",X"0A",X"0C",X"05",X"00",X"0A",
		X"0E",X"05",X"24",X"0A",X"0C",X"05",X"00",X"0A",X"0A",X"05",X"22",X"0A",X"11",X"0A",X"00",X"0A",
		X"13",X"0A",X"00",X"0A",X"11",X"0A",X"00",X"0A",X"0A",X"05",X"00",X"0A",X"11",X"0A",X"00",X"0A",
		X"13",X"0A",X"00",X"0A",X"11",X"0A",X"00",X"0A",X"0A",X"05",X"00",X"0A",X"05",X"0C",X"00",X"0A",
		X"05",X"0C",X"00",X"0A",X"05",X"0C",X"00",X"0A",X"05",X"0C",X"1D",X"0A",X"00",X"00",X"00",X"0A",
		X"00",X"00",X"22",X"0A",X"00",X"00",X"00",X"0A",X"0A",X"05",X"26",X"0A",X"11",X"0A",X"00",X"0A",
		X"13",X"0A",X"00",X"0A",X"11",X"0A",X"00",X"0A",X"0A",X"05",X"26",X"0A",X"11",X"0A",X"00",X"0A",
		X"13",X"0A",X"00",X"0A",X"11",X"0A",X"00",X"0A",X"0A",X"05",X"26",X"0A",X"11",X"0A",X"00",X"0A",
		X"13",X"0A",X"00",X"0A",X"11",X"01",X"24",X"0A",X"0A",X"05",X"00",X"0A",X"11",X"0A",X"26",X"0A",
		X"13",X"0A",X"24",X"0A",X"11",X"0A",X"26",X"0A",X"0A",X"05",X"24",X"0A",X"11",X"0A",X"22",X"0A",
		X"13",X"0A",X"00",X"0A",X"11",X"0A",X"00",X"0A",X"0A",X"05",X"00",X"0A",X"11",X"0A",X"00",X"0A",
		X"13",X"0A",X"00",X"0A",X"11",X"0A",X"00",X"0A",X"0A",X"05",X"00",X"0A",X"11",X"0A",X"00",X"0A",
		X"13",X"0A",X"00",X"0A",X"11",X"0A",X"00",X"0A",X"0A",X"05",X"1D",X"0A",X"11",X"0A",X"00",X"0A",
		X"13",X"0A",X"22",X"0A",X"11",X"0A",X"00",X"0A",X"0A",X"05",X"26",X"0A",X"11",X"0A",X"00",X"0A",
		X"13",X"0A",X"00",X"0A",X"11",X"0A",X"00",X"0A",X"0A",X"05",X"22",X"0A",X"11",X"0A",X"00",X"0A",
		X"13",X"0A",X"26",X"0A",X"11",X"0A",X"00",X"0A",X"0A",X"05",X"29",X"0A",X"11",X"0A",X"00",X"0A",
		X"13",X"0A",X"00",X"0A",X"11",X"0A",X"2B",X"0A",X"0A",X"05",X"00",X"0A",X"11",X"0A",X"29",X"0A",
		X"13",X"0A",X"27",X"0A",X"11",X"0A",X"26",X"0A",X"05",X"0C",X"24",X"0A",X"0C",X"05",X"00",X"0A",
		X"0E",X"05",X"00",X"0A",X"0C",X"05",X"00",X"0A",X"05",X"0C",X"00",X"0A",X"0C",X"05",X"00",X"0A",
		X"0E",X"05",X"00",X"0A",X"0C",X"05",X"00",X"0A",X"0C",X"05",X"00",X"0A",X"0C",X"05",X"00",X"0A",
		X"0E",X"05",X"00",X"0A",X"0C",X"05",X"00",X"0A",X"05",X"0C",X"29",X"0A",X"0C",X"05",X"00",X"0A",
		X"0E",X"05",X"27",X"0A",X"0C",X"05",X"00",X"0A",X"0A",X"05",X"26",X"0A",X"11",X"0A",X"00",X"0A",
		X"13",X"0A",X"00",X"0A",X"11",X"0A",X"00",X"0A",X"0A",X"05",X"26",X"0A",X"11",X"0A",X"00",X"0A",
		X"13",X"0A",X"24",X"0A",X"11",X"0A",X"00",X"0A",X"0A",X"05",X"22",X"0A",X"11",X"0A",X"00",X"0A",
		X"13",X"0A",X"00",X"0A",X"11",X"0A",X"24",X"0A",X"0A",X"05",X"00",X"0A",X"11",X"0A",X"26",X"0A",
		X"13",X"0A",X"00",X"0A",X"11",X"0A",X"29",X"0A",X"03",X"0A",X"00",X"0A",X"0A",X"03",X"27",X"0A",
		X"0C",X"03",X"00",X"0A",X"0A",X"03",X"00",X"0A",X"03",X"0A",X"00",X"0A",X"0A",X"03",X"00",X"0A",
		X"0C",X"03",X"00",X"0A",X"0A",X"03",X"00",X"0A",X"03",X"0A",X"00",X"0A",X"0A",X"03",X"00",X"0A",
		X"0C",X"03",X"00",X"0A",X"0A",X"03",X"00",X"0A",X"03",X"0A",X"21",X"0A",X"0A",X"03",X"00",X"0A",
		X"0C",X"03",X"1F",X"0A",X"0A",X"03",X"00",X"0A",X"0A",X"05",X"1D",X"0A",X"11",X"0A",X"00",X"0A",
		X"13",X"0A",X"00",X"0A",X"11",X"0A",X"00",X"0A",X"0A",X"05",X"21",X"0A",X"11",X"0A",X"00",X"0A",
		X"13",X"0A",X"22",X"0A",X"11",X"0A",X"00",X"0A",X"05",X"0C",X"24",X"0A",X"0C",X"05",X"00",X"0A",
		X"0E",X"05",X"00",X"0A",X"0C",X"05",X"00",X"0A",X"05",X"0C",X"26",X"0A",X"0C",X"05",X"00",X"0A",
		X"0E",X"05",X"24",X"0A",X"0C",X"05",X"00",X"0A",X"0A",X"05",X"22",X"0A",X"11",X"0A",X"00",X"0A",
		X"13",X"0A",X"00",X"0A",X"11",X"0A",X"00",X"0A",X"0A",X"05",X"00",X"0A",X"11",X"0A",X"00",X"0A",
		X"13",X"0A",X"00",X"0A",X"11",X"0A",X"00",X"0A",X"0A",X"05",X"00",X"0A",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"1D",X"0A",X"1A",X"1D",X"22",X"14",X"1A",X"1D",X"22",X"1E",X"1A",X"1D",X"22",X"0A",
		X"1A",X"1D",X"26",X"14",X"21",X"1D",X"24",X"14",X"22",X"1F",X"1B",X"1E",X"21",X"1D",X"24",X"0A",
		X"21",X"1D",X"26",X"14",X"21",X"1D",X"24",X"0A",X"1A",X"1D",X"22",X"0A",X"1A",X"1D",X"22",X"1E",
		X"1A",X"1D",X"26",X"0A",X"1A",X"1D",X"29",X"14",X"22",X"27",X"2B",X"14",X"22",X"27",X"2B",X"3C",
		X"26",X"22",X"29",X"14",X"22",X"1D",X"26",X"1E",X"22",X"1D",X"26",X"0A",X"1D",X"1A",X"22",X"14",
		X"21",X"1D",X"24",X"14",X"1F",X"1A",X"22",X"1E",X"21",X"1D",X"24",X"0A",X"21",X"1D",X"26",X"14",
		X"21",X"1D",X"24",X"0A",X"1F",X"1A",X"22",X"0A",X"1A",X"16",X"1F",X"1E",X"1B",X"16",X"1F",X"0A",
		X"18",X"15",X"1D",X"14",X"1D",X"1A",X"22",X"14",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"15",X"FE",X"FE",X"FE",X"40",
		X"FE",X"FE",X"FE",X"01",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"DB",X"46",X"E0",X"E0",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",
		X"DB",X"DB",X"E0",X"E0",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"46",X"E0",X"E0",X"DB",X"DB",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"DB",X"46",X"E0",X"E0",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",
		X"DB",X"DB",X"E0",X"DF",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"46",X"E0",X"E0",X"DB",X"DB",X"E0",
		X"E0",X"E0",X"82",X"E0",X"E0",X"50",X"46",X"E0",X"E0",X"50",X"DB",X"40",X"DB",X"DB",X"DB",X"DB",
		X"DB",X"46",X"E0",X"E0",X"50",X"5B",X"5A",X"5B",X"DB",X"DB",X"46",X"4A",X"E0",X"50",X"DB",X"E0",
		X"E0",X"E0",X"82",X"E0",X"E0",X"50",X"46",X"E0",X"E0",X"50",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",
		X"DB",X"46",X"E0",X"E0",X"50",X"5A",X"5B",X"5A",X"DB",X"DB",X"46",X"4B",X"49",X"50",X"DB",X"E0",
		X"E0",X"E0",X"82",X"E0",X"DF",X"FB",X"F9",X"DF",X"DF",X"50",X"DB",X"DB",X"DB",X"5A",X"46",X"E4",
		X"FE",X"F9",X"DF",X"DF",X"50",X"5B",X"5A",X"5B",X"DB",X"DB",X"46",X"E0",X"E0",X"50",X"DB",X"E0",
		X"C0",X"E0",X"82",X"E0",X"FF",X"FF",X"FF",X"FF",X"FF",X"50",X"0F",X"DB",X"5A",X"5B",X"46",X"E0",
		X"FF",X"FF",X"FF",X"FF",X"50",X"DB",X"5B",X"12",X"DB",X"DB",X"46",X"E0",X"E0",X"50",X"DB",X"E0",
		X"E0",X"E0",X"82",X"E0",X"DE",X"FA",X"FC",X"DE",X"DE",X"50",X"DB",X"DB",X"5B",X"5A",X"46",X"E0",
		X"DE",X"FA",X"DE",X"DE",X"50",X"DB",X"DB",X"DB",X"DB",X"DB",X"46",X"E0",X"E0",X"50",X"DB",X"E0",
		X"E0",X"E0",X"82",X"4A",X"E0",X"50",X"46",X"E9",X"E9",X"50",X"DB",X"DB",X"5A",X"5B",X"46",X"E0",
		X"E0",X"46",X"4A",X"E0",X"50",X"DB",X"DB",X"DB",X"12",X"DB",X"46",X"4A",X"E0",X"50",X"DB",X"E0",
		X"E0",X"E0",X"83",X"4B",X"49",X"50",X"46",X"E9",X"E9",X"E8",X"DB",X"DB",X"5B",X"5A",X"46",X"E0",
		X"E0",X"46",X"4B",X"49",X"50",X"0D",X"DB",X"DB",X"DB",X"DB",X"46",X"4B",X"49",X"50",X"DB",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"EC",X"F0",X"E9",X"E9",X"C9",X"DB",X"5A",X"5B",X"46",X"E0",
		X"E0",X"46",X"E0",X"DF",X"FB",X"FE",X"FE",X"FE",X"FE",X"FE",X"F9",X"DF",X"DF",X"50",X"DB",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"DB",X"F1",X"E9",X"E9",X"C9",X"DA",X"5B",X"5A",X"46",X"E0",
		X"E0",X"46",X"E0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"50",X"DB",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"DB",X"EC",X"F0",X"E9",X"E9",X"C9",X"DB",X"5B",X"46",X"E0",
		X"E0",X"46",X"4A",X"DE",X"FA",X"FD",X"FC",X"DE",X"DE",X"FA",X"FC",X"DE",X"DE",X"50",X"DB",X"E0",
		X"E0",X"E0",X"55",X"51",X"57",X"50",X"DB",X"DB",X"F1",X"E9",X"E9",X"C9",X"DA",X"5A",X"46",X"E0",
		X"E0",X"46",X"4B",X"49",X"DB",X"DB",X"46",X"4B",X"49",X"50",X"46",X"4A",X"E0",X"50",X"DB",X"E0",
		X"E0",X"E0",X"56",X"52",X"E0",X"50",X"DB",X"41",X"EC",X"F0",X"E9",X"E9",X"C9",X"5B",X"46",X"E0",
		X"DF",X"FB",X"DF",X"DF",X"DB",X"12",X"EE",X"E0",X"E0",X"50",X"46",X"4B",X"49",X"50",X"DB",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"0F",X"DB",X"DB",X"F1",X"E9",X"E9",X"C9",X"DA",X"46",X"E0",
		X"FF",X"FF",X"FF",X"FF",X"DB",X"ED",X"EF",X"E0",X"E0",X"50",X"46",X"E0",X"E0",X"50",X"DB",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"DB",X"DB",X"DB",X"EC",X"F0",X"E9",X"E9",X"C9",X"46",X"E5",
		X"FD",X"FD",X"FD",X"FD",X"DB",X"EE",X"E0",X"E0",X"E0",X"50",X"46",X"E0",X"E0",X"50",X"DB",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"DB",X"DB",X"DB",X"DB",X"F1",X"E9",X"E9",X"C9",X"DA",X"DB",
		X"0C",X"DB",X"DB",X"13",X"ED",X"EF",X"E0",X"E0",X"5D",X"DB",X"46",X"E0",X"E0",X"50",X"DB",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"DB",X"DB",X"DB",X"DB",X"EC",X"F0",X"E9",X"E9",X"C9",X"DB",
		X"DB",X"DB",X"DB",X"DB",X"EE",X"E0",X"E0",X"E0",X"5E",X"DB",X"46",X"E0",X"E0",X"50",X"DB",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"DB",X"0D",X"DB",X"DB",X"DB",X"F1",X"E9",X"E9",X"C9",X"DA",
		X"DB",X"DB",X"DB",X"ED",X"EF",X"E0",X"E0",X"5D",X"5C",X"DB",X"46",X"E0",X"E0",X"50",X"DB",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"DB",X"DB",X"DB",X"DB",X"DB",X"EC",X"F0",X"E9",X"E9",X"C9",
		X"DB",X"DB",X"0F",X"EE",X"E0",X"E0",X"E0",X"5E",X"DB",X"DB",X"46",X"E0",X"E0",X"50",X"DB",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"DB",X"DB",X"DB",X"13",X"DB",X"DB",X"F1",X"E9",X"E9",X"C9",
		X"DA",X"DB",X"ED",X"EF",X"E0",X"E0",X"5D",X"5C",X"47",X"DB",X"46",X"E0",X"E0",X"50",X"DB",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"DB",X"DB",X"DB",X"DB",X"DB",X"12",X"EC",X"F0",X"E9",X"E9",
		X"C9",X"0E",X"46",X"E0",X"E0",X"E0",X"5E",X"DB",X"48",X"DB",X"46",X"E0",X"E0",X"50",X"DB",X"E0",
		X"E0",X"E0",X"81",X"4A",X"E0",X"50",X"DB",X"DB",X"0D",X"44",X"DB",X"DB",X"DB",X"F1",X"E9",X"E9",
		X"C9",X"DA",X"46",X"4A",X"E0",X"5D",X"5C",X"DB",X"DB",X"13",X"46",X"4A",X"E0",X"50",X"DB",X"E0",
		X"E0",X"E0",X"82",X"4B",X"49",X"50",X"0F",X"DB",X"DB",X"45",X"DB",X"DB",X"DB",X"46",X"E9",X"E9",
		X"E7",X"DB",X"46",X"4B",X"49",X"5E",X"0E",X"DB",X"DB",X"DB",X"46",X"4B",X"49",X"50",X"DB",X"E0",
		X"E0",X"E0",X"82",X"E0",X"DF",X"FB",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"F9",X"DF",X"DF",
		X"FB",X"FE",X"F9",X"DF",X"DF",X"FB",X"FE",X"FE",X"FE",X"FE",X"F9",X"DF",X"DF",X"50",X"DB",X"E0",
		X"E0",X"E0",X"82",X"E0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"50",X"DB",X"E0",
		X"E0",X"E0",X"82",X"E0",X"DE",X"FA",X"FC",X"DE",X"DE",X"FA",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",
		X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FC",X"DE",X"DE",X"50",X"DB",X"E0",
		X"E0",X"E0",X"82",X"4A",X"E0",X"50",X"46",X"E0",X"E0",X"50",X"DB",X"40",X"DB",X"DB",X"13",X"DB",
		X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"12",X"DB",X"46",X"E0",X"E0",X"50",X"DB",X"E0",
		X"E0",X"E0",X"83",X"4B",X"49",X"50",X"46",X"E0",X"E0",X"50",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",
		X"DB",X"0D",X"DB",X"41",X"DB",X"DB",X"DB",X"DB",X"DB",X"0F",X"46",X"E0",X"E0",X"50",X"DB",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"12",X"DB",X"DB",X"DB",
		X"DB",X"DB",X"DB",X"DB",X"DB",X"12",X"DB",X"DB",X"DB",X"DB",X"46",X"DB",X"DB",X"DB",X"13",X"E0",
		X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",
		X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"E0",
		X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",
		X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"DB",X"DB",X"DB",X"46",X"E0",X"E0",X"50",X"DB",X"DB",X"DB",
		X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"DB",X"DB",X"DB",X"46",X"E0",X"E0",X"50",X"DB",X"DB",X"DB",
		X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"46",X"DB",X"DB",X"DB",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"DB",X"DB",X"DB",X"46",X"E0",X"E0",X"50",X"DB",X"45",X"DB",
		X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"0F",X"DB",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"DB",X"DB",X"0D",X"46",X"4A",X"E0",X"50",X"DB",X"DB",X"DB",
		X"DB",X"DB",X"DB",X"12",X"DB",X"DB",X"DB",X"46",X"E4",X"FE",X"FE",X"F9",X"DF",X"DF",X"50",X"E0",
		X"E0",X"E0",X"81",X"4A",X"E0",X"50",X"DB",X"DB",X"DB",X"46",X"4B",X"49",X"50",X"0C",X"DB",X"DB",
		X"DB",X"DB",X"DB",X"DB",X"41",X"DB",X"DB",X"46",X"E0",X"FF",X"FF",X"FF",X"FF",X"FF",X"50",X"E0",
		X"E0",X"E0",X"82",X"4B",X"49",X"50",X"0D",X"DB",X"DB",X"46",X"E0",X"E0",X"50",X"DB",X"DB",X"DB",
		X"0F",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"46",X"E0",X"DE",X"FA",X"FC",X"DE",X"DE",X"50",X"E0",
		X"E0",X"E0",X"82",X"E0",X"DF",X"FB",X"FE",X"FE",X"FE",X"F9",X"DF",X"DF",X"FB",X"FE",X"FE",X"FE",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"F9",X"DF",X"DF",X"50",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"82",X"E0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"50",X"46",X"4A",X"E0",X"50",X"E0",
		X"E0",X"E0",X"82",X"E0",X"DE",X"FA",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FC",X"DE",X"DE",X"FA",
		X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FC",X"DE",X"DE",X"50",X"46",X"4B",X"49",X"50",X"E0",
		X"E0",X"E0",X"82",X"4A",X"E0",X"50",X"DB",X"DB",X"12",X"DB",X"DB",X"40",X"46",X"4A",X"E0",X"5A",
		X"DB",X"DB",X"5A",X"5A",X"DB",X"DB",X"DB",X"46",X"4A",X"E0",X"50",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"83",X"4B",X"49",X"50",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"46",X"4B",X"49",X"5B",
		X"5A",X"5A",X"5B",X"5B",X"5A",X"DB",X"DB",X"46",X"4B",X"49",X"50",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"12",X"DB",X"DB",X"DB",X"DB",X"DB",X"46",X"E0",X"E0",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"46",X"4A",X"E0",X"50",X"E0",
		X"E0",X"E0",X"55",X"51",X"57",X"50",X"DB",X"DB",X"DB",X"DB",X"0F",X"DB",X"46",X"E0",X"E0",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"46",X"4B",X"49",X"50",X"E0",
		X"E0",X"E0",X"56",X"52",X"E0",X"50",X"44",X"DB",X"DB",X"DB",X"DB",X"DB",X"46",X"E0",X"E0",X"5B",
		X"5A",X"5B",X"5A",X"5B",X"5A",X"5B",X"5A",X"46",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"45",X"DB",X"DB",X"DB",X"DB",X"EA",X"F6",X"E0",X"E0",X"5A",
		X"5B",X"5A",X"5B",X"DB",X"5B",X"5A",X"5B",X"46",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"DB",X"DB",X"12",X"DB",X"EA",X"F6",X"E0",X"E0",X"F7",X"5B",
		X"DB",X"5B",X"DB",X"0E",X"DB",X"5B",X"DB",X"46",X"4A",X"E0",X"50",X"46",X"4A",X"E0",X"50",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"DB",X"DB",X"DB",X"EA",X"F6",X"E0",X"E0",X"F7",X"DB",X"DB",
		X"13",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"46",X"4B",X"49",X"50",X"46",X"4B",X"49",X"50",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"DB",X"DB",X"EA",X"F6",X"E0",X"E0",X"F7",X"46",X"E4",X"FE",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"DB",X"46",X"E0",X"E0",X"50",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"0F",X"EA",X"F6",X"E0",X"E0",X"F7",X"DB",X"46",X"E0",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"50",X"46",X"E0",X"E0",X"50",X"46",X"4A",X"E0",X"50",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"EA",X"F6",X"E0",X"E0",X"F7",X"DB",X"DB",X"46",X"E0",X"DE",
		X"FA",X"FD",X"FD",X"FC",X"DE",X"DE",X"50",X"46",X"E0",X"E0",X"50",X"46",X"4B",X"49",X"50",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"46",X"E0",X"E0",X"F7",X"DB",X"DB",X"DB",X"46",X"E0",X"E0",
		X"50",X"12",X"DB",X"46",X"E0",X"E0",X"50",X"46",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"81",X"4A",X"E0",X"50",X"46",X"4A",X"E0",X"50",X"DB",X"13",X"DB",X"46",X"E0",X"E0",
		X"50",X"DB",X"DB",X"46",X"4A",X"E0",X"50",X"46",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"82",X"4B",X"49",X"50",X"46",X"4B",X"49",X"50",X"40",X"DB",X"DB",X"46",X"E0",X"E0",
		X"50",X"DB",X"DB",X"46",X"4B",X"49",X"50",X"46",X"E0",X"E0",X"50",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"82",X"E0",X"DF",X"FB",X"F9",X"DF",X"DF",X"50",X"DB",X"DB",X"DB",X"46",X"E0",X"E0",
		X"50",X"DB",X"0F",X"46",X"E0",X"E0",X"50",X"46",X"E0",X"E0",X"50",X"46",X"4A",X"E0",X"50",X"E0",
		X"E0",X"E0",X"82",X"E0",X"FF",X"FF",X"FF",X"FF",X"FF",X"50",X"DB",X"46",X"DB",X"46",X"BE",X"BF",
		X"50",X"DB",X"E4",X"F9",X"DF",X"DF",X"FB",X"F9",X"DF",X"DF",X"50",X"46",X"4B",X"49",X"50",X"E0",
		X"E0",X"E0",X"82",X"E0",X"DE",X"FA",X"FC",X"DE",X"DE",X"50",X"DB",X"46",X"FB",X"FB",X"FB",X"5A",
		X"DB",X"46",X"E0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"50",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"82",X"E0",X"E0",X"50",X"46",X"E0",X"E0",X"50",X"DB",X"46",X"FB",X"FB",X"FB",X"5B",
		X"5A",X"46",X"E0",X"DE",X"FA",X"FD",X"FD",X"FD",X"FD",X"FD",X"46",X"E4",X"DF",X"DF",X"50",X"E0",
		X"E0",X"E0",X"82",X"E0",X"E0",X"50",X"46",X"E0",X"E0",X"50",X"DB",X"46",X"FB",X"FB",X"FB",X"5A",
		X"5B",X"46",X"4A",X"E0",X"50",X"12",X"DB",X"DB",X"44",X"DB",X"46",X"E0",X"FF",X"FF",X"50",X"E0",
		X"E0",X"E0",X"82",X"E0",X"E0",X"50",X"46",X"E0",X"E0",X"50",X"12",X"46",X"E0",X"E0",X"E0",X"5B",
		X"5A",X"46",X"4B",X"49",X"50",X"DB",X"DB",X"DB",X"45",X"DB",X"46",X"E0",X"DE",X"FA",X"DB",X"E0",
		X"E0",X"E0",X"82",X"E0",X"E0",X"50",X"46",X"E0",X"E0",X"50",X"DB",X"46",X"5B",X"5A",X"5B",X"5A",
		X"5B",X"46",X"E0",X"E0",X"50",X"DB",X"13",X"DB",X"DB",X"DB",X"46",X"E0",X"E0",X"50",X"DB",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"DB",X"46",X"E0",X"E0",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",
		X"DB",X"46",X"E0",X"E0",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"46",X"E0",X"E0",X"DB",X"DB",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"DB",X"46",X"E0",X"E0",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",
		X"DB",X"46",X"E0",X"E0",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"46",X"E0",X"E0",X"DB",X"DB",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"DB",X"DB",X"DB",X"DB",X"46",X"E0",X"E0",X"DB",X"DB",X"DB",X"DB",
		X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"46",X"E0",X"E0",X"DB",X"46",X"E0",X"E0",X"DB",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"DB",X"DB",X"DB",X"DB",X"46",X"E0",X"E0",X"DB",X"DB",X"DB",X"DB",
		X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"46",X"E0",X"E0",X"DB",X"46",X"E0",X"E0",X"DB",X"E0",
		X"E0",X"E0",X"81",X"4A",X"E0",X"50",X"DB",X"DB",X"13",X"46",X"E0",X"E0",X"50",X"DB",X"12",X"DB",
		X"DB",X"DB",X"DB",X"DB",X"DB",X"13",X"DB",X"46",X"E0",X"E0",X"BF",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"82",X"4B",X"49",X"50",X"0F",X"DB",X"DB",X"46",X"E0",X"E0",X"50",X"DB",X"DB",X"DB",
		X"DB",X"DB",X"0C",X"DB",X"DB",X"DB",X"DB",X"46",X"E0",X"E0",X"BF",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"82",X"E0",X"DF",X"FB",X"FE",X"FE",X"FE",X"F9",X"DF",X"DF",X"FB",X"FE",X"FE",X"FE",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"F9",X"DF",X"DF",X"FB",X"F9",X"DF",X"DF",X"50",X"E0",
		X"E0",X"E0",X"82",X"E0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"50",X"E0",
		X"E0",X"E0",X"82",X"E0",X"DE",X"FA",X"FD",X"FD",X"FD",X"FC",X"DE",X"DE",X"FA",X"FD",X"FD",X"FC",
		X"DE",X"DE",X"FA",X"FD",X"FD",X"FD",X"FD",X"FC",X"DE",X"DE",X"FA",X"FC",X"DE",X"DE",X"50",X"E0",
		X"E0",X"E0",X"82",X"E0",X"E0",X"50",X"DB",X"DB",X"DB",X"46",X"E0",X"E0",X"50",X"DB",X"0D",X"46",
		X"E0",X"E0",X"50",X"DB",X"DB",X"DB",X"DB",X"46",X"4A",X"E0",X"BF",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"82",X"E0",X"E0",X"50",X"DB",X"12",X"DB",X"46",X"4A",X"E0",X"50",X"DB",X"DB",X"46",
		X"E0",X"E0",X"50",X"DB",X"13",X"DB",X"47",X"46",X"4B",X"49",X"BF",X"46",X"4A",X"E0",X"50",X"E0",
		X"E0",X"E0",X"82",X"E0",X"E0",X"50",X"DB",X"DB",X"DB",X"46",X"4B",X"49",X"50",X"DB",X"44",X"46",
		X"4A",X"E0",X"50",X"DB",X"DB",X"DB",X"48",X"46",X"E0",X"E0",X"BF",X"46",X"4B",X"49",X"50",X"E0",
		X"E0",X"E0",X"82",X"E0",X"E0",X"50",X"DB",X"DB",X"12",X"46",X"E0",X"E0",X"50",X"DB",X"45",X"46",
		X"4B",X"49",X"50",X"DB",X"DB",X"DB",X"12",X"46",X"E0",X"E0",X"BF",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"82",X"E0",X"E0",X"50",X"0D",X"DB",X"DB",X"46",X"E0",X"E0",X"50",X"12",X"DB",X"46",
		X"E0",X"E0",X"50",X"DB",X"DB",X"DB",X"DB",X"46",X"4A",X"E0",X"BF",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"82",X"E0",X"DF",X"FB",X"FE",X"FE",X"FE",X"F9",X"DF",X"DF",X"50",X"DB",X"0F",X"46",
		X"E0",X"E0",X"50",X"DB",X"DB",X"DB",X"DB",X"46",X"4B",X"49",X"BF",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"82",X"E0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"50",X"DB",X"12",X"46",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"BF",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"82",X"E0",X"DE",X"FA",X"FD",X"FD",X"FD",X"FC",X"DE",X"DE",X"50",X"DB",X"DB",X"46",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"BF",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"82",X"4A",X"E0",X"50",X"13",X"DB",X"DB",X"46",X"E0",X"E0",X"50",X"DB",X"DB",X"46",
		X"E0",X"E0",X"DB",X"5A",X"DB",X"5A",X"5B",X"46",X"E0",X"E0",X"BF",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"83",X"4B",X"49",X"50",X"DB",X"40",X"DB",X"46",X"E0",X"E0",X"50",X"12",X"EA",X"F6",
		X"E0",X"E0",X"DB",X"5B",X"5A",X"5B",X"5A",X"46",X"4A",X"E0",X"BF",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"DB",X"DB",X"DB",X"46",X"E0",X"E0",X"50",X"EA",X"F6",X"E0",
		X"E0",X"F7",X"3A",X"5A",X"5B",X"5A",X"5B",X"46",X"4B",X"49",X"BF",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"DB",X"DB",X"DB",X"46",X"4A",X"E0",X"EA",X"F6",X"E0",X"E0",
		X"F7",X"DB",X"3B",X"E0",X"E0",X"E0",X"DB",X"46",X"E0",X"E0",X"BF",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"DB",X"DB",X"12",X"46",X"4B",X"49",X"F6",X"E0",X"E0",X"F7",
		X"DB",X"DB",X"3C",X"E0",X"E0",X"E0",X"DB",X"DC",X"E0",X"E0",X"BF",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"DB",X"DB",X"DB",X"46",X"E0",X"E0",X"E0",X"E0",X"F7",X"DB",
		X"DB",X"DB",X"3D",X"E0",X"E0",X"E0",X"DB",X"46",X"E0",X"E0",X"BF",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"DB",X"DB",X"DB",X"46",X"E0",X"E0",X"E0",X"F7",X"DB",X"DB",
		X"DB",X"DB",X"3E",X"E0",X"E0",X"E0",X"DB",X"46",X"E0",X"E0",X"BF",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"DB",X"0D",X"DB",X"46",X"E0",X"E0",X"F7",X"DB",X"12",X"DB",
		X"DB",X"DB",X"3F",X"46",X"4A",X"E0",X"DB",X"46",X"4A",X"E0",X"BF",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"DB",X"DB",X"DB",X"46",X"E0",X"E0",X"DB",X"DB",X"DB",X"DB",
		X"DB",X"0F",X"DB",X"46",X"4B",X"49",X"13",X"46",X"4B",X"49",X"BF",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"DB",X"5A",X"DB",X"46",X"E0",X"DF",X"FB",X"FE",X"FE",X"FE",
		X"FE",X"FE",X"FE",X"F9",X"DF",X"DF",X"FB",X"F9",X"DF",X"DF",X"BF",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"5A",X"5B",X"DB",X"46",X"E0",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"50",X"5B",X"5A",X"DB",X"46",X"E0",X"DE",X"FA",X"FD",X"FD",X"FD",
		X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FC",X"DE",X"DE",X"BF",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"55",X"51",X"57",X"50",X"5A",X"5B",X"DB",X"46",X"E0",X"E0",X"50",X"DB",X"DB",X"DB",
		X"DB",X"DB",X"12",X"DB",X"DB",X"DB",X"0D",X"46",X"E0",X"E0",X"BF",X"46",X"4A",X"E0",X"50",X"E0",
		X"E0",X"E0",X"56",X"52",X"E0",X"5A",X"5B",X"DB",X"DB",X"46",X"E0",X"E0",X"50",X"DB",X"0F",X"DB",
		X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"46",X"E0",X"E0",X"BF",X"46",X"4B",X"49",X"50",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"5B",X"5A",X"DB",X"DB",X"46",X"E0",X"E0",X"50",X"DB",X"DB",X"DB",
		X"DB",X"DB",X"DB",X"DB",X"40",X"DB",X"DB",X"46",X"DB",X"DB",X"DB",X"46",X"E0",X"E0",X"50",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"DB",X"DB",X"DB",X"DB",X"46",X"E0",X"E0",X"DB",X"DB",X"DB",X"DB",
		X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"BF",X"46",X"E0",X"E0",X"DB",X"E0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"DB",X"DB",X"DB",X"DB",X"46",X"E0",X"E0",X"DB",X"DB",X"DB",X"DB",
		X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"DB",X"BF",X"46",X"E0",X"E0",X"DB",X"E0",
		X"FF",X"FE",X"FD",X"FC",X"E5",X"E5",X"EE",X"ED",X"EC",X"E5",X"3F",X"FB",X"FA",X"F9",X"F8",X"F4",
		X"F2",X"F0",X"EB",X"EA",X"E9",X"3F",X"E5",X"F7",X"F6",X"F5",X"F3",X"F1",X"EF",X"E8",X"E7",X"E6",
		X"3F",X"E4",X"E3",X"E2",X"E1",X"E2",X"E0",X"DF",X"E2",X"3F",X"D9",X"D8",X"D7",X"D6",X"D5",X"91",
		X"D4",X"D3",X"91",X"D2",X"D1",X"D0",X"CF",X"CE",X"CD",X"CC",X"CB",X"CA",X"C9",X"C8",X"C7",X"C6",
		X"C5",X"C4",X"C3",X"C2",X"3F",X"C1",X"C0",X"BF",X"BE",X"BD",X"91",X"BC",X"BB",X"BA",X"B9",X"B8",
		X"B7",X"B6",X"B5",X"B4",X"B3",X"B2",X"B1",X"B0",X"AF",X"AE",X"BC",X"AD",X"AC",X"AB",X"AA",X"3F",
		X"A9",X"A8",X"A7",X"A6",X"A5",X"91",X"A4",X"A3",X"A2",X"A1",X"A0",X"9F",X"9E",X"9D",X"9C",X"9B",
		X"9A",X"99",X"98",X"97",X"96",X"95",X"94",X"93",X"B3",X"92",X"3F",X"DE",X"91",X"DD",X"DC",X"DB",
		X"DA",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"8A",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",
		X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"8F",X"3F",X"8C",X"90",X"90",X"90",X"90",
		X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",
		X"90",X"90",X"90",X"90",X"8D",X"3F",X"85",X"84",X"83",X"82",X"81",X"80",X"7F",X"91",X"91",X"3F",
		X"91",X"54",X"89",X"88",X"87",X"86",X"91",X"91",X"91",X"3F",X"7E",X"7D",X"7C",X"7B",X"7A",X"91",
		X"91",X"91",X"91",X"3F",X"79",X"78",X"77",X"76",X"75",X"74",X"91",X"91",X"91",X"3F",X"73",X"72",
		X"71",X"70",X"6F",X"6E",X"6D",X"6C",X"6B",X"3F",X"91",X"91",X"6A",X"69",X"68",X"67",X"66",X"91",
		X"91",X"3F",X"91",X"65",X"64",X"63",X"62",X"91",X"91",X"91",X"91",X"3F",X"61",X"60",X"5F",X"5E",
		X"5D",X"91",X"91",X"91",X"91",X"3F",X"5A",X"59",X"91",X"58",X"57",X"3F",X"5C",X"3F",X"5B",X"3F",
		X"56",X"3F",X"55",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0A",X"00",X"00",X"0A",X"0A",X"00",X"00",X"0A",X"0E",X"00",X"00",X"0A",X"0A",X"00",X"00",X"0A",
		X"11",X"00",X"00",X"0A",X"0A",X"00",X"00",X"0A",X"13",X"00",X"00",X"0A",X"0A",X"00",X"00",X"0A",
		X"14",X"00",X"00",X"0A",X"0A",X"00",X"1C",X"0A",X"13",X"00",X"1D",X"0A",X"0A",X"00",X"00",X"0A",
		X"11",X"00",X"22",X"0A",X"0A",X"00",X"00",X"0A",X"0F",X"00",X"24",X"0A",X"0E",X"09",X"00",X"0A",
		X"0A",X"0A",X"26",X"0A",X"0A",X"16",X"00",X"0A",X"0E",X"0A",X"00",X"0A",X"0A",X"16",X"26",X"0A",
		X"11",X"0A",X"00",X"0A",X"0A",X"16",X"00",X"0A",X"13",X"0A",X"00",X"0A",X"0A",X"16",X"00",X"0A",
		X"14",X"0A",X"00",X"0A",X"0A",X"16",X"26",X"0A",X"13",X"0A",X"00",X"0A",X"0A",X"16",X"26",X"0A",
		X"11",X"0A",X"25",X"0A",X"0A",X"16",X"26",X"0A",X"0F",X"0A",X"00",X"0A",X"0E",X"09",X"00",X"0A",
		X"0A",X"0A",X"22",X"0A",X"0A",X"16",X"00",X"0A",X"0E",X"0A",X"00",X"0A",X"0A",X"16",X"22",X"0A",
		X"11",X"0A",X"00",X"0A",X"0A",X"16",X"00",X"0A",X"13",X"0A",X"00",X"0A",X"0A",X"16",X"00",X"0A",
		X"14",X"0A",X"00",X"0A",X"0A",X"16",X"00",X"0A",X"13",X"0A",X"22",X"0A",X"0A",X"16",X"00",X"0A",
		X"11",X"0A",X"24",X"0A",X"0A",X"16",X"00",X"0A",X"0F",X"0A",X"26",X"0A",X"0E",X"02",X"00",X"0A",
		X"03",X"03",X"27",X"0A",X"03",X"0F",X"00",X"0A",X"07",X"03",X"00",X"0A",X"03",X"0F",X"2B",X"0A",
		X"0A",X"03",X"00",X"0A",X"03",X"0F",X"00",X"0A",X"0C",X"03",X"00",X"0A",X"03",X"0F",X"00",X"0A",
		X"0D",X"03",X"00",X"0A",X"03",X"0F",X"2B",X"0A",X"0C",X"03",X"00",X"0A",X"03",X"0F",X"2B",X"0A",
		X"0A",X"03",X"29",X"0A",X"03",X"0F",X"27",X"0A",X"08",X"03",X"00",X"0A",X"07",X"09",X"00",X"0A",
		X"0A",X"0A",X"26",X"0A",X"0A",X"16",X"00",X"0A",X"0E",X"0A",X"00",X"0A",X"0A",X"16",X"22",X"0A",
		X"11",X"0A",X"00",X"0A",X"0A",X"16",X"00",X"0A",X"13",X"0A",X"00",X"0A",X"0A",X"16",X"00",X"0A",
		X"14",X"0A",X"00",X"0A",X"0A",X"16",X"21",X"0A",X"13",X"0A",X"22",X"0A",X"0A",X"16",X"00",X"0A",
		X"11",X"0A",X"24",X"0A",X"0A",X"16",X"00",X"0A",X"0F",X"0A",X"26",X"0A",X"0E",X"02",X"00",X"0A",
		X"03",X"03",X"27",X"0A",X"03",X"0F",X"00",X"0A",X"07",X"03",X"00",X"0A",X"03",X"0F",X"2B",X"0A",
		X"0A",X"03",X"00",X"0A",X"03",X"0F",X"00",X"0A",X"0C",X"03",X"00",X"0A",X"03",X"0F",X"00",X"0A",
		X"0D",X"03",X"00",X"0A",X"03",X"0F",X"2B",X"0A",X"0C",X"03",X"00",X"0A",X"03",X"0F",X"2B",X"0A",
		X"0A",X"03",X"29",X"0A",X"03",X"0F",X"27",X"0A",X"08",X"03",X"00",X"0A",X"07",X"09",X"00",X"0A",
		X"0A",X"0A",X"26",X"0A",X"0A",X"16",X"00",X"0A",X"0E",X"0A",X"00",X"0A",X"0A",X"16",X"22",X"0A",
		X"11",X"0A",X"00",X"0A",X"0A",X"16",X"00",X"0A",X"13",X"0A",X"00",X"0A",X"0A",X"16",X"00",X"0A",
		X"14",X"0A",X"00",X"0A",X"0A",X"16",X"00",X"0A",X"13",X"0A",X"1D",X"0A",X"0A",X"16",X"00",X"0A",
		X"11",X"0A",X"22",X"0A",X"0A",X"16",X"00",X"0A",X"0F",X"0A",X"24",X"0A",X"0E",X"09",X"00",X"0A",
		X"0A",X"0A",X"26",X"0A",X"0A",X"16",X"00",X"0A",X"0E",X"0A",X"00",X"0A",X"0A",X"16",X"26",X"0A",
		X"11",X"0A",X"00",X"0A",X"0A",X"16",X"00",X"0A",X"0F",X"0A",X"27",X"0A",X"0E",X"04",X"00",X"0A",
		X"05",X"05",X"24",X"0A",X"05",X"11",X"00",X"0A",X"09",X"05",X"24",X"0A",X"05",X"11",X"00",X"0A",
		X"0C",X"05",X"00",X"0A",X"05",X"11",X"26",X"0A",X"0A",X"05",X"00",X"0A",X"09",X"09",X"22",X"0A",
		X"0A",X"0A",X"00",X"0A",X"0A",X"16",X"00",X"0A",X"0E",X"0A",X"00",X"0A",X"0A",X"16",X"00",X"0A",
		X"11",X"0A",X"00",X"0A",X"11",X"16",X"00",X"0A",X"0D",X"0A",X"00",X"0A",X"0E",X"16",X"00",X"0A",
		X"0A",X"0A",X"00",X"0A",X"0A",X"00",X"1C",X"0A",X"13",X"00",X"1D",X"0A",X"0A",X"00",X"00",X"0A",
		X"11",X"00",X"22",X"0A",X"0A",X"00",X"00",X"0A",X"0F",X"00",X"24",X"0A",X"0E",X"09",X"00",X"0A",
		X"0A",X"0A",X"26",X"0A",X"0A",X"16",X"00",X"0A",X"0E",X"0A",X"00",X"0A",X"0A",X"16",X"26",X"0A",
		X"11",X"0A",X"00",X"0A",X"0A",X"16",X"00",X"0A",X"13",X"0A",X"00",X"0A",X"0A",X"16",X"00",X"0A",
		X"14",X"0A",X"00",X"0A",X"0A",X"16",X"26",X"0A",X"13",X"0A",X"00",X"0A",X"0A",X"16",X"26",X"0A",
		X"11",X"0A",X"25",X"0A",X"0A",X"16",X"26",X"0A",X"0F",X"0A",X"00",X"0A",X"0E",X"09",X"00",X"0A",
		X"0A",X"0A",X"22",X"0A",X"0A",X"16",X"00",X"0A",X"0E",X"0A",X"00",X"0A",X"0A",X"16",X"22",X"0A",
		X"11",X"0A",X"00",X"0A",X"0A",X"16",X"00",X"0A",X"13",X"0A",X"00",X"0A",X"0A",X"16",X"00",X"0A",
		X"14",X"0A",X"00",X"0A",X"0A",X"16",X"00",X"0A",X"13",X"0A",X"22",X"0A",X"0A",X"16",X"00",X"0A",
		X"11",X"0A",X"24",X"0A",X"0A",X"16",X"00",X"0A",X"0F",X"0A",X"26",X"0A",X"0E",X"02",X"00",X"0A",
		X"03",X"03",X"27",X"0A",X"03",X"0F",X"00",X"0A",X"07",X"03",X"00",X"0A",X"03",X"0F",X"2B",X"0A",
		X"0A",X"03",X"00",X"0A",X"03",X"0F",X"00",X"0A",X"0C",X"03",X"00",X"0A",X"03",X"0F",X"00",X"0A",
		X"0D",X"03",X"00",X"0A",X"03",X"0F",X"2B",X"0A",X"0C",X"03",X"00",X"0A",X"03",X"0F",X"2B",X"0A",
		X"0A",X"03",X"29",X"0A",X"03",X"0F",X"27",X"0A",X"08",X"03",X"00",X"0A",X"07",X"09",X"00",X"0A",
		X"0A",X"0A",X"26",X"0A",X"0A",X"16",X"00",X"0A",X"0E",X"0A",X"00",X"0A",X"0A",X"16",X"22",X"0A",
		X"11",X"0A",X"00",X"0A",X"0A",X"16",X"00",X"0A",X"13",X"0A",X"00",X"0A",X"0A",X"16",X"00",X"0A",
		X"14",X"0A",X"00",X"0A",X"0A",X"16",X"21",X"0A",X"13",X"0A",X"22",X"0A",X"0A",X"16",X"00",X"0A",
		X"11",X"0A",X"24",X"0A",X"0A",X"16",X"00",X"0A",X"0F",X"0A",X"26",X"0A",X"0E",X"02",X"00",X"0A",
		X"03",X"03",X"27",X"0A",X"03",X"0F",X"00",X"0A",X"07",X"03",X"00",X"0A",X"03",X"0F",X"2B",X"0A",
		X"0A",X"03",X"00",X"0A",X"03",X"0F",X"00",X"0A",X"0C",X"03",X"00",X"0A",X"03",X"0F",X"00",X"0A",
		X"0D",X"03",X"00",X"0A",X"03",X"0F",X"2B",X"0A",X"0C",X"03",X"00",X"0A",X"03",X"0F",X"2B",X"0A",
		X"0A",X"03",X"29",X"0A",X"03",X"0F",X"27",X"0A",X"08",X"03",X"00",X"0A",X"07",X"09",X"00",X"0A",
		X"0A",X"0A",X"26",X"0A",X"0A",X"16",X"00",X"0A",X"0E",X"0A",X"00",X"0A",X"0A",X"16",X"22",X"0A",
		X"11",X"0A",X"00",X"0A",X"0A",X"16",X"00",X"0A",X"13",X"0A",X"00",X"0A",X"0A",X"16",X"00",X"0A",
		X"14",X"0A",X"00",X"0A",X"0A",X"16",X"00",X"0A",X"13",X"0A",X"1D",X"0A",X"0A",X"16",X"00",X"0A",
		X"11",X"0A",X"22",X"0A",X"0A",X"16",X"00",X"0A",X"0F",X"0A",X"24",X"0A",X"0E",X"09",X"00",X"0A",
		X"0A",X"0A",X"26",X"0A",X"0A",X"16",X"00",X"0A",X"0E",X"0A",X"00",X"0A",X"0A",X"16",X"26",X"0A",
		X"11",X"0A",X"00",X"0A",X"0A",X"16",X"00",X"0A",X"0F",X"0A",X"27",X"0A",X"0E",X"04",X"00",X"0A",
		X"05",X"05",X"24",X"0A",X"05",X"11",X"00",X"0A",X"09",X"05",X"24",X"0A",X"05",X"11",X"00",X"0A",
		X"0C",X"05",X"00",X"0A",X"05",X"11",X"26",X"0A",X"0A",X"05",X"00",X"0A",X"09",X"09",X"22",X"0A",
		X"0A",X"0A",X"00",X"0A",X"0A",X"16",X"00",X"0A",X"0E",X"0A",X"00",X"0A",X"0A",X"16",X"00",X"0A",
		X"11",X"0A",X"00",X"0A",X"11",X"16",X"00",X"0A",X"0D",X"0A",X"00",X"0A",X"0E",X"16",X"00",X"0A",
		X"0A",X"0A",X"00",X"0A",X"00",X"00",X"00",X"FF",X"12",X"12",X"12",X"01",X"00",X"00",X"00",X"28",
		X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3A",X"ED",X"61",X"FE",X"01",X"C8",X"3A",X"7C",X"61",X"FE",X"00",X"C2",X"31",X"55",X"DD",X"21",
		X"76",X"61",X"AF",X"7D",X"47",X"DD",X"7E",X"00",X"80",X"27",X"DD",X"77",X"00",X"7C",X"47",X"DD",
		X"7E",X"01",X"88",X"27",X"DD",X"77",X"01",X"DD",X"7E",X"02",X"CE",X"00",X"27",X"DD",X"77",X"02",
		X"C9",X"DD",X"21",X"79",X"61",X"18",X"DB",X"FD",X"7E",X"02",X"47",X"DD",X"7E",X"02",X"CD",X"4E",
		X"55",X"FD",X"7E",X"03",X"47",X"DD",X"7E",X"03",X"CD",X"4E",X"55",X"3E",X"01",X"C9",X"4F",X"C6",
		X"0B",X"B8",X"38",X"07",X"79",X"D6",X"08",X"B8",X"30",X"01",X"C9",X"F1",X"AF",X"C9",X"DD",X"21",
		X"80",X"65",X"FD",X"21",X"09",X"60",X"18",X"1A",X"DD",X"21",X"94",X"65",X"FD",X"21",X"38",X"60",
		X"3A",X"99",X"60",X"18",X"10",X"DD",X"21",X"98",X"65",X"FD",X"21",X"78",X"60",X"3A",X"9A",X"60",
		X"18",X"03",X"3A",X"0D",X"60",X"32",X"98",X"60",X"CD",X"8C",X"55",X"C9",X"CD",X"AC",X"55",X"CD",
		X"9A",X"55",X"FD",X"75",X"00",X"FD",X"74",X"01",X"C9",X"C9",X"DD",X"7E",X"03",X"C6",X"10",X"CB",
		X"3F",X"CB",X"3F",X"CB",X"3F",X"85",X"6F",X"7C",X"CE",X"00",X"67",X"C9",X"DD",X"7E",X"02",X"C6",
		X"07",X"2F",X"CB",X"3F",X"C3",X"CD",X"5B",X"00",X"47",X"11",X"20",X"00",X"21",X"00",X"40",X"19",
		X"10",X"FD",X"3A",X"98",X"60",X"FE",X"01",X"C8",X"FE",X"02",X"20",X"05",X"7C",X"C6",X"04",X"67",
		X"C9",X"FE",X"03",X"C0",X"7C",X"C6",X"08",X"67",X"C9",X"01",X"E0",X"FF",X"1A",X"FE",X"3F",X"C8",
		X"D6",X"30",X"77",X"E5",X"7C",X"C6",X"08",X"67",X"3E",X"00",X"77",X"E1",X"13",X"09",X"18",X"E9",
		X"01",X"E0",X"FF",X"1A",X"FE",X"3F",X"C8",X"77",X"E5",X"7C",X"C6",X"08",X"67",X"08",X"77",X"08",
		X"E1",X"13",X"09",X"18",X"EB",X"11",X"20",X"00",X"06",X"1C",X"77",X"19",X"10",X"FC",X"C9",X"DD",
		X"21",X"76",X"61",X"21",X"E1",X"92",X"CD",X"3C",X"56",X"DD",X"21",X"79",X"61",X"21",X"61",X"90",
		X"CD",X"3C",X"56",X"DD",X"21",X"E8",X"61",X"21",X"01",X"92",X"06",X"01",X"CD",X"41",X"56",X"DD",
		X"21",X"E9",X"61",X"21",X"C1",X"91",X"06",X"01",X"CD",X"41",X"56",X"C9",X"06",X"03",X"11",X"20",
		X"00",X"DD",X"7E",X"00",X"CD",X"4D",X"56",X"DD",X"23",X"19",X"10",X"F5",X"C9",X"F5",X"E6",X"0F",
		X"77",X"19",X"F1",X"CB",X"0F",X"CB",X"0F",X"CB",X"0F",X"CB",X"0F",X"E6",X"0F",X"77",X"C9",X"ED",
		X"52",X"06",X"11",X"CD",X"6A",X"56",X"CD",X"75",X"56",X"C9",X"78",X"77",X"E5",X"7C",X"C6",X"08",
		X"67",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"50",X"4C",X"41",X"59",X"45",X"52",X"10",X"31",X"3F",X"43",X"52",X"45",X"44",X"49",X"54",X"3F",
		X"10",X"10",X"10",X"48",X"49",X"47",X"48",X"10",X"53",X"43",X"4F",X"52",X"45",X"10",X"10",X"10",
		X"3F",X"47",X"41",X"4D",X"45",X"10",X"4F",X"56",X"45",X"52",X"10",X"3F",X"10",X"10",X"10",X"10",
		X"10",X"49",X"4E",X"53",X"45",X"52",X"54",X"10",X"43",X"30",X"49",X"4E",X"53",X"10",X"10",X"10",
		X"10",X"10",X"3F",X"10",X"10",X"10",X"10",X"10",X"50",X"55",X"53",X"48",X"10",X"53",X"54",X"41",
		X"52",X"54",X"10",X"42",X"55",X"54",X"54",X"4F",X"4E",X"10",X"10",X"10",X"10",X"10",X"3F",X"10",
		X"4F",X"4E",X"45",X"10",X"50",X"4C",X"41",X"59",X"45",X"52",X"10",X"4F",X"4E",X"4C",X"59",X"10",
		X"10",X"3F",X"4F",X"4E",X"45",X"10",X"4F",X"52",X"10",X"54",X"57",X"4F",X"10",X"50",X"4C",X"41",
		X"59",X"45",X"52",X"53",X"3F",X"42",X"4F",X"4E",X"55",X"53",X"3F",X"56",X"41",X"4C",X"41",X"44",
		X"4F",X"4E",X"10",X"41",X"55",X"54",X"4F",X"4D",X"41",X"54",X"49",X"4F",X"4E",X"3F",X"10",X"10",
		X"10",X"10",X"10",X"10",X"4D",X"4F",X"56",X"45",X"10",X"4A",X"4F",X"59",X"53",X"54",X"49",X"43",
		X"4B",X"10",X"10",X"10",X"10",X"10",X"3F",X"10",X"10",X"54",X"4F",X"10",X"44",X"49",X"53",X"50",
		X"4C",X"41",X"59",X"10",X"59",X"4F",X"55",X"52",X"10",X"4E",X"41",X"4D",X"45",X"10",X"3F",X"53",
		X"43",X"4F",X"52",X"45",X"3F",X"4E",X"41",X"4D",X"45",X"3F",X"50",X"4C",X"41",X"59",X"45",X"52",
		X"10",X"31",X"3F",X"50",X"4C",X"41",X"59",X"45",X"52",X"10",X"32",X"3F",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"3F",X"10",X"10",X"45",X"4E",X"44",X"10",X"42",X"59",X"10",X"41",X"43",
		X"54",X"49",X"4F",X"4E",X"10",X"42",X"55",X"54",X"54",X"4F",X"4E",X"10",X"10",X"10",X"3F",X"43",
		X"4F",X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"10",X"31",X"39",X"38",X"32",X"3F",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"3F",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"3F",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"3F",X"4A",X"45",X"55",X"10",X"4C",X"45",
		X"10",X"42",X"41",X"47",X"4E",X"41",X"52",X"44",X"3F",X"42",X"52",X"49",X"53",X"53",X"45",X"10",
		X"4A",X"41",X"43",X"51",X"55",X"45",X"53",X"3F",X"37",X"31",X"35",X"33",X"30",X"10",X"43",X"48",
		X"41",X"4C",X"4F",X"4E",X"10",X"53",X"55",X"52",X"10",X"53",X"41",X"4F",X"4E",X"45",X"3F",X"46",
		X"52",X"41",X"4E",X"43",X"45",X"3F",X"4A",X"4F",X"55",X"45",X"55",X"52",X"10",X"31",X"3F",X"43",
		X"52",X"45",X"44",X"49",X"54",X"3F",X"4D",X"45",X"49",X"4C",X"4C",X"45",X"55",X"52",X"53",X"10",
		X"53",X"43",X"4F",X"52",X"45",X"53",X"3F",X"4A",X"45",X"55",X"10",X"46",X"49",X"4E",X"49",X"10",
		X"10",X"3F",X"49",X"4E",X"54",X"52",X"4F",X"44",X"55",X"49",X"53",X"45",X"5A",X"10",X"56",X"4F",
		X"53",X"10",X"50",X"49",X"45",X"43",X"45",X"53",X"3F",X"41",X"50",X"50",X"55",X"59",X"45",X"5A",
		X"10",X"53",X"55",X"52",X"10",X"4C",X"45",X"10",X"42",X"4F",X"55",X"54",X"4F",X"4E",X"10",X"53",
		X"54",X"41",X"52",X"54",X"3F",X"31",X"10",X"4A",X"4F",X"55",X"45",X"55",X"52",X"10",X"53",X"45",
		X"55",X"4C",X"45",X"4D",X"45",X"4E",X"54",X"3F",X"10",X"10",X"31",X"10",X"4F",X"55",X"10",X"32",
		X"10",X"4A",X"4F",X"55",X"45",X"55",X"52",X"53",X"10",X"10",X"3F",X"42",X"4F",X"4E",X"55",X"53",
		X"3F",X"56",X"41",X"4C",X"41",X"44",X"4F",X"4E",X"10",X"41",X"55",X"54",X"4F",X"4D",X"41",X"54",
		X"49",X"4F",X"4E",X"3F",X"55",X"54",X"49",X"4C",X"49",X"53",X"45",X"5A",X"10",X"4C",X"45",X"10",
		X"4D",X"41",X"4E",X"49",X"50",X"55",X"4C",X"41",X"54",X"45",X"55",X"52",X"3F",X"50",X"4F",X"55",
		X"52",X"10",X"49",X"4E",X"53",X"43",X"52",X"49",X"52",X"45",X"10",X"56",X"4F",X"54",X"52",X"45",
		X"10",X"4E",X"4F",X"4D",X"3F",X"53",X"43",X"4F",X"52",X"45",X"3F",X"4E",X"4F",X"4D",X"10",X"3F",
		X"4A",X"4F",X"55",X"45",X"55",X"52",X"10",X"31",X"3F",X"4A",X"4F",X"55",X"45",X"55",X"52",X"10",
		X"32",X"3F",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"3F",X"10",X"10",X"10",X"41",X"43",
		X"54",X"49",X"4F",X"4E",X"10",X"50",X"4F",X"55",X"52",X"10",X"46",X"49",X"4E",X"49",X"52",X"10",
		X"10",X"10",X"10",X"10",X"3F",X"43",X"4F",X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"10",X"31",
		X"39",X"38",X"32",X"3F",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"3F",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"3F",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"3F",
		X"80",X"40",X"20",X"10",X"40",X"A4",X"E0",X"40",X"A9",X"90",X"43",X"24",X"A0",X"43",X"30",X"B0",
		X"43",X"35",X"B0",X"43",X"3D",X"D0",X"40",X"D4",X"D0",X"41",X"54",X"E0",X"41",X"5D",X"D0",X"41",
		X"D4",X"90",X"44",X"E4",X"E0",X"44",X"EC",X"B0",X"44",X"FA",X"D0",X"44",X"BE",X"D0",X"47",X"09",
		X"D0",X"48",X"A4",X"E0",X"49",X"A4",X"E0",X"48",X"AC",X"F0",X"49",X"AC",X"D0",X"48",X"B2",X"70",
		X"48",X"BA",X"F0",X"48",X"BE",X"D0",X"4B",X"2C",X"E0",X"4B",X"3A",X"D0",X"31",X"A4",X"E0",X"31",
		X"F0",X"E0",X"31",X"FA",X"D0",X"36",X"D0",X"D0",X"37",X"70",X"D0",X"D0",X"78",X"B0",X"46",X"7E",
		X"D0",X"46",X"C4",X"E0",X"48",X"E4",X"E0",X"48",X"87",X"60",X"48",X"8B",X"50",X"48",X"EB",X"E0",
		X"4A",X"27",X"E0",X"4A",X"2B",X"90",X"48",X"F4",X"D0",X"48",X"94",X"60",X"48",X"9B",X"50",X"49",
		X"D1",X"60",X"49",X"D4",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"58",X"93",X"02",X"A8",X"91",X"01",X"12",X"91",
		X"01",X"98",X"90",X"01",X"2E",X"93",X"01",X"36",X"93",X"01",X"C8",X"91",X"02",X"4C",X"92",X"02",
		X"CA",X"90",X"02",X"CD",X"90",X"02",X"91",X"90",X"02",X"9C",X"90",X"02",X"62",X"90",X"03",X"65",
		X"91",X"03",X"69",X"91",X"03",X"15",X"92",X"03",X"99",X"92",X"03",X"39",X"91",X"03",X"F1",X"F2",
		X"F3",X"F4",X"F5",X"F6",X"F7",X"1F",X"1F",X"1F",X"FF",X"09",X"00",X"1F",X"1F",X"1F",X"FF",X"02",
		X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"20",X"00",X"00",X"03",X"00",X"00",X"00",X"15",
		X"1B",X"00",X"00",X"0C",X"1B",X"00",X"00",X"0C",X"1B",X"00",X"00",X"0C",X"1C",X"00",X"00",X"0C",
		X"1B",X"00",X"00",X"0C",X"00",X"00",X"00",X"0C",X"1F",X"00",X"00",X"16",X"20",X"00",X"00",X"0C",
		X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"FF",X"24",X"19",X"00",X"0C",X"20",X"1A",X"00",X"0C",
		X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"FF",X"1B",X"00",X"00",X"0C",X"20",X"00",X"00",X"0C",
		X"24",X"00",X"00",X"0C",X"27",X"00",X"00",X"0C",X"24",X"00",X"00",X"0C",X"00",X"00",X"00",X"0C",
		X"00",X"00",X"00",X"FF",X"1B",X"00",X"00",X"0C",X"20",X"00",X"00",X"0C",X"24",X"00",X"00",X"0C",
		X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"FF",X"1B",X"0F",X"00",X"02",X"18",X"0E",X"00",X"0C",
		X"14",X"0E",X"00",X"0C",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"FF",X"7F",X"75",X"CE",X"99",
		X"C0",X"8B",X"C4",X"82",X"65",X"96",X"01",X"9E",X"65",X"8B",X"B4",X"8D",X"B0",X"CB",X"3F",X"CB",
		X"3F",X"FE",X"00",X"CA",X"C2",X"55",X"C3",X"B8",X"55",X"20",X"00",X"00",X"02",X"00",X"00",X"00",
		X"08",X"1B",X"00",X"00",X"0F",X"1B",X"00",X"00",X"08",X"1B",X"00",X"00",X"08",X"1C",X"00",X"00",
		X"08",X"00",X"00",X"00",X"08",X"1B",X"00",X"00",X"08",X"00",X"00",X"00",X"08",X"1F",X"00",X"00",
		X"20",X"20",X"00",X"00",X"0F",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"FF",X"FF",X"08",X"00",
		X"3A",X"F5",X"61",X"FE",X"00",X"C2",X"68",X"05",X"3A",X"CF",X"61",X"FE",X"00",X"C2",X"68",X"05",
		X"C3",X"5B",X"05",X"26",X"3A",X"F5",X"61",X"FE",X"00",X"C2",X"52",X"06",X"3A",X"CF",X"61",X"FE",
		X"00",X"C2",X"52",X"06",X"C3",X"45",X"06",X"05",X"50",X"50",X"49",X"60",X"46",X"44",X"0C",X"04",
		X"3A",X"59",X"61",X"FE",X"01",X"C8",X"3A",X"5E",X"61",X"FE",X"01",X"C8",X"0A",X"D9",X"FE",X"00",
		X"C3",X"AE",X"23",X"FF",X"58",X"93",X"02",X"A8",X"91",X"01",X"12",X"91",X"01",X"98",X"90",X"01",
		X"DC",X"91",X"01",X"36",X"93",X"01",X"71",X"90",X"01",X"4C",X"92",X"02",X"CA",X"90",X"02",X"C5",
		X"90",X"02",X"91",X"90",X"02",X"9C",X"90",X"02",X"71",X"93",X"03",X"85",X"92",X"03",X"C9",X"91",
		X"03",X"15",X"92",X"03",X"99",X"92",X"03",X"F9",X"90",X"03",X"FF",X"10",X"FF",X"FF",X"FF",X"FF",
		X"3A",X"54",X"60",X"FE",X"00",X"C8",X"CD",X"00",X"55",X"C9",X"C3",X"46",X"5E",X"FE",X"01",X"C8",
		X"DD",X"21",X"44",X"5D",X"FD",X"21",X"80",X"65",X"11",X"04",X"00",X"3A",X"88",X"62",X"FE",X"00",
		X"CC",X"2A",X"5D",X"3A",X"88",X"62",X"FE",X"00",X"28",X"05",X"DD",X"19",X"3D",X"18",X"F7",X"DD",
		X"7E",X"03",X"FE",X"FF",X"28",X"3C",X"FE",X"FE",X"CA",X"1C",X"5D",X"47",X"3A",X"26",X"60",X"E6",
		X"07",X"B0",X"32",X"26",X"60",X"FD",X"7E",X"02",X"DD",X"BE",X"00",X"C0",X"FD",X"7E",X"03",X"DD",
		X"BE",X"01",X"C0",X"3A",X"0D",X"60",X"DD",X"BE",X"02",X"C0",X"3A",X"88",X"62",X"3C",X"32",X"88",
		X"62",X"3A",X"26",X"60",X"E6",X"80",X"FE",X"80",X"C8",X"3A",X"26",X"60",X"E6",X"07",X"32",X"26",
		X"60",X"C9",X"3E",X"10",X"32",X"97",X"65",X"32",X"9B",X"65",X"3E",X"D0",X"32",X"96",X"65",X"3E",
		X"E0",X"C3",X"38",X"5E",X"3A",X"87",X"65",X"FE",X"11",X"C0",X"18",X"CE",X"3A",X"8A",X"65",X"FE",
		X"7F",X"C0",X"3A",X"19",X"60",X"FE",X"01",X"C0",X"18",X"C0",X"21",X"C2",X"91",X"22",X"C4",X"61",
		X"22",X"FA",X"61",X"3E",X"01",X"32",X"C6",X"61",X"32",X"FC",X"61",X"3E",X"03",X"32",X"99",X"60",
		X"32",X"9A",X"60",X"C9",X"3C",X"E0",X"01",X"10",X"3C",X"70",X"01",X"20",X"28",X"70",X"01",X"08",
		X"28",X"70",X"01",X"80",X"28",X"70",X"01",X"00",X"28",X"70",X"01",X"00",X"28",X"70",X"01",X"00",
		X"39",X"70",X"01",X"10",X"3C",X"11",X"01",X"20",X"85",X"10",X"01",X"10",X"85",X"10",X"01",X"80",
		X"85",X"10",X"01",X"00",X"85",X"10",X"01",X"00",X"85",X"10",X"01",X"00",X"56",X"10",X"01",X"08",
		X"7D",X"10",X"01",X"10",X"7D",X"10",X"01",X"80",X"7D",X"10",X"01",X"00",X"7D",X"10",X"01",X"00",
		X"7D",X"10",X"01",X"00",X"6C",X"10",X"02",X"10",X"6C",X"10",X"02",X"80",X"6C",X"10",X"02",X"00",
		X"6C",X"10",X"02",X"00",X"6C",X"10",X"02",X"00",X"8C",X"10",X"02",X"10",X"8C",X"10",X"02",X"FF",
		X"98",X"10",X"02",X"10",X"98",X"88",X"02",X"00",X"38",X"88",X"02",X"08",X"38",X"88",X"02",X"80",
		X"38",X"88",X"02",X"00",X"38",X"88",X"02",X"00",X"38",X"88",X"02",X"00",X"38",X"88",X"02",X"00",
		X"38",X"88",X"02",X"00",X"38",X"88",X"02",X"00",X"38",X"88",X"02",X"00",X"38",X"88",X"02",X"00",
		X"38",X"88",X"02",X"00",X"38",X"88",X"02",X"00",X"38",X"88",X"02",X"00",X"38",X"88",X"02",X"00",
		X"5B",X"88",X"02",X"10",X"5C",X"C0",X"02",X"40",X"40",X"C0",X"02",X"08",X"44",X"C0",X"02",X"10",
		X"40",X"C0",X"02",X"08",X"44",X"C0",X"02",X"10",X"40",X"C0",X"02",X"08",X"59",X"C0",X"02",X"10",
		X"5C",X"E0",X"02",X"40",X"7D",X"E0",X"02",X"10",X"7D",X"E0",X"02",X"80",X"7D",X"E0",X"02",X"FE",
		X"7D",X"E0",X"02",X"80",X"B9",X"E0",X"02",X"00",X"B4",X"C8",X"02",X"20",X"B8",X"C8",X"02",X"10",
		X"FF",X"FF",X"FF",X"10",X"60",X"FF",X"FF",X"FF",X"32",X"9A",X"65",X"3E",X"03",X"32",X"99",X"60",
		X"32",X"9A",X"60",X"C3",X"14",X"5D",X"3A",X"54",X"60",X"FE",X"01",X"C8",X"3A",X"26",X"60",X"E6",
		X"07",X"32",X"26",X"60",X"C3",X"A0",X"5C",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3E",X"0A",X"32",X"7D",X"62",X"0E",X"01",X"C9",X"FF",X"32",X"ED",X"61",X"3E",X"0A",X"32",X"7D",
		X"62",X"C3",X"C9",X"38",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
