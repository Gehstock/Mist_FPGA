-- generated with romgen by MikeJ
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ROM_SND_0 is
  port (
    CLK         : in    std_logic;
    ADDR        : in    std_logic_vector(10 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_SND_0 is


  type ROM_ARRAY is array(0 to 2047) of std_logic_vector(7 downto 0);
  constant ROM : ROM_ARRAY := (
    x"C3",x"CE",x"01",x"01",x"F7",x"00",x"01",x"DC", -- 0x0000
    x"00",x"01",x"15",x"01",x"01",x"F7",x"00",x"01", -- 0x0008
    x"DC",x"00",x"01",x"D0",x"00",x"01",x"F7",x"00", -- 0x0010
    x"01",x"DC",x"00",x"01",x"D0",x"00",x"01",x"B9", -- 0x0018
    x"00",x"01",x"DC",x"00",x"01",x"D0",x"00",x"01", -- 0x0020
    x"00",x"00",x"01",x"68",x"00",x"FF",x"FF",x"FF", -- 0x0028
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0030
    x"08",x"D9",x"3E",x"0E",x"D3",x"40",x"DB",x"80", -- 0x0038
    x"B7",x"28",x"32",x"57",x"E6",x"0F",x"20",x"3B", -- 0x0040
    x"7A",x"FE",x"10",x"28",x"3E",x"FE",x"20",x"28", -- 0x0048
    x"43",x"FE",x"30",x"28",x"48",x"FE",x"40",x"28", -- 0x0050
    x"4D",x"FE",x"50",x"28",x"52",x"FE",x"60",x"28", -- 0x0058
    x"57",x"FE",x"70",x"28",x"5C",x"FE",x"80",x"28", -- 0x0060
    x"61",x"FE",x"90",x"28",x"66",x"FE",x"A0",x"28", -- 0x0068
    x"6B",x"D9",x"08",x"FB",x"C9",x"06",x"06",x"21", -- 0x0070
    x"00",x"80",x"77",x"23",x"05",x"20",x"FB",x"D9", -- 0x0078
    x"08",x"FB",x"C9",x"7A",x"CD",x"01",x"01",x"D9", -- 0x0080
    x"08",x"FB",x"C9",x"3E",x"11",x"CD",x"01",x"01", -- 0x0088
    x"D9",x"08",x"FB",x"C9",x"3E",x"11",x"CD",x"E5", -- 0x0090
    x"00",x"D9",x"08",x"FB",x"C9",x"3E",x"12",x"CD", -- 0x0098
    x"01",x"01",x"D9",x"08",x"FB",x"C9",x"3E",x"12", -- 0x00A0
    x"CD",x"E5",x"00",x"D9",x"08",x"FB",x"C9",x"3E", -- 0x00A8
    x"13",x"CD",x"01",x"01",x"D9",x"08",x"FB",x"C9", -- 0x00B0
    x"3E",x"13",x"CD",x"E5",x"00",x"D9",x"08",x"FB", -- 0x00B8
    x"C9",x"3E",x"14",x"CD",x"01",x"01",x"D9",x"08", -- 0x00C0
    x"FB",x"C9",x"3E",x"14",x"CD",x"E5",x"00",x"D9", -- 0x00C8
    x"08",x"FB",x"C9",x"3E",x"15",x"CD",x"01",x"01", -- 0x00D0
    x"D9",x"08",x"FB",x"C9",x"3E",x"15",x"CD",x"E5", -- 0x00D8
    x"00",x"D9",x"08",x"FB",x"C9",x"CD",x"99",x"01", -- 0x00E0
    x"B7",x"C8",x"FE",x"01",x"28",x"09",x"FE",x"02", -- 0x00E8
    x"28",x"0A",x"AF",x"32",x"04",x"80",x"C9",x"AF", -- 0x00F0
    x"32",x"00",x"80",x"C9",x"AF",x"32",x"02",x"80", -- 0x00F8
    x"C9",x"32",x"06",x"80",x"CD",x"99",x"01",x"B7", -- 0x0100
    x"C0",x"AF",x"CD",x"99",x"01",x"B7",x"20",x"41", -- 0x0108
    x"3A",x"00",x"80",x"CD",x"BC",x"01",x"32",x"07", -- 0x0110
    x"80",x"3A",x"02",x"80",x"CD",x"BC",x"01",x"32", -- 0x0118
    x"08",x"80",x"3A",x"04",x"80",x"CD",x"BC",x"01", -- 0x0120
    x"32",x"09",x"80",x"3A",x"06",x"80",x"CD",x"BC", -- 0x0128
    x"01",x"32",x"0A",x"80",x"3A",x"07",x"80",x"21", -- 0x0130
    x"08",x"80",x"BE",x"FA",x"6E",x"01",x"3A",x"09", -- 0x0138
    x"80",x"BE",x"FA",x"8D",x"01",x"3A",x"0A",x"80", -- 0x0140
    x"BE",x"F8",x"21",x"02",x"80",x"CD",x"C5",x"01", -- 0x0148
    x"C9",x"FE",x"01",x"28",x"0B",x"FE",x"02",x"28", -- 0x0150
    x"0E",x"3A",x"06",x"80",x"32",x"04",x"80",x"C9", -- 0x0158
    x"3A",x"06",x"80",x"32",x"00",x"80",x"C9",x"3A", -- 0x0160
    x"06",x"80",x"32",x"02",x"80",x"C9",x"21",x"09", -- 0x0168
    x"80",x"BE",x"FA",x"81",x"01",x"3A",x"0A",x"80", -- 0x0170
    x"BE",x"F8",x"21",x"04",x"80",x"CD",x"C5",x"01", -- 0x0178
    x"C9",x"21",x"0A",x"80",x"BE",x"F0",x"21",x"00", -- 0x0180
    x"80",x"CD",x"C5",x"01",x"C9",x"21",x"0A",x"80", -- 0x0188
    x"BE",x"F0",x"21",x"04",x"80",x"CD",x"C5",x"01", -- 0x0190
    x"C9",x"06",x"00",x"21",x"00",x"80",x"BE",x"28", -- 0x0198
    x"0C",x"23",x"23",x"BE",x"28",x"0C",x"23",x"23", -- 0x01A0
    x"BE",x"28",x"0C",x"AF",x"C9",x"23",x"70",x"3E", -- 0x01A8
    x"01",x"C9",x"23",x"70",x"3E",x"02",x"C9",x"23", -- 0x01B0
    x"70",x"3E",x"03",x"C9",x"21",x"A1",x"04",x"5F", -- 0x01B8
    x"16",x"00",x"19",x"7E",x"C9",x"3A",x"06",x"80", -- 0x01C0
    x"77",x"3E",x"00",x"23",x"77",x"C9",x"06",x"00", -- 0x01C8
    x"21",x"00",x"80",x"70",x"23",x"7C",x"FE",x"84", -- 0x01D0
    x"20",x"F9",x"31",x"00",x"84",x"ED",x"56",x"3E", -- 0x01D8
    x"07",x"D3",x"40",x"3E",x"3F",x"32",x"0C",x"80", -- 0x01E0
    x"D3",x"80",x"CD",x"FA",x"03",x"CD",x"02",x"04", -- 0x01E8
    x"CD",x"0A",x"04",x"FB",x"3E",x"0F",x"D3",x"40", -- 0x01F0
    x"DB",x"80",x"E6",x"80",x"20",x"F6",x"3E",x"0F", -- 0x01F8
    x"D3",x"40",x"DB",x"80",x"E6",x"80",x"28",x"F6", -- 0x0200
    x"F3",x"3E",x"01",x"32",x"0B",x"80",x"3A",x"01", -- 0x0208
    x"80",x"B7",x"28",x"34",x"3A",x"00",x"80",x"CD", -- 0x0210
    x"2B",x"03",x"FB",x"00",x"00",x"00",x"F3",x"3E", -- 0x0218
    x"02",x"32",x"0B",x"80",x"3A",x"03",x"80",x"B7", -- 0x0220
    x"28",x"26",x"3A",x"02",x"80",x"CD",x"2B",x"03", -- 0x0228
    x"FB",x"00",x"00",x"00",x"F3",x"3E",x"03",x"32", -- 0x0230
    x"0B",x"80",x"3A",x"05",x"80",x"B7",x"28",x"18", -- 0x0238
    x"3A",x"04",x"80",x"CD",x"2B",x"03",x"18",x"AB", -- 0x0240
    x"3A",x"00",x"80",x"CD",x"60",x"02",x"18",x"CA", -- 0x0248
    x"3A",x"02",x"80",x"CD",x"60",x"02",x"18",x"D8", -- 0x0250
    x"3A",x"04",x"80",x"CD",x"60",x"02",x"18",x"93", -- 0x0258
    x"FE",x"01",x"28",x"5C",x"FE",x"02",x"28",x"5D", -- 0x0260
    x"FE",x"03",x"28",x"5E",x"FE",x"04",x"28",x"5F", -- 0x0268
    x"FE",x"05",x"28",x"60",x"FE",x"06",x"28",x"61", -- 0x0270
    x"FE",x"07",x"28",x"62",x"FE",x"08",x"28",x"63", -- 0x0278
    x"FE",x"09",x"28",x"64",x"FE",x"0A",x"28",x"65", -- 0x0280
    x"FE",x"0B",x"28",x"66",x"FE",x"0C",x"28",x"67", -- 0x0288
    x"FE",x"0D",x"28",x"68",x"FE",x"0E",x"28",x"69", -- 0x0290
    x"FE",x"11",x"28",x"6A",x"FE",x"12",x"28",x"6B", -- 0x0298
    x"FE",x"13",x"28",x"6C",x"FE",x"14",x"28",x"6D", -- 0x02A0
    x"FE",x"15",x"28",x"6E",x"CD",x"B7",x"04",x"3A", -- 0x02A8
    x"0B",x"80",x"FE",x"01",x"28",x"69",x"FE",x"02", -- 0x02B0
    x"28",x"6B",x"3E",x"01",x"32",x"05",x"80",x"C9", -- 0x02B8
    x"CD",x"2A",x"05",x"18",x"EA",x"CD",x"90",x"05", -- 0x02C0
    x"18",x"E5",x"CD",x"D8",x"05",x"18",x"E0",x"CD", -- 0x02C8
    x"3A",x"06",x"18",x"DB",x"CD",x"F7",x"08",x"18", -- 0x02D0
    x"D6",x"CD",x"68",x"09",x"18",x"D1",x"CD",x"53", -- 0x02D8
    x"0F",x"18",x"CC",x"CD",x"AE",x"09",x"18",x"C7", -- 0x02E0
    x"CD",x"38",x"0A",x"18",x"C2",x"CD",x"0F",x"0B", -- 0x02E8
    x"18",x"BD",x"CD",x"78",x"0B",x"18",x"B8",x"CD", -- 0x02F0
    x"A3",x"0B",x"18",x"B3",x"CD",x"05",x"0C",x"18", -- 0x02F8
    x"AE",x"CD",x"BA",x"07",x"18",x"A9",x"CD",x"6E", -- 0x0300
    x"0C",x"18",x"A4",x"CD",x"CE",x"0C",x"18",x"9F", -- 0x0308
    x"CD",x"32",x"0E",x"18",x"9A",x"CD",x"F5",x"0E", -- 0x0310
    x"18",x"95",x"CD",x"24",x"0F",x"18",x"90",x"3E", -- 0x0318
    x"01",x"32",x"01",x"80",x"C9",x"3E",x"01",x"32", -- 0x0320
    x"03",x"80",x"C9",x"FE",x"01",x"28",x"49",x"FE", -- 0x0328
    x"02",x"28",x"4A",x"FE",x"03",x"28",x"4B",x"FE", -- 0x0330
    x"04",x"28",x"4C",x"FE",x"05",x"28",x"4D",x"FE", -- 0x0338
    x"06",x"28",x"4E",x"FE",x"07",x"28",x"4F",x"FE", -- 0x0340
    x"08",x"28",x"50",x"FE",x"09",x"28",x"6A",x"FE", -- 0x0348
    x"0A",x"28",x"4D",x"FE",x"0B",x"28",x"4E",x"FE", -- 0x0350
    x"0C",x"28",x"4F",x"FE",x"0D",x"28",x"50",x"FE", -- 0x0358
    x"0E",x"28",x"51",x"FE",x"11",x"28",x"57",x"FE", -- 0x0360
    x"12",x"28",x"58",x"FE",x"13",x"28",x"59",x"FE", -- 0x0368
    x"14",x"28",x"5A",x"FE",x"15",x"28",x"5B",x"C9", -- 0x0370
    x"CD",x"4D",x"05",x"18",x"58",x"CD",x"A4",x"05", -- 0x0378
    x"18",x"53",x"CD",x"EF",x"05",x"18",x"4E",x"CD", -- 0x0380
    x"67",x"06",x"18",x"49",x"CD",x"21",x"09",x"18", -- 0x0388
    x"44",x"CD",x"7C",x"09",x"18",x"3F",x"CD",x"76", -- 0x0390
    x"0F",x"18",x"3A",x"CD",x"D0",x"09",x"18",x"35", -- 0x0398
    x"CD",x"2C",x"0B",x"18",x"30",x"CD",x"8C",x"0B", -- 0x03A0
    x"18",x"2B",x"CD",x"BA",x"0B",x"18",x"26",x"CD", -- 0x03A8
    x"22",x"0C",x"18",x"21",x"CD",x"E0",x"07",x"18", -- 0x03B0
    x"1C",x"CD",x"5E",x"0A",x"18",x"17",x"CD",x"8C", -- 0x03B8
    x"0C",x"18",x"12",x"CD",x"E3",x"0C",x"18",x"0D", -- 0x03C0
    x"CD",x"5E",x"0E",x"18",x"08",x"CD",x"21",x"0F", -- 0x03C8
    x"18",x"03",x"CD",x"50",x"0F",x"B7",x"C8",x"3A", -- 0x03D0
    x"0B",x"80",x"FE",x"01",x"28",x"0C",x"FE",x"02", -- 0x03D8
    x"28",x"10",x"AF",x"32",x"04",x"80",x"32",x"05", -- 0x03E0
    x"80",x"C9",x"AF",x"32",x"00",x"80",x"32",x"01", -- 0x03E8
    x"80",x"C9",x"AF",x"32",x"02",x"80",x"32",x"03", -- 0x03F0
    x"80",x"C9",x"3E",x"08",x"D3",x"40",x"AF",x"D3", -- 0x03F8
    x"80",x"C9",x"3E",x"09",x"D3",x"40",x"AF",x"D3", -- 0x0400
    x"80",x"C9",x"3E",x"0A",x"D3",x"40",x"AF",x"D3", -- 0x0408
    x"80",x"C9",x"3A",x"0B",x"80",x"FE",x"01",x"28", -- 0x0410
    x"14",x"FE",x"02",x"28",x"14",x"06",x"04",x"78", -- 0x0418
    x"D3",x"40",x"7D",x"D3",x"80",x"04",x"78",x"D3", -- 0x0420
    x"40",x"7C",x"D3",x"80",x"C9",x"06",x"00",x"18", -- 0x0428
    x"EE",x"06",x"02",x"18",x"EA",x"3A",x"0B",x"80", -- 0x0430
    x"FE",x"01",x"28",x"14",x"FE",x"02",x"28",x"14", -- 0x0438
    x"06",x"04",x"78",x"D3",x"40",x"DB",x"80",x"6F", -- 0x0440
    x"04",x"78",x"D3",x"40",x"DB",x"80",x"67",x"C9", -- 0x0448
    x"06",x"00",x"18",x"EE",x"06",x"02",x"18",x"EA", -- 0x0450
    x"3A",x"0B",x"80",x"FE",x"01",x"28",x"0C",x"FE", -- 0x0458
    x"02",x"28",x"0E",x"06",x"FB",x"1E",x"20",x"CD", -- 0x0460
    x"77",x"04",x"C9",x"06",x"FE",x"1E",x"08",x"18", -- 0x0468
    x"F6",x"06",x"FD",x"1E",x"10",x"18",x"F0",x"3E", -- 0x0470
    x"07",x"D3",x"40",x"3A",x"0C",x"80",x"A0",x"B3", -- 0x0478
    x"32",x"0C",x"80",x"D3",x"80",x"C9",x"3A",x"0B", -- 0x0480
    x"80",x"FE",x"01",x"28",x"0C",x"FE",x"02",x"28", -- 0x0488
    x"0C",x"3E",x"0A",x"D3",x"40",x"78",x"D3",x"80", -- 0x0490
    x"C9",x"3E",x"08",x"18",x"F6",x"3E",x"09",x"18", -- 0x0498
    x"F2",x"00",x"0B",x"06",x"01",x"0C",x"08",x"04", -- 0x04A0
    x"09",x"07",x"0A",x"05",x"03",x"02",x"0D",x"0E", -- 0x04A8
    x"0F",x"10",x"11",x"12",x"13",x"14",x"15",x"3A", -- 0x04B0
    x"0B",x"80",x"FE",x"01",x"28",x"0D",x"FE",x"02", -- 0x04B8
    x"28",x"12",x"06",x"24",x"CD",x"DD",x"04",x"CD", -- 0x04C0
    x"0A",x"04",x"C9",x"06",x"09",x"CD",x"DD",x"04", -- 0x04C8
    x"CD",x"FA",x"03",x"C9",x"06",x"12",x"CD",x"DD", -- 0x04D0
    x"04",x"CD",x"02",x"04",x"C9",x"3E",x"07",x"D3", -- 0x04D8
    x"40",x"3A",x"0C",x"80",x"B0",x"32",x"0C",x"80", -- 0x04E0
    x"D3",x"80",x"C9",x"3A",x"0B",x"80",x"FE",x"01", -- 0x04E8
    x"28",x"0C",x"FE",x"02",x"28",x"0E",x"06",x"DF", -- 0x04F0
    x"1E",x"04",x"CD",x"77",x"04",x"C9",x"06",x"F7", -- 0x04F8
    x"1E",x"01",x"18",x"F6",x"06",x"EF",x"1E",x"02", -- 0x0500
    x"18",x"F0",x"D3",x"40",x"78",x"D3",x"80",x"C9", -- 0x0508
    x"3A",x"0B",x"80",x"FE",x"01",x"28",x"0B",x"FE", -- 0x0510
    x"02",x"28",x"0B",x"3E",x"0A",x"D3",x"40",x"DB", -- 0x0518
    x"80",x"C9",x"3E",x"08",x"18",x"F7",x"3E",x"09", -- 0x0520
    x"18",x"F3",x"3E",x"02",x"32",x"10",x"80",x"21", -- 0x0528
    x"00",x"01",x"22",x"11",x"80",x"3E",x"01",x"32", -- 0x0530
    x"13",x"80",x"AF",x"32",x"14",x"80",x"21",x"C0", -- 0x0538
    x"00",x"CD",x"12",x"04",x"CD",x"58",x"04",x"06", -- 0x0540
    x"0F",x"CD",x"86",x"04",x"C9",x"21",x"10",x"80", -- 0x0548
    x"35",x"20",x"0A",x"3E",x"02",x"77",x"CD",x"35", -- 0x0550
    x"04",x"2B",x"CD",x"12",x"04",x"3A",x"14",x"80", -- 0x0558
    x"FE",x"00",x"28",x"15",x"21",x"13",x"80",x"35", -- 0x0560
    x"20",x"0D",x"3E",x"01",x"77",x"CD",x"10",x"05", -- 0x0568
    x"3D",x"28",x"1A",x"47",x"CD",x"86",x"04",x"AF", -- 0x0570
    x"C9",x"2A",x"11",x"80",x"2B",x"7C",x"B5",x"28", -- 0x0578
    x"05",x"22",x"11",x"80",x"18",x"F1",x"3E",x"01", -- 0x0580
    x"32",x"14",x"80",x"18",x"EA",x"3E",x"FF",x"C9", -- 0x0588
    x"3E",x"10",x"32",x"16",x"80",x"21",x"80",x"00", -- 0x0590
    x"CD",x"12",x"04",x"CD",x"58",x"04",x"06",x"0F", -- 0x0598
    x"CD",x"86",x"04",x"C9",x"21",x"16",x"80",x"35", -- 0x05A0
    x"28",x"1A",x"CD",x"35",x"04",x"11",x"04",x"00", -- 0x05A8
    x"19",x"11",x"00",x"01",x"7C",x"BA",x"20",x"07", -- 0x05B0
    x"7D",x"BB",x"20",x"03",x"21",x"80",x"00",x"CD", -- 0x05B8
    x"12",x"04",x"AF",x"C9",x"3E",x"10",x"32",x"16", -- 0x05C0
    x"80",x"CD",x"10",x"05",x"3D",x"28",x"06",x"47", -- 0x05C8
    x"CD",x"86",x"04",x"18",x"D5",x"3E",x"FF",x"C9", -- 0x05D0
    x"3E",x"01",x"32",x"18",x"80",x"3E",x"08",x"32", -- 0x05D8
    x"19",x"80",x"AF",x"32",x"1A",x"80",x"CD",x"58", -- 0x05E0
    x"04",x"06",x"00",x"CD",x"86",x"04",x"C9",x"3A", -- 0x05E8
    x"1A",x"80",x"FE",x"00",x"28",x"24",x"FE",x"01", -- 0x05F0
    x"28",x"31",x"CD",x"35",x"04",x"01",x"40",x"00", -- 0x05F8
    x"B7",x"ED",x"42",x"CD",x"12",x"04",x"21",x"19", -- 0x0600
    x"80",x"35",x"20",x"0C",x"36",x"08",x"CD",x"10", -- 0x0608
    x"05",x"3D",x"28",x"23",x"47",x"CD",x"86",x"04", -- 0x0610
    x"AF",x"C9",x"21",x"00",x"04",x"CD",x"12",x"04", -- 0x0618
    x"06",x"0F",x"CD",x"86",x"04",x"21",x"1A",x"80", -- 0x0620
    x"34",x"18",x"ED",x"21",x"18",x"80",x"35",x"20", -- 0x0628
    x"E7",x"21",x"1A",x"80",x"34",x"18",x"E1",x"3E", -- 0x0630
    x"FF",x"C9",x"3E",x"0B",x"32",x"1C",x"80",x"32", -- 0x0638
    x"1D",x"80",x"21",x"18",x"07",x"22",x"1E",x"80", -- 0x0640
    x"AF",x"32",x"20",x"80",x"32",x"21",x"80",x"21", -- 0x0648
    x"8A",x"00",x"CD",x"12",x"04",x"CD",x"58",x"04", -- 0x0650
    x"06",x"0F",x"CD",x"86",x"04",x"3E",x"0E",x"32", -- 0x0658
    x"04",x"80",x"AF",x"32",x"05",x"80",x"C9",x"3A", -- 0x0660
    x"20",x"80",x"FE",x"01",x"28",x"14",x"FE",x"02", -- 0x0668
    x"28",x"24",x"3A",x"21",x"80",x"FE",x"44",x"28", -- 0x0670
    x"3E",x"E6",x"01",x"20",x"49",x"CD",x"F0",x"06", -- 0x0678
    x"AF",x"C9",x"CD",x"10",x"05",x"C6",x"05",x"FE", -- 0x0680
    x"0F",x"20",x"05",x"21",x"20",x"80",x"36",x"00", -- 0x0688
    x"47",x"CD",x"86",x"04",x"18",x"EA",x"CD",x"10", -- 0x0690
    x"05",x"D6",x"05",x"20",x"05",x"21",x"20",x"80", -- 0x0698
    x"36",x"00",x"47",x"CD",x"86",x"04",x"3A",x"20", -- 0x06A0
    x"80",x"FE",x"00",x"20",x"D3",x"3A",x"21",x"80", -- 0x06A8
    x"FE",x"44",x"20",x"CC",x"3E",x"FF",x"C9",x"CD", -- 0x06B0
    x"04",x"07",x"B7",x"20",x"02",x"18",x"C1",x"21", -- 0x06B8
    x"20",x"80",x"36",x"02",x"18",x"BA",x"CD",x"CB", -- 0x06C0
    x"06",x"18",x"B5",x"CD",x"04",x"07",x"B7",x"C8", -- 0x06C8
    x"ED",x"5B",x"1E",x"80",x"1A",x"32",x"1D",x"80", -- 0x06D0
    x"13",x"1A",x"6F",x"13",x"1A",x"67",x"13",x"ED", -- 0x06D8
    x"53",x"1E",x"80",x"CD",x"12",x"04",x"21",x"21", -- 0x06E0
    x"80",x"34",x"21",x"20",x"80",x"36",x"01",x"C9", -- 0x06E8
    x"CD",x"04",x"07",x"B7",x"C8",x"3E",x"01",x"32", -- 0x06F0
    x"1D",x"80",x"21",x"21",x"80",x"34",x"21",x"20", -- 0x06F8
    x"80",x"36",x"02",x"C9",x"21",x"1C",x"80",x"35", -- 0x0700
    x"20",x"0C",x"3E",x"0B",x"77",x"21",x"1D",x"80", -- 0x0708
    x"35",x"20",x"03",x"3E",x"FF",x"C9",x"AF",x"C9", -- 0x0710
    x"01",x"8A",x"00",x"01",x"8A",x"00",x"0B",x"8A", -- 0x0718
    x"00",x"01",x"8A",x"00",x"01",x"8A",x"00",x"03", -- 0x0720
    x"8A",x"00",x"03",x"A5",x"00",x"03",x"D0",x"00", -- 0x0728
    x"03",x"A5",x"00",x"03",x"8A",x"00",x"03",x"A5", -- 0x0730
    x"00",x"03",x"8A",x"00",x"03",x"68",x"00",x"03", -- 0x0738
    x"8A",x"00",x"03",x"A5",x"00",x"03",x"D0",x"00", -- 0x0740
    x"03",x"A5",x"00",x"03",x"8A",x"00",x"03",x"A5", -- 0x0748
    x"00",x"03",x"8A",x"00",x"03",x"68",x"00",x"0B", -- 0x0750
    x"8A",x"00",x"01",x"8A",x"00",x"01",x"8A",x"00", -- 0x0758
    x"0B",x"8A",x"00",x"01",x"8A",x"00",x"01",x"8A", -- 0x0760
    x"00",x"0B",x"8A",x"00",x"01",x"8A",x"00",x"01", -- 0x0768
    x"8A",x"00",x"0B",x"8A",x"00",x"01",x"8A",x"00", -- 0x0770
    x"01",x"8A",x"00",x"20",x"8A",x"00",x"01",x"8A", -- 0x0778
    x"00",x"01",x"8A",x"00",x"03",x"8A",x"00",x"03", -- 0x0780
    x"8A",x"00",x"03",x"8A",x"00",x"01",x"8A",x"00", -- 0x0788
    x"01",x"8A",x"00",x"03",x"8A",x"00",x"03",x"8A", -- 0x0790
    x"00",x"03",x"8A",x"00",x"01",x"8A",x"00",x"01", -- 0x0798
    x"8A",x"00",x"03",x"8A",x"00",x"03",x"8A",x"00", -- 0x07A0
    x"03",x"8A",x"00",x"01",x"8A",x"00",x"01",x"8A", -- 0x07A8
    x"00",x"03",x"8A",x"00",x"03",x"8A",x"00",x"20", -- 0x07B0
    x"8A",x"00",x"3E",x"0B",x"32",x"22",x"80",x"3E", -- 0x07B8
    x"0D",x"32",x"23",x"80",x"21",x"91",x"08",x"22", -- 0x07C0
    x"24",x"80",x"AF",x"32",x"26",x"80",x"32",x"27", -- 0x07C8
    x"80",x"21",x"15",x"01",x"CD",x"12",x"04",x"CD", -- 0x07D0
    x"58",x"04",x"06",x"0F",x"CD",x"86",x"04",x"C9", -- 0x07D8
    x"3A",x"26",x"80",x"FE",x"01",x"28",x"14",x"FE", -- 0x07E0
    x"02",x"28",x"24",x"3A",x"27",x"80",x"FE",x"44", -- 0x07E8
    x"28",x"3E",x"E6",x"01",x"20",x"49",x"CD",x"69", -- 0x07F0
    x"08",x"AF",x"C9",x"CD",x"10",x"05",x"C6",x"05"  -- 0x07F8
  );

begin

  p_rom : process
  begin
    wait until rising_edge(CLK);
     DATA <= ROM(to_integer(unsigned(ADDR)));
  end process;
end RTL;
