library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity botanic_program is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of botanic_program is
	type rom is array(0 to  24575) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"F3",X"C3",X"B3",X"03",X"00",X"FF",X"00",X"FF",X"D3",X"08",X"00",X"DB",X"0C",X"C9",X"00",X"FF",
		X"AF",X"32",X"05",X"A0",X"C9",X"00",X"FF",X"00",X"3E",X"01",X"32",X"05",X"A0",X"C9",X"FF",X"00",
		X"C9",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"F5",X"C5",X"D5",X"E5",X"08",X"D9",X"F5",X"C5",
		X"D5",X"E5",X"DD",X"E5",X"FD",X"E5",X"AF",X"32",X"00",X"A0",X"32",X"03",X"A0",X"F3",X"3A",X"00",
		X"B8",X"3A",X"0C",X"71",X"FE",X"00",X"28",X"16",X"3D",X"32",X"0C",X"71",X"FE",X"00",X"20",X"0E",
		X"32",X"06",X"A0",X"3E",X"0A",X"D3",X"08",X"AF",X"D3",X"09",X"3C",X"32",X"06",X"A0",X"3A",X"CC",
		X"70",X"B7",X"C2",X"A0",X"01",X"3A",X"01",X"75",X"FE",X"00",X"CA",X"D7",X"00",X"3A",X"04",X"75",
		X"3D",X"32",X"04",X"75",X"20",X"51",X"D7",X"3E",X"08",X"D3",X"08",X"AF",X"D3",X"09",X"DF",X"DD",
		X"2A",X"15",X"75",X"DD",X"7E",X"00",X"FE",X"FF",X"20",X"07",X"AF",X"32",X"01",X"75",X"C3",X"D7",
		X"00",X"DD",X"7E",X"02",X"32",X"04",X"75",X"D7",X"3E",X"07",X"D3",X"08",X"3E",X"38",X"D3",X"09",
		X"AF",X"D3",X"08",X"DD",X"7E",X"01",X"D3",X"09",X"3E",X"01",X"D3",X"08",X"DD",X"7E",X"00",X"D3",
		X"09",X"DF",X"DD",X"23",X"DD",X"23",X"DD",X"23",X"DD",X"22",X"15",X"75",X"D7",X"3E",X"08",X"D3",
		X"08",X"3A",X"12",X"75",X"D3",X"09",X"DF",X"3A",X"02",X"75",X"FE",X"00",X"CA",X"3A",X"01",X"3A",
		X"05",X"75",X"3D",X"32",X"05",X"75",X"20",X"52",X"D7",X"3E",X"09",X"D3",X"08",X"AF",X"D3",X"09",
		X"DF",X"DD",X"2A",X"17",X"75",X"DD",X"7E",X"00",X"FE",X"FF",X"20",X"07",X"AF",X"32",X"02",X"75",
		X"C3",X"3A",X"01",X"DD",X"7E",X"02",X"32",X"05",X"75",X"D7",X"3E",X"07",X"D3",X"08",X"3E",X"38",
		X"D3",X"09",X"3E",X"02",X"D3",X"08",X"DD",X"7E",X"01",X"D3",X"09",X"3E",X"03",X"D3",X"08",X"DD",
		X"7E",X"00",X"D3",X"09",X"DF",X"DD",X"23",X"DD",X"23",X"DD",X"23",X"DD",X"22",X"17",X"75",X"D7",
		X"3E",X"09",X"D3",X"08",X"3A",X"13",X"75",X"D3",X"09",X"DF",X"3A",X"03",X"75",X"FE",X"00",X"CA",
		X"9D",X"01",X"3A",X"06",X"75",X"3D",X"32",X"06",X"75",X"20",X"52",X"D7",X"3E",X"0A",X"D3",X"08",
		X"AF",X"D3",X"09",X"DF",X"DD",X"2A",X"19",X"75",X"DD",X"7E",X"00",X"FE",X"FF",X"20",X"07",X"AF",
		X"32",X"03",X"75",X"C3",X"9D",X"01",X"DD",X"7E",X"02",X"32",X"06",X"75",X"D7",X"3E",X"07",X"D3",
		X"08",X"3E",X"38",X"D3",X"09",X"3E",X"04",X"D3",X"08",X"DD",X"7E",X"01",X"D3",X"09",X"3E",X"05",
		X"D3",X"08",X"DD",X"7E",X"00",X"D3",X"09",X"DF",X"DD",X"23",X"DD",X"23",X"DD",X"23",X"DD",X"22",
		X"19",X"75",X"D7",X"3E",X"0A",X"D3",X"08",X"3A",X"14",X"75",X"D3",X"09",X"DF",X"CD",X"E4",X"44",
		X"21",X"49",X"70",X"3A",X"94",X"70",X"BE",X"28",X"06",X"AF",X"32",X"03",X"98",X"18",X"0E",X"06",
		X"04",X"21",X"0A",X"74",X"11",X"00",X"98",X"7E",X"12",X"13",X"23",X"10",X"FA",X"21",X"49",X"70",
		X"3A",X"9F",X"70",X"BE",X"28",X"06",X"AF",X"32",X"07",X"98",X"18",X"0E",X"06",X"04",X"21",X"0E",
		X"74",X"11",X"04",X"98",X"7E",X"12",X"13",X"23",X"10",X"FA",X"21",X"49",X"70",X"3A",X"AA",X"70",
		X"BE",X"28",X"06",X"AF",X"32",X"0B",X"98",X"18",X"0E",X"06",X"04",X"21",X"12",X"74",X"11",X"08",
		X"98",X"7E",X"12",X"13",X"23",X"10",X"FA",X"21",X"49",X"70",X"3A",X"87",X"70",X"BE",X"28",X"06",
		X"AF",X"32",X"0F",X"98",X"18",X"0E",X"06",X"04",X"21",X"16",X"74",X"11",X"0C",X"98",X"7E",X"12",
		X"13",X"23",X"10",X"FA",X"21",X"49",X"70",X"3A",X"88",X"70",X"BE",X"28",X"06",X"AF",X"32",X"13",
		X"98",X"18",X"0E",X"06",X"04",X"21",X"1A",X"74",X"11",X"10",X"98",X"7E",X"12",X"13",X"23",X"10",
		X"FA",X"21",X"49",X"70",X"3A",X"89",X"70",X"BE",X"28",X"06",X"AF",X"32",X"17",X"98",X"18",X"0E",
		X"06",X"04",X"21",X"1E",X"74",X"11",X"14",X"98",X"7E",X"12",X"13",X"23",X"10",X"FA",X"06",X"08",
		X"21",X"22",X"74",X"11",X"18",X"98",X"7E",X"12",X"23",X"13",X"10",X"FA",X"3A",X"31",X"70",X"32",
		X"02",X"A0",X"32",X"01",X"A0",X"CD",X"01",X"03",X"CD",X"BB",X"02",X"CD",X"1E",X"03",X"CD",X"80",
		X"03",X"3E",X"01",X"32",X"00",X"A0",X"32",X"03",X"A0",X"ED",X"56",X"FD",X"E1",X"DD",X"E1",X"E1",
		X"D1",X"C1",X"F1",X"D9",X"08",X"E1",X"D1",X"C1",X"F1",X"FB",X"C9",X"AF",X"32",X"06",X"A0",X"3E",
		X"06",X"D3",X"08",X"3E",X"18",X"D3",X"09",X"3E",X"07",X"D3",X"08",X"3E",X"1F",X"D3",X"09",X"3E",
		X"0A",X"D3",X"08",X"3E",X"0F",X"D3",X"09",X"3E",X"08",X"D3",X"08",X"AF",X"D3",X"09",X"3E",X"09",
		X"D3",X"08",X"AF",X"D3",X"09",X"3E",X"01",X"32",X"06",X"A0",X"C9",X"AF",X"32",X"05",X"A0",X"3E",
		X"0E",X"CF",X"32",X"32",X"70",X"3E",X"0F",X"CF",X"32",X"33",X"70",X"3A",X"F4",X"70",X"FE",X"01",
		X"C2",X"F6",X"02",X"3A",X"6F",X"70",X"FE",X"01",X"C2",X"F6",X"02",X"3A",X"33",X"70",X"2F",X"E6",
		X"F8",X"5F",X"3A",X"32",X"70",X"2F",X"E6",X"07",X"B3",X"2F",X"32",X"32",X"70",X"3E",X"01",X"32",
		X"05",X"A0",X"32",X"31",X"70",X"C9",X"3E",X"00",X"32",X"31",X"70",X"3E",X"01",X"32",X"05",X"A0",
		X"C9",X"3A",X"00",X"A8",X"2F",X"E6",X"03",X"FE",X"03",X"28",X"07",X"C6",X"03",X"32",X"34",X"70",
		X"18",X"05",X"3E",X"02",X"32",X"34",X"70",X"00",X"3E",X"06",X"32",X"35",X"70",X"C9",X"3A",X"05",
		X"70",X"FE",X"09",X"C8",X"3A",X"32",X"70",X"2F",X"21",X"36",X"70",X"5F",X"AE",X"73",X"A3",X"CB",
		X"47",X"28",X"05",X"F5",X"CD",X"3E",X"03",X"F1",X"CB",X"4F",X"C4",X"73",X"03",X"C9",X"3A",X"00",
		X"A8",X"2F",X"CB",X"57",X"28",X"16",X"3E",X"01",X"32",X"11",X"75",X"21",X"04",X"70",X"7E",X"FE",
		X"09",X"20",X"03",X"36",X"00",X"23",X"34",X"21",X"FE",X"70",X"34",X"C9",X"3A",X"37",X"70",X"FE",
		X"01",X"20",X"06",X"AF",X"32",X"37",X"70",X"18",X"DD",X"3E",X"01",X"32",X"37",X"70",X"C9",X"21",
		X"FE",X"70",X"34",X"3A",X"00",X"A8",X"2F",X"CB",X"57",X"28",X"CB",X"CD",X"46",X"03",X"18",X"C6",
		X"3A",X"FF",X"70",X"3D",X"32",X"FF",X"70",X"F5",X"FE",X"09",X"C2",X"91",X"03",X"AF",X"32",X"04",
		X"A0",X"F1",X"C0",X"3E",X"12",X"32",X"FF",X"70",X"21",X"FE",X"70",X"7E",X"FE",X"00",X"C8",X"3E",
		X"01",X"32",X"04",X"A0",X"35",X"C9",X"00",X"01",X"01",X"01",X"00",X"01",X"01",X"01",X"01",X"01",
		X"00",X"01",X"31",X"3E",X"FF",X"21",X"00",X"70",X"77",X"BE",X"C2",X"98",X"04",X"4F",X"3A",X"00",
		X"B8",X"79",X"23",X"4F",X"3E",X"78",X"BC",X"79",X"C2",X"B8",X"03",X"FE",X"FF",X"C2",X"D4",X"03",
		X"AF",X"C3",X"B5",X"03",X"31",X"FF",X"77",X"AF",X"32",X"01",X"A0",X"32",X"02",X"A0",X"21",X"00",
		X"70",X"06",X"00",X"70",X"23",X"7C",X"FE",X"78",X"20",X"F9",X"21",X"00",X"98",X"06",X"20",X"36",
		X"00",X"23",X"10",X"FB",X"21",X"0B",X"70",X"06",X"05",X"0E",X"02",X"71",X"7D",X"C6",X"06",X"6F",
		X"10",X"F9",X"3A",X"00",X"A8",X"2F",X"E6",X"80",X"FE",X"80",X"C2",X"17",X"04",X"3E",X"01",X"32",
		X"F4",X"70",X"3E",X"12",X"32",X"FF",X"70",X"06",X"46",X"21",X"0A",X"72",X"36",X"10",X"23",X"10",
		X"FB",X"06",X"2A",X"21",X"6E",X"04",X"11",X"0A",X"72",X"7E",X"D6",X"30",X"12",X"23",X"13",X"10",
		X"F8",X"AF",X"32",X"05",X"A0",X"06",X"C8",X"3E",X"07",X"D3",X"08",X"3E",X"38",X"D3",X"09",X"10",
		X"F6",X"3E",X"01",X"32",X"05",X"A0",X"3E",X"07",X"32",X"11",X"75",X"3E",X"01",X"32",X"0C",X"71",
		X"CD",X"8B",X"02",X"ED",X"56",X"3E",X"01",X"32",X"00",X"A0",X"FB",X"CD",X"E0",X"40",X"11",X"1F",
		X"43",X"21",X"1F",X"8B",X"0E",X"0E",X"CD",X"71",X"41",X"CD",X"A3",X"13",X"18",X"6D",X"48",X"45",
		X"4E",X"4B",X"40",X"53",X"50",X"49",X"54",X"53",X"40",X"40",X"40",X"40",X"4A",X"4F",X"53",X"45",
		X"50",X"40",X"4D",X"5D",X"40",X"50",X"45",X"54",X"49",X"54",X"4A",X"4F",X"53",X"45",X"50",X"40",
		X"4D",X"4F",X"52",X"49",X"4C",X"4C",X"41",X"53",X"21",X"6F",X"8A",X"11",X"20",X"00",X"3E",X"01",
		X"32",X"03",X"A0",X"97",X"36",X"12",X"ED",X"52",X"36",X"11",X"ED",X"52",X"36",X"14",X"ED",X"52",
		X"36",X"10",X"ED",X"52",X"36",X"10",X"ED",X"52",X"36",X"22",X"ED",X"52",X"36",X"11",X"ED",X"52",
		X"36",X"1D",X"21",X"6F",X"9A",X"11",X"20",X"00",X"0E",X"0C",X"06",X"08",X"71",X"3A",X"00",X"B8",
		X"97",X"ED",X"52",X"10",X"F7",X"3A",X"00",X"B8",X"C3",X"D5",X"04",X"AF",X"32",X"31",X"70",X"32",
		X"6F",X"70",X"3E",X"01",X"32",X"CC",X"70",X"21",X"02",X"70",X"36",X"16",X"23",X"36",X"16",X"21",
		X"00",X"06",X"22",X"E6",X"70",X"21",X"00",X"B0",X"22",X"E8",X"70",X"3E",X"03",X"32",X"30",X"70",
		X"CD",X"E0",X"40",X"CD",X"00",X"41",X"CD",X"AC",X"3E",X"CD",X"27",X"41",X"0E",X"15",X"CD",X"4E",
		X"3E",X"CD",X"6A",X"3F",X"CD",X"77",X"08",X"CD",X"0E",X"09",X"CD",X"6F",X"05",X"3A",X"05",X"70",
		X"FE",X"00",X"20",X"6C",X"3A",X"04",X"70",X"FE",X"00",X"C2",X"90",X"05",X"2A",X"E8",X"70",X"2B",
		X"22",X"E8",X"70",X"7C",X"B5",X"C2",X"17",X"05",X"21",X"00",X"B0",X"22",X"E8",X"70",X"3A",X"30",
		X"70",X"3D",X"32",X"30",X"70",X"C2",X"17",X"05",X"3E",X"03",X"32",X"30",X"70",X"AF",X"32",X"0D",
		X"74",X"32",X"11",X"74",X"32",X"15",X"74",X"32",X"19",X"74",X"32",X"1D",X"74",X"32",X"21",X"74",
		X"32",X"25",X"74",X"32",X"29",X"74",X"32",X"22",X"74",X"32",X"26",X"74",X"C3",X"FD",X"2E",X"2A",
		X"E6",X"70",X"2B",X"22",X"E6",X"70",X"7C",X"B5",X"C0",X"3A",X"02",X"70",X"3C",X"FE",X"1F",X"20",
		X"02",X"3E",X"10",X"32",X"02",X"70",X"21",X"00",X"04",X"22",X"E6",X"70",X"CD",X"00",X"41",X"C9",
		X"AF",X"32",X"CC",X"70",X"32",X"0D",X"74",X"32",X"11",X"74",X"32",X"15",X"74",X"32",X"19",X"74",
		X"32",X"1D",X"74",X"32",X"21",X"74",X"32",X"25",X"74",X"32",X"29",X"74",X"32",X"22",X"74",X"32",
		X"26",X"74",X"06",X"3C",X"21",X"0A",X"73",X"36",X"00",X"23",X"10",X"FB",X"06",X"3C",X"21",X"6E",
		X"73",X"36",X"00",X"23",X"10",X"FB",X"21",X"39",X"07",X"22",X"FA",X"70",X"CD",X"E0",X"40",X"CD",
		X"2D",X"3F",X"DD",X"21",X"AC",X"88",X"0E",X"38",X"06",X"13",X"CD",X"F1",X"3D",X"CD",X"9A",X"3F",
		X"CD",X"75",X"3F",X"CD",X"09",X"06",X"3A",X"32",X"70",X"2F",X"CB",X"57",X"C2",X"4A",X"07",X"3A",
		X"05",X"70",X"FE",X"00",X"20",X"07",X"3A",X"04",X"70",X"FE",X"01",X"28",X"E0",X"3A",X"33",X"70",
		X"2F",X"CB",X"57",X"C2",X"64",X"07",X"C3",X"DD",X"05",X"3A",X"F9",X"70",X"FE",X"00",X"C0",X"ED",
		X"4B",X"FA",X"70",X"3A",X"32",X"70",X"2F",X"21",X"FC",X"70",X"5F",X"AE",X"73",X"A3",X"CB",X"5F",
		X"C2",X"49",X"06",X"CB",X"67",X"C2",X"44",X"06",X"CB",X"6F",X"C2",X"3F",X"06",X"CB",X"77",X"C2",
		X"3A",X"06",X"CB",X"7F",X"C8",X"1E",X"08",X"C3",X"4B",X"06",X"1E",X"D3",X"C3",X"4B",X"06",X"1E",
		X"3E",X"C3",X"4B",X"06",X"1E",X"38",X"C3",X"4B",X"06",X"1E",X"09",X"0A",X"FE",X"C9",X"CA",X"61",
		X"06",X"BB",X"C2",X"5B",X"06",X"03",X"ED",X"43",X"FA",X"70",X"C9",X"3E",X"01",X"32",X"F9",X"70",
		X"C9",X"CD",X"E0",X"40",X"DD",X"21",X"D3",X"06",X"21",X"04",X"8B",X"CD",X"B7",X"06",X"DD",X"21",
		X"E4",X"06",X"21",X"26",X"8A",X"CD",X"B7",X"06",X"DD",X"21",X"E7",X"06",X"21",X"C8",X"8A",X"CD",
		X"B7",X"06",X"DD",X"21",X"F5",X"06",X"21",X"CA",X"8A",X"CD",X"B7",X"06",X"DD",X"21",X"03",X"07",
		X"21",X"CC",X"8A",X"CD",X"B7",X"06",X"DD",X"21",X"0E",X"07",X"21",X"CE",X"8A",X"CD",X"B7",X"06",
		X"DD",X"21",X"1D",X"07",X"21",X"D0",X"8A",X"CD",X"B7",X"06",X"DD",X"21",X"2C",X"07",X"21",X"D3",
		X"8A",X"CD",X"B7",X"06",X"C3",X"B4",X"06",X"01",X"20",X"00",X"11",X"00",X"10",X"DD",X"7E",X"00",
		X"FE",X"FF",X"C8",X"3D",X"3D",X"77",X"E5",X"19",X"36",X"0C",X"E1",X"97",X"ED",X"42",X"DD",X"23",
		X"C3",X"BD",X"06",X"0F",X"12",X"15",X"21",X"22",X"2B",X"24",X"1B",X"19",X"1A",X"26",X"12",X"03",
		X"0B",X"0A",X"05",X"FF",X"14",X"2B",X"FF",X"1B",X"26",X"1B",X"25",X"13",X"12",X"22",X"13",X"1E",
		X"13",X"1F",X"21",X"25",X"FF",X"22",X"24",X"21",X"19",X"24",X"13",X"1F",X"13",X"16",X"21",X"24",
		X"17",X"25",X"FF",X"1A",X"17",X"20",X"1D",X"12",X"25",X"22",X"1B",X"26",X"25",X"FF",X"1C",X"21",
		X"25",X"17",X"22",X"12",X"1F",X"2F",X"12",X"22",X"17",X"26",X"1B",X"26",X"FF",X"1C",X"21",X"25",
		X"17",X"22",X"12",X"1F",X"21",X"24",X"1B",X"1E",X"1E",X"13",X"25",X"FF",X"21",X"15",X"26",X"27",
		X"14",X"24",X"17",X"12",X"03",X"0B",X"0A",X"05",X"FF",X"08",X"D3",X"08",X"3E",X"38",X"D3",X"09",
		X"3E",X"08",X"D3",X"08",X"3E",X"D3",X"D3",X"09",X"08",X"C9",X"3E",X"02",X"32",X"11",X"75",X"AF",
		X"32",X"5D",X"70",X"3E",X"01",X"32",X"F9",X"70",X"3A",X"34",X"70",X"32",X"70",X"70",X"CD",X"83",
		X"07",X"C3",X"91",X"07",X"3E",X"02",X"32",X"11",X"75",X"3E",X"01",X"32",X"5D",X"70",X"32",X"F9",
		X"70",X"3A",X"34",X"70",X"32",X"70",X"70",X"32",X"71",X"70",X"CD",X"83",X"07",X"CD",X"83",X"07",
		X"C3",X"91",X"07",X"21",X"04",X"70",X"AF",X"BE",X"28",X"02",X"35",X"C9",X"36",X"09",X"23",X"35",
		X"C9",X"3A",X"00",X"A8",X"2F",X"E6",X"18",X"FE",X"00",X"28",X"13",X"FE",X"10",X"28",X"1A",X"FE",
		X"08",X"28",X"21",X"CD",X"3F",X"08",X"3E",X"02",X"32",X"66",X"73",X"C3",X"81",X"30",X"CD",X"CF",
		X"07",X"3E",X"03",X"32",X"66",X"73",X"C3",X"81",X"30",X"CD",X"07",X"08",X"3E",X"03",X"32",X"66",
		X"73",X"C3",X"81",X"30",X"CD",X"3F",X"08",X"3E",X"03",X"32",X"66",X"73",X"C3",X"81",X"30",X"21",
		X"28",X"23",X"22",X"50",X"73",X"22",X"46",X"73",X"21",X"F8",X"2A",X"22",X"48",X"73",X"21",X"F8",
		X"2A",X"22",X"4C",X"73",X"22",X"4E",X"73",X"3E",X"1A",X"32",X"61",X"73",X"32",X"B2",X"70",X"3E",
		X"1A",X"32",X"AF",X"70",X"32",X"65",X"73",X"3E",X"18",X"32",X"55",X"73",X"3E",X"1A",X"32",X"5A",
		X"73",X"3E",X"1C",X"32",X"5F",X"73",X"C9",X"21",X"34",X"21",X"22",X"50",X"73",X"22",X"46",X"73",
		X"21",X"04",X"29",X"22",X"48",X"73",X"21",X"F8",X"2A",X"22",X"4C",X"73",X"22",X"4E",X"73",X"3E",
		X"18",X"32",X"61",X"73",X"32",X"B2",X"70",X"3E",X"18",X"32",X"AF",X"70",X"32",X"65",X"73",X"3E",
		X"16",X"32",X"55",X"73",X"3E",X"18",X"32",X"5A",X"73",X"3E",X"1A",X"32",X"5F",X"73",X"C9",X"21",
		X"40",X"1F",X"22",X"50",X"73",X"22",X"46",X"73",X"21",X"10",X"27",X"22",X"48",X"73",X"21",X"F8",
		X"2A",X"22",X"4C",X"73",X"22",X"4E",X"73",X"3E",X"16",X"32",X"61",X"73",X"32",X"B2",X"70",X"3E",
		X"16",X"32",X"AF",X"70",X"32",X"65",X"73",X"3E",X"14",X"32",X"55",X"73",X"3E",X"16",X"32",X"5A",
		X"73",X"3E",X"18",X"32",X"5F",X"73",X"C9",X"AF",X"32",X"94",X"70",X"32",X"9F",X"70",X"32",X"AA",
		X"70",X"32",X"87",X"70",X"32",X"87",X"70",X"32",X"88",X"70",X"32",X"89",X"70",X"32",X"49",X"70",
		X"32",X"DA",X"70",X"32",X"E5",X"70",X"3E",X"20",X"32",X"0A",X"74",X"32",X"1A",X"74",X"3C",X"32",
		X"0E",X"74",X"32",X"1E",X"74",X"3C",X"32",X"12",X"74",X"32",X"22",X"74",X"3C",X"32",X"16",X"74",
		X"32",X"26",X"74",X"3E",X"2C",X"32",X"0B",X"74",X"32",X"0F",X"74",X"32",X"13",X"74",X"32",X"17",
		X"74",X"3E",X"24",X"32",X"1B",X"74",X"32",X"1F",X"74",X"32",X"23",X"74",X"32",X"27",X"74",X"3E",
		X"78",X"32",X"0C",X"74",X"32",X"1C",X"74",X"3E",X"D8",X"32",X"0D",X"74",X"32",X"1D",X"74",X"21",
		X"F7",X"09",X"22",X"D4",X"70",X"21",X"23",X"0C",X"22",X"DF",X"70",X"21",X"01",X"00",X"22",X"D6",
		X"70",X"22",X"E1",X"70",X"22",X"D8",X"70",X"22",X"E3",X"70",X"AF",X"32",X"DA",X"70",X"32",X"E5",
		X"70",X"32",X"D0",X"70",X"32",X"D2",X"70",X"32",X"DB",X"70",X"32",X"DD",X"70",X"C9",X"CD",X"1A",
		X"09",X"CD",X"6B",X"09",X"CD",X"47",X"0B",X"C3",X"97",X"0B",X"3A",X"DA",X"70",X"B7",X"C0",X"2A",
		X"D6",X"70",X"2B",X"22",X"D6",X"70",X"7C",X"B5",X"C0",X"21",X"00",X"03",X"22",X"D6",X"70",X"CD",
		X"A7",X"09",X"32",X"0C",X"74",X"32",X"14",X"74",X"C6",X"10",X"32",X"10",X"74",X"3D",X"32",X"18",
		X"74",X"AF",X"32",X"D0",X"70",X"CD",X"C5",X"09",X"32",X"0D",X"74",X"32",X"11",X"74",X"C6",X"10",
		X"32",X"15",X"74",X"32",X"19",X"74",X"AF",X"32",X"D2",X"70",X"2A",X"D4",X"70",X"7E",X"32",X"D0",
		X"70",X"23",X"7E",X"32",X"D2",X"70",X"23",X"22",X"D4",X"70",X"C9",X"3A",X"DA",X"70",X"B7",X"C2",
		X"E5",X"09",X"2A",X"D8",X"70",X"2B",X"22",X"D8",X"70",X"7C",X"B5",X"C0",X"21",X"74",X"01",X"22",
		X"D8",X"70",X"3A",X"0A",X"74",X"FE",X"20",X"28",X"16",X"FE",X"24",X"28",X"16",X"3E",X"20",X"32",
		X"0A",X"74",X"3C",X"32",X"0E",X"74",X"3C",X"32",X"12",X"74",X"3C",X"32",X"16",X"74",X"C9",X"3E",
		X"24",X"18",X"EC",X"3E",X"28",X"18",X"E8",X"3A",X"0C",X"74",X"5F",X"3A",X"D0",X"70",X"FE",X"03",
		X"CA",X"DE",X"09",X"FE",X"00",X"28",X"08",X"FE",X"01",X"28",X"06",X"7B",X"D6",X"03",X"C9",X"7B",
		X"C9",X"7B",X"C6",X"03",X"C9",X"3A",X"0D",X"74",X"5F",X"3A",X"D2",X"70",X"FE",X"00",X"28",X"08",
		X"FE",X"01",X"28",X"06",X"7B",X"D6",X"03",X"C9",X"7B",X"C9",X"7B",X"C6",X"03",X"C9",X"DD",X"E1",
		X"3E",X"01",X"32",X"DA",X"70",X"2A",X"D8",X"70",X"2B",X"7C",X"B5",X"20",X"06",X"CD",X"82",X"09",
		X"21",X"B0",X"03",X"22",X"D8",X"70",X"C9",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"01",X"02",X"01",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"01",
		X"02",X"01",X"02",X"01",X"02",X"01",X"02",X"01",X"01",X"01",X"01",X"01",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"01",X"02",X"01",X"02",X"01",X"02",X"01",X"02",X"01",X"02",X"01",X"02",X"01",
		X"02",X"01",X"02",X"01",X"02",X"01",X"02",X"01",X"02",X"01",X"02",X"01",X"02",X"01",X"02",X"01",
		X"02",X"01",X"02",X"01",X"02",X"01",X"02",X"01",X"01",X"01",X"02",X"01",X"02",X"01",X"02",X"01",
		X"02",X"01",X"01",X"01",X"02",X"01",X"02",X"01",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"01",
		X"02",X"01",X"02",X"01",X"02",X"01",X"01",X"01",X"02",X"01",X"02",X"01",X"02",X"01",X"01",X"01",
		X"02",X"01",X"02",X"01",X"02",X"01",X"02",X"02",X"01",X"02",X"01",X"02",X"01",X"02",X"01",X"02",
		X"02",X"02",X"01",X"02",X"01",X"02",X"01",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"01",X"02",X"01",X"02",X"01",X"02",X"01",X"02",X"02",X"02",X"01",X"02",X"01",X"01",X"01",X"02",
		X"01",X"02",X"01",X"02",X"02",X"01",X"01",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"01",
		X"01",X"02",X"02",X"02",X"02",X"02",X"02",X"01",X"01",X"02",X"01",X"02",X"01",X"02",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"01",X"01",X"02",X"01",X"01",X"01",X"01",X"01",X"01",
		X"02",X"01",X"01",X"00",X"01",X"00",X"01",X"01",X"02",X"01",X"02",X"01",X"02",X"01",X"02",X"01",
		X"02",X"02",X"01",X"01",X"01",X"02",X"01",X"02",X"01",X"02",X"01",X"02",X"01",X"02",X"01",X"02",
		X"01",X"02",X"01",X"02",X"01",X"02",X"01",X"01",X"01",X"02",X"02",X"02",X"01",X"02",X"01",X"02",
		X"01",X"02",X"01",X"02",X"01",X"01",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"00",X"00",X"00",X"01",X"00",X"00",X"02",X"00",X"00",X"01",X"02",X"02",X"02",X"02",X"02",
		X"01",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"01",X"02",X"02",X"01",X"02",
		X"02",X"02",X"02",X"02",X"03",X"03",X"03",X"3A",X"E5",X"70",X"B7",X"C0",X"2A",X"E1",X"70",X"2B",
		X"22",X"E1",X"70",X"7C",X"B5",X"C0",X"21",X"70",X"02",X"22",X"E1",X"70",X"CD",X"D3",X"0B",X"32",
		X"1C",X"74",X"32",X"24",X"74",X"C6",X"10",X"32",X"20",X"74",X"32",X"28",X"74",X"AF",X"32",X"DB",
		X"70",X"CD",X"F1",X"0B",X"32",X"1D",X"74",X"32",X"21",X"74",X"C6",X"10",X"32",X"25",X"74",X"32",
		X"29",X"74",X"AF",X"32",X"DD",X"70",X"2A",X"DF",X"70",X"7E",X"32",X"DB",X"70",X"23",X"7E",X"32",
		X"DD",X"70",X"23",X"22",X"DF",X"70",X"C9",X"3A",X"E5",X"70",X"B7",X"C2",X"11",X"0C",X"2A",X"E3",
		X"70",X"2B",X"22",X"E3",X"70",X"7C",X"B5",X"C0",X"21",X"70",X"01",X"22",X"E3",X"70",X"3A",X"1A",
		X"74",X"FE",X"20",X"28",X"16",X"FE",X"24",X"28",X"16",X"3E",X"20",X"32",X"1A",X"74",X"3C",X"32",
		X"1E",X"74",X"3C",X"32",X"22",X"74",X"3C",X"32",X"26",X"74",X"C9",X"3E",X"24",X"18",X"EC",X"3E",
		X"28",X"18",X"E8",X"3A",X"1C",X"74",X"5F",X"3A",X"DB",X"70",X"FE",X"03",X"CA",X"0A",X"0C",X"FE",
		X"00",X"28",X"08",X"FE",X"01",X"28",X"06",X"7B",X"D6",X"03",X"C9",X"7B",X"C9",X"7B",X"C6",X"03",
		X"C9",X"3A",X"1D",X"74",X"5F",X"3A",X"DD",X"70",X"FE",X"00",X"28",X"08",X"FE",X"01",X"28",X"06",
		X"7B",X"D6",X"03",X"C9",X"7B",X"C9",X"7B",X"C6",X"03",X"C9",X"DD",X"E1",X"3E",X"01",X"32",X"E5",
		X"70",X"2A",X"E3",X"70",X"2B",X"7C",X"B5",X"20",X"06",X"CD",X"AE",X"0B",X"21",X"00",X"03",X"22",
		X"E3",X"70",X"C9",X"01",X"02",X"01",X"02",X"01",X"02",X"01",X"02",X"01",X"02",X"01",X"02",X"01",
		X"01",X"01",X"01",X"01",X"02",X"01",X"02",X"01",X"02",X"01",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"01",X"02",X"01",X"02",X"02",X"01",X"02",X"01",X"02",X"01",X"02",X"01",
		X"02",X"01",X"02",X"01",X"02",X"01",X"02",X"01",X"02",X"01",X"02",X"01",X"02",X"01",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"01",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"01",X"02",
		X"02",X"02",X"02",X"02",X"02",X"01",X"02",X"01",X"02",X"01",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"01",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"01",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"02",X"01",X"02",X"01",X"02",X"01",X"02",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"02",X"01",X"01",X"01",X"01",X"02",X"01",X"01",X"01",X"01",X"01",X"01",
		X"02",X"02",X"01",X"01",X"02",X"01",X"02",X"01",X"02",X"01",X"02",X"02",X"01",X"01",X"02",X"01",
		X"02",X"01",X"02",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"01",X"02",X"01",X"02",
		X"01",X"02",X"02",X"02",X"01",X"01",X"01",X"02",X"01",X"02",X"01",X"02",X"02",X"02",X"01",X"00",
		X"01",X"00",X"01",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"01",X"01",X"02",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"02",X"01",X"01",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"02",X"02",X"01",X"02",X"01",X"02",X"01",X"02",X"01",X"02",X"01",X"02",X"00",X"00",X"00",
		X"01",X"00",X"00",X"01",X"00",X"00",X"01",X"00",X"02",X"00",X"02",X"00",X"01",X"00",X"02",X"00",
		X"02",X"01",X"02",X"01",X"02",X"01",X"02",X"02",X"02",X"01",X"01",X"01",X"02",X"01",X"02",X"01",
		X"03",X"03",X"03",X"ED",X"5F",X"FE",X"0C",X"30",X"04",X"21",X"C1",X"0D",X"C9",X"FE",X"18",X"30",
		X"04",X"21",X"FD",X"0D",X"C9",X"FE",X"24",X"30",X"04",X"21",X"39",X"0E",X"C9",X"FE",X"30",X"30",
		X"04",X"21",X"75",X"0E",X"C9",X"FE",X"3C",X"30",X"04",X"21",X"B1",X"0E",X"C9",X"FE",X"48",X"30",
		X"04",X"21",X"ED",X"0E",X"C9",X"FE",X"54",X"30",X"04",X"21",X"29",X"0F",X"C9",X"FE",X"60",X"30",
		X"04",X"21",X"65",X"0F",X"C9",X"FE",X"6C",X"30",X"04",X"21",X"A1",X"0F",X"C9",X"21",X"DD",X"0F",
		X"C9",X"E2",X"E2",X"E6",X"F9",X"DE",X"E2",X"E6",X"E6",X"CE",X"DE",X"CE",X"CA",X"E6",X"E6",X"DE",
		X"CE",X"DA",X"DA",X"DA",X"C6",X"E2",X"E6",X"DE",X"E6",X"CA",X"F9",X"E6",X"E6",X"E6",X"DE",X"E2",
		X"E2",X"D2",X"E6",X"CA",X"E2",X"E6",X"E2",X"D6",X"DE",X"D2",X"D6",X"D2",X"D6",X"CA",X"E2",X"E2",
		X"E2",X"E2",X"CA",X"E2",X"E6",X"E6",X"D6",X"DE",X"E2",X"E2",X"CA",X"E6",X"DE",X"F9",X"E6",X"E6",
		X"E6",X"C6",X"E2",X"E2",X"E2",X"E6",X"DE",X"E2",X"E6",X"DA",X"D6",X"DE",X"CE",X"CE",X"C6",X"DA",
		X"C6",X"CE",X"E6",X"DE",X"E6",X"DE",X"E2",X"DE",X"DE",X"E6",X"DE",X"CE",X"DE",X"E6",X"DE",X"DE",
		X"E2",X"E6",X"DE",X"E6",X"DE",X"D2",X"D6",X"D6",X"D6",X"CA",X"E2",X"D2",X"DE",X"CA",X"DE",X"F9",
		X"DE",X"E6",X"E6",X"DE",X"F9",X"DE",X"E6",X"D2",X"C6",X"E2",X"D6",X"E2",X"E6",X"DE",X"E2",X"E2",
		X"DE",X"DE",X"DE",X"E2",X"C6",X"E6",X"E6",X"DE",X"CE",X"DA",X"DA",X"DA",X"C6",X"D2",X"C6",X"DE",
		X"E6",X"DE",X"E2",X"E6",X"E6",X"E2",X"F9",X"E2",X"CA",X"E6",X"E6",X"DE",X"D2",X"E6",X"E6",X"D2",
		X"C6",X"D2",X"D6",X"D6",X"D6",X"CA",X"E2",X"D2",X"E6",X"E6",X"F9",X"E2",X"E6",X"CA",X"E6",X"F9",
		X"E2",X"CA",X"E6",X"E6",X"DE",X"E2",X"E6",X"B2",X"E6",X"DE",X"E2",X"E6",X"E6",X"E6",X"DE",X"E2",
		X"E6",X"B2",X"E6",X"DE",X"CE",X"DA",X"DA",X"DA",X"C6",X"E2",X"E6",X"DE",X"E6",X"DE",X"E2",X"E2",
		X"E2",X"E6",X"F9",X"E2",X"E6",X"E6",X"E6",X"DE",X"E2",X"D2",X"E6",X"CA",X"DE",X"D2",X"D6",X"D6",
		X"D6",X"CA",X"E2",X"E6",X"E6",X"CE",X"CA",X"E2",X"D2",X"C6",X"E6",X"DE",X"E2",X"E6",X"E6",X"E6",
		X"DE",X"E2",X"CE",X"E6",X"E2",X"CA",X"E2",X"E6",X"E6",X"DE",X"DE",X"E2",X"E2",X"E2",X"F9",X"DE",
		X"CE",X"DA",X"CE",X"DA",X"C6",X"E2",X"DE",X"E6",X"E6",X"DE",X"F9",X"E6",X"E6",X"D2",X"C6",X"E2",
		X"E6",X"E6",X"E6",X"DE",X"E2",X"F9",X"E6",X"E2",X"DE",X"D2",X"D6",X"D6",X"D6",X"CA",X"D2",X"DE",
		X"DE",X"DE",X"DE",X"D2",X"E6",X"E6",X"D2",X"DE",X"E2",X"DA",X"E6",X"C6",X"DE",X"E2",X"E6",X"F9",
		X"E6",X"DE",X"E2",X"DE",X"DE",X"E6",X"CA",X"E2",X"F9",X"E6",X"E6",X"DE",X"CE",X"DA",X"DA",X"B2",
		X"C6",X"E2",X"E6",X"E6",X"CA",X"DE",X"E2",X"D6",X"E6",X"DE",X"DE",X"E2",X"CA",X"E6",X"E6",X"C6",
		X"E2",X"E6",X"E6",X"E6",X"C6",X"D2",X"B2",X"D6",X"B2",X"CA",X"E2",X"E6",X"E6",X"E6",X"DE",X"D2",
		X"E6",X"DE",X"E6",X"DE",X"F9",X"E6",X"E2",X"E6",X"DE",X"E2",X"E6",X"DE",X"DE",X"DE",X"E2",X"E6",
		X"E2",X"E2",X"DE",X"D2",X"DE",X"E6",X"E6",X"DE",X"CE",X"DA",X"DA",X"CE",X"C6",X"E2",X"E6",X"DE",
		X"E6",X"DE",X"E2",X"CA",X"E6",X"DE",X"DE",X"E2",X"D6",X"E6",X"D6",X"DE",X"E2",X"DA",X"E6",X"CA",
		X"DE",X"D2",X"D6",X"D6",X"B2",X"CA",X"E2",X"E2",X"E2",X"E2",X"CA",X"E2",X"E6",X"E2",X"E6",X"DE",
		X"E2",X"E2",X"E6",X"D2",X"DE",X"E2",X"E6",X"E6",X"E6",X"DE",X"CE",X"E6",X"D6",X"E6",X"DE",X"E2",
		X"E6",X"DE",X"E6",X"CA",X"CE",X"DA",X"CE",X"C6",X"C6",X"CE",X"E6",X"E6",X"E6",X"CA",X"E2",X"E6",
		X"E6",X"E2",X"CA",X"D2",X"E2",X"DE",X"E6",X"F9",X"E2",X"DA",X"E6",X"CE",X"CA",X"D2",X"D2",X"D6",
		X"D2",X"CA",X"E2",X"E6",X"E2",X"E6",X"DE",X"D2",X"E2",X"E6",X"E2",X"CA",X"E2",X"DE",X"E6",X"D6",
		X"DE",X"E2",X"E6",X"E2",X"DE",X"DE",X"F9",X"D6",X"DE",X"E6",X"F9",X"E2",X"E6",X"DE",X"E6",X"C6",
		X"CE",X"B2",X"DA",X"DA",X"C6",X"E2",X"DE",X"E6",X"F9",X"DE",X"F9",X"DE",X"E6",X"E6",X"DE",X"E2",
		X"F9",X"DE",X"E6",X"DE",X"E2",X"E6",X"E6",X"E2",X"F9",X"D2",X"D6",X"D6",X"D6",X"CA",X"D2",X"E6",
		X"F9",X"E6",X"F9",X"E2",X"E2",X"E6",X"E6",X"DE",X"E2",X"E6",X"CA",X"E6",X"CA",X"E2",X"E6",X"E2",
		X"F9",X"DE",X"E2",X"E6",X"E6",X"E6",X"DE",X"E2",X"DE",X"DE",X"DE",X"DE",X"CE",X"DA",X"DA",X"DA",
		X"C6",X"E2",X"E6",X"D2",X"E6",X"DE",X"F9",X"E6",X"F9",X"E6",X"DE",X"E2",X"E6",X"E6",X"E6",X"CA",
		X"E2",X"CA",X"E6",X"D2",X"DE",X"D2",X"D6",X"D6",X"D6",X"CA",X"E2",X"E6",X"DE",X"E6",X"DE",X"D2",
		X"E6",X"DE",X"DE",X"DE",X"F9",X"E6",X"E2",X"E6",X"DE",X"CD",X"E0",X"40",X"CD",X"B2",X"10",X"0E",
		X"12",X"CD",X"4E",X"3E",X"11",X"88",X"42",X"21",X"E1",X"8A",X"0E",X"0B",X"CD",X"71",X"41",X"11",
		X"9A",X"42",X"21",X"F2",X"8A",X"0E",X"09",X"CD",X"71",X"41",X"11",X"AB",X"42",X"21",X"F4",X"8A",
		X"0E",X"09",X"CD",X"71",X"41",X"11",X"BC",X"42",X"21",X"56",X"8A",X"0E",X"09",X"CD",X"71",X"41",
		X"11",X"3B",X"42",X"21",X"FA",X"8A",X"0E",X"08",X"CD",X"71",X"41",X"3E",X"07",X"32",X"F0",X"70",
		X"21",X"50",X"00",X"22",X"EC",X"70",X"21",X"00",X"18",X"22",X"EE",X"70",X"2A",X"EC",X"70",X"2B",
		X"7D",X"B4",X"CA",X"AF",X"10",X"22",X"EC",X"70",X"3A",X"05",X"70",X"FE",X"00",X"C2",X"90",X"05",
		X"3A",X"04",X"70",X"FE",X"00",X"C2",X"90",X"05",X"2A",X"EE",X"70",X"2B",X"22",X"EE",X"70",X"7C",
		X"B5",X"20",X"E5",X"21",X"00",X"18",X"22",X"EE",X"70",X"3A",X"F0",X"70",X"EE",X"0F",X"32",X"F0",
		X"70",X"21",X"1A",X"99",X"11",X"20",X"00",X"06",X"10",X"77",X"19",X"10",X"FC",X"18",X"BD",X"C3",
		X"DB",X"04",X"CD",X"54",X"41",X"CD",X"6A",X"3F",X"11",X"79",X"42",X"21",X"44",X"8B",X"0E",X"07",
		X"CD",X"71",X"41",X"FD",X"21",X"AE",X"9A",X"DD",X"21",X"27",X"70",X"21",X"AE",X"8A",X"11",X"20",
		X"00",X"06",X"05",X"C5",X"E5",X"FD",X"E5",X"06",X"06",X"DD",X"7E",X"00",X"77",X"FD",X"36",X"00",
		X"0C",X"DD",X"2B",X"19",X"FD",X"19",X"10",X"F1",X"FD",X"E1",X"E1",X"C1",X"2B",X"2B",X"FD",X"2B",
		X"FD",X"2B",X"10",X"DF",X"FD",X"21",X"AE",X"98",X"DD",X"21",X"4F",X"72",X"21",X"AE",X"88",X"11",
		X"20",X"00",X"06",X"05",X"C5",X"E5",X"FD",X"E5",X"06",X"0E",X"DD",X"7E",X"00",X"77",X"FD",X"36",
		X"00",X"0C",X"DD",X"2B",X"19",X"FD",X"19",X"10",X"F1",X"FD",X"E1",X"E1",X"C1",X"2B",X"2B",X"FD",
		X"2B",X"FD",X"2B",X"10",X"DF",X"C9",X"CD",X"B2",X"10",X"11",X"E2",X"42",X"21",X"10",X"8B",X"0E",
		X"09",X"CD",X"71",X"41",X"11",X"F5",X"42",X"21",X"31",X"8B",X"0E",X"09",X"CD",X"71",X"41",X"11",
		X"C2",X"42",X"21",X"73",X"8A",X"0E",X"05",X"CD",X"71",X"41",X"11",X"CA",X"42",X"21",X"17",X"8B",
		X"0E",X"05",X"CD",X"71",X"41",X"11",X"DC",X"42",X"21",X"5B",X"8A",X"0E",X"05",X"CD",X"71",X"41",
		X"11",X"0A",X"43",X"21",X"3D",X"8B",X"0E",X"09",X"CD",X"71",X"41",X"3E",X"FF",X"32",X"15",X"8A",
		X"AF",X"32",X"19",X"8A",X"3C",X"32",X"57",X"8A",X"3C",X"32",X"D7",X"89",X"3E",X"15",X"32",X"15",
		X"9A",X"3E",X"35",X"32",X"19",X"9A",X"32",X"57",X"9A",X"32",X"D7",X"99",X"C9",X"16",X"01",X"DD",
		X"21",X"0A",X"70",X"2A",X"F1",X"70",X"06",X"06",X"4E",X"DD",X"7E",X"00",X"B9",X"DA",X"B9",X"11",
		X"C2",X"A8",X"11",X"2B",X"DD",X"23",X"10",X"F0",X"14",X"7A",X"FE",X"06",X"C8",X"AF",X"B8",X"CA",
		X"93",X"11",X"DD",X"23",X"10",X"FC",X"C3",X"93",X"11",X"00",X"7A",X"32",X"F3",X"70",X"FE",X"01",
		X"CA",X"D5",X"11",X"FE",X"02",X"CA",X"ED",X"11",X"FE",X"03",X"CA",X"02",X"12",X"FE",X"04",X"CA",
		X"14",X"12",X"C3",X"23",X"12",X"CD",X"42",X"12",X"CD",X"59",X"12",X"CD",X"70",X"12",X"CD",X"87",
		X"12",X"21",X"0A",X"72",X"CD",X"3A",X"12",X"11",X"0A",X"70",X"C3",X"2C",X"12",X"CD",X"42",X"12",
		X"CD",X"59",X"12",X"CD",X"70",X"12",X"21",X"18",X"72",X"CD",X"3A",X"12",X"11",X"10",X"70",X"C3",
		X"2C",X"12",X"CD",X"42",X"12",X"CD",X"59",X"12",X"21",X"26",X"72",X"CD",X"3A",X"12",X"11",X"16",
		X"70",X"C3",X"2C",X"12",X"CD",X"42",X"12",X"21",X"34",X"72",X"CD",X"3A",X"12",X"11",X"1C",X"70",
		X"C3",X"2C",X"12",X"21",X"42",X"72",X"CD",X"3A",X"12",X"11",X"22",X"70",X"2A",X"F1",X"70",X"06",
		X"06",X"7E",X"12",X"2B",X"13",X"10",X"FA",X"C3",X"9E",X"12",X"06",X"0E",X"36",X"10",X"23",X"10",
		X"FB",X"C9",X"21",X"1C",X"70",X"11",X"22",X"70",X"01",X"06",X"00",X"ED",X"B0",X"21",X"34",X"72",
		X"11",X"42",X"72",X"01",X"0E",X"00",X"ED",X"B0",X"C9",X"21",X"16",X"70",X"11",X"1C",X"70",X"01",
		X"06",X"00",X"ED",X"B0",X"21",X"26",X"72",X"11",X"34",X"72",X"01",X"0E",X"00",X"ED",X"B0",X"C9",
		X"21",X"10",X"70",X"11",X"16",X"70",X"01",X"06",X"00",X"ED",X"B0",X"21",X"18",X"72",X"11",X"26",
		X"72",X"01",X"0E",X"00",X"ED",X"B0",X"C9",X"21",X"0A",X"70",X"11",X"10",X"70",X"01",X"06",X"00",
		X"ED",X"B0",X"21",X"0A",X"72",X"11",X"18",X"72",X"01",X"0E",X"00",X"ED",X"B0",X"C9",X"CD",X"26",
		X"11",X"3A",X"F3",X"70",X"FE",X"01",X"CA",X"F0",X"12",X"FE",X"02",X"CA",X"E2",X"12",X"FE",X"03",
		X"CA",X"D4",X"12",X"FE",X"04",X"CA",X"C6",X"12",X"21",X"4E",X"8A",X"FD",X"21",X"42",X"72",X"DD",
		X"21",X"8D",X"88",X"C3",X"FB",X"12",X"21",X"4C",X"8A",X"FD",X"21",X"34",X"72",X"DD",X"21",X"8B",
		X"88",X"C3",X"FB",X"12",X"21",X"4A",X"8A",X"FD",X"21",X"26",X"72",X"DD",X"21",X"89",X"8A",X"C3",
		X"FB",X"12",X"21",X"48",X"8A",X"FD",X"21",X"18",X"72",X"DD",X"21",X"87",X"88",X"C3",X"FB",X"12",
		X"21",X"46",X"8A",X"FD",X"21",X"0A",X"72",X"DD",X"21",X"85",X"88",X"E5",X"FD",X"E5",X"0E",X"38",
		X"06",X"0E",X"CD",X"A2",X"3D",X"FD",X"E1",X"E1",X"3E",X"FA",X"32",X"F6",X"70",X"0E",X"00",X"06",
		X"11",X"11",X"20",X"00",X"70",X"FD",X"70",X"00",X"CD",X"87",X"13",X"3A",X"F6",X"70",X"3D",X"FE",
		X"00",X"28",X"7E",X"32",X"F6",X"70",X"3A",X"32",X"70",X"2F",X"CB",X"67",X"20",X"12",X"CB",X"5F",
		X"20",X"1E",X"CB",X"6F",X"20",X"29",X"CB",X"77",X"20",X"38",X"CB",X"7F",X"C0",X"C3",X"18",X"13",
		X"00",X"05",X"3E",X"0F",X"B8",X"DA",X"4A",X"13",X"06",X"2D",X"70",X"FD",X"70",X"00",X"18",X"C8",
		X"00",X"04",X"3E",X"2E",X"B8",X"30",X"02",X"06",X"10",X"70",X"FD",X"70",X"00",X"18",X"B9",X"79",
		X"FE",X"0D",X"28",X"B4",X"0C",X"97",X"ED",X"52",X"FD",X"23",X"06",X"11",X"70",X"FD",X"70",X"00",
		X"18",X"A6",X"79",X"FE",X"00",X"CA",X"18",X"13",X"0D",X"3E",X"10",X"FD",X"77",X"00",X"77",X"19",
		X"FD",X"2B",X"FD",X"46",X"00",X"18",X"91",X"C5",X"01",X"00",X"15",X"0B",X"F5",X"3A",X"32",X"70",
		X"2F",X"CB",X"7F",X"CA",X"99",X"13",X"01",X"00",X"00",X"CD",X"75",X"3F",X"F1",X"78",X"B1",X"20",
		X"EA",X"C1",X"C9",X"0E",X"0A",X"DD",X"21",X"40",X"88",X"DD",X"E5",X"11",X"00",X"10",X"06",X"09",
		X"DD",X"36",X"00",X"05",X"DD",X"36",X"01",X"03",X"DD",X"36",X"02",X"03",X"DD",X"36",X"03",X"05",
		X"DD",X"36",X"20",X"04",X"DD",X"36",X"23",X"04",X"DD",X"36",X"40",X"04",X"DD",X"36",X"43",X"04",
		X"DD",X"36",X"60",X"05",X"DD",X"36",X"61",X"03",X"DD",X"36",X"62",X"03",X"DD",X"36",X"63",X"05",
		X"DD",X"E5",X"DD",X"19",X"DD",X"36",X"00",X"30",X"DD",X"36",X"01",X"30",X"DD",X"36",X"02",X"30",
		X"DD",X"36",X"03",X"30",X"DD",X"36",X"20",X"30",X"DD",X"36",X"23",X"30",X"DD",X"36",X"40",X"30",
		X"DD",X"36",X"43",X"30",X"DD",X"36",X"60",X"30",X"DD",X"36",X"61",X"30",X"DD",X"36",X"62",X"30",
		X"DD",X"36",X"63",X"30",X"DD",X"E1",X"D5",X"11",X"60",X"00",X"DD",X"19",X"D1",X"10",X"91",X"DD",
		X"E1",X"DD",X"23",X"DD",X"23",X"DD",X"23",X"0D",X"C2",X"A9",X"13",X"3E",X"12",X"0E",X"12",X"DD",
		X"21",X"8D",X"89",X"CD",X"77",X"14",X"3E",X"38",X"0E",X"08",X"CD",X"77",X"14",X"3E",X"12",X"0E",
		X"17",X"DD",X"21",X"ED",X"89",X"CD",X"77",X"14",X"3E",X"36",X"0E",X"06",X"CD",X"77",X"14",X"3E",
		X"12",X"0E",X"22",X"DD",X"21",X"4D",X"8A",X"CD",X"77",X"14",X"3E",X"3B",X"0E",X"0B",X"CD",X"77",
		X"14",X"16",X"05",X"01",X"FF",X"FF",X"0B",X"78",X"B1",X"C2",X"66",X"14",X"0B",X"78",X"B1",X"C2",
		X"6C",X"14",X"15",X"C2",X"66",X"14",X"C9",X"11",X"00",X"10",X"DD",X"77",X"00",X"DD",X"77",X"01",
		X"DD",X"77",X"06",X"DD",X"77",X"07",X"DD",X"77",X"20",X"DD",X"77",X"21",X"DD",X"77",X"26",X"DD",
		X"77",X"27",X"DD",X"71",X"2A",X"DD",X"77",X"FB",X"DD",X"77",X"FA",X"DD",X"77",X"1A",X"DD",X"77",
		X"1B",X"DD",X"19",X"C9",X"CD",X"B0",X"14",X"CD",X"B0",X"18",X"CD",X"DA",X"14",X"C3",X"6F",X"15",
		X"3A",X"5E",X"70",X"FE",X"01",X"C8",X"3A",X"72",X"70",X"FE",X"00",X"CA",X"0B",X"15",X"2A",X"4A",
		X"73",X"2B",X"22",X"4A",X"73",X"7C",X"B5",X"20",X"31",X"AF",X"32",X"20",X"74",X"32",X"21",X"74",
		X"32",X"72",X"70",X"2A",X"4C",X"73",X"22",X"4E",X"73",X"C9",X"3A",X"5E",X"70",X"FE",X"01",X"CA",
		X"EE",X"14",X"3A",X"01",X"75",X"FE",X"01",X"C8",X"3E",X"06",X"32",X"11",X"75",X"C9",X"3A",X"01",
		X"75",X"FE",X"01",X"C8",X"3E",X"04",X"32",X"11",X"75",X"C9",X"7D",X"CB",X"7F",X"28",X"06",X"3E",
		X"04",X"32",X"1F",X"74",X"C9",X"3E",X"00",X"32",X"1F",X"74",X"C9",X"2A",X"4E",X"73",X"2B",X"22",
		X"4E",X"73",X"7C",X"B5",X"C0",X"3A",X"49",X"70",X"32",X"89",X"70",X"3A",X"CC",X"70",X"FE",X"01",
		X"C2",X"2A",X"15",X"3E",X"30",X"06",X"26",X"C3",X"54",X"15",X"ED",X"5F",X"FE",X"1E",X"D2",X"38",
		X"15",X"3E",X"30",X"06",X"24",X"C3",X"54",X"15",X"FE",X"3C",X"D2",X"44",X"15",X"3E",X"60",X"06",
		X"25",X"C3",X"54",X"15",X"FE",X"5A",X"D2",X"50",X"15",X"3E",X"90",X"06",X"26",X"C3",X"54",X"15",
		X"3E",X"C0",X"06",X"25",X"32",X"21",X"74",X"32",X"20",X"74",X"21",X"1E",X"74",X"70",X"2A",X"48",
		X"73",X"22",X"4A",X"73",X"3E",X"01",X"32",X"72",X"70",X"3E",X"08",X"32",X"1F",X"74",X"C9",X"3A",
		X"6F",X"70",X"B7",X"C2",X"B1",X"15",X"21",X"A0",X"9B",X"CD",X"01",X"16",X"3A",X"BE",X"70",X"B7",
		X"20",X"1D",X"06",X"06",X"21",X"79",X"70",X"11",X"C5",X"70",X"4E",X"1A",X"B9",X"38",X"06",X"C0",
		X"2B",X"13",X"10",X"F6",X"C9",X"3E",X"01",X"32",X"BE",X"70",X"AF",X"32",X"BF",X"70",X"C9",X"21",
		X"CA",X"70",X"11",X"74",X"70",X"06",X"06",X"1A",X"77",X"2B",X"13",X"10",X"FA",X"CD",X"EC",X"15",
		X"C9",X"21",X"40",X"99",X"CD",X"01",X"16",X"3A",X"BF",X"70",X"B7",X"20",X"1D",X"06",X"06",X"21",
		X"80",X"70",X"11",X"C5",X"70",X"4E",X"1A",X"B9",X"38",X"06",X"C0",X"2B",X"13",X"10",X"F6",X"C9",
		X"3E",X"01",X"32",X"BF",X"70",X"AF",X"32",X"BE",X"70",X"C9",X"21",X"CA",X"70",X"11",X"7B",X"70",
		X"06",X"06",X"1A",X"77",X"13",X"2B",X"10",X"FA",X"CD",X"EC",X"15",X"C9",X"21",X"A1",X"89",X"11",
		X"CA",X"70",X"06",X"06",X"1A",X"77",X"7D",X"C6",X"20",X"30",X"01",X"24",X"6F",X"1B",X"10",X"F4",
		X"C9",X"3A",X"EB",X"70",X"3D",X"32",X"EB",X"70",X"C0",X"97",X"11",X"20",X"00",X"06",X"09",X"3A",
		X"EA",X"70",X"77",X"ED",X"52",X"10",X"FB",X"3A",X"EA",X"70",X"EE",X"0C",X"32",X"EA",X"70",X"3E",
		X"FF",X"32",X"EB",X"70",X"C9",X"00",X"3A",X"AF",X"70",X"3D",X"32",X"AF",X"70",X"C0",X"3A",X"65",
		X"73",X"32",X"AF",X"70",X"CD",X"AB",X"16",X"21",X"19",X"74",X"3A",X"AE",X"70",X"B7",X"20",X"2E",
		X"34",X"3E",X"FE",X"BE",X"28",X"34",X"2B",X"34",X"3E",X"FE",X"BE",X"28",X"2D",X"3A",X"49",X"70",
		X"5F",X"3A",X"87",X"70",X"BB",X"C0",X"3A",X"24",X"74",X"BE",X"C0",X"3A",X"25",X"74",X"23",X"BE",
		X"30",X"06",X"3E",X"01",X"32",X"AE",X"70",X"C9",X"3E",X"02",X"32",X"AE",X"70",X"C9",X"3A",X"AE",
		X"70",X"FE",X"01",X"28",X"30",X"34",X"3E",X"FE",X"BE",X"C0",X"3A",X"87",X"70",X"FE",X"02",X"28",
		X"11",X"3C",X"32",X"87",X"70",X"AF",X"32",X"18",X"74",X"32",X"AE",X"70",X"ED",X"5F",X"32",X"19",
		X"74",X"C9",X"3A",X"16",X"74",X"EE",X"02",X"32",X"16",X"74",X"3A",X"17",X"74",X"EE",X"08",X"32",
		X"17",X"74",X"AF",X"18",X"DD",X"35",X"AF",X"BE",X"C0",X"18",X"CF",X"3A",X"B6",X"70",X"3D",X"20",
		X"0B",X"3A",X"16",X"74",X"EE",X"01",X"32",X"16",X"74",X"3A",X"B5",X"70",X"32",X"B6",X"70",X"C9",
		X"06",X"20",X"AF",X"10",X"FD",X"C9",X"3A",X"B2",X"70",X"3D",X"32",X"B2",X"70",X"FE",X"00",X"C2",
		X"A1",X"17",X"3A",X"61",X"73",X"32",X"B2",X"70",X"3A",X"C4",X"70",X"FE",X"00",X"CA",X"E5",X"16",
		X"3D",X"32",X"C4",X"70",X"C9",X"3A",X"B3",X"70",X"FE",X"00",X"CA",X"32",X"17",X"FE",X"08",X"28",
		X"09",X"21",X"1D",X"74",X"34",X"21",X"B3",X"70",X"35",X"C9",X"21",X"49",X"70",X"3A",X"88",X"70",
		X"BE",X"C2",X"2B",X"17",X"3A",X"B1",X"70",X"5F",X"16",X"00",X"21",X"26",X"18",X"19",X"7E",X"21",
		X"E2",X"89",X"19",X"FE",X"00",X"20",X"04",X"36",X"F8",X"18",X"0A",X"FE",X"01",X"20",X"04",X"36",
		X"F6",X"18",X"02",X"36",X"F7",X"11",X"00",X"10",X"19",X"36",X"12",X"21",X"B1",X"70",X"34",X"C3",
		X"F1",X"16",X"3A",X"B4",X"70",X"FE",X"00",X"28",X"3B",X"FE",X"08",X"28",X"09",X"21",X"1D",X"74",
		X"35",X"21",X"B4",X"70",X"35",X"C9",X"3A",X"B1",X"70",X"5F",X"16",X"00",X"21",X"26",X"18",X"19",
		X"7E",X"21",X"E2",X"89",X"19",X"FE",X"00",X"20",X"04",X"36",X"10",X"18",X"0A",X"FE",X"01",X"20",
		X"04",X"36",X"F9",X"18",X"02",X"36",X"FA",X"11",X"00",X"10",X"19",X"36",X"11",X"21",X"B1",X"70",
		X"35",X"C3",X"3D",X"17",X"2A",X"BA",X"70",X"7E",X"23",X"22",X"BA",X"70",X"FE",X"33",X"28",X"1A",
		X"FE",X"01",X"C2",X"8B",X"17",X"3E",X"08",X"32",X"B4",X"70",X"C9",X"FE",X"00",X"C2",X"96",X"17",
		X"3E",X"08",X"32",X"B3",X"70",X"C9",X"32",X"B2",X"70",X"C9",X"21",X"44",X"18",X"22",X"BA",X"70",
		X"C9",X"3A",X"BC",X"70",X"3D",X"20",X"0B",X"3A",X"1A",X"74",X"EE",X"01",X"32",X"1A",X"74",X"3A",
		X"BD",X"70",X"32",X"BC",X"70",X"C9",X"3A",X"C0",X"70",X"FE",X"01",X"C2",X"EC",X"17",X"11",X"26",
		X"18",X"21",X"E2",X"89",X"DD",X"21",X"E2",X"99",X"06",X"1C",X"1A",X"FE",X"00",X"20",X"04",X"36",
		X"10",X"18",X"0A",X"FE",X"01",X"20",X"04",X"36",X"F9",X"18",X"02",X"36",X"FA",X"DD",X"36",X"00",
		X"11",X"23",X"13",X"DD",X"23",X"10",X"E3",X"AF",X"32",X"C0",X"70",X"C9",X"3A",X"C1",X"70",X"FE",
		X"01",X"C0",X"3A",X"B1",X"70",X"FE",X"00",X"28",X"28",X"DD",X"21",X"E2",X"99",X"11",X"26",X"18",
		X"21",X"E2",X"89",X"47",X"1A",X"FE",X"00",X"20",X"04",X"36",X"F8",X"18",X"0A",X"FE",X"01",X"20",
		X"04",X"36",X"F6",X"18",X"02",X"36",X"F7",X"DD",X"36",X"00",X"12",X"DD",X"23",X"23",X"13",X"10",
		X"E3",X"AF",X"32",X"C1",X"70",X"C9",X"00",X"01",X"02",X"00",X"00",X"00",X"00",X"01",X"02",X"00",
		X"00",X"00",X"00",X"01",X"02",X"00",X"00",X"00",X"00",X"01",X"02",X"00",X"00",X"00",X"00",X"01",
		X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"0A",X"00",X"00",X"00",X"00",X"00",X"01",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"14",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"0A",X"01",X"01",X"01",X"01",
		X"00",X"01",X"01",X"01",X"00",X"01",X"01",X"01",X"00",X"01",X"01",X"01",X"01",X"01",X"0A",X"01",
		X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"01",X"01",X"01",X"00",X"01",X"00",X"01",X"01",X"14",
		X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"01",X"01",X"00",X"01",X"14",X"33",
		X"3A",X"00",X"A8",X"2F",X"E6",X"20",X"FE",X"20",X"CA",X"2D",X"19",X"3A",X"CC",X"70",X"FE",X"01",
		X"C8",X"3A",X"5E",X"70",X"FE",X"01",X"C8",X"3A",X"66",X"73",X"FE",X"00",X"C8",X"3A",X"32",X"70",
		X"2F",X"CB",X"7F",X"C8",X"3A",X"66",X"73",X"3D",X"32",X"66",X"73",X"3E",X"01",X"32",X"5E",X"70",
		X"21",X"AC",X"03",X"E7",X"CD",X"28",X"1F",X"3E",X"24",X"32",X"23",X"74",X"32",X"27",X"74",X"AF",
		X"32",X"0B",X"74",X"3E",X"05",X"32",X"0F",X"74",X"32",X"13",X"74",X"21",X"00",X"10",X"22",X"46",
		X"73",X"3E",X"04",X"32",X"11",X"75",X"CD",X"14",X"19",X"3A",X"66",X"73",X"FE",X"00",X"C8",X"47",
		X"3E",X"FE",X"18",X"04",X"3E",X"10",X"06",X"03",X"21",X"BF",X"8A",X"DD",X"21",X"BF",X"9A",X"11",
		X"20",X"00",X"77",X"DD",X"36",X"00",X"18",X"19",X"DD",X"19",X"10",X"F6",X"C9",X"3A",X"CC",X"70",
		X"FE",X"01",X"C8",X"3A",X"32",X"70",X"2F",X"CB",X"7F",X"CA",X"50",X"19",X"3A",X"0B",X"71",X"FE",
		X"00",X"C8",X"3A",X"67",X"73",X"3D",X"3D",X"3D",X"32",X"0A",X"71",X"AF",X"32",X"0B",X"71",X"C9",
		X"3A",X"0B",X"71",X"FE",X"01",X"C8",X"CD",X"14",X"19",X"3A",X"67",X"73",X"32",X"0A",X"71",X"3E",
		X"01",X"32",X"0B",X"71",X"C9",X"3A",X"54",X"73",X"3D",X"32",X"54",X"73",X"C0",X"3A",X"55",X"73",
		X"32",X"54",X"73",X"CD",X"EF",X"1B",X"3A",X"8C",X"70",X"FE",X"01",X"CA",X"48",X"1A",X"3A",X"92",
		X"70",X"FE",X"00",X"CA",X"22",X"1A",X"CD",X"E8",X"19",X"3A",X"5E",X"70",X"FE",X"01",X"CA",X"A1",
		X"19",X"3A",X"49",X"70",X"21",X"94",X"70",X"BE",X"CA",X"A1",X"19",X"DA",X"29",X"1B",X"C3",X"5D",
		X"1B",X"3A",X"0C",X"74",X"FE",X"30",X"C2",X"B6",X"19",X"3A",X"94",X"70",X"FE",X"00",X"C2",X"B6",
		X"19",X"3E",X"01",X"32",X"8F",X"70",X"3A",X"0C",X"74",X"FE",X"C0",X"C2",X"CB",X"19",X"3A",X"94",
		X"70",X"FE",X"02",X"C2",X"CB",X"19",X"3E",X"01",X"32",X"90",X"70",X"3A",X"0D",X"74",X"FE",X"18",
		X"C2",X"DB",X"19",X"3E",X"01",X"32",X"8D",X"70",X"C3",X"E5",X"19",X"FE",X"D8",X"C2",X"E5",X"19",
		X"3E",X"01",X"32",X"8E",X"70",X"C3",X"95",X"1A",X"3A",X"95",X"70",X"FE",X"FF",X"CA",X"1C",X"1A",
		X"FE",X"00",X"C2",X"FD",X"19",X"3E",X"01",X"32",X"8F",X"70",X"C3",X"1C",X"1A",X"FE",X"05",X"C2",
		X"0A",X"1A",X"3E",X"01",X"32",X"90",X"70",X"C3",X"1C",X"1A",X"FE",X"0A",X"C2",X"17",X"1A",X"3E",
		X"01",X"32",X"8D",X"70",X"C3",X"1C",X"1A",X"3E",X"01",X"32",X"8E",X"70",X"3E",X"FF",X"32",X"95",
		X"70",X"C9",X"3A",X"0C",X"74",X"FE",X"FF",X"CA",X"3B",X"1A",X"FE",X"00",X"C2",X"7B",X"1A",X"3E",
		X"FD",X"32",X"0C",X"74",X"21",X"94",X"70",X"35",X"C3",X"7B",X"1A",X"00",X"3E",X"02",X"32",X"0C",
		X"74",X"21",X"94",X"70",X"34",X"C3",X"7B",X"1A",X"AF",X"32",X"8C",X"70",X"3A",X"93",X"70",X"32",
		X"95",X"70",X"FE",X"00",X"20",X"08",X"3E",X"05",X"32",X"93",X"70",X"C3",X"7B",X"1A",X"FE",X"05",
		X"20",X"07",X"AF",X"32",X"93",X"70",X"C3",X"7B",X"1A",X"FE",X"0A",X"C2",X"76",X"1A",X"3E",X"0F",
		X"32",X"93",X"70",X"C3",X"7B",X"1A",X"3E",X"0A",X"32",X"93",X"70",X"21",X"0A",X"74",X"0E",X"14",
		X"3A",X"93",X"70",X"FE",X"00",X"CA",X"A0",X"1B",X"FE",X"05",X"CA",X"B0",X"1B",X"FE",X"0A",X"CA",
		X"C0",X"1B",X"C3",X"CF",X"1B",X"AF",X"32",X"92",X"70",X"3A",X"24",X"74",X"21",X"0C",X"74",X"BE",
		X"C2",X"15",X"1B",X"21",X"25",X"74",X"3A",X"0D",X"74",X"BE",X"DA",X"E1",X"1A",X"3A",X"5E",X"70",
		X"FE",X"01",X"CA",X"E9",X"1A",X"3A",X"8D",X"70",X"FE",X"01",X"CA",X"C5",X"1A",X"3E",X"0A",X"32",
		X"93",X"70",X"C3",X"7B",X"1A",X"3A",X"8F",X"70",X"FE",X"01",X"CA",X"D3",X"1A",X"32",X"93",X"70",
		X"C3",X"7B",X"1A",X"3A",X"90",X"70",X"FE",X"01",X"C8",X"3E",X"05",X"32",X"93",X"70",X"C3",X"7B",
		X"1A",X"3A",X"5E",X"70",X"FE",X"01",X"CA",X"B5",X"1A",X"3A",X"8E",X"70",X"FE",X"01",X"CA",X"F9",
		X"1A",X"3E",X"0F",X"32",X"93",X"70",X"C3",X"7B",X"1A",X"3A",X"90",X"70",X"FE",X"01",X"CA",X"09",
		X"1B",X"3E",X"05",X"32",X"93",X"70",X"C3",X"7B",X"1A",X"3A",X"8F",X"70",X"FE",X"01",X"C8",X"32",
		X"93",X"70",X"C3",X"7B",X"1A",X"21",X"0D",X"74",X"3A",X"25",X"74",X"BE",X"C2",X"93",X"1B",X"21",
		X"24",X"74",X"3A",X"0C",X"74",X"BE",X"DA",X"5D",X"1B",X"3A",X"5E",X"70",X"FE",X"01",X"CA",X"65",
		X"1B",X"3A",X"8F",X"70",X"FE",X"01",X"CA",X"3F",X"1B",X"32",X"93",X"70",X"C3",X"7B",X"1A",X"3A",
		X"8D",X"70",X"FE",X"01",X"CA",X"4F",X"1B",X"3E",X"0A",X"32",X"93",X"70",X"C3",X"7B",X"1A",X"3A",
		X"8E",X"70",X"FE",X"01",X"C8",X"3E",X"0F",X"32",X"93",X"70",X"C3",X"7B",X"1A",X"3A",X"5E",X"70",
		X"FE",X"01",X"CA",X"31",X"1B",X"3A",X"90",X"70",X"FE",X"01",X"CA",X"75",X"1B",X"3E",X"05",X"32",
		X"93",X"70",X"C3",X"7B",X"1A",X"3A",X"8E",X"70",X"FE",X"01",X"CA",X"85",X"1B",X"3E",X"0F",X"32",
		X"93",X"70",X"C3",X"7B",X"1A",X"3A",X"8D",X"70",X"FE",X"01",X"C8",X"3E",X"0A",X"32",X"93",X"70",
		X"C3",X"7B",X"1A",X"3A",X"25",X"74",X"21",X"0D",X"74",X"BE",X"DA",X"AD",X"1A",X"C3",X"E1",X"1A",
		X"7E",X"E6",X"01",X"0C",X"0C",X"B1",X"F6",X"80",X"77",X"CD",X"DE",X"1B",X"23",X"23",X"35",X"C9",
		X"7E",X"E6",X"01",X"0C",X"0C",X"B1",X"E6",X"3F",X"77",X"CD",X"DE",X"1B",X"23",X"23",X"34",X"C9",
		X"7E",X"E6",X"01",X"B1",X"E6",X"3F",X"77",X"CD",X"DE",X"1B",X"23",X"23",X"23",X"35",X"C9",X"7E",
		X"E6",X"01",X"B1",X"F6",X"C0",X"77",X"CD",X"DE",X"1B",X"23",X"23",X"23",X"34",X"C9",X"3A",X"52",
		X"73",X"3D",X"20",X"07",X"7E",X"EE",X"01",X"77",X"3A",X"53",X"73",X"32",X"52",X"73",X"C9",X"3A",
		X"93",X"70",X"FE",X"0A",X"CA",X"04",X"1C",X"FE",X"0F",X"CA",X"22",X"1C",X"FE",X"00",X"CA",X"40",
		X"1C",X"C3",X"5E",X"1C",X"3A",X"0D",X"74",X"06",X"05",X"21",X"98",X"1C",X"BE",X"CA",X"17",X"1D",
		X"23",X"10",X"F9",X"06",X"05",X"21",X"9D",X"1C",X"BE",X"CA",X"B8",X"1E",X"23",X"10",X"F9",X"C3",
		X"79",X"1C",X"3A",X"0D",X"74",X"06",X"05",X"21",X"8E",X"1C",X"BE",X"CA",X"17",X"1D",X"23",X"10",
		X"F9",X"06",X"05",X"21",X"93",X"1C",X"BE",X"CA",X"48",X"1E",X"23",X"10",X"F9",X"C3",X"79",X"1C",
		X"3A",X"0C",X"74",X"06",X"04",X"21",X"86",X"1C",X"BE",X"CA",X"17",X"1D",X"23",X"10",X"F9",X"06",
		X"04",X"21",X"8A",X"1C",X"BE",X"CA",X"68",X"1D",X"23",X"10",X"F9",X"C3",X"79",X"1C",X"3A",X"0C",
		X"74",X"06",X"04",X"21",X"7E",X"1C",X"BE",X"CA",X"17",X"1D",X"23",X"10",X"F9",X"06",X"04",X"21",
		X"82",X"1C",X"BE",X"CA",X"D8",X"1D",X"23",X"10",X"F9",X"AF",X"32",X"92",X"70",X"C9",X"20",X"50",
		X"80",X"B0",X"30",X"60",X"90",X"C0",X"D0",X"A0",X"70",X"40",X"C0",X"90",X"60",X"30",X"08",X"38",
		X"68",X"98",X"C8",X"18",X"48",X"78",X"A8",X"D8",X"28",X"58",X"88",X"B8",X"E8",X"18",X"48",X"78",
		X"A8",X"D8",X"ED",X"5B",X"93",X"70",X"16",X"00",X"21",X"EF",X"1C",X"19",X"06",X"05",X"3A",X"0D",
		X"74",X"0E",X"00",X"BE",X"CA",X"BB",X"1C",X"0C",X"23",X"10",X"F8",X"21",X"03",X"1D",X"19",X"06",
		X"05",X"3A",X"0C",X"74",X"BE",X"CA",X"D0",X"1C",X"23",X"0C",X"0C",X"0C",X"0C",X"0C",X"10",X"F4",
		X"79",X"32",X"8A",X"70",X"21",X"F6",X"72",X"3A",X"94",X"70",X"C6",X"01",X"47",X"11",X"14",X"00",
		X"19",X"10",X"FD",X"ED",X"5B",X"8A",X"70",X"16",X"00",X"19",X"7E",X"32",X"8B",X"70",X"C9",X"18",
		X"48",X"78",X"A8",X"D8",X"18",X"48",X"78",X"A8",X"D8",X"28",X"58",X"88",X"B8",X"E8",X"08",X"38",
		X"68",X"98",X"C8",X"D0",X"A0",X"70",X"40",X"00",X"B0",X"80",X"50",X"20",X"00",X"C0",X"90",X"60",
		X"30",X"00",X"C0",X"90",X"60",X"30",X"00",X"CD",X"A2",X"1C",X"3A",X"93",X"70",X"FE",X"00",X"20",
		X"06",X"21",X"5C",X"1D",X"C3",X"3E",X"1D",X"FE",X"05",X"20",X"06",X"21",X"58",X"1D",X"C3",X"3E",
		X"1D",X"FE",X"0A",X"20",X"06",X"21",X"60",X"1D",X"C3",X"3E",X"1D",X"21",X"64",X"1D",X"3A",X"8B",
		X"70",X"06",X"04",X"BE",X"CA",X"4F",X"1D",X"23",X"10",X"F9",X"AF",X"32",X"8C",X"70",X"C9",X"3E",
		X"01",X"32",X"92",X"70",X"32",X"8C",X"70",X"C9",X"C6",X"CE",X"DA",X"B2",X"CA",X"D2",X"D6",X"B2",
		X"C6",X"CA",X"DE",X"F9",X"CE",X"D2",X"E2",X"F9",X"3A",X"0C",X"74",X"21",X"8A",X"1C",X"06",X"05",
		X"BE",X"28",X"04",X"23",X"10",X"FA",X"C9",X"3E",X"01",X"32",X"92",X"70",X"AF",X"32",X"8D",X"70",
		X"32",X"8E",X"70",X"32",X"8F",X"70",X"32",X"90",X"70",X"3A",X"8B",X"70",X"FE",X"00",X"C8",X"FE",
		X"C6",X"C2",X"9D",X"1D",X"3E",X"01",X"32",X"8E",X"70",X"32",X"8F",X"70",X"C9",X"FE",X"CE",X"C2",
		X"AB",X"1D",X"3E",X"01",X"32",X"8D",X"70",X"32",X"8F",X"70",X"C9",X"FE",X"DA",X"C2",X"B6",X"1D",
		X"3E",X"01",X"32",X"8F",X"70",X"C9",X"FE",X"DE",X"C2",X"C1",X"1D",X"3E",X"01",X"32",X"8E",X"70",
		X"C9",X"FE",X"E2",X"C2",X"CC",X"1D",X"3E",X"01",X"32",X"8D",X"70",X"C9",X"FE",X"F9",X"C0",X"3E",
		X"01",X"32",X"8D",X"70",X"32",X"8E",X"70",X"C9",X"3A",X"0C",X"74",X"21",X"8A",X"1C",X"06",X"05",
		X"BE",X"28",X"04",X"23",X"10",X"FA",X"C9",X"3E",X"01",X"32",X"92",X"70",X"AF",X"32",X"8D",X"70",
		X"32",X"8E",X"70",X"32",X"8F",X"70",X"32",X"90",X"70",X"3A",X"8B",X"70",X"FE",X"00",X"C8",X"FE",
		X"CA",X"C2",X"0D",X"1E",X"3E",X"01",X"32",X"8E",X"70",X"32",X"90",X"70",X"C9",X"FE",X"D2",X"C2",
		X"1B",X"1E",X"3E",X"01",X"32",X"8D",X"70",X"32",X"90",X"70",X"C9",X"FE",X"D6",X"C2",X"26",X"1E",
		X"3E",X"01",X"32",X"90",X"70",X"C9",X"FE",X"DE",X"C2",X"31",X"1E",X"3E",X"01",X"32",X"8E",X"70",
		X"C9",X"FE",X"E2",X"C2",X"3C",X"1E",X"3E",X"01",X"32",X"8D",X"70",X"C9",X"FE",X"F9",X"C0",X"3E",
		X"01",X"32",X"8D",X"70",X"32",X"8E",X"70",X"C9",X"3A",X"0D",X"74",X"21",X"93",X"1C",X"06",X"05",
		X"BE",X"28",X"04",X"23",X"10",X"FA",X"C9",X"3E",X"01",X"32",X"92",X"70",X"AF",X"32",X"8D",X"70",
		X"32",X"8E",X"70",X"32",X"8F",X"70",X"32",X"90",X"70",X"3A",X"8B",X"70",X"FE",X"00",X"C8",X"FE",
		X"C6",X"C2",X"7D",X"1E",X"3E",X"01",X"32",X"8F",X"70",X"32",X"8E",X"70",X"C9",X"FE",X"CA",X"C2",
		X"8B",X"1E",X"3E",X"01",X"32",X"90",X"70",X"32",X"8E",X"70",X"C9",X"FE",X"D6",X"C2",X"96",X"1E",
		X"3E",X"01",X"32",X"90",X"70",X"C9",X"FE",X"DA",X"C2",X"A1",X"1E",X"3E",X"01",X"32",X"8F",X"70",
		X"C9",X"FE",X"DE",X"C2",X"AC",X"1E",X"3E",X"01",X"32",X"8E",X"70",X"C9",X"FE",X"B2",X"C0",X"3E",
		X"01",X"32",X"8F",X"70",X"32",X"90",X"70",X"C9",X"3A",X"0D",X"74",X"21",X"93",X"1C",X"06",X"05",
		X"BE",X"28",X"04",X"23",X"10",X"FA",X"C9",X"3E",X"01",X"32",X"92",X"70",X"AF",X"32",X"8D",X"70",
		X"32",X"8E",X"70",X"32",X"8F",X"70",X"32",X"90",X"70",X"3A",X"8B",X"70",X"FE",X"00",X"C8",X"FE",
		X"CE",X"C2",X"ED",X"1E",X"3E",X"01",X"32",X"8F",X"70",X"32",X"8D",X"70",X"C9",X"FE",X"D2",X"C2",
		X"FB",X"1E",X"3E",X"01",X"32",X"90",X"70",X"32",X"8D",X"70",X"C9",X"FE",X"D6",X"C2",X"06",X"1F",
		X"3E",X"01",X"32",X"90",X"70",X"C9",X"FE",X"DA",X"C2",X"11",X"1F",X"3E",X"01",X"32",X"8F",X"70",
		X"C9",X"FE",X"E2",X"C2",X"1C",X"1F",X"3E",X"01",X"32",X"8D",X"70",X"C9",X"FE",X"B2",X"C0",X"3E",
		X"01",X"32",X"8F",X"70",X"32",X"90",X"70",X"C9",X"00",X"3A",X"93",X"70",X"FE",X"00",X"20",X"08",
		X"3E",X"05",X"32",X"93",X"70",X"C3",X"55",X"1F",X"FE",X"05",X"20",X"07",X"AF",X"32",X"93",X"70",
		X"C3",X"55",X"1F",X"FE",X"0A",X"C2",X"50",X"1F",X"3E",X"0F",X"32",X"93",X"70",X"C3",X"55",X"1F",
		X"3E",X"0A",X"32",X"93",X"70",X"3A",X"9E",X"70",X"FE",X"00",X"20",X"08",X"3E",X"05",X"32",X"9E",
		X"70",X"C3",X"81",X"1F",X"FE",X"05",X"20",X"07",X"AF",X"32",X"9E",X"70",X"C3",X"81",X"1F",X"FE",
		X"0A",X"C2",X"7C",X"1F",X"3E",X"0F",X"32",X"9E",X"70",X"C3",X"81",X"1F",X"3E",X"0A",X"32",X"9E",
		X"70",X"3A",X"A9",X"70",X"FE",X"00",X"20",X"06",X"3E",X"05",X"32",X"A9",X"70",X"C9",X"FE",X"05",
		X"20",X"05",X"AF",X"32",X"A9",X"70",X"C9",X"FE",X"0A",X"C2",X"A2",X"1F",X"3E",X"0F",X"32",X"A9",
		X"70",X"C9",X"3E",X"0A",X"32",X"A9",X"70",X"C9",X"3A",X"58",X"73",X"3D",X"32",X"58",X"73",X"C0",
		X"3A",X"5A",X"73",X"32",X"58",X"73",X"CD",X"31",X"22",X"3A",X"98",X"70",X"FE",X"01",X"CA",X"8A",
		X"20",X"3A",X"9D",X"70",X"FE",X"00",X"CA",X"64",X"20",X"CD",X"2A",X"20",X"3A",X"5E",X"70",X"FE",
		X"01",X"28",X"10",X"3A",X"49",X"70",X"21",X"9F",X"70",X"BE",X"CA",X"E3",X"1F",X"DA",X"6B",X"21",
		X"C3",X"9F",X"21",X"3A",X"10",X"74",X"FE",X"30",X"C2",X"F8",X"1F",X"3A",X"9F",X"70",X"FE",X"00",
		X"C2",X"F8",X"1F",X"3E",X"01",X"32",X"9B",X"70",X"3A",X"10",X"74",X"FE",X"C0",X"C2",X"0D",X"20",
		X"3A",X"9F",X"70",X"FE",X"02",X"C2",X"0D",X"20",X"3E",X"01",X"32",X"9C",X"70",X"3A",X"11",X"74",
		X"FE",X"18",X"C2",X"1D",X"20",X"3E",X"01",X"32",X"99",X"70",X"C3",X"27",X"20",X"FE",X"D8",X"C2",
		X"27",X"20",X"3E",X"01",X"32",X"9A",X"70",X"C3",X"D7",X"20",X"3A",X"A0",X"70",X"FE",X"FF",X"CA",
		X"5E",X"20",X"FE",X"00",X"C2",X"3F",X"20",X"3E",X"01",X"32",X"9B",X"70",X"C3",X"5E",X"20",X"FE",
		X"05",X"C2",X"4C",X"20",X"3E",X"01",X"32",X"9C",X"70",X"C3",X"5E",X"20",X"FE",X"0A",X"C2",X"59",
		X"20",X"3E",X"01",X"32",X"99",X"70",X"C3",X"5E",X"20",X"3E",X"01",X"32",X"9A",X"70",X"3E",X"FF",
		X"32",X"A0",X"70",X"C9",X"3A",X"10",X"74",X"FE",X"FF",X"CA",X"7D",X"20",X"FE",X"00",X"C2",X"BD",
		X"20",X"3E",X"FD",X"32",X"10",X"74",X"21",X"9F",X"70",X"35",X"C3",X"BD",X"20",X"00",X"3E",X"02",
		X"32",X"10",X"74",X"21",X"9F",X"70",X"34",X"C3",X"BD",X"20",X"AF",X"32",X"98",X"70",X"3A",X"9E",
		X"70",X"32",X"A0",X"70",X"FE",X"00",X"20",X"08",X"3E",X"05",X"32",X"9E",X"70",X"C3",X"BD",X"20",
		X"FE",X"05",X"20",X"07",X"AF",X"32",X"9E",X"70",X"C3",X"BD",X"20",X"FE",X"0A",X"C2",X"B8",X"20",
		X"3E",X"0F",X"32",X"9E",X"70",X"C3",X"BD",X"20",X"3E",X"0A",X"32",X"9E",X"70",X"21",X"0E",X"74",
		X"0E",X"1C",X"3A",X"9E",X"70",X"FE",X"00",X"CA",X"E2",X"21",X"FE",X"05",X"CA",X"F2",X"21",X"FE",
		X"0A",X"CA",X"02",X"22",X"C3",X"11",X"22",X"AF",X"32",X"9D",X"70",X"3A",X"24",X"74",X"21",X"10",
		X"74",X"BE",X"C2",X"57",X"21",X"21",X"25",X"74",X"3A",X"11",X"74",X"BE",X"DA",X"23",X"21",X"3A",
		X"5E",X"70",X"FE",X"01",X"CA",X"2B",X"21",X"3A",X"99",X"70",X"FE",X"01",X"CA",X"07",X"21",X"3E",
		X"0A",X"32",X"9E",X"70",X"C3",X"BD",X"20",X"3A",X"9B",X"70",X"FE",X"01",X"CA",X"15",X"21",X"32",
		X"9E",X"70",X"C3",X"BD",X"20",X"3A",X"9C",X"70",X"FE",X"01",X"C8",X"3E",X"05",X"32",X"9E",X"70",
		X"C3",X"BD",X"20",X"3A",X"5E",X"70",X"FE",X"01",X"CA",X"F7",X"20",X"3A",X"9A",X"70",X"FE",X"01",
		X"CA",X"3B",X"21",X"3E",X"0F",X"32",X"9E",X"70",X"C3",X"BD",X"20",X"3A",X"9C",X"70",X"FE",X"01",
		X"CA",X"4B",X"21",X"3E",X"05",X"32",X"9E",X"70",X"C3",X"BD",X"20",X"3A",X"9B",X"70",X"FE",X"01",
		X"C8",X"32",X"9E",X"70",X"C3",X"BD",X"20",X"21",X"11",X"74",X"3A",X"25",X"74",X"BE",X"C2",X"D5",
		X"21",X"21",X"24",X"74",X"3A",X"10",X"74",X"BE",X"DA",X"9F",X"21",X"3A",X"5E",X"70",X"FE",X"01",
		X"CA",X"A7",X"21",X"3A",X"9B",X"70",X"FE",X"01",X"CA",X"81",X"21",X"32",X"9E",X"70",X"C3",X"BD",
		X"20",X"3A",X"99",X"70",X"FE",X"01",X"CA",X"91",X"21",X"3E",X"0A",X"32",X"9E",X"70",X"C3",X"BD",
		X"20",X"3A",X"9A",X"70",X"FE",X"01",X"C8",X"3E",X"0F",X"32",X"9E",X"70",X"C3",X"BD",X"20",X"3A",
		X"5E",X"70",X"FE",X"01",X"CA",X"73",X"21",X"3A",X"9C",X"70",X"FE",X"01",X"CA",X"B7",X"21",X"3E",
		X"05",X"32",X"9E",X"70",X"C3",X"BD",X"20",X"3A",X"9A",X"70",X"FE",X"01",X"CA",X"C7",X"21",X"3E",
		X"0F",X"32",X"9E",X"70",X"C3",X"BD",X"20",X"3A",X"99",X"70",X"FE",X"01",X"C8",X"3E",X"0A",X"32",
		X"9E",X"70",X"C3",X"BD",X"20",X"3A",X"10",X"74",X"21",X"24",X"74",X"BE",X"DA",X"9F",X"21",X"C3",
		X"6B",X"21",X"7E",X"E6",X"01",X"0C",X"0C",X"B1",X"F6",X"80",X"77",X"CD",X"20",X"22",X"23",X"23",
		X"35",X"C9",X"7E",X"E6",X"01",X"0C",X"0C",X"B1",X"E6",X"3F",X"77",X"CD",X"20",X"22",X"23",X"23",
		X"34",X"C9",X"7E",X"E6",X"01",X"B1",X"E6",X"3F",X"77",X"CD",X"20",X"22",X"23",X"23",X"23",X"35",
		X"C9",X"7E",X"E6",X"01",X"B1",X"F6",X"C0",X"77",X"CD",X"20",X"22",X"23",X"23",X"23",X"34",X"C9",
		X"3A",X"56",X"73",X"3D",X"20",X"07",X"7E",X"EE",X"01",X"77",X"3A",X"57",X"73",X"32",X"56",X"73",
		X"C9",X"3A",X"9E",X"70",X"FE",X"0A",X"CA",X"46",X"22",X"FE",X"0F",X"CA",X"64",X"22",X"FE",X"00",
		X"CA",X"82",X"22",X"C3",X"A0",X"22",X"3A",X"11",X"74",X"06",X"05",X"21",X"98",X"1C",X"BE",X"CA",
		X"0D",X"23",X"23",X"10",X"F9",X"06",X"05",X"21",X"9D",X"1C",X"BE",X"CA",X"9E",X"24",X"23",X"10",
		X"F9",X"C3",X"BB",X"22",X"3A",X"11",X"74",X"06",X"05",X"21",X"8E",X"1C",X"BE",X"CA",X"0D",X"23",
		X"23",X"10",X"F9",X"06",X"05",X"21",X"93",X"1C",X"BE",X"CA",X"2E",X"24",X"23",X"10",X"F9",X"C3",
		X"BB",X"22",X"3A",X"10",X"74",X"06",X"04",X"21",X"86",X"1C",X"BE",X"CA",X"0D",X"23",X"23",X"10",
		X"F9",X"06",X"04",X"21",X"8A",X"1C",X"BE",X"CA",X"4E",X"23",X"23",X"10",X"F9",X"C3",X"BB",X"22",
		X"3A",X"10",X"74",X"06",X"04",X"21",X"7E",X"1C",X"BE",X"CA",X"0D",X"23",X"23",X"10",X"F9",X"06",
		X"04",X"21",X"82",X"1C",X"BE",X"CA",X"BE",X"23",X"23",X"10",X"F9",X"AF",X"32",X"9D",X"70",X"C9",
		X"ED",X"5B",X"9E",X"70",X"16",X"00",X"21",X"EF",X"1C",X"19",X"06",X"05",X"3A",X"11",X"74",X"0E",
		X"00",X"BE",X"CA",X"D9",X"22",X"0C",X"23",X"10",X"F8",X"21",X"03",X"1D",X"19",X"06",X"05",X"3A",
		X"10",X"74",X"BE",X"CA",X"EE",X"22",X"23",X"0C",X"0C",X"0C",X"0C",X"0C",X"10",X"F4",X"79",X"32",
		X"96",X"70",X"21",X"F6",X"72",X"3A",X"9F",X"70",X"C6",X"01",X"47",X"11",X"14",X"00",X"19",X"10",
		X"FD",X"ED",X"5B",X"96",X"70",X"16",X"00",X"19",X"7E",X"32",X"97",X"70",X"C9",X"CD",X"C0",X"22",
		X"3A",X"9E",X"70",X"FE",X"00",X"20",X"06",X"21",X"5C",X"1D",X"C3",X"34",X"23",X"FE",X"05",X"20",
		X"06",X"21",X"58",X"1D",X"C3",X"34",X"23",X"FE",X"0A",X"20",X"06",X"21",X"60",X"1D",X"C3",X"34",
		X"23",X"21",X"64",X"1D",X"3A",X"97",X"70",X"06",X"04",X"BE",X"CA",X"45",X"23",X"23",X"10",X"F9",
		X"AF",X"32",X"98",X"70",X"C9",X"3E",X"01",X"32",X"9D",X"70",X"32",X"98",X"70",X"C9",X"3A",X"10",
		X"74",X"21",X"8A",X"1C",X"06",X"05",X"BE",X"28",X"04",X"23",X"10",X"FA",X"C9",X"3E",X"01",X"32",
		X"9D",X"70",X"AF",X"32",X"99",X"70",X"32",X"9A",X"70",X"32",X"9B",X"70",X"32",X"9C",X"70",X"3A",
		X"97",X"70",X"FE",X"00",X"C8",X"FE",X"C6",X"C2",X"83",X"23",X"3E",X"01",X"32",X"9A",X"70",X"32",
		X"9B",X"70",X"C9",X"FE",X"CE",X"C2",X"91",X"23",X"3E",X"01",X"32",X"99",X"70",X"32",X"9B",X"70",
		X"C9",X"FE",X"DA",X"C2",X"9C",X"23",X"3E",X"01",X"32",X"9B",X"70",X"C9",X"FE",X"DE",X"C2",X"A7",
		X"23",X"3E",X"01",X"32",X"9A",X"70",X"C9",X"FE",X"E2",X"C2",X"B2",X"23",X"3E",X"01",X"32",X"99",
		X"70",X"C9",X"FE",X"F9",X"C0",X"3E",X"01",X"32",X"99",X"70",X"32",X"9A",X"70",X"C9",X"3A",X"10",
		X"74",X"21",X"8A",X"1C",X"06",X"05",X"BE",X"28",X"04",X"23",X"10",X"FA",X"C9",X"3E",X"01",X"32",
		X"9D",X"70",X"AF",X"32",X"99",X"70",X"32",X"9A",X"70",X"32",X"9B",X"70",X"32",X"9C",X"70",X"3A",
		X"97",X"70",X"FE",X"00",X"C8",X"FE",X"CA",X"C2",X"F3",X"23",X"3E",X"01",X"32",X"9A",X"70",X"32",
		X"9C",X"70",X"C9",X"FE",X"D2",X"C2",X"01",X"24",X"3E",X"01",X"32",X"99",X"70",X"32",X"9C",X"70",
		X"C9",X"FE",X"D6",X"C2",X"0C",X"24",X"3E",X"01",X"32",X"9C",X"70",X"C9",X"FE",X"DE",X"C2",X"17",
		X"24",X"3E",X"01",X"32",X"9A",X"70",X"C9",X"FE",X"E2",X"C2",X"22",X"24",X"3E",X"01",X"32",X"99",
		X"70",X"C9",X"FE",X"F9",X"C0",X"3E",X"01",X"32",X"99",X"70",X"32",X"9A",X"70",X"C9",X"3A",X"11",
		X"74",X"21",X"93",X"1C",X"06",X"05",X"BE",X"28",X"04",X"23",X"10",X"FA",X"C9",X"3E",X"01",X"32",
		X"9D",X"70",X"AF",X"32",X"99",X"70",X"32",X"9A",X"70",X"32",X"9B",X"70",X"32",X"9C",X"70",X"3A",
		X"97",X"70",X"FE",X"00",X"C8",X"FE",X"C6",X"C2",X"63",X"24",X"3E",X"01",X"32",X"9B",X"70",X"32",
		X"9A",X"70",X"C9",X"FE",X"CA",X"C2",X"71",X"24",X"3E",X"01",X"32",X"9C",X"70",X"32",X"9A",X"70",
		X"C9",X"FE",X"D6",X"C2",X"7C",X"24",X"3E",X"01",X"32",X"9C",X"70",X"C9",X"FE",X"DA",X"C2",X"87",
		X"24",X"3E",X"01",X"32",X"9B",X"70",X"C9",X"FE",X"DE",X"C2",X"92",X"24",X"3E",X"01",X"32",X"9A",
		X"70",X"C9",X"FE",X"B2",X"C0",X"3E",X"01",X"32",X"9B",X"70",X"32",X"9C",X"70",X"C9",X"3A",X"11",
		X"74",X"21",X"93",X"1C",X"06",X"05",X"BE",X"28",X"04",X"23",X"10",X"FA",X"C9",X"3E",X"01",X"32",
		X"9D",X"70",X"AF",X"32",X"99",X"70",X"32",X"9A",X"70",X"32",X"9B",X"70",X"32",X"9C",X"70",X"3A",
		X"97",X"70",X"FE",X"00",X"C8",X"FE",X"CE",X"C2",X"D3",X"24",X"3E",X"01",X"32",X"9B",X"70",X"32",
		X"99",X"70",X"C9",X"FE",X"D2",X"C2",X"E1",X"24",X"3E",X"01",X"32",X"9C",X"70",X"32",X"99",X"70",
		X"C9",X"FE",X"D6",X"C2",X"EC",X"24",X"3E",X"01",X"32",X"9C",X"70",X"C9",X"FE",X"DA",X"C2",X"F7",
		X"24",X"3E",X"01",X"32",X"9B",X"70",X"C9",X"FE",X"E2",X"C2",X"02",X"25",X"3E",X"01",X"32",X"99",
		X"70",X"C9",X"FE",X"B2",X"C0",X"3E",X"01",X"32",X"9B",X"70",X"32",X"9C",X"70",X"C9",X"3A",X"5E",
		X"73",X"3D",X"32",X"5E",X"73",X"C0",X"3A",X"5F",X"73",X"32",X"5E",X"73",X"CD",X"4F",X"28",X"3A",
		X"A3",X"70",X"FE",X"01",X"CA",X"F1",X"25",X"3A",X"A8",X"70",X"FE",X"00",X"CA",X"CB",X"25",X"CD",
		X"91",X"25",X"3A",X"5E",X"70",X"FE",X"01",X"CA",X"4A",X"25",X"3A",X"49",X"70",X"21",X"AA",X"70",
		X"BE",X"CA",X"4A",X"25",X"DA",X"D2",X"26",X"C3",X"06",X"27",X"3A",X"14",X"74",X"FE",X"30",X"C2",
		X"5F",X"25",X"3A",X"AA",X"70",X"FE",X"00",X"C2",X"5F",X"25",X"3E",X"01",X"32",X"A6",X"70",X"3A",
		X"14",X"74",X"FE",X"C0",X"C2",X"74",X"25",X"3A",X"AA",X"70",X"FE",X"02",X"C2",X"74",X"25",X"3E",
		X"01",X"32",X"A7",X"70",X"3A",X"15",X"74",X"FE",X"18",X"C2",X"84",X"25",X"3E",X"01",X"32",X"A4",
		X"70",X"C3",X"8E",X"25",X"FE",X"D8",X"C2",X"8E",X"25",X"3E",X"01",X"32",X"A5",X"70",X"C3",X"3E",
		X"26",X"3A",X"AB",X"70",X"FE",X"FF",X"CA",X"C5",X"25",X"FE",X"00",X"C2",X"A6",X"25",X"3E",X"01",
		X"32",X"A6",X"70",X"C3",X"C5",X"25",X"FE",X"05",X"C2",X"B3",X"25",X"3E",X"01",X"32",X"A7",X"70",
		X"C3",X"C5",X"25",X"FE",X"0A",X"C2",X"C0",X"25",X"3E",X"01",X"32",X"A4",X"70",X"C3",X"C5",X"25",
		X"3E",X"01",X"32",X"A5",X"70",X"3E",X"FF",X"32",X"AB",X"70",X"C9",X"3A",X"14",X"74",X"FE",X"FF",
		X"CA",X"E4",X"25",X"FE",X"00",X"C2",X"24",X"26",X"3E",X"FD",X"32",X"14",X"74",X"21",X"AA",X"70",
		X"35",X"C3",X"24",X"26",X"00",X"3E",X"02",X"32",X"14",X"74",X"21",X"AA",X"70",X"34",X"C3",X"24",
		X"26",X"AF",X"32",X"A3",X"70",X"3A",X"A9",X"70",X"32",X"AB",X"70",X"FE",X"00",X"20",X"08",X"3E",
		X"05",X"32",X"A9",X"70",X"C3",X"24",X"26",X"FE",X"05",X"20",X"07",X"AF",X"32",X"A9",X"70",X"C3",
		X"24",X"26",X"FE",X"0A",X"C2",X"1F",X"26",X"3E",X"0F",X"32",X"A9",X"70",X"C3",X"24",X"26",X"3E",
		X"0A",X"32",X"A9",X"70",X"21",X"12",X"74",X"0E",X"0C",X"3A",X"A9",X"70",X"FE",X"00",X"CA",X"00",
		X"28",X"FE",X"05",X"CA",X"10",X"28",X"FE",X"0A",X"CA",X"20",X"28",X"C3",X"2F",X"28",X"AF",X"32",
		X"A8",X"70",X"3A",X"24",X"74",X"21",X"14",X"74",X"BE",X"C2",X"BE",X"26",X"21",X"25",X"74",X"3A",
		X"15",X"74",X"BE",X"DA",X"8A",X"26",X"3A",X"5E",X"70",X"FE",X"01",X"CA",X"92",X"26",X"3A",X"A4",
		X"70",X"FE",X"01",X"CA",X"6E",X"26",X"3E",X"0A",X"32",X"A9",X"70",X"C3",X"24",X"26",X"3A",X"A6",
		X"70",X"FE",X"01",X"CA",X"7C",X"26",X"32",X"A9",X"70",X"C3",X"24",X"26",X"3A",X"A7",X"70",X"FE",
		X"01",X"C8",X"3E",X"05",X"32",X"A9",X"70",X"C3",X"24",X"26",X"3A",X"5E",X"70",X"FE",X"01",X"CA",
		X"5E",X"26",X"3A",X"A5",X"70",X"FE",X"01",X"CA",X"A2",X"26",X"3E",X"0F",X"32",X"A9",X"70",X"C3",
		X"24",X"26",X"3A",X"A7",X"70",X"FE",X"01",X"CA",X"B2",X"26",X"3E",X"05",X"32",X"A9",X"70",X"C3",
		X"24",X"26",X"3A",X"A6",X"70",X"FE",X"01",X"C8",X"32",X"A9",X"70",X"C3",X"24",X"26",X"21",X"15",
		X"74",X"3A",X"25",X"74",X"BE",X"C2",X"3C",X"27",X"21",X"24",X"74",X"3A",X"14",X"74",X"BE",X"DA",
		X"06",X"27",X"3A",X"5E",X"70",X"FE",X"01",X"CA",X"0E",X"27",X"3A",X"A6",X"70",X"FE",X"01",X"CA",
		X"E8",X"26",X"32",X"A9",X"70",X"C3",X"24",X"26",X"3A",X"A4",X"70",X"FE",X"01",X"CA",X"F8",X"26",
		X"3E",X"0A",X"32",X"A9",X"70",X"C3",X"24",X"26",X"3A",X"A5",X"70",X"FE",X"01",X"C8",X"3E",X"0F",
		X"32",X"A9",X"70",X"C3",X"24",X"26",X"3A",X"5E",X"70",X"FE",X"01",X"CA",X"DA",X"26",X"3A",X"A7",
		X"70",X"FE",X"01",X"CA",X"1E",X"27",X"3E",X"05",X"32",X"A9",X"70",X"C3",X"24",X"26",X"3A",X"A5",
		X"70",X"FE",X"01",X"CA",X"2E",X"27",X"3E",X"0F",X"32",X"A9",X"70",X"C3",X"24",X"26",X"3A",X"A4",
		X"70",X"FE",X"01",X"C8",X"3E",X"0A",X"32",X"A9",X"70",X"C3",X"24",X"26",X"3A",X"A9",X"70",X"FE",
		X"00",X"C2",X"6F",X"27",X"3A",X"A4",X"70",X"FE",X"01",X"CA",X"54",X"27",X"3E",X"0A",X"32",X"A9",
		X"70",X"C3",X"24",X"26",X"3A",X"A5",X"70",X"FE",X"01",X"CA",X"64",X"27",X"3E",X"0F",X"32",X"A9",
		X"70",X"C3",X"24",X"26",X"3A",X"A6",X"70",X"FE",X"01",X"CA",X"F1",X"25",X"C3",X"24",X"26",X"3A",
		X"A9",X"70",X"FE",X"05",X"C2",X"A2",X"27",X"3A",X"A5",X"70",X"FE",X"01",X"CA",X"87",X"27",X"3E",
		X"0F",X"32",X"A9",X"70",X"C3",X"24",X"26",X"3A",X"A4",X"70",X"FE",X"01",X"CA",X"97",X"27",X"3E",
		X"0A",X"32",X"A9",X"70",X"C3",X"24",X"26",X"3A",X"A7",X"70",X"FE",X"01",X"CA",X"F1",X"25",X"C3",
		X"24",X"26",X"3A",X"A9",X"70",X"FE",X"0F",X"C2",X"D5",X"27",X"3A",X"A7",X"70",X"FE",X"01",X"CA",
		X"BA",X"27",X"3E",X"05",X"32",X"A9",X"70",X"C3",X"24",X"26",X"3A",X"A6",X"70",X"FE",X"01",X"CA",
		X"CA",X"27",X"3E",X"00",X"32",X"A9",X"70",X"C3",X"24",X"26",X"3A",X"A5",X"70",X"FE",X"01",X"CA",
		X"F1",X"25",X"C3",X"24",X"26",X"3A",X"A6",X"70",X"FE",X"01",X"CA",X"E5",X"27",X"3E",X"00",X"32",
		X"A9",X"70",X"C3",X"24",X"26",X"3A",X"A7",X"70",X"FE",X"01",X"CA",X"F5",X"27",X"3E",X"05",X"32",
		X"A9",X"70",X"C3",X"24",X"26",X"3A",X"A4",X"70",X"FE",X"01",X"CA",X"F1",X"25",X"C3",X"24",X"26",
		X"7E",X"E6",X"01",X"0C",X"0C",X"B1",X"F6",X"80",X"77",X"CD",X"3E",X"28",X"23",X"23",X"35",X"C9",
		X"7E",X"E6",X"01",X"0C",X"0C",X"B1",X"E6",X"3F",X"77",X"CD",X"3E",X"28",X"23",X"23",X"34",X"C9",
		X"7E",X"E6",X"01",X"B1",X"E6",X"3F",X"77",X"CD",X"3E",X"28",X"23",X"23",X"23",X"35",X"C9",X"7E",
		X"E6",X"01",X"B1",X"F6",X"C0",X"77",X"CD",X"3E",X"28",X"23",X"23",X"23",X"34",X"C9",X"3A",X"5C",
		X"73",X"3D",X"20",X"07",X"7E",X"EE",X"01",X"77",X"3A",X"5D",X"73",X"32",X"5C",X"73",X"C9",X"3A",
		X"A9",X"70",X"FE",X"0A",X"CA",X"64",X"28",X"FE",X"0F",X"CA",X"82",X"28",X"FE",X"00",X"CA",X"A0",
		X"28",X"C3",X"BE",X"28",X"3A",X"15",X"74",X"06",X"05",X"21",X"98",X"1C",X"BE",X"CA",X"2B",X"29",
		X"23",X"10",X"F9",X"06",X"05",X"21",X"9D",X"1C",X"BE",X"CA",X"BC",X"2A",X"23",X"10",X"F9",X"C3",
		X"D9",X"28",X"3A",X"15",X"74",X"06",X"05",X"21",X"8E",X"1C",X"BE",X"CA",X"2B",X"29",X"23",X"10",
		X"F9",X"06",X"05",X"21",X"93",X"1C",X"BE",X"CA",X"4C",X"2A",X"23",X"10",X"F9",X"C3",X"D9",X"28",
		X"3A",X"14",X"74",X"06",X"04",X"21",X"86",X"1C",X"BE",X"CA",X"2B",X"29",X"23",X"10",X"F9",X"06",
		X"04",X"21",X"8A",X"1C",X"BE",X"CA",X"6C",X"29",X"23",X"10",X"F9",X"C3",X"D9",X"28",X"3A",X"14",
		X"74",X"06",X"04",X"21",X"7E",X"1C",X"BE",X"CA",X"2B",X"29",X"23",X"10",X"F9",X"06",X"04",X"21",
		X"82",X"1C",X"BE",X"CA",X"DC",X"29",X"23",X"10",X"F9",X"AF",X"32",X"A8",X"70",X"C9",X"ED",X"5B",
		X"A9",X"70",X"16",X"00",X"21",X"EF",X"1C",X"19",X"06",X"05",X"3A",X"15",X"74",X"0E",X"00",X"BE",
		X"CA",X"F7",X"28",X"0C",X"23",X"10",X"F8",X"21",X"03",X"1D",X"19",X"06",X"05",X"3A",X"14",X"74",
		X"BE",X"CA",X"0C",X"29",X"23",X"0C",X"0C",X"0C",X"0C",X"0C",X"10",X"F4",X"79",X"32",X"A1",X"70",
		X"21",X"F6",X"72",X"3A",X"AA",X"70",X"C6",X"01",X"47",X"11",X"14",X"00",X"19",X"10",X"FD",X"ED",
		X"5B",X"A1",X"70",X"16",X"00",X"19",X"7E",X"32",X"A2",X"70",X"C9",X"CD",X"DE",X"28",X"3A",X"A9",
		X"70",X"FE",X"00",X"20",X"06",X"21",X"5C",X"1D",X"C3",X"52",X"29",X"FE",X"05",X"20",X"06",X"21",
		X"58",X"1D",X"C3",X"52",X"29",X"FE",X"0A",X"20",X"06",X"21",X"60",X"1D",X"C3",X"52",X"29",X"21",
		X"64",X"1D",X"3A",X"A2",X"70",X"06",X"04",X"BE",X"CA",X"63",X"29",X"23",X"10",X"F9",X"AF",X"32",
		X"A3",X"70",X"C9",X"3E",X"01",X"32",X"A8",X"70",X"32",X"A3",X"70",X"C9",X"3A",X"14",X"74",X"21",
		X"8A",X"1C",X"06",X"05",X"BE",X"28",X"04",X"23",X"10",X"FA",X"C9",X"3E",X"01",X"32",X"A8",X"70",
		X"AF",X"32",X"A4",X"70",X"32",X"A5",X"70",X"32",X"A6",X"70",X"32",X"A7",X"70",X"3A",X"A2",X"70",
		X"FE",X"00",X"C8",X"FE",X"C6",X"C2",X"A1",X"29",X"3E",X"01",X"32",X"A5",X"70",X"32",X"A6",X"70",
		X"C9",X"FE",X"CE",X"C2",X"AF",X"29",X"3E",X"01",X"32",X"A4",X"70",X"32",X"A6",X"70",X"C9",X"FE",
		X"DA",X"C2",X"BA",X"29",X"3E",X"01",X"32",X"A6",X"70",X"C9",X"FE",X"DE",X"C2",X"C5",X"29",X"3E",
		X"01",X"32",X"A5",X"70",X"C9",X"FE",X"E2",X"C2",X"D0",X"29",X"3E",X"01",X"32",X"A4",X"70",X"C9",
		X"FE",X"F9",X"C0",X"3E",X"01",X"32",X"A4",X"70",X"32",X"A5",X"70",X"C9",X"3A",X"14",X"74",X"21",
		X"8A",X"1C",X"06",X"05",X"BE",X"28",X"04",X"23",X"10",X"FA",X"C9",X"3E",X"01",X"32",X"A8",X"70",
		X"AF",X"32",X"A4",X"70",X"32",X"A5",X"70",X"32",X"A6",X"70",X"32",X"A7",X"70",X"3A",X"A2",X"70",
		X"FE",X"00",X"C8",X"FE",X"CA",X"C2",X"11",X"2A",X"3E",X"01",X"32",X"A5",X"70",X"32",X"A7",X"70",
		X"C9",X"FE",X"D2",X"C2",X"1F",X"2A",X"3E",X"01",X"32",X"A4",X"70",X"32",X"A7",X"70",X"C9",X"FE",
		X"D6",X"C2",X"2A",X"2A",X"3E",X"01",X"32",X"A7",X"70",X"C9",X"FE",X"DE",X"C2",X"35",X"2A",X"3E",
		X"01",X"32",X"A5",X"70",X"C9",X"FE",X"E2",X"C2",X"40",X"2A",X"3E",X"01",X"32",X"A4",X"70",X"C9",
		X"FE",X"F9",X"C0",X"3E",X"01",X"32",X"A4",X"70",X"32",X"A5",X"70",X"C9",X"3A",X"15",X"74",X"21",
		X"93",X"1C",X"06",X"05",X"BE",X"28",X"04",X"23",X"10",X"FA",X"C9",X"3E",X"01",X"32",X"A8",X"70",
		X"AF",X"32",X"A4",X"70",X"32",X"A5",X"70",X"32",X"A6",X"70",X"32",X"A7",X"70",X"3A",X"A2",X"70",
		X"FE",X"00",X"C8",X"FE",X"C6",X"C2",X"81",X"2A",X"3E",X"01",X"32",X"A6",X"70",X"32",X"A5",X"70",
		X"C9",X"FE",X"CA",X"C2",X"8F",X"2A",X"3E",X"01",X"32",X"A7",X"70",X"32",X"A5",X"70",X"C9",X"FE",
		X"D6",X"C2",X"9A",X"2A",X"3E",X"01",X"32",X"A7",X"70",X"C9",X"FE",X"DA",X"C2",X"A5",X"2A",X"3E",
		X"01",X"32",X"A6",X"70",X"C9",X"FE",X"DE",X"C2",X"B0",X"2A",X"3E",X"01",X"32",X"A5",X"70",X"C9",
		X"FE",X"B2",X"C0",X"3E",X"01",X"32",X"A6",X"70",X"32",X"A7",X"70",X"C9",X"3A",X"15",X"74",X"21",
		X"93",X"1C",X"06",X"05",X"BE",X"28",X"04",X"23",X"10",X"FA",X"C9",X"3E",X"01",X"32",X"A8",X"70",
		X"AF",X"32",X"A4",X"70",X"32",X"A5",X"70",X"32",X"A6",X"70",X"32",X"A7",X"70",X"3A",X"A2",X"70",
		X"FE",X"00",X"C8",X"FE",X"CE",X"C2",X"F1",X"2A",X"3E",X"01",X"32",X"A6",X"70",X"32",X"A4",X"70",
		X"C9",X"FE",X"D2",X"C2",X"FF",X"2A",X"3E",X"01",X"32",X"A7",X"70",X"32",X"A4",X"70",X"C9",X"FE",
		X"D6",X"C2",X"0A",X"2B",X"3E",X"01",X"32",X"A7",X"70",X"C9",X"FE",X"DA",X"C2",X"15",X"2B",X"3E",
		X"01",X"32",X"A6",X"70",X"C9",X"FE",X"E2",X"C2",X"20",X"2B",X"3E",X"01",X"32",X"A4",X"70",X"C9",
		X"FE",X"B2",X"C0",X"3E",X"01",X"32",X"A6",X"70",X"32",X"A7",X"70",X"C9",X"3A",X"59",X"70",X"3D",
		X"32",X"59",X"70",X"C0",X"3A",X"0A",X"71",X"32",X"59",X"70",X"3A",X"CC",X"70",X"FE",X"01",X"CA",
		X"2D",X"2F",X"CD",X"48",X"2B",X"C3",X"9C",X"2B",X"3A",X"54",X"70",X"FE",X"01",X"CA",X"65",X"2B",
		X"3A",X"39",X"70",X"FE",X"01",X"CA",X"61",X"2B",X"FE",X"02",X"CA",X"61",X"2B",X"CD",X"6C",X"2B",
		X"C9",X"CD",X"84",X"2B",X"C9",X"CD",X"84",X"2B",X"CD",X"6C",X"2B",X"C9",X"3A",X"32",X"70",X"2F",
		X"CB",X"5F",X"CA",X"7B",X"2B",X"3E",X"03",X"32",X"57",X"70",X"C9",X"CB",X"67",X"C8",X"3E",X"04",
		X"32",X"57",X"70",X"C9",X"3A",X"32",X"70",X"2F",X"CB",X"6F",X"CA",X"93",X"2B",X"3E",X"01",X"32",
		X"57",X"70",X"C9",X"CB",X"77",X"C8",X"3E",X"02",X"32",X"57",X"70",X"C9",X"3A",X"53",X"70",X"FE",
		X"00",X"C0",X"3A",X"57",X"70",X"FE",X"03",X"CA",X"B7",X"2B",X"FE",X"04",X"CA",X"14",X"2C",X"FE",
		X"02",X"CA",X"CD",X"2C",X"C3",X"72",X"2C",X"00",X"3A",X"50",X"70",X"FE",X"00",X"C2",X"10",X"2C",
		X"3E",X"01",X"32",X"51",X"70",X"32",X"52",X"70",X"CD",X"9C",X"2E",X"CD",X"11",X"2E",X"3A",X"01",
		X"70",X"C6",X"04",X"E6",X"FE",X"4F",X"3A",X"22",X"74",X"E6",X"01",X"B1",X"F6",X"80",X"32",X"22",
		X"74",X"3A",X"00",X"70",X"FE",X"04",X"CC",X"28",X"2D",X"21",X"24",X"74",X"35",X"7E",X"C6",X"10",
		X"32",X"28",X"74",X"3A",X"01",X"70",X"C6",X"06",X"E6",X"FE",X"4F",X"3A",X"26",X"74",X"E6",X"01",
		X"B1",X"F6",X"80",X"32",X"26",X"74",X"3E",X"01",X"32",X"00",X"70",X"3E",X"03",X"32",X"39",X"70",
		X"CD",X"37",X"2D",X"C9",X"00",X"3A",X"4F",X"70",X"FE",X"00",X"C2",X"6E",X"2C",X"3E",X"01",X"32",
		X"51",X"70",X"32",X"52",X"70",X"CD",X"9C",X"2E",X"CD",X"D2",X"2D",X"3A",X"01",X"70",X"C6",X"04",
		X"E6",X"FE",X"4F",X"3A",X"22",X"74",X"E6",X"01",X"B1",X"E6",X"3F",X"32",X"22",X"74",X"3A",X"00",
		X"70",X"FE",X"04",X"CC",X"28",X"2D",X"21",X"24",X"74",X"34",X"7E",X"D6",X"10",X"21",X"28",X"74",
		X"77",X"3A",X"01",X"70",X"C6",X"06",X"E6",X"FE",X"4F",X"3A",X"26",X"74",X"E6",X"01",X"B1",X"E6",
		X"3F",X"32",X"26",X"74",X"3E",X"01",X"32",X"00",X"70",X"3E",X"04",X"32",X"39",X"70",X"CD",X"37",
		X"2D",X"C9",X"00",X"3A",X"51",X"70",X"FE",X"00",X"C2",X"C9",X"2C",X"3E",X"01",X"32",X"50",X"70",
		X"32",X"4F",X"70",X"CD",X"50",X"2E",X"CD",X"54",X"2D",X"3A",X"01",X"70",X"E6",X"FE",X"4F",X"3A",
		X"22",X"74",X"E6",X"01",X"B1",X"E6",X"3F",X"32",X"22",X"74",X"3A",X"00",X"70",X"FE",X"01",X"CC",
		X"28",X"2D",X"21",X"25",X"74",X"35",X"7E",X"C6",X"10",X"32",X"29",X"74",X"3A",X"01",X"70",X"C6",
		X"02",X"E6",X"FE",X"4F",X"3A",X"26",X"74",X"E6",X"01",X"B1",X"E6",X"3F",X"32",X"26",X"74",X"3E",
		X"04",X"32",X"00",X"70",X"3E",X"01",X"32",X"39",X"70",X"CD",X"37",X"2D",X"C9",X"00",X"3A",X"52",
		X"70",X"FE",X"00",X"C2",X"24",X"2D",X"3E",X"01",X"32",X"50",X"70",X"32",X"4F",X"70",X"CD",X"50",
		X"2E",X"CD",X"93",X"2D",X"3A",X"01",X"70",X"E6",X"FE",X"4F",X"3A",X"22",X"74",X"E6",X"01",X"B1",
		X"F6",X"C0",X"32",X"22",X"74",X"3A",X"00",X"70",X"FE",X"01",X"CC",X"28",X"2D",X"21",X"25",X"74",
		X"34",X"7E",X"D6",X"0F",X"32",X"29",X"74",X"3A",X"01",X"70",X"C6",X"02",X"E6",X"FE",X"4F",X"3A",
		X"26",X"74",X"E6",X"01",X"B1",X"F6",X"C0",X"32",X"26",X"74",X"3E",X"04",X"32",X"00",X"70",X"3E",
		X"02",X"32",X"39",X"70",X"CD",X"37",X"2D",X"C9",X"F5",X"3A",X"24",X"74",X"32",X"28",X"74",X"3A",
		X"25",X"74",X"32",X"29",X"74",X"F1",X"C9",X"3A",X"45",X"70",X"3D",X"20",X"13",X"3A",X"22",X"74",
		X"EE",X"01",X"32",X"22",X"74",X"3A",X"26",X"74",X"EE",X"01",X"32",X"26",X"74",X"3A",X"58",X"70",
		X"32",X"45",X"70",X"C9",X"3A",X"24",X"74",X"4F",X"21",X"E2",X"2E",X"06",X"04",X"16",X"00",X"7E",
		X"23",X"B9",X"28",X"07",X"3E",X"05",X"82",X"57",X"10",X"F5",X"C9",X"7A",X"32",X"43",X"70",X"21",
		X"E6",X"2E",X"3A",X"25",X"74",X"4F",X"06",X"05",X"16",X"00",X"7E",X"23",X"B9",X"28",X"09",X"14",
		X"10",X"F8",X"3E",X"00",X"32",X"42",X"70",X"C9",X"3A",X"43",X"70",X"82",X"32",X"3A",X"70",X"3E",
		X"01",X"18",X"F1",X"3A",X"24",X"74",X"4F",X"21",X"E2",X"2E",X"06",X"04",X"16",X"00",X"7E",X"23",
		X"B9",X"28",X"07",X"3E",X"05",X"82",X"57",X"10",X"F5",X"C9",X"7A",X"32",X"43",X"70",X"21",X"EB",
		X"2E",X"3A",X"25",X"74",X"4F",X"06",X"05",X"16",X"00",X"7E",X"23",X"B9",X"28",X"09",X"14",X"10",
		X"F8",X"3E",X"00",X"32",X"42",X"70",X"C9",X"3A",X"43",X"70",X"82",X"32",X"3A",X"70",X"3E",X"01",
		X"18",X"F1",X"3A",X"25",X"74",X"4F",X"21",X"F0",X"2E",X"06",X"05",X"16",X"00",X"7E",X"23",X"B9",
		X"28",X"04",X"14",X"10",X"F8",X"C9",X"7A",X"32",X"43",X"70",X"21",X"F9",X"2E",X"3A",X"24",X"74",
		X"4F",X"06",X"04",X"16",X"00",X"7E",X"23",X"B9",X"28",X"0C",X"3E",X"05",X"82",X"57",X"10",X"F5",
		X"3E",X"00",X"32",X"42",X"70",X"C9",X"3A",X"43",X"70",X"82",X"32",X"3A",X"70",X"3E",X"01",X"18",
		X"F1",X"3A",X"25",X"74",X"4F",X"21",X"F0",X"2E",X"06",X"05",X"16",X"00",X"7E",X"23",X"B9",X"28",
		X"04",X"14",X"10",X"F8",X"C9",X"7A",X"32",X"43",X"70",X"21",X"F5",X"2E",X"3A",X"24",X"74",X"4F",
		X"06",X"04",X"16",X"00",X"7E",X"23",X"B9",X"28",X"0C",X"3E",X"05",X"82",X"57",X"10",X"F5",X"3E",
		X"00",X"32",X"42",X"70",X"C9",X"3A",X"43",X"70",X"82",X"32",X"3A",X"70",X"3E",X"01",X"18",X"F1",
		X"21",X"25",X"74",X"7E",X"FE",X"10",X"CA",X"98",X"2E",X"FE",X"F0",X"CA",X"9A",X"2E",X"3A",X"24",
		X"74",X"FE",X"29",X"38",X"1C",X"FE",X"37",X"38",X"1A",X"FE",X"59",X"38",X"14",X"FE",X"67",X"38",
		X"16",X"FE",X"89",X"38",X"0C",X"FE",X"97",X"38",X"12",X"FE",X"B9",X"38",X"04",X"FE",X"C7",X"38",
		X"0E",X"00",X"C9",X"3E",X"30",X"18",X"0A",X"3E",X"60",X"18",X"06",X"3E",X"90",X"18",X"02",X"3E",
		X"C0",X"32",X"24",X"74",X"32",X"28",X"74",X"C9",X"34",X"C9",X"35",X"C9",X"3A",X"25",X"74",X"FE",
		X"11",X"38",X"24",X"FE",X"1F",X"38",X"22",X"FE",X"41",X"38",X"1C",X"FE",X"4F",X"38",X"1E",X"FE",
		X"71",X"38",X"14",X"FE",X"7F",X"38",X"1A",X"FE",X"A1",X"38",X"0C",X"FE",X"AF",X"38",X"16",X"FE",
		X"D1",X"38",X"04",X"FE",X"DF",X"38",X"12",X"00",X"C9",X"3E",X"18",X"18",X"0E",X"3E",X"48",X"18",
		X"0A",X"3E",X"78",X"18",X"06",X"3E",X"A8",X"18",X"02",X"3E",X"D8",X"32",X"25",X"74",X"32",X"29",
		X"74",X"C9",X"C0",X"90",X"60",X"30",X"26",X"56",X"86",X"B6",X"E6",X"00",X"3A",X"6A",X"9A",X"CA",
		X"18",X"48",X"78",X"A8",X"D8",X"CE",X"9E",X"6E",X"3E",X"B2",X"82",X"52",X"22",X"CD",X"CF",X"07",
		X"21",X"81",X"2F",X"22",X"CD",X"70",X"AF",X"32",X"5D",X"70",X"3E",X"01",X"32",X"70",X"70",X"32",
		X"CC",X"70",X"3E",X"0C",X"32",X"67",X"73",X"32",X"0A",X"71",X"CD",X"E0",X"40",X"CD",X"2D",X"3F",
		X"06",X"3C",X"21",X"0A",X"73",X"36",X"00",X"23",X"10",X"FB",X"C3",X"81",X"30",X"3A",X"04",X"70",
		X"FE",X"00",X"20",X"2F",X"3A",X"CF",X"70",X"FE",X"00",X"CA",X"43",X"2F",X"3D",X"32",X"CF",X"70",
		X"C3",X"9C",X"2B",X"3A",X"54",X"70",X"FE",X"00",X"CA",X"9C",X"2B",X"3E",X"08",X"32",X"CF",X"70",
		X"2A",X"CD",X"70",X"7E",X"FE",X"FF",X"CA",X"63",X"2F",X"32",X"57",X"70",X"23",X"22",X"CD",X"70",
		X"C3",X"9C",X"2B",X"DD",X"E1",X"AF",X"32",X"0D",X"74",X"32",X"11",X"74",X"32",X"15",X"74",X"32",
		X"19",X"74",X"32",X"1D",X"74",X"32",X"21",X"74",X"32",X"25",X"74",X"32",X"29",X"74",X"C3",X"19",
		X"10",X"01",X"01",X"01",X"04",X"02",X"04",X"02",X"03",X"04",X"04",X"02",X"02",X"03",X"04",X"01",
		X"04",X"02",X"04",X"04",X"01",X"04",X"02",X"04",X"04",X"04",X"01",X"03",X"03",X"04",X"04",X"01",
		X"01",X"01",X"03",X"03",X"03",X"02",X"03",X"01",X"03",X"03",X"02",X"03",X"01",X"03",X"02",X"03",
		X"02",X"04",X"02",X"02",X"01",X"01",X"02",X"04",X"02",X"04",X"01",X"01",X"02",X"01",X"04",X"03",
		X"03",X"04",X"04",X"03",X"02",X"02",X"01",X"01",X"02",X"02",X"03",X"04",X"01",X"01",X"03",X"04",
		X"04",X"03",X"02",X"01",X"02",X"01",X"02",X"01",X"01",X"FF",X"21",X"42",X"88",X"22",X"00",X"71",
		X"22",X"04",X"71",X"21",X"5F",X"88",X"22",X"02",X"71",X"21",X"A2",X"8B",X"22",X"06",X"71",X"06",
		X"10",X"C5",X"CD",X"05",X"30",X"CD",X"1D",X"30",X"CD",X"3B",X"30",X"CD",X"59",X"30",X"CD",X"77",
		X"30",X"C1",X"10",X"ED",X"C9",X"11",X"00",X"10",X"06",X"1E",X"2A",X"04",X"71",X"36",X"10",X"E5",
		X"19",X"36",X"00",X"E1",X"23",X"10",X"F6",X"23",X"23",X"22",X"04",X"71",X"C9",X"2A",X"06",X"71",
		X"E5",X"06",X"1E",X"11",X"00",X"10",X"36",X"10",X"E5",X"19",X"36",X"00",X"E1",X"23",X"10",X"F6",
		X"E1",X"01",X"20",X"00",X"97",X"ED",X"42",X"22",X"06",X"71",X"C9",X"06",X"1C",X"11",X"00",X"10",
		X"2A",X"00",X"71",X"E5",X"36",X"10",X"E5",X"19",X"36",X"00",X"E1",X"C5",X"01",X"20",X"00",X"09",
		X"C1",X"10",X"F1",X"E1",X"23",X"22",X"00",X"71",X"C9",X"2A",X"02",X"71",X"E5",X"06",X"1C",X"11",
		X"00",X"10",X"36",X"10",X"E5",X"19",X"36",X"00",X"E1",X"C5",X"01",X"20",X"00",X"09",X"C1",X"10",
		X"F1",X"E1",X"2B",X"22",X"02",X"71",X"C9",X"01",X"80",X"05",X"0B",X"78",X"B1",X"C2",X"7A",X"30",
		X"C9",X"00",X"3E",X"08",X"32",X"58",X"70",X"32",X"45",X"70",X"32",X"53",X"73",X"32",X"52",X"73",
		X"32",X"57",X"73",X"32",X"56",X"73",X"32",X"5D",X"73",X"32",X"5C",X"73",X"3E",X"05",X"32",X"B5",
		X"70",X"32",X"B6",X"70",X"3E",X"10",X"32",X"01",X"70",X"CD",X"73",X"0D",X"22",X"62",X"73",X"3E",
		X"04",X"32",X"0B",X"74",X"3E",X"08",X"32",X"0F",X"74",X"32",X"13",X"74",X"AF",X"32",X"17",X"74",
		X"32",X"AC",X"70",X"32",X"AD",X"70",X"32",X"6F",X"70",X"21",X"74",X"70",X"06",X"0F",X"36",X"00",
		X"23",X"10",X"FB",X"AF",X"32",X"BE",X"70",X"32",X"BF",X"70",X"06",X"07",X"21",X"C5",X"70",X"36",
		X"00",X"23",X"10",X"FB",X"3A",X"CC",X"70",X"FE",X"00",X"20",X"08",X"3E",X"09",X"32",X"67",X"73",
		X"32",X"0A",X"71",X"3E",X"10",X"32",X"68",X"73",X"32",X"5B",X"70",X"3E",X"14",X"32",X"73",X"70",
		X"3E",X"30",X"32",X"68",X"70",X"3E",X"07",X"32",X"EA",X"70",X"21",X"44",X"18",X"22",X"BA",X"70",
		X"3E",X"02",X"32",X"88",X"70",X"3E",X"7D",X"32",X"1C",X"74",X"3E",X"0A",X"32",X"1D",X"74",X"3E",
		X"58",X"32",X"1A",X"74",X"3E",X"08",X"32",X"1B",X"74",X"3E",X"FF",X"32",X"64",X"73",X"3E",X"90",
		X"32",X"BC",X"70",X"32",X"BD",X"70",X"3E",X"30",X"32",X"68",X"70",X"06",X"06",X"21",X"0A",X"70",
		X"11",X"C5",X"70",X"7E",X"12",X"13",X"23",X"10",X"FA",X"3E",X"18",X"32",X"0D",X"74",X"32",X"0C",
		X"74",X"32",X"11",X"74",X"32",X"10",X"74",X"3E",X"01",X"32",X"94",X"70",X"32",X"AA",X"70",X"3E",
		X"02",X"32",X"9F",X"70",X"3E",X"48",X"32",X"15",X"74",X"3E",X"C0",X"32",X"14",X"74",X"3E",X"2C",
		X"32",X"B9",X"70",X"32",X"16",X"74",X"AF",X"32",X"AE",X"70",X"32",X"C2",X"70",X"32",X"C3",X"70",
		X"32",X"69",X"73",X"32",X"07",X"75",X"32",X"49",X"70",X"21",X"00",X"10",X"22",X"69",X"70",X"22",
		X"6B",X"70",X"22",X"6D",X"70",X"22",X"B7",X"70",X"22",X"84",X"70",X"3E",X"01",X"32",X"50",X"70",
		X"32",X"4F",X"70",X"21",X"0A",X"73",X"11",X"6E",X"73",X"01",X"63",X"00",X"ED",X"B0",X"AF",X"32",
		X"F7",X"70",X"32",X"F8",X"70",X"3A",X"CC",X"70",X"FE",X"00",X"28",X"09",X"21",X"39",X"0E",X"22",
		X"62",X"73",X"C3",X"5B",X"35",X"CD",X"73",X"0D",X"22",X"62",X"73",X"C3",X"5B",X"35",X"00",X"00",
		X"AF",X"32",X"56",X"70",X"CD",X"3D",X"35",X"CD",X"F2",X"31",X"CD",X"25",X"16",X"CD",X"F1",X"54",
		X"CD",X"F2",X"38",X"CD",X"A4",X"14",X"CD",X"7F",X"3C",X"CD",X"B6",X"17",X"CD",X"0E",X"32",X"C3",
		X"CF",X"31",X"C3",X"38",X"34",X"CD",X"C6",X"16",X"C3",X"98",X"34",X"CD",X"0E",X"25",X"C3",X"CF",
		X"34",X"CD",X"A8",X"1F",X"C3",X"06",X"35",X"CD",X"65",X"19",X"CD",X"2C",X"2B",X"C9",X"3A",X"6F",
		X"70",X"FE",X"01",X"CA",X"36",X"32",X"3A",X"F7",X"70",X"FE",X"01",X"C8",X"3A",X"35",X"70",X"47",
		X"3A",X"78",X"70",X"B8",X"C0",X"3A",X"70",X"70",X"3C",X"32",X"70",X"70",X"47",X"CD",X"EB",X"36",
		X"3E",X"01",X"32",X"F7",X"70",X"C9",X"3A",X"F8",X"70",X"FE",X"01",X"C8",X"3A",X"35",X"70",X"47",
		X"3A",X"7F",X"70",X"B8",X"C0",X"3A",X"71",X"70",X"3C",X"32",X"71",X"70",X"47",X"CD",X"EB",X"36",
		X"3E",X"01",X"32",X"F8",X"70",X"C9",X"00",X"21",X"67",X"73",X"34",X"34",X"34",X"34",X"3E",X"01",
		X"32",X"56",X"70",X"CD",X"3D",X"35",X"CD",X"F2",X"31",X"CD",X"2C",X"2B",X"CD",X"25",X"16",X"CD",
		X"F1",X"54",X"CD",X"F2",X"38",X"CD",X"A4",X"14",X"CD",X"B6",X"17",X"CD",X"E4",X"44",X"CD",X"0E",
		X"32",X"CD",X"F9",X"32",X"3A",X"24",X"74",X"FE",X"A8",X"C2",X"5E",X"32",X"3A",X"25",X"74",X"FE",
		X"D8",X"C2",X"5E",X"32",X"21",X"67",X"73",X"35",X"35",X"35",X"35",X"3E",X"11",X"32",X"22",X"74",
		X"3E",X"13",X"32",X"26",X"74",X"3E",X"A8",X"32",X"24",X"74",X"32",X"28",X"74",X"3E",X"D0",X"32",
		X"25",X"74",X"3E",X"E0",X"32",X"29",X"74",X"3E",X"01",X"32",X"C0",X"70",X"CD",X"B6",X"17",X"AF",
		X"32",X"0D",X"74",X"32",X"11",X"74",X"32",X"15",X"74",X"32",X"19",X"74",X"32",X"1D",X"74",X"32",
		X"21",X"74",X"CD",X"AD",X"33",X"CD",X"8C",X"33",X"CD",X"77",X"08",X"3E",X"05",X"32",X"11",X"75",
		X"21",X"00",X"E8",X"22",X"E8",X"70",X"CD",X"0E",X"09",X"2A",X"E8",X"70",X"2B",X"22",X"E8",X"70",
		X"7C",X"B5",X"C2",X"E6",X"32",X"CD",X"F9",X"33",X"C9",X"DD",X"21",X"39",X"89",X"DD",X"36",X"E0",
		X"F0",X"DD",X"36",X"E1",X"F1",X"DD",X"36",X"FF",X"EF",X"DD",X"36",X"FE",X"EE",X"DD",X"36",X"00",
		X"EA",X"DD",X"36",X"01",X"EB",X"DD",X"36",X"1F",X"F3",X"DD",X"36",X"1E",X"F2",X"DD",X"36",X"20",
		X"EC",X"DD",X"36",X"21",X"ED",X"DD",X"36",X"40",X"F4",X"DD",X"36",X"41",X"F5",X"DD",X"21",X"39",
		X"99",X"DD",X"E5",X"06",X"02",X"DD",X"36",X"00",X"14",X"DD",X"36",X"20",X"14",X"DD",X"23",X"10",
		X"F4",X"DD",X"E1",X"DD",X"36",X"E0",X"13",X"DD",X"36",X"E1",X"13",X"DD",X"36",X"FF",X"13",X"DD",
		X"36",X"FE",X"13",X"DD",X"36",X"1F",X"13",X"DD",X"36",X"1E",X"13",X"DD",X"36",X"40",X"13",X"DD",
		X"36",X"41",X"13",X"DD",X"21",X"3B",X"89",X"DD",X"36",X"00",X"DE",X"DD",X"36",X"01",X"DF",X"DD",
		X"36",X"20",X"E0",X"DD",X"36",X"21",X"E1",X"DD",X"21",X"3B",X"99",X"DD",X"36",X"00",X"11",X"DD",
		X"36",X"01",X"11",X"DD",X"36",X"20",X"11",X"DD",X"36",X"21",X"11",X"C9",X"DD",X"21",X"39",X"89",
		X"DD",X"36",X"01",X"10",X"DD",X"36",X"21",X"10",X"DD",X"36",X"00",X"0E",X"DD",X"36",X"20",X"0F",
		X"DD",X"21",X"39",X"99",X"DD",X"36",X"00",X"34",X"DD",X"36",X"20",X"34",X"C9",X"3E",X"1C",X"32",
		X"0A",X"74",X"3E",X"28",X"32",X"0B",X"74",X"3A",X"49",X"70",X"32",X"94",X"70",X"3E",X"A8",X"32",
		X"0C",X"74",X"3E",X"B8",X"32",X"0D",X"74",X"3E",X"08",X"32",X"11",X"75",X"01",X"00",X"A0",X"CD",
		X"16",X"3C",X"3E",X"1D",X"32",X"0A",X"74",X"3E",X"09",X"32",X"11",X"75",X"01",X"00",X"A0",X"CD",
		X"16",X"3C",X"3E",X"1E",X"32",X"0A",X"74",X"3E",X"0A",X"32",X"11",X"75",X"01",X"FF",X"FF",X"CD",
		X"16",X"3C",X"CD",X"16",X"3C",X"CD",X"16",X"3C",X"C9",X"3E",X"10",X"32",X"01",X"70",X"3E",X"04",
		X"32",X"0B",X"74",X"3E",X"08",X"32",X"0F",X"74",X"32",X"13",X"74",X"AF",X"32",X"17",X"74",X"32",
		X"22",X"74",X"32",X"26",X"74",X"32",X"1D",X"74",X"3E",X"58",X"32",X"1A",X"74",X"3E",X"08",X"32",
		X"1B",X"74",X"3E",X"2C",X"32",X"B9",X"70",X"32",X"16",X"74",X"3E",X"28",X"32",X"23",X"74",X"32",
		X"27",X"74",X"3E",X"02",X"32",X"88",X"70",X"C9",X"3A",X"63",X"70",X"FE",X"00",X"CA",X"F5",X"31",
		X"2A",X"B7",X"70",X"2B",X"22",X"B7",X"70",X"7C",X"B5",X"C2",X"F8",X"31",X"AF",X"32",X"63",X"70",
		X"21",X"00",X"10",X"22",X"B7",X"70",X"21",X"88",X"70",X"3E",X"01",X"32",X"C0",X"70",X"AF",X"32",
		X"B1",X"70",X"32",X"B4",X"70",X"32",X"B3",X"70",X"21",X"44",X"18",X"22",X"BA",X"70",X"3E",X"25",
		X"32",X"61",X"73",X"32",X"B2",X"70",X"3E",X"02",X"32",X"88",X"70",X"3E",X"7D",X"32",X"1C",X"74",
		X"3E",X"0A",X"32",X"1D",X"74",X"3E",X"58",X"32",X"1A",X"74",X"3E",X"08",X"32",X"1B",X"74",X"3A",
		X"64",X"73",X"32",X"C4",X"70",X"C3",X"F8",X"31",X"3A",X"61",X"70",X"FE",X"00",X"CA",X"FB",X"31",
		X"2A",X"6D",X"70",X"2B",X"22",X"6D",X"70",X"7C",X"B5",X"C2",X"FE",X"31",X"AF",X"32",X"61",X"70",
		X"21",X"00",X"10",X"22",X"6D",X"70",X"21",X"AA",X"70",X"3E",X"60",X"32",X"14",X"74",X"3A",X"49",
		X"70",X"FE",X"02",X"28",X"05",X"3C",X"77",X"C3",X"FE",X"31",X"3D",X"77",X"C3",X"FE",X"31",X"3A",
		X"60",X"70",X"FE",X"00",X"CA",X"01",X"32",X"2A",X"6B",X"70",X"2B",X"22",X"6B",X"70",X"7C",X"B5",
		X"C2",X"04",X"32",X"AF",X"32",X"60",X"70",X"21",X"00",X"10",X"22",X"6B",X"70",X"21",X"9F",X"70",
		X"3E",X"60",X"32",X"10",X"74",X"3A",X"49",X"70",X"FE",X"02",X"28",X"05",X"3C",X"77",X"C3",X"04",
		X"32",X"3D",X"77",X"C3",X"04",X"32",X"3A",X"5F",X"70",X"FE",X"00",X"CA",X"07",X"32",X"2A",X"69",
		X"70",X"2B",X"22",X"69",X"70",X"7C",X"B5",X"C2",X"0A",X"32",X"AF",X"32",X"5F",X"70",X"21",X"00",
		X"10",X"22",X"69",X"70",X"21",X"94",X"70",X"3E",X"60",X"32",X"0C",X"74",X"3A",X"49",X"70",X"FE",
		X"02",X"28",X"05",X"3C",X"77",X"C3",X"0A",X"32",X"3D",X"77",X"C3",X"0A",X"32",X"3A",X"64",X"70",
		X"FE",X"00",X"C8",X"2A",X"84",X"70",X"2B",X"22",X"84",X"70",X"7C",X"B5",X"C0",X"AF",X"32",X"64",
		X"70",X"32",X"21",X"74",X"21",X"00",X"10",X"22",X"84",X"70",X"C9",X"3A",X"CC",X"70",X"FE",X"01",
		X"28",X"3A",X"CD",X"DA",X"2F",X"3A",X"07",X"75",X"FE",X"00",X"28",X"05",X"3E",X"0D",X"32",X"11",
		X"75",X"11",X"18",X"42",X"21",X"B0",X"8A",X"0E",X"05",X"CD",X"71",X"41",X"DD",X"21",X"2F",X"89",
		X"06",X"0C",X"0E",X"38",X"CD",X"A2",X"3D",X"01",X"FF",X"FF",X"CD",X"16",X"3C",X"CD",X"16",X"3C",
		X"CD",X"16",X"3C",X"CD",X"16",X"3C",X"CD",X"16",X"3C",X"CD",X"DA",X"2F",X"CD",X"2E",X"38",X"CD",
		X"4A",X"37",X"21",X"70",X"70",X"35",X"46",X"3E",X"FF",X"B8",X"20",X"01",X"34",X"CD",X"EB",X"36",
		X"CD",X"06",X"19",X"3A",X"C2",X"70",X"CD",X"BF",X"35",X"CD",X"72",X"2C",X"C3",X"CE",X"31",X"3C",
		X"47",X"3A",X"CC",X"70",X"FE",X"01",X"C8",X"78",X"21",X"7F",X"88",X"11",X"20",X"00",X"36",X"FD",
		X"19",X"10",X"FB",X"47",X"21",X"7F",X"98",X"36",X"18",X"19",X"10",X"FB",X"C9",X"00",X"3E",X"01",
		X"32",X"07",X"75",X"3A",X"70",X"70",X"FE",X"00",X"CC",X"08",X"36",X"AF",X"32",X"1D",X"74",X"3A",
		X"71",X"70",X"FE",X"00",X"CA",X"FD",X"35",X"CD",X"30",X"37",X"C3",X"18",X"36",X"3A",X"70",X"70",
		X"FE",X"00",X"CA",X"AC",X"36",X"C3",X"5B",X"35",X"11",X"E5",X"41",X"CD",X"BF",X"36",X"21",X"79",
		X"70",X"22",X"F1",X"70",X"CD",X"8D",X"11",X"C9",X"CD",X"DA",X"2F",X"3E",X"0D",X"32",X"11",X"75",
		X"11",X"0B",X"42",X"21",X"B0",X"8A",X"0E",X"05",X"CD",X"71",X"41",X"DD",X"21",X"2F",X"89",X"06",
		X"0C",X"0E",X"38",X"CD",X"A2",X"3D",X"01",X"FF",X"FF",X"CD",X"16",X"3C",X"CD",X"16",X"3C",X"CD",
		X"16",X"3C",X"CD",X"16",X"3C",X"CD",X"16",X"3C",X"CD",X"DA",X"2F",X"CD",X"2E",X"38",X"CD",X"4A",
		X"37",X"21",X"71",X"70",X"35",X"46",X"3E",X"FF",X"B8",X"20",X"01",X"34",X"CD",X"EB",X"36",X"CD",
		X"06",X"19",X"3A",X"C3",X"70",X"CD",X"BF",X"35",X"CD",X"72",X"2C",X"C3",X"CE",X"31",X"00",X"3A",
		X"71",X"70",X"FE",X"00",X"CC",X"98",X"36",X"AF",X"32",X"1D",X"74",X"3A",X"70",X"70",X"FE",X"00",
		X"CA",X"8D",X"36",X"CD",X"30",X"37",X"AF",X"32",X"31",X"70",X"C3",X"5B",X"35",X"3A",X"71",X"70",
		X"FE",X"00",X"CA",X"AC",X"36",X"C3",X"18",X"36",X"11",X"EF",X"41",X"CD",X"BF",X"36",X"21",X"80",
		X"70",X"22",X"F1",X"70",X"CD",X"8D",X"11",X"AF",X"32",X"31",X"70",X"C9",X"3A",X"05",X"70",X"FE",
		X"00",X"C2",X"90",X"05",X"3A",X"04",X"70",X"FE",X"00",X"C2",X"90",X"05",X"C3",X"19",X"10",X"3E",
		X"03",X"32",X"11",X"75",X"21",X"90",X"8A",X"CD",X"71",X"41",X"11",X"31",X"42",X"21",X"8F",X"8A",
		X"CD",X"71",X"41",X"DD",X"21",X"6E",X"89",X"06",X"09",X"0E",X"39",X"CD",X"F1",X"3D",X"16",X"0C",
		X"01",X"FF",X"FF",X"CD",X"16",X"3C",X"15",X"C2",X"E0",X"36",X"C9",X"DD",X"21",X"5F",X"8B",X"FD",
		X"21",X"5F",X"9B",X"FD",X"36",X"E0",X"06",X"DD",X"36",X"E0",X"10",X"FD",X"36",X"00",X"06",X"DD",
		X"36",X"00",X"10",X"FD",X"36",X"20",X"06",X"DD",X"36",X"20",X"10",X"FD",X"36",X"40",X"06",X"DD",
		X"36",X"40",X"10",X"FD",X"36",X"40",X"06",X"DD",X"36",X"60",X"10",X"FD",X"36",X"60",X"06",X"97",
		X"B8",X"C8",X"97",X"21",X"BF",X"8B",X"11",X"20",X"00",X"36",X"0C",X"ED",X"52",X"10",X"FA",X"C9",
		X"06",X"63",X"21",X"0A",X"73",X"11",X"6E",X"73",X"4E",X"1A",X"77",X"79",X"12",X"23",X"13",X"10",
		X"F7",X"3A",X"6F",X"70",X"EE",X"01",X"32",X"6F",X"70",X"C9",X"CD",X"F7",X"37",X"CD",X"C4",X"3F",
		X"21",X"0A",X"73",X"0E",X"00",X"06",X"14",X"7E",X"FE",X"00",X"C2",X"65",X"37",X"C3",X"C1",X"37",
		X"23",X"0C",X"10",X"F3",X"C9",X"C5",X"E5",X"F5",X"DD",X"21",X"4B",X"5A",X"79",X"87",X"5F",X"16",
		X"00",X"DD",X"19",X"DD",X"66",X"00",X"DD",X"6E",X"01",X"E5",X"DD",X"E1",X"F1",X"DD",X"77",X"21",
		X"3C",X"DD",X"77",X"22",X"3C",X"DD",X"77",X"41",X"3C",X"DD",X"77",X"42",X"DD",X"36",X"00",X"00",
		X"DD",X"36",X"03",X"00",X"DD",X"36",X"60",X"00",X"DD",X"36",X"63",X"00",X"DD",X"36",X"01",X"F9",
		X"DD",X"36",X"02",X"FA",X"DD",X"36",X"20",X"B3",X"DD",X"36",X"40",X"B4",X"DD",X"36",X"61",X"F9",
		X"DD",X"36",X"62",X"FA",X"DD",X"36",X"23",X"B3",X"DD",X"36",X"43",X"B4",X"E1",X"C1",X"C3",X"60",
		X"37",X"C5",X"E5",X"DD",X"21",X"4B",X"5A",X"79",X"87",X"5F",X"16",X"00",X"DD",X"19",X"DD",X"66",
		X"00",X"DD",X"6E",X"01",X"E5",X"DD",X"E1",X"06",X"04",X"3E",X"A2",X"11",X"20",X"00",X"DD",X"77",
		X"00",X"3C",X"DD",X"77",X"01",X"3C",X"DD",X"77",X"02",X"3C",X"DD",X"77",X"03",X"3C",X"DD",X"19",
		X"10",X"EC",X"E1",X"C1",X"C3",X"60",X"37",X"DD",X"21",X"A2",X"98",X"06",X"04",X"00",X"3E",X"11",
		X"C5",X"CD",X"0D",X"38",X"11",X"40",X"00",X"DD",X"19",X"C1",X"10",X"F1",X"C9",X"06",X"04",X"C5",
		X"06",X"04",X"DD",X"77",X"00",X"DD",X"77",X"06",X"DD",X"77",X"0C",X"DD",X"77",X"12",X"DD",X"77",
		X"18",X"DD",X"23",X"10",X"ED",X"11",X"1C",X"00",X"DD",X"19",X"C1",X"10",X"E2",X"C9",X"3E",X"18",
		X"32",X"0D",X"74",X"32",X"0C",X"74",X"32",X"11",X"74",X"32",X"10",X"74",X"3E",X"01",X"32",X"94",
		X"70",X"32",X"AA",X"70",X"2A",X"50",X"73",X"22",X"46",X"73",X"AF",X"32",X"5E",X"70",X"32",X"0B",
		X"71",X"3E",X"02",X"32",X"9F",X"70",X"3E",X"48",X"32",X"15",X"74",X"3E",X"C0",X"32",X"14",X"74",
		X"3E",X"10",X"32",X"01",X"70",X"3E",X"C0",X"32",X"25",X"74",X"3E",X"30",X"32",X"24",X"74",X"32",
		X"28",X"74",X"3E",X"D0",X"32",X"29",X"74",X"3E",X"28",X"32",X"23",X"74",X"32",X"27",X"74",X"3E",
		X"04",X"32",X"0B",X"74",X"3E",X"08",X"32",X"0F",X"74",X"32",X"13",X"74",X"3E",X"FF",X"32",X"73",
		X"70",X"3E",X"01",X"32",X"50",X"70",X"32",X"4F",X"70",X"32",X"52",X"70",X"AF",X"32",X"51",X"70",
		X"32",X"49",X"70",X"32",X"53",X"70",X"32",X"54",X"70",X"32",X"39",X"70",X"32",X"57",X"70",X"32",
		X"46",X"70",X"32",X"B1",X"70",X"32",X"B4",X"70",X"32",X"B3",X"70",X"21",X"44",X"18",X"22",X"BA",
		X"70",X"3E",X"0A",X"32",X"1D",X"74",X"3E",X"7D",X"32",X"1C",X"74",X"21",X"44",X"18",X"22",X"BA",
		X"70",X"3E",X"30",X"32",X"68",X"70",X"21",X"A0",X"9B",X"11",X"20",X"00",X"06",X"09",X"97",X"36",
		X"07",X"ED",X"52",X"10",X"FA",X"21",X"40",X"99",X"06",X"09",X"97",X"36",X"07",X"ED",X"52",X"10",
		X"FA",X"C9",X"1E",X"00",X"3A",X"5E",X"70",X"FE",X"00",X"28",X"41",X"2A",X"46",X"73",X"2B",X"22",
		X"46",X"73",X"CD",X"A9",X"3A",X"7C",X"B5",X"20",X"33",X"AF",X"32",X"5E",X"70",X"2A",X"50",X"73",
		X"22",X"46",X"73",X"3E",X"30",X"32",X"68",X"70",X"3E",X"28",X"32",X"23",X"74",X"32",X"27",X"74",
		X"3E",X"04",X"32",X"0B",X"74",X"3E",X"08",X"32",X"0F",X"74",X"32",X"13",X"74",X"AF",X"32",X"55",
		X"70",X"3E",X"06",X"32",X"11",X"75",X"3A",X"B9",X"70",X"32",X"16",X"74",X"3A",X"94",X"70",X"21",
		X"49",X"70",X"BE",X"C2",X"69",X"3A",X"3A",X"5F",X"70",X"FE",X"00",X"C2",X"69",X"3A",X"21",X"0C",
		X"74",X"01",X"24",X"74",X"0A",X"C6",X"0A",X"BE",X"DA",X"70",X"39",X"D6",X"14",X"BE",X"D2",X"70",
		X"39",X"23",X"03",X"0A",X"C6",X"0A",X"BE",X"DA",X"70",X"39",X"D6",X"14",X"BE",X"DA",X"93",X"3A",
		X"1C",X"3A",X"9F",X"70",X"21",X"49",X"70",X"BE",X"C2",X"70",X"3A",X"3A",X"60",X"70",X"FE",X"00",
		X"C2",X"70",X"3A",X"21",X"10",X"74",X"01",X"24",X"74",X"0A",X"C6",X"0A",X"BE",X"DA",X"A4",X"39",
		X"D6",X"14",X"BE",X"30",X"0F",X"23",X"03",X"0A",X"C6",X"0A",X"BE",X"DA",X"A4",X"39",X"D6",X"14",
		X"BE",X"DA",X"93",X"3A",X"1C",X"3A",X"AA",X"70",X"21",X"49",X"70",X"BE",X"C2",X"77",X"3A",X"3A",
		X"61",X"70",X"FE",X"00",X"C2",X"77",X"3A",X"21",X"14",X"74",X"01",X"24",X"74",X"0A",X"C6",X"0A",
		X"BE",X"DA",X"D8",X"39",X"D6",X"14",X"BE",X"30",X"0F",X"23",X"03",X"0A",X"C6",X"0A",X"BE",X"DA",
		X"D8",X"39",X"D6",X"14",X"BE",X"DA",X"93",X"3A",X"1C",X"3A",X"87",X"70",X"21",X"49",X"70",X"BE",
		X"C2",X"7E",X"3A",X"21",X"18",X"74",X"01",X"24",X"74",X"0A",X"C6",X"0A",X"BE",X"38",X"15",X"D6",
		X"14",X"BE",X"D2",X"04",X"3A",X"23",X"03",X"0A",X"C6",X"0A",X"BE",X"DA",X"04",X"3A",X"D6",X"14",
		X"BE",X"DA",X"86",X"3B",X"1C",X"3A",X"88",X"70",X"21",X"49",X"70",X"BE",X"C2",X"85",X"3A",X"3A",
		X"63",X"70",X"FE",X"00",X"C2",X"85",X"3A",X"21",X"1C",X"74",X"01",X"24",X"74",X"0A",X"C6",X"0A",
		X"BE",X"38",X"12",X"D6",X"14",X"BE",X"30",X"0D",X"23",X"03",X"0A",X"C6",X"0A",X"BE",X"38",X"05",
		X"D6",X"14",X"BE",X"38",X"5E",X"1C",X"3A",X"89",X"70",X"21",X"49",X"70",X"BE",X"C2",X"8C",X"3A",
		X"3A",X"64",X"70",X"FE",X"00",X"C2",X"8C",X"3A",X"21",X"20",X"74",X"01",X"24",X"74",X"0A",X"C6",
		X"0D",X"BE",X"38",X"14",X"D6",X"1A",X"BE",X"30",X"0F",X"23",X"03",X"0A",X"C6",X"0D",X"BE",X"DA",
		X"68",X"3A",X"D6",X"1A",X"BE",X"DA",X"F9",X"3A",X"C9",X"06",X"07",X"10",X"FE",X"C3",X"70",X"39",
		X"06",X"07",X"10",X"FE",X"C3",X"A4",X"39",X"06",X"07",X"10",X"FE",X"C3",X"D8",X"39",X"06",X"07",
		X"10",X"FE",X"C3",X"04",X"3A",X"06",X"07",X"10",X"FE",X"C3",X"35",X"3A",X"06",X"07",X"10",X"FE",
		X"C3",X"68",X"3A",X"3A",X"5E",X"70",X"FE",X"00",X"CA",X"86",X"3B",X"FE",X"01",X"CA",X"A1",X"3A",
		X"C9",X"3E",X"0B",X"32",X"11",X"75",X"C3",X"0A",X"3B",X"3E",X"0A",X"BC",X"30",X"01",X"C9",X"3A",
		X"73",X"70",X"3D",X"32",X"73",X"70",X"C0",X"3E",X"FF",X"32",X"73",X"70",X"3A",X"23",X"74",X"FE",
		X"24",X"20",X"0D",X"E5",X"21",X"12",X"75",X"35",X"23",X"35",X"E1",X"3E",X"01",X"32",X"55",X"70",
		X"3A",X"23",X"74",X"EE",X"0C",X"32",X"23",X"74",X"3A",X"27",X"74",X"EE",X"0C",X"32",X"27",X"74",
		X"3A",X"0B",X"74",X"EE",X"04",X"32",X"0B",X"74",X"3A",X"0F",X"74",X"EE",X"0D",X"32",X"0F",X"74",
		X"3A",X"13",X"74",X"EE",X"0D",X"32",X"13",X"74",X"C9",X"3E",X"01",X"32",X"5E",X"70",X"3E",X"04",
		X"32",X"11",X"75",X"D5",X"E5",X"CD",X"28",X"1F",X"E1",X"D1",X"2B",X"2B",X"2B",X"3A",X"68",X"70",
		X"77",X"3C",X"32",X"68",X"70",X"16",X"00",X"21",X"5F",X"70",X"19",X"36",X"01",X"3E",X"24",X"32",
		X"23",X"74",X"32",X"27",X"74",X"AF",X"32",X"0B",X"74",X"3E",X"05",X"32",X"0F",X"74",X"32",X"13",
		X"74",X"3A",X"6F",X"70",X"FE",X"00",X"28",X"05",X"21",X"7E",X"70",X"18",X"03",X"21",X"77",X"70",
		X"3A",X"68",X"70",X"3D",X"FE",X"30",X"28",X"1D",X"FE",X"31",X"28",X"20",X"FE",X"32",X"28",X"23",
		X"FE",X"33",X"28",X"26",X"06",X"03",X"CD",X"F0",X"3E",X"2B",X"06",X"02",X"CD",X"F0",X"3E",X"3E",
		X"34",X"32",X"68",X"70",X"C9",X"06",X"02",X"2B",X"CD",X"F0",X"3E",X"C9",X"06",X"04",X"2B",X"CD",
		X"F0",X"3E",X"C9",X"06",X"08",X"2B",X"CD",X"F0",X"3E",X"C9",X"06",X"01",X"CD",X"F0",X"3E",X"2B",
		X"06",X"06",X"CD",X"F0",X"3E",X"C9",X"CD",X"1C",X"3C",X"3E",X"0C",X"32",X"11",X"75",X"3A",X"24",
		X"74",X"D6",X"10",X"32",X"28",X"74",X"3A",X"25",X"74",X"32",X"29",X"74",X"16",X"03",X"3E",X"08",
		X"32",X"22",X"74",X"3E",X"0A",X"32",X"26",X"74",X"3A",X"56",X"70",X"FE",X"00",X"CA",X"B3",X"3B",
		X"CD",X"3B",X"3C",X"CD",X"13",X"3C",X"CD",X"02",X"3C",X"15",X"20",X"F7",X"16",X"03",X"3E",X"09",
		X"32",X"22",X"74",X"3E",X"0B",X"32",X"26",X"74",X"3A",X"56",X"70",X"FE",X"00",X"CA",X"D3",X"3B",
		X"CD",X"57",X"3C",X"CD",X"13",X"3C",X"CD",X"02",X"3C",X"15",X"20",X"F7",X"3A",X"56",X"70",X"FE",
		X"00",X"CA",X"F2",X"3B",X"CD",X"5D",X"3C",X"DD",X"E1",X"DD",X"E1",X"21",X"67",X"73",X"35",X"35",
		X"35",X"35",X"01",X"FF",X"FF",X"CD",X"16",X"3C",X"CD",X"16",X"3C",X"AF",X"32",X"0D",X"74",X"C3",
		X"63",X"3C",X"3A",X"22",X"74",X"EE",X"40",X"32",X"22",X"74",X"3A",X"26",X"74",X"EE",X"40",X"32",
		X"26",X"74",X"C9",X"01",X"00",X"30",X"0B",X"78",X"B1",X"20",X"FB",X"C9",X"CD",X"13",X"3C",X"AF",
		X"32",X"0C",X"74",X"32",X"10",X"74",X"32",X"14",X"74",X"32",X"18",X"74",X"32",X"1C",X"74",X"32",
		X"20",X"74",X"3E",X"01",X"32",X"C0",X"70",X"CD",X"B6",X"17",X"C9",X"00",X"3E",X"1C",X"32",X"0A",
		X"74",X"3E",X"28",X"32",X"0B",X"74",X"3A",X"49",X"70",X"32",X"94",X"70",X"3E",X"A8",X"32",X"0C",
		X"74",X"3E",X"B8",X"32",X"0D",X"74",X"C9",X"3E",X"1D",X"32",X"0A",X"74",X"C9",X"3E",X"1F",X"32",
		X"0A",X"74",X"C9",X"AF",X"32",X"25",X"74",X"32",X"29",X"74",X"DD",X"E1",X"3A",X"CC",X"70",X"FE",
		X"01",X"CA",X"65",X"2F",X"3A",X"6F",X"70",X"FE",X"00",X"CA",X"DD",X"35",X"C3",X"6E",X"36",X"3A",
		X"6F",X"70",X"FE",X"01",X"28",X"09",X"3A",X"AC",X"70",X"FE",X"3C",X"CA",X"B5",X"3C",X"C9",X"3A",
		X"AD",X"70",X"FE",X"3C",X"C0",X"CD",X"56",X"32",X"CD",X"D5",X"3C",X"CD",X"E9",X"3C",X"AF",X"32",
		X"AD",X"70",X"21",X"71",X"70",X"34",X"DD",X"E1",X"CD",X"73",X"0D",X"22",X"62",X"73",X"21",X"C3",
		X"70",X"34",X"C3",X"18",X"36",X"CD",X"56",X"32",X"CD",X"D5",X"3C",X"CD",X"E9",X"3C",X"AF",X"32",
		X"AC",X"70",X"21",X"70",X"70",X"34",X"DD",X"E1",X"CD",X"73",X"0D",X"22",X"62",X"73",X"21",X"C2",
		X"70",X"34",X"C3",X"5B",X"35",X"21",X"0A",X"73",X"06",X"3C",X"36",X"00",X"23",X"10",X"FB",X"3A",
		X"33",X"70",X"2F",X"CB",X"4F",X"C0",X"DD",X"E1",X"C9",X"3A",X"6F",X"70",X"FE",X"00",X"20",X"0A",
		X"3A",X"C2",X"70",X"FE",X"0A",X"D2",X"88",X"3D",X"18",X"08",X"3A",X"C3",X"70",X"FE",X"0A",X"D2",
		X"88",X"3D",X"97",X"2A",X"50",X"73",X"11",X"F4",X"01",X"ED",X"52",X"22",X"50",X"73",X"22",X"46",
		X"73",X"97",X"2A",X"48",X"73",X"ED",X"52",X"22",X"48",X"73",X"97",X"2A",X"4C",X"73",X"ED",X"52",
		X"22",X"4C",X"73",X"22",X"4E",X"73",X"21",X"55",X"73",X"7E",X"FE",X"06",X"28",X"02",X"35",X"35",
		X"21",X"5A",X"73",X"7E",X"FE",X"08",X"28",X"02",X"35",X"35",X"21",X"5F",X"73",X"FE",X"08",X"28",
		X"02",X"35",X"35",X"3A",X"68",X"73",X"FE",X"02",X"28",X"08",X"3D",X"3D",X"32",X"68",X"73",X"32",
		X"5B",X"70",X"21",X"61",X"73",X"7E",X"FE",X"04",X"28",X"02",X"35",X"35",X"3A",X"64",X"73",X"D6",
		X"14",X"32",X"64",X"73",X"21",X"65",X"73",X"7E",X"FE",X"06",X"28",X"02",X"35",X"35",X"3A",X"69",
		X"73",X"FE",X"01",X"28",X"06",X"3C",X"32",X"69",X"73",X"18",X"0D",X"21",X"67",X"73",X"7E",X"FE",
		X"04",X"28",X"05",X"35",X"AF",X"32",X"69",X"73",X"AF",X"32",X"0D",X"74",X"32",X"11",X"74",X"32",
		X"15",X"74",X"32",X"19",X"74",X"32",X"1D",X"74",X"32",X"21",X"74",X"32",X"25",X"74",X"32",X"29",
		X"74",X"C9",X"DD",X"E5",X"FD",X"E1",X"11",X"00",X"10",X"FD",X"19",X"DD",X"36",X"00",X"0B",X"DD",
		X"36",X"01",X"09",X"DD",X"36",X"02",X"0D",X"FD",X"71",X"00",X"FD",X"71",X"01",X"FD",X"71",X"02",
		X"11",X"20",X"00",X"DD",X"19",X"FD",X"19",X"DD",X"36",X"00",X"06",X"DD",X"36",X"02",X"08",X"FD",
		X"71",X"00",X"FD",X"71",X"02",X"DD",X"19",X"FD",X"19",X"10",X"EC",X"FD",X"71",X"00",X"FD",X"71",
		X"01",X"FD",X"71",X"02",X"DD",X"36",X"00",X"0A",X"DD",X"36",X"01",X"07",X"DD",X"36",X"02",X"0C",
		X"C9",X"DD",X"E5",X"FD",X"E1",X"11",X"00",X"10",X"FD",X"19",X"DD",X"36",X"00",X"0B",X"DD",X"36",
		X"01",X"09",X"DD",X"36",X"02",X"09",X"DD",X"36",X"03",X"0D",X"FD",X"71",X"00",X"FD",X"71",X"01",
		X"FD",X"71",X"02",X"FD",X"71",X"03",X"11",X"20",X"00",X"DD",X"19",X"FD",X"19",X"DD",X"36",X"00",
		X"06",X"DD",X"36",X"03",X"08",X"FD",X"71",X"00",X"FD",X"71",X"03",X"DD",X"19",X"FD",X"19",X"10",
		X"EC",X"FD",X"71",X"00",X"FD",X"71",X"01",X"FD",X"71",X"02",X"FD",X"71",X"03",X"DD",X"36",X"00",
		X"0A",X"DD",X"36",X"01",X"07",X"DD",X"36",X"02",X"07",X"DD",X"36",X"03",X"0C",X"C9",X"06",X"1F",
		X"21",X"40",X"98",X"11",X"40",X"88",X"CD",X"93",X"3E",X"06",X"1F",X"21",X"A0",X"9B",X"11",X"A0",
		X"8B",X"CD",X"93",X"3E",X"21",X"40",X"98",X"11",X"40",X"88",X"06",X"1B",X"3E",X"9C",X"CD",X"9C",
		X"3E",X"06",X"1B",X"21",X"5E",X"98",X"11",X"5E",X"88",X"3E",X"9C",X"CD",X"9C",X"3E",X"21",X"40",
		X"88",X"36",X"A0",X"21",X"5E",X"88",X"36",X"9D",X"21",X"A0",X"8B",X"36",X"9F",X"21",X"BE",X"8B",
		X"36",X"9E",X"C9",X"3E",X"A1",X"71",X"12",X"23",X"13",X"10",X"FA",X"C9",X"71",X"12",X"F5",X"7D",
		X"C6",X"20",X"30",X"02",X"24",X"14",X"6F",X"5F",X"F1",X"10",X"F1",X"C9",X"3E",X"40",X"06",X"08",
		X"21",X"8E",X"99",X"11",X"8E",X"89",X"CD",X"D1",X"3E",X"3E",X"94",X"06",X"04",X"21",X"B8",X"99",
		X"11",X"B8",X"89",X"CD",X"D1",X"3E",X"3E",X"98",X"32",X"58",X"8A",X"3E",X"18",X"32",X"58",X"9A",
		X"C9",X"36",X"18",X"12",X"F5",X"7D",X"C6",X"20",X"30",X"02",X"24",X"14",X"6F",X"5F",X"F1",X"3C",
		X"10",X"EF",X"3A",X"00",X"A8",X"E6",X"20",X"FE",X"20",X"C0",X"3E",X"44",X"32",X"8E",X"89",X"C9",
		X"00",X"E5",X"7E",X"80",X"77",X"7E",X"FE",X"0A",X"38",X"0C",X"D6",X"0A",X"77",X"23",X"7E",X"FE",
		X"10",X"28",X"03",X"34",X"18",X"EF",X"06",X"06",X"11",X"20",X"00",X"21",X"E1",X"8A",X"DD",X"21",
		X"74",X"70",X"DD",X"7E",X"00",X"77",X"DD",X"23",X"19",X"10",X"F7",X"06",X"06",X"21",X"81",X"88",
		X"DD",X"23",X"DD",X"7E",X"00",X"77",X"DD",X"23",X"19",X"10",X"F7",X"E1",X"C9",X"CD",X"E0",X"40",
		X"21",X"A0",X"8B",X"11",X"E5",X"41",X"0E",X"07",X"CD",X"71",X"41",X"21",X"40",X"89",X"11",X"EF",
		X"41",X"0E",X"07",X"CD",X"71",X"41",X"21",X"81",X"8B",X"11",X"4C",X"42",X"0E",X"0C",X"CD",X"71",
		X"41",X"21",X"21",X"89",X"11",X"4C",X"42",X"0E",X"0C",X"CD",X"71",X"41",X"11",X"72",X"42",X"21",
		X"40",X"8A",X"0E",X"09",X"CD",X"71",X"41",X"CD",X"85",X"3F",X"21",X"9F",X"89",X"11",X"00",X"42",
		X"0E",X"0C",X"CD",X"71",X"41",X"3A",X"04",X"70",X"32",X"7F",X"88",X"3A",X"05",X"70",X"FE",X"00",
		X"C8",X"32",X"9F",X"88",X"C9",X"21",X"A1",X"89",X"11",X"0F",X"70",X"06",X"06",X"1A",X"77",X"7D",
		X"C6",X"20",X"30",X"01",X"24",X"6F",X"1B",X"10",X"F4",X"C9",X"21",X"2D",X"8A",X"11",X"AC",X"41",
		X"0E",X"05",X"CD",X"71",X"41",X"3A",X"05",X"70",X"FE",X"00",X"20",X"07",X"3A",X"04",X"70",X"FE",
		X"01",X"28",X"05",X"11",X"B2",X"41",X"18",X"03",X"11",X"D3",X"41",X"21",X"0E",X"8B",X"0E",X"05",
		X"CD",X"71",X"41",X"C9",X"00",X"DD",X"21",X"43",X"98",X"FD",X"21",X"43",X"88",X"06",X"05",X"C5",
		X"06",X"0E",X"DD",X"E5",X"FD",X"E5",X"FD",X"36",X"00",X"F9",X"FD",X"36",X"01",X"FA",X"FD",X"36",
		X"20",X"FB",X"FD",X"36",X"21",X"FC",X"DD",X"36",X"00",X"11",X"DD",X"36",X"01",X"11",X"DD",X"36",
		X"20",X"11",X"DD",X"36",X"21",X"11",X"11",X"40",X"00",X"DD",X"19",X"FD",X"19",X"10",X"D7",X"FD",
		X"E1",X"DD",X"E1",X"11",X"06",X"00",X"DD",X"19",X"FD",X"19",X"C1",X"10",X"C2",X"DD",X"21",X"C3",
		X"98",X"FD",X"21",X"C3",X"88",X"06",X"04",X"C5",X"06",X"0E",X"DD",X"E5",X"FD",X"E5",X"FD",X"36",
		X"00",X"B2",X"FD",X"36",X"01",X"B3",X"FD",X"36",X"20",X"B4",X"FD",X"36",X"21",X"B5",X"DD",X"36",
		X"00",X"11",X"DD",X"36",X"01",X"11",X"DD",X"36",X"20",X"11",X"DD",X"36",X"21",X"11",X"11",X"02",
		X"00",X"DD",X"19",X"FD",X"19",X"10",X"D7",X"FD",X"E1",X"DD",X"E1",X"11",X"C0",X"00",X"DD",X"19",
		X"FD",X"19",X"C1",X"10",X"C2",X"C9",X"DD",X"21",X"A3",X"88",X"06",X"05",X"C5",X"06",X"06",X"1A",
		X"CD",X"7B",X"40",X"13",X"DD",X"23",X"DD",X"23",X"DD",X"23",X"DD",X"23",X"DD",X"23",X"10",X"EF",
		X"D5",X"11",X"82",X"00",X"DD",X"19",X"D1",X"C1",X"10",X"E2",X"C9",X"DD",X"77",X"00",X"3C",X"DD",
		X"77",X"01",X"3C",X"DD",X"77",X"20",X"3C",X"DD",X"77",X"21",X"C9",X"CD",X"C4",X"3F",X"DD",X"21",
		X"A2",X"88",X"FD",X"21",X"A2",X"98",X"06",X"04",X"3E",X"A2",X"0E",X"11",X"C5",X"CD",X"AB",X"40",
		X"11",X"40",X"00",X"DD",X"19",X"FD",X"19",X"C1",X"10",X"EE",X"C9",X"06",X"04",X"C5",X"06",X"04",
		X"DD",X"77",X"00",X"FD",X"71",X"00",X"DD",X"77",X"06",X"FD",X"71",X"06",X"DD",X"77",X"0C",X"FD",
		X"71",X"0C",X"DD",X"77",X"12",X"FD",X"71",X"12",X"DD",X"77",X"18",X"FD",X"71",X"18",X"3C",X"DD",
		X"23",X"FD",X"23",X"10",X"DB",X"11",X"1C",X"00",X"DD",X"19",X"FD",X"19",X"C1",X"10",X"CE",X"C9",
		X"21",X"40",X"88",X"11",X"40",X"98",X"AF",X"36",X"10",X"12",X"23",X"13",X"7C",X"FE",X"8B",X"20",
		X"F5",X"7D",X"FE",X"C0",X"20",X"F0",X"21",X"1F",X"43",X"7E",X"FE",X"49",X"C8",X"DD",X"E1",X"C9",
		X"11",X"82",X"99",X"21",X"82",X"89",X"0E",X"00",X"06",X"08",X"3A",X"02",X"70",X"71",X"12",X"23",
		X"13",X"0C",X"10",X"F9",X"7D",X"FE",X"6A",X"C8",X"C6",X"18",X"30",X"01",X"24",X"6F",X"7B",X"C6",
		X"18",X"30",X"01",X"14",X"5F",X"18",X"E1",X"11",X"F1",X"98",X"21",X"F1",X"88",X"0E",X"48",X"06",
		X"04",X"3A",X"03",X"70",X"71",X"12",X"23",X"13",X"0C",X"10",X"F9",X"7D",X"FE",X"35",X"20",X"05",
		X"7C",X"FE",X"8B",X"C8",X"7D",X"C6",X"1C",X"30",X"01",X"24",X"6F",X"7B",X"C6",X"1C",X"30",X"01",
		X"14",X"5F",X"18",X"DB",X"21",X"42",X"88",X"11",X"42",X"98",X"0E",X"1C",X"AF",X"06",X"1E",X"36",
		X"10",X"12",X"23",X"13",X"10",X"F9",X"23",X"23",X"13",X"13",X"0D",X"79",X"FE",X"00",X"20",X"ED",
		X"C9",X"3A",X"00",X"A8",X"E6",X"20",X"FE",X"20",X"28",X"08",X"E5",X"EB",X"11",X"B2",X"01",X"19",
		X"EB",X"E1",X"1A",X"FE",X"3F",X"CA",X"9D",X"41",X"D6",X"30",X"77",X"06",X"10",X"E5",X"7C",X"80",
		X"67",X"71",X"E1",X"7D",X"DE",X"20",X"6F",X"30",X"01",X"25",X"13",X"18",X"E5",X"DD",X"21",X"AB",
		X"42",X"DD",X"7E",X"03",X"FE",X"49",X"C8",X"21",X"70",X"70",X"34",X"C9",X"50",X"55",X"53",X"48",
		X"40",X"3F",X"4F",X"4E",X"45",X"40",X"4F",X"52",X"40",X"40",X"54",X"57",X"4F",X"40",X"50",X"4C",
		X"41",X"59",X"45",X"52",X"53",X"3F",X"53",X"54",X"41",X"52",X"54",X"40",X"42",X"55",X"54",X"54",
		X"4F",X"4E",X"3F",X"40",X"4F",X"4E",X"4C",X"59",X"40",X"4F",X"4E",X"45",X"40",X"40",X"50",X"4C",
		X"41",X"59",X"45",X"52",X"3F",X"50",X"4C",X"41",X"59",X"45",X"52",X"40",X"31",X"40",X"3F",X"50",
		X"4C",X"41",X"59",X"45",X"52",X"40",X"32",X"40",X"3F",X"43",X"52",X"45",X"44",X"49",X"54",X"3F",
		X"43",X"52",X"45",X"44",X"49",X"54",X"53",X"40",X"40",X"40",X"3F",X"50",X"4C",X"41",X"59",X"45",
		X"52",X"40",X"40",X"40",X"54",X"57",X"4F",X"3F",X"50",X"4C",X"41",X"59",X"45",X"52",X"40",X"40",
		X"40",X"4F",X"4E",X"45",X"3F",X"52",X"45",X"41",X"44",X"59",X"40",X"54",X"4F",X"40",X"47",X"4F",
		X"3F",X"47",X"41",X"4D",X"45",X"40",X"4F",X"56",X"45",X"52",X"3F",X"40",X"40",X"49",X"4E",X"53",
		X"45",X"52",X"54",X"40",X"40",X"43",X"4F",X"49",X"4E",X"40",X"40",X"3F",X"30",X"30",X"30",X"30",
		X"30",X"30",X"3F",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",
		X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",
		X"40",X"3F",X"52",X"45",X"43",X"4F",X"52",X"44",X"3F",X"53",X"43",X"4F",X"52",X"45",X"40",X"40",
		X"40",X"4E",X"41",X"4D",X"45",X"40",X"40",X"3F",X"40",X"40",X"40",X"48",X"49",X"47",X"48",X"40",
		X"40",X"53",X"43",X"4F",X"52",X"45",X"40",X"40",X"40",X"3F",X"3D",X"40",X"43",X"4F",X"50",X"59",
		X"52",X"49",X"47",X"48",X"54",X"40",X"31",X"39",X"38",X"33",X"3F",X"42",X"59",X"40",X"49",X"54",
		X"49",X"53",X"41",X"40",X"50",X"41",X"4C",X"41",X"4D",X"4F",X"53",X"3F",X"53",X"50",X"41",X"49",
		X"4E",X"3F",X"40",X"57",X"52",X"49",X"54",X"45",X"40",X"3F",X"49",X"4E",X"43",X"52",X"5D",X"40",
		X"40",X"40",X"40",X"40",X"40",X"40",X"44",X"45",X"43",X"52",X"5D",X"3F",X"45",X"52",X"41",X"53",
		X"45",X"3F",X"40",X"40",X"4D",X"4F",X"56",X"45",X"40",X"4A",X"4F",X"59",X"53",X"54",X"49",X"43",
		X"4B",X"40",X"40",X"40",X"3F",X"54",X"4F",X"40",X"44",X"49",X"53",X"50",X"4C",X"41",X"59",X"40",
		X"59",X"4F",X"55",X"52",X"40",X"4E",X"41",X"4D",X"45",X"3F",X"45",X"4E",X"44",X"40",X"42",X"59",
		X"40",X"41",X"43",X"54",X"49",X"4F",X"4E",X"40",X"42",X"55",X"54",X"54",X"4F",X"4E",X"3F",X"49",
		X"40",X"54",X"40",X"49",X"40",X"53",X"40",X"41",X"40",X"40",X"50",X"41",X"4C",X"41",X"4D",X"4F",
		X"53",X"3F",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"50",X"55",
		X"4C",X"53",X"45",X"3F",X"55",X"4E",X"4F",X"40",X"4F",X"40",X"44",X"4F",X"53",X"40",X"4A",X"55",
		X"47",X"41",X"44",X"4F",X"52",X"45",X"53",X"3F",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",
		X"40",X"40",X"40",X"40",X"3F",X"40",X"53",X"4F",X"4C",X"4F",X"40",X"55",X"4E",X"40",X"40",X"4A",
		X"55",X"47",X"41",X"44",X"4F",X"52",X"3F",X"4A",X"55",X"47",X"41",X"44",X"4F",X"52",X"40",X"31",
		X"3F",X"4A",X"55",X"47",X"41",X"44",X"4F",X"52",X"40",X"32",X"3F",X"43",X"52",X"45",X"44",X"49",
		X"54",X"3F",X"43",X"52",X"45",X"44",X"49",X"54",X"53",X"40",X"40",X"40",X"3F",X"4A",X"55",X"47",
		X"41",X"44",X"4F",X"52",X"40",X"40",X"44",X"4F",X"53",X"3F",X"4A",X"55",X"47",X"41",X"44",X"4F",
		X"52",X"40",X"40",X"55",X"4E",X"4F",X"3F",X"40",X"40",X"40",X"4C",X"49",X"53",X"54",X"4F",X"40",
		X"40",X"40",X"3F",X"47",X"41",X"4D",X"45",X"40",X"4F",X"56",X"45",X"52",X"3F",X"49",X"4E",X"53",
		X"45",X"52",X"54",X"45",X"40",X"40",X"4D",X"4F",X"4E",X"45",X"44",X"41",X"53",X"3F",X"30",X"30",
		X"30",X"30",X"30",X"30",X"3F",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",
		X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",
		X"40",X"40",X"40",X"3F",X"52",X"45",X"43",X"4F",X"52",X"44",X"3F",X"50",X"55",X"4E",X"54",X"4F",
		X"53",X"40",X"40",X"4E",X"4F",X"4D",X"42",X"52",X"45",X"3F",X"4D",X"45",X"4A",X"4F",X"52",X"45",
		X"53",X"40",X"4A",X"55",X"47",X"41",X"44",X"4F",X"52",X"45",X"53",X"3F",X"3D",X"40",X"43",X"4F",
		X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"40",X"31",X"39",X"38",X"33",X"3F",X"42",X"59",X"40",
		X"49",X"54",X"49",X"53",X"41",X"40",X"50",X"41",X"4C",X"41",X"4D",X"4F",X"53",X"3F",X"53",X"50",
		X"41",X"49",X"4E",X"3F",X"40",X"47",X"52",X"41",X"42",X"41",X"40",X"3F",X"49",X"4E",X"43",X"52",
		X"5D",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"44",X"45",X"43",X"52",X"5D",X"3F",X"42",X"4F",
		X"52",X"52",X"41",X"3F",X"4D",X"4F",X"56",X"45",X"52",X"40",X"50",X"41",X"4C",X"41",X"4E",X"43",
		X"41",X"40",X"50",X"41",X"52",X"41",X"3F",X"40",X"49",X"4E",X"54",X"52",X"4F",X"44",X"55",X"43",
		X"49",X"52",X"40",X"40",X"4E",X"4F",X"4D",X"42",X"52",X"45",X"40",X"3F",X"46",X"49",X"4E",X"5C",
		X"40",X"42",X"4F",X"54",X"4F",X"4E",X"40",X"44",X"45",X"40",X"41",X"43",X"43",X"49",X"4F",X"4E",
		X"3F",X"49",X"40",X"54",X"40",X"49",X"40",X"53",X"40",X"41",X"40",X"40",X"50",X"41",X"4C",X"41",
		X"4D",X"4F",X"53",X"3F",X"3A",X"11",X"75",X"FE",X"00",X"C8",X"3A",X"11",X"75",X"FE",X"01",X"CA",
		X"33",X"45",X"FE",X"02",X"CA",X"49",X"45",X"FE",X"03",X"CA",X"7D",X"45",X"FE",X"04",X"CA",X"B1",
		X"45",X"FE",X"05",X"CA",X"D8",X"45",X"FE",X"06",X"CA",X"10",X"46",X"FE",X"07",X"CA",X"46",X"46",
		X"FE",X"08",X"CA",X"69",X"46",X"FE",X"09",X"CA",X"7F",X"46",X"FE",X"0A",X"CA",X"87",X"46",X"FE",
		X"0B",X"CA",X"AD",X"46",X"FE",X"0C",X"CA",X"C3",X"46",X"FE",X"0D",X"CA",X"F5",X"46",X"AF",X"32",
		X"11",X"75",X"C9",X"21",X"02",X"50",X"22",X"19",X"75",X"3E",X"0F",X"32",X"14",X"75",X"3E",X"01",
		X"32",X"03",X"75",X"32",X"06",X"75",X"C3",X"2E",X"45",X"21",X"A0",X"52",X"22",X"15",X"75",X"21",
		X"EC",X"52",X"22",X"17",X"75",X"21",X"38",X"53",X"22",X"19",X"75",X"3E",X"0F",X"32",X"12",X"75",
		X"32",X"13",X"75",X"32",X"14",X"75",X"3E",X"01",X"32",X"01",X"75",X"32",X"02",X"75",X"32",X"03",
		X"75",X"32",X"04",X"75",X"32",X"05",X"75",X"32",X"06",X"75",X"C3",X"2E",X"45",X"21",X"E8",X"4E",
		X"22",X"15",X"75",X"21",X"79",X"4F",X"22",X"17",X"75",X"21",X"B6",X"4F",X"22",X"19",X"75",X"3E",
		X"0F",X"32",X"12",X"75",X"32",X"13",X"75",X"32",X"14",X"75",X"3E",X"01",X"32",X"01",X"75",X"32",
		X"02",X"75",X"32",X"03",X"75",X"32",X"04",X"75",X"32",X"05",X"75",X"32",X"06",X"75",X"C3",X"2E",
		X"45",X"21",X"CB",X"4B",X"22",X"15",X"75",X"21",X"E8",X"4D",X"22",X"17",X"75",X"3E",X"0D",X"32",
		X"12",X"75",X"3E",X"0B",X"32",X"13",X"75",X"3E",X"01",X"32",X"01",X"75",X"32",X"02",X"75",X"32",
		X"04",X"75",X"32",X"05",X"75",X"C3",X"2E",X"45",X"21",X"42",X"50",X"22",X"15",X"75",X"21",X"9A",
		X"50",X"22",X"17",X"75",X"21",X"9D",X"51",X"22",X"19",X"75",X"3E",X"0E",X"32",X"12",X"75",X"3E",
		X"0F",X"32",X"13",X"75",X"3E",X"0F",X"32",X"14",X"75",X"3E",X"01",X"32",X"01",X"75",X"32",X"02",
		X"75",X"32",X"03",X"75",X"32",X"04",X"75",X"32",X"05",X"75",X"32",X"06",X"75",X"C3",X"2E",X"45",
		X"21",X"45",X"47",X"22",X"15",X"75",X"21",X"02",X"49",X"22",X"17",X"75",X"21",X"62",X"4A",X"22",
		X"19",X"75",X"3E",X"0A",X"32",X"12",X"75",X"3E",X"09",X"32",X"13",X"75",X"32",X"14",X"75",X"3E",
		X"01",X"32",X"01",X"75",X"32",X"02",X"75",X"32",X"03",X"75",X"32",X"04",X"75",X"32",X"05",X"75",
		X"32",X"06",X"75",X"C3",X"2E",X"45",X"21",X"29",X"47",X"22",X"19",X"75",X"22",X"17",X"75",X"22",
		X"15",X"75",X"3E",X"01",X"32",X"01",X"75",X"32",X"02",X"75",X"32",X"03",X"75",X"32",X"04",X"75",
		X"32",X"05",X"75",X"32",X"06",X"75",X"C3",X"2E",X"45",X"21",X"29",X"47",X"22",X"15",X"75",X"3E",
		X"01",X"32",X"01",X"75",X"32",X"04",X"75",X"21",X"2D",X"47",X"11",X"31",X"47",X"18",X"0E",X"21",
		X"35",X"47",X"11",X"39",X"47",X"18",X"06",X"21",X"3D",X"47",X"11",X"41",X"47",X"22",X"19",X"75",
		X"ED",X"53",X"17",X"75",X"3E",X"01",X"32",X"03",X"75",X"32",X"02",X"75",X"32",X"06",X"75",X"32",
		X"06",X"75",X"3E",X"0E",X"32",X"14",X"75",X"32",X"13",X"75",X"C3",X"2E",X"45",X"21",X"84",X"53",
		X"22",X"19",X"75",X"3E",X"01",X"32",X"03",X"75",X"32",X"06",X"75",X"3E",X"0F",X"32",X"14",X"75",
		X"C3",X"2E",X"45",X"21",X"A6",X"53",X"22",X"19",X"75",X"21",X"29",X"47",X"22",X"17",X"75",X"22",
		X"15",X"75",X"3E",X"01",X"32",X"03",X"75",X"32",X"02",X"75",X"32",X"01",X"75",X"32",X"06",X"75",
		X"32",X"04",X"75",X"32",X"05",X"75",X"3E",X"0F",X"32",X"14",X"75",X"AF",X"32",X"13",X"75",X"32",
		X"12",X"75",X"C3",X"2E",X"45",X"21",X"0D",X"54",X"22",X"15",X"75",X"21",X"59",X"54",X"22",X"17",
		X"75",X"21",X"A5",X"54",X"22",X"19",X"75",X"3E",X"0D",X"32",X"12",X"75",X"32",X"13",X"75",X"32",
		X"14",X"75",X"3E",X"01",X"32",X"01",X"75",X"32",X"02",X"75",X"32",X"03",X"75",X"32",X"04",X"75",
		X"32",X"05",X"75",X"32",X"06",X"75",X"C3",X"2E",X"45",X"00",X"00",X"01",X"FF",X"00",X"F5",X"12",
		X"FF",X"00",X"F4",X"12",X"FF",X"00",X"AD",X"12",X"FF",X"00",X"AC",X"12",X"FF",X"00",X"74",X"24",
		X"FF",X"00",X"73",X"24",X"FF",X"00",X"C2",X"06",X"00",X"D9",X"06",X"00",X"E7",X"06",X"00",X"D9",
		X"06",X"00",X"B8",X"18",X"00",X"A3",X"06",X"00",X"B8",X"06",X"00",X"C2",X"06",X"00",X"B8",X"06",
		X"00",X"92",X"18",X"00",X"89",X"06",X"00",X"92",X"06",X"00",X"9A",X"06",X"00",X"92",X"06",X"00",
		X"61",X"06",X"00",X"6D",X"06",X"00",X"74",X"06",X"00",X"6D",X"06",X"00",X"61",X"06",X"00",X"6D",
		X"06",X"00",X"74",X"06",X"00",X"6D",X"06",X"00",X"5C",X"18",X"00",X"6D",X"0C",X"00",X"5C",X"0C",
		X"00",X"61",X"0C",X"00",X"6D",X"0C",X"00",X"7B",X"0C",X"00",X"6D",X"0C",X"00",X"61",X"0C",X"00",
		X"6D",X"0C",X"00",X"7B",X"0C",X"00",X"6D",X"0C",X"00",X"61",X"0C",X"00",X"6D",X"0C",X"00",X"7B",
		X"0C",X"00",X"82",X"0C",X"00",X"92",X"18",X"00",X"92",X"0C",X"00",X"89",X"0C",X"00",X"7B",X"0C",
		X"00",X"7B",X"0C",X"00",X"6D",X"06",X"00",X"7B",X"06",X"00",X"89",X"06",X"00",X"92",X"06",X"00",
		X"A3",X"18",X"00",X"92",X"0C",X"00",X"89",X"0C",X"00",X"7B",X"0C",X"00",X"7B",X"0C",X"00",X"6D",
		X"06",X"00",X"7B",X"06",X"00",X"89",X"06",X"00",X"92",X"06",X"00",X"A3",X"18",X"00",X"B8",X"0C",
		X"00",X"A3",X"0C",X"00",X"92",X"0C",X"00",X"92",X"0C",X"00",X"89",X"06",X"00",X"92",X"06",X"00",
		X"A3",X"06",X"00",X"B8",X"06",X"00",X"C2",X"18",X"00",X"B8",X"0C",X"00",X"A3",X"0C",X"00",X"92",
		X"0C",X"00",X"92",X"0C",X"00",X"89",X"06",X"00",X"92",X"06",X"00",X"A3",X"06",X"00",X"B8",X"06",
		X"00",X"C2",X"18",X"00",X"C2",X"06",X"00",X"D9",X"06",X"00",X"E7",X"06",X"00",X"D9",X"06",X"00",
		X"B8",X"18",X"00",X"A3",X"06",X"00",X"B8",X"06",X"00",X"C2",X"06",X"00",X"B8",X"06",X"00",X"92",
		X"18",X"00",X"89",X"06",X"00",X"92",X"06",X"00",X"9A",X"06",X"00",X"92",X"06",X"00",X"61",X"06",
		X"00",X"6D",X"06",X"00",X"74",X"06",X"00",X"6D",X"06",X"00",X"61",X"06",X"00",X"6D",X"06",X"00",
		X"74",X"06",X"00",X"6D",X"06",X"00",X"5C",X"18",X"00",X"6D",X"0C",X"00",X"5C",X"0C",X"00",X"61",
		X"0C",X"00",X"6D",X"0C",X"00",X"7B",X"0C",X"00",X"6D",X"0C",X"00",X"61",X"0C",X"00",X"6D",X"0C",
		X"00",X"7B",X"0C",X"00",X"6D",X"0C",X"00",X"61",X"0C",X"00",X"6D",X"0C",X"00",X"7B",X"0C",X"00",
		X"82",X"0C",X"00",X"92",X"18",X"00",X"92",X"0C",X"00",X"89",X"0C",X"00",X"7B",X"0C",X"00",X"7B",
		X"0C",X"00",X"6D",X"06",X"00",X"7B",X"06",X"00",X"89",X"06",X"00",X"92",X"06",X"00",X"A3",X"18",
		X"00",X"92",X"0C",X"00",X"89",X"0C",X"00",X"7B",X"0C",X"00",X"7B",X"0C",X"00",X"6D",X"06",X"00",
		X"7B",X"06",X"00",X"89",X"06",X"00",X"92",X"06",X"00",X"A3",X"18",X"00",X"B8",X"0C",X"00",X"A3",
		X"0C",X"00",X"92",X"0C",X"00",X"92",X"0C",X"00",X"89",X"06",X"00",X"92",X"06",X"00",X"A3",X"06",
		X"00",X"B8",X"06",X"00",X"C2",X"18",X"00",X"B8",X"0C",X"00",X"A3",X"0C",X"00",X"92",X"0C",X"00",
		X"92",X"0C",X"00",X"89",X"06",X"00",X"92",X"06",X"00",X"A3",X"06",X"00",X"B8",X"06",X"00",X"C2",
		X"18",X"FF",X"00",X"00",X"18",X"00",X"00",X"0C",X"00",X"92",X"0C",X"00",X"00",X"0C",X"00",X"92",
		X"0C",X"00",X"00",X"0C",X"00",X"92",X"0C",X"00",X"00",X"0C",X"00",X"92",X"0C",X"00",X"00",X"0C",
		X"00",X"92",X"0C",X"00",X"00",X"0C",X"00",X"92",X"0C",X"00",X"00",X"0C",X"00",X"92",X"0C",X"00",
		X"00",X"0C",X"00",X"92",X"0C",X"00",X"00",X"0C",X"00",X"C2",X"0C",X"00",X"00",X"0C",X"00",X"C2",
		X"0C",X"00",X"00",X"0C",X"00",X"C2",X"0C",X"00",X"00",X"0C",X"00",X"C2",X"0C",X"00",X"00",X"0C",
		X"00",X"C2",X"0C",X"00",X"00",X"0C",X"00",X"C2",X"0C",X"00",X"00",X"30",X"00",X"00",X"0C",X"00",
		X"F5",X"0C",X"00",X"00",X"0C",X"00",X"F5",X"0C",X"00",X"00",X"0C",X"00",X"F5",X"0C",X"00",X"00",
		X"0C",X"00",X"F5",X"0C",X"00",X"00",X"0C",X"00",X"F5",X"0C",X"00",X"00",X"0C",X"00",X"F5",X"0C",
		X"00",X"00",X"0C",X"00",X"F5",X"0C",X"00",X"00",X"0C",X"00",X"F5",X"0C",X"00",X"00",X"0C",X"00",
		X"92",X"0C",X"00",X"00",X"0C",X"00",X"92",X"0C",X"00",X"00",X"0C",X"00",X"92",X"0C",X"00",X"00",
		X"0C",X"00",X"92",X"0C",X"00",X"00",X"0C",X"00",X"92",X"0C",X"00",X"00",X"0C",X"00",X"92",X"0C",
		X"00",X"00",X"30",X"00",X"00",X"0C",X"00",X"92",X"0C",X"00",X"00",X"0C",X"00",X"92",X"0C",X"00",
		X"00",X"0C",X"00",X"92",X"0C",X"00",X"00",X"0C",X"00",X"92",X"0C",X"00",X"00",X"0C",X"00",X"92",
		X"0C",X"00",X"00",X"0C",X"00",X"92",X"0C",X"00",X"00",X"0C",X"00",X"92",X"0C",X"00",X"00",X"0C",
		X"00",X"92",X"0C",X"00",X"00",X"0C",X"00",X"C2",X"0C",X"00",X"00",X"0C",X"00",X"C2",X"0C",X"00",
		X"00",X"0C",X"00",X"C2",X"0C",X"00",X"00",X"0C",X"00",X"C2",X"0C",X"00",X"00",X"0C",X"00",X"C2",
		X"0C",X"00",X"00",X"0C",X"00",X"C2",X"0C",X"00",X"00",X"30",X"00",X"00",X"0C",X"00",X"F5",X"0C",
		X"00",X"00",X"0C",X"00",X"F5",X"0C",X"00",X"00",X"0C",X"00",X"F5",X"0C",X"00",X"00",X"0C",X"00",
		X"F5",X"0C",X"00",X"00",X"0C",X"00",X"F5",X"0C",X"00",X"00",X"0C",X"00",X"F5",X"0C",X"00",X"00",
		X"0C",X"00",X"F5",X"0C",X"00",X"00",X"0C",X"00",X"F5",X"0C",X"00",X"00",X"0C",X"00",X"92",X"0C",
		X"00",X"00",X"0C",X"00",X"92",X"0C",X"00",X"00",X"0C",X"00",X"92",X"0C",X"00",X"00",X"0C",X"00",
		X"92",X"0C",X"00",X"00",X"0C",X"00",X"92",X"0C",X"00",X"00",X"0C",X"00",X"92",X"0C",X"00",X"00",
		X"18",X"FF",X"00",X"00",X"18",X"00",X"D9",X"0C",X"00",X"B8",X"0C",X"00",X"D9",X"0C",X"00",X"B8",
		X"0C",X"00",X"D9",X"0C",X"00",X"B8",X"0C",X"00",X"D9",X"0C",X"00",X"B8",X"0C",X"00",X"D9",X"0C",
		X"00",X"B8",X"0C",X"00",X"D9",X"0C",X"00",X"B8",X"0C",X"00",X"D9",X"0C",X"00",X"B8",X"0C",X"00",
		X"D9",X"0C",X"00",X"B8",X"0C",X"01",X"23",X"0C",X"00",X"F5",X"0C",X"01",X"23",X"0C",X"00",X"F5",
		X"0C",X"01",X"23",X"0C",X"00",X"F5",X"0C",X"01",X"23",X"0C",X"00",X"F5",X"0C",X"01",X"35",X"0C",
		X"01",X"04",X"0C",X"01",X"35",X"0C",X"01",X"04",X"0C",X"01",X"23",X"18",X"00",X"00",X"18",X"01",
		X"70",X"0C",X"01",X"23",X"0C",X"01",X"70",X"0C",X"01",X"23",X"0C",X"01",X"48",X"0C",X"01",X"13",
		X"0C",X"01",X"48",X"0C",X"01",X"13",X"0C",X"01",X"70",X"0C",X"01",X"23",X"0C",X"01",X"70",X"0C",
		X"01",X"23",X"0C",X"01",X"48",X"0C",X"01",X"13",X"0C",X"01",X"48",X"0C",X"01",X"13",X"0C",X"00",
		X"D9",X"0C",X"00",X"B8",X"0C",X"00",X"D9",X"0C",X"00",X"B8",X"0C",X"00",X"E7",X"0C",X"00",X"C2",
		X"0C",X"00",X"E7",X"0C",X"00",X"C2",X"0C",X"00",X"D9",X"0C",X"00",X"B8",X"0C",X"00",X"D9",X"0C",
		X"00",X"B8",X"0C",X"00",X"E7",X"18",X"00",X"00",X"18",X"00",X"D9",X"0C",X"00",X"B8",X"0C",X"00",
		X"D9",X"0C",X"00",X"B8",X"0C",X"00",X"D9",X"0C",X"00",X"B8",X"0C",X"00",X"D9",X"0C",X"00",X"B8",
		X"0C",X"00",X"D9",X"0C",X"00",X"B8",X"0C",X"00",X"D9",X"0C",X"00",X"B8",X"0C",X"00",X"D9",X"0C",
		X"00",X"B8",X"0C",X"00",X"D9",X"0C",X"00",X"B8",X"0C",X"01",X"23",X"0C",X"00",X"F5",X"0C",X"01",
		X"23",X"0C",X"00",X"F5",X"0C",X"01",X"23",X"0C",X"00",X"F5",X"0C",X"01",X"23",X"0C",X"00",X"F5",
		X"0C",X"01",X"35",X"0C",X"01",X"04",X"0C",X"01",X"35",X"0C",X"01",X"04",X"0C",X"01",X"23",X"18",
		X"00",X"00",X"18",X"01",X"70",X"0C",X"01",X"23",X"0C",X"01",X"70",X"0C",X"01",X"23",X"0C",X"01",
		X"48",X"0C",X"01",X"13",X"0C",X"01",X"48",X"0C",X"01",X"13",X"0C",X"01",X"70",X"0C",X"01",X"23",
		X"0C",X"01",X"70",X"0C",X"01",X"23",X"0C",X"01",X"48",X"0C",X"01",X"13",X"0C",X"01",X"48",X"0C",
		X"01",X"13",X"0C",X"00",X"D9",X"0C",X"00",X"B8",X"0C",X"00",X"D9",X"0C",X"00",X"B8",X"0C",X"00",
		X"E7",X"0C",X"00",X"C2",X"0C",X"00",X"E7",X"0C",X"00",X"C2",X"0C",X"00",X"D9",X"0C",X"00",X"B8",
		X"0C",X"00",X"D9",X"0C",X"00",X"B8",X"0C",X"00",X"00",X"18",X"FF",X"01",X"70",X"04",X"00",X"00",
		X"02",X"01",X"13",X"04",X"00",X"00",X"02",X"00",X"D9",X"10",X"00",X"00",X"02",X"00",X"D9",X"04",
		X"00",X"00",X"02",X"00",X"D9",X"0A",X"00",X"00",X"02",X"01",X"70",X"04",X"00",X"00",X"02",X"01",
		X"13",X"04",X"00",X"00",X"02",X"00",X"D9",X"10",X"00",X"00",X"02",X"00",X"D9",X"04",X"00",X"00",
		X"02",X"00",X"D9",X"0A",X"00",X"00",X"02",X"01",X"70",X"04",X"00",X"00",X"02",X"01",X"13",X"04",
		X"00",X"00",X"02",X"00",X"D9",X"10",X"00",X"00",X"02",X"00",X"D9",X"04",X"00",X"00",X"02",X"00",
		X"D9",X"0A",X"00",X"00",X"02",X"00",X"F5",X"04",X"00",X"00",X"02",X"00",X"D9",X"04",X"00",X"00",
		X"02",X"00",X"A3",X"16",X"00",X"00",X"02",X"00",X"B8",X"16",X"00",X"00",X"02",X"00",X"CE",X"10",
		X"00",X"00",X"02",X"01",X"70",X"04",X"00",X"00",X"02",X"01",X"70",X"10",X"00",X"00",X"02",X"00",
		X"CE",X"04",X"00",X"00",X"02",X"00",X"D9",X"10",X"00",X"00",X"02",X"01",X"13",X"04",X"00",X"00",
		X"02",X"01",X"13",X"10",X"00",X"00",X"02",X"00",X"D9",X"04",X"00",X"00",X"02",X"00",X"F5",X"0A",
		X"00",X"00",X"02",X"00",X"D9",X"04",X"00",X"00",X"02",X"00",X"F5",X"04",X"00",X"00",X"02",X"01",
		X"13",X"0A",X"00",X"00",X"02",X"01",X"23",X"04",X"00",X"00",X"02",X"01",X"13",X"04",X"00",X"00",
		X"02",X"00",X"F5",X"22",X"00",X"00",X"02",X"01",X"70",X"04",X"00",X"00",X"02",X"01",X"13",X"04",
		X"00",X"00",X"02",X"00",X"D9",X"10",X"00",X"00",X"02",X"00",X"D9",X"04",X"00",X"00",X"02",X"00",
		X"D9",X"0A",X"00",X"00",X"02",X"01",X"70",X"04",X"00",X"00",X"02",X"01",X"13",X"04",X"00",X"00",
		X"02",X"00",X"D9",X"10",X"00",X"00",X"02",X"00",X"D9",X"04",X"00",X"00",X"02",X"00",X"D9",X"0A",
		X"00",X"00",X"02",X"01",X"70",X"04",X"00",X"00",X"02",X"01",X"13",X"04",X"00",X"00",X"02",X"00",
		X"D9",X"10",X"00",X"00",X"02",X"00",X"D9",X"04",X"00",X"00",X"02",X"00",X"D9",X"0A",X"00",X"00",
		X"02",X"00",X"F5",X"04",X"00",X"00",X"02",X"00",X"D9",X"04",X"00",X"00",X"02",X"00",X"A3",X"16",
		X"00",X"00",X"02",X"00",X"B8",X"16",X"00",X"00",X"02",X"00",X"CE",X"10",X"00",X"00",X"02",X"01",
		X"70",X"04",X"00",X"00",X"02",X"01",X"70",X"10",X"00",X"00",X"02",X"00",X"CE",X"04",X"00",X"00",
		X"02",X"00",X"D9",X"10",X"00",X"00",X"02",X"01",X"13",X"04",X"00",X"00",X"02",X"01",X"13",X"10",
		X"00",X"00",X"02",X"00",X"D9",X"04",X"00",X"00",X"02",X"00",X"F5",X"0A",X"00",X"00",X"02",X"00",
		X"D9",X"04",X"00",X"00",X"02",X"00",X"F5",X"04",X"00",X"00",X"02",X"01",X"13",X"0A",X"00",X"00",
		X"02",X"01",X"23",X"04",X"00",X"00",X"02",X"00",X"F5",X"04",X"00",X"00",X"02",X"01",X"13",X"16",
		X"00",X"00",X"02",X"01",X"13",X"10",X"00",X"00",X"02",X"01",X"13",X"04",X"00",X"00",X"02",X"01",
		X"13",X"16",X"00",X"00",X"02",X"01",X"23",X"10",X"00",X"00",X"02",X"01",X"13",X"04",X"00",X"00",
		X"02",X"00",X"F5",X"16",X"00",X"00",X"02",X"01",X"13",X"10",X"00",X"00",X"02",X"00",X"F5",X"04",
		X"00",X"00",X"02",X"00",X"D9",X"16",X"00",X"00",X"02",X"00",X"F5",X"10",X"00",X"00",X"02",X"00",
		X"D9",X"04",X"00",X"00",X"02",X"00",X"CE",X"0A",X"00",X"00",X"02",X"00",X"D9",X"04",X"00",X"00",
		X"02",X"00",X"F5",X"04",X"00",X"00",X"02",X"01",X"13",X"0A",X"00",X"00",X"02",X"00",X"D9",X"0A",
		X"00",X"00",X"02",X"00",X"F5",X"0A",X"00",X"00",X"02",X"00",X"B8",X"04",X"00",X"00",X"02",X"00",
		X"B8",X"04",X"00",X"00",X"02",X"00",X"B8",X"0A",X"00",X"00",X"02",X"01",X"70",X"04",X"00",X"00",
		X"02",X"01",X"13",X"04",X"00",X"00",X"02",X"FF",X"00",X"00",X"0C",X"01",X"13",X"16",X"00",X"00",
		X"02",X"01",X"13",X"16",X"00",X"00",X"02",X"01",X"13",X"16",X"00",X"00",X"02",X"01",X"13",X"16",
		X"00",X"00",X"02",X"01",X"13",X"16",X"00",X"00",X"02",X"01",X"13",X"16",X"00",X"00",X"02",X"01",
		X"13",X"16",X"00",X"00",X"02",X"01",X"13",X"16",X"00",X"00",X"02",X"01",X"23",X"16",X"00",X"00",
		X"02",X"01",X"23",X"16",X"00",X"00",X"02",X"01",X"13",X"16",X"00",X"00",X"02",X"00",X"D9",X"16",
		X"00",X"00",X"02",X"00",X"CE",X"16",X"00",X"00",X"02",X"00",X"D9",X"16",X"00",X"00",X"02",X"01",
		X"23",X"16",X"00",X"00",X"02",X"01",X"23",X"16",X"00",X"00",X"02",X"01",X"13",X"16",X"00",X"00",
		X"02",X"01",X"13",X"16",X"00",X"00",X"02",X"01",X"13",X"16",X"00",X"00",X"02",X"01",X"13",X"16",
		X"00",X"00",X"02",X"01",X"13",X"16",X"00",X"00",X"02",X"01",X"13",X"16",X"00",X"00",X"02",X"01",
		X"13",X"16",X"00",X"00",X"02",X"01",X"13",X"16",X"00",X"00",X"02",X"01",X"23",X"16",X"00",X"00",
		X"02",X"01",X"23",X"16",X"00",X"00",X"02",X"01",X"13",X"16",X"00",X"00",X"02",X"00",X"D9",X"16",
		X"00",X"00",X"02",X"00",X"CE",X"16",X"00",X"00",X"02",X"00",X"D9",X"16",X"00",X"00",X"02",X"00",
		X"D9",X"16",X"00",X"00",X"02",X"00",X"D9",X"10",X"00",X"00",X"02",X"00",X"D9",X"04",X"00",X"00",
		X"02",X"00",X"D9",X"16",X"00",X"00",X"02",X"00",X"00",X"18",X"01",X"23",X"16",X"00",X"00",X"02",
		X"01",X"70",X"16",X"00",X"00",X"02",X"01",X"23",X"16",X"00",X"00",X"02",X"01",X"70",X"16",X"00",
		X"00",X"02",X"00",X"F5",X"16",X"00",X"00",X"02",X"01",X"70",X"16",X"00",X"00",X"02",X"01",X"23",
		X"16",X"00",X"00",X"02",X"00",X"00",X"18",X"FF",X"00",X"B8",X"0A",X"00",X"00",X"02",X"00",X"D9",
		X"0A",X"00",X"00",X"02",X"00",X"F5",X"0A",X"00",X"00",X"02",X"00",X"B8",X"0A",X"00",X"00",X"02",
		X"00",X"D9",X"0A",X"00",X"00",X"02",X"00",X"F5",X"0A",X"00",X"00",X"02",X"00",X"B8",X"0A",X"00",
		X"00",X"02",X"00",X"D9",X"0A",X"00",X"00",X"02",X"00",X"A3",X"0A",X"00",X"00",X"02",X"00",X"D9",
		X"0A",X"00",X"00",X"02",X"00",X"F5",X"0A",X"00",X"00",X"02",X"00",X"A3",X"0A",X"00",X"00",X"02",
		X"00",X"D9",X"0A",X"00",X"00",X"02",X"00",X"F5",X"0A",X"00",X"00",X"02",X"00",X"A3",X"0A",X"00",
		X"00",X"02",X"00",X"F5",X"0A",X"00",X"00",X"02",X"00",X"B8",X"16",X"00",X"00",X"02",X"00",X"92",
		X"0A",X"00",X"00",X"02",X"00",X"B8",X"0A",X"00",X"00",X"02",X"00",X"D9",X"16",X"00",X"00",X"02",
		X"00",X"F5",X"16",X"00",X"00",X"02",X"00",X"00",X"18",X"00",X"C2",X"16",X"00",X"00",X"02",X"00",
		X"B8",X"16",X"00",X"00",X"02",X"00",X"00",X"18",X"FF",X"00",X"F5",X"16",X"00",X"00",X"02",X"00",
		X"00",X"18",X"00",X"00",X"18",X"00",X"F5",X"16",X"00",X"00",X"02",X"00",X"F5",X"16",X"00",X"00",
		X"02",X"00",X"00",X"18",X"00",X"00",X"18",X"00",X"00",X"18",X"00",X"F5",X"16",X"00",X"00",X"02",
		X"00",X"00",X"48",X"00",X"00",X"18",X"00",X"F5",X"16",X"00",X"00",X"02",X"00",X"F5",X"16",X"00",
		X"00",X"02",X"00",X"00",X"18",X"FF",X"01",X"23",X"16",X"00",X"00",X"02",X"01",X"23",X"16",X"00",
		X"00",X"02",X"01",X"23",X"16",X"00",X"00",X"02",X"01",X"23",X"16",X"00",X"00",X"02",X"01",X"13",
		X"16",X"00",X"00",X"02",X"01",X"13",X"16",X"00",X"00",X"02",X"01",X"13",X"16",X"00",X"00",X"02",
		X"01",X"13",X"16",X"00",X"00",X"02",X"01",X"23",X"16",X"00",X"00",X"02",X"00",X"00",X"48",X"00",
		X"00",X"18",X"01",X"13",X"16",X"00",X"00",X"02",X"01",X"23",X"16",X"00",X"00",X"02",X"00",X"00",
		X"18",X"FF",X"03",X"B3",X"01",X"00",X"00",X"01",X"02",X"C5",X"01",X"00",X"00",X"01",X"02",X"32",
		X"01",X"00",X"00",X"01",X"01",X"D9",X"01",X"00",X"00",X"01",X"01",X"62",X"01",X"00",X"00",X"01",
		X"01",X"19",X"01",X"00",X"00",X"01",X"00",X"EE",X"01",X"00",X"00",X"01",X"00",X"B1",X"01",X"00",
		X"00",X"01",X"00",X"8D",X"01",X"00",X"00",X"01",X"00",X"76",X"01",X"00",X"00",X"01",X"00",X"59",
		X"01",X"FF",X"00",X"F5",X"18",X"00",X"7B",X"30",X"00",X"92",X"06",X"00",X"A3",X"06",X"00",X"92",
		X"06",X"00",X"89",X"06",X"00",X"7B",X"18",X"00",X"92",X"18",X"00",X"B8",X"18",X"00",X"5C",X"30",
		X"00",X"6D",X"06",X"00",X"7B",X"06",X"00",X"6D",X"06",X"00",X"61",X"06",X"00",X"5C",X"18",X"00",
		X"6D",X"18",X"00",X"89",X"18",X"00",X"7B",X"30",X"00",X"92",X"06",X"00",X"A3",X"06",X"00",X"92",
		X"06",X"00",X"89",X"06",X"00",X"7B",X"18",X"00",X"92",X"18",X"00",X"B8",X"18",X"00",X"A3",X"18",
		X"00",X"B8",X"18",X"00",X"C2",X"18",X"00",X"B8",X"18",X"FF",X"00",X"00",X"18",X"01",X"23",X"0A",
		X"00",X"00",X"02",X"01",X"23",X"0A",X"00",X"00",X"02",X"01",X"23",X"0A",X"00",X"00",X"02",X"01",
		X"23",X"0A",X"00",X"00",X"02",X"01",X"23",X"0A",X"00",X"00",X"02",X"01",X"23",X"0A",X"00",X"00",
		X"02",X"01",X"23",X"0A",X"00",X"00",X"02",X"01",X"23",X"0A",X"00",X"00",X"02",X"01",X"23",X"0A",
		X"00",X"00",X"02",X"01",X"23",X"0A",X"00",X"00",X"02",X"01",X"23",X"0A",X"00",X"00",X"02",X"01",
		X"23",X"0A",X"00",X"00",X"02",X"00",X"D9",X"0A",X"00",X"00",X"02",X"00",X"D9",X"0A",X"00",X"00",
		X"02",X"00",X"D9",X"0A",X"00",X"00",X"02",X"00",X"D9",X"0A",X"00",X"00",X"02",X"00",X"D9",X"0A",
		X"00",X"00",X"02",X"00",X"D9",X"0A",X"00",X"00",X"02",X"00",X"D9",X"0A",X"00",X"00",X"02",X"00",
		X"D9",X"0A",X"00",X"00",X"02",X"00",X"D9",X"0A",X"00",X"00",X"02",X"00",X"D9",X"0A",X"00",X"00",
		X"02",X"00",X"D9",X"0A",X"00",X"00",X"02",X"00",X"D9",X"0A",X"00",X"00",X"02",X"01",X"23",X"0A",
		X"00",X"00",X"02",X"01",X"23",X"0A",X"00",X"00",X"02",X"01",X"23",X"0A",X"00",X"00",X"02",X"01",
		X"23",X"0A",X"00",X"00",X"02",X"01",X"23",X"0A",X"00",X"00",X"02",X"01",X"23",X"0A",X"00",X"00",
		X"02",X"01",X"23",X"0A",X"00",X"00",X"02",X"01",X"23",X"0A",X"00",X"00",X"02",X"01",X"23",X"0A",
		X"00",X"00",X"02",X"01",X"23",X"0A",X"00",X"00",X"02",X"01",X"23",X"0A",X"00",X"00",X"02",X"01",
		X"23",X"0A",X"00",X"00",X"02",X"00",X"C2",X"0A",X"00",X"00",X"02",X"00",X"C2",X"0A",X"00",X"00",
		X"02",X"00",X"89",X"0A",X"00",X"00",X"02",X"00",X"89",X"0A",X"00",X"00",X"02",X"00",X"A3",X"0A",
		X"00",X"00",X"02",X"00",X"A3",X"0A",X"00",X"00",X"02",X"01",X"70",X"18",X"FF",X"00",X"00",X"18",
		X"01",X"70",X"0A",X"00",X"00",X"02",X"01",X"70",X"0A",X"00",X"00",X"02",X"01",X"70",X"0A",X"00",
		X"00",X"02",X"01",X"70",X"0A",X"00",X"00",X"02",X"01",X"70",X"0A",X"00",X"00",X"02",X"01",X"70",
		X"0A",X"00",X"00",X"02",X"01",X"70",X"0A",X"00",X"00",X"02",X"01",X"70",X"0A",X"00",X"00",X"02",
		X"01",X"70",X"0A",X"00",X"00",X"02",X"01",X"70",X"0A",X"00",X"00",X"02",X"01",X"70",X"0A",X"00",
		X"00",X"02",X"01",X"70",X"0A",X"00",X"00",X"02",X"01",X"13",X"0A",X"00",X"00",X"02",X"01",X"13",
		X"0A",X"00",X"00",X"02",X"01",X"13",X"0A",X"00",X"00",X"02",X"01",X"13",X"0A",X"00",X"00",X"02",
		X"01",X"13",X"0A",X"00",X"00",X"02",X"01",X"13",X"0A",X"00",X"00",X"02",X"01",X"13",X"0A",X"00",
		X"00",X"02",X"01",X"13",X"0A",X"00",X"00",X"02",X"01",X"13",X"0A",X"00",X"00",X"02",X"01",X"13",
		X"0A",X"00",X"00",X"02",X"01",X"13",X"0A",X"00",X"00",X"02",X"01",X"13",X"0A",X"00",X"00",X"02",
		X"01",X"70",X"0A",X"00",X"00",X"02",X"01",X"70",X"0A",X"00",X"00",X"02",X"01",X"70",X"0A",X"00",
		X"00",X"02",X"01",X"70",X"0A",X"00",X"00",X"02",X"01",X"70",X"0A",X"00",X"00",X"02",X"01",X"70",
		X"0A",X"00",X"00",X"02",X"01",X"70",X"0A",X"00",X"00",X"02",X"01",X"70",X"0A",X"00",X"00",X"02",
		X"01",X"70",X"0A",X"00",X"00",X"02",X"01",X"70",X"0A",X"00",X"00",X"02",X"01",X"70",X"0A",X"00",
		X"00",X"02",X"01",X"70",X"0A",X"00",X"00",X"02",X"00",X"F5",X"0A",X"00",X"00",X"02",X"00",X"F5",
		X"0A",X"00",X"00",X"02",X"00",X"A3",X"0A",X"00",X"00",X"02",X"00",X"A3",X"0A",X"00",X"00",X"02",
		X"00",X"C2",X"0A",X"00",X"00",X"02",X"00",X"C2",X"0A",X"00",X"00",X"02",X"01",X"23",X"18",X"FF",
		X"00",X"89",X"0E",X"00",X"00",X"02",X"00",X"89",X"06",X"00",X"00",X"02",X"00",X"89",X"06",X"00",
		X"00",X"02",X"00",X"89",X"2E",X"00",X"00",X"02",X"00",X"89",X"06",X"00",X"00",X"02",X"00",X"89",
		X"06",X"00",X"00",X"02",X"00",X"89",X"0E",X"00",X"00",X"02",X"00",X"B8",X"0E",X"00",X"00",X"02",
		X"00",X"89",X"0E",X"00",X"00",X"02",X"00",X"6D",X"0E",X"00",X"00",X"02",X"00",X"5C",X"16",X"00",
		X"00",X"02",X"00",X"7B",X"06",X"00",X"00",X"02",X"00",X"7B",X"40",X"FF",X"00",X"B8",X"0E",X"00",
		X"00",X"02",X"00",X"B8",X"06",X"00",X"00",X"02",X"00",X"B8",X"06",X"00",X"00",X"02",X"00",X"B8",
		X"2E",X"00",X"00",X"02",X"00",X"B8",X"06",X"00",X"00",X"02",X"00",X"B8",X"06",X"00",X"00",X"02",
		X"00",X"B8",X"0E",X"00",X"00",X"02",X"00",X"D9",X"0E",X"00",X"00",X"02",X"00",X"B8",X"0E",X"00",
		X"00",X"02",X"00",X"89",X"0E",X"00",X"00",X"02",X"00",X"7B",X"16",X"00",X"00",X"02",X"00",X"92",
		X"06",X"00",X"00",X"02",X"00",X"92",X"40",X"FF",X"00",X"D9",X"0E",X"00",X"00",X"02",X"00",X"D9",
		X"06",X"00",X"00",X"02",X"00",X"D9",X"06",X"00",X"00",X"02",X"00",X"D9",X"2E",X"00",X"00",X"02",
		X"00",X"D9",X"06",X"00",X"00",X"02",X"00",X"D9",X"06",X"00",X"00",X"02",X"00",X"D9",X"0E",X"00",
		X"00",X"02",X"01",X"13",X"0E",X"00",X"00",X"02",X"00",X"D9",X"0E",X"00",X"00",X"02",X"00",X"B8",
		X"0E",X"00",X"00",X"02",X"00",X"92",X"16",X"00",X"00",X"02",X"00",X"B8",X"06",X"00",X"00",X"02",
		X"00",X"B8",X"40",X"FF",X"01",X"23",X"01",X"01",X"04",X"01",X"00",X"D9",X"01",X"00",X"C2",X"01",
		X"00",X"9A",X"01",X"00",X"74",X"01",X"00",X"61",X"01",X"00",X"39",X"01",X"00",X"61",X"01",X"00",
		X"92",X"01",X"00",X"C2",X"01",X"FF",X"00",X"78",X"02",X"00",X"6E",X"02",X"00",X"69",X"02",X"00",
		X"64",X"02",X"00",X"5F",X"02",X"00",X"5A",X"02",X"00",X"60",X"02",X"00",X"6B",X"02",X"00",X"77",
		X"02",X"00",X"82",X"02",X"00",X"8C",X"02",X"00",X"96",X"02",X"00",X"A0",X"02",X"00",X"AA",X"02",
		X"00",X"9F",X"02",X"00",X"95",X"02",X"00",X"85",X"02",X"00",X"78",X"02",X"00",X"82",X"02",X"00",
		X"8C",X"02",X"00",X"96",X"02",X"00",X"9F",X"02",X"00",X"B4",X"02",X"00",X"BE",X"02",X"00",X"D2",
		X"02",X"00",X"F0",X"02",X"01",X"04",X"02",X"01",X"18",X"02",X"01",X"36",X"02",X"01",X"54",X"02",
		X"01",X"7C",X"02",X"01",X"9A",X"02",X"01",X"D6",X"02",X"02",X"08",X"02",X"FF",X"00",X"89",X"0A",
		X"00",X"00",X"02",X"00",X"89",X"04",X"00",X"00",X"02",X"00",X"89",X"04",X"00",X"00",X"02",X"00",
		X"89",X"22",X"00",X"00",X"02",X"00",X"89",X"04",X"00",X"00",X"02",X"00",X"89",X"04",X"00",X"00",
		X"02",X"00",X"89",X"0A",X"00",X"00",X"02",X"00",X"B8",X"0A",X"00",X"00",X"02",X"00",X"89",X"0A",
		X"00",X"00",X"02",X"00",X"6D",X"0A",X"00",X"00",X"02",X"00",X"5C",X"10",X"00",X"00",X"02",X"00",
		X"7B",X"04",X"00",X"00",X"02",X"00",X"7B",X"30",X"FF",X"00",X"B8",X"0A",X"00",X"00",X"02",X"00",
		X"B8",X"04",X"00",X"00",X"02",X"00",X"B8",X"04",X"00",X"00",X"02",X"00",X"B8",X"22",X"00",X"00",
		X"02",X"00",X"B8",X"04",X"00",X"00",X"02",X"00",X"B8",X"04",X"00",X"00",X"02",X"00",X"B8",X"0A",
		X"00",X"00",X"02",X"00",X"D9",X"0A",X"00",X"00",X"02",X"00",X"B8",X"0A",X"00",X"00",X"02",X"00",
		X"89",X"0A",X"00",X"00",X"02",X"00",X"7B",X"10",X"00",X"00",X"02",X"00",X"92",X"04",X"00",X"00",
		X"02",X"00",X"92",X"30",X"FF",X"00",X"D9",X"0A",X"00",X"00",X"02",X"00",X"D9",X"04",X"00",X"00",
		X"02",X"00",X"D9",X"04",X"00",X"00",X"02",X"00",X"D9",X"22",X"00",X"00",X"02",X"00",X"D9",X"04",
		X"00",X"00",X"02",X"00",X"D9",X"04",X"00",X"00",X"02",X"00",X"D9",X"0A",X"00",X"00",X"02",X"01",
		X"13",X"0A",X"00",X"00",X"02",X"00",X"D9",X"0A",X"00",X"00",X"02",X"00",X"B8",X"0A",X"00",X"00",
		X"02",X"00",X"92",X"10",X"00",X"00",X"02",X"00",X"B8",X"04",X"00",X"00",X"02",X"00",X"B8",X"30",
		X"FF",X"CD",X"FD",X"54",X"CD",X"37",X"5A",X"CD",X"49",X"57",X"C3",X"68",X"56",X"3A",X"46",X"70",
		X"FE",X"00",X"CA",X"30",X"55",X"3A",X"5B",X"70",X"3D",X"32",X"5B",X"70",X"28",X"01",X"C9",X"3A",
		X"68",X"73",X"32",X"5B",X"70",X"3A",X"46",X"70",X"DD",X"2A",X"47",X"70",X"FE",X"04",X"CA",X"87",
		X"55",X"FE",X"03",X"CA",X"9C",X"55",X"FE",X"02",X"CA",X"B1",X"55",X"FE",X"01",X"CA",X"C6",X"55",
		X"3A",X"42",X"70",X"FE",X"01",X"C0",X"21",X"0A",X"73",X"ED",X"5B",X"3A",X"70",X"16",X"00",X"19",
		X"CD",X"4F",X"56",X"19",X"7E",X"FE",X"00",X"C0",X"3E",X"01",X"32",X"53",X"70",X"21",X"4B",X"5A",
		X"3A",X"3A",X"70",X"87",X"5F",X"16",X"00",X"19",X"56",X"23",X"5E",X"ED",X"53",X"47",X"70",X"3E",
		X"04",X"32",X"46",X"70",X"DD",X"2A",X"47",X"70",X"DD",X"36",X"01",X"BE",X"DD",X"36",X"02",X"BF",
		X"DD",X"36",X"21",X"C0",X"DD",X"36",X"22",X"C1",X"3A",X"CC",X"70",X"FE",X"01",X"C8",X"3E",X"06",
		X"32",X"0C",X"71",X"CD",X"8B",X"02",X"C9",X"DD",X"36",X"61",X"C4",X"DD",X"36",X"62",X"C5",X"DD",
		X"36",X"41",X"C2",X"DD",X"36",X"42",X"C3",X"21",X"46",X"70",X"35",X"C9",X"DD",X"36",X"20",X"BA",
		X"DD",X"36",X"40",X"BC",X"DD",X"36",X"21",X"BB",X"DD",X"36",X"41",X"BD",X"21",X"46",X"70",X"35",
		X"C9",X"DD",X"36",X"23",X"B7",X"DD",X"36",X"43",X"B9",X"DD",X"36",X"22",X"B6",X"DD",X"36",X"42",
		X"B8",X"21",X"46",X"70",X"35",X"C9",X"2A",X"62",X"73",X"CD",X"4F",X"56",X"19",X"ED",X"5B",X"3A",
		X"70",X"16",X"00",X"19",X"7E",X"F5",X"21",X"0A",X"73",X"ED",X"5B",X"3A",X"70",X"16",X"00",X"19",
		X"CD",X"4F",X"56",X"19",X"F1",X"77",X"DD",X"2A",X"47",X"70",X"DD",X"77",X"21",X"3C",X"DD",X"77",
		X"22",X"3C",X"DD",X"77",X"41",X"3C",X"DD",X"77",X"42",X"DD",X"36",X"00",X"00",X"DD",X"36",X"03",
		X"00",X"DD",X"36",X"60",X"00",X"DD",X"36",X"63",X"00",X"DD",X"36",X"01",X"F9",X"DD",X"36",X"02",
		X"FA",X"DD",X"36",X"20",X"B3",X"DD",X"36",X"40",X"B4",X"DD",X"36",X"61",X"F9",X"DD",X"36",X"62",
		X"FA",X"DD",X"36",X"23",X"B3",X"DD",X"36",X"43",X"B4",X"21",X"46",X"70",X"35",X"AF",X"32",X"53",
		X"70",X"3A",X"6F",X"70",X"FE",X"00",X"C2",X"43",X"56",X"21",X"AC",X"70",X"34",X"21",X"76",X"70",
		X"C3",X"4A",X"56",X"21",X"AD",X"70",X"34",X"21",X"7D",X"70",X"06",X"02",X"C3",X"F0",X"3E",X"3A",
		X"49",X"70",X"FE",X"00",X"C2",X"5B",X"56",X"11",X"00",X"00",X"C9",X"FE",X"01",X"C2",X"64",X"56",
		X"11",X"14",X"00",X"C9",X"11",X"28",X"00",X"C9",X"3A",X"24",X"74",X"FE",X"E9",X"CA",X"76",X"56",
		X"FE",X"08",X"CA",X"A1",X"56",X"C9",X"3E",X"09",X"32",X"24",X"74",X"21",X"49",X"70",X"3E",X"01",
		X"BE",X"20",X"03",X"32",X"C1",X"70",X"34",X"00",X"CD",X"4F",X"56",X"21",X"0A",X"73",X"19",X"0E",
		X"00",X"06",X"14",X"7E",X"FE",X"00",X"C2",X"B7",X"56",X"C3",X"13",X"57",X"23",X"0C",X"10",X"F3",
		X"C9",X"3E",X"E8",X"32",X"24",X"74",X"21",X"49",X"70",X"3E",X"02",X"BE",X"20",X"05",X"3E",X"01",
		X"32",X"C0",X"70",X"35",X"C3",X"87",X"56",X"C5",X"E5",X"F5",X"DD",X"21",X"4B",X"5A",X"79",X"87",
		X"5F",X"16",X"00",X"DD",X"19",X"DD",X"66",X"00",X"DD",X"6E",X"01",X"E5",X"DD",X"E1",X"F1",X"DD",
		X"77",X"21",X"3C",X"DD",X"77",X"22",X"3C",X"DD",X"77",X"41",X"3C",X"DD",X"77",X"42",X"DD",X"36",
		X"00",X"00",X"DD",X"36",X"03",X"00",X"DD",X"36",X"60",X"00",X"DD",X"36",X"63",X"00",X"DD",X"36",
		X"01",X"F9",X"DD",X"36",X"02",X"FA",X"DD",X"36",X"20",X"B3",X"DD",X"36",X"40",X"B4",X"DD",X"36",
		X"61",X"F9",X"DD",X"36",X"62",X"FA",X"DD",X"36",X"23",X"B3",X"DD",X"36",X"43",X"B4",X"E1",X"C1",
		X"C3",X"9C",X"56",X"C5",X"E5",X"DD",X"21",X"4B",X"5A",X"79",X"87",X"5F",X"16",X"00",X"DD",X"19",
		X"DD",X"66",X"00",X"DD",X"6E",X"01",X"E5",X"DD",X"E1",X"06",X"04",X"3E",X"A2",X"11",X"20",X"00",
		X"DD",X"77",X"00",X"3C",X"DD",X"77",X"01",X"3C",X"DD",X"77",X"02",X"3C",X"DD",X"77",X"03",X"3C",
		X"DD",X"19",X"10",X"EC",X"E1",X"C1",X"C3",X"9C",X"56",X"3A",X"39",X"70",X"FE",X"01",X"CA",X"5E",
		X"57",X"FE",X"02",X"CA",X"A2",X"57",X"FE",X"03",X"CA",X"E6",X"57",X"C3",X"21",X"58",X"3A",X"25",
		X"74",X"06",X"05",X"21",X"80",X"5A",X"BE",X"CA",X"5B",X"58",X"23",X"10",X"F9",X"FE",X"18",X"38",
		X"29",X"FE",X"1D",X"DA",X"D6",X"59",X"FE",X"48",X"38",X"20",X"FE",X"4D",X"DA",X"D6",X"59",X"FE",
		X"78",X"38",X"17",X"FE",X"7D",X"DA",X"D6",X"59",X"FE",X"A8",X"38",X"0E",X"FE",X"AD",X"DA",X"D6",
		X"59",X"FE",X"D8",X"38",X"05",X"FE",X"DD",X"DA",X"D6",X"59",X"AF",X"32",X"52",X"70",X"32",X"54",
		X"70",X"C9",X"3A",X"25",X"74",X"06",X"05",X"21",X"7B",X"5A",X"BE",X"CA",X"71",X"58",X"23",X"10",
		X"F9",X"FE",X"13",X"38",X"29",X"FE",X"19",X"DA",X"75",X"59",X"FE",X"43",X"38",X"20",X"FE",X"49",
		X"DA",X"75",X"59",X"FE",X"73",X"38",X"17",X"FE",X"79",X"DA",X"75",X"59",X"FE",X"A3",X"38",X"0E",
		X"FE",X"A9",X"DA",X"75",X"59",X"FE",X"D3",X"38",X"05",X"FE",X"D9",X"DA",X"75",X"59",X"AF",X"32",
		X"51",X"70",X"32",X"54",X"70",X"C9",X"3A",X"24",X"74",X"06",X"04",X"21",X"77",X"5A",X"BE",X"CA",
		X"87",X"58",X"23",X"10",X"F9",X"FE",X"2F",X"38",X"20",X"FE",X"35",X"DA",X"B3",X"58",X"FE",X"5F",
		X"38",X"17",X"FE",X"65",X"DA",X"B3",X"58",X"FE",X"8F",X"38",X"0E",X"FE",X"95",X"DA",X"B3",X"58",
		X"FE",X"BF",X"38",X"05",X"FE",X"C5",X"DA",X"B3",X"58",X"AF",X"32",X"4F",X"70",X"32",X"54",X"70",
		X"C9",X"3A",X"24",X"74",X"06",X"04",X"21",X"73",X"5A",X"BE",X"28",X"71",X"23",X"10",X"FA",X"FE",
		X"2B",X"38",X"20",X"FE",X"31",X"DA",X"14",X"59",X"FE",X"5F",X"38",X"17",X"FE",X"61",X"DA",X"14",
		X"59",X"FE",X"8B",X"38",X"0E",X"FE",X"91",X"DA",X"14",X"59",X"FE",X"BB",X"38",X"05",X"FE",X"C1",
		X"DA",X"14",X"59",X"AF",X"32",X"50",X"70",X"32",X"54",X"70",X"C9",X"CD",X"37",X"5A",X"21",X"8D",
		X"5A",X"06",X"04",X"BE",X"CA",X"6B",X"58",X"23",X"10",X"F9",X"C9",X"3E",X"01",X"32",X"51",X"70",
		X"C9",X"CD",X"37",X"5A",X"21",X"91",X"5A",X"06",X"04",X"BE",X"CA",X"81",X"58",X"23",X"10",X"F9",
		X"C9",X"3E",X"01",X"32",X"52",X"70",X"C9",X"CD",X"37",X"5A",X"21",X"89",X"5A",X"06",X"04",X"BE",
		X"CA",X"97",X"58",X"23",X"10",X"F9",X"C9",X"3E",X"01",X"32",X"50",X"70",X"C9",X"CD",X"37",X"5A",
		X"21",X"85",X"5A",X"06",X"04",X"BE",X"CA",X"AD",X"58",X"23",X"10",X"F9",X"C9",X"3E",X"01",X"32",
		X"4F",X"70",X"C9",X"CD",X"37",X"5A",X"FE",X"C6",X"C2",X"C7",X"58",X"AF",X"32",X"51",X"70",X"3E",
		X"01",X"32",X"50",X"70",X"C3",X"0E",X"59",X"FE",X"CE",X"C2",X"D8",X"58",X"AF",X"32",X"52",X"70",
		X"3E",X"01",X"32",X"50",X"70",X"C3",X"0E",X"59",X"FE",X"DA",X"C2",X"EC",X"58",X"AF",X"32",X"51",
		X"70",X"32",X"52",X"70",X"3E",X"01",X"32",X"50",X"70",X"C3",X"0E",X"59",X"FE",X"DE",X"C2",X"F8",
		X"58",X"AF",X"32",X"51",X"70",X"C3",X"0E",X"59",X"FE",X"E2",X"C2",X"04",X"59",X"AF",X"32",X"52",
		X"70",X"C3",X"0E",X"59",X"FE",X"E6",X"C0",X"AF",X"32",X"51",X"70",X"32",X"52",X"70",X"3E",X"01",
		X"32",X"54",X"70",X"C9",X"CD",X"37",X"5A",X"FE",X"CA",X"C2",X"28",X"59",X"AF",X"32",X"51",X"70",
		X"3E",X"01",X"32",X"4F",X"70",X"C3",X"6F",X"59",X"FE",X"D2",X"C2",X"39",X"59",X"AF",X"32",X"52",
		X"70",X"3E",X"01",X"32",X"4F",X"70",X"C3",X"6F",X"59",X"FE",X"D6",X"C2",X"4D",X"59",X"AF",X"32",
		X"51",X"70",X"32",X"52",X"70",X"3E",X"01",X"32",X"4F",X"70",X"C3",X"6F",X"59",X"FE",X"DE",X"C2",
		X"59",X"59",X"AF",X"32",X"51",X"70",X"C3",X"6F",X"59",X"FE",X"E2",X"C2",X"65",X"59",X"AF",X"32",
		X"52",X"70",X"C3",X"6F",X"59",X"FE",X"E6",X"C0",X"AF",X"32",X"51",X"70",X"32",X"52",X"70",X"3E",
		X"01",X"32",X"54",X"70",X"C9",X"CD",X"37",X"5A",X"FE",X"C6",X"C2",X"89",X"59",X"AF",X"32",X"4F",
		X"70",X"3E",X"01",X"32",X"52",X"70",X"C3",X"D0",X"59",X"FE",X"CA",X"C2",X"9A",X"59",X"AF",X"32",
		X"50",X"70",X"3E",X"01",X"32",X"52",X"70",X"C3",X"D0",X"59",X"FE",X"D6",X"C2",X"A6",X"59",X"AF",
		X"32",X"50",X"70",X"C3",X"D0",X"59",X"FE",X"DA",X"C2",X"B2",X"59",X"AF",X"32",X"4F",X"70",X"C3",
		X"D0",X"59",X"FE",X"DE",X"C2",X"C6",X"59",X"AF",X"32",X"4F",X"70",X"32",X"50",X"70",X"3E",X"01",
		X"32",X"52",X"70",X"C3",X"D0",X"59",X"FE",X"E6",X"C0",X"AF",X"32",X"4F",X"70",X"32",X"50",X"70",
		X"3E",X"01",X"32",X"54",X"70",X"C9",X"CD",X"37",X"5A",X"FE",X"CE",X"C2",X"EA",X"59",X"AF",X"32",
		X"4F",X"70",X"3E",X"01",X"32",X"51",X"70",X"C3",X"31",X"5A",X"FE",X"D2",X"C2",X"FB",X"59",X"AF",
		X"32",X"50",X"70",X"3E",X"01",X"32",X"51",X"70",X"C3",X"31",X"5A",X"FE",X"D6",X"C2",X"07",X"5A",
		X"AF",X"32",X"50",X"70",X"C3",X"31",X"5A",X"FE",X"DA",X"C2",X"13",X"5A",X"AF",X"32",X"4F",X"70",
		X"C3",X"31",X"5A",X"FE",X"E2",X"C2",X"27",X"5A",X"AF",X"32",X"4F",X"70",X"32",X"50",X"70",X"3E",
		X"01",X"32",X"51",X"70",X"C3",X"31",X"5A",X"FE",X"E6",X"C0",X"AF",X"32",X"50",X"70",X"32",X"4F",
		X"70",X"3E",X"01",X"32",X"54",X"70",X"C9",X"00",X"21",X"0A",X"73",X"ED",X"5B",X"3A",X"70",X"16",
		X"00",X"19",X"CD",X"4F",X"56",X"19",X"7E",X"32",X"4E",X"70",X"C9",X"88",X"A2",X"88",X"A8",X"88",
		X"AE",X"88",X"B4",X"88",X"BA",X"89",X"62",X"89",X"68",X"89",X"6E",X"89",X"74",X"89",X"7A",X"8A",
		X"22",X"8A",X"28",X"8A",X"2E",X"8A",X"34",X"8A",X"3A",X"8A",X"E2",X"8A",X"E8",X"8A",X"EE",X"8A",
		X"F4",X"8A",X"FA",X"24",X"54",X"84",X"B4",X"CC",X"9C",X"6C",X"3C",X"0C",X"3C",X"6C",X"9C",X"CC",
		X"24",X"54",X"84",X"B4",X"E4",X"C6",X"CE",X"DA",X"B2",X"CA",X"D2",X"D6",X"B2",X"C6",X"CA",X"DE",
		X"F9",X"CE",X"D2",X"E2",X"F9",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"08",X"FF",X"00",X"FF",X"08",X"FF",X"08",X"FF",X"00",X"FF",X"00",X"FF",X"08",X"FF",
		X"DF",X"08",X"FF",X"00",X"FF",X"08",X"FF",X"00",X"FF",X"00",X"FF",X"08",X"FF",X"08",X"FF",X"08",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"08",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"80",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"08",X"FF",X"00",X"FF",X"08",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"08",X"FF",X"00",X"FF",X"08",X"FF",X"00",X"FF",X"08",X"FF",X"00",X"FF",X"08",X"FF",X"00",X"FF",
		X"FF",X"08",X"7F",X"00",X"FF",X"08",X"FF",X"00",X"FF",X"00",X"FF",X"08",X"F7",X"08",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"08",X"FF",X"00",X"FF",X"08",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"08",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"10",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"04",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"80",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"08",X"FF",X"00",X"FF",X"80",X"FF",X"00",X"FF",X"00",
		X"08",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"08",X"FF",X"00",X"FF",X"08",X"FF",X"00",X"FF",X"08",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FB",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"08",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"08",X"FF",X"08",
		X"08",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"08",X"FF",X"00",X"FF",X"08",X"FF",X"00",X"EF",X"08",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"EF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"08",X"FF",
		X"FF",X"00",X"FF",X"00",X"F7",X"08",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"F7",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"08",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FB",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"08",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"08",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"08",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"7F",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"F7",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
