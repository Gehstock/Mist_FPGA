library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity travusa_spr_bit1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of travusa_spr_bit1 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"01",X"03",X"0F",X"3A",X"00",X"00",X"80",X"D6",X"81",X"23",X"49",X"81",
		X"12",X"02",X"00",X"00",X"01",X"00",X"00",X"00",X"81",X"03",X"06",X"01",X"07",X"9E",X"00",X"00",
		X"00",X"00",X"00",X"18",X"0C",X"36",X"C8",X"64",X"00",X"00",X"00",X"00",X"00",X"1E",X"34",X"B0",
		X"76",X"7F",X"DE",X"DC",X"98",X"00",X"00",X"00",X"00",X"04",X"1E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"0F",X"3F",X"00",X"00",X"00",X"80",X"D6",X"8F",X"23",X"49",
		X"1A",X"02",X"00",X"00",X"01",X"00",X"00",X"00",X"81",X"81",X"03",X"06",X"01",X"9F",X"07",X"00",
		X"00",X"00",X"00",X"00",X"1E",X"4D",X"96",X"C8",X"00",X"00",X"00",X"00",X"1E",X"E0",X"7C",X"B0",
		X"64",X"76",X"7F",X"DE",X"DC",X"18",X"00",X"00",X"20",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"06",X"01",X"4D",X"00",X"00",X"0F",X"00",X"0C",X"F3",X"80",X"80",
		X"1B",X"03",X"02",X"02",X"00",X"00",X"00",X"00",X"02",X"51",X"80",X"80",X"02",X"0D",X"00",X"00",
		X"00",X"00",X"E4",X"3E",X"3F",X"38",X"AC",X"68",X"00",X"00",X"00",X"BC",X"06",X"E0",X"1C",X"64",
		X"21",X"9D",X"C6",X"F4",X"F0",X"80",X"00",X"00",X"B2",X"00",X"04",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"02",X"36",X"03",X"01",X"21",X"00",X"00",X"1F",X"00",X"B1",X"EE",X"91",X"08",
		X"0E",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"02",X"20",X"C2",X"01",X"11",X"03",X"27",X"1E",
		X"00",X"08",X"CC",X"0F",X"FE",X"33",X"18",X"EC",X"00",X"00",X"20",X"BC",X"2E",X"C0",X"78",X"0C",
		X"79",X"03",X"9E",X"4E",X"78",X"60",X"00",X"00",X"E4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"07",X"0B",X"41",X"01",X"00",X"00",X"1F",X"00",X"B1",X"EE",X"91",X"08",
		X"0E",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"02",X"20",X"C2",X"01",X"11",X"03",X"27",X"1E",
		X"00",X"08",X"CC",X"0F",X"FE",X"33",X"18",X"EC",X"00",X"C0",X"00",X"BC",X"0E",X"C0",X"78",X"0C",
		X"79",X"03",X"9E",X"4E",X"78",X"60",X"00",X"00",X"E4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"01",X"01",X"01",X"06",X"06",X"04",X"98",X"A8",X"80",X"80",X"40",X"A3",X"C0",X"18",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"01",X"03",X"0F",X"3A",X"00",X"00",X"82",X"D5",X"80",X"28",X"52",X"98",
		X"12",X"02",X"00",X"00",X"01",X"00",X"00",X"00",X"90",X"00",X"01",X"00",X"05",X"9F",X"03",X"00",
		X"00",X"00",X"00",X"18",X"9C",X"C6",X"64",X"52",X"00",X"00",X"00",X"00",X"00",X"1E",X"34",X"B0",
		X"5B",X"DF",X"BE",X"BC",X"D8",X"80",X"00",X"00",X"20",X"04",X"1E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"01",X"03",X"0F",X"5A",X"00",X"00",X"82",X"D5",X"80",X"28",X"52",X"98",
		X"12",X"02",X"00",X"00",X"01",X"00",X"00",X"00",X"90",X"00",X"01",X"00",X"05",X"9F",X"03",X"00",
		X"00",X"00",X"00",X"18",X"9C",X"C6",X"64",X"52",X"00",X"00",X"00",X"00",X"00",X"1E",X"34",X"B0",
		X"5B",X"DF",X"BE",X"BC",X"D8",X"80",X"00",X"00",X"20",X"04",X"1E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"01",X"03",X"0F",X"3A",X"00",X"00",X"80",X"D7",X"80",X"21",X"44",X"90",
		X"12",X"02",X"00",X"00",X"01",X"00",X"00",X"00",X"80",X"01",X"03",X"00",X"07",X"9F",X"03",X"00",
		X"00",X"00",X"00",X"18",X"0C",X"9E",X"C8",X"A4",X"00",X"00",X"00",X"00",X"00",X"1E",X"34",X"B0",
		X"B6",X"BF",X"6E",X"5C",X"D8",X"80",X"00",X"00",X"20",X"04",X"1E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"01",X"03",X"07",X"4A",X"00",X"00",X"80",X"D7",X"80",X"20",X"44",X"90",
		X"0A",X"02",X"00",X"00",X"01",X"00",X"00",X"00",X"80",X"01",X"03",X"00",X"07",X"9F",X"03",X"00",
		X"00",X"00",X"00",X"18",X"0C",X"9E",X"C8",X"A4",X"00",X"00",X"00",X"00",X"00",X"1E",X"34",X"B0",
		X"B6",X"BF",X"6E",X"5C",X"D8",X"80",X"00",X"00",X"20",X"04",X"1E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"01",X"03",X"0F",X"1A",X"00",X"00",X"82",X"D5",X"80",X"28",X"52",X"98",
		X"12",X"02",X"00",X"00",X"01",X"00",X"00",X"00",X"90",X"00",X"01",X"00",X"05",X"9F",X"03",X"00",
		X"00",X"00",X"00",X"18",X"9C",X"C6",X"64",X"52",X"00",X"00",X"00",X"00",X"00",X"1E",X"34",X"B0",
		X"5B",X"DF",X"BE",X"BC",X"D8",X"80",X"00",X"00",X"20",X"04",X"1E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"03",X"00",X"00",X"00",X"CC",X"B3",X"80",X"28",X"52",
		X"0E",X"1A",X"3A",X"10",X"00",X"01",X"00",X"00",X"98",X"80",X"00",X"00",X"00",X"01",X"9F",X"07",
		X"00",X"00",X"00",X"18",X"1C",X"96",X"4A",X"64",X"00",X"00",X"00",X"00",X"00",X"1E",X"34",X"B0",
		X"52",X"5B",X"DF",X"B6",X"6E",X"CC",X"80",X"00",X"20",X"04",X"1E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"03",X"06",X"07",X"06",X"0F",X"2F",X"80",X"02",X"00",X"40",X"08",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"08",X"7F",X"1E",X"00",X"00",X"00",X"00",X"30",X"C0",X"60",X"70",
		X"87",X"E7",X"73",X"5F",X"5F",X"DF",X"BA",X"23",X"A4",X"08",X"10",X"40",X"00",X"00",X"00",X"00",
		X"2D",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"06",X"0C",X"52",X"40",X"C0",
		X"00",X"00",X"00",X"01",X"02",X"01",X"06",X"79",X"00",X"40",X"80",X"60",X"E0",X"C4",X"58",X"10",
		X"24",X"C2",X"0F",X"C7",X"AE",X"5D",X"5B",X"58",X"00",X"00",X"00",X"00",X"80",X"00",X"80",X"80",
		X"01",X"01",X"01",X"01",X"01",X"06",X"06",X"0C",X"88",X"A8",X"80",X"80",X"40",X"A3",X"C0",X"18",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"70",X"D0",X"60",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"01",X"03",X"07",X"4A",X"00",X"00",X"80",X"D6",X"81",X"23",X"49",X"81",
		X"0A",X"02",X"00",X"00",X"01",X"00",X"00",X"00",X"81",X"03",X"06",X"01",X"07",X"9E",X"00",X"00",
		X"00",X"00",X"00",X"18",X"0C",X"36",X"C8",X"64",X"00",X"00",X"00",X"00",X"00",X"1E",X"34",X"B0",
		X"76",X"7F",X"DE",X"DC",X"98",X"00",X"00",X"00",X"00",X"04",X"1E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"20",X"00",X"43",X"6B",X"35",X"08",X"BC",X"C0",X"00",X"40",X"80",X"00",X"00",X"80",X"60",
		X"F6",X"63",X"03",X"1F",X"0E",X"14",X"02",X"01",X"90",X"08",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"01",X"01",X"01",X"06",X"06",X"04",X"98",X"A8",X"80",X"80",X"40",X"A3",X"C0",X"18",
		X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"00",X"00",
		X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"10",X"00",X"08",X"08",X"00",X"00",X"00",X"08",X"08",
		X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"00",X"00",X"00",
		X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"00",X"04",X"04",X"00",X"00",X"00",X"08",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"00",X"60",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"40",X"5E",X"58",X"50",X"40",X"00",X"C0",X"3E",X"00",X"20",X"00",X"00",X"00",
		X"40",X"00",X"03",X"7F",X"7C",X"60",X"60",X"60",X"00",X"3C",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"20",X"33",X"7A",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",
		X"30",X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"30",X"CF",X"00",X"00",X"00",X"04",X"0E",X"00",X"00",X"80",X"3E",X"C0",X"00",X"00",X"00",
		X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"02",
		X"00",X"00",X"43",X"00",X"7F",X"40",X"40",X"40",X"00",X"C0",X"3E",X"00",X"7E",X"00",X"00",X"00",
		X"00",X"03",X"7C",X"20",X"00",X"00",X"00",X"20",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"7F",X"F8",X"CF",X"A2",X"B2",X"FA",X"00",X"00",X"C3",X"10",X"FF",X"0F",X"EF",X"EF",
		X"B2",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"EF",X"EF",X"EF",X"EE",X"EB",X"06",X"09",X"0A",
		X"00",X"30",X"CF",X"0E",X"FE",X"F8",X"E0",X"EE",X"00",X"00",X"80",X"3A",X"C0",X"00",X"00",X"00",
		X"E7",X"E7",X"E7",X"E7",X"E7",X"E7",X"A7",X"67",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",
		X"F2",X"F2",X"F2",X"F2",X"F3",X"F2",X"F3",X"B2",X"0A",X"09",X"06",X"0B",X"BE",X"EF",X"FF",X"EF",
		X"FB",X"B2",X"A3",X"CF",X"F8",X"7F",X"00",X"00",X"FF",X"4F",X"5F",X"FF",X"10",X"C3",X"00",X"00",
		X"67",X"A7",X"E7",X"E7",X"E7",X"E7",X"E7",X"E7",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"E0",X"F8",X"FE",X"0E",X"CF",X"30",X"00",X"00",X"00",X"00",X"C0",X"3A",X"80",X"00",X"00",
		X"20",X"00",X"00",X"00",X"20",X"7C",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",
		X"40",X"40",X"40",X"7F",X"00",X"43",X"00",X"00",X"00",X"00",X"00",X"7E",X"00",X"3E",X"C0",X"00",
		X"00",X"00",X"00",X"01",X"06",X"1B",X"36",X"27",X"00",X"00",X"00",X"00",X"06",X"0F",X"D0",X"00",
		X"5F",X"5F",X"4F",X"C0",X"80",X"80",X"80",X"80",X"FC",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"BF",X"00",X"1B",X"00",X"00",X"08",X"34",X"60",X"FB",X"01",X"DE",
		X"0E",X"00",X"86",X"C4",X"E0",X"C0",X"C0",X"C0",X"F0",X"00",X"86",X"0A",X"06",X"06",X"06",X"06",
		X"00",X"00",X"00",X"78",X"1C",X"3E",X"03",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"39",X"89",X"81",X"81",X"81",X"81",X"81",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"6F",X"77",X"FF",
		X"00",X"00",X"01",X"03",X"01",X"01",X"01",X"01",X"A0",X"E0",X"C0",X"C3",X"C7",X"DF",X"EF",X"9F",
		X"00",X"00",X"00",X"00",X"C0",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"26",X"FE",X"F2",X"FA",X"E2",X"E2",X"E2",X"F8",X"00",X"69",X"FD",X"FD",X"FD",X"FD",X"FD",
		X"00",X"00",X"00",X"00",X"F8",X"00",X"02",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0D",X"11",X"C9",X"A1",X"40",X"08",X"08",X"08",X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"38",X"20",X"20",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"21",X"2B",X"8E",X"38",X"70",X"01",X"07",X"5F",
		X"00",X"00",X"00",X"48",X"0F",X"79",X"04",X"0E",X"00",X"00",X"00",X"00",X"FC",X"F8",X"01",X"F8",
		X"8F",X"8C",X"C4",X"06",X"06",X"06",X"86",X"86",X"09",X"45",X"05",X"05",X"05",X"09",X"FB",X"E3",
		X"00",X"00",X"00",X"AA",X"00",X"8F",X"85",X"40",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"00",X"00",X"00",X"80",X"80",
		X"00",X"01",X"03",X"40",X"5E",X"58",X"50",X"40",X"00",X"00",X"3E",X"00",X"20",X"00",X"00",X"00",
		X"40",X"00",X"03",X"7F",X"7C",X"60",X"60",X"60",X"00",X"3C",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"20",X"33",X"7A",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",
		X"30",X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"CF",X"00",X"00",X"00",X"04",X"0E",X"00",X"00",X"80",X"3E",X"C4",X"00",X"00",X"00",
		X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"02",
		X"00",X"01",X"43",X"00",X"7F",X"40",X"40",X"40",X"00",X"00",X"3E",X"00",X"7E",X"00",X"00",X"00",
		X"00",X"03",X"7C",X"20",X"00",X"00",X"00",X"20",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"7F",X"F8",X"CD",X"A3",X"B3",X"F9",X"00",X"00",X"C3",X"10",X"B7",X"FF",X"FF",X"F7",
		X"B3",X"F9",X"FB",X"F9",X"FB",X"FA",X"FA",X"FA",X"FF",X"F7",X"FF",X"F6",X"FB",X"06",X"09",X"0A",
		X"00",X"40",X"CF",X"0E",X"FE",X"F8",X"E0",X"EE",X"00",X"00",X"80",X"3A",X"C0",X"00",X"00",X"00",
		X"E7",X"E7",X"E7",X"E7",X"E7",X"E7",X"E7",X"67",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",
		X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"FA",X"B2",X"0A",X"09",X"06",X"0B",X"0E",X"0F",X"0F",X"0F",
		X"FA",X"B2",X"A2",X"CF",X"F8",X"7F",X"00",X"00",X"8F",X"CF",X"0F",X"FF",X"10",X"C3",X"00",X"00",
		X"67",X"E7",X"E7",X"E7",X"E7",X"E7",X"E7",X"E7",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"E0",X"F8",X"FE",X"0E",X"CF",X"40",X"00",X"00",X"00",X"00",X"C0",X"3A",X"80",X"00",X"00",
		X"20",X"00",X"00",X"00",X"20",X"7C",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",
		X"40",X"40",X"40",X"7F",X"00",X"43",X"01",X"00",X"00",X"00",X"00",X"7E",X"00",X"3E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"06",X"1B",X"36",X"27",X"00",X"00",X"00",X"C0",X"06",X"0F",X"D0",X"00",
		X"5F",X"5F",X"4F",X"C0",X"80",X"80",X"80",X"80",X"FC",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"BF",X"00",X"1B",X"00",X"00",X"06",X"34",X"60",X"FB",X"01",X"DE",
		X"0E",X"00",X"86",X"C4",X"E0",X"C0",X"C0",X"C0",X"F0",X"00",X"86",X"0A",X"06",X"06",X"06",X"06",
		X"00",X"00",X"00",X"78",X"1C",X"3E",X"03",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"39",X"89",X"81",X"81",X"81",X"81",X"81",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"6F",X"77",X"FF",
		X"00",X"00",X"01",X"03",X"01",X"01",X"01",X"01",X"A0",X"E0",X"C0",X"C3",X"C7",X"DF",X"EF",X"9F",
		X"00",X"00",X"00",X"00",X"C0",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"26",X"FE",X"F2",X"FA",X"E2",X"E2",X"E2",X"F8",X"00",X"69",X"FD",X"FD",X"FD",X"FD",X"FD",
		X"00",X"00",X"00",X"00",X"F8",X"00",X"02",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0D",X"11",X"C9",X"A1",X"40",X"08",X"08",X"08",X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"38",X"0C",X"14",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"10",X"1B",X"8E",X"18",X"58",X"01",X"07",X"5F",
		X"00",X"00",X"00",X"A8",X"0F",X"79",X"04",X"0E",X"00",X"00",X"00",X"01",X"FC",X"F8",X"01",X"78",
		X"8F",X"8C",X"C4",X"06",X"06",X"06",X"86",X"86",X"09",X"45",X"05",X"05",X"05",X"09",X"FB",X"E3",
		X"00",X"00",X"00",X"75",X"00",X"8F",X"85",X"40",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"00",X"00",X"00",X"80",X"80",
		X"00",X"08",X"1A",X"08",X"00",X"14",X"16",X"05",X"00",X"30",X"FF",X"00",X"84",X"00",X"3F",X"98",
		X"10",X"10",X"08",X"08",X"08",X"08",X"18",X"18",X"FB",X"BC",X"98",X"F8",X"B8",X"98",X"F8",X"F8",
		X"18",X"18",X"4F",X"1F",X"1F",X"5F",X"9E",X"1C",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",
		X"9C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1E",X"3E",X"7F",X"7F",X"7F",X"7F",X"3F",X"07",X"00",
		X"18",X"18",X"00",X"08",X"00",X"00",X"10",X"10",X"F8",X"F8",X"98",X"18",X"E8",X"18",X"18",X"08",
		X"01",X"12",X"10",X"00",X"08",X"1A",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"30",X"00",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1C",X"1C",X"1C",X"00",X"F0",X"FE",X"FF",X"FF",X"7F",X"7F",X"3E",
		X"1C",X"1E",X"5F",X"1F",X"1F",X"4F",X"18",X"18",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",
		X"C0",X"C0",X"FF",X"FF",X"FF",X"7F",X"3F",X"1F",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"1F",X"1F",X"1F",X"FF",X"FF",X"FF",X"FE",X"7E",X"FF",X"FF",X"FF",X"E0",X"80",X"00",X"0E",X"1E",
		X"C5",X"C0",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"FE",X"00",X"FF",X"FF",X"FF",X"31",X"31",X"31",
		X"FE",X"FE",X"FF",X"FF",X"7E",X"3E",X"1E",X"1E",X"31",X"31",X"F1",X"F1",X"31",X"31",X"30",X"30",
		X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0E",X"0E",X"3C",X"78",X"70",X"60",X"41",X"03",X"07",X"0E",
		X"1F",X"1F",X"3F",X"FF",X"FF",X"FF",X"C0",X"C0",X"00",X"80",X"E0",X"FF",X"FF",X"FF",X"00",X"00",
		X"1E",X"36",X"66",X"C6",X"C6",X"86",X"0E",X"0E",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",
		X"1E",X"3E",X"FE",X"FF",X"FF",X"FF",X"C0",X"C5",X"30",X"30",X"31",X"FF",X"FF",X"FF",X"00",X"FE",
		X"DD",X"C0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"5E",X"00",X"FF",X"FF",X"FF",X"F1",X"F1",X"F1",
		X"FF",X"FF",X"FF",X"81",X"00",X"00",X"00",X"00",X"F1",X"F1",X"F1",X"F1",X"F1",X"71",X"71",X"31",
		X"DF",X"C0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"D6",X"06",X"F8",X"FA",X"FA",X"18",X"1A",X"1A",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"18",X"1A",X"1A",X"18",X"1A",X"1A",X"18",X"1A",
		X"7C",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FC",X"31",X"31",X"31",X"31",X"31",X"30",X"38",X"38",
		X"00",X"00",X"00",X"FF",X"FF",X"FF",X"C0",X"DD",X"3C",X"7E",X"FF",X"FF",X"FF",X"FF",X"00",X"5E",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"1A",X"18",X"1A",X"1A",X"18",X"1A",X"1A",X"18",
		X"00",X"00",X"80",X"FF",X"FF",X"FF",X"C0",X"DF",X"1A",X"1A",X"18",X"FA",X"FA",X"F8",X"06",X"D6",
		X"00",X"08",X"1A",X"08",X"00",X"10",X"14",X"03",X"00",X"80",X"FF",X"00",X"84",X"00",X"7F",X"D8",
		X"1C",X"1C",X"08",X"08",X"08",X"08",X"18",X"18",X"FB",X"FC",X"D8",X"F8",X"F8",X"D8",X"F8",X"F8",
		X"18",X"18",X"00",X"08",X"00",X"00",X"10",X"11",X"F8",X"F8",X"D8",X"58",X"E8",X"58",X"58",X"08",
		X"02",X"10",X"10",X"00",X"08",X"1A",X"08",X"00",X"40",X"40",X"00",X"00",X"00",X"FF",X"80",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"0F",X"00",X"00",X"00",X"8E",X"D1",X"80",X"20",X"04",
		X"3A",X"12",X"02",X"00",X"00",X"01",X"00",X"00",X"80",X"90",X"01",X"03",X"01",X"07",X"8F",X"00",
		X"00",X"00",X"00",X"2C",X"77",X"19",X"88",X"C8",X"00",X"00",X"00",X"00",X"3E",X"F8",X"3C",X"B0",
		X"A5",X"BF",X"BE",X"6C",X"46",X"9C",X"18",X"00",X"20",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"5C",X"23",
		X"02",X"05",X"06",X"0D",X"5D",X"12",X"01",X"00",X"00",X"04",X"00",X"10",X"01",X"03",X"0F",X"9F",
		X"00",X"00",X"00",X"03",X"37",X"F8",X"40",X"8C",X"00",X"00",X"38",X"D0",X"78",X"30",X"80",X"0C",
		X"47",X"F6",X"B6",X"BE",X"A2",X"64",X"C6",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"0C",
		X"00",X"00",X"00",X"01",X"07",X"07",X"26",X"1E",X"30",X"1F",X"1C",X"11",X"80",X"00",X"04",X"80",
		X"00",X"00",X"00",X"03",X"2E",X"E1",X"CE",X"F1",X"00",X"20",X"F0",X"90",X"20",X"E0",X"C8",X"10",
		X"D0",X"4E",X"9F",X"8D",X"5B",X"F7",X"B2",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"34",X"02",X"00",X"01",X"00",X"00",X"00",X"00",X"31",X"03",X"00",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"0C",
		X"00",X"00",X"00",X"01",X"03",X"0F",X"06",X"5E",X"30",X"1F",X"1C",X"11",X"80",X"00",X"04",X"80",
		X"14",X"02",X"00",X"01",X"00",X"00",X"00",X"00",X"31",X"03",X"00",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0C",X"C0",X"D8",X"0C",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"07",X"2E",X"02",X"04",X"00",X"08",X"08",
		X"00",X"00",X"00",X"3F",X"1F",X"80",X"9D",X"3A",X"00",X"00",X"00",X"C9",X"F3",X"00",X"3C",X"DF",
		X"54",X"60",X"80",X"40",X"21",X"12",X"0F",X"7F",X"3B",X"3C",X"23",X"A0",X"E8",X"C0",X"C0",X"00",
		X"00",X"40",X"40",X"40",X"8C",X"FC",X"F8",X"9C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"8C",X"C4",X"60",X"B0",X"5C",X"20",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"20",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"20",X"00",X"40",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"03",X"36",X"30",X"02",X"02",X"02",X"20",X"F0",X"A8",X"20",X"27",X"00",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"12",X"0A",X"0B",X"0A",X"19",X"1A",X"19",X"1A",X"E0",X"E0",X"F8",X"EC",X"06",X"0E",X"03",X"07",
		X"19",X"1A",X"1B",X"1A",X"11",X"00",X"00",X"00",X"07",X"83",X"43",X"85",X"D9",X"61",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"00",X"00",X"00",X"00",X"00",X"84",X"8E",X"8C",
		X"03",X"36",X"34",X"0E",X"0B",X"1B",X"09",X"03",X"18",X"34",X"68",X"D0",X"D0",X"A0",X"A0",X"A0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"65",X"43",X"01",X"02",X"15",X"00",X"01",
		X"02",X"0C",X"3A",X"74",X"E8",X"14",X"28",X"30",X"3E",X"CF",X"70",X"7F",X"78",X"60",X"28",X"20",
		X"60",X"70",X"0C",X"81",X"83",X"06",X"0C",X"80",X"E0",X"70",X"E0",X"E0",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"06",X"0F",X"2E",X"70",X"00",X"00",X"20",X"60",X"00",X"F8",X"7C",X"00",
		X"8F",X"33",X"1C",X"1F",X"1E",X"18",X"0A",X"08",X"80",X"F2",X"3F",X"C2",X"00",X"00",X"00",X"00",
		X"80",X"8A",X"04",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"33",X"2F",X"1C",X"70",X"00",X"00",X"40",X"C0",X"C0",X"0E",X"1E",X"78",
		X"23",X"07",X"8E",X"A9",X"A7",X"6E",X"5C",X"5C",X"E0",X"80",X"00",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"02",X"02",X"05",X"1D",X"1D",X"8F",X"1E",X"39",X"A6",X"9C",X"B8",X"70",X"70",
		X"3A",X"3A",X"74",X"76",X"E8",X"AC",X"18",X"0C",X"38",X"0C",X"14",X"0C",X"04",X"1C",X"1C",X"19",
		X"83",X"03",X"07",X"07",X"06",X"C6",X"2C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"08",X"00",X"00",X"80",X"01",X"C0",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1D",X"3A",X"2B",X"06",X"03",X"01",X"20",X"40",
		X"06",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"7F",X"47",X"44",X"48",X"30",X"00",X"00",
		X"6A",X"AA",X"98",X"94",X"50",X"52",X"35",X"3A",X"00",X"F8",X"9C",X"74",X"0E",X"07",X"03",X"83",
		X"19",X"1D",X"1D",X"0E",X"0C",X"04",X"00",X"00",X"D4",X"B8",X"F0",X"00",X"1E",X"0D",X"0C",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"20",X"00",X"00",X"70",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"38",X"A0",X"80",X"11",X"10",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"06",X"16",X"16",X"16",X"04",X"00",X"E0",X"60",X"C0",X"C0",X"C0",X"C8",X"C0",
		X"04",X"34",X"24",X"04",X"05",X"02",X"02",X"02",X"D0",X"C0",X"E0",X"EA",X"A8",X"AB",X"63",X"51",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"10",X"18",X"08",X"0C",X"84",X"D6",
		X"00",X"00",X"03",X"03",X"00",X"00",X"00",X"00",X"C6",X"67",X"23",X"11",X"18",X"28",X"27",X"01",
		X"40",X"64",X"6A",X"75",X"37",X"1B",X"8A",X"88",X"00",X"00",X"AC",X"7F",X"C7",X"01",X"01",X"01",
		X"70",X"1A",X"07",X"03",X"01",X"00",X"00",X"00",X"A2",X"5A",X"3E",X"D8",X"E0",X"F0",X"20",X"10",
		X"00",X"30",X"08",X"04",X"80",X"C4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"0A",X"22",X"70",X"68",X"C8",X"C4",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"18",X"0B",X"03",X"30",X"20",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"0C",X"0A",X"75",X"34",X"0A",X"0C",X"00",X"00",X"40",X"03",X"0B",X"0B",X"03",X"40",X"80",X"00",
		X"0F",X"18",X"10",X"13",X"10",X"18",X"10",X"13",X"F8",X"0C",X"04",X"F4",X"04",X"0C",X"04",X"F4",
		X"10",X"78",X"40",X"40",X"60",X"39",X"0E",X"03",X"07",X"01",X"01",X"03",X"E7",X"04",X"0C",X"F8",
		X"0F",X"18",X"10",X"13",X"10",X"18",X"10",X"13",X"F8",X"0C",X"04",X"F4",X"04",X"0C",X"04",X"F4",
		X"10",X"68",X"4F",X"4E",X"42",X"40",X"40",X"7F",X"04",X"03",X"01",X"01",X"F1",X"99",X"8B",X"8E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"00",X"00",X"00",X"00",X"04",X"00",X"09",X"08",X"42",X"80",X"0F",X"71",X"9C",X"4D",X"D4",
		X"03",X"07",X"0B",X"00",X"02",X"00",X"00",X"00",X"8F",X"5D",X"FC",X"7A",X"A8",X"10",X"40",X"10",
		X"00",X"A3",X"4C",X"36",X"BC",X"00",X"C4",X"EA",X"C0",X"C0",X"10",X"A8",X"85",X"A0",X"55",X"A8",
		X"B5",X"0E",X"15",X"19",X"1A",X"00",X"10",X"00",X"49",X"08",X"60",X"8A",X"00",X"00",X"00",X"20",
		X"04",X"00",X"00",X"00",X"02",X"04",X"00",X"43",X"08",X"40",X"98",X"2C",X"00",X"53",X"EE",X"D0",
		X"0E",X"18",X"0C",X"02",X"01",X"00",X"00",X"08",X"A2",X"67",X"14",X"C2",X"F0",X"18",X"20",X"10",
		X"00",X"03",X"24",X"0E",X"B8",X"83",X"1E",X"28",X"20",X"C8",X"10",X"08",X"D5",X"6D",X"16",X"36",
		X"E1",X"0F",X"15",X"1E",X"19",X"1A",X"04",X"20",X"C0",X"5C",X"C3",X"60",X"0A",X"00",X"80",X"00",
		X"02",X"00",X"00",X"00",X"30",X"37",X"53",X"7E",X"08",X"00",X"88",X"40",X"E4",X"C3",X"13",X"AB",
		X"F4",X"78",X"7E",X"6A",X"70",X"70",X"61",X"61",X"7E",X"F4",X"EB",X"45",X"2B",X"7E",X"E9",X"E7",
		X"08",X"01",X"00",X"81",X"1A",X"01",X"4F",X"D4",X"00",X"00",X"00",X"40",X"30",X"5E",X"62",X"DC",
		X"91",X"36",X"42",X"84",X"1D",X"FB",X"E2",X"88",X"92",X"82",X"2C",X"40",X"90",X"20",X"CE",X"DC",
		X"63",X"62",X"73",X"70",X"65",X"71",X"70",X"F4",X"73",X"21",X"D8",X"53",X"25",X"01",X"DC",X"36",
		X"74",X"50",X"37",X"30",X"00",X"00",X"00",X"00",X"10",X"09",X"87",X"C4",X"41",X"80",X"00",X"08",
		X"C9",X"7A",X"D3",X"EC",X"90",X"7A",X"BE",X"F7",X"D4",X"E6",X"51",X"04",X"01",X"0D",X"1C",X"02",
		X"70",X"4D",X"11",X"00",X"01",X"00",X"01",X"00",X"91",X"68",X"28",X"16",X"40",X"00",X"00",X"00",
		X"02",X"00",X"00",X"00",X"31",X"37",X"52",X"7C",X"08",X"00",X"98",X"61",X"E5",X"5F",X"BD",X"61",
		X"F4",X"78",X"7D",X"68",X"70",X"74",X"61",X"63",X"C2",X"80",X"49",X"47",X"27",X"3C",X"30",X"42",
		X"08",X"01",X"04",X"89",X"D3",X"20",X"5A",X"64",X"00",X"00",X"00",X"40",X"13",X"28",X"70",X"EC",
		X"A1",X"C2",X"42",X"85",X"1A",X"F3",X"E4",X"88",X"C0",X"00",X"F0",X"90",X"28",X"90",X"2E",X"1C",
		X"6E",X"66",X"70",X"72",X"6B",X"7D",X"78",X"F6",X"52",X"21",X"10",X"43",X"CC",X"2D",X"FF",X"56",
		X"75",X"50",X"37",X"30",X"00",X"00",X"00",X"00",X"1B",X"A9",X"A4",X"B6",X"59",X"95",X"00",X"00",
		X"07",X"02",X"60",X"40",X"92",X"7F",X"2E",X"87",X"DC",X"EE",X"75",X"1E",X"00",X"45",X"1E",X"40",
		X"11",X"4C",X"24",X"1E",X"01",X"00",X"01",X"00",X"B0",X"A8",X"20",X"32",X"C0",X"40",X"02",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"1E",X"00",X"00",X"86",X"B3",X"01",X"00",X"8C",X"18",
		X"0E",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"93",X"0F",X"01",X"80",X"98",X"00",X"00",
		X"00",X"00",X"00",X"00",X"90",X"59",X"B2",X"95",X"00",X"00",X"00",X"00",X"14",X"00",X"64",X"B0",
		X"B7",X"A2",X"4D",X"9A",X"10",X"00",X"00",X"00",X"20",X"04",X"00",X"14",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"03",X"0C",X"3E",X"00",X"00",X"00",X"80",X"BE",X"0F",X"00",X"8C",
		X"1A",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"18",X"10",X"93",X"0F",X"81",X"98",X"00",X"00",
		X"00",X"00",X"00",X"00",X"22",X"90",X"40",X"B6",X"00",X"00",X"00",X"00",X"14",X"C0",X"64",X"B0",
		X"95",X"B7",X"A6",X"4C",X"88",X"18",X"10",X"00",X"20",X"04",X"14",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"02",X"4D",X"00",X"00",X"00",X"00",X"00",X"80",X"9E",X"4F",
		X"18",X"02",X"02",X"02",X"00",X"00",X"00",X"00",X"10",X"8C",X"08",X"90",X"11",X"97",X"00",X"00",
		X"00",X"00",X"08",X"00",X"04",X"23",X"10",X"82",X"00",X"00",X"00",X"00",X"14",X"80",X"F4",X"70",
		X"45",X"B7",X"96",X"B4",X"E4",X"88",X"00",X"00",X"B0",X"04",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"42",X"01",X"0E",X"00",X"00",X"00",X"00",X"00",X"82",X"C6",X"09",
		X"00",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"0F",X"9E",X"10",X"8C",X"38",X"10",X"11",X"0B",
		X"00",X"00",X"05",X"18",X"0C",X"43",X"20",X"02",X"00",X"00",X"80",X"60",X"14",X"00",X"C4",X"34",
		X"85",X"77",X"96",X"B0",X"B0",X"E0",X"80",X"00",X"88",X"38",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"02",X"21",X"0E",X"00",X"00",X"00",X"00",X"00",X"82",X"C6",X"09",
		X"00",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"0F",X"9E",X"10",X"8C",X"38",X"10",X"11",X"0B",
		X"00",X"00",X"05",X"18",X"0C",X"43",X"20",X"02",X"00",X"00",X"80",X"60",X"14",X"00",X"C4",X"34",
		X"85",X"77",X"96",X"B0",X"B0",X"E0",X"80",X"00",X"88",X"38",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"2E",X"00",X"00",X"86",X"B3",X"01",X"00",X"8C",X"18",
		X"0E",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"93",X"0F",X"01",X"80",X"98",X"00",X"00",
		X"00",X"00",X"00",X"00",X"90",X"59",X"B2",X"95",X"00",X"00",X"00",X"00",X"14",X"00",X"64",X"70",
		X"B7",X"A2",X"4D",X"9A",X"10",X"00",X"00",X"00",X"20",X"04",X"00",X"14",X"00",X"00",X"00",X"00",
		X"07",X"0C",X"18",X"10",X"13",X"10",X"18",X"10",X"FC",X"06",X"02",X"02",X"F2",X"06",X"02",X"02",
		X"13",X"10",X"60",X"40",X"40",X"40",X"73",X"1E",X"F2",X"07",X"01",X"01",X"01",X"03",X"FE",X"00",
		X"3F",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",
		X"00",X"00",X"18",X"20",X"00",X"40",X"00",X"00",X"30",X"38",X"18",X"1C",X"1D",X"0D",X"0E",X"0E",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"30",X"1F",X"1F",X"0E",X"0E",X"1C",X"1C",X"3C",X"78",X"F8",X"F0",
		X"27",X"20",X"20",X"20",X"20",X"20",X"3F",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"C0",X"C0",X"40",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",
		X"0F",X"18",X"10",X"13",X"10",X"18",X"10",X"11",X"F4",X"02",X"02",X"F2",X"06",X"02",X"02",X"F6",
		X"30",X"60",X"40",X"40",X"5E",X"52",X"53",X"71",X"02",X"02",X"72",X"02",X"02",X"02",X"06",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"80",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"10",X"DC",X"DC",
		X"00",X"80",X"FF",X"FF",X"00",X"00",X"C0",X"C0",X"00",X"10",X"DC",X"DC",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"06",X"06",X"06",
		X"00",X"00",X"00",X"7F",X"7F",X"7F",X"00",X"00",X"06",X"06",X"06",X"FE",X"FE",X"FE",X"00",X"00",
		X"FF",X"DF",X"C0",X"C0",X"00",X"80",X"FF",X"F8",X"FC",X"FC",X"00",X"00",X"00",X"00",X"FC",X"E0",
		X"03",X"8E",X"FF",X"FF",X"00",X"80",X"FF",X"FF",X"80",X"00",X"FC",X"FC",X"00",X"00",X"FC",X"FC",
		X"00",X"00",X"00",X"00",X"01",X"0F",X"7F",X"7D",X"00",X"00",X"06",X"3E",X"FE",X"FE",X"FC",X"E0",
		X"7C",X"7F",X"0F",X"01",X"00",X"00",X"00",X"00",X"E0",X"E0",X"F8",X"FE",X"3E",X"06",X"00",X"00",
		X"00",X"00",X"BF",X"C0",X"C0",X"C0",X"FF",X"7F",X"00",X"00",X"F8",X"04",X"04",X"04",X"F8",X"F8",
		X"00",X"00",X"BE",X"C1",X"C1",X"C1",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"FC",
		X"00",X"40",X"7F",X"7F",X"7F",X"6F",X"60",X"60",X"00",X"00",X"FC",X"FE",X"FE",X"FE",X"0E",X"0E",
		X"60",X"60",X"60",X"7F",X"7F",X"3F",X"00",X"00",X"0E",X"0E",X"0E",X"FE",X"FE",X"FE",X"02",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"C0",X"F0",X"3C",X"1F",X"80",X"FF",X"FF",X"00",X"0C",X"30",X"C0",X"00",X"80",X"FC",X"FC",
		X"00",X"40",X"79",X"79",X"79",X"79",X"61",X"61",X"00",X"00",X"FC",X"FE",X"FE",X"FE",X"8E",X"8E",
		X"60",X"60",X"60",X"7F",X"7F",X"3F",X"00",X"00",X"0E",X"0E",X"06",X"FE",X"FE",X"FE",X"02",X"00",
		X"00",X"00",X"B0",X"C0",X"C0",X"C0",X"FF",X"7F",X"00",X"20",X"38",X"3C",X"0C",X"04",X"F8",X"F8",
		X"00",X"80",X"C0",X"C1",X"C1",X"C1",X"FF",X"FF",X"00",X"00",X"04",X"04",X"04",X"04",X"FC",X"FC",
		X"00",X"80",X"FF",X"FF",X"03",X"81",X"FF",X"FF",X"00",X"00",X"FC",X"00",X"00",X"00",X"FC",X"FC",
		X"00",X"00",X"B0",X"C0",X"C0",X"C0",X"FF",X"7F",X"00",X"20",X"38",X"3C",X"0C",X"04",X"F8",X"F8",
		X"00",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"21",X"18",X"0C",
		X"00",X"00",X"03",X"07",X"07",X"03",X"00",X"00",X"0C",X"04",X"C6",X"E6",X"4C",X"E9",X"00",X"00",
		X"00",X"00",X"40",X"00",X"80",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"8F",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"10",X"40",X"7C",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
		X"03",X"00",X"03",X"07",X"07",X"03",X"00",X"00",X"F0",X"38",X"DC",X"EC",X"48",X"E9",X"00",X"00",
		X"00",X"00",X"00",X"00",X"40",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"8F",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
		X"00",X"08",X"02",X"0F",X"0F",X"13",X"A0",X"40",X"00",X"08",X"80",X"E0",X"30",X"D9",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"0F",X"07",X"03",X"01",X"03",X"01",X"08",X"80",X"E0",X"70",X"F9",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"80",X"8F",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0B",X"0F",X"07",X"03",X"01",X"00",X"01",X"08",X"80",X"E0",X"70",X"F9",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"06",X"0F",X"0F",X"1B",X"10",X"32",X"24",X"08",X"80",X"E0",X"B0",X"D9",X"00",X"80",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"80",X"8C",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"00",X"00",X"01",
		X"03",X"07",X"07",X"03",X"00",X"00",X"00",X"00",X"CB",X"E7",X"4E",X"EC",X"E9",X"00",X"00",X"00",
		X"08",X"18",X"30",X"60",X"40",X"40",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"87",X"80",X"8C",X"0F",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"07",X"07",X"03",X"00",X"00",X"00",X"00",X"C9",X"E3",X"4F",X"EE",X"E9",X"00",X"00",X"00",
		X"00",X"00",X"0C",X"0C",X"10",X"20",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"87",X"80",X"8C",X"0F",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"17",X"1F",X"1F",X"0B",X"0F",X"0D",X"06",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"7F",X"7F",X"71",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"07",X"0F",X"1E",X"1D",X"1F",
		X"05",X"06",X"02",X"03",X"03",X"01",X"01",X"00",X"E0",X"E0",X"F0",X"7F",X"3F",X"DF",X"E0",X"7F",
		X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"F9",X"FF",X"FF",X"CF",X"F0",X"1F",X"00",X"00",
		X"73",X"30",X"30",X"39",X"39",X"19",X"19",X"1F",X"FF",X"1F",X"00",X"E0",X"FF",X"C3",X"C0",X"C0",
		X"1F",X"00",X"03",X"07",X"07",X"07",X"06",X"04",X"C0",X"00",X"FF",X"FF",X"FF",X"40",X"FF",X"C1",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"FE",X"FE",X"EE",X"E7",X"67",X"67",X"73",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"FF",
		X"00",X"80",X"80",X"C0",X"C0",X"E0",X"F0",X"78",X"7F",X"5E",X"7C",X"7E",X"2E",X"3F",X"3F",X"17",
		X"BC",X"DF",X"EF",X"73",X"3C",X"1F",X"07",X"00",X"1F",X"1F",X"FE",X"FF",X"7D",X"83",X"FF",X"FE",
		X"1B",X"0B",X"0D",X"0D",X"FD",X"FE",X"FE",X"06",X"8F",X"80",X"C0",X"C0",X"C0",X"F0",X"FF",X"FF",
		X"FC",X"0F",X"00",X"E0",X"E0",X"60",X"E0",X"E0",X"1F",X"F0",X"3F",X"00",X"0F",X"3F",X"3C",X"7B",
		X"07",X"00",X"00",X"80",X"FE",X"FF",X"FF",X"83",X"99",X"DD",X"CC",X"6E",X"7E",X"F6",X"F6",X"F6",
		X"FE",X"C7",X"FF",X"FF",X"7F",X"C1",X"FA",X"1B",X"0E",X"FC",X"00",X"FC",X"FF",X"FF",X"07",X"FC",
		X"FC",X"FE",X"FE",X"07",X"07",X"FF",X"1F",X"00",X"FE",X"FF",X"7F",X"7F",X"3F",X"BF",X"9F",X"1F",
		X"00",X"00",X"80",X"FE",X"FF",X"FF",X"83",X"FE",X"1F",X"0F",X"0F",X"07",X"E7",X"F3",X"FB",X"3B",
		X"40",X"60",X"30",X"38",X"1C",X"1E",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"07",X"07",X"07",X"03",X"03",X"01",X"01",X"00",X"80",X"C0",X"E0",X"F0",X"F8",X"F8",X"FC",X"FE",
		X"EF",X"F7",X"3B",X"1D",X"0E",X"07",X"03",X"01",X"87",X"C7",X"E7",X"F3",X"F3",X"79",X"FD",X"BC",
		X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"FE",X"DE",X"7E",X"6E",X"3E",X"3C",X"10",X"00",
		X"F6",X"03",X"03",X"01",X"01",X"00",X"C0",X"FE",X"6F",X"6F",X"EF",X"EF",X"EF",X"EF",X"EF",X"6C",
		X"FF",X"7F",X"C3",X"FF",X"F0",X"FC",X"7E",X"9F",X"6C",X"2D",X"A1",X"A1",X"3F",X"1F",X"0F",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"7F",X"77",X"37",X"23",X"F3",X"F3",X"F7",X"E7",X"E7",X"EF",X"EF",X"EE",
		X"23",X"03",X"01",X"01",X"C1",X"E0",X"E0",X"74",X"EE",X"EC",X"EC",X"ED",X"ED",X"ED",X"EC",X"EC",
		X"00",X"00",X"80",X"80",X"C0",X"C0",X"E0",X"F0",X"2E",X"2C",X"2C",X"21",X"21",X"3F",X"00",X"00",
		X"F0",X"F8",X"F8",X"FD",X"FD",X"FF",X"FF",X"FF",X"00",X"80",X"80",X"83",X"C6",X"CC",X"E8",X"F9",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"21",X"21",X"3F",X"3F",X"21",X"21",X"2C",X"2C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2E",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2E",X"2E",X"2C",X"2C",X"2C",X"2C",X"2F",X"2F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2F",X"2F",X"2F",X"2F",X"2F",X"2E",X"2C",X"2C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"06",X"04",X"0C",X"09",X"09",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1B",X"13",X"13",X"37",X"27",X"27",X"2F",X"2E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2C",X"2C",X"21",X"21",X"3F",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2F",X"2F",X"2E",X"2E",X"2E",X"2C",X"2C",X"2D",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"2C",X"2C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2C",X"2D",X"21",X"21",X"3F",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"20",X"20",X"2F",X"2F",X"2F",X"2F",X"2F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2E",X"2C",X"2C",X"2D",X"2D",X"2D",X"2C",X"2C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"06",X"0C",X"08",X"19",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"13",X"13",X"37",X"27",X"27",X"2F",X"2F",X"2E",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"F8",X"F0",X"F0",X"E0",X"C0",X"C0",X"80",
		X"FF",X"7F",X"7E",X"3C",X"3C",X"18",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"01",X"00",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"80",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"03",X"00",X"F8",X"FF",X"F8",X"F8",X"FC",
		X"FF",X"FF",X"FF",X"FF",X"E0",X"80",X"0F",X"39",X"FF",X"FF",X"FF",X"FF",X"7F",X"1F",X"07",X"C3",
		X"60",X"C0",X"C0",X"E0",X"E0",X"F0",X"1F",X"00",X"71",X"38",X"2C",X"26",X"23",X"21",X"C1",X"7F",
		X"3F",X"00",X"80",X"FE",X"03",X"00",X"00",X"00",X"FF",X"FF",X"03",X"00",X"F8",X"2F",X"20",X"20",
		X"00",X"00",X"FF",X"80",X"00",X"3F",X"FF",X"FF",X"20",X"00",X"F8",X"0F",X"01",X"E0",X"FC",X"FF",
		X"FE",X"03",X"00",X"00",X"00",X"80",X"F0",X"1F",X"00",X"F8",X"2F",X"20",X"20",X"20",X"20",X"C0",
		X"00",X"C0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"01",X"00",X"FC",X"FF",X"FF",X"FF",X"FF",
		X"40",X"C0",X"80",X"F0",X"1F",X"00",X"C0",X"FF",X"20",X"20",X"20",X"20",X"C0",X"7F",X"01",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"80",X"80",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"1F",X"F0",X"80",X"07",X"3F",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"FC",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FC",X"E0",X"81",X"0F",X"38",X"60",X"FF",X"FF",X"03",X"00",X"F8",X"2F",X"20",X"20",
		X"C0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"01",X"00",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"80",X"FE",X"03",X"00",X"00",X"00",X"00",X"FF",X"03",X"00",X"F8",X"2F",X"20",X"20",X"20",
		X"07",X"1C",X"70",X"40",X"C0",X"80",X"80",X"80",X"A0",X"27",X"24",X"24",X"25",X"24",X"24",X"27",
		X"00",X"00",X"00",X"00",X"00",X"F0",X"1F",X"00",X"21",X"20",X"20",X"20",X"20",X"20",X"C0",X"7F",
		X"00",X"C0",X"7E",X"03",X"00",X"00",X"00",X"00",X"FF",X"03",X"00",X"F8",X"2F",X"20",X"20",X"20",
		X"F0",X"1F",X"00",X"C0",X"FE",X"FE",X"F0",X"C0",X"20",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",
		X"60",X"C0",X"80",X"80",X"80",X"F0",X"1F",X"00",X"71",X"38",X"2C",X"26",X"23",X"21",X"C1",X"7F",
		X"C0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"FF",X"80",X"00",X"3F",X"FF",X"FF",X"20",X"00",X"F8",X"0F",X"01",X"E0",X"FC",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"E0",X"80",X"0F",X"39",X"FF",X"FF",X"FF",X"FF",X"7F",X"1F",X"07",X"C3",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"9F",X"1F",X"1E",X"FE",X"FF",X"FF",X"FF",X"FF",X"C0",X"00",X"1F",X"00",X"C0",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"07",X"00",X"E0",X"3F",X"00",X"00",X"FF",X"FF",X"FF",X"3F",X"00",X"80",X"FE",X"03",
		X"98",X"C8",X"CC",X"E4",X"E4",X"F6",X"F2",X"F2",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"FF",
		X"FB",X"FA",X"78",X"78",X"39",X"3B",X"BF",X"9F",X"80",X"00",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"0F",X"00",X"E0",X"3F",X"00",X"FF",X"FF",X"FF",X"FF",X"3F",X"00",X"80",X"FE",
		X"00",X"00",X"00",X"00",X"C0",X"60",X"30",X"10",X"03",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
		X"0F",X"00",X"E0",X"3F",X"00",X"00",X"00",X"00",X"FF",X"3F",X"00",X"80",X"FE",X"03",X"00",X"00",
		X"00",X"FC",X"07",X"00",X"F0",X"FF",X"FF",X"FF",X"00",X"00",X"F0",X"1F",X"00",X"C0",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"07",X"F0",X"1E",X"03",X"00",X"00",X"00",X"00",X"F0",
		X"00",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"00",X"C0",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"FC",X"07",X"00",X"F0",X"FF",X"FF",X"FF",X"00",X"00",X"E0",X"3E",X"03",X"80",X"F8",X"FF",
		X"FF",X"FF",X"FF",X"1F",X"01",X"C0",X"7C",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"00",X"80",
		X"DA",X"1B",X"18",X"F8",X"FF",X"FF",X"FF",X"FF",X"00",X"F0",X"1F",X"00",X"C0",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"0F",X"00",X"E0",X"3F",X"00",X"00",X"FF",X"FF",X"FF",X"3F",X"00",X"80",X"FE",X"03",
		X"00",X"FC",X"07",X"00",X"F0",X"7F",X"3E",X"3C",X"01",X"01",X"E1",X"21",X"21",X"A0",X"20",X"20",
		X"9C",X"99",X"D9",X"5B",X"5A",X"5A",X"5A",X"5A",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"07",X"00",X"E0",X"3F",X"00",X"00",X"FF",X"FF",X"FF",X"3F",X"00",X"80",X"FE",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
		X"FB",X"FA",X"78",X"78",X"39",X"3B",X"BF",X"9F",X"80",X"00",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"9F",X"1F",X"1E",X"FE",X"FF",X"FF",X"FF",X"FF",X"C0",X"00",X"1F",X"00",X"C0",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"C0",X"60",X"30",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
		X"98",X"C8",X"CC",X"E4",X"E4",X"F6",X"F2",X"F2",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"FF",
		X"0F",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"34",X"84",X"84",X"FC",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"7F",X"01",X"00",X"FC",X"FF",X"30",X"FC",X"84",X"84",X"34",X"34",X"74",X"F4",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"03",X"00",X"F8",X"F4",X"F4",X"F4",X"F4",X"F4",X"F4",X"74",X"34",
		X"3F",X"7F",X"71",X"20",X"04",X"8E",X"FC",X"F0",X"88",X"CC",X"E4",X"E4",X"F4",X"74",X"74",X"F4",
		X"01",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"F4",X"F4",X"F4",X"E4",X"E4",X"C4",X"8C",X"18",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"03",X"F4",X"F4",X"F4",X"F4",X"F4",X"F4",X"F4",X"F4",
		X"00",X"F8",X"0F",X"01",X"7F",X"C0",X"80",X"1E",X"74",X"34",X"34",X"84",X"84",X"FC",X"30",X"18",
		X"FF",X"FF",X"FF",X"03",X"00",X"F8",X"0F",X"01",X"F4",X"F4",X"F4",X"F4",X"74",X"34",X"34",X"84",
		X"00",X"00",X"00",X"C0",X"7F",X"01",X"00",X"FC",X"84",X"FC",X"FC",X"84",X"84",X"34",X"34",X"74",
		X"3F",X"0F",X"87",X"E3",X"31",X"19",X"0C",X"04",X"90",X"D8",X"C8",X"C8",X"E8",X"EC",X"E4",X"E4",
		X"C6",X"7E",X"00",X"00",X"FC",X"FF",X"FF",X"FF",X"F4",X"74",X"74",X"74",X"74",X"F4",X"F4",X"F4",
		X"0F",X"01",X"00",X"00",X"C0",X"70",X"1C",X"06",X"34",X"84",X"84",X"FC",X"00",X"00",X"00",X"00",
		X"C3",X"F1",X"F8",X"FC",X"FE",X"FF",X"FF",X"FF",X"00",X"80",X"C0",X"40",X"60",X"20",X"30",X"90",
		X"00",X"00",X"C0",X"7F",X"01",X"00",X"FC",X"FF",X"B4",X"B4",X"B4",X"B4",X"B4",X"34",X"34",X"F4",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"03",X"00",X"F8",X"F4",X"F4",X"F4",X"F4",X"F4",X"F4",X"74",X"34",
		X"00",X"7C",X"0F",X"03",X"E1",X"38",X"0C",X"06",X"04",X"04",X"F4",X"F4",X"F4",X"F4",X"F4",X"74",
		X"02",X"03",X"01",X"01",X"01",X"00",X"00",X"00",X"74",X"74",X"34",X"34",X"B4",X"B4",X"B4",X"B4",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"03",X"00",X"F8",X"F4",X"F4",X"F4",X"F4",X"F4",X"F4",X"74",X"34",
		X"0F",X"01",X"00",X"00",X"00",X"00",X"FF",X"01",X"34",X"84",X"84",X"FC",X"00",X"00",X"00",X"FC",
		X"01",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"F4",X"F4",X"F4",X"E4",X"E4",X"C4",X"8C",X"18",
		X"00",X"00",X"FF",X"7F",X"01",X"00",X"FC",X"FF",X"30",X"FC",X"84",X"84",X"34",X"34",X"74",X"F4",
		X"00",X"00",X"00",X"00",X"7F",X"C0",X"80",X"1E",X"00",X"00",X"00",X"00",X"80",X"E0",X"30",X"18",
		X"3F",X"7F",X"71",X"20",X"04",X"8E",X"FC",X"F0",X"88",X"CC",X"E4",X"E4",X"F4",X"74",X"74",X"F4",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"0C",X"1A",X"67",X"7E",X"23",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"07",X"10",X"70",X"60",X"00",X"00",X"00",X"00",X"80",X"40",X"20",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"02",X"20",X"23",X"7E",X"27",X"1A",X"0C",X"06",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"00",X"00",X"00",X"00",X"01",X"08",X"15",X"AA",
		X"15",X"B0",X"E0",X"06",X"0F",X"16",X"10",X"16",X"FF",X"FF",X"5D",X"2B",X"05",X"80",X"40",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"40",X"A8",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"F8",X"54",X"A0",X"FC",X"A9",X"00",X"00",X"00",X"00",X"00",X"03",X"08",X"80",X"E0",X"00",
		X"01",X"1E",X"15",X"05",X"06",X"E0",X"B0",X"05",X"60",X"C0",X"40",X"15",X"2B",X"5D",X"FF",X"57",
		X"E0",X"3C",X"07",X"00",X"00",X"00",X"00",X"00",X"AA",X"00",X"80",X"F0",X"1F",X"01",X"00",X"00",
		X"00",X"14",X"AD",X"FD",X"F4",X"54",X"A8",X"F0",X"00",X"80",X"E0",X"F0",X"04",X"00",X"00",X"00",
		X"70",X"A8",X"00",X"00",X"00",X"F0",X"1E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"0C",X"1A",X"67",X"7E",X"23",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"F7",X"F0",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"60",X"30",X"10",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"02",X"20",X"23",X"7E",X"27",X"1A",X"0C",X"06",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"02",X"15",X"AA",X"55",
		X"16",X"B0",X"E0",X"06",X"0F",X"16",X"10",X"16",X"00",X"00",X"20",X"14",X"1A",X"8F",X"47",X"E7",
		X"00",X"00",X"00",X"08",X"24",X"BC",X"58",X"A4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"0A",X"5B",X"F7",X"F0",X"00",X"00",X"00",X"03",X"08",X"80",X"E0",X"00",
		X"01",X"1E",X"15",X"05",X"06",X"E0",X"B0",X"FA",X"67",X"C7",X"4F",X"0A",X"14",X"20",X"00",X"A8",
		X"1F",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"FF",X"7F",X"0F",X"00",X"00",X"00",X"00",
		X"F0",X"E7",X"53",X"03",X"08",X"00",X"02",X"00",X"00",X"80",X"E0",X"F0",X"04",X"00",X"00",X"00",
		X"8C",X"54",X"FC",X"FC",X"F8",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"18",X"10",X"13",X"10",X"18",X"10",X"13",X"FE",X"02",X"02",X"F2",X"06",X"02",X"02",X"F2",
		X"30",X"60",X"40",X"40",X"4E",X"46",X"6F",X"38",X"03",X"01",X"01",X"01",X"79",X"D9",X"93",X"1E",
		X"FF",X"FF",X"C0",X"DF",X"DF",X"DF",X"DF",X"DF",X"FE",X"FC",X"00",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"DF",X"DF",X"DF",X"DF",X"DF",X"C0",X"80",X"00",X"F8",X"F8",X"F8",X"F8",X"F8",X"00",X"00",X"00",
		X"FF",X"FF",X"C0",X"DF",X"DF",X"DF",X"DF",X"DF",X"FE",X"FC",X"00",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"DF",X"DF",X"DF",X"DF",X"DF",X"C0",X"80",X"00",X"F8",X"F8",X"F8",X"F8",X"F8",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
