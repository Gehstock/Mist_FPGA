library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity spr1_rom is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of spr1_rom is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"EE",X"1D",X"22",X"00",X"88",X"D1",X"40",X"00",X"80",X"58",X"C0",X"00",
		X"08",X"D0",X"84",X"10",X"80",X"B4",X"F3",X"30",X"80",X"E9",X"7B",X"52",X"C0",X"78",X"D7",X"70",
		X"A4",X"69",X"0F",X"70",X"E0",X"F0",X"09",X"52",X"62",X"52",X"0F",X"30",X"62",X"30",X"06",X"00",
		X"22",X"30",X"00",X"00",X"22",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"80",X"00",X"80",X"10",X"80",X"10",
		X"C0",X"30",X"48",X"30",X"84",X"34",X"F3",X"52",X"A4",X"E9",X"7B",X"70",X"E0",X"78",X"D7",X"70",
		X"68",X"78",X"0F",X"52",X"E2",X"D2",X"09",X"70",X"A2",X"70",X"0F",X"30",X"22",X"21",X"06",X"00",
		X"22",X"30",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"22",X"00",X"30",X"00",X"10",X"00",X"12",X"80",X"10",
		X"00",X"70",X"48",X"30",X"E2",X"E1",X"F3",X"30",X"E2",X"F8",X"7B",X"52",X"E2",X"5A",X"D7",X"70",
		X"2A",X"78",X"0F",X"52",X"A2",X"D2",X"09",X"70",X"88",X"F0",X"0F",X"30",X"88",X"94",X"06",X"00",
		X"88",X"C0",X"00",X"00",X"88",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"30",X"00",X"00",X"A4",X"52",X"00",X"00",X"F0",X"70",X"00",
		X"80",X"B4",X"07",X"00",X"C0",X"E9",X"0D",X"00",X"22",X"6E",X"0D",X"00",X"00",X"EE",X"07",X"00",
		X"4A",X"7C",X"21",X"00",X"C2",X"D2",X"70",X"00",X"00",X"E0",X"B4",X"12",X"E6",X"B4",X"E1",X"12",
		X"E6",X"E1",X"30",X"00",X"22",X"80",X"E1",X"00",X"22",X"00",X"FC",X"33",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"30",X"00",X"00",X"D2",X"61",X"00",X"A2",X"F0",X"70",X"00",
		X"C0",X"A5",X"07",X"00",X"00",X"F8",X"0D",X"00",X"00",X"6E",X"0D",X"00",X"00",X"EE",X"07",X"00",
		X"00",X"4C",X"21",X"00",X"00",X"C4",X"70",X"00",X"00",X"F0",X"D2",X"12",X"80",X"B4",X"78",X"12",
		X"80",X"F0",X"61",X"00",X"00",X"96",X"30",X"00",X"00",X"C0",X"FE",X"11",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"30",X"00",X"22",X"B4",X"61",X"00",X"C0",X"F0",X"70",X"00",
		X"80",X"A5",X"07",X"00",X"00",X"F8",X"0D",X"00",X"00",X"6E",X"0D",X"00",X"00",X"EE",X"07",X"00",
		X"00",X"6C",X"E1",X"12",X"00",X"F0",X"78",X"12",X"4A",X"78",X"52",X"00",X"C2",X"D2",X"F0",X"00",
		X"00",X"E0",X"ED",X"33",X"00",X"E0",X"00",X"00",X"00",X"EE",X"33",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"11",X"22",X"00",X"88",X"11",X"40",X"00",X"80",X"10",X"C0",X"00",X"08",X"30",X"84",X"10",
		X"80",X"70",X"F3",X"30",X"80",X"DA",X"7B",X"52",X"C0",X"78",X"D7",X"70",X"A4",X"69",X"0F",X"70",
		X"E0",X"F0",X"09",X"52",X"62",X"52",X"0F",X"30",X"62",X"30",X"06",X"00",X"22",X"34",X"00",X"00",
		X"2A",X"3C",X"00",X"00",X"08",X"0F",X"00",X"00",X"08",X"0F",X"00",X"00",X"00",X"07",X"00",X"00",
		X"00",X"00",X"00",X"11",X"00",X"00",X"80",X"00",X"00",X"00",X"80",X"10",X"80",X"30",X"48",X"30",
		X"48",X"70",X"F3",X"52",X"E0",X"DA",X"7B",X"70",X"A4",X"78",X"D7",X"70",X"E0",X"69",X"0F",X"52",
		X"E2",X"F0",X"09",X"70",X"A2",X"61",X"0F",X"30",X"22",X"30",X"06",X"00",X"22",X"34",X"00",X"00",
		X"08",X"3C",X"00",X"00",X"08",X"0F",X"00",X"00",X"08",X"0F",X"00",X"00",X"00",X"07",X"00",X"00",
		X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"40",X"E2",X"10",X"00",X"60",X"E2",X"61",X"80",X"70",
		X"E2",X"F0",X"F3",X"52",X"6A",X"DA",X"7B",X"70",X"A2",X"78",X"D7",X"52",X"C0",X"78",X"0F",X"30",
		X"68",X"D2",X"09",X"30",X"E0",X"60",X"0F",X"10",X"62",X"60",X"06",X"00",X"22",X"68",X"00",X"00",
		X"22",X"69",X"01",X"00",X"22",X"0F",X"01",X"00",X"00",X"0F",X"01",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"10",X"00",X"00",X"D2",X"21",X"00",X"80",X"F0",X"30",X"00",
		X"C0",X"5A",X"03",X"00",X"68",X"7C",X"06",X"00",X"11",X"3F",X"06",X"00",X"00",X"7F",X"03",X"00",
		X"00",X"2E",X"10",X"07",X"00",X"F0",X"38",X"0F",X"80",X"D2",X"D2",X"1E",X"F3",X"78",X"F0",X"1E",
		X"7B",X"F0",X"10",X"07",X"11",X"48",X"70",X"00",X"11",X"80",X"FE",X"11",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"F0",X"10",X"00",X"80",X"69",X"30",X"00",X"D1",X"F0",X"30",X"00",
		X"68",X"5A",X"03",X"00",X"80",X"7C",X"06",X"00",X"00",X"3F",X"06",X"00",X"00",X"7F",X"03",X"00",
		X"00",X"2E",X"10",X"07",X"00",X"F0",X"38",X"0F",X"80",X"D2",X"F0",X"1E",X"80",X"78",X"D2",X"1E",
		X"80",X"E1",X"30",X"07",X"00",X"D2",X"10",X"00",X"00",X"E0",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"11",X"00",X"00",X"00",X"E0",X"70",X"00",X"00",X"C0",X"A5",X"10",X"00",X"80",X"F0",X"30",X"00",
		X"80",X"5A",X"03",X"00",X"00",X"7C",X"06",X"00",X"00",X"3F",X"06",X"00",X"00",X"7F",X"03",X"07",
		X"00",X"3E",X"18",X"0F",X"80",X"F0",X"F0",X"1E",X"80",X"D2",X"E1",X"1E",X"48",X"F0",X"10",X"07",
		X"C0",X"D2",X"21",X"00",X"C0",X"B0",X"70",X"00",X"CC",X"77",X"FC",X"33",X"00",X"00",X"00",X"00",
		X"EE",X"11",X"00",X"00",X"88",X"11",X"22",X"00",X"80",X"10",X"40",X"00",X"80",X"30",X"C0",X"00",
		X"80",X"61",X"84",X"10",X"80",X"F0",X"F3",X"21",X"C0",X"E9",X"F3",X"70",X"E0",X"78",X"D7",X"61",
		X"52",X"69",X"0F",X"70",X"62",X"B4",X"09",X"52",X"22",X"E0",X"0F",X"30",X"22",X"C0",X"16",X"00",
		X"22",X"00",X"70",X"00",X"00",X"00",X"2C",X"00",X"00",X"00",X"0C",X"01",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"80",X"00",
		X"80",X"70",X"80",X"10",X"6A",X"D2",X"48",X"30",X"E2",X"F0",X"F3",X"52",X"6A",X"DA",X"7B",X"70",
		X"A2",X"78",X"D7",X"70",X"22",X"5A",X"0F",X"52",X"00",X"F0",X"09",X"70",X"08",X"A1",X"0F",X"30",
		X"0C",X"80",X"16",X"00",X"00",X"80",X"10",X"00",X"00",X"08",X"03",X"00",X"00",X"00",X"02",X"00",
		X"00",X"07",X"00",X"00",X"00",X"03",X"00",X"22",X"62",X"30",X"00",X"40",X"E2",X"30",X"00",X"60",
		X"6A",X"70",X"80",X"70",X"E2",X"D2",X"F3",X"52",X"A2",X"F8",X"7B",X"70",X"80",X"5A",X"D7",X"52",
		X"E2",X"78",X"0F",X"30",X"6A",X"D2",X"09",X"30",X"E2",X"70",X"0F",X"10",X"A2",X"10",X"06",X"00",
		X"A2",X"10",X"00",X"00",X"08",X"01",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"30",X"00",X"00",X"20",X"52",X"00",X"00",X"5A",X"70",X"0C",
		X"80",X"F0",X"07",X"06",X"C0",X"E9",X"0D",X"16",X"22",X"6E",X"0D",X"30",X"00",X"EE",X"87",X"10",
		X"00",X"6A",X"E1",X"00",X"00",X"F0",X"D2",X"00",X"80",X"F0",X"70",X"00",X"F3",X"A5",X"21",X"00",
		X"F3",X"F0",X"10",X"00",X"11",X"C0",X"21",X"00",X"11",X"80",X"FE",X"11",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"70",X"00",X"00",X"A4",X"D2",X"00",X"44",X"F0",X"F0",X"00",
		X"80",X"5A",X"1E",X"00",X"00",X"E0",X"1B",X"01",X"00",X"CC",X"0B",X"0D",X"00",X"CC",X"1F",X"34",
		X"00",X"E8",X"C3",X"34",X"00",X"F0",X"70",X"00",X"00",X"5A",X"D2",X"00",X"00",X"F0",X"78",X"00",
		X"00",X"5A",X"18",X"01",X"00",X"E0",X"00",X"01",X"00",X"EE",X"33",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"F0",X"00",X"00",X"A2",X"5A",X"30",X"00",X"00",X"F0",X"70",X"00",
		X"00",X"B4",X"07",X"00",X"00",X"E8",X"0D",X"00",X"00",X"6E",X"0D",X"00",X"00",X"EE",X"07",X"00",
		X"00",X"6A",X"21",X"00",X"01",X"F0",X"70",X"00",X"C3",X"5A",X"52",X"00",X"C3",X"F0",X"F0",X"12",
		X"80",X"E1",X"D2",X"16",X"C0",X"30",X"70",X"04",X"CC",X"77",X"FF",X"11",X"00",X"00",X"00",X"00",
		X"EE",X"11",X"00",X"00",X"88",X"1F",X"22",X"00",X"80",X"1E",X"41",X"00",X"80",X"3C",X"C1",X"00",
		X"80",X"69",X"85",X"10",X"80",X"F0",X"F3",X"21",X"C0",X"E9",X"F3",X"70",X"E0",X"78",X"D7",X"61",
		X"A4",X"69",X"0F",X"70",X"62",X"B4",X"09",X"52",X"22",X"E0",X"0F",X"30",X"22",X"C0",X"16",X"00",
		X"22",X"00",X"70",X"00",X"00",X"00",X"2C",X"00",X"00",X"00",X"0C",X"01",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"01",X"11",X"00",X"0E",X"83",X"00",
		X"80",X"78",X"83",X"10",X"6A",X"D2",X"4B",X"30",X"E2",X"F0",X"F3",X"52",X"6A",X"DA",X"7B",X"70",
		X"A2",X"78",X"D7",X"70",X"22",X"5A",X"0F",X"52",X"00",X"F0",X"09",X"70",X"08",X"A1",X"0F",X"30",
		X"0C",X"80",X"16",X"00",X"00",X"80",X"10",X"00",X"00",X"08",X"03",X"00",X"00",X"00",X"02",X"00",
		X"00",X"07",X"00",X"00",X"00",X"03",X"00",X"22",X"62",X"38",X"03",X"40",X"E2",X"3C",X"07",X"60",
		X"6A",X"78",X"87",X"70",X"E2",X"D2",X"F3",X"52",X"A2",X"F8",X"7B",X"70",X"80",X"5A",X"D7",X"52",
		X"E2",X"78",X"0F",X"30",X"6A",X"D2",X"09",X"30",X"E2",X"70",X"0F",X"10",X"A2",X"10",X"06",X"00",
		X"A2",X"10",X"00",X"00",X"08",X"01",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"30",X"00",X"00",X"E0",X"52",X"00",X"00",X"5A",X"70",X"0C",
		X"80",X"F0",X"07",X"06",X"C0",X"E9",X"0D",X"16",X"22",X"6E",X"0D",X"30",X"0C",X"EF",X"87",X"10",
		X"0E",X"6D",X"E1",X"00",X"0E",X"F0",X"D2",X"00",X"86",X"F0",X"70",X"00",X"F3",X"A5",X"21",X"00",
		X"F3",X"F0",X"10",X"00",X"11",X"C0",X"21",X"00",X"11",X"80",X"FE",X"11",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"70",X"00",X"00",X"A4",X"D2",X"00",X"44",X"F0",X"F0",X"00",
		X"80",X"5A",X"1E",X"00",X"00",X"E0",X"1B",X"01",X"08",X"CF",X"0B",X"0D",X"0C",X"CF",X"1F",X"34",
		X"0C",X"E9",X"C3",X"34",X"0C",X"F0",X"70",X"00",X"08",X"5A",X"D2",X"00",X"00",X"F0",X"78",X"00",
		X"00",X"5A",X"18",X"01",X"00",X"E0",X"00",X"01",X"00",X"EE",X"33",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"F0",X"00",X"00",X"A2",X"5A",X"30",X"00",X"00",X"F0",X"70",X"00",
		X"00",X"B4",X"07",X"00",X"08",X"E9",X"0D",X"00",X"0C",X"6F",X"0D",X"00",X"0C",X"EF",X"07",X"00",
		X"0C",X"6D",X"B1",X"00",X"09",X"F0",X"70",X"00",X"C3",X"5A",X"52",X"00",X"C3",X"F0",X"F0",X"12",
		X"80",X"E1",X"D2",X"16",X"C0",X"30",X"70",X"04",X"CC",X"77",X"FF",X"11",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"EE",X"11",X"00",X"00",X"88",X"11",X"22",X"00",X"80",X"10",X"40",X"00",
		X"08",X"10",X"C0",X"00",X"80",X"30",X"84",X"10",X"80",X"52",X"F3",X"30",X"48",X"F8",X"7B",X"52",
		X"E0",X"78",X"D7",X"70",X"E0",X"69",X"0F",X"70",X"62",X"F0",X"09",X"52",X"22",X"52",X"0F",X"30",
		X"22",X"30",X"06",X"00",X"22",X"30",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"07",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",
		X"00",X"70",X"80",X"00",X"80",X"D2",X"80",X"10",X"6A",X"F0",X"48",X"30",X"E2",X"D2",X"F3",X"52",
		X"E2",X"F8",X"7B",X"70",X"A2",X"69",X"D7",X"70",X"22",X"78",X"0F",X"52",X"00",X"30",X"09",X"70",
		X"00",X"30",X"0F",X"30",X"00",X"30",X"06",X"00",X"00",X"03",X"00",X"00",X"00",X"07",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"62",X"00",X"00",X"00",X"E2",X"00",X"00",X"00",
		X"6A",X"10",X"00",X"22",X"E2",X"30",X"00",X"40",X"A2",X"61",X"00",X"60",X"80",X"B4",X"80",X"70",
		X"C0",X"E1",X"F3",X"52",X"C0",X"F8",X"7B",X"70",X"C4",X"69",X"D7",X"52",X"44",X"78",X"0F",X"30",
		X"44",X"30",X"09",X"30",X"44",X"30",X"0F",X"10",X"00",X"03",X"06",X"00",X"00",X"07",X"00",X"00",
		X"00",X"00",X"00",X"00",X"EE",X"11",X"00",X"00",X"88",X"11",X"22",X"00",X"80",X"1C",X"40",X"00",
		X"80",X"1E",X"C1",X"00",X"80",X"2D",X"85",X"10",X"80",X"78",X"F3",X"30",X"C0",X"E9",X"7B",X"52",
		X"E0",X"78",X"D7",X"70",X"A4",X"69",X"0F",X"70",X"62",X"F0",X"09",X"52",X"22",X"52",X"0F",X"30",
		X"22",X"30",X"06",X"00",X"22",X"30",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"07",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"01",X"11",
		X"00",X"78",X"83",X"00",X"80",X"D2",X"83",X"10",X"6A",X"F0",X"4B",X"30",X"E2",X"D2",X"F3",X"52",
		X"E2",X"F8",X"7B",X"70",X"A2",X"69",X"D7",X"70",X"22",X"78",X"0F",X"52",X"00",X"30",X"09",X"70",
		X"00",X"30",X"0F",X"30",X"00",X"30",X"06",X"00",X"00",X"03",X"00",X"00",X"00",X"07",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"62",X"00",X"00",X"00",X"E2",X"00",X"00",X"00",
		X"6A",X"1C",X"01",X"22",X"E2",X"3C",X"03",X"40",X"A2",X"69",X"03",X"60",X"80",X"B4",X"83",X"70",
		X"C0",X"E1",X"F3",X"52",X"C0",X"F8",X"7B",X"70",X"C4",X"69",X"D7",X"52",X"44",X"78",X"0F",X"30",
		X"44",X"30",X"09",X"30",X"44",X"30",X"0F",X"10",X"00",X"03",X"06",X"00",X"00",X"07",X"00",X"00",
		X"00",X"06",X"22",X"00",X"00",X"0F",X"40",X"00",X"00",X"0F",X"C0",X"00",X"00",X"16",X"84",X"10",
		X"00",X"30",X"F3",X"30",X"A6",X"F8",X"7B",X"52",X"E2",X"5A",X"D7",X"70",X"6A",X"78",X"0F",X"70",
		X"A2",X"F0",X"09",X"52",X"A2",X"A5",X"0F",X"30",X"80",X"D0",X"06",X"00",X"80",X"D0",X"00",X"00",
		X"88",X"1D",X"00",X"00",X"88",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"1D",X"00",X"22",X"88",X"D1",X"00",X"40",X"80",X"58",X"00",X"60",X"80",X"D0",X"80",X"70",
		X"80",X"E1",X"F3",X"52",X"80",X"BC",X"7B",X"70",X"C0",X"69",X"D7",X"52",X"A4",X"78",X"0F",X"30",
		X"E0",X"E1",X"09",X"30",X"62",X"70",X"0F",X"10",X"62",X"30",X"06",X"00",X"22",X"30",X"00",X"00",
		X"22",X"03",X"03",X"00",X"00",X"08",X"07",X"00",X"00",X"08",X"07",X"00",X"00",X"00",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"10",X"00",X"00",X"D2",X"21",X"00",X"80",X"F0",X"30",X"00",
		X"C0",X"5A",X"03",X"00",X"68",X"7C",X"06",X"00",X"11",X"3F",X"06",X"00",X"00",X"7F",X"03",X"00",
		X"06",X"2E",X"F0",X"01",X"0F",X"E0",X"D2",X"23",X"0F",X"B4",X"30",X"22",X"86",X"F0",X"D2",X"33",
		X"00",X"68",X"F0",X"33",X"00",X"C2",X"00",X"00",X"00",X"EE",X"33",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"E0",X"70",X"00",X"00",X"D1",X"A5",X"10",X"00",X"80",X"F0",X"30",X"00",
		X"80",X"5A",X"03",X"00",X"00",X"7C",X"06",X"06",X"00",X"3F",X"06",X"0F",X"00",X"7F",X"03",X"0F",
		X"A5",X"3E",X"10",X"06",X"E1",X"D2",X"30",X"00",X"00",X"F0",X"F0",X"01",X"F3",X"A5",X"E1",X"01",
		X"F3",X"F0",X"10",X"00",X"11",X"48",X"70",X"00",X"11",X"80",X"FE",X"11",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"EE",X"11",X"00",X"00",X"60",X"44",X"00",X"00",X"A4",X"80",X"00",X"00",
		X"E0",X"E3",X"00",X"00",X"4A",X"6B",X"00",X"00",X"4A",X"C2",X"00",X"00",X"68",X"C3",X"00",X"00",
		X"68",X"4B",X"00",X"00",X"4A",X"C2",X"00",X"00",X"4A",X"A7",X"00",X"00",X"E0",X"63",X"00",X"00",
		X"A4",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"EE",X"11",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"79",X"10",X"44",X"00",X"C0",X"30",X"44",X"08",X"49",X"70",X"C4",X"90",X"90",X"52",
		X"4C",X"B0",X"B0",X"70",X"C0",X"52",X"12",X"00",X"80",X"F0",X"38",X"33",X"00",X"5A",X"3C",X"67",
		X"00",X"F0",X"12",X"07",X"80",X"5A",X"1E",X"07",X"E0",X"F0",X"1E",X"07",X"A4",X"69",X"12",X"07",
		X"E2",X"90",X"3C",X"67",X"22",X"00",X"38",X"33",X"22",X"00",X"30",X"00",X"22",X"00",X"03",X"00",
		X"00",X"CC",X"77",X"00",X"00",X"00",X"60",X"00",X"84",X"10",X"F0",X"00",X"84",X"21",X"D2",X"00",
		X"80",X"F0",X"E0",X"10",X"00",X"DE",X"B4",X"10",X"00",X"8F",X"F1",X"21",X"0A",X"0C",X"A5",X"30",
		X"4A",X"0F",X"E1",X"10",X"68",X"0F",X"A5",X"21",X"48",X"0C",X"E1",X"30",X"00",X"8F",X"B5",X"10",
		X"00",X"CE",X"F0",X"00",X"00",X"E0",X"30",X"00",X"CC",X"F3",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"48",X"00",X"00",X"22",X"C0",X"00",X"00",X"22",
		X"48",X"F3",X"70",X"66",X"0C",X"E7",X"B4",X"74",X"02",X"87",X"E1",X"65",X"0E",X"87",X"B4",X"54",
		X"0E",X"87",X"61",X"00",X"02",X"87",X"70",X"00",X"0C",X"E7",X"A5",X"00",X"48",X"F3",X"F0",X"10",
		X"C0",X"00",X"68",X"10",X"84",X"00",X"C0",X"32",X"C0",X"00",X"88",X"33",X"0C",X"00",X"FF",X"11",
		X"0C",X"CC",X"33",X"00",X"C0",X"C0",X"00",X"00",X"48",X"48",X"00",X"00",X"C0",X"C0",X"00",X"00",
		X"48",X"F3",X"10",X"00",X"0C",X"E7",X"21",X"07",X"02",X"87",X"30",X"05",X"0E",X"87",X"01",X"05",
		X"0E",X"87",X"10",X"05",X"02",X"87",X"21",X"05",X"0C",X"E7",X"30",X"07",X"48",X"F3",X"10",X"00",
		X"C0",X"48",X"00",X"00",X"84",X"C0",X"00",X"00",X"C0",X"C0",X"00",X"00",X"0C",X"CC",X"33",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"FF",X"11",X"00",X"CC",X"FF",X"3B",X"01",
		X"88",X"F7",X"3F",X"03",X"00",X"F3",X"36",X"03",X"88",X"73",X"36",X"03",X"CC",X"73",X"7E",X"01",
		X"CC",X"73",X"FE",X"00",X"88",X"73",X"7E",X"01",X"00",X"73",X"3E",X"03",X"88",X"73",X"36",X"03",
		X"CC",X"73",X"36",X"03",X"88",X"73",X"3A",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"FF",X"33",X"00",X"CC",X"FF",X"77",X"03",
		X"88",X"F1",X"7E",X"07",X"EE",X"30",X"7C",X"04",X"CC",X"10",X"6C",X"04",X"88",X"10",X"EC",X"03",
		X"88",X"10",X"EC",X"11",X"CC",X"10",X"EC",X"03",X"EE",X"10",X"6C",X"07",X"88",X"10",X"6C",X"04",
		X"CC",X"10",X"6C",X"04",X"EE",X"10",X"64",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"0C",X"01",X"08",X"0F",X"0E",X"03",
		X"08",X"09",X"17",X"02",X"00",X"8F",X"3F",X"01",X"88",X"FF",X"FF",X"33",X"CC",X"F1",X"F0",X"30",
		X"CC",X"30",X"00",X"00",X"CC",X"F1",X"F0",X"30",X"CC",X"FF",X"FF",X"33",X"CC",X"FF",X"FF",X"33",
		X"CC",X"DD",X"BB",X"33",X"88",X"88",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"07",X"0C",X"01",X"08",X"09",X"06",X"02",X"08",X"09",X"17",X"02",
		X"00",X"8F",X"3F",X"01",X"88",X"FF",X"FF",X"33",X"CC",X"F1",X"F0",X"30",X"CC",X"30",X"00",X"00",
		X"CC",X"10",X"00",X"00",X"CC",X"10",X"00",X"00",X"CC",X"30",X"00",X"00",X"CC",X"F1",X"F0",X"30",
		X"CC",X"FF",X"FF",X"33",X"CC",X"66",X"66",X"33",X"44",X"22",X"44",X"22",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0C",X"00",X"88",X"AA",X"1F",X"01",X"CC",X"FF",X"13",X"01",X"88",X"FF",X"13",X"01",
		X"EE",X"FF",X"3F",X"11",X"CC",X"F1",X"F8",X"1F",X"EE",X"30",X"C0",X"19",X"E6",X"10",X"80",X"3A",
		X"F3",X"00",X"00",X"FC",X"71",X"00",X"00",X"E8",X"31",X"00",X"00",X"C8",X"31",X"00",X"00",X"C0",
		X"30",X"00",X"00",X"80",X"10",X"00",X"00",X"80",X"10",X"00",X"00",X"80",X"10",X"00",X"00",X"80",
		X"00",X"0E",X"F7",X"F0",X"00",X"02",X"F1",X"00",X"00",X"8A",X"30",X"00",X"0E",X"F7",X"10",X"00",
		X"03",X"E3",X"00",X"00",X"03",X"61",X"00",X"00",X"0E",X"31",X"00",X"00",X"EE",X"31",X"00",X"00",
		X"EE",X"31",X"00",X"00",X"CC",X"31",X"00",X"00",X"EE",X"71",X"00",X"01",X"CC",X"F3",X"00",X"00",
		X"EE",X"F7",X"10",X"00",X"44",X"FF",X"30",X"00",X"00",X"DD",X"F1",X"10",X"00",X"00",X"FF",X"F0",
		X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"C2",X"18",X"0F",X"00",X"C2",X"78",X"78",X"01",
		X"C2",X"B4",X"F0",X"01",X"C2",X"F0",X"F0",X"01",X"C2",X"F3",X"F0",X"01",X"C0",X"F3",X"87",X"01",
		X"C2",X"F3",X"84",X"01",X"C2",X"F3",X"84",X"01",X"C2",X"B7",X"F0",X"01",X"82",X"B7",X"78",X"01",
		X"02",X"3F",X"3C",X"00",X"00",X"3B",X"07",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"70",X"0F",X"01",X"86",X"F0",X"E1",X"03",
		X"0C",X"78",X"F0",X"12",X"08",X"E1",X"F0",X"12",X"80",X"FE",X"F0",X"12",X"80",X"FE",X"1F",X"12",
		X"80",X"F8",X"19",X"12",X"08",X"F8",X"19",X"12",X"0E",X"C8",X"F1",X"12",X"08",X"89",X"F1",X"03",
		X"00",X"8B",X"79",X"01",X"00",X"88",X"1F",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"08",X"F0",X"00",X"00",X"08",X"F0",X"1E",X"00",
		X"08",X"F0",X"69",X"03",X"08",X"F0",X"F0",X"12",X"08",X"F7",X"F0",X"16",X"88",X"F7",X"F0",X"34",
		X"88",X"F1",X"3C",X"25",X"88",X"F1",X"34",X"24",X"88",X"F1",X"34",X"24",X"88",X"D1",X"E1",X"34",
		X"88",X"11",X"C3",X"16",X"88",X"00",X"0E",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"0F",X"0F",X"00",
		X"0C",X"F0",X"78",X"01",X"84",X"78",X"C3",X"03",X"84",X"78",X"C0",X"12",X"84",X"78",X"C0",X"12",
		X"0C",X"F0",X"F0",X"03",X"80",X"E1",X"3C",X"01",X"80",X"FC",X"FF",X"33",X"C0",X"FC",X"FF",X"77",
		X"E0",X"F0",X"F0",X"00",X"C0",X"F0",X"70",X"00",X"0C",X"07",X"0F",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"0F",X"0F",X"00",X"0C",X"F0",X"78",X"01",
		X"84",X"78",X"C3",X"03",X"84",X"78",X"C0",X"12",X"84",X"78",X"C0",X"12",X"0C",X"F8",X"FF",X"33",
		X"80",X"ED",X"FF",X"77",X"E0",X"FC",X"70",X"00",X"C0",X"FC",X"30",X"01",X"C0",X"D2",X"38",X"01",
		X"80",X"C3",X"1E",X"00",X"08",X"01",X"04",X"00",X"08",X"00",X"04",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"0F",X"01",X"00",X"87",X"F0",X"03",X"00",X"E1",X"81",X"12",
		X"08",X"E1",X"81",X"12",X"08",X"F0",X"87",X"12",X"08",X"F0",X"F0",X"03",X"80",X"E1",X"78",X"01",
		X"C0",X"F0",X"F0",X"00",X"C0",X"FC",X"F0",X"00",X"C0",X"FC",X"70",X"00",X"E0",X"FC",X"FF",X"11",
		X"0C",X"8F",X"FF",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"40",X"60",X"00",X"84",X"D0",X"E0",X"00",X"84",X"F1",X"F4",X"10",
		X"84",X"FB",X"FD",X"30",X"8C",X"FE",X"FF",X"31",X"8C",X"9F",X"FE",X"73",X"80",X"1F",X"3F",X"77",
		X"8A",X"3F",X"2F",X"67",X"86",X"7A",X"2F",X"47",X"02",X"7F",X"07",X"46",X"02",X"EA",X"07",X"46",
		X"02",X"00",X"1E",X"23",X"00",X"00",X"8E",X"11",X"00",X"00",X"06",X"00",X"00",X"00",X"07",X"00",
		X"00",X"00",X"00",X"00",X"80",X"40",X"60",X"00",X"82",X"D0",X"E0",X"00",X"86",X"F1",X"F4",X"10",
		X"82",X"FB",X"FD",X"30",X"8A",X"FE",X"F0",X"31",X"8A",X"9F",X"FE",X"73",X"80",X"9F",X"3F",X"77",
		X"8C",X"97",X"3F",X"67",X"84",X"9F",X"3F",X"47",X"04",X"9F",X"36",X"46",X"04",X"8E",X"37",X"46",
		X"04",X"06",X"3E",X"23",X"00",X"06",X"EE",X"11",X"00",X"07",X"00",X"00",X"08",X"03",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"40",X"60",X"00",X"84",X"D0",X"E0",X"00",X"84",X"F1",X"F4",X"07",
		X"84",X"FB",X"1F",X"0F",X"8C",X"7E",X"0F",X"3D",X"8C",X"1F",X"CF",X"3F",X"80",X"1F",X"3F",X"7F",
		X"8A",X"F7",X"3F",X"67",X"86",X"FD",X"3F",X"47",X"02",X"FF",X"36",X"46",X"02",X"EA",X"37",X"46",
		X"02",X"00",X"3E",X"23",X"00",X"00",X"EE",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"C8",X"FF",X"00",X"00",X"FC",X"1F",X"11",X"80",X"FE",X"03",X"23",
		X"C0",X"7F",X"03",X"23",X"E8",X"7F",X"0F",X"0F",X"E0",X"FE",X"3F",X"0F",X"80",X"FB",X"0F",X"18",
		X"C0",X"7F",X"8F",X"00",X"E0",X"3D",X"E7",X"00",X"80",X"3F",X"FD",X"00",X"C8",X"FD",X"77",X"00",
		X"E0",X"F6",X"31",X"00",X"0C",X"07",X"02",X"00",X"00",X"00",X"0F",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"C8",X"FF",X"00",X"00",X"FC",X"1F",X"11",X"80",X"FE",X"03",X"23",
		X"C0",X"7F",X"03",X"23",X"E8",X"7F",X"0F",X"23",X"E0",X"FE",X"FF",X"33",X"80",X"FB",X"FB",X"10",
		X"C0",X"F0",X"FE",X"00",X"E0",X"3E",X"0F",X"07",X"80",X"3F",X"0F",X"0F",X"C8",X"FD",X"77",X"0C",
		X"E0",X"F6",X"31",X"08",X"08",X"00",X"0F",X"01",X"0C",X"07",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"08",X"8F",X"FF",X"00",X"08",X"ED",X"1F",X"11",X"08",X"EF",X"03",X"33",
		X"C0",X"4F",X"03",X"23",X"E8",X"4F",X"0F",X"23",X"E0",X"8F",X"FF",X"33",X"80",X"9F",X"FB",X"10",
		X"C0",X"1F",X"FE",X"00",X"E0",X"3E",X"F7",X"00",X"80",X"3F",X"FD",X"00",X"C8",X"FD",X"77",X"00",
		X"E0",X"F6",X"31",X"00",X"0C",X"07",X"02",X"00",X"00",X"00",X"0F",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"02",X"70",X"0E",X"03",X"0E",X"F0",X"D2",X"16",
		X"02",X"F0",X"E1",X"34",X"02",X"F0",X"F0",X"34",X"02",X"F6",X"F0",X"34",X"00",X"F6",X"3C",X"25",
		X"08",X"F6",X"30",X"25",X"08",X"F6",X"30",X"25",X"08",X"F6",X"E1",X"34",X"08",X"66",X"E1",X"16",
		X"08",X"66",X"C3",X"03",X"00",X"66",X"0E",X"01",X"00",X"EE",X"00",X"00",X"00",X"AA",X"11",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"08",X"E0",X"0E",X"03",X"08",X"F0",X"D2",X"16",
		X"08",X"F0",X"E1",X"34",X"08",X"F0",X"F0",X"34",X"08",X"F6",X"F0",X"34",X"00",X"F6",X"3C",X"25",
		X"02",X"F6",X"30",X"25",X"0E",X"F6",X"30",X"25",X"02",X"F6",X"E1",X"34",X"02",X"66",X"E1",X"16",
		X"02",X"66",X"C3",X"03",X"00",X"66",X"0E",X"01",X"00",X"EE",X"00",X"00",X"00",X"AA",X"11",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"02",X"F0",X"00",X"00",X"0E",X"F0",X"1E",X"00",
		X"02",X"F0",X"69",X"03",X"02",X"F0",X"F0",X"12",X"02",X"F6",X"F0",X"16",X"00",X"F6",X"F0",X"34",
		X"08",X"F6",X"3C",X"25",X"08",X"F6",X"34",X"24",X"08",X"F6",X"34",X"24",X"08",X"E6",X"E1",X"34",
		X"08",X"66",X"C3",X"16",X"00",X"66",X"0E",X"03",X"00",X"EE",X"00",X"00",X"00",X"AA",X"11",X"00",
		X"80",X"10",X"00",X"00",X"84",X"16",X"00",X"00",X"84",X"2D",X"00",X"00",X"84",X"78",X"00",X"00",
		X"84",X"78",X"00",X"00",X"8C",X"79",X"00",X"00",X"8C",X"79",X"00",X"00",X"88",X"5B",X"00",X"00",
		X"88",X"5B",X"00",X"00",X"8C",X"5B",X"00",X"00",X"8C",X"59",X"00",X"00",X"8C",X"59",X"00",X"00",
		X"8C",X"79",X"00",X"00",X"8C",X"79",X"00",X"00",X"8C",X"3D",X"00",X"00",X"88",X"07",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"20",X"00",X"00",X"42",X"20",X"00",
		X"00",X"03",X"30",X"00",X"80",X"90",X"16",X"00",X"C0",X"C0",X"0F",X"00",X"0C",X"C0",X"0F",X"01",
		X"08",X"90",X"0F",X"00",X"80",X"B0",X"16",X"00",X"00",X"30",X"30",X"00",X"00",X"43",X"30",X"00",
		X"00",X"42",X"20",X"00",X"00",X"E0",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"00",
		X"00",X"CC",X"77",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"CC",X"00",X"88",X"55",X"44",X"00",
		X"44",X"77",X"00",X"00",X"CC",X"DD",X"00",X"00",X"CC",X"FF",X"00",X"00",X"44",X"BB",X"00",X"00",
		X"88",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"0F",X"03",X"00",X"08",X"0F",X"01",X"00",X"80",X"0F",X"00",X"00",X"C0",X"1E",X"00",X"00",
		X"C0",X"3E",X"00",X"00",X"80",X"4F",X"00",X"00",X"40",X"CF",X"01",X"00",X"E0",X"3F",X"03",X"00",
		X"E0",X"0E",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
