library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_PGM_0 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_PGM_0 is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"AF",X"32",X"01",X"70",X"C3",X"59",X"1A",X"FF",X"3A",X"07",X"40",X"0F",X"D0",X"33",X"33",X"C9",
		X"77",X"23",X"10",X"FC",X"C9",X"FF",X"FF",X"21",X"77",X"23",X"10",X"FC",X"0D",X"20",X"F9",X"C9",
		X"85",X"6F",X"3E",X"00",X"8C",X"67",X"7E",X"C9",X"87",X"E1",X"5F",X"16",X"00",X"19",X"5E",X"23",
		X"56",X"EB",X"E9",X"FF",X"FF",X"FF",X"FF",X"FF",X"AF",X"32",X"01",X"70",X"C3",X"00",X"00",X"F5",
		X"E5",X"D5",X"C5",X"DD",X"E5",X"3A",X"0D",X"40",X"4F",X"06",X"00",X"21",X"C0",X"43",X"09",X"7E",
		X"FE",X"08",X"D2",X"49",X"03",X"3E",X"08",X"96",X"47",X"DD",X"21",X"80",X"43",X"11",X"E0",X"FF",
		X"C3",X"41",X"03",X"C3",X"8E",X"16",X"F5",X"C5",X"D5",X"E5",X"DD",X"E5",X"FD",X"E5",X"AF",X"32",
		X"01",X"70",X"3A",X"1A",X"40",X"A7",X"C2",X"D1",X"1B",X"21",X"20",X"40",X"11",X"00",X"58",X"01",
		X"80",X"00",X"ED",X"B0",X"3A",X"00",X"78",X"3A",X"15",X"40",X"32",X"16",X"40",X"3A",X"13",X"40",
		X"32",X"15",X"40",X"2A",X"10",X"40",X"22",X"13",X"40",X"3A",X"00",X"70",X"32",X"12",X"40",X"3A",
		X"00",X"68",X"32",X"11",X"40",X"3A",X"00",X"60",X"32",X"10",X"40",X"CB",X"77",X"C2",X"00",X"00",
		X"21",X"5F",X"42",X"35",X"CD",X"F3",X"18",X"CD",X"35",X"19",X"CD",X"80",X"19",X"CD",X"F9",X"16",
		X"CD",X"9C",X"18",X"CD",X"C4",X"18",X"21",X"D8",X"00",X"E5",X"3A",X"05",X"40",X"EF",X"E6",X"00",
		X"56",X"01",X"F2",X"03",X"36",X"05",X"7B",X"07",X"FD",X"E1",X"DD",X"E1",X"E1",X"D1",X"C1",X"3E",
		X"01",X"32",X"01",X"70",X"F1",X"C9",X"2A",X"0B",X"40",X"06",X"20",X"3E",X"10",X"D7",X"22",X"0B",
		X"40",X"21",X"08",X"40",X"35",X"C0",X"2D",X"36",X"01",X"2D",X"36",X"00",X"2D",X"36",X"01",X"AF",
		X"32",X"0A",X"40",X"3A",X"11",X"40",X"07",X"07",X"E6",X"03",X"32",X"00",X"40",X"3A",X"12",X"40",
		X"E6",X"04",X"0F",X"0F",X"32",X"1F",X"40",X"11",X"1B",X"05",X"CD",X"46",X"06",X"3A",X"10",X"40",
		X"E6",X"20",X"07",X"07",X"07",X"32",X"0F",X"40",X"3A",X"00",X"70",X"E6",X"03",X"21",X"52",X"01",
		X"E7",X"32",X"AC",X"40",X"CD",X"95",X"05",X"3E",X"01",X"32",X"40",X"53",X"3E",X"25",X"32",X"20",
		X"53",X"3E",X"20",X"32",X"00",X"53",X"11",X"04",X"06",X"CD",X"F2",X"08",X"11",X"03",X"05",X"C3",
		X"F2",X"08",X"FF",X"40",X"50",X"70",X"CD",X"0D",X"09",X"CD",X"8E",X"09",X"21",X"D7",X"03",X"E5",
		X"3A",X"0A",X"40",X"EF",X"8C",X"01",X"BE",X"01",X"C6",X"01",X"E1",X"01",X"18",X"02",X"3F",X"02",
		X"67",X"02",X"8E",X"02",X"C6",X"01",X"9D",X"02",X"D1",X"02",X"2E",X"03",X"E8",X"02",X"FD",X"02",
		X"14",X"06",X"61",X"06",X"D8",X"06",X"2E",X"03",X"22",X"03",X"00",X"00",X"11",X"01",X"07",X"CD",
		X"F2",X"08",X"11",X"00",X"06",X"CD",X"F2",X"08",X"3E",X"01",X"32",X"07",X"40",X"32",X"04",X"70",
		X"32",X"02",X"70",X"32",X"03",X"70",X"21",X"0A",X"40",X"34",X"AF",X"32",X"19",X"40",X"32",X"0D",
		X"40",X"32",X"0E",X"40",X"32",X"06",X"40",X"21",X"05",X"01",X"22",X"08",X"40",X"C9",X"3E",X"01",
		X"32",X"19",X"40",X"C3",X"36",X"03",X"21",X"00",X"41",X"06",X"80",X"AF",X"D7",X"32",X"5F",X"42",
		X"32",X"24",X"42",X"21",X"02",X"50",X"22",X"0B",X"40",X"21",X"09",X"40",X"36",X"20",X"2C",X"34",
		X"C9",X"2A",X"0B",X"40",X"06",X"1C",X"3E",X"10",X"D7",X"11",X"04",X"00",X"19",X"22",X"0B",X"40",
		X"21",X"09",X"40",X"35",X"C0",X"2C",X"34",X"21",X"40",X"04",X"22",X"08",X"40",X"AF",X"06",X"30",
		X"21",X"00",X"42",X"D7",X"32",X"06",X"70",X"32",X"07",X"70",X"32",X"18",X"40",X"3E",X"01",X"CD",
		X"A1",X"27",X"21",X"B5",X"1D",X"C3",X"98",X"05",X"C3",X"20",X"29",X"21",X"08",X"40",X"35",X"C0",
		X"36",X"50",X"2C",X"16",X"06",X"7E",X"82",X"5F",X"CD",X"F2",X"08",X"35",X"C0",X"2C",X"34",X"CD",
		X"3A",X"29",X"22",X"08",X"40",X"21",X"A0",X"42",X"AF",X"47",X"D7",X"C3",X"3B",X"39",X"C9",X"CD",
		X"63",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"CD",X"67",X"03",X"21",X"08",X"40",X"35",X"C0",
		X"36",X"D2",X"2C",X"CD",X"62",X"39",X"EB",X"21",X"41",X"42",X"34",X"EB",X"35",X"C0",X"36",X"D2",
		X"2C",X"34",X"AF",X"32",X"58",X"40",X"C9",X"CD",X"63",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CD",X"67",X"03",X"21",X"09",X"40",X"35",X"C0",X"2C",X"34",X"AF",X"32",X"58",X"40",X"21",X"40",
		X"11",X"22",X"08",X"40",X"21",X"41",X"42",X"34",X"11",X"11",X"06",X"C3",X"F2",X"08",X"CD",X"63",
		X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"CD",X"67",X"03",X"C3",X"E0",X"1F",X"CD",X"63",X"03",
		X"2A",X"0B",X"40",X"06",X"1C",X"3E",X"10",X"D7",X"11",X"04",X"00",X"19",X"22",X"0B",X"40",X"21",
		X"09",X"40",X"35",X"C0",X"2C",X"34",X"21",X"A0",X"42",X"AF",X"47",X"D7",X"21",X"60",X"40",X"06",
		X"40",X"D7",X"21",X"40",X"04",X"22",X"08",X"40",X"CD",X"95",X"05",X"11",X"00",X"06",X"C3",X"F2",
		X"08",X"11",X"01",X"07",X"CD",X"F2",X"08",X"11",X"00",X"06",X"CD",X"F2",X"08",X"21",X"0A",X"40",
		X"34",X"21",X"60",X"10",X"22",X"08",X"40",X"C9",X"21",X"00",X"41",X"06",X"80",X"AF",X"D7",X"32",
		X"5F",X"42",X"32",X"38",X"42",X"21",X"09",X"40",X"36",X"40",X"C3",X"93",X"05",X"11",X"1B",X"05",
		X"CD",X"46",X"06",X"EB",X"11",X"18",X"42",X"01",X"08",X"00",X"ED",X"B0",X"AF",X"32",X"5F",X"42",
		X"3C",X"32",X"1D",X"42",X"21",X"0A",X"40",X"34",X"2C",X"36",X"96",X"21",X"40",X"06",X"22",X"45",
		X"42",X"C9",X"3E",X"01",X"32",X"0A",X"40",X"21",X"03",X"03",X"22",X"08",X"40",X"C9",X"21",X"09",
		X"40",X"35",X"C0",X"2C",X"34",X"C9",X"21",X"08",X"40",X"35",X"C0",X"36",X"3C",X"2C",X"C3",X"31",
		X"03",X"DD",X"36",X"18",X"01",X"DD",X"19",X"10",X"F8",X"DD",X"E1",X"C1",X"D1",X"E1",X"F1",X"CA",
		X"E8",X"2D",X"DD",X"36",X"18",X"01",X"DD",X"19",X"C3",X"E0",X"2D",X"3A",X"0D",X"40",X"4F",X"C3",
		X"CC",X"15",X"C9",X"AF",X"C3",X"72",X"09",X"3A",X"41",X"42",X"A7",X"C8",X"3D",X"C8",X"47",X"3A",
		X"5F",X"42",X"4F",X"E6",X"3F",X"28",X"49",X"FE",X"20",X"C0",X"79",X"07",X"07",X"E6",X"03",X"4F",
		X"87",X"81",X"5F",X"16",X"00",X"21",X"9A",X"03",X"00",X"11",X"AD",X"51",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"CD",X"AF",X"03",X"10",X"FB",X"C9",X"10",X"02",X"00",X"10",X"03",X"00",
		X"10",X"04",X"00",X"10",X"05",X"00",X"01",X"00",X"00",X"12",X"19",X"17",X"10",X"06",X"00",X"0E",
		X"03",X"7E",X"12",X"23",X"7B",X"D6",X"20",X"5F",X"0D",X"C2",X"B1",X"03",X"C6",X"63",X"5F",X"C9",
		X"21",X"AD",X"51",X"11",X"E0",X"FF",X"0E",X"03",X"3E",X"10",X"77",X"19",X"0D",X"C2",X"CA",X"03",
		X"7D",X"C6",X"63",X"6F",X"10",X"F0",X"C9",X"3A",X"02",X"40",X"A7",X"C8",X"21",X"05",X"40",X"34",
		X"2C",X"2C",X"36",X"00",X"AF",X"32",X"0A",X"40",X"32",X"C2",X"41",X"32",X"DF",X"41",X"32",X"B0",
		X"40",X"C9",X"CD",X"98",X"39",X"CD",X"8E",X"09",X"21",X"92",X"04",X"E5",X"3A",X"0A",X"40",X"EF",
		X"08",X"04",X"30",X"04",X"43",X"04",X"73",X"04",X"21",X"95",X"1D",X"CD",X"98",X"05",X"21",X"60",
		X"40",X"06",X"40",X"AF",X"D7",X"21",X"60",X"42",X"D7",X"06",X"40",X"D7",X"CD",X"CE",X"1E",X"32",
		X"B0",X"40",X"21",X"02",X"50",X"22",X"0B",X"40",X"21",X"09",X"40",X"36",X"10",X"2C",X"34",X"C9",
		X"21",X"19",X"40",X"35",X"C2",X"73",X"04",X"21",X"0A",X"40",X"34",X"21",X"00",X"41",X"06",X"80",
		X"AF",X"D7",X"C9",X"2A",X"0B",X"40",X"06",X"1C",X"3E",X"10",X"D7",X"11",X"04",X"00",X"19",X"06",
		X"1C",X"D7",X"19",X"22",X"0B",X"40",X"21",X"09",X"40",X"35",X"C0",X"CD",X"EA",X"1F",X"32",X"06",
		X"70",X"32",X"07",X"70",X"32",X"18",X"40",X"11",X"02",X"07",X"CD",X"F2",X"08",X"11",X"01",X"06",
		X"CD",X"F2",X"08",X"3A",X"5F",X"42",X"E6",X"20",X"28",X"11",X"3A",X"02",X"40",X"A7",X"C8",X"47",
		X"3E",X"01",X"32",X"00",X"60",X"05",X"C8",X"32",X"01",X"60",X"C9",X"32",X"00",X"60",X"32",X"01",
		X"60",X"C9",X"3A",X"11",X"40",X"CB",X"47",X"20",X"59",X"CB",X"4F",X"C8",X"3A",X"02",X"40",X"FE",
		X"02",X"D8",X"D6",X"02",X"32",X"02",X"40",X"21",X"1B",X"05",X"11",X"A0",X"41",X"01",X"20",X"00",
		X"ED",X"B0",X"3A",X"1F",X"40",X"0F",X"DC",X"0F",X"05",X"21",X"00",X"01",X"CD",X"3B",X"36",X"21",
		X"1B",X"05",X"11",X"80",X"41",X"01",X"20",X"00",X"ED",X"B0",X"3A",X"1F",X"40",X"0F",X"DC",X"15",
		X"05",X"AF",X"32",X"0A",X"40",X"3E",X"03",X"32",X"05",X"40",X"3E",X"01",X"32",X"06",X"40",X"32",
		X"D1",X"41",X"11",X"04",X"06",X"CD",X"F2",X"08",X"11",X"00",X"04",X"CD",X"F2",X"08",X"1C",X"C3",
		X"F2",X"08",X"3A",X"02",X"40",X"A7",X"28",X"11",X"3D",X"32",X"02",X"40",X"21",X"A0",X"41",X"06",
		X"20",X"AF",X"D7",X"21",X"00",X"00",X"C3",X"BC",X"04",X"3E",X"01",X"32",X"05",X"40",X"C9",X"3E",
		X"05",X"32",X"B5",X"41",X"C9",X"3E",X"05",X"32",X"95",X"41",X"C9",X"00",X"00",X"00",X"00",X"88",
		X"11",X"50",X"0A",X"A0",X"05",X"A0",X"05",X"50",X"0A",X"88",X"11",X"3C",X"14",X"00",X"00",X"00",
		X"03",X"00",X"0F",X"00",X"00",X"00",X"CD",X"0D",X"09",X"CD",X"8E",X"09",X"3A",X"0A",X"40",X"EF",
		X"50",X"05",X"83",X"05",X"A5",X"05",X"05",X"06",X"14",X"06",X"61",X"06",X"D8",X"06",X"3D",X"07",
		X"21",X"00",X"41",X"06",X"80",X"AF",X"32",X"00",X"60",X"CD",X"AF",X"39",X"D7",X"32",X"5F",X"42",
		X"21",X"00",X"42",X"06",X"17",X"D7",X"2C",X"06",X"18",X"D7",X"21",X"60",X"42",X"06",X"20",X"D7",
		X"3E",X"01",X"32",X"26",X"42",X"21",X"0A",X"40",X"34",X"2D",X"36",X"20",X"21",X"00",X"50",X"22",
		X"0B",X"40",X"C9",X"2A",X"0B",X"40",X"06",X"20",X"3E",X"10",X"D7",X"22",X"0B",X"40",X"21",X"09",
		X"40",X"35",X"C0",X"2C",X"34",X"21",X"75",X"1D",X"11",X"21",X"40",X"06",X"20",X"7E",X"12",X"23",
		X"1C",X"1C",X"10",X"F9",X"C9",X"11",X"80",X"41",X"CD",X"46",X"06",X"EB",X"11",X"18",X"42",X"01",
		X"08",X"00",X"ED",X"B0",X"AF",X"32",X"5F",X"42",X"32",X"20",X"42",X"32",X"06",X"70",X"32",X"07",
		X"70",X"32",X"18",X"40",X"21",X"0A",X"40",X"34",X"2D",X"36",X"96",X"21",X"80",X"06",X"22",X"45",
		X"42",X"3A",X"06",X"40",X"0F",X"D0",X"3A",X"0E",X"40",X"0F",X"38",X"20",X"11",X"00",X"05",X"CD",
		X"F2",X"08",X"1E",X"02",X"CD",X"F2",X"08",X"14",X"CD",X"F2",X"08",X"1E",X"04",X"CD",X"F2",X"08",
		X"11",X"03",X"07",X"CD",X"F2",X"08",X"11",X"00",X"07",X"C3",X"F2",X"08",X"11",X"03",X"05",X"CD",
		X"F2",X"08",X"C3",X"E2",X"05",X"21",X"09",X"40",X"35",X"C0",X"36",X"14",X"2C",X"34",X"11",X"82",
		X"06",X"C3",X"F2",X"08",X"21",X"09",X"40",X"35",X"C0",X"36",X"0A",X"2C",X"34",X"21",X"01",X"00",
		X"22",X"00",X"42",X"3E",X"80",X"32",X"02",X"42",X"21",X"CA",X"15",X"11",X"4A",X"42",X"01",X"10",
		X"00",X"ED",X"B0",X"AF",X"32",X"54",X"40",X"32",X"56",X"40",X"11",X"03",X"07",X"CD",X"F2",X"08",
		X"11",X"00",X"02",X"C3",X"F2",X"08",X"CD",X"16",X"38",X"06",X"10",X"0E",X"01",X"1A",X"A1",X"28",
		X"0B",X"36",X"01",X"23",X"CB",X"01",X"30",X"F5",X"13",X"10",X"F2",X"C9",X"36",X"00",X"C3",X"53",
		X"06",X"C3",X"08",X"36",X"CD",X"98",X"08",X"CD",X"74",X"0A",X"CD",X"AA",X"0C",X"CD",X"A5",X"0B",
		X"CD",X"32",X"0A",X"CD",X"F2",X"0A",X"CD",X"5E",X"0B",X"CD",X"0E",X"12",X"CD",X"85",X"12",X"CD",
		X"E5",X"08",X"CD",X"F3",X"13",X"CD",X"2B",X"13",X"CD",X"C8",X"13",X"CD",X"DA",X"14",X"CD",X"D4",
		X"12",X"CD",X"0E",X"13",X"CD",X"8D",X"16",X"CD",X"FC",X"14",X"CD",X"3C",X"15",X"00",X"00",X"00",
		X"CD",X"DB",X"15",X"CD",X"08",X"16",X"CD",X"1E",X"16",X"CD",X"9F",X"16",X"CD",X"6F",X"16",X"CD",
		X"92",X"19",X"3A",X"08",X"42",X"2A",X"00",X"42",X"B4",X"B5",X"0F",X"D8",X"3A",X"25",X"42",X"0F",
		X"D0",X"21",X"60",X"42",X"11",X"05",X"00",X"06",X"07",X"AF",X"B6",X"19",X"10",X"FC",X"0F",X"D8",
		X"21",X"09",X"40",X"35",X"C0",X"C3",X"E6",X"28",X"21",X"0A",X"40",X"3A",X"1D",X"42",X"A7",X"20",
		X"20",X"3A",X"B5",X"41",X"A7",X"28",X"3B",X"3A",X"0E",X"40",X"A7",X"28",X"35",X"34",X"2D",X"36",
		X"82",X"3A",X"06",X"40",X"0F",X"D0",X"11",X"02",X"06",X"CD",X"F2",X"08",X"1E",X"00",X"C3",X"F2",
		X"08",X"3A",X"B5",X"41",X"A7",X"28",X"0B",X"3A",X"0E",X"40",X"A7",X"28",X"05",X"34",X"2D",X"36",
		X"50",X"C9",X"3A",X"06",X"40",X"0F",X"30",X"05",X"36",X"04",X"C3",X"0E",X"07",X"36",X"0E",X"C3",
		X"0E",X"07",X"3A",X"06",X"40",X"0F",X"30",X"E5",X"3E",X"01",X"32",X"05",X"40",X"AF",X"32",X"06",
		X"40",X"32",X"0A",X"40",X"CD",X"B9",X"1C",X"11",X"00",X"06",X"C3",X"F2",X"08",X"21",X"09",X"40",
		X"35",X"C0",X"2C",X"AF",X"77",X"32",X"22",X"42",X"32",X"2B",X"42",X"11",X"80",X"41",X"CD",X"64",
		X"07",X"21",X"18",X"42",X"01",X"08",X"00",X"ED",X"B0",X"3E",X"01",X"32",X"0D",X"40",X"3E",X"04",
		X"32",X"05",X"40",X"C9",X"CD",X"BB",X"37",X"06",X"10",X"0E",X"01",X"AF",X"CB",X"46",X"28",X"01",
		X"B1",X"23",X"CB",X"01",X"30",X"F6",X"12",X"13",X"10",X"F1",X"C9",X"CD",X"0D",X"09",X"CD",X"8E",
		X"09",X"3A",X"0A",X"40",X"EF",X"50",X"05",X"83",X"05",X"95",X"07",X"05",X"06",X"14",X"06",X"61",
		X"06",X"E8",X"07",X"18",X"08",X"11",X"A0",X"41",X"CD",X"46",X"06",X"EB",X"11",X"18",X"42",X"01",
		X"08",X"00",X"ED",X"B0",X"AF",X"32",X"5F",X"42",X"32",X"20",X"42",X"3A",X"0F",X"40",X"A7",X"28",
		X"09",X"32",X"18",X"40",X"32",X"06",X"70",X"32",X"07",X"70",X"21",X"0A",X"40",X"34",X"2D",X"36",
		X"96",X"21",X"60",X"08",X"22",X"45",X"42",X"3A",X"06",X"40",X"0F",X"D0",X"11",X"03",X"05",X"CD",
		X"F2",X"08",X"11",X"03",X"06",X"CD",X"F2",X"08",X"1C",X"CD",X"F2",X"08",X"11",X"03",X"07",X"CD",
		X"F2",X"08",X"11",X"00",X"07",X"C3",X"F2",X"08",X"21",X"0A",X"40",X"3A",X"1D",X"42",X"A7",X"20",
		X"1B",X"3A",X"95",X"41",X"A7",X"CA",X"22",X"07",X"34",X"2D",X"36",X"82",X"3A",X"06",X"40",X"0F",
		X"D0",X"11",X"03",X"06",X"CD",X"F2",X"08",X"1E",X"00",X"C3",X"F2",X"08",X"3A",X"95",X"41",X"A7",
		X"CA",X"12",X"07",X"34",X"2D",X"36",X"50",X"C9",X"21",X"09",X"40",X"35",X"C0",X"2C",X"AF",X"77",
		X"00",X"00",X"00",X"3E",X"03",X"32",X"05",X"40",X"11",X"A0",X"41",X"CD",X"64",X"07",X"21",X"18",
		X"42",X"01",X"08",X"00",X"C3",X"90",X"38",X"21",X"00",X"42",X"CB",X"46",X"28",X"39",X"2C",X"2C",
		X"3A",X"06",X"40",X"0F",X"D2",X"92",X"08",X"3A",X"18",X"40",X"0F",X"38",X"3F",X"3A",X"10",X"40",
		X"47",X"CB",X"5F",X"28",X"06",X"7E",X"FE",X"17",X"38",X"01",X"35",X"CB",X"50",X"28",X"06",X"7E",
		X"FE",X"E9",X"30",X"01",X"34",X"7E",X"2F",X"C6",X"80",X"0E",X"06",X"21",X"50",X"40",X"06",X"04",
		X"77",X"2C",X"71",X"2C",X"10",X"FA",X"C9",X"2C",X"CB",X"46",X"20",X"06",X"2C",X"36",X"00",X"C3",
		X"65",X"08",X"2C",X"7E",X"2F",X"C6",X"80",X"0E",X"07",X"C3",X"6B",X"08",X"3A",X"11",X"40",X"C3",
		X"50",X"08",X"3A",X"3F",X"42",X"C3",X"50",X"08",X"CD",X"BC",X"08",X"2A",X"09",X"42",X"3A",X"18",
		X"40",X"0F",X"38",X"0D",X"7D",X"2F",X"C6",X"FC",X"32",X"9F",X"40",X"7C",X"2F",X"32",X"9D",X"40",
		X"C9",X"7D",X"3D",X"32",X"9F",X"40",X"7C",X"2F",X"32",X"9D",X"40",X"C9",X"21",X"08",X"42",X"CB",
		X"46",X"23",X"28",X"0F",X"7E",X"D6",X"06",X"77",X"D6",X"0E",X"D6",X"0C",X"D0",X"3E",X"01",X"32",
		X"0B",X"42",X"C9",X"36",X"CC",X"2C",X"3A",X"00",X"42",X"CB",X"47",X"28",X"05",X"3A",X"02",X"42",
		X"77",X"C9",X"36",X"00",X"C9",X"C3",X"D5",X"28",X"0F",X"D0",X"AF",X"32",X"0B",X"42",X"32",X"08",
		X"42",X"C9",X"E5",X"26",X"40",X"3A",X"A0",X"40",X"6F",X"CB",X"7E",X"28",X"0E",X"72",X"2C",X"73",
		X"2C",X"7D",X"FE",X"C0",X"30",X"02",X"3E",X"C0",X"32",X"A0",X"40",X"E1",X"C9",X"21",X"08",X"42",
		X"CB",X"46",X"28",X"2A",X"2C",X"7E",X"D6",X"22",X"FE",X"50",X"30",X"22",X"2C",X"3A",X"0E",X"42",
		X"96",X"ED",X"44",X"47",X"C6",X"02",X"E6",X"0F",X"FE",X"03",X"30",X"12",X"78",X"0F",X"0F",X"0F",
		X"0F",X"E6",X"0F",X"5F",X"16",X"00",X"21",X"F0",X"41",X"19",X"CB",X"46",X"20",X"4A",X"2A",X"0E",
		X"42",X"ED",X"5B",X"10",X"42",X"3A",X"0D",X"42",X"A7",X"20",X"12",X"CB",X"7C",X"20",X"04",X"7D",
		X"BB",X"30",X"2A",X"3A",X"5F",X"42",X"E6",X"03",X"C0",X"23",X"C3",X"6C",X"09",X"CB",X"7C",X"28",
		X"04",X"7D",X"BA",X"38",X"1E",X"3A",X"5F",X"42",X"E6",X"03",X"C0",X"2B",X"22",X"0E",X"42",X"7D",
		X"ED",X"44",X"21",X"28",X"40",X"06",X"09",X"77",X"2C",X"2C",X"10",X"FB",X"C9",X"3E",X"01",X"32",
		X"0D",X"42",X"C9",X"AF",X"32",X"0D",X"42",X"C9",X"2A",X"0E",X"42",X"C3",X"6F",X"09",X"AF",X"11",
		X"E8",X"41",X"12",X"1C",X"12",X"1C",X"0E",X"06",X"21",X"23",X"41",X"06",X"0A",X"AF",X"B6",X"2C",
		X"10",X"FC",X"12",X"1C",X"7D",X"C6",X"06",X"6F",X"0D",X"C2",X"9B",X"09",X"AF",X"12",X"1C",X"12",
		X"1C",X"12",X"1C",X"21",X"23",X"41",X"0E",X"0A",X"D5",X"11",X"10",X"00",X"06",X"06",X"AF",X"B6",
		X"19",X"10",X"FC",X"D1",X"12",X"1C",X"7D",X"D6",X"5F",X"6F",X"0D",X"C2",X"B8",X"09",X"21",X"FC",
		X"41",X"06",X"0A",X"1E",X"22",X"CB",X"46",X"20",X"09",X"2D",X"7B",X"C6",X"10",X"5F",X"10",X"F5",
		X"1E",X"22",X"21",X"F3",X"41",X"06",X"0A",X"16",X"E0",X"CB",X"46",X"20",X"09",X"2C",X"7A",X"D6",
		X"10",X"57",X"10",X"F5",X"16",X"E0",X"ED",X"53",X"10",X"42",X"21",X"EA",X"41",X"0E",X"01",X"06",
		X"04",X"AF",X"B6",X"2C",X"10",X"FC",X"A9",X"32",X"21",X"42",X"A9",X"B6",X"2C",X"B6",X"A9",X"32",
		X"20",X"42",X"21",X"C0",X"42",X"11",X"20",X"00",X"06",X"07",X"AF",X"B6",X"19",X"10",X"FC",X"A9",
		X"32",X"26",X"42",X"A9",X"21",X"A1",X"42",X"06",X"08",X"B6",X"19",X"10",X"FC",X"A9",X"32",X"25",
		X"42",X"C9",X"3A",X"00",X"42",X"0F",X"D0",X"3A",X"08",X"42",X"0F",X"D8",X"3A",X"06",X"40",X"0F",
		X"30",X"26",X"3A",X"18",X"40",X"0F",X"38",X"15",X"3A",X"13",X"40",X"2F",X"47",X"3A",X"10",X"40",
		X"A0",X"E6",X"10",X"C8",X"3E",X"01",X"32",X"08",X"42",X"32",X"CC",X"41",X"C9",X"3A",X"14",X"40",
		X"2F",X"47",X"3A",X"11",X"40",X"C3",X"50",X"0A",X"3A",X"5F",X"42",X"E6",X"1F",X"C0",X"3E",X"01",
		X"32",X"08",X"42",X"C9",X"DD",X"21",X"60",X"42",X"FD",X"21",X"81",X"40",X"06",X"07",X"DD",X"CB",
		X"00",X"46",X"28",X"27",X"DD",X"7E",X"01",X"C6",X"02",X"DD",X"77",X"01",X"C6",X"04",X"38",X"1B",
		X"DD",X"6E",X"02",X"DD",X"66",X"03",X"DD",X"5E",X"04",X"CB",X"13",X"9F",X"57",X"19",X"DD",X"75",
		X"02",X"DD",X"74",X"03",X"7C",X"C6",X"10",X"FE",X"20",X"30",X"0A",X"AF",X"DD",X"77",X"00",X"DD",
		X"77",X"01",X"DD",X"77",X"03",X"3A",X"18",X"40",X"0F",X"38",X"21",X"DD",X"7E",X"01",X"2F",X"3D",
		X"FD",X"77",X"02",X"DD",X"7E",X"03",X"2F",X"4F",X"78",X"FE",X"05",X"38",X"01",X"0C",X"FD",X"71",
		X"00",X"11",X"05",X"00",X"DD",X"19",X"1D",X"FD",X"19",X"10",X"A3",X"C9",X"DD",X"7E",X"01",X"D6",
		X"04",X"FD",X"77",X"02",X"DD",X"7E",X"03",X"2F",X"4F",X"78",X"FE",X"05",X"38",X"E0",X"0D",X"C3",
		X"CE",X"0A",X"21",X"08",X"42",X"CB",X"46",X"C8",X"23",X"7E",X"FE",X"68",X"D0",X"D6",X"1E",X"D8",
		X"06",X"06",X"D6",X"04",X"D8",X"D6",X"08",X"38",X"03",X"10",X"F7",X"C9",X"23",X"3A",X"0E",X"42",
		X"96",X"ED",X"44",X"4F",X"E6",X"0F",X"D6",X"02",X"FE",X"0B",X"D0",X"04",X"79",X"E6",X"F0",X"80",
		X"0F",X"0F",X"0F",X"0F",X"5F",X"16",X"00",X"21",X"00",X"41",X"19",X"CB",X"46",X"C8",X"72",X"16",
		X"01",X"5D",X"CD",X"F2",X"08",X"7A",X"32",X"0B",X"42",X"32",X"A1",X"42",X"AF",X"32",X"A2",X"42",
		X"2A",X"09",X"42",X"22",X"A3",X"42",X"16",X"03",X"7B",X"FE",X"50",X"18",X"0C",X"E6",X"70",X"0F",
		X"0F",X"0F",X"0F",X"D6",X"04",X"5F",X"C3",X"F2",X"08",X"1E",X"00",X"C3",X"F2",X"08",X"3A",X"00",
		X"42",X"0F",X"D0",X"DD",X"21",X"60",X"42",X"11",X"05",X"00",X"06",X"07",X"CD",X"74",X"0B",X"DD",
		X"19",X"10",X"F9",X"C9",X"DD",X"CB",X"00",X"46",X"C8",X"DD",X"7E",X"01",X"C6",X"2F",X"93",X"38",
		X"10",X"D6",X"09",X"D0",X"3A",X"02",X"42",X"DD",X"96",X"03",X"83",X"FE",X"0B",X"D0",X"C3",X"9B",
		X"0B",X"3A",X"02",X"42",X"DD",X"96",X"03",X"C6",X"02",X"BB",X"D0",X"DD",X"36",X"00",X"00",X"3E",
		X"01",X"32",X"04",X"42",X"C9",X"3A",X"18",X"40",X"0F",X"38",X"2E",X"DD",X"21",X"A0",X"42",X"FD",
		X"21",X"60",X"40",X"06",X"03",X"0E",X"07",X"CD",X"07",X"0C",X"11",X"20",X"00",X"DD",X"19",X"11",
		X"04",X"00",X"FD",X"19",X"10",X"F1",X"06",X"05",X"0C",X"CD",X"07",X"0C",X"11",X"20",X"00",X"DD",
		X"19",X"11",X"04",X"00",X"FD",X"19",X"10",X"F1",X"C9",X"DD",X"21",X"A0",X"42",X"FD",X"21",X"60",
		X"40",X"06",X"03",X"0E",X"09",X"CD",X"07",X"0C",X"11",X"20",X"00",X"DD",X"19",X"11",X"04",X"00",
		X"FD",X"19",X"10",X"F1",X"06",X"05",X"0D",X"CD",X"07",X"0C",X"11",X"20",X"00",X"DD",X"19",X"11",
		X"04",X"00",X"FD",X"19",X"10",X"F1",X"C9",X"DD",X"CB",X"00",X"46",X"CA",X"7F",X"0C",X"DD",X"7E",
		X"16",X"FD",X"77",X"02",X"DD",X"7E",X"03",X"D6",X"08",X"FD",X"77",X"03",X"DD",X"7E",X"04",X"2F",
		X"91",X"FD",X"77",X"00",X"DD",X"7E",X"05",X"A7",X"F2",X"3F",X"0C",X"FE",X"FA",X"FA",X"69",X"0C",
		X"2F",X"C6",X"12",X"F6",X"40",X"DD",X"86",X"0F",X"FD",X"77",X"01",X"FD",X"34",X"03",X"C9",X"FE",
		X"06",X"F2",X"55",X"0C",X"C6",X"11",X"F6",X"C0",X"DD",X"86",X"0F",X"FD",X"77",X"01",X"FD",X"34",
		X"03",X"FD",X"34",X"00",X"C9",X"FE",X"0C",X"F2",X"77",X"0C",X"2F",X"C6",X"1E",X"F6",X"80",X"DD",
		X"86",X"0F",X"FD",X"77",X"01",X"FD",X"34",X"00",X"C9",X"FE",X"F4",X"FA",X"7B",X"0C",X"C6",X"1D",
		X"DD",X"86",X"0F",X"FD",X"77",X"01",X"C9",X"D6",X"18",X"18",X"AC",X"C6",X"18",X"18",X"A8",X"DD",
		X"CB",X"01",X"46",X"CA",X"A1",X"0C",X"FD",X"36",X"02",X"07",X"DD",X"7E",X"03",X"D6",X"08",X"FD",
		X"77",X"03",X"DD",X"7E",X"04",X"2F",X"91",X"FD",X"77",X"00",X"DD",X"7E",X"12",X"FD",X"77",X"01",
		X"C9",X"FD",X"36",X"03",X"F8",X"FD",X"36",X"00",X"F8",X"C9",X"DD",X"21",X"A0",X"42",X"11",X"20",
		X"00",X"06",X"08",X"D9",X"CD",X"BD",X"0C",X"D9",X"DD",X"19",X"10",X"F7",X"C9",X"DD",X"CB",X"01",
		X"46",X"C2",X"CB",X"10",X"DD",X"CB",X"00",X"46",X"C8",X"DD",X"7E",X"02",X"EF",X"ED",X"0C",X"58",
		X"0D",X"B8",X"0D",X"12",X"0E",X"52",X"0E",X"80",X"0E",X"EE",X"0E",X"23",X"0F",X"4D",X"0F",X"96",
		X"0F",X"06",X"10",X"75",X"10",X"78",X"10",X"82",X"10",X"A9",X"10",X"BF",X"10",X"DD",X"36",X"17",
		X"00",X"3E",X"01",X"32",X"C2",X"41",X"CD",X"2E",X"11",X"DD",X"5E",X"07",X"16",X"01",X"CD",X"F2",
		X"08",X"7B",X"E6",X"70",X"21",X"D5",X"1D",X"0F",X"0F",X"0F",X"5F",X"16",X"00",X"19",X"7E",X"DD",
		X"77",X"16",X"23",X"7E",X"DD",X"77",X"18",X"7B",X"FE",X"0E",X"00",X"00",X"DD",X"36",X"0F",X"00",
		X"DD",X"36",X"10",X"03",X"DD",X"36",X"11",X"0C",X"DD",X"36",X"13",X"00",X"DD",X"34",X"02",X"DD",
		X"CB",X"06",X"46",X"20",X"05",X"DD",X"36",X"05",X"0C",X"C9",X"DD",X"36",X"05",X"F4",X"C9",X"DD",
		X"36",X"0F",X"18",X"AF",X"DD",X"CB",X"20",X"46",X"28",X"01",X"3C",X"DD",X"CB",X"40",X"46",X"28",
		X"01",X"3C",X"32",X"2A",X"42",X"C3",X"20",X"0D",X"DD",X"6E",X"13",X"26",X"1E",X"DD",X"7E",X"03",
		X"00",X"DD",X"77",X"03",X"2C",X"DD",X"CB",X"06",X"46",X"20",X"24",X"DD",X"7E",X"04",X"00",X"DD",
		X"77",X"04",X"C6",X"07",X"FE",X"0E",X"38",X"3B",X"2C",X"DD",X"75",X"13",X"DD",X"35",X"10",X"C0",
		X"DD",X"36",X"10",X"04",X"DD",X"35",X"05",X"DD",X"35",X"11",X"C0",X"DD",X"34",X"02",X"C9",X"DD",
		X"7E",X"04",X"00",X"DD",X"77",X"04",X"C6",X"07",X"FE",X"0E",X"38",X"17",X"2C",X"DD",X"75",X"13",
		X"DD",X"35",X"10",X"C0",X"DD",X"36",X"10",X"04",X"DD",X"34",X"05",X"DD",X"35",X"11",X"C0",X"DD",
		X"34",X"02",X"C9",X"DD",X"36",X"02",X"05",X"C9",X"DD",X"34",X"03",X"DD",X"7E",X"07",X"E6",X"70",
		X"FE",X"60",X"28",X"43",X"3A",X"02",X"42",X"47",X"DD",X"7E",X"04",X"90",X"38",X"28",X"1F",X"C6",
		X"10",X"FE",X"30",X"30",X"02",X"3E",X"30",X"FE",X"70",X"38",X"02",X"3E",X"70",X"DD",X"77",X"19",
		X"DD",X"96",X"04",X"ED",X"44",X"DD",X"77",X"09",X"AF",X"DD",X"77",X"1A",X"DD",X"77",X"1B",X"DD",
		X"77",X"1C",X"DD",X"34",X"02",X"C9",X"1F",X"D6",X"10",X"FE",X"D0",X"38",X"02",X"3E",X"D0",X"FE",
		X"90",X"30",X"DA",X"3E",X"90",X"18",X"D6",X"3A",X"C0",X"42",X"0F",X"30",X"B7",X"3A",X"D9",X"42",
		X"18",X"CB",X"DD",X"34",X"03",X"CD",X"52",X"11",X"DD",X"7E",X"09",X"DD",X"86",X"19",X"DD",X"77",
		X"04",X"C6",X"07",X"FE",X"0E",X"38",X"24",X"DD",X"7E",X"03",X"C6",X"48",X"38",X"20",X"3A",X"00",
		X"42",X"0F",X"D0",X"CD",X"97",X"11",X"3A",X"2B",X"42",X"0F",X"D8",X"2A",X"13",X"42",X"DD",X"7E",
		X"03",X"BC",X"CA",X"C7",X"11",X"C6",X"19",X"2D",X"20",X"F7",X"C9",X"DD",X"34",X"02",X"DD",X"34",
		X"02",X"C9",X"3A",X"5F",X"42",X"E6",X"01",X"3C",X"DD",X"86",X"03",X"DD",X"77",X"03",X"D6",X"06",
		X"FE",X"03",X"38",X"18",X"CD",X"52",X"11",X"DD",X"7E",X"19",X"A7",X"FA",X"77",X"0E",X"DD",X"86",
		X"09",X"38",X"09",X"DD",X"77",X"04",X"C9",X"DD",X"86",X"09",X"38",X"F7",X"DD",X"34",X"02",X"C9",
		X"DD",X"36",X"03",X"08",X"DD",X"34",X"17",X"DD",X"36",X"05",X"00",X"DD",X"7E",X"07",X"E6",X"70",
		X"FE",X"70",X"28",X"2D",X"3A",X"00",X"42",X"0F",X"30",X"23",X"3A",X"24",X"42",X"A7",X"20",X"06",
		X"3A",X"21",X"42",X"A7",X"28",X"17",X"DD",X"7E",X"04",X"1F",X"4F",X"CD",X"DC",X"16",X"E6",X"1F",
		X"81",X"C6",X"20",X"DD",X"77",X"04",X"DD",X"36",X"10",X"28",X"DD",X"34",X"02",X"DD",X"34",X"02",
		X"C9",X"3A",X"2A",X"42",X"A7",X"20",X"12",X"DD",X"36",X"00",X"00",X"3A",X"1E",X"42",X"3C",X"FE",
		X"03",X"38",X"02",X"3E",X"02",X"32",X"1E",X"42",X"C9",X"AF",X"DD",X"CB",X"20",X"46",X"28",X"01",
		X"3C",X"DD",X"CB",X"40",X"46",X"28",X"01",X"3C",X"32",X"2A",X"42",X"C3",X"94",X"0E",X"DD",X"46",
		X"03",X"04",X"CD",X"2E",X"11",X"DD",X"7E",X"03",X"DD",X"70",X"03",X"90",X"28",X"14",X"FE",X"19",
		X"D0",X"E6",X"01",X"C0",X"DD",X"CB",X"06",X"46",X"20",X"04",X"DD",X"34",X"05",X"C9",X"DD",X"35",
		X"05",X"C9",X"DD",X"36",X"00",X"00",X"26",X"41",X"DD",X"6E",X"07",X"16",X"00",X"36",X"01",X"5D",
		X"C3",X"F2",X"08",X"DD",X"34",X"03",X"3A",X"02",X"42",X"DD",X"96",X"04",X"ED",X"44",X"17",X"5F",
		X"9F",X"57",X"CB",X"13",X"CB",X"12",X"DD",X"66",X"04",X"DD",X"6E",X"09",X"A7",X"ED",X"52",X"DD",
		X"74",X"04",X"DD",X"75",X"09",X"DD",X"35",X"10",X"C0",X"DD",X"34",X"02",X"C9",X"DD",X"34",X"03",
		X"DD",X"7E",X"03",X"D6",X"60",X"FE",X"40",X"30",X"09",X"DD",X"7E",X"04",X"D6",X"60",X"FE",X"40",
		X"38",X"0C",X"CD",X"C4",X"0D",X"DD",X"36",X"18",X"03",X"DD",X"36",X"10",X"64",X"C9",X"DD",X"34",
		X"02",X"DD",X"34",X"02",X"DD",X"36",X"10",X"03",X"DD",X"36",X"11",X"0C",X"DD",X"36",X"05",X"00",
		X"DD",X"36",X"13",X"00",X"3A",X"02",X"42",X"DD",X"96",X"04",X"38",X"05",X"DD",X"36",X"06",X"00",
		X"C9",X"DD",X"36",X"06",X"01",X"C9",X"DD",X"34",X"03",X"CD",X"52",X"11",X"DD",X"7E",X"17",X"FE",
		X"04",X"28",X"48",X"30",X"4D",X"DD",X"7E",X"09",X"DD",X"86",X"19",X"DD",X"77",X"04",X"C6",X"07",
		X"FE",X"0E",X"38",X"29",X"DD",X"7E",X"03",X"C6",X"40",X"38",X"27",X"DD",X"35",X"10",X"28",X"27",
		X"3A",X"00",X"42",X"0F",X"D0",X"CD",X"97",X"11",X"3A",X"2B",X"42",X"0F",X"D8",X"2A",X"13",X"42",
		X"DD",X"7E",X"03",X"BC",X"CA",X"C7",X"11",X"C6",X"19",X"2D",X"20",X"F7",X"C9",X"DD",X"36",X"02",
		X"05",X"C9",X"DD",X"36",X"02",X"04",X"C9",X"DD",X"35",X"02",X"C9",X"3A",X"5F",X"42",X"E6",X"01",
		X"28",X"B3",X"3A",X"02",X"42",X"DD",X"96",X"09",X"38",X"06",X"DD",X"34",X"09",X"C3",X"A5",X"0F",
		X"DD",X"35",X"09",X"C3",X"A5",X"0F",X"DD",X"6E",X"13",X"26",X"1E",X"DD",X"7E",X"03",X"00",X"DD",
		X"77",X"03",X"2C",X"DD",X"CB",X"06",X"46",X"20",X"2E",X"DD",X"7E",X"04",X"00",X"DD",X"77",X"04",
		X"2C",X"DD",X"75",X"13",X"DD",X"35",X"10",X"C0",X"DD",X"36",X"10",X"04",X"DD",X"35",X"05",X"DD",
		X"35",X"11",X"C0",X"DD",X"34",X"02",X"DD",X"36",X"10",X"03",X"DD",X"36",X"11",X"0C",X"DD",X"36",
		X"05",X"0C",X"DD",X"36",X"13",X"00",X"C9",X"DD",X"7E",X"04",X"00",X"DD",X"77",X"04",X"2C",X"DD",
		X"75",X"13",X"DD",X"35",X"10",X"C0",X"DD",X"36",X"10",X"04",X"DD",X"34",X"05",X"DD",X"35",X"11",
		X"C0",X"DD",X"34",X"02",X"DD",X"36",X"10",X"03",X"DD",X"36",X"11",X"0C",X"DD",X"36",X"05",X"F4",
		X"DD",X"36",X"13",X"00",X"C9",X"C3",X"58",X"0D",X"DD",X"34",X"03",X"DD",X"36",X"02",X"08",X"C3",
		X"62",X"0F",X"FD",X"CB",X"18",X"46",X"28",X"0C",X"FD",X"CB",X"08",X"46",X"20",X"06",X"C3",X"0F",
		X"1E",X"CA",X"AA",X"15",X"FD",X"19",X"10",X"EA",X"C9",X"FE",X"04",X"C2",X"3D",X"2D",X"3A",X"0D",
		X"40",X"4F",X"06",X"00",X"21",X"C0",X"43",X"09",X"34",X"C3",X"46",X"2D",X"DD",X"36",X"1F",X"00",
		X"CA",X"46",X"2D",X"C3",X"9E",X"10",X"3A",X"0D",X"40",X"4F",X"06",X"00",X"21",X"AA",X"43",X"09",
		X"7E",X"C9",X"21",X"C0",X"43",X"09",X"7E",X"A7",X"C3",X"FA",X"26",X"DD",X"7E",X"02",X"EF",X"D7",
		X"10",X"F9",X"10",X"24",X"11",X"2D",X"11",X"DD",X"36",X"10",X"04",X"DD",X"36",X"11",X"04",X"DD",
		X"36",X"12",X"1C",X"DD",X"34",X"02",X"DD",X"7E",X"07",X"FE",X"70",X"00",X"00",X"3E",X"07",X"32",
		X"DF",X"41",X"C9",X"3E",X"17",X"32",X"DF",X"41",X"C9",X"DD",X"35",X"10",X"C0",X"DD",X"36",X"10",
		X"04",X"DD",X"34",X"12",X"DD",X"35",X"11",X"C0",X"DD",X"7E",X"07",X"FE",X"70",X"00",X"00",X"DD",
		X"36",X"01",X"00",X"C9",X"DD",X"36",X"10",X"32",X"3A",X"2D",X"42",X"C6",X"20",X"DD",X"77",X"12",
		X"DD",X"34",X"02",X"C9",X"DD",X"35",X"10",X"C0",X"DD",X"36",X"01",X"00",X"C9",X"C9",X"DD",X"7E",
		X"07",X"E6",X"70",X"0F",X"4F",X"0F",X"81",X"ED",X"44",X"C6",X"7C",X"DD",X"77",X"03",X"DD",X"7E",
		X"07",X"E6",X"0F",X"07",X"07",X"07",X"07",X"C6",X"07",X"4F",X"3A",X"0E",X"42",X"81",X"DD",X"77",
		X"04",X"C9",X"DD",X"7E",X"18",X"E6",X"03",X"3C",X"47",X"DD",X"66",X"19",X"DD",X"6E",X"1A",X"DD",
		X"56",X"1B",X"DD",X"5E",X"1C",X"7D",X"4C",X"87",X"30",X"01",X"25",X"82",X"57",X"3E",X"00",X"8C",
		X"FE",X"80",X"20",X"01",X"79",X"67",X"4D",X"ED",X"44",X"87",X"30",X"01",X"2D",X"83",X"5F",X"3E",
		X"00",X"8D",X"FE",X"80",X"20",X"01",X"79",X"6F",X"10",X"DB",X"DD",X"74",X"19",X"DD",X"75",X"1A",
		X"DD",X"72",X"1B",X"DD",X"73",X"1C",X"C9",X"3E",X"F0",X"DD",X"96",X"03",X"57",X"3A",X"02",X"42",
		X"DD",X"96",X"04",X"38",X"07",X"CD",X"B7",X"11",X"DD",X"77",X"05",X"C9",X"ED",X"44",X"CD",X"B7",
		X"11",X"ED",X"44",X"DD",X"77",X"05",X"C9",X"CD",X"E8",X"16",X"79",X"A7",X"F2",X"C1",X"11",X"3E",
		X"80",X"07",X"07",X"07",X"E6",X"07",X"C9",X"11",X"05",X"00",X"21",X"60",X"42",X"06",X"07",X"CB",
		X"46",X"28",X"04",X"19",X"10",X"F9",X"C9",X"36",X"01",X"23",X"DD",X"7E",X"03",X"77",X"3E",X"F0",
		X"96",X"57",X"23",X"23",X"DD",X"7E",X"04",X"77",X"23",X"3A",X"02",X"42",X"DD",X"96",X"04",X"38",
		X"05",X"CD",X"FF",X"11",X"77",X"C9",X"ED",X"44",X"CD",X"FF",X"11",X"ED",X"44",X"77",X"C9",X"CD",
		X"E8",X"16",X"CD",X"DC",X"16",X"E6",X"1F",X"81",X"C6",X"06",X"F0",X"3E",X"7F",X"C9",X"3A",X"08",
		X"42",X"0F",X"D0",X"DD",X"21",X"C0",X"42",X"11",X"20",X"00",X"06",X"07",X"D9",X"CD",X"26",X"12",
		X"D9",X"DD",X"19",X"10",X"F7",X"C9",X"DD",X"CB",X"00",X"46",X"C8",X"2A",X"09",X"42",X"DD",X"7E",
		X"03",X"95",X"C6",X"03",X"FE",X"09",X"D0",X"DD",X"7E",X"04",X"94",X"C6",X"05",X"FE",X"0C",X"D0",
		X"3E",X"01",X"32",X"0B",X"42",X"DD",X"36",X"00",X"00",X"DD",X"36",X"01",X"01",X"DD",X"36",X"02",
		X"00",X"11",X"00",X"03",X"C3",X"F2",X"08",X"DD",X"7E",X"07",X"B9",X"DA",X"F2",X"08",X"08",X"D6",
		X"10",X"10",X"F7",X"21",X"01",X"F0",X"22",X"2B",X"42",X"3A",X"2A",X"42",X"FE",X"02",X"CC",X"79",
		X"12",X"32",X"2D",X"42",X"83",X"5F",X"C3",X"F2",X"08",X"DD",X"CB",X"20",X"46",X"C0",X"DD",X"CB",
		X"40",X"46",X"C0",X"3C",X"C9",X"3A",X"00",X"42",X"0F",X"D0",X"DD",X"21",X"C0",X"42",X"11",X"20",
		X"00",X"06",X"07",X"D9",X"CD",X"9D",X"12",X"D9",X"DD",X"19",X"10",X"F7",X"C9",X"DD",X"CB",X"00",
		X"46",X"C8",X"DD",X"7E",X"03",X"C6",X"31",X"D6",X"05",X"38",X"16",X"D6",X"0C",X"D0",X"3A",X"02",
		X"42",X"DD",X"96",X"04",X"C6",X"0A",X"FE",X"15",X"D0",X"3E",X"01",X"32",X"04",X"42",X"C3",X"45",
		X"12",X"3A",X"02",X"42",X"DD",X"96",X"04",X"C6",X"07",X"FE",X"0F",X"D0",X"3E",X"01",X"32",X"04",
		X"42",X"C3",X"45",X"12",X"21",X"04",X"42",X"CB",X"46",X"C8",X"36",X"00",X"21",X"00",X"01",X"22",
		X"00",X"42",X"21",X"09",X"04",X"22",X"05",X"42",X"11",X"05",X"02",X"CD",X"F2",X"08",X"3A",X"1A",
		X"42",X"A7",X"28",X"01",X"3D",X"32",X"1A",X"42",X"21",X"1D",X"42",X"35",X"7E",X"FE",X"06",X"38",
		X"02",X"36",X"05",X"3A",X"06",X"40",X"0F",X"D0",X"3E",X"01",X"32",X"03",X"68",X"C9",X"3A",X"01",
		X"42",X"0F",X"D0",X"21",X"05",X"42",X"35",X"C0",X"36",X"09",X"23",X"16",X"02",X"5E",X"CD",X"F2",
		X"08",X"35",X"C0",X"AF",X"32",X"01",X"42",X"CD",X"34",X"39",X"C9",X"C9",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DD",X"21",X"C0",X"42",
		X"DD",X"CB",X"00",X"46",X"C2",X"51",X"13",X"DD",X"CB",X"01",X"46",X"C2",X"51",X"13",X"C3",X"A7",
		X"14",X"C5",X"06",X"00",X"0E",X"20",X"DD",X"09",X"00",X"00",X"C1",X"3A",X"B5",X"43",X"3C",X"32",
		X"B5",X"43",X"C3",X"98",X"13",X"C3",X"40",X"13",X"36",X"41",X"27",X"41",X"28",X"41",X"39",X"41",
		X"47",X"41",X"48",X"41",X"57",X"41",X"58",X"41",X"66",X"41",X"69",X"41",X"77",X"41",X"78",X"41",
		X"23",X"41",X"34",X"41",X"45",X"41",X"2C",X"41",X"3B",X"41",X"4A",X"41",X"73",X"41",X"64",X"41",
		X"55",X"41",X"7C",X"41",X"6B",X"41",X"5A",X"41",X"FE",X"08",X"C2",X"40",X"13",X"AF",X"32",X"B5",
		X"43",X"C9",X"00",X"21",X"C9",X"41",X"7E",X"3D",X"C2",X"B5",X"13",X"77",X"21",X"20",X"00",X"22",
		X"CA",X"41",X"C3",X"D6",X"27",X"23",X"7E",X"A7",X"CA",X"D6",X"27",X"CD",X"8E",X"18",X"C3",X"16",
		X"17",X"00",X"16",X"01",X"5D",X"C3",X"F2",X"08",X"2A",X"0E",X"42",X"ED",X"5B",X"10",X"42",X"CB",
		X"7C",X"28",X"0B",X"7D",X"92",X"FE",X"1C",X"30",X"11",X"AF",X"32",X"15",X"42",X"C9",X"7B",X"95",
		X"FE",X"08",X"30",X"06",X"3E",X"01",X"32",X"15",X"42",X"C9",X"CD",X"DC",X"16",X"E6",X"01",X"32",
		X"15",X"42",X"C9",X"3A",X"20",X"42",X"0F",X"D8",X"3A",X"00",X"42",X"0F",X"D0",X"3A",X"28",X"42",
		X"0F",X"D0",X"AF",X"32",X"28",X"42",X"32",X"B1",X"43",X"32",X"B2",X"43",X"32",X"B7",X"43",X"32",
		X"B5",X"43",X"3A",X"B6",X"43",X"CB",X"47",X"C2",X"20",X"14",X"CD",X"2B",X"14",X"C3",X"23",X"14",
		X"CD",X"64",X"14",X"3A",X"B6",X"43",X"3C",X"32",X"B6",X"43",X"C9",X"3A",X"B3",X"43",X"5F",X"3A",
		X"B1",X"43",X"83",X"4F",X"06",X"00",X"21",X"68",X"13",X"09",X"09",X"5E",X"23",X"56",X"EB",X"CB",
		X"46",X"C4",X"A0",X"14",X"3A",X"B1",X"43",X"3C",X"32",X"B1",X"43",X"FE",X"04",X"CA",X"54",X"14",
		X"00",X"C3",X"2B",X"14",X"3A",X"B7",X"43",X"A7",X"00",X"00",X"00",X"3A",X"B3",X"43",X"C6",X"04",
		X"C3",X"C6",X"14",X"C9",X"3A",X"B4",X"43",X"5F",X"3A",X"B2",X"43",X"83",X"4F",X"06",X"00",X"21",
		X"80",X"13",X"09",X"09",X"5E",X"23",X"56",X"EB",X"CB",X"46",X"C4",X"A0",X"14",X"3A",X"B2",X"43",
		X"3C",X"32",X"B2",X"43",X"FE",X"03",X"CA",X"8D",X"14",X"00",X"C3",X"64",X"14",X"3A",X"B7",X"43",
		X"A7",X"00",X"00",X"00",X"3A",X"B4",X"43",X"C6",X"03",X"C3",X"D0",X"14",X"00",X"00",X"00",X"C9",
		X"3A",X"15",X"42",X"4F",X"C3",X"38",X"13",X"36",X"00",X"DD",X"36",X"00",X"01",X"DD",X"36",X"02",
		X"00",X"DD",X"71",X"06",X"DD",X"75",X"07",X"3A",X"B7",X"43",X"3C",X"00",X"32",X"B7",X"43",X"16",
		X"01",X"5D",X"C3",X"F2",X"08",X"00",X"FE",X"0C",X"C2",X"CC",X"14",X"AF",X"32",X"B3",X"43",X"C9",
		X"FE",X"0C",X"C2",X"D6",X"14",X"AF",X"32",X"B4",X"43",X"C9",X"3A",X"00",X"42",X"0F",X"D0",X"3A",
		X"2B",X"42",X"0F",X"D8",X"21",X"18",X"42",X"35",X"C0",X"36",X"3C",X"23",X"35",X"C0",X"36",X"14",
		X"23",X"7E",X"FE",X"07",X"C8",X"30",X"02",X"34",X"C9",X"36",X"07",X"C9",X"3A",X"00",X"42",X"0F",
		X"D0",X"3A",X"20",X"42",X"0F",X"D8",X"3A",X"2B",X"42",X"0F",X"D8",X"2A",X"1A",X"42",X"7C",X"FE",
		X"02",X"30",X"01",X"AF",X"85",X"E6",X"0F",X"06",X"01",X"21",X"4A",X"42",X"11",X"CA",X"15",X"35",
		X"28",X"05",X"AF",X"32",X"28",X"42",X"C9",X"0E",X"00",X"1A",X"77",X"23",X"13",X"35",X"CC",X"C6",
		X"15",X"10",X"F8",X"79",X"A7",X"C8",X"3E",X"01",X"32",X"28",X"42",X"C9",X"3A",X"00",X"42",X"0F",
		X"D0",X"3A",X"EF",X"41",X"0F",X"D0",X"3A",X"2B",X"42",X"0F",X"D8",X"3A",X"06",X"40",X"0F",X"30",
		X"3D",X"21",X"45",X"42",X"35",X"C0",X"36",X"3C",X"3A",X"21",X"42",X"0F",X"38",X"2C",X"23",X"35",
		X"C0",X"34",X"2A",X"77",X"41",X"7C",X"85",X"E6",X"03",X"4F",X"2A",X"1A",X"42",X"7C",X"85",X"C8",
		X"0F",X"0F",X"E6",X"03",X"2F",X"C6",X"0A",X"91",X"32",X"46",X"42",X"07",X"07",X"32",X"2F",X"42",
		X"07",X"32",X"4A",X"42",X"3E",X"01",X"32",X"2E",X"42",X"C9",X"3E",X"04",X"18",X"ED",X"21",X"45",
		X"42",X"35",X"C0",X"36",X"78",X"23",X"35",X"C0",X"36",X"05",X"3E",X"5A",X"32",X"2F",X"42",X"3E",
		X"2D",X"32",X"4A",X"42",X"3E",X"01",X"32",X"2E",X"42",X"C9",X"FD",X"74",X"04",X"FD",X"75",X"07",
		X"FD",X"36",X"18",X"00",X"FD",X"36",X"05",X"20",X"C3",X"C5",X"31",X"DD",X"7E",X"00",X"FE",X"04",
		X"C2",X"DA",X"36",X"C3",X"02",X"18",X"1A",X"77",X"0C",X"C9",X"03",X"2F",X"06",X"00",X"C3",X"C2",
		X"10",X"65",X"4F",X"49",X"43",X"3D",X"3B",X"35",X"2B",X"29",X"25",X"21",X"E8",X"41",X"06",X"04",
		X"3A",X"1B",X"42",X"A7",X"20",X"16",X"1E",X"01",X"16",X"84",X"CB",X"46",X"20",X"09",X"23",X"CB",
		X"46",X"20",X"04",X"23",X"1C",X"10",X"F3",X"ED",X"53",X"13",X"42",X"C9",X"1E",X"02",X"16",X"9D",
		X"18",X"E8",X"1E",X"03",X"16",X"B6",X"18",X"E2",X"3A",X"20",X"42",X"0F",X"D0",X"3A",X"25",X"42",
		X"0F",X"D0",X"3A",X"22",X"42",X"0F",X"D8",X"C3",X"6D",X"39",X"22",X"22",X"42",X"C9",X"21",X"22",
		X"42",X"CB",X"46",X"C8",X"C3",X"00",X"28",X"2B",X"36",X"00",X"11",X"1B",X"05",X"CD",X"46",X"06",
		X"AF",X"32",X"1A",X"42",X"32",X"5F",X"42",X"21",X"01",X"00",X"22",X"0E",X"42",X"2A",X"1B",X"42",
		X"24",X"7D",X"FE",X"07",X"28",X"03",X"30",X"22",X"3C",X"6F",X"22",X"1B",X"42",X"11",X"00",X"07",
		X"CD",X"F2",X"08",X"C9",X"1E",X"42",X"A7",X"C8",X"21",X"77",X"41",X"36",X"01",X"3D",X"32",X"1E",
		X"42",X"C8",X"23",X"36",X"01",X"AF",X"32",X"1E",X"42",X"C9",X"3E",X"07",X"C3",X"49",X"16",X"21",
		X"2B",X"42",X"CB",X"46",X"C8",X"3A",X"24",X"42",X"A7",X"20",X"0B",X"3A",X"21",X"42",X"A7",X"20",
		X"05",X"3A",X"26",X"42",X"0F",X"D0",X"23",X"35",X"C0",X"2B",X"36",X"00",X"C9",X"3A",X"07",X"40",
		X"0F",X"D8",X"21",X"DF",X"41",X"7E",X"A7",X"C8",X"0F",X"0F",X"00",X"00",X"00",X"35",X"C9",X"3A",
		X"07",X"40",X"0F",X"D8",X"21",X"23",X"41",X"11",X"06",X"00",X"4B",X"3E",X"01",X"06",X"0A",X"86",
		X"2C",X"10",X"FC",X"19",X"0D",X"C2",X"AD",X"16",X"21",X"00",X"68",X"06",X"03",X"3D",X"28",X"14",
		X"36",X"01",X"2C",X"10",X"F8",X"FE",X"02",X"38",X"05",X"AF",X"32",X"24",X"42",X"C9",X"3E",X"01",
		X"32",X"24",X"42",X"C9",X"36",X"00",X"2C",X"10",X"FB",X"C3",X"C5",X"16",X"3A",X"1E",X"40",X"47",
		X"87",X"87",X"80",X"3C",X"32",X"1E",X"40",X"C9",X"0E",X"00",X"06",X"08",X"BA",X"38",X"01",X"92",
		X"3F",X"CB",X"11",X"CB",X"1A",X"10",X"F5",X"C9",X"C9",X"C3",X"AC",X"27",X"00",X"3D",X"32",X"C1",
		X"41",X"CD",X"4B",X"17",X"CD",X"D4",X"17",X"CD",X"1D",X"18",X"CD",X"61",X"17",X"CD",X"53",X"18",
		X"CD",X"7A",X"18",X"CD",X"27",X"17",X"3A",X"C0",X"41",X"32",X"06",X"68",X"0F",X"32",X"07",X"68",
		X"3A",X"C1",X"41",X"32",X"00",X"78",X"C9",X"3A",X"CC",X"41",X"3D",X"C2",X"37",X"17",X"32",X"CC",
		X"41",X"3E",X"08",X"32",X"CE",X"41",X"C9",X"3A",X"CE",X"41",X"A7",X"CA",X"47",X"17",X"3D",X"32",
		X"CE",X"41",X"3A",X"07",X"40",X"EE",X"01",X"32",X"05",X"68",X"C9",X"3A",X"D1",X"41",X"3D",X"C0",
		X"32",X"D1",X"41",X"3C",X"32",X"D2",X"41",X"32",X"D6",X"41",X"21",X"68",X"1E",X"22",X"D3",X"41",
		X"C9",X"21",X"D2",X"41",X"CD",X"70",X"17",X"21",X"CF",X"41",X"CD",X"70",X"17",X"21",X"CD",X"41",
		X"7E",X"A7",X"C8",X"EB",X"3E",X"02",X"32",X"C0",X"41",X"3A",X"D5",X"41",X"32",X"C1",X"41",X"3A",
		X"D6",X"41",X"3D",X"C2",X"A6",X"17",X"2A",X"D3",X"41",X"7E",X"FE",X"E0",X"28",X"1C",X"23",X"22",
		X"D3",X"41",X"47",X"E6",X"1F",X"21",X"AD",X"17",X"E7",X"32",X"D5",X"41",X"78",X"E6",X"E0",X"07",
		X"07",X"07",X"21",X"CC",X"17",X"E7",X"32",X"D6",X"41",X"C9",X"AF",X"12",X"C9",X"FF",X"00",X"E1",
		X"55",X"5F",X"68",X"70",X"80",X"8E",X"9A",X"A0",X"AA",X"B4",X"B8",X"C0",X"C7",X"CD",X"D0",X"D5",
		X"DA",X"DC",X"E0",X"0C",X"35",X"87",X"A5",X"C4",X"D3",X"CA",X"E3",X"E6",X"01",X"02",X"04",X"08",
		X"10",X"20",X"40",X"00",X"3A",X"06",X"40",X"0F",X"D0",X"21",X"C2",X"41",X"7E",X"3D",X"C2",X"E9",
		X"17",X"77",X"21",X"02",X"A0",X"22",X"C3",X"41",X"C9",X"3A",X"26",X"42",X"0F",X"D8",X"3A",X"C4",
		X"41",X"32",X"C1",X"41",X"3C",X"32",X"C4",X"41",X"FE",X"E0",X"20",X"05",X"C6",X"80",X"32",X"C4",
		X"41",X"C9",X"DD",X"36",X"04",X"FF",X"DD",X"36",X"07",X"FF",X"DD",X"36",X"00",X"00",X"DD",X"36",
		X"18",X"01",X"C3",X"D6",X"36",X"DD",X"36",X"00",X"00",X"00",X"C3",X"33",X"2D",X"3A",X"06",X"40",
		X"0F",X"D0",X"3A",X"DF",X"41",X"FE",X"06",X"C2",X"3E",X"18",X"3A",X"CD",X"41",X"0F",X"D8",X"3E",
		X"01",X"32",X"CF",X"41",X"32",X"D6",X"41",X"21",X"BD",X"1E",X"22",X"D3",X"41",X"C9",X"FE",X"16",
		X"C0",X"C3",X"18",X"24",X"41",X"3C",X"32",X"CD",X"41",X"32",X"D6",X"41",X"21",X"DF",X"1E",X"22",
		X"D3",X"41",X"C9",X"2A",X"C7",X"41",X"CB",X"45",X"CA",X"62",X"18",X"21",X"00",X"80",X"22",X"C7",
		X"41",X"C9",X"7C",X"A7",X"C8",X"3D",X"32",X"C8",X"41",X"E6",X"04",X"CA",X"70",X"18",X"3E",X"81",
		X"3D",X"32",X"C1",X"41",X"3E",X"01",X"32",X"C0",X"41",X"C9",X"21",X"C9",X"41",X"7E",X"3D",X"C2",
		X"8A",X"18",X"77",X"21",X"20",X"00",X"22",X"CA",X"41",X"C9",X"23",X"7E",X"A7",X"C8",X"35",X"23",
		X"7E",X"C6",X"04",X"77",X"32",X"C1",X"41",X"AF",X"32",X"C0",X"41",X"C9",X"3A",X"D0",X"41",X"A7",
		X"28",X"08",X"AF",X"32",X"D0",X"41",X"3E",X"0F",X"18",X"0C",X"3A",X"5F",X"42",X"C6",X"01",X"D0",
		X"3A",X"1F",X"42",X"A7",X"C8",X"3D",X"32",X"1F",X"42",X"06",X"04",X"21",X"04",X"60",X"77",X"23",
		X"0F",X"10",X"FB",X"C9",X"3A",X"B0",X"40",X"0F",X"D0",X"2A",X"B1",X"40",X"7E",X"E6",X"07",X"20",
		X"1B",X"EB",X"2A",X"B3",X"40",X"7E",X"FE",X"3F",X"28",X"11",X"23",X"22",X"B3",X"40",X"D6",X"30",
		X"2A",X"B5",X"40",X"77",X"01",X"E0",X"FF",X"09",X"22",X"B5",X"40",X"EB",X"35",X"C0",X"AF",X"32",
		X"B0",X"40",X"C9",X"3A",X"00",X"40",X"FE",X"03",X"28",X"21",X"21",X"10",X"40",X"7E",X"2C",X"2C",
		X"2C",X"B6",X"2C",X"2C",X"2F",X"A6",X"2C",X"A6",X"CB",X"7F",X"20",X"16",X"E6",X"03",X"C8",X"21",
		X"04",X"40",X"34",X"CB",X"47",X"C8",X"E6",X"02",X"C8",X"34",X"C9",X"21",X"00",X"09",X"22",X"01",
		X"40",X"C9",X"21",X"02",X"40",X"7E",X"FE",X"63",X"D0",X"34",X"3E",X"01",X"32",X"C9",X"41",X"11",
		X"01",X"07",X"C3",X"F2",X"08",X"21",X"03",X"40",X"7E",X"A7",X"20",X"3C",X"2C",X"B6",X"C8",X"35",
		X"2D",X"36",X"0F",X"3A",X"00",X"40",X"FE",X"03",X"C8",X"3D",X"28",X"1C",X"21",X"02",X"40",X"3D",
		X"CC",X"53",X"19",X"7E",X"FE",X"63",X"C8",X"30",X"0C",X"34",X"3E",X"01",X"32",X"C9",X"41",X"11",
		X"01",X"07",X"C3",X"F2",X"08",X"36",X"63",X"C9",X"21",X"01",X"40",X"CB",X"46",X"28",X"06",X"36",
		X"00",X"2C",X"C3",X"53",X"19",X"36",X"01",X"C9",X"0F",X"0F",X"0F",X"32",X"03",X"60",X"35",X"C9",
		X"3A",X"02",X"40",X"FE",X"09",X"30",X"06",X"3E",X"00",X"00",X"00",X"00",X"C9",X"AF",X"00",X"00",
		X"00",X"C9",X"3A",X"5F",X"42",X"C6",X"09",X"E6",X"1F",X"C0",X"3A",X"07",X"40",X"0F",X"D0",X"3A",
		X"00",X"42",X"0F",X"D0",X"DD",X"21",X"C0",X"42",X"06",X"00",X"D9",X"11",X"20",X"00",X"06",X"07",
		X"D9",X"DD",X"66",X"03",X"DD",X"6E",X"04",X"DD",X"4E",X"1A",X"CD",X"16",X"1A",X"D9",X"DD",X"19",
		X"10",X"EE",X"DD",X"21",X"60",X"42",X"11",X"05",X"00",X"06",X"07",X"D9",X"DD",X"66",X"01",X"DD",
		X"6E",X"03",X"DD",X"4E",X"04",X"CD",X"16",X"1A",X"D9",X"DD",X"19",X"10",X"EE",X"D9",X"3A",X"02",
		X"42",X"4F",X"3A",X"0E",X"42",X"C6",X"80",X"91",X"CB",X"2F",X"CB",X"2F",X"CB",X"2F",X"CB",X"2F",
		X"CB",X"2F",X"80",X"CB",X"2F",X"4F",X"CD",X"DC",X"16",X"41",X"87",X"9F",X"20",X"01",X"3C",X"80",
		X"C6",X"01",X"FA",X"12",X"1A",X"FE",X"02",X"30",X"05",X"AF",X"32",X"3F",X"42",X"C9",X"3E",X"04",
		X"18",X"F8",X"3E",X"08",X"18",X"F4",X"DD",X"CB",X"00",X"46",X"C8",X"7C",X"D6",X"80",X"D8",X"1E",
		X"00",X"D6",X"34",X"38",X"04",X"1C",X"D6",X"34",X"D0",X"3A",X"02",X"42",X"95",X"D6",X"40",X"FE",
		X"80",X"D0",X"E6",X"60",X"6F",X"79",X"E6",X"80",X"B5",X"0F",X"0F",X"0F",X"0F",X"B3",X"5F",X"16",
		X"00",X"21",X"49",X"1A",X"19",X"7E",X"80",X"47",X"C9",X"02",X"03",X"FE",X"02",X"FF",X"FE",X"00",
		X"FF",X"00",X"01",X"01",X"02",X"02",X"FE",X"FE",X"03",X"21",X"00",X"50",X"06",X"04",X"3E",X"10",
		X"77",X"2C",X"C2",X"60",X"1A",X"24",X"3A",X"00",X"78",X"10",X"F3",X"21",X"00",X"58",X"AF",X"77",
		X"2C",X"C2",X"6F",X"1A",X"AF",X"21",X"00",X"60",X"06",X"04",X"77",X"23",X"10",X"FC",X"3C",X"06",
		X"04",X"77",X"23",X"10",X"FC",X"AF",X"06",X"08",X"21",X"00",X"68",X"77",X"23",X"10",X"FC",X"06",
		X"08",X"21",X"01",X"70",X"77",X"23",X"10",X"FC",X"3D",X"32",X"00",X"78",X"0E",X"20",X"21",X"00",
		X"40",X"06",X"04",X"79",X"C6",X"2F",X"77",X"2C",X"C2",X"A4",X"1A",X"3C",X"24",X"10",X"F5",X"21",
		X"00",X"40",X"06",X"04",X"79",X"C6",X"2F",X"BE",X"20",X"45",X"2C",X"C2",X"B5",X"1A",X"3C",X"24",
		X"10",X"F3",X"3A",X"00",X"78",X"0D",X"C2",X"9E",X"1A",X"31",X"00",X"44",X"0E",X"20",X"21",X"00",
		X"50",X"06",X"04",X"79",X"C6",X"2F",X"77",X"2C",X"C2",X"D4",X"1A",X"3C",X"24",X"10",X"F5",X"3A",
		X"00",X"78",X"21",X"00",X"50",X"06",X"04",X"79",X"C6",X"2F",X"BE",X"20",X"16",X"2C",X"C2",X"E8",
		X"1A",X"3C",X"24",X"10",X"F3",X"3A",X"00",X"78",X"0D",X"C2",X"CE",X"1A",X"C3",X"74",X"1B",X"3E",
		X"01",X"18",X"05",X"CD",X"61",X"1B",X"3E",X"02",X"32",X"F3",X"51",X"11",X"31",X"1B",X"21",X"33",
		X"52",X"01",X"20",X"00",X"D9",X"06",X"07",X"D9",X"1A",X"77",X"09",X"13",X"D9",X"10",X"F8",X"AF",
		X"32",X"01",X"70",X"3A",X"00",X"78",X"3A",X"00",X"60",X"E6",X"40",X"C2",X"1F",X"1B",X"C3",X"00",
		X"00",X"1D",X"11",X"22",X"10",X"14",X"11",X"12",X"4F",X"3A",X"00",X"60",X"47",X"3A",X"00",X"68",
		X"A0",X"E6",X"04",X"28",X"10",X"79",X"E6",X"0F",X"32",X"D3",X"51",X"79",X"0F",X"0F",X"0F",X"0F",
		X"E6",X"0F",X"32",X"F3",X"51",X"11",X"5A",X"1B",X"18",X"B4",X"1D",X"1F",X"22",X"10",X"14",X"11",
		X"12",X"21",X"00",X"50",X"06",X"04",X"3E",X"10",X"77",X"2C",X"C2",X"68",X"1B",X"24",X"3A",X"00",
		X"78",X"10",X"F3",X"C9",X"CD",X"61",X"1B",X"21",X"00",X"00",X"06",X"28",X"AF",X"86",X"2C",X"C2",
		X"7D",X"1B",X"24",X"4F",X"3A",X"00",X"78",X"79",X"10",X"F3",X"AF",X"C2",X"38",X"1B",X"21",X"00",
		X"40",X"06",X"C0",X"D7",X"3D",X"06",X"40",X"D7",X"AF",X"D7",X"D7",X"06",X"C0",X"D7",X"32",X"01",
		X"70",X"32",X"05",X"70",X"32",X"06",X"70",X"32",X"07",X"70",X"32",X"18",X"40",X"3A",X"00",X"78",
		X"3E",X"20",X"32",X"08",X"40",X"3E",X"03",X"32",X"1A",X"40",X"21",X"C0",X"C0",X"22",X"A0",X"40",
		X"3E",X"01",X"32",X"04",X"70",X"32",X"02",X"70",X"32",X"03",X"70",X"32",X"01",X"70",X"C3",X"00",
		X"20",X"21",X"D8",X"00",X"E5",X"3D",X"CA",X"3E",X"1C",X"3D",X"CA",X"2C",X"1D",X"3D",X"C2",X"00",
		X"00",X"21",X"00",X"58",X"3A",X"1E",X"40",X"77",X"C6",X"2F",X"2C",X"C2",X"E7",X"1B",X"3A",X"1E",
		X"40",X"BE",X"20",X"3C",X"C6",X"2F",X"2C",X"C2",X"F1",X"1B",X"3A",X"00",X"78",X"CD",X"DC",X"16",
		X"21",X"08",X"40",X"35",X"C0",X"AF",X"21",X"00",X"58",X"47",X"D7",X"3E",X"01",X"32",X"06",X"40",
		X"32",X"1A",X"40",X"32",X"00",X"60",X"32",X"01",X"60",X"00",X"00",X"00",X"32",X"26",X"42",X"32",
		X"5F",X"42",X"32",X"38",X"42",X"3E",X"1F",X"32",X"13",X"52",X"3E",X"1B",X"32",X"F3",X"51",X"C9",
		X"21",X"00",X"58",X"AF",X"77",X"2C",X"C2",X"34",X"1C",X"3E",X"03",X"C3",X"08",X"1B",X"CD",X"F9",
		X"16",X"CD",X"8D",X"16",X"3A",X"00",X"78",X"3A",X"00",X"60",X"47",X"E6",X"83",X"28",X"05",X"3E",
		X"01",X"32",X"C9",X"41",X"3A",X"00",X"68",X"4F",X"E6",X"03",X"28",X"05",X"3E",X"16",X"32",X"DF",
		X"41",X"78",X"B1",X"E6",X"0C",X"28",X"05",X"3E",X"06",X"32",X"DF",X"41",X"78",X"B1",X"E6",X"10",
		X"28",X"05",X"3E",X"01",X"32",X"CC",X"41",X"3A",X"00",X"68",X"07",X"07",X"E6",X"03",X"CD",X"D3",
		X"1C",X"3A",X"00",X"70",X"E6",X"03",X"C6",X"04",X"CD",X"D3",X"1C",X"3A",X"00",X"70",X"0F",X"0F",
		X"E6",X"01",X"C6",X"08",X"CD",X"D3",X"1C",X"3A",X"00",X"60",X"E6",X"40",X"C0",X"AF",X"32",X"06",
		X"40",X"3E",X"02",X"32",X"1A",X"40",X"21",X"10",X"30",X"22",X"08",X"40",X"21",X"00",X"50",X"22",
		X"0B",X"40",X"AF",X"21",X"00",X"60",X"06",X"04",X"D7",X"3E",X"01",X"21",X"04",X"60",X"06",X"04",
		X"D7",X"AF",X"06",X"08",X"21",X"00",X"68",X"D7",X"06",X"05",X"21",X"01",X"70",X"D7",X"3D",X"32",
		X"00",X"78",X"C9",X"47",X"87",X"87",X"80",X"5F",X"16",X"00",X"21",X"FA",X"1C",X"19",X"06",X"02",
		X"5E",X"23",X"56",X"23",X"D5",X"10",X"F9",X"46",X"D9",X"E1",X"D1",X"01",X"E0",X"FF",X"D9",X"D9",
		X"1A",X"D6",X"30",X"77",X"13",X"09",X"D9",X"10",X"F6",X"C9",X"12",X"1F",X"D6",X"52",X"10",X"22",
		X"1F",X"D6",X"52",X"10",X"32",X"1F",X"D6",X"52",X"10",X"42",X"1F",X"D6",X"52",X"10",X"52",X"1F",
		X"D8",X"52",X"0A",X"5C",X"1F",X"D8",X"52",X"0A",X"66",X"1F",X"D8",X"52",X"0A",X"70",X"1F",X"D8",
		X"52",X"0A",X"7A",X"1F",X"DA",X"52",X"0A",X"84",X"1F",X"DA",X"52",X"0A",X"21",X"08",X"40",X"3A",
		X"00",X"78",X"7E",X"A7",X"CA",X"55",X"1D",X"D9",X"2A",X"0B",X"40",X"06",X"10",X"36",X"30",X"23",
		X"36",X"32",X"23",X"10",X"F8",X"06",X"10",X"36",X"34",X"23",X"36",X"36",X"23",X"10",X"F8",X"22",
		X"0B",X"40",X"D9",X"35",X"C0",X"23",X"7E",X"A7",X"28",X"02",X"35",X"C0",X"3A",X"00",X"60",X"E6",
		X"40",X"C0",X"21",X"00",X"50",X"22",X"0B",X"40",X"3E",X"20",X"32",X"08",X"40",X"AF",X"32",X"1A",
		X"40",X"32",X"05",X"40",X"C9",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",
		X"06",X"01",X"02",X"02",X"06",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",
		X"04",X"02",X"02",X"02",X"02",X"02",X"00",X"00",X"04",X"05",X"06",X"02",X"02",X"07",X"07",X"07",
		X"00",X"04",X"00",X"04",X"04",X"00",X"04",X"04",X"00",X"04",X"04",X"00",X"04",X"04",X"00",X"04",
		X"04",X"00",X"02",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"01",X"00",X"03",X"00",
		X"02",X"00",X"02",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"21",X"C0",X"43",X"09",X"7E",X"FE",X"02",X"D8",X"DD",X"21",X"A0",X"42",X"C3",X"1E",X"34",X"FD",
		X"CB",X"1F",X"46",X"C2",X"94",X"10",X"3C",X"FE",X"02",X"C3",X"91",X"10",X"3A",X"A4",X"43",X"E6",
		X"03",X"83",X"5F",X"C3",X"F2",X"08",X"DD",X"36",X"00",X"00",X"DD",X"36",X"04",X"FF",X"DD",X"36",
		X"07",X"FF",X"C9",X"DD",X"77",X"04",X"FE",X"F0",X"D2",X"26",X"1E",X"FE",X"10",X"DA",X"26",X"1E",
		X"C3",X"FB",X"2F",X"DD",X"77",X"19",X"3A",X"A9",X"43",X"FE",X"01",X"C2",X"BB",X"33",X"3A",X"0D",
		X"40",X"4F",X"06",X"00",X"21",X"C0",X"43",X"09",X"7E",X"07",X"07",X"07",X"DD",X"77",X"19",X"C3",
		X"BB",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"8A",X"8E",X"8A",X"8E",X"90",X"8D",X"90",X"8D",
		X"8A",X"8E",X"8A",X"8E",X"90",X"8D",X"90",X"8D",X"8A",X"8E",X"90",X"8D",X"8A",X"8E",X"90",X"8D",
		X"8A",X"8E",X"8B",X"8C",X"4A",X"4A",X"2A",X"2E",X"4A",X"4E",X"2A",X"2E",X"4A",X"4E",X"00",X"4A",
		X"2E",X"2A",X"4E",X"2A",X"4E",X"4A",X"2E",X"2A",X"4E",X"4A",X"2E",X"4E",X"0E",X"E0",X"FD",X"36",
		X"00",X"04",X"3A",X"0D",X"40",X"4F",X"06",X"00",X"21",X"AA",X"43",X"09",X"34",X"C9",X"05",X"06",
		X"07",X"08",X"09",X"0A",X"02",X"03",X"05",X"06",X"07",X"08",X"09",X"0A",X"E0",X"15",X"15",X"15",
		X"02",X"02",X"02",X"02",X"15",X"15",X"15",X"02",X"02",X"02",X"15",X"15",X"15",X"E0",X"21",X"00",
		X"68",X"06",X"08",X"77",X"23",X"10",X"FC",X"32",X"38",X"42",X"C9",X"0F",X"10",X"0F",X"E0",X"21",
		X"A3",X"43",X"34",X"CB",X"56",X"C8",X"36",X"00",X"21",X"00",X"50",X"C3",X"7A",X"29",X"21",X"A3",
		X"43",X"34",X"CB",X"56",X"C8",X"36",X"00",X"3A",X"A0",X"43",X"C3",X"9A",X"29",X"DD",X"66",X"04",
		X"DD",X"6E",X"07",X"06",X"08",X"AF",X"FD",X"21",X"A0",X"42",X"11",X"20",X"00",X"C3",X"82",X"10",
		X"3C",X"E0",X"31",X"40",X"43",X"4F",X"49",X"4E",X"40",X"31",X"40",X"43",X"52",X"45",X"44",X"49",
		X"54",X"40",X"32",X"40",X"43",X"4F",X"49",X"4E",X"53",X"40",X"31",X"40",X"43",X"52",X"45",X"44",
		X"49",X"54",X"31",X"40",X"43",X"4F",X"49",X"4E",X"40",X"32",X"40",X"43",X"52",X"45",X"44",X"49",
		X"54",X"53",X"46",X"52",X"45",X"45",X"40",X"50",X"4C",X"41",X"59",X"40",X"40",X"40",X"40",X"40",
		X"40",X"40",X"42",X"4F",X"4E",X"55",X"53",X"40",X"4E",X"4F",X"4E",X"45",X"42",X"4F",X"4E",X"55",
		X"53",X"40",X"34",X"30",X"30",X"30",X"42",X"4F",X"4E",X"55",X"53",X"40",X"35",X"30",X"30",X"30",
		X"42",X"4F",X"4E",X"55",X"53",X"40",X"37",X"30",X"30",X"30",X"47",X"41",X"4C",X"41",X"58",X"49",
		X"50",X"40",X"40",X"33",X"47",X"41",X"4C",X"41",X"58",X"49",X"50",X"40",X"40",X"35",X"00",X"00",
		X"3A",X"91",X"24",X"FE",X"49",X"C2",X"00",X"00",X"3A",X"77",X"23",X"FE",X"8F",X"C2",X"00",X"00",
		X"21",X"88",X"02",X"AF",X"06",X"06",X"AE",X"23",X"10",X"FC",X"FE",X"3F",X"C2",X"00",X"00",X"DD",
		X"CB",X"1B",X"46",X"C3",X"50",X"35",X"32",X"A1",X"43",X"32",X"A2",X"43",X"CD",X"0D",X"09",X"C9",
		X"3A",X"0D",X"40",X"4F",X"06",X"00",X"21",X"C0",X"43",X"09",X"7E",X"A7",X"CA",X"D8",X"1F",X"FA",
		X"D8",X"1F",X"DD",X"6E",X"01",X"C3",X"AF",X"2E",X"DD",X"36",X"18",X"01",X"C9",X"FF",X"FF",X"FF",
		X"3A",X"DE",X"42",X"0F",X"D2",X"36",X"03",X"C3",X"AC",X"25",X"2C",X"34",X"AF",X"21",X"20",X"40",
		X"06",X"20",X"C3",X"77",X"09",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"21",X"A2",X"40",X"06",X"1E",X"36",X"00",X"23",X"10",X"FB",X"26",X"40",X"3A",X"A1",X"40",X"6F",
		X"7E",X"87",X"30",X"05",X"CD",X"67",X"20",X"18",X"F1",X"E6",X"0F",X"4F",X"06",X"00",X"36",X"FF",
		X"2C",X"5E",X"36",X"FF",X"2C",X"7D",X"FE",X"C0",X"30",X"02",X"3E",X"C0",X"32",X"A1",X"40",X"7B",
		X"21",X"3D",X"20",X"09",X"5E",X"23",X"56",X"21",X"0A",X"20",X"E5",X"EB",X"E9",X"55",X"20",X"5E",
		X"20",X"5F",X"21",X"A6",X"21",X"F7",X"21",X"2A",X"22",X"EA",X"22",X"AF",X"24",X"E4",X"7B",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"CD",X"E1",X"20",X"CD",X"04",X"21",X"C3",X"31",X"21",X"CD",X"E1",
		X"20",X"DA",X"78",X"25",X"C3",X"9C",X"25",X"3A",X"5F",X"42",X"47",X"E6",X"0F",X"28",X"2D",X"21",
		X"20",X"41",X"85",X"6F",X"3A",X"38",X"42",X"0F",X"D8",X"0E",X"10",X"06",X"06",X"C5",X"E5",X"7D",
		X"CB",X"46",X"20",X"05",X"CD",X"5E",X"20",X"18",X"0B",X"CD",X"E1",X"20",X"0E",X"00",X"CD",X"1D",
		X"21",X"CD",X"31",X"21",X"E1",X"C1",X"7D",X"81",X"6F",X"10",X"E2",X"C9",X"3A",X"06",X"40",X"A7",
		X"28",X"05",X"32",X"AB",X"40",X"18",X"05",X"3A",X"AB",X"40",X"A7",X"C8",X"3A",X"0D",X"40",X"CD",
		X"4E",X"21",X"11",X"E0",X"FF",X"CB",X"60",X"28",X"14",X"3E",X"10",X"77",X"19",X"77",X"19",X"77",
		X"3A",X"0E",X"40",X"A7",X"C8",X"3A",X"0D",X"40",X"EE",X"01",X"CD",X"4E",X"21",X"3C",X"77",X"19",
		X"36",X"25",X"19",X"36",X"20",X"CB",X"60",X"C0",X"3A",X"06",X"40",X"A7",X"C0",X"32",X"AB",X"40",
		X"C9",X"47",X"E6",X"0F",X"0F",X"0F",X"4F",X"E6",X"03",X"67",X"79",X"E6",X"C0",X"6F",X"78",X"0F",
		X"0F",X"0F",X"0F",X"E6",X"07",X"4F",X"1F",X"F5",X"89",X"2F",X"E6",X"0F",X"85",X"6F",X"11",X"00",
		X"50",X"19",X"F1",X"C9",X"F5",X"78",X"FE",X"70",X"18",X"04",X"06",X"80",X"F1",X"C9",X"E6",X"0F",
		X"47",X"3A",X"5F",X"42",X"E6",X"0F",X"0E",X"00",X"B8",X"30",X"01",X"0D",X"F1",X"F5",X"78",X"FE",
		X"70",X"00",X"00",X"3A",X"5F",X"42",X"0F",X"0F",X"0F",X"0F",X"80",X"81",X"E6",X"03",X"47",X"F1",
		X"C9",X"EB",X"38",X"09",X"21",X"57",X"21",X"78",X"E7",X"EB",X"C3",X"9E",X"25",X"78",X"A7",X"C3",
		X"46",X"21",X"3E",X"A4",X"18",X"04",X"21",X"5B",X"21",X"E7",X"EB",X"C3",X"7A",X"25",X"21",X"40",
		X"53",X"A7",X"C8",X"21",X"E0",X"50",X"C9",X"41",X"35",X"41",X"31",X"44",X"38",X"44",X"3C",X"A7",
		X"28",X"39",X"3D",X"28",X"22",X"3D",X"87",X"87",X"87",X"87",X"2F",X"E6",X"30",X"C6",X"C0",X"21",
		X"D8",X"51",X"CD",X"7A",X"25",X"21",X"DA",X"51",X"CD",X"7A",X"25",X"21",X"18",X"52",X"CD",X"7A",
		X"25",X"21",X"1A",X"52",X"C3",X"7A",X"25",X"21",X"D8",X"51",X"11",X"1C",X"00",X"0E",X"04",X"06",
		X"04",X"36",X"40",X"23",X"10",X"FB",X"19",X"0D",X"20",X"F5",X"C9",X"CD",X"87",X"21",X"3E",X"60",
		X"21",X"FA",X"51",X"C3",X"7A",X"25",X"4F",X"CF",X"CD",X"89",X"22",X"79",X"81",X"81",X"4F",X"06",
		X"00",X"21",X"C9",X"22",X"09",X"A7",X"06",X"03",X"1A",X"8E",X"27",X"12",X"13",X"23",X"10",X"F8",
		X"1B",X"D5",X"1B",X"1A",X"21",X"AC",X"40",X"BE",X"D4",X"95",X"22",X"13",X"3A",X"0D",X"40",X"CD",
		X"4F",X"22",X"D1",X"21",X"AA",X"40",X"06",X"03",X"1A",X"BE",X"D8",X"20",X"05",X"1B",X"2B",X"10",
		X"F7",X"C9",X"CD",X"89",X"22",X"21",X"A8",X"40",X"06",X"03",X"1A",X"77",X"13",X"23",X"10",X"FA",
		X"1B",X"DD",X"21",X"41",X"52",X"18",X"63",X"FE",X"03",X"30",X"26",X"F5",X"21",X"A2",X"40",X"11",
		X"AD",X"40",X"A7",X"28",X"0E",X"21",X"A5",X"40",X"11",X"AE",X"40",X"3D",X"28",X"05",X"21",X"A8",
		X"40",X"5D",X"54",X"36",X"00",X"23",X"36",X"00",X"23",X"36",X"00",X"EB",X"36",X"00",X"F1",X"18",
		X"09",X"3D",X"F5",X"CD",X"F7",X"21",X"F1",X"C8",X"18",X"F7",X"FE",X"03",X"30",X"18",X"A7",X"11",
		X"A4",X"40",X"28",X"1B",X"3D",X"20",X"0A",X"3A",X"0E",X"40",X"A7",X"C8",X"11",X"A7",X"40",X"18",
		X"0E",X"11",X"AA",X"40",X"18",X"AB",X"3D",X"F5",X"CD",X"2A",X"22",X"F1",X"C8",X"18",X"F7",X"DD",
		X"21",X"81",X"53",X"A7",X"28",X"04",X"DD",X"21",X"21",X"51",X"21",X"E0",X"FF",X"EB",X"06",X"03",
		X"0E",X"04",X"7E",X"0F",X"0F",X"0F",X"0F",X"CD",X"72",X"22",X"7E",X"CD",X"72",X"22",X"2B",X"10",
		X"F1",X"C9",X"E6",X"0F",X"28",X"04",X"0E",X"00",X"18",X"07",X"79",X"A7",X"28",X"03",X"3E",X"10",
		X"0D",X"C6",X"00",X"DD",X"77",X"00",X"DD",X"19",X"C9",X"11",X"A2",X"40",X"3A",X"0D",X"40",X"A7",
		X"C8",X"11",X"A5",X"40",X"C9",X"3A",X"0D",X"40",X"21",X"AD",X"40",X"85",X"6F",X"CB",X"46",X"C0",
		X"36",X"01",X"3E",X"01",X"32",X"C7",X"41",X"21",X"1D",X"42",X"34",X"46",X"21",X"9E",X"53",X"0E",
		X"05",X"3A",X"00",X"42",X"A7",X"28",X"03",X"05",X"28",X"08",X"3E",X"66",X"CD",X"88",X"25",X"0D",
		X"10",X"F8",X"0D",X"F8",X"CD",X"86",X"25",X"18",X"F9",X"20",X"00",X"00",X"30",X"00",X"00",X"40",
		X"00",X"00",X"50",X"00",X"00",X"00",X"01",X"00",X"00",X"02",X"00",X"00",X"03",X"00",X"00",X"04",
		X"00",X"00",X"05",X"00",X"00",X"36",X"01",X"C3",X"95",X"37",X"21",X"55",X"23",X"87",X"F5",X"E6",
		X"3F",X"5F",X"16",X"00",X"19",X"5E",X"23",X"56",X"EB",X"5E",X"23",X"56",X"23",X"EB",X"01",X"E0",
		X"FF",X"F1",X"38",X"0E",X"FA",X"1C",X"23",X"1A",X"D6",X"30",X"FE",X"0F",X"C8",X"77",X"13",X"09",
		X"18",X"F5",X"1A",X"FE",X"3F",X"C8",X"36",X"40",X"13",X"09",X"18",X"F6",X"22",X"B5",X"40",X"EB",
		X"22",X"B3",X"40",X"7B",X"E6",X"1F",X"47",X"87",X"C6",X"20",X"6F",X"26",X"40",X"22",X"B1",X"40",
		X"E5",X"CB",X"3B",X"CB",X"3B",X"7A",X"E6",X"03",X"0F",X"0F",X"B3",X"E6",X"F8",X"4F",X"21",X"00",
		X"50",X"78",X"85",X"6F",X"11",X"20",X"00",X"43",X"36",X"10",X"19",X"10",X"FB",X"E1",X"71",X"3E",
		X"01",X"32",X"B0",X"40",X"C9",X"7B",X"23",X"88",X"23",X"9E",X"23",X"AB",X"23",X"B8",X"23",X"C4",
		X"23",X"CF",X"23",X"EA",X"23",X"F9",X"23",X"09",X"24",X"1D",X"24",X"29",X"24",X"3A",X"24",X"4B",
		X"24",X"5C",X"24",X"6D",X"24",X"7E",X"24",X"8F",X"24",X"96",X"24",X"96",X"52",X"47",X"41",X"4D",
		X"45",X"40",X"40",X"4F",X"56",X"45",X"52",X"3F",X"0F",X"53",X"50",X"55",X"53",X"48",X"40",X"53",
		X"45",X"4C",X"45",X"43",X"54",X"40",X"42",X"55",X"54",X"54",X"4F",X"4E",X"40",X"3F",X"94",X"52",
		X"50",X"4C",X"41",X"59",X"45",X"52",X"40",X"30",X"4E",X"45",X"3F",X"94",X"52",X"50",X"4C",X"41",
		X"59",X"45",X"52",X"40",X"54",X"57",X"4F",X"3F",X"60",X"52",X"54",X"4F",X"50",X"40",X"53",X"43",
		X"4F",X"52",X"45",X"3F",X"BF",X"53",X"43",X"52",X"45",X"44",X"49",X"54",X"40",X"40",X"3F",X"75",
		X"53",X"40",X"42",X"4F",X"4E",X"55",X"53",X"40",X"53",X"48",X"49",X"50",X"40",X"46",X"4F",X"52",
		X"40",X"40",X"40",X"30",X"30",X"40",X"50",X"54",X"53",X"3F",X"AB",X"52",X"50",X"4F",X"49",X"4E",
		X"54",X"40",X"53",X"59",X"53",X"54",X"45",X"4D",X"3F",X"28",X"52",X"53",X"54",X"52",X"49",X"4B",
		X"45",X"53",X"40",X"42",X"41",X"43",X"4B",X"40",X"3F",X"46",X"53",X"54",X"48",X"45",X"40",X"47",
		X"41",X"4C",X"41",X"58",X"59",X"40",X"45",X"4D",X"50",X"49",X"52",X"45",X"3F",X"63",X"52",X"41",
		X"54",X"54",X"45",X"4E",X"54",X"49",X"4F",X"4E",X"3F",X"8D",X"52",X"8E",X"8E",X"8E",X"8E",X"8E",
		X"8E",X"40",X"40",X"32",X"30",X"40",X"50",X"54",X"53",X"3F",X"90",X"52",X"8E",X"8E",X"8E",X"8E",
		X"8E",X"8E",X"40",X"40",X"33",X"30",X"40",X"50",X"54",X"53",X"3F",X"93",X"52",X"8E",X"8E",X"8E",
		X"8E",X"8E",X"8E",X"40",X"40",X"34",X"30",X"40",X"50",X"54",X"53",X"3F",X"96",X"52",X"8E",X"8E",
		X"8E",X"8E",X"8E",X"8E",X"40",X"40",X"35",X"30",X"40",X"50",X"54",X"53",X"3F",X"99",X"52",X"8E",
		X"8E",X"8E",X"8E",X"8E",X"8E",X"40",X"31",X"30",X"30",X"40",X"50",X"54",X"53",X"3F",X"9C",X"52",
		X"8E",X"8E",X"8E",X"8E",X"8E",X"8E",X"40",X"42",X"49",X"47",X"40",X"50",X"54",X"53",X"3F",X"3F",
		X"52",X"49",X"52",X"45",X"4D",X"3F",X"7F",X"53",X"46",X"52",X"45",X"45",X"40",X"50",X"4C",X"41",
		X"59",X"3F",X"3F",X"7F",X"53",X"46",X"52",X"45",X"45",X"40",X"50",X"4C",X"41",X"59",X"3F",X"A7",
		X"28",X"63",X"3D",X"28",X"2B",X"3D",X"28",X"08",X"3A",X"1D",X"42",X"47",X"CF",X"C3",X"AC",X"22",
		X"3A",X"AC",X"40",X"FE",X"FF",X"C8",X"3E",X"06",X"CD",X"EA",X"22",X"3A",X"AC",X"40",X"E6",X"0F",
		X"32",X"55",X"51",X"3A",X"AC",X"40",X"E6",X"F0",X"0F",X"0F",X"0F",X"0F",X"32",X"75",X"51",X"C9",
		X"3A",X"06",X"40",X"0F",X"D8",X"3A",X"11",X"40",X"E6",X"C0",X"FE",X"C0",X"3E",X"12",X"CA",X"EA",
		X"22",X"3E",X"05",X"CD",X"EA",X"22",X"3A",X"02",X"40",X"FE",X"63",X"38",X"02",X"3E",X"63",X"CD",
		X"5E",X"25",X"47",X"E6",X"F0",X"28",X"07",X"0F",X"0F",X"0F",X"0F",X"32",X"DF",X"52",X"78",X"E6",
		X"0F",X"32",X"BF",X"52",X"C9",X"CF",X"3A",X"20",X"42",X"A7",X"28",X"05",X"3E",X"01",X"32",X"D0",
		X"41",X"3A",X"1C",X"42",X"3C",X"FE",X"30",X"38",X"02",X"3E",X"30",X"CD",X"5E",X"25",X"F5",X"21",
		X"7E",X"50",X"E6",X"F0",X"28",X"10",X"0F",X"0F",X"0F",X"0F",X"47",X"0E",X"10",X"3E",X"68",X"CD",
		X"7A",X"25",X"0D",X"0D",X"10",X"F7",X"F1",X"E6",X"0F",X"47",X"11",X"1F",X"00",X"28",X"08",X"3E",
		X"6C",X"CD",X"95",X"25",X"0D",X"10",X"F8",X"0D",X"F8",X"CD",X"93",X"25",X"18",X"F9",X"47",X"E6",
		X"0F",X"C6",X"00",X"27",X"4F",X"78",X"E6",X"F0",X"28",X"0B",X"0F",X"0F",X"0F",X"0F",X"47",X"AF",
		X"C6",X"16",X"27",X"10",X"FB",X"81",X"27",X"C9",X"3E",X"2C",X"D5",X"11",X"1F",X"00",X"CD",X"95",
		X"25",X"CD",X"95",X"25",X"D1",X"C9",X"3E",X"2E",X"D5",X"11",X"DF",X"FF",X"CD",X"95",X"25",X"C6",
		X"FC",X"18",X"EE",X"3E",X"2C",X"77",X"3C",X"23",X"77",X"3C",X"19",X"C9",X"3E",X"2C",X"D5",X"11",
		X"20",X"00",X"77",X"C6",X"02",X"19",X"77",X"D1",X"C9",X"3A",X"0D",X"40",X"4F",X"06",X"00",X"21",
		X"C0",X"43",X"09",X"3A",X"A9",X"43",X"36",X"10",X"FE",X"02",X"20",X"02",X"36",X"08",X"CD",X"18",
		X"2E",X"C9",X"C0",X"EB",X"3A",X"0D",X"40",X"4F",X"06",X"00",X"21",X"C0",X"43",X"09",X"7E",X"07",
		X"EB",X"C6",X"0F",X"77",X"C3",X"5F",X"32",X"28",X"0A",X"DD",X"7E",X"02",X"A7",X"CA",X"BA",X"32",
		X"C3",X"CB",X"32",X"DD",X"7E",X"02",X"A7",X"CA",X"CB",X"32",X"C3",X"BA",X"32",X"DD",X"7E",X"02",
		X"EE",X"01",X"DD",X"77",X"02",X"C3",X"CB",X"32",X"DD",X"7E",X"02",X"EE",X"01",X"DD",X"77",X"02",
		X"C3",X"BA",X"32",X"21",X"AA",X"43",X"09",X"36",X"00",X"C3",X"F4",X"35",X"DD",X"7E",X"04",X"D6",
		X"08",X"C9",X"36",X"00",X"21",X"1C",X"50",X"06",X"20",X"11",X"20",X"00",X"36",X"5E",X"19",X"10",
		X"FB",X"C9",X"21",X"BE",X"43",X"34",X"7E",X"FE",X"10",X"20",X"15",X"21",X"A0",X"42",X"06",X"00",
		X"AF",X"D7",X"21",X"1C",X"50",X"06",X"20",X"11",X"20",X"00",X"36",X"40",X"19",X"10",X"FB",X"C9",
		X"FE",X"20",X"20",X"20",X"01",X"57",X"26",X"21",X"AE",X"52",X"11",X"E0",X"FF",X"0A",X"A7",X"28",
		X"05",X"77",X"19",X"03",X"18",X"F7",X"C9",X"1E",X"15",X"28",X"24",X"10",X"20",X"11",X"24",X"24",
		X"15",X"22",X"1E",X"00",X"FE",X"80",X"20",X"08",X"01",X"0C",X"37",X"C3",X"47",X"26",X"D7",X"C9",
		X"FE",X"C0",X"C0",X"36",X"00",X"21",X"22",X"42",X"C3",X"78",X"37",X"7F",X"7E",X"00",X"00",X"00",
		X"3A",X"0D",X"40",X"4F",X"06",X"00",X"21",X"AA",X"43",X"09",X"3E",X"07",X"96",X"57",X"21",X"C0",
		X"43",X"09",X"7E",X"92",X"4F",X"DD",X"21",X"A0",X"42",X"C9",X"CD",X"46",X"37",X"0D",X"F8",X"DD",
		X"36",X"18",X"00",X"C9",X"0F",X"0F",X"E6",X"07",X"32",X"62",X"40",X"3E",X"24",X"32",X"61",X"40",
		X"3E",X"78",X"32",X"60",X"40",X"3E",X"7F",X"32",X"63",X"40",X"C3",X"4C",X"28",X"DD",X"CB",X"08",
		X"46",X"C2",X"35",X"2E",X"DD",X"36",X"04",X"00",X"DD",X"36",X"07",X"00",X"C3",X"31",X"2E",X"3A",
		X"BF",X"43",X"A7",X"C2",X"D2",X"35",X"7E",X"FE",X"02",X"C2",X"D2",X"35",X"35",X"3E",X"01",X"C3",
		X"FC",X"36",X"C9",X"21",X"A0",X"42",X"06",X"00",X"AF",X"D7",X"32",X"BF",X"43",X"21",X"1C",X"50",
		X"C9",X"CD",X"F8",X"39",X"3E",X"01",X"32",X"BF",X"43",X"C9",X"C2",X"95",X"37",X"C3",X"E5",X"22",
		X"2A",X"C7",X"41",X"CB",X"45",X"CA",X"11",X"27",X"21",X"00",X"80",X"22",X"C7",X"41",X"C3",X"D3",
		X"27",X"7C",X"A7",X"CA",X"D3",X"27",X"CD",X"65",X"18",X"C3",X"16",X"17",X"00",X"36",X"C3",X"C9",
		X"FE",X"01",X"20",X"05",X"36",X"01",X"C3",X"CA",X"27",X"FE",X"02",X"20",X"05",X"36",X"02",X"C3",
		X"CA",X"27",X"FE",X"03",X"20",X"05",X"36",X"03",X"C3",X"CA",X"27",X"36",X"00",X"C3",X"CA",X"27",
		X"C4",X"92",X"3A",X"3A",X"B9",X"43",X"C3",X"3E",X"3A",X"3A",X"5F",X"42",X"0F",X"0F",X"0F",X"85",
		X"3A",X"07",X"40",X"0F",X"D2",X"C4",X"3A",X"1E",X"00",X"C3",X"C4",X"3A",X"00",X"00",X"00",X"20",
		X"C4",X"67",X"27",X"3A",X"B9",X"43",X"C9",X"5F",X"16",X"00",X"21",X"18",X"3B",X"19",X"19",X"5E",
		X"23",X"56",X"EB",X"C3",X"81",X"3A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CB",X"7D",X"CA",X"A0",X"2A",X"C3",X"6B",X"2A",X"CB",X"75",X"CA",X"F1",X"2A",X"C3",X"CC",X"2A",
		X"CD",X"63",X"03",X"3A",X"AB",X"43",X"C9",X"CD",X"D3",X"2B",X"21",X"B5",X"1D",X"CD",X"98",X"05",
		X"C9",X"32",X"38",X"42",X"06",X"10",X"AF",X"21",X"A0",X"43",X"D7",X"C9",X"3A",X"0D",X"40",X"4F",
		X"06",X"00",X"21",X"A1",X"43",X"09",X"7E",X"A7",X"20",X"07",X"AF",X"32",X"C0",X"41",X"C3",X"FD",
		X"16",X"3A",X"A9",X"43",X"21",X"BD",X"43",X"C3",X"20",X"27",X"CD",X"27",X"17",X"CD",X"BA",X"3A",
		X"C3",X"00",X"27",X"C3",X"A3",X"13",X"CD",X"00",X"3A",X"C9",X"00",X"00",X"27",X"17",X"CD",X"BA",
		X"3A",X"CD",X"00",X"3A",X"C9",X"32",X"B8",X"43",X"3E",X"01",X"32",X"BC",X"43",X"C9",X"3A",X"BC",
		X"43",X"0F",X"DA",X"48",X"3A",X"3E",X"FF",X"32",X"00",X"78",X"AF",X"32",X"BC",X"43",X"C9",X"00",
		X"23",X"35",X"7E",X"FE",X"FF",X"20",X"06",X"11",X"01",X"02",X"C3",X"BD",X"28",X"FE",X"F0",X"20",
		X"1A",X"3E",X"01",X"32",X"04",X"68",X"3E",X"27",X"32",X"2D",X"52",X"3E",X"11",X"32",X"0D",X"52",
		X"3E",X"22",X"32",X"ED",X"51",X"3E",X"20",X"32",X"CD",X"51",X"C9",X"FE",X"D0",X"30",X"34",X"FE",
		X"81",X"38",X"24",X"2F",X"32",X"00",X"78",X"2F",X"32",X"63",X"40",X"0F",X"0F",X"E6",X"07",X"32",
		X"62",X"40",X"3E",X"18",X"32",X"61",X"40",X"3E",X"78",X"32",X"60",X"40",X"3E",X"00",X"32",X"06",
		X"00",X"3E",X"00",X"32",X"07",X"68",X"C9",X"FE",X"31",X"38",X"08",X"2F",X"32",X"00",X"78",X"00",
		X"C3",X"A4",X"26",X"FE",X"30",X"20",X"13",X"3E",X"FF",X"32",X"00",X"78",X"AF",X"32",X"60",X"40",
		X"32",X"61",X"40",X"32",X"62",X"40",X"32",X"63",X"40",X"C9",X"FE",X"10",X"20",X"13",X"AF",X"32",
		X"04",X"68",X"3E",X"10",X"32",X"2D",X"52",X"32",X"0D",X"52",X"32",X"ED",X"51",X"32",X"CD",X"51",
		X"C9",X"FE",X"05",X"20",X"06",X"11",X"00",X"02",X"C3",X"C9",X"28",X"A7",X"C0",X"C3",X"D9",X"39",
		X"3A",X"08",X"42",X"2A",X"00",X"42",X"B4",X"B5",X"0F",X"30",X"06",X"21",X"22",X"42",X"C3",X"EE",
		X"28",X"C3",X"F6",X"28",X"CB",X"46",X"C8",X"23",X"35",X"C0",X"C3",X"27",X"16",X"AF",X"32",X"00",
		X"42",X"3E",X"01",X"32",X"08",X"42",X"C3",X"A8",X"39",X"3E",X"01",X"CD",X"12",X"29",X"AF",X"32",
		X"08",X"42",X"C3",X"03",X"29",X"3A",X"00",X"42",X"0F",X"38",X"05",X"3A",X"01",X"42",X"0F",X"D0",
		X"3A",X"0B",X"42",X"C3",X"E8",X"08",X"3A",X"23",X"42",X"A7",X"C0",X"2C",X"34",X"C9",X"3E",X"01",
		X"32",X"A0",X"43",X"C3",X"21",X"16",X"3A",X"A0",X"43",X"A7",X"C2",X"AB",X"28",X"21",X"22",X"42",
		X"C3",X"B4",X"28",X"AF",X"32",X"A0",X"43",X"3E",X"80",X"32",X"02",X"42",X"32",X"0A",X"42",X"C3",
		X"F2",X"08",X"3A",X"08",X"42",X"32",X"00",X"42",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"CD",X"A0",X"39",X"4F",X"06",X"00",X"21",X"49",X"29",X"09",X"09",X"5E",X"23",X"56",X"00",X"00",
		X"00",X"00",X"EB",X"E9",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"10",X"21",X"A0",X"43",X"AF",
		X"D7",X"21",X"20",X"06",X"C9",X"00",X"C3",X"1B",X"02",X"61",X"29",X"77",X"29",X"97",X"29",X"D4",
		X"29",X"61",X"2A",X"C6",X"2A",X"03",X"2B",X"76",X"2B",X"90",X"2B",X"A6",X"2B",X"46",X"29",X"FF",
		X"FF",X"06",X"1C",X"00",X"21",X"24",X"40",X"0E",X"06",X"77",X"23",X"71",X"23",X"10",X"FA",X"3E",
		X"02",X"32",X"A0",X"43",X"C3",X"D3",X"2B",X"C3",X"DF",X"1E",X"3A",X"A0",X"43",X"4F",X"06",X"00",
		X"09",X"11",X"20",X"00",X"43",X"36",X"6E",X"19",X"10",X"FB",X"3A",X"A0",X"43",X"3C",X"32",X"A0",
		X"43",X"FE",X"1E",X"C0",X"C3",X"D3",X"2B",X"C3",X"EE",X"1E",X"00",X"00",X"00",X"00",X"21",X"00",
		X"50",X"3A",X"A0",X"43",X"4F",X"06",X"00",X"09",X"11",X"20",X"00",X"43",X"36",X"40",X"19",X"10",
		X"FB",X"3A",X"A0",X"43",X"3D",X"32",X"A0",X"43",X"FE",X"01",X"C0",X"CD",X"D3",X"2B",X"AF",X"06",
		X"03",X"21",X"A0",X"43",X"77",X"23",X"10",X"FC",X"06",X"07",X"21",X"A4",X"43",X"77",X"23",X"C6",
		X"20",X"10",X"FA",X"C9",X"2A",X"A1",X"43",X"23",X"22",X"A1",X"43",X"CB",X"6D",X"CA",X"F2",X"29",
		X"CD",X"B0",X"2B",X"3A",X"A0",X"43",X"3C",X"32",X"A0",X"43",X"FE",X"08",X"C2",X"F2",X"29",X"C3",
		X"D3",X"2B",X"3A",X"A0",X"43",X"4F",X"00",X"00",X"06",X"00",X"0D",X"F8",X"CD",X"02",X"2A",X"C3",
		X"FA",X"29",X"21",X"60",X"40",X"09",X"09",X"09",X"09",X"EB",X"21",X"A4",X"43",X"00",X"09",X"7E",
		X"34",X"34",X"C5",X"4F",X"06",X"00",X"21",X"00",X"2C",X"09",X"7E",X"4F",X"12",X"23",X"13",X"13",
		X"13",X"7E",X"12",X"47",X"1B",X"00",X"78",X"A9",X"E6",X"07",X"12",X"1B",X"E6",X"01",X"F6",X"24",
		X"12",X"C1",X"C9",X"21",X"60",X"40",X"09",X"09",X"09",X"09",X"EB",X"21",X"A4",X"43",X"09",X"7E",
		X"34",X"34",X"C5",X"4F",X"06",X"00",X"21",X"00",X"2C",X"09",X"7E",X"4F",X"23",X"13",X"13",X"13",
		X"7E",X"47",X"1B",X"00",X"78",X"A9",X"E6",X"07",X"12",X"1B",X"E6",X"01",X"F6",X"24",X"12",X"C1",
		X"C9",X"2A",X"A1",X"43",X"23",X"22",X"A1",X"43",X"C3",X"80",X"27",X"CD",X"B0",X"2B",X"CD",X"CE",
		X"2B",X"3A",X"A3",X"43",X"FE",X"08",X"C2",X"82",X"2A",X"CD",X"B7",X"2B",X"CD",X"BC",X"2B",X"C3",
		X"D3",X"2B",X"3A",X"A3",X"43",X"3D",X"CD",X"D8",X"2B",X"21",X"F0",X"2B",X"09",X"5E",X"23",X"56",
		X"21",X"60",X"40",X"09",X"09",X"73",X"23",X"23",X"23",X"72",X"3A",X"A2",X"43",X"E6",X"03",X"C0",
		X"3A",X"A3",X"43",X"4F",X"0D",X"06",X"00",X"0C",X"3E",X"07",X"00",X"B9",X"CA",X"B5",X"2A",X"CD",
		X"02",X"2A",X"C3",X"A7",X"2A",X"06",X"00",X"0E",X"FF",X"0C",X"3A",X"A3",X"43",X"B9",X"C8",X"7E",
		X"CD",X"33",X"2A",X"C3",X"B9",X"2A",X"CD",X"C1",X"2B",X"C3",X"88",X"27",X"CD",X"B0",X"2B",X"CD",
		X"CE",X"2B",X"7E",X"FE",X"08",X"C2",X"DB",X"2A",X"C3",X"D3",X"2B",X"3A",X"A3",X"43",X"4F",X"0D",
		X"06",X"00",X"21",X"61",X"40",X"09",X"09",X"09",X"09",X"23",X"36",X"00",X"2B",X"3E",X"29",X"81",
		X"77",X"3A",X"A3",X"43",X"3D",X"4F",X"06",X"00",X"0C",X"3E",X"07",X"B9",X"C8",X"CD",X"33",X"2A",
		X"C3",X"F8",X"2A",X"3A",X"A3",X"43",X"C3",X"DD",X"2B",X"AF",X"32",X"A3",X"43",X"CD",X"19",X"2B",
		X"CD",X"C1",X"2B",X"CB",X"7D",X"C8",X"C3",X"D3",X"2B",X"3A",X"A0",X"43",X"4F",X"06",X"00",X"21",
		X"60",X"40",X"09",X"09",X"09",X"09",X"46",X"E5",X"D1",X"23",X"23",X"23",X"4E",X"CD",X"3A",X"2B",
		X"CD",X"C9",X"2B",X"3E",X"07",X"BE",X"C3",X"E6",X"2B",X"C9",X"78",X"FE",X"7C",X"C2",X"4B",X"2B",
		X"79",X"FE",X"C5",X"C2",X"47",X"2B",X"C9",X"CD",X"6A",X"2B",X"C9",X"79",X"FE",X"C5",X"C2",X"55",
		X"2B",X"CD",X"5C",X"2B",X"C9",X"CD",X"5C",X"2B",X"CD",X"6A",X"2B",X"C9",X"78",X"FE",X"7C",X"DA",
		X"66",X"2B",X"05",X"78",X"12",X"C9",X"04",X"78",X"12",X"C9",X"79",X"FE",X"C5",X"DA",X"73",X"2B",
		X"0D",X"71",X"C9",X"0C",X"71",X"C9",X"21",X"60",X"40",X"AF",X"06",X"20",X"77",X"23",X"10",X"FC",
		X"21",X"10",X"04",X"22",X"05",X"42",X"11",X"05",X"02",X"CD",X"F2",X"08",X"CD",X"D3",X"2B",X"C9",
		X"21",X"05",X"42",X"35",X"C0",X"36",X"10",X"23",X"16",X"02",X"5E",X"CD",X"F2",X"08",X"35",X"C0",
		X"CD",X"B0",X"2B",X"C3",X"D3",X"2B",X"CD",X"C1",X"2B",X"CB",X"5D",X"C8",X"CD",X"97",X"27",X"C9",
		X"21",X"00",X"00",X"22",X"A1",X"43",X"C9",X"AF",X"32",X"A0",X"43",X"C9",X"AF",X"32",X"A3",X"43",
		X"C9",X"2A",X"A1",X"43",X"23",X"22",X"A1",X"43",X"C9",X"21",X"A0",X"43",X"34",X"C9",X"21",X"A3",
		X"43",X"34",X"C9",X"21",X"AB",X"43",X"34",X"C9",X"07",X"4F",X"06",X"00",X"C9",X"CD",X"CE",X"2B",
		X"CB",X"47",X"C8",X"C3",X"09",X"2B",X"C2",X"19",X"2B",X"C3",X"B7",X"2B",X"FF",X"FF",X"FF",X"FF",
		X"40",X"70",X"50",X"70",X"60",X"70",X"70",X"70",X"80",X"70",X"90",X"70",X"B0",X"70",X"00",X"00",
		X"B7",X"28",X"B1",X"2D",X"A6",X"2E",X"A3",X"30",X"9A",X"33",X"93",X"3E",X"88",X"42",X"81",X"49",
		X"79",X"54",X"72",X"5D",X"67",X"60",X"64",X"65",X"59",X"6A",X"52",X"6F",X"49",X"6E",X"38",X"6B",
		X"32",X"68",X"29",X"61",X"22",X"5E",X"1A",X"53",X"19",X"4C",X"19",X"41",X"18",X"38",X"19",X"34",
		X"22",X"32",X"29",X"2F",X"32",X"2C",X"38",X"29",X"47",X"28",X"52",X"2B",X"5A",X"30",X"60",X"3E",
		X"6B",X"44",X"70",X"4D",X"73",X"52",X"78",X"5B",X"7D",X"84",X"80",X"8F",X"83",X"92",X"8A",X"9D",
		X"8D",X"B2",X"92",X"B7",X"95",X"B9",X"A7",X"BA",X"A7",X"BA",X"A7",X"BA",X"A7",X"BA",X"A7",X"BA",
		X"B1",X"C0",X"BA",X"C3",X"D2",X"C5",X"DB",X"CA",X"C4",X"C7",X"C9",X"C2",X"E0",X"BF",X"E3",X"B6",
		X"E4",X"B1",X"E8",X"AE",X"E3",X"A8",X"DA",X"A5",X"D2",X"A2",X"CB",X"9F",X"C0",X"9B",X"BE",X"9F",
		X"AA",X"9A",X"A1",X"97",X"98",X"93",X"93",X"90",X"8C",X"8D",X"85",X"8A",X"7C",X"87",X"73",X"8E",
		X"68",X"92",X"65",X"9F",X"5C",X"A2",X"53",X"AF",X"4C",X"B4",X"46",X"BD",X"2E",X"C2",X"33",X"C2",
		X"2F",X"C8",X"22",X"C9",X"18",X"C5",X"13",X"C2",X"13",X"BF",X"13",X"B6",X"13",X"AD",X"18",X"A4",
		X"20",X"9F",X"2A",X"96",X"2F",X"8D",X"32",X"8D",X"3A",X"8B",X"44",X"8B",X"48",X"89",X"50",X"8A",
		X"59",X"86",X"62",X"85",X"6B",X"84",X"74",X"83",X"7E",X"82",X"80",X"81",X"8F",X"7D",X"94",X"79",
		X"99",X"72",X"99",X"6F",X"99",X"6F",X"99",X"6F",X"A0",X"6B",X"A3",X"6B",X"A4",X"69",X"A7",X"69",
		X"AE",X"69",X"B2",X"62",X"BB",X"5F",X"BE",X"5A",X"D4",X"57",X"D7",X"54",X"DA",X"50",X"D7",X"4D",
		X"D4",X"48",X"AE",X"43",X"AE",X"41",X"AE",X"3E",X"AD",X"3A",X"BA",X"34",X"B9",X"31",X"B7",X"28",
		X"2A",X"A4",X"43",X"23",X"22",X"A4",X"43",X"C3",X"A3",X"2D",X"3A",X"0D",X"40",X"4F",X"06",X"00",
		X"21",X"C2",X"43",X"09",X"09",X"09",X"06",X"08",X"DD",X"21",X"A0",X"42",X"11",X"20",X"00",X"DD",
		X"CB",X"08",X"46",X"CA",X"2B",X"2D",X"DD",X"7E",X"04",X"77",X"23",X"DD",X"19",X"10",X"F0",X"21",
		X"A0",X"42",X"C9",X"DD",X"36",X"1C",X"00",X"C3",X"5B",X"2D",X"C3",X"99",X"10",X"DD",X"CB",X"1F",
		X"46",X"C3",X"AC",X"10",X"00",X"00",X"3A",X"0D",X"40",X"4F",X"06",X"00",X"21",X"C0",X"43",X"09",
		X"18",X"31",X"DD",X"36",X"00",X"00",X"DD",X"36",X"18",X"00",X"C9",X"3A",X"A9",X"43",X"FE",X"01",
		X"CA",X"46",X"2D",X"DD",X"7E",X"00",X"C3",X"3A",X"2D",X"D2",X"E7",X"35",X"21",X"C0",X"43",X"09",
		X"7E",X"FE",X"04",X"DA",X"E7",X"35",X"C5",X"CD",X"46",X"2D",X"C1",X"21",X"AA",X"43",X"09",X"34",
		X"C3",X"CF",X"26",X"EB",X"21",X"AA",X"43",X"09",X"7E",X"A7",X"28",X"01",X"3C",X"EB",X"86",X"FE",
		X"09",X"38",X"04",X"35",X"C3",X"52",X"2D",X"35",X"C9",X"D3",X"52",X"E5",X"52",X"8F",X"53",X"A4",
		X"53",X"E7",X"53",X"21",X"A8",X"43",X"7E",X"A7",X"C2",X"E8",X"2D",X"36",X"01",X"CD",X"E3",X"26",
		X"06",X"20",X"11",X"20",X"00",X"36",X"5E",X"19",X"10",X"FB",X"CD",X"20",X"38",X"35",X"CD",X"18",
		X"2E",X"3A",X"0D",X"40",X"4F",X"06",X"00",X"21",X"A6",X"43",X"09",X"7E",X"32",X"A9",X"43",X"21",
		X"AA",X"43",X"09",X"46",X"DD",X"21",X"80",X"43",X"CD",X"E8",X"39",X"78",X"B7",X"C3",X"3F",X"00",
		X"7E",X"CD",X"F1",X"26",X"DD",X"19",X"10",X"F8",X"3A",X"A9",X"43",X"4F",X"06",X"00",X"21",X"FC",
		X"2D",X"09",X"09",X"5E",X"23",X"56",X"21",X"06",X"2E",X"E5",X"EB",X"E9",X"18",X"2E",X"4A",X"2E",
		X"41",X"30",X"1C",X"32",X"49",X"2E",X"CD",X"89",X"34",X"CD",X"57",X"33",X"CD",X"39",X"35",X"3A",
		X"A9",X"43",X"FE",X"04",X"00",X"C3",X"72",X"37",X"06",X"08",X"DD",X"21",X"A0",X"42",X"11",X"20",
		X"00",X"DD",X"36",X"00",X"00",X"DD",X"36",X"01",X"00",X"DD",X"36",X"02",X"00",X"C3",X"BD",X"26",
		X"00",X"DD",X"36",X"18",X"00",X"DD",X"36",X"1B",X"00",X"DD",X"36",X"1C",X"00",X"DD",X"36",X"1F",
		X"00",X"DD",X"19",X"10",X"DC",X"C3",X"00",X"38",X"34",X"C9",X"DD",X"21",X"A0",X"42",X"11",X"20",
		X"00",X"06",X"08",X"D9",X"CD",X"80",X"2E",X"D9",X"DD",X"19",X"10",X"F7",X"CD",X"60",X"2E",X"C9",
		X"DD",X"21",X"A0",X"42",X"11",X"20",X"00",X"06",X"08",X"3E",X"01",X"DD",X"A6",X"18",X"00",X"00",
		X"00",X"DD",X"19",X"10",X"F6",X"CB",X"47",X"C8",X"C3",X"53",X"36",X"CD",X"A9",X"25",X"00",X"C9",
		X"CD",X"9B",X"2E",X"DD",X"7E",X"00",X"EF",X"AC",X"2E",X"C8",X"2E",X"38",X"2F",X"58",X"2F",X"8C",
		X"2F",X"BE",X"2F",X"E3",X"2F",X"09",X"30",X"FF",X"FF",X"FF",X"FF",X"DD",X"CB",X"08",X"46",X"C2",
		X"AA",X"2E",X"DD",X"CB",X"18",X"46",X"C2",X"83",X"36",X"C9",X"F1",X"C9",X"C3",X"C0",X"1F",X"DD",
		X"66",X"02",X"23",X"DD",X"75",X"01",X"DD",X"74",X"02",X"C3",X"CB",X"39",X"DD",X"36",X"01",X"00",
		X"DD",X"36",X"02",X"00",X"DD",X"34",X"00",X"C9",X"DD",X"34",X"01",X"DD",X"7E",X"01",X"FE",X"04",
		X"C0",X"DD",X"36",X"01",X"00",X"DD",X"7E",X"02",X"D9",X"80",X"D9",X"E6",X"07",X"47",X"DD",X"7E",
		X"03",X"2F",X"10",X"FD",X"DD",X"77",X"03",X"A7",X"CA",X"F2",X"2E",X"DD",X"36",X"05",X"24",X"C3",
		X"F6",X"2E",X"DD",X"36",X"05",X"25",X"DD",X"7E",X"02",X"D9",X"80",X"D9",X"E6",X"07",X"DD",X"77",
		X"06",X"D9",X"78",X"CD",X"C3",X"39",X"4F",X"06",X"00",X"21",X"28",X"2F",X"09",X"09",X"7E",X"DD",
		X"77",X"04",X"23",X"7E",X"DD",X"77",X"07",X"DD",X"34",X"02",X"DD",X"7E",X"02",X"FE",X"10",X"C0",
		X"DD",X"36",X"02",X"00",X"DD",X"34",X"00",X"C9",X"40",X"40",X"60",X"50",X"60",X"40",X"70",X"30",
		X"90",X"30",X"A0",X"40",X"A0",X"50",X"C0",X"40",X"DD",X"36",X"05",X"12",X"DD",X"36",X"06",X"01",
		X"DD",X"36",X"0C",X"00",X"D9",X"78",X"D9",X"CB",X"07",X"CB",X"07",X"CB",X"07",X"CB",X"07",X"C6",
		X"40",X"DD",X"77",X"0D",X"DD",X"34",X"00",X"C9",X"CD",X"53",X"37",X"CB",X"07",X"4F",X"06",X"00",
		X"21",X"00",X"3E",X"09",X"5E",X"23",X"56",X"DD",X"7E",X"04",X"83",X"DD",X"77",X"04",X"DD",X"7E",
		X"07",X"82",X"DD",X"77",X"07",X"DD",X"34",X"0C",X"DD",X"7E",X"0C",X"FE",X"40",X"C2",X"84",X"2F",
		X"DD",X"36",X"0C",X"00",X"DD",X"35",X"0D",X"C0",X"DD",X"34",X"00",X"C9",X"DD",X"7E",X"04",X"FE",
		X"80",X"D2",X"9A",X"2F",X"DD",X"35",X"04",X"C3",X"9D",X"2F",X"DD",X"34",X"04",X"CD",X"6A",X"37",
		X"DD",X"7E",X"04",X"FE",X"E8",X"CA",X"B6",X"2F",X"FE",X"18",X"CA",X"B6",X"2F",X"DD",X"7E",X"07",
		X"FE",X"78",X"D2",X"B6",X"2F",X"C9",X"DD",X"36",X"0D",X"05",X"DD",X"34",X"00",X"C9",X"DD",X"35",
		X"0D",X"C0",X"3A",X"02",X"42",X"DD",X"46",X"04",X"90",X"C3",X"49",X"36",X"00",X"00",X"00",X"DD",
		X"34",X"11",X"CB",X"2F",X"CB",X"2F",X"CB",X"2F",X"CB",X"2F",X"00",X"00",X"DD",X"77",X"10",X"DD",
		X"34",X"00",X"C9",X"DD",X"34",X"07",X"DD",X"34",X"07",X"DD",X"7E",X"10",X"DD",X"CB",X"11",X"46",
		X"C2",X"F5",X"2F",X"00",X"00",X"DD",X"86",X"04",X"C3",X"33",X"1E",X"DD",X"7E",X"07",X"FE",X"70",
		X"D8",X"DD",X"36",X"0C",X"00",X"DD",X"34",X"00",X"C9",X"CD",X"53",X"37",X"CB",X"07",X"4F",X"06",
		X"00",X"21",X"80",X"3E",X"09",X"5E",X"23",X"56",X"7B",X"DD",X"CB",X"11",X"46",X"C2",X"22",X"30",
		X"ED",X"44",X"5F",X"DD",X"7E",X"04",X"83",X"DD",X"77",X"04",X"DD",X"7E",X"07",X"82",X"CD",X"70",
		X"36",X"DD",X"7E",X"04",X"FE",X"F0",X"D2",X"3C",X"30",X"FE",X"10",X"D0",X"C3",X"26",X"1E",X"00",
		X"C9",X"DD",X"21",X"A0",X"42",X"11",X"20",X"00",X"06",X"08",X"D9",X"CD",X"5D",X"30",X"D9",X"DD",
		X"19",X"10",X"F7",X"CD",X"58",X"32",X"CD",X"02",X"34",X"CD",X"60",X"2E",X"C9",X"CD",X"9B",X"2E",
		X"DD",X"7E",X"00",X"EF",X"AC",X"2E",X"C8",X"2E",X"72",X"30",X"B1",X"30",X"D1",X"31",X"FF",X"FF",
		X"FF",X"FF",X"DD",X"36",X"05",X"0E",X"DD",X"36",X"06",X"02",X"D9",X"78",X"D9",X"E6",X"01",X"DD",
		X"77",X"09",X"21",X"00",X"3C",X"DD",X"75",X"0A",X"DD",X"74",X"0B",X"D9",X"78",X"D9",X"CB",X"07",
		X"CB",X"07",X"CB",X"07",X"CB",X"07",X"DD",X"77",X"0C",X"DD",X"36",X"0D",X"50",X"CD",X"D1",X"38",
		X"00",X"DD",X"36",X"0F",X"05",X"DD",X"36",X"12",X"00",X"DD",X"36",X"13",X"00",X"DD",X"34",X"00",
		X"C9",X"C3",X"8C",X"36",X"DD",X"34",X"0C",X"DD",X"34",X"0C",X"4F",X"06",X"00",X"DD",X"7E",X"0C",
		X"A7",X"C2",X"CC",X"30",X"DD",X"7E",X"0B",X"EE",X"01",X"DD",X"77",X"0B",X"DD",X"6E",X"0A",X"DD",
		X"66",X"0B",X"09",X"5E",X"23",X"56",X"DD",X"73",X"10",X"DD",X"72",X"11",X"3A",X"A9",X"43",X"FE",
		X"02",X"CA",X"0C",X"31",X"DD",X"7E",X"0C",X"CB",X"0F",X"0F",X"0F",X"DD",X"CB",X"0C",X"7E",X"C3",
		X"F4",X"30",X"EE",X"0F",X"E6",X"07",X"47",X"CB",X"07",X"CB",X"07",X"CB",X"07",X"E6",X"C0",X"4F",
		X"78",X"E6",X"07",X"B1",X"C6",X"28",X"DD",X"77",X"05",X"C3",X"1F",X"31",X"DD",X"7E",X"0C",X"CB",
		X"0F",X"CB",X"0F",X"CB",X"0F",X"D9",X"80",X"D9",X"E6",X"01",X"C6",X"0E",X"C3",X"B6",X"39",X"DD",
		X"CB",X"09",X"46",X"CA",X"2E",X"31",X"DD",X"7E",X"10",X"ED",X"44",X"DD",X"77",X"10",X"DD",X"CB",
		X"12",X"46",X"CA",X"3D",X"31",X"DD",X"7E",X"10",X"ED",X"44",X"DD",X"77",X"10",X"DD",X"7E",X"10",
		X"DD",X"86",X"04",X"F5",X"00",X"00",X"DD",X"CB",X"13",X"46",X"CA",X"55",X"31",X"DD",X"7E",X"11",
		X"ED",X"44",X"DD",X"77",X"11",X"DD",X"7E",X"11",X"DD",X"86",X"07",X"FE",X"20",X"DA",X"6B",X"31",
		X"FE",X"B0",X"D2",X"6B",X"31",X"DD",X"77",X"07",X"C3",X"73",X"31",X"DD",X"7E",X"13",X"EE",X"01",
		X"DD",X"77",X"13",X"F1",X"FE",X"D0",X"30",X"0B",X"FE",X"30",X"38",X"07",X"DD",X"77",X"04",X"C3",
		X"8B",X"31",X"00",X"DD",X"7E",X"12",X"EE",X"01",X"DD",X"77",X"12",X"DD",X"35",X"0D",X"C0",X"DD",
		X"36",X"0D",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"3A",X"0D",X"40",X"4F",X"06",X"00",X"21",X"AA",X"43",X"09",X"7E",X"FE",X"03",
		X"D0",X"C3",X"FD",X"1E",X"00",X"FD",X"36",X"06",X"05",X"FD",X"36",X"14",X"01",X"C3",X"9E",X"1E",
		X"C9",X"00",X"00",X"00",X"00",X"DD",X"34",X"07",X"00",X"DD",X"34",X"07",X"DD",X"7E",X"07",X"FE",
		X"B0",X"D8",X"DD",X"36",X"18",X"01",X"DD",X"36",X"17",X"03",X"00",X"00",X"00",X"DD",X"36",X"08",
		X"01",X"D9",X"78",X"D9",X"E6",X"03",X"DD",X"77",X"16",X"DD",X"36",X"05",X"20",X"DD",X"36",X"06",
		X"05",X"DD",X"36",X"07",X"E8",X"D9",X"78",X"D9",X"CB",X"07",X"CB",X"07",X"CB",X"07",X"CB",X"07",
		X"DD",X"86",X"16",X"DD",X"77",X"15",X"00",X"DD",X"36",X"00",X"00",X"C9",X"DD",X"21",X"A0",X"42",
		X"11",X"20",X"00",X"06",X"08",X"D9",X"CD",X"38",X"32",X"D9",X"DD",X"19",X"10",X"F7",X"CD",X"58",
		X"32",X"CD",X"02",X"34",X"CD",X"60",X"2E",X"C9",X"CD",X"9B",X"2E",X"DD",X"7E",X"00",X"EF",X"AC",
		X"2E",X"C8",X"2E",X"4D",X"32",X"B1",X"30",X"D1",X"31",X"FF",X"FF",X"FF",X"FF",X"DD",X"36",X"05",
		X"28",X"DD",X"36",X"06",X"04",X"C3",X"7A",X"30",X"21",X"AC",X"43",X"35",X"C3",X"C2",X"25",X"3A",
		X"0D",X"40",X"4F",X"06",X"00",X"21",X"AA",X"43",X"09",X"7E",X"A7",X"C8",X"DD",X"21",X"A0",X"42",
		X"11",X"20",X"00",X"06",X"08",X"D9",X"CD",X"7F",X"32",X"D9",X"DD",X"19",X"10",X"F7",X"C9",X"DD",
		X"7E",X"08",X"A7",X"C8",X"DD",X"6E",X"15",X"DD",X"66",X"16",X"45",X"7C",X"CB",X"0F",X"CB",X"0F",
		X"CB",X"0F",X"E6",X"60",X"4F",X"7D",X"CB",X"0F",X"CB",X"0F",X"CB",X"0F",X"E6",X"1F",X"B1",X"5F",
		X"16",X"00",X"21",X"80",X"3F",X"19",X"4E",X"78",X"E6",X"07",X"47",X"3E",X"01",X"05",X"FA",X"B6",
		X"32",X"CB",X"07",X"C3",X"AD",X"32",X"A1",X"C3",X"D7",X"25",X"DD",X"7E",X"04",X"FE",X"E0",X"D2",
		X"ED",X"25",X"DD",X"34",X"04",X"DD",X"34",X"04",X"C3",X"D9",X"32",X"DD",X"7E",X"04",X"FE",X"20",
		X"DA",X"F8",X"25",X"DD",X"35",X"04",X"DD",X"35",X"04",X"DD",X"7E",X"04",X"CB",X"0F",X"E6",X"03",
		X"4F",X"06",X"00",X"21",X"53",X"33",X"09",X"7E",X"DD",X"77",X"05",X"79",X"FE",X"00",X"C2",X"2C",
		X"33",X"CD",X"22",X"39",X"DD",X"7E",X"17",X"E6",X"0F",X"C2",X"2C",X"33",X"3A",X"02",X"42",X"E6",
		X"01",X"C6",X"01",X"CD",X"2B",X"39",X"DD",X"7E",X"04",X"E6",X"F8",X"21",X"FC",X"4F",X"5F",X"16",
		X"00",X"19",X"19",X"19",X"19",X"36",X"5F",X"3A",X"02",X"42",X"DD",X"96",X"04",X"C6",X"0A",X"FE",
		X"15",X"D2",X"3D",X"33",X"3A",X"00",X"42",X"32",X"04",X"42",X"18",X"11",X"DD",X"7E",X"04",X"E6",
		X"F8",X"21",X"FC",X"4F",X"5F",X"16",X"00",X"19",X"19",X"19",X"C3",X"DD",X"38",X"DD",X"6E",X"15",
		X"DD",X"66",X"16",X"23",X"CB",X"54",X"CA",X"4C",X"33",X"21",X"00",X"00",X"DD",X"75",X"15",X"DD",
		X"74",X"16",X"C9",X"21",X"20",X"22",X"20",X"3A",X"A9",X"43",X"A7",X"C8",X"DD",X"21",X"A0",X"42",
		X"11",X"20",X"00",X"06",X"08",X"D9",X"CD",X"6F",X"33",X"D9",X"DD",X"19",X"10",X"F7",X"C9",X"DD",
		X"7E",X"00",X"FE",X"03",X"D8",X"DD",X"7E",X"08",X"A7",X"C0",X"DD",X"CB",X"18",X"46",X"C0",X"DD",
		X"6E",X"19",X"DD",X"66",X"1A",X"7C",X"E6",X"00",X"67",X"2B",X"DD",X"75",X"19",X"DD",X"74",X"1A",
		X"7C",X"B5",X"C0",X"DD",X"7E",X"15",X"E6",X"30",X"CB",X"0F",X"47",X"3A",X"1C",X"42",X"CB",X"07",
		X"CB",X"07",X"CB",X"07",X"E6",X"70",X"4F",X"3A",X"02",X"42",X"E6",X"03",X"CB",X"07",X"CB",X"07",
		X"CB",X"07",X"CB",X"07",X"C6",X"80",X"91",X"80",X"C3",X"43",X"1E",X"DD",X"36",X"1A",X"00",X"DD",
		X"7E",X"07",X"FE",X"60",X"D8",X"FE",X"A0",X"D0",X"11",X"05",X"00",X"21",X"60",X"42",X"06",X"07",
		X"CB",X"46",X"CA",X"D9",X"33",X"19",X"10",X"F8",X"C9",X"36",X"01",X"23",X"DD",X"7E",X"07",X"77",
		X"3E",X"F0",X"96",X"57",X"23",X"23",X"CD",X"0C",X"26",X"77",X"23",X"3A",X"02",X"42",X"DD",X"96",
		X"04",X"DA",X"F9",X"33",X"CD",X"FF",X"11",X"77",X"C9",X"ED",X"44",X"CD",X"FF",X"11",X"ED",X"44",
		X"77",X"C9",X"2A",X"AD",X"43",X"23",X"22",X"AD",X"43",X"CB",X"4C",X"CA",X"4E",X"34",X"21",X"00",
		X"00",X"22",X"AD",X"43",X"CD",X"B6",X"10",X"FE",X"01",X"D8",X"C3",X"00",X"1E",X"00",X"11",X"20",
		X"00",X"06",X"08",X"D9",X"CD",X"2D",X"34",X"D9",X"DD",X"19",X"10",X"F7",X"C9",X"DD",X"CB",X"18",
		X"46",X"C8",X"DD",X"CB",X"1B",X"46",X"C0",X"DD",X"CB",X"08",X"46",X"C0",X"DD",X"36",X"05",X"15",
		X"DD",X"36",X"06",X"00",X"DD",X"36",X"1F",X"01",X"CD",X"3D",X"37",X"00",X"F1",X"C9",X"DD",X"2A",
		X"AF",X"43",X"DD",X"7E",X"1F",X"FE",X"01",X"C0",X"CB",X"44",X"C3",X"9A",X"36",X"DD",X"7E",X"0C",
		X"FE",X"40",X"DA",X"6C",X"34",X"DD",X"36",X"0C",X"00",X"C3",X"6F",X"34",X"DD",X"34",X"0C",X"DD",
		X"7E",X"0C",X"4F",X"06",X"00",X"21",X"00",X"3F",X"09",X"09",X"7E",X"DD",X"77",X"04",X"23",X"7E",
		X"DD",X"77",X"07",X"C9",X"C3",X"A4",X"36",X"00",X"C9",X"21",X"A4",X"42",X"11",X"60",X"40",X"06",
		X"08",X"7E",X"ED",X"44",X"12",X"23",X"13",X"7E",X"12",X"23",X"13",X"7E",X"12",X"23",X"13",X"7E",
		X"00",X"00",X"12",X"13",X"C5",X"01",X"1D",X"00",X"09",X"C1",X"05",X"C2",X"91",X"34",X"3A",X"08",
		X"42",X"0F",X"D0",X"DD",X"21",X"A0",X"42",X"11",X"20",X"00",X"06",X"08",X"D9",X"CD",X"C6",X"34",
		X"D9",X"DD",X"19",X"10",X"F7",X"C9",X"DD",X"CB",X"18",X"46",X"CA",X"D2",X"34",X"DD",X"CB",X"1F",
		X"46",X"C8",X"DD",X"CB",X"1B",X"46",X"C0",X"DD",X"CB",X"08",X"46",X"C0",X"3A",X"A9",X"43",X"A7",
		X"C8",X"DD",X"7E",X"00",X"FE",X"03",X"D8",X"2A",X"09",X"42",X"DD",X"7E",X"07",X"95",X"C6",X"18",
		X"FE",X"0C",X"D0",X"DD",X"7E",X"04",X"94",X"C6",X"00",X"FE",X"10",X"D0",X"3E",X"01",X"32",X"0B",
		X"42",X"3A",X"A9",X"43",X"FE",X"03",X"C2",X"2C",X"35",X"DD",X"7E",X"00",X"FE",X"03",X"C3",X"30",
		X"37",X"DD",X"7E",X"04",X"94",X"C6",X"FE",X"FE",X"04",X"D0",X"DD",X"7E",X"05",X"E6",X"3F",X"FE",
		X"28",X"C8",X"00",X"00",X"FE",X"2C",X"00",X"00",X"00",X"00",X"00",X"C8",X"C3",X"EF",X"38",X"00",
		X"DD",X"36",X"1B",X"01",X"C3",X"BD",X"36",X"00",X"C9",X"DD",X"21",X"A0",X"42",X"11",X"20",X"00",
		X"06",X"08",X"D9",X"CD",X"4C",X"35",X"D9",X"DD",X"19",X"10",X"F7",X"C9",X"C3",X"90",X"1F",X"00",
		X"C8",X"DD",X"7E",X"1C",X"EF",X"5B",X"35",X"9A",X"35",X"FF",X"FF",X"DD",X"36",X"1D",X"04",X"DD",
		X"36",X"1E",X"04",X"DD",X"36",X"05",X"1C",X"DD",X"34",X"1C",X"DD",X"CB",X"1F",X"46",X"CA",X"7B",
		X"35",X"00",X"00",X"00",X"00",X"11",X"05",X"03",X"C3",X"1C",X"1E",X"3A",X"A9",X"43",X"FE",X"01",
		X"CA",X"91",X"35",X"DD",X"7E",X"00",X"FE",X"04",X"C3",X"EB",X"36",X"11",X"04",X"03",X"C3",X"F2",
		X"08",X"3A",X"A9",X"43",X"5F",X"16",X"03",X"C3",X"F2",X"08",X"DD",X"35",X"1D",X"C0",X"DD",X"36",
		X"1D",X"04",X"DD",X"34",X"05",X"DD",X"35",X"1E",X"C0",X"DD",X"36",X"1B",X"00",X"C3",X"1C",X"37",
		X"FE",X"02",X"CA",X"BA",X"35",X"FE",X"03",X"C2",X"E7",X"35",X"DD",X"7E",X"00",X"FE",X"03",X"C2",
		X"E7",X"35",X"3A",X"0D",X"40",X"4F",X"06",X"00",X"21",X"AA",X"43",X"09",X"7E",X"FE",X"03",X"C3",
		X"69",X"2D",X"DD",X"36",X"05",X"20",X"DD",X"36",X"06",X"05",X"DD",X"36",X"14",X"01",X"DD",X"36",
		X"00",X"04",X"DD",X"36",X"18",X"00",X"C9",X"DD",X"36",X"04",X"FF",X"DD",X"36",X"07",X"FF",X"C3",
		X"15",X"18",X"00",X"C9",X"3A",X"0D",X"40",X"4F",X"06",X"00",X"21",X"A1",X"43",X"09",X"36",X"01",
		X"00",X"00",X"00",X"00",X"00",X"C9",X"00",X"00",X"3A",X"0D",X"40",X"4F",X"06",X"00",X"21",X"A1",
		X"43",X"09",X"7E",X"A7",X"C3",X"A2",X"38",X"CD",X"37",X"08",X"C3",X"64",X"06",X"CD",X"37",X"08",
		X"CD",X"98",X"08",X"CD",X"74",X"0A",X"CD",X"32",X"0A",X"CD",X"5E",X"0B",X"CD",X"E5",X"08",X"CD",
		X"D4",X"12",X"CD",X"0E",X"13",X"00",X"00",X"00",X"C3",X"00",X"2D",X"22",X"0D",X"40",X"21",X"A0",
		X"43",X"AF",X"06",X"10",X"77",X"23",X"10",X"FC",X"C9",X"DD",X"36",X"11",X"00",X"D2",X"D2",X"2F",
		X"C3",X"CD",X"2F",X"DD",X"21",X"A0",X"42",X"11",X"20",X"00",X"06",X"08",X"AF",X"DD",X"B6",X"1B",
		X"DD",X"19",X"10",X"F9",X"CB",X"47",X"C0",X"C3",X"7B",X"2E",X"3A",X"02",X"42",X"C6",X"80",X"C9",
		X"DD",X"77",X"07",X"DD",X"34",X"0C",X"DD",X"7E",X"0C",X"FE",X"40",X"C2",X"82",X"36",X"DD",X"36",
		X"0C",X"00",X"C9",X"DD",X"7E",X"05",X"FE",X"24",X"C8",X"C3",X"AA",X"2E",X"DD",X"35",X"0F",X"C0",
		X"DD",X"36",X"0F",X"05",X"DD",X"7E",X"0C",X"C3",X"B4",X"30",X"C2",X"84",X"34",X"7D",X"E6",X"03",
		X"C0",X"C3",X"5D",X"34",X"DD",X"36",X"1F",X"00",X"DD",X"36",X"04",X"FF",X"DD",X"36",X"07",X"FF",
		X"C9",X"DD",X"34",X"00",X"34",X"C9",X"D2",X"E7",X"35",X"34",X"C3",X"D2",X"35",X"DD",X"36",X"1C",
		X"00",X"DD",X"CB",X"1F",X"46",X"C8",X"CD",X"80",X"26",X"00",X"11",X"20",X"00",X"06",X"08",X"DD",
		X"CB",X"08",X"46",X"CA",X"BB",X"15",X"CD",X"9A",X"26",X"00",X"DD",X"19",X"10",X"F1",X"3A",X"0D",
		X"40",X"4F",X"06",X"00",X"21",X"AA",X"43",X"09",X"C3",X"12",X"26",X"C2",X"91",X"35",X"3A",X"0D",
		X"40",X"4F",X"06",X"00",X"21",X"AA",X"43",X"09",X"35",X"C3",X"8B",X"35",X"32",X"BF",X"43",X"DD",
		X"36",X"04",X"FF",X"DD",X"36",X"07",X"FF",X"DD",X"36",X"18",X"01",X"C9",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"00",X"25",X"F9",X"C9",X"DD",X"CB",X"1F",X"46",
		X"C2",X"29",X"37",X"3A",X"A9",X"43",X"C3",X"B0",X"35",X"AF",X"32",X"BF",X"43",X"C3",X"E7",X"35",
		X"C2",X"2C",X"35",X"DD",X"CB",X"1F",X"46",X"C2",X"2C",X"35",X"C3",X"11",X"35",X"DD",X"22",X"AF",
		X"43",X"DD",X"36",X"00",X"03",X"C9",X"DD",X"CB",X"08",X"86",X"DD",X"36",X"04",X"FF",X"DD",X"36",
		X"07",X"FF",X"C9",X"DD",X"7E",X"0C",X"CB",X"0F",X"CB",X"0F",X"CB",X"0F",X"D9",X"80",X"D9",X"E6",
		X"03",X"C6",X"11",X"DD",X"77",X"05",X"DD",X"7E",X"0C",X"C9",X"DD",X"36",X"05",X"12",X"DD",X"34",
		X"07",X"C9",X"C2",X"5B",X"03",X"C3",X"22",X"26",X"00",X"00",X"00",X"3A",X"0D",X"40",X"4F",X"06",
		X"00",X"21",X"A1",X"43",X"09",X"36",X"00",X"CD",X"97",X"38",X"09",X"36",X"00",X"AF",X"32",X"A8",
		X"43",X"C3",X"F3",X"37",X"C9",X"3A",X"08",X"42",X"2A",X"00",X"42",X"B4",X"B5",X"0F",X"D8",X"00",
		X"00",X"00",X"00",X"00",X"21",X"60",X"42",X"11",X"05",X"00",X"06",X"07",X"AF",X"B6",X"19",X"10",
		X"FC",X"0F",X"D8",X"21",X"09",X"40",X"35",X"C0",X"C3",X"68",X"38",X"21",X"00",X"00",X"22",X"AD",
		X"43",X"22",X"A4",X"43",X"AF",X"32",X"A8",X"43",X"32",X"AC",X"43",X"21",X"A0",X"42",X"06",X"00",
		X"36",X"00",X"23",X"10",X"FB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"CD",X"E8",X"37",X"C3",X"4A",X"38",X"C9",X"21",X"60",X"40",X"AF",X"06",X"20",X"77",X"23",
		X"10",X"FC",X"C9",X"32",X"A9",X"43",X"21",X"22",X"42",X"CD",X"28",X"16",X"C3",X"C1",X"38",X"09",
		X"21",X"00",X"00",X"22",X"AF",X"43",X"21",X"A9",X"43",X"34",X"3A",X"0D",X"40",X"4F",X"06",X"00",
		X"21",X"A6",X"43",X"09",X"34",X"C9",X"3A",X"0E",X"40",X"A7",X"20",X"13",X"21",X"00",X"41",X"C9",
		X"3A",X"0D",X"40",X"4F",X"06",X"00",X"21",X"A6",X"43",X"09",X"35",X"21",X"A9",X"43",X"C9",X"3A",
		X"0D",X"40",X"4F",X"06",X"00",X"21",X"A1",X"43",X"09",X"7E",X"A7",X"CA",X"1C",X"38",X"21",X"00",
		X"41",X"AF",X"06",X"10",X"77",X"23",X"10",X"FC",X"18",X"3E",X"3A",X"0E",X"40",X"A7",X"CA",X"64",
		X"38",X"3A",X"0D",X"40",X"EE",X"00",X"4F",X"06",X"00",X"21",X"A1",X"43",X"09",X"7E",X"A7",X"CA",
		X"64",X"38",X"18",X"24",X"21",X"00",X"41",X"C9",X"2C",X"34",X"21",X"00",X"00",X"22",X"AD",X"43",
		X"22",X"A4",X"43",X"AF",X"32",X"A8",X"43",X"32",X"AC",X"43",X"CD",X"0A",X"2D",X"06",X"00",X"36",
		X"00",X"23",X"10",X"FB",X"CD",X"E8",X"37",X"C9",X"EB",X"11",X"10",X"00",X"19",X"EB",X"F1",X"C9",
		X"ED",X"B0",X"AF",X"32",X"0D",X"40",X"C9",X"21",X"A6",X"43",X"09",X"36",X"00",X"21",X"AA",X"43",
		X"09",X"C9",X"C2",X"AC",X"38",X"AF",X"32",X"02",X"60",X"C3",X"17",X"36",X"3E",X"01",X"32",X"02",
		X"60",X"C3",X"1D",X"36",X"DD",X"36",X"02",X"00",X"DD",X"36",X"04",X"00",X"DD",X"36",X"07",X"00",
		X"C9",X"21",X"1C",X"50",X"06",X"20",X"11",X"20",X"00",X"36",X"10",X"19",X"10",X"FB",X"C3",X"E8",
		X"37",X"3A",X"02",X"42",X"D9",X"80",X"D9",X"E6",X"07",X"DD",X"77",X"0E",X"C9",X"19",X"36",X"5E",
		X"11",X"E0",X"FF",X"19",X"36",X"5E",X"11",X"40",X"00",X"19",X"36",X"5E",X"C3",X"3D",X"33",X"DD",
		X"7E",X"05",X"FE",X"15",X"C2",X"FF",X"38",X"21",X"B9",X"43",X"36",X"20",X"C3",X"1B",X"39",X"FE",
		X"20",X"C2",X"0D",X"39",X"21",X"B9",X"43",X"36",X"08",X"C3",X"1B",X"39",X"00",X"3A",X"A9",X"43",
		X"FE",X"03",X"C2",X"17",X"39",X"3E",X"04",X"21",X"B9",X"43",X"77",X"DD",X"36",X"18",X"01",X"C3",
		X"30",X"35",X"DD",X"35",X"17",X"21",X"B9",X"43",X"36",X"10",X"C9",X"DD",X"77",X"17",X"21",X"B9",
		X"43",X"36",X"40",X"C9",X"32",X"03",X"68",X"32",X"08",X"42",X"C9",X"32",X"41",X"42",X"21",X"4A",
		X"39",X"11",X"60",X"40",X"01",X"18",X"00",X"ED",X"B0",X"C9",X"40",X"20",X"00",X"64",X"40",X"21",
		X"01",X"7C",X"40",X"22",X"02",X"94",X"40",X"23",X"04",X"AC",X"40",X"26",X"05",X"C4",X"40",X"27",
		X"00",X"DC",X"3A",X"41",X"42",X"C6",X"4B",X"5F",X"16",X"06",X"C3",X"F2",X"08",X"3A",X"08",X"42",
		X"2A",X"00",X"42",X"B4",X"B5",X"0F",X"DA",X"92",X"39",X"3A",X"25",X"42",X"0F",X"D2",X"92",X"39",
		X"21",X"60",X"42",X"11",X"05",X"00",X"06",X"07",X"AF",X"B6",X"19",X"10",X"FC",X"0F",X"DA",X"92",
		X"39",X"C9",X"21",X"01",X"00",X"C3",X"1A",X"16",X"AF",X"32",X"02",X"60",X"CD",X"B6",X"1F",X"C9",
		X"AF",X"32",X"02",X"60",X"CD",X"90",X"27",X"C9",X"AF",X"32",X"0A",X"42",X"C3",X"F2",X"08",X"32",
		X"01",X"60",X"32",X"02",X"60",X"C9",X"DD",X"77",X"05",X"DD",X"7E",X"10",X"07",X"DD",X"77",X"10",
		X"C3",X"1F",X"31",X"D9",X"21",X"A5",X"43",X"AE",X"E6",X"07",X"C9",X"D9",X"78",X"D9",X"07",X"07",
		X"07",X"07",X"47",X"7D",X"B8",X"D8",X"C3",X"BC",X"2E",X"3A",X"0D",X"40",X"4F",X"06",X"00",X"21",
		X"C0",X"43",X"09",X"36",X"10",X"C3",X"03",X"26",X"3A",X"0D",X"40",X"5F",X"16",X"00",X"21",X"C2",
		X"43",X"19",X"19",X"19",X"11",X"E0",X"FF",X"C9",X"DD",X"77",X"04",X"23",X"CD",X"E2",X"31",X"C9",
		X"00",X"00",X"00",X"00",X"00",X"3A",X"07",X"40",X"0F",X"D8",X"AF",X"32",X"B8",X"43",X"3A",X"B9",
		X"43",X"CB",X"67",X"C4",X"65",X"3A",X"3A",X"B9",X"43",X"CB",X"47",X"3E",X"00",X"CD",X"60",X"27",
		X"00",X"CB",X"4F",X"3E",X"01",X"CD",X"60",X"27",X"00",X"CB",X"57",X"3E",X"02",X"CD",X"60",X"27",
		X"00",X"CB",X"5F",X"3E",X"03",X"CD",X"60",X"27",X"00",X"CB",X"6F",X"C3",X"40",X"27",X"CB",X"77",
		X"C4",X"A6",X"3A",X"C3",X"EE",X"27",X"00",X"00",X"3A",X"B8",X"43",X"32",X"06",X"68",X"0F",X"32",
		X"07",X"68",X"2A",X"BA",X"43",X"7E",X"32",X"00",X"78",X"23",X"22",X"BA",X"43",X"7E",X"A7",X"C0",
		X"C3",X"F5",X"27",X"00",X"00",X"21",X"68",X"3B",X"22",X"BA",X"43",X"3A",X"B9",X"43",X"CB",X"A7",
		X"32",X"B9",X"43",X"3E",X"02",X"CD",X"E5",X"27",X"C9",X"21",X"18",X"3B",X"85",X"5E",X"23",X"56",
		X"EB",X"22",X"BA",X"43",X"3A",X"B9",X"43",X"E6",X"F0",X"32",X"B9",X"43",X"3E",X"02",X"CD",X"E5",
		X"27",X"C9",X"21",X"19",X"3B",X"22",X"BA",X"43",X"3A",X"B9",X"43",X"CB",X"AF",X"32",X"B9",X"43",
		X"3E",X"02",X"CD",X"E5",X"27",X"C9",X"21",X"58",X"3B",X"22",X"BA",X"43",X"3A",X"B9",X"43",X"CB",
		X"B7",X"32",X"B9",X"43",X"3E",X"02",X"CD",X"E5",X"27",X"C9",X"3A",X"BD",X"43",X"5E",X"C3",X"50",
		X"27",X"00",X"00",X"00",X"21",X"20",X"3B",X"16",X"00",X"19",X"46",X"21",X"00",X"68",X"CB",X"40",
		X"CC",X"0A",X"3B",X"C4",X"11",X"3B",X"CB",X"48",X"CC",X"0A",X"3B",X"C4",X"11",X"3B",X"CB",X"50",
		X"CC",X"0A",X"3B",X"C4",X"11",X"3B",X"21",X"04",X"60",X"CB",X"58",X"CC",X"0A",X"3B",X"C4",X"11",
		X"3B",X"CB",X"60",X"CC",X"0A",X"3B",X"C4",X"11",X"3B",X"CB",X"68",X"CC",X"0A",X"3B",X"C4",X"11",
		X"3B",X"CB",X"70",X"CC",X"0A",X"3B",X"C4",X"11",X"3B",X"C9",X"F5",X"3E",X"00",X"77",X"23",X"F1",
		X"C9",X"F5",X"3E",X"01",X"77",X"23",X"F1",X"C9",X"95",X"3B",X"B0",X"3B",X"E0",X"3B",X"40",X"3E",
		X"00",X"32",X"22",X"15",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"E0",X"E1",X"DC",X"F0",X"F1",X"EE",X"EF",X"EB",X"EC",X"E9",X"EA",X"E6",X"E7",X"E4",X"E5",X"E2",
		X"E3",X"E1",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"CE",X"C3",X"CE",X"C3",X"CE",X"C3",X"CE",X"C3",
		X"CE",X"C3",X"CE",X"C0",X"00",X"FF",X"FF",X"FF",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",
		X"E1",X"FF",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"00",X"FF",X"FF",X"E0",X"E1",X"DC",X"F0",
		X"F1",X"EE",X"EB",X"EC",X"E9",X"EA",X"E6",X"E7",X"E4",X"E5",X"E2",X"E3",X"E1",X"E0",X"E1",X"DC",
		X"F0",X"F1",X"EE",X"EF",X"00",X"80",X"70",X"D0",X"8E",X"E0",X"87",X"55",X"FF",X"FF",X"40",X"68",
		X"70",X"DC",X"D5",X"CD",X"CD",X"8E",X"8F",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"E0",X"E0",X"E0",X"D1",X"D1",X"D1",X"E0",X"E0",X"E0",X"D1",X"D1",X"D1",X"E0",X"E0",X"E0",X"D1",
		X"D1",X"D1",X"E0",X"E0",X"E0",X"D1",X"D1",X"D1",X"E0",X"E0",X"E0",X"D1",X"D1",X"D1",X"E0",X"E0",
		X"E0",X"D1",X"D1",X"D1",X"E0",X"E0",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"DC",X"DC",X"DC",X"DC",X"DC",X"DC",X"E0",X"E0",X"DC",X"DC",X"D1",X"C0",X"C2",X"C1",X"C3",X"C4",
		X"C2",X"C0",X"C3",X"C2",X"C2",X"C2",X"C2",X"C2",X"C2",X"C2",X"C2",X"00",X"FF",X"FF",X"FF",X"FF",
		X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"01",X"01",X"02",X"00",X"02",X"00",X"01",X"01",
		X"02",X"00",X"02",X"01",X"02",X"01",X"02",X"01",X"02",X"01",X"02",X"02",X"02",X"01",X"02",X"02",
		X"02",X"02",X"02",X"02",X"01",X"02",X"02",X"02",X"01",X"02",X"01",X"02",X"01",X"02",X"01",X"02",
		X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"01",X"01",X"00",X"02",X"00",X"02",X"00",X"02",
		X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"FF",X"01",X"00",X"02",X"00",X"02",X"FF",X"01",
		X"00",X"02",X"FF",X"02",X"FF",X"02",X"FF",X"02",X"FF",X"02",X"FF",X"02",X"FF",X"02",X"FE",X"02",
		X"FE",X"02",X"FE",X"02",X"FE",X"01",X"FE",X"01",X"FE",X"01",X"FE",X"01",X"FE",X"01",X"FE",X"01",
		X"FE",X"00",X"FF",X"00",X"FE",X"00",X"FE",X"00",X"FF",X"01",X"FE",X"00",X"FE",X"00",X"FE",X"00",
		X"FE",X"00",X"FE",X"00",X"FE",X"00",X"FE",X"00",X"FF",X"FF",X"FE",X"00",X"FE",X"00",X"FF",X"FF",
		X"FE",X"00",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FE",X"FE",X"FF",X"FE",X"FE",
		X"FE",X"FE",X"FE",X"FE",X"FF",X"FE",X"FE",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",
		X"00",X"FE",X"FF",X"FF",X"00",X"FE",X"00",X"FE",X"FF",X"FF",X"00",X"FE",X"00",X"FE",X"00",X"FE",
		X"00",X"FE",X"00",X"FE",X"00",X"FE",X"00",X"FE",X"01",X"FF",X"00",X"FE",X"00",X"FE",X"01",X"FF",
		X"00",X"FE",X"01",X"FE",X"01",X"FE",X"01",X"FE",X"01",X"FE",X"02",X"FE",X"01",X"FE",X"02",X"FF",
		X"02",X"FE",X"02",X"FE",X"02",X"FF",X"02",X"FE",X"02",X"FF",X"02",X"FF",X"02",X"FF",X"02",X"FF",
		X"02",X"00",X"01",X"FF",X"02",X"00",X"02",X"00",X"01",X"FF",X"02",X"00",X"02",X"00",X"02",X"00",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"03",X"02",X"03",X"02",X"02",X"01",X"03",X"01",
		X"03",X"01",X"03",X"00",X"03",X"01",X"03",X"00",X"03",X"00",X"04",X"00",X"04",X"00",X"02",X"02",
		X"FD",X"02",X"FD",X"01",X"FD",X"01",X"FD",X"01",X"FD",X"01",X"FD",X"01",X"FD",X"01",X"FD",X"01",
		X"FD",X"01",X"FD",X"01",X"FD",X"00",X"FD",X"00",X"00",X"03",X"00",X"04",X"00",X"03",X"FD",X"02",
		X"FD",X"01",X"FD",X"01",X"FC",X"01",X"FC",X"01",X"FC",X"00",X"FC",X"00",X"02",X"02",X"02",X"03",
		X"03",X"02",X"03",X"02",X"03",X"01",X"04",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"02",X"FF",
		X"02",X"FE",X"03",X"00",X"03",X"02",X"02",X"02",X"02",X"02",X"03",X"02",X"03",X"01",X"04",X"01",
		X"04",X"00",X"03",X"01",X"FE",X"02",X"FC",X"02",X"FC",X"02",X"FC",X"02",X"FC",X"01",X"FC",X"01",
		X"FC",X"01",X"FC",X"01",X"FC",X"00",X"FC",X"02",X"FC",X"02",X"FD",X"02",X"FD",X"02",X"FD",X"02",
		X"FC",X"02",X"FD",X"01",X"FC",X"00",X"00",X"04",X"00",X"04",X"00",X"04",X"02",X"02",X"03",X"02",
		X"02",X"02",X"03",X"02",X"03",X"03",X"03",X"03",X"03",X"01",X"05",X"01",X"05",X"00",X"04",X"00",
		X"04",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"05",X"00",X"05",X"00",X"04",X"01",X"04",X"01",
		X"04",X"02",X"03",X"04",X"02",X"04",X"01",X"03",X"01",X"04",X"00",X"04",X"FF",X"04",X"FD",X"04",
		X"FD",X"02",X"FD",X"01",X"FD",X"01",X"FD",X"00",X"FD",X"FF",X"FD",X"FF",X"FC",X"00",X"FD",X"02",
		X"FD",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"FD",X"04",X"FD",X"02",X"FD",X"03",
		X"FD",X"03",X"FD",X"03",X"FD",X"03",X"FD",X"03",X"FD",X"03",X"02",X"03",X"03",X"04",X"02",X"03",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"01",X"FF",X"00",X"FF",X"01",X"FF",X"01",X"FF",X"01",X"00",X"01",
		X"00",X"01",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"01",X"01",X"01",X"00",
		X"01",X"00",X"01",X"00",X"01",X"FF",X"01",X"00",X"01",X"FF",X"01",X"FF",X"01",X"FF",X"01",X"FF",
		X"01",X"FF",X"01",X"FF",X"01",X"FF",X"01",X"FF",X"01",X"FF",X"01",X"00",X"01",X"FF",X"01",X"00",
		X"01",X"00",X"01",X"00",X"01",X"01",X"01",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"01",
		X"00",X"01",X"00",X"01",X"FF",X"01",X"FF",X"01",X"FF",X"01",X"FF",X"00",X"FF",X"01",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FC",X"04",X"FD",X"03",X"FD",X"03",X"FD",X"03",X"FD",X"02",X"FD",X"01",X"FC",X"01",X"FC",X"00",
		X"FC",X"FF",X"FD",X"FE",X"FD",X"FE",X"FE",X"FD",X"FE",X"FD",X"FE",X"FD",X"FE",X"FD",X"FE",X"FC",
		X"00",X"FC",X"01",X"FC",X"04",X"FD",X"04",X"FF",X"04",X"00",X"02",X"02",X"03",X"03",X"02",X"03",
		X"01",X"04",X"00",X"04",X"FE",X"03",X"FE",X"03",X"FD",X"02",X"FD",X"02",X"FD",X"02",X"FD",X"02",
		X"FC",X"03",X"FC",X"03",X"FB",X"02",X"FB",X"02",X"FA",X"02",X"FB",X"01",X"FB",X"02",X"FB",X"02",
		X"FA",X"02",X"FB",X"02",X"FB",X"02",X"FB",X"02",X"FB",X"02",X"FB",X"01",X"FB",X"02",X"FB",X"02",
		X"FA",X"01",X"FA",X"01",X"FA",X"01",X"FA",X"01",X"FA",X"01",X"F9",X"01",X"F9",X"01",X"F9",X"01",
		X"F8",X"01",X"F8",X"01",X"F8",X"00",X"F8",X"00",X"F8",X"00",X"F8",X"00",X"F8",X"00",X"F8",X"00",
		X"D0",X"1F",X"CA",X"1E",X"C5",X"1E",X"C1",X"1F",X"BD",X"21",X"B9",X"24",X"B6",X"27",X"B4",X"2A",
		X"B3",X"2E",X"B3",X"32",X"B4",X"36",X"B6",X"39",X"BA",X"3A",X"BE",X"39",X"C0",X"36",X"CF",X"32",
		X"BB",X"30",X"B7",X"2F",X"B3",X"2E",X"AF",X"2C",X"AB",X"2A",X"A8",X"27",X"A3",X"24",X"9E",X"22",
		X"98",X"21",X"91",X"21",X"89",X"21",X"59",X"21",X"59",X"20",X"59",X"20",X"56",X"20",X"51",X"20",
		X"4D",X"23",X"49",X"26",X"45",X"2A",X"41",X"2E",X"3D",X"32",X"39",X"36",X"35",X"39",X"31",X"3B",
		X"2E",X"3E",X"29",X"40",X"26",X"3D",X"24",X"39",X"26",X"36",X"2A",X"32",X"2F",X"30",X"36",X"30",
		X"3D",X"30",X"45",X"30",X"4D",X"30",X"55",X"30",X"5D",X"30",X"65",X"31",X"6D",X"32",X"75",X"33",
		X"7D",X"34",X"85",X"35",X"CC",X"35",X"D4",X"34",X"DA",X"32",X"DC",X"2D",X"DA",X"28",X"D6",X"23",
		X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"00",X"00",X"00",X"55",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
