library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity defender_sound is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of defender_sound is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"EF",X"0F",X"8E",X"00",X"7F",X"CE",X"84",X"00",X"6F",X"01",X"6F",X"03",X"86",X"FF",X"A7",X"00",
		X"6F",X"02",X"86",X"07",X"A7",X"01",X"A7",X"03",X"97",X"1C",X"7F",X"00",X"20",X"0E",X"20",X"FE",
		X"CE",X"FA",X"D0",X"C6",X"1C",X"BD",X"F9",X"94",X"BD",X"F8",X"EB",X"39",X"CE",X"FA",X"0C",X"C6",
		X"1C",X"BD",X"F9",X"94",X"BD",X"F8",X"EB",X"39",X"CE",X"FA",X"28",X"C6",X"1C",X"BD",X"F9",X"94",
		X"BD",X"F8",X"EB",X"39",X"CE",X"FA",X"44",X"C6",X"1C",X"BD",X"F9",X"94",X"BD",X"F8",X"EB",X"39",
		X"CE",X"FA",X"60",X"C6",X"1C",X"BD",X"F9",X"94",X"BD",X"F8",X"EB",X"39",X"CE",X"FA",X"7C",X"C6",
		X"1C",X"BD",X"F9",X"94",X"BD",X"F8",X"EB",X"39",X"CE",X"FA",X"98",X"C6",X"1C",X"BD",X"F9",X"94",
		X"BD",X"F8",X"EB",X"39",X"CE",X"FA",X"B4",X"C6",X"1C",X"BD",X"F9",X"94",X"BD",X"F8",X"EB",X"39",
		X"CE",X"FB",X"08",X"C6",X"1C",X"BD",X"F9",X"94",X"BD",X"F8",X"EB",X"39",X"CE",X"FB",X"24",X"C6",
		X"1C",X"BD",X"F9",X"94",X"BD",X"F8",X"EB",X"39",X"CE",X"FB",X"40",X"C6",X"1C",X"BD",X"F9",X"94",
		X"BD",X"F8",X"EB",X"CE",X"00",X"00",X"DF",X"22",X"CE",X"FB",X"5C",X"C6",X"1C",X"BD",X"F9",X"94",
		X"BD",X"F8",X"EB",X"39",X"CE",X"FB",X"78",X"C6",X"1C",X"BD",X"F9",X"94",X"BD",X"F8",X"EB",X"39",
		X"CE",X"FA",X"EC",X"C6",X"1C",X"BD",X"F9",X"94",X"BD",X"F8",X"EB",X"39",X"CE",X"00",X"01",X"DF",
		X"00",X"CE",X"10",X"00",X"DF",X"02",X"7F",X"84",X"00",X"DE",X"00",X"08",X"DF",X"00",X"09",X"26",
		X"FD",X"73",X"84",X"00",X"DE",X"02",X"09",X"26",X"FD",X"20",X"EB",X"DF",X"24",X"CE",X"F9",X"90",
		X"DF",X"26",X"86",X"80",X"D6",X"03",X"2A",X"09",X"D6",X"1D",X"54",X"54",X"54",X"5C",X"5A",X"26",
		X"FD",X"7A",X"00",X"08",X"27",X"4C",X"7A",X"00",X"09",X"27",X"4C",X"7A",X"00",X"0A",X"27",X"4C",
		X"7A",X"00",X"0B",X"26",X"DF",X"D6",X"03",X"27",X"DB",X"C4",X"7F",X"D7",X"0B",X"D6",X"1D",X"58",
		X"DB",X"1D",X"CB",X"0B",X"D7",X"1D",X"7A",X"00",X"1B",X"26",X"0E",X"D6",X"0F",X"D7",X"1B",X"DE",
		X"26",X"09",X"8C",X"F9",X"89",X"27",X"4E",X"DF",X"26",X"D6",X"1D",X"2B",X"06",X"D4",X"07",X"C4",
		X"7F",X"20",X"05",X"D4",X"07",X"C4",X"7F",X"50",X"36",X"1B",X"16",X"32",X"DE",X"26",X"AD",X"00",
		X"20",X"A2",X"CE",X"00",X"00",X"20",X"08",X"CE",X"00",X"01",X"20",X"03",X"CE",X"00",X"02",X"6D",
		X"18",X"27",X"12",X"6A",X"18",X"26",X"0E",X"E6",X"0C",X"E7",X"18",X"E6",X"00",X"EB",X"10",X"E1",
		X"14",X"27",X"12",X"E7",X"00",X"E6",X"00",X"E7",X"08",X"AB",X"04",X"60",X"04",X"16",X"DE",X"26",
		X"AD",X"00",X"7E",X"F8",X"F4",X"DE",X"24",X"39",X"54",X"54",X"54",X"54",X"54",X"54",X"54",X"54",
		X"F7",X"84",X"00",X"39",X"36",X"A6",X"00",X"DF",X"24",X"DE",X"22",X"A7",X"00",X"08",X"DF",X"22",
		X"DE",X"24",X"08",X"5A",X"26",X"EF",X"32",X"39",X"8E",X"00",X"7F",X"CE",X"F9",X"90",X"DF",X"26",
		X"B6",X"84",X"02",X"CE",X"00",X"00",X"DF",X"22",X"C6",X"AF",X"D7",X"1E",X"0E",X"84",X"1F",X"27",
		X"16",X"81",X"00",X"23",X"FE",X"81",X"11",X"22",X"FE",X"4A",X"48",X"CE",X"FB",X"94",X"8D",X"0B",
		X"EE",X"00",X"AD",X"00",X"7C",X"00",X"1F",X"96",X"20",X"27",X"FE",X"DF",X"24",X"9B",X"25",X"97",
		X"25",X"96",X"24",X"89",X"00",X"97",X"24",X"DE",X"24",X"39",X"0F",X"CE",X"FF",X"FF",X"5F",X"0C",
		X"E9",X"00",X"09",X"8C",X"F8",X"00",X"26",X"F8",X"E1",X"00",X"27",X"01",X"3E",X"CE",X"F9",X"90",
		X"DF",X"26",X"CE",X"00",X"00",X"DF",X"22",X"BD",X"F8",X"B4",X"20",X"F1",X"00",X"00",X"00",X"40",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"18",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"18",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"60",X"40",X"45",X"00",X"18",X"40",X"40",X"00",X"FF",X"40",X"45",X"00",X"18",
		X"20",X"20",X"00",X"60",X"02",X"05",X"00",X"FF",X"00",X"00",X"00",X"80",X"20",X"20",X"00",X"60",
		X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"70",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"C0",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"01",X"01",X"00",X"00",X"3F",X"3F",X"00",X"00",
		X"01",X"01",X"00",X"00",X"20",X"20",X"00",X"00",X"01",X"02",X"00",X"00",X"31",X"31",X"00",X"00",
		X"20",X"20",X"00",X"00",X"03",X"00",X"00",X"04",X"3F",X"00",X"00",X"3F",X"03",X"00",X"00",X"04",
		X"FF",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"A0",
		X"04",X"01",X"01",X"00",X"1F",X"1F",X"1F",X"00",X"04",X"01",X"01",X"00",X"02",X"02",X"02",X"00",
		X"04",X"02",X"00",X"00",X"40",X"40",X"40",X"00",X"02",X"02",X"02",X"00",X"04",X"01",X"01",X"00",
		X"10",X"10",X"10",X"00",X"04",X"01",X"01",X"00",X"08",X"08",X"FF",X"00",X"04",X"02",X"00",X"00",
		X"AC",X"FF",X"00",X"00",X"08",X"08",X"FF",X"00",X"01",X"01",X"01",X"00",X"1F",X"1F",X"1F",X"00",
		X"01",X"01",X"01",X"00",X"08",X"08",X"FF",X"00",X"05",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"08",X"08",X"FF",X"00",X"30",X"00",X"00",X"00",X"7F",X"00",X"00",X"00",X"30",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"7F",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"40",X"00",X"00",X"04",X"3F",X"00",X"00",X"1F",X"40",X"00",X"00",X"04",X"FF",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"80",X"02",X"00",X"00",X"03",
		X"3F",X"00",X"00",X"3F",X"02",X"00",X"00",X"03",X"FF",X"00",X"00",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"80",X"40",X"00",X"00",X"00",X"7F",X"00",X"00",X"00",
		X"40",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"00",X"00",X"00",X"F8",X"2C",X"F8",X"20",X"F8",X"74",X"F8",X"5C",X"F8",X"80",X"F8",X"2C",
		X"F8",X"2C",X"F8",X"44",X"F8",X"50",X"F8",X"5C",X"F8",X"CC",X"F8",X"68",X"F8",X"38",X"F8",X"44",
		X"F8",X"C0",X"F8",X"8C",X"F8",X"98",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F9",X"A8",X"F8",X"01",X"F9",X"EA",X"F8",X"01");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
