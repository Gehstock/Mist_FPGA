library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity prom_ic40 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of prom_ic40 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"24",X"18",X"7E",X"18",X"24",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"24",X"42",X"42",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"3E",X"00",X"00",X"00",X"3E",X"00",X"00",X"00",X"00",X"00",X"F0",
		X"00",X"00",X"00",X"7C",X"00",X"00",X"00",X"00",X"00",X"7C",X"00",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"00",X"00",X"00",X"F0",X"00",X"00",
		X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"00",
		X"00",X"F0",X"00",X"00",X"00",X"00",X"7C",X"00",X"00",X"00",X"00",X"00",X"7C",X"00",X"00",X"00",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"3E",X"00",X"00",X"00",X"3E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"00",X"00",X"00",X"00",X"FC",X"00",X"FC",X"00",X"00",X"00",X"00",X"C0",X"00",X"DC",
		X"C0",X"00",X"00",X"00",X"FC",X"00",X"00",X"00",X"FC",X"00",X"00",X"00",X"C0",X"00",X"DC",X"00",
		X"00",X"00",X"FC",X"00",X"00",X"00",X"00",X"00",X"FC",X"00",X"00",X"C0",X"00",X"DC",X"00",X"C0",
		X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"00",X"C0",X"00",X"DC",X"00",X"C0",X"00",
		X"00",X"C0",X"00",X"DC",X"00",X"C0",X"00",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",
		X"C0",X"00",X"DC",X"00",X"C0",X"00",X"00",X"FC",X"00",X"00",X"00",X"00",X"00",X"FC",X"00",X"00",
		X"00",X"DC",X"00",X"C0",X"00",X"00",X"00",X"FC",X"00",X"00",X"00",X"FC",X"00",X"00",X"00",X"C0",
		X"DC",X"00",X"C0",X"00",X"00",X"00",X"00",X"FC",X"00",X"FC",X"00",X"00",X"00",X"00",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"00",X"00",X"00",
		X"00",X"00",X"00",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"00",X"00",X"00",X"00",X"0F",X"0F",X"00",X"00",
		X"00",X"00",X"0F",X"0F",X"00",X"00",X"00",X"00",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",
		X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7E",X"CC",X"01",X"00",X"01",X"CC",X"7E",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",
		X"01",X"00",X"01",X"1C",X"0E",X"FF",X"3E",X"00",X"00",X"00",X"00",X"00",X"3E",X"FF",X"0E",X"1C",
		X"01",X"1C",X"0E",X"07",X"0F",X"3E",X"FC",X"00",X"FC",X"3E",X"0F",X"07",X"0E",X"1C",X"01",X"00",
		X"0E",X"FF",X"3E",X"00",X"00",X"00",X"00",X"00",X"3E",X"FF",X"0E",X"1C",X"01",X"00",X"01",X"1C",
		X"FF",X"1C",X"01",X"00",X"01",X"1C",X"FF",X"00",X"AA",X"82",X"C6",X"C6",X"C6",X"82",X"82",X"82",
		X"FF",X"38",X"80",X"00",X"80",X"38",X"FF",X"00",X"82",X"82",X"82",X"C6",X"C6",X"C6",X"82",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0C",X"00",X"00",X"00",X"0C",X"00",X"00",X"1E",X"0C",X"01",X"00",X"01",X"00",X"1E",X"00",
		X"01",X"06",X"0C",X"18",X"10",X"20",X"00",X"00",X"00",X"00",X"04",X"08",X"1A",X"33",X"60",X"80",
		X"60",X"30",X"18",X"08",X"04",X"00",X"00",X"00",X"00",X"20",X"10",X"58",X"CC",X"06",X"01",X"00",
		X"80",X"01",X"06",X"CC",X"58",X"10",X"20",X"00",X"00",X"00",X"00",X"04",X"08",X"18",X"30",X"60",
		X"60",X"33",X"1A",X"08",X"04",X"00",X"00",X"00",X"00",X"20",X"10",X"18",X"0C",X"06",X"01",X"00",
		X"03",X"03",X"03",X"06",X"0E",X"1C",X"F8",X"E0",X"E0",X"F8",X"1C",X"0E",X"06",X"03",X"03",X"03",
		X"C6",X"82",X"82",X"82",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"AA",X"82",X"C6",X"C6",
		X"C0",X"C0",X"C0",X"60",X"70",X"38",X"1F",X"07",X"07",X"1F",X"38",X"70",X"60",X"C0",X"C0",X"C0",
		X"00",X"00",X"00",X"00",X"0A",X"11",X"11",X"0E",X"00",X"00",X"00",X"80",X"3C",X"80",X"00",X"00",
		X"F0",X"F8",X"3C",X"0C",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"00",X"C0",
		X"90",X"00",X"20",X"70",X"70",X"38",X"18",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",
		X"18",X"1C",X"0C",X"0C",X"1C",X"18",X"10",X"00",X"00",X"00",X"00",X"00",X"88",X"E4",X"C0",X"08",
		X"40",X"20",X"08",X"30",X"60",X"C0",X"80",X"00",X"80",X"40",X"60",X"30",X"18",X"04",X"00",X"00",
		X"00",X"00",X"08",X"30",X"60",X"C0",X"80",X"00",X"80",X"40",X"60",X"30",X"18",X"04",X"10",X"20",
		X"F0",X"C0",X"10",X"00",X"10",X"C0",X"F0",X"00",X"F0",X"80",X"02",X"07",X"02",X"80",X"F0",X"00",
		X"C6",X"C6",X"82",X"AA",X"00",X"00",X"00",X"00",X"10",X"38",X"10",X"00",X"82",X"82",X"82",X"C6",
		X"00",X"C0",X"C0",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"C0",X"E0",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"38",X"1C",X"1C",X"0E",X"0E",X"04",X"00",
		X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"1C",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"0F",X"1C",X"00",
		X"02",X"04",X"0C",X"18",X"30",X"40",X"00",X"00",X"04",X"08",X"20",X"18",X"0C",X"06",X"02",X"01",
		X"02",X"04",X"0C",X"18",X"30",X"40",X"10",X"09",X"00",X"00",X"20",X"18",X"0C",X"06",X"02",X"01",
		X"0F",X"01",X"40",X"E0",X"40",X"01",X"0F",X"00",X"0F",X"03",X"08",X"00",X"08",X"03",X"0F",X"00",
		X"7A",X"F9",X"D0",X"83",X"87",X"03",X"03",X"1E",X"1E",X"07",X"03",X"87",X"83",X"D0",X"F9",X"7A",
		X"02",X"00",X"01",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"01",X"00",X"02",X"00",
		X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",
		X"28",X"70",X"60",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"20",X"10",X"00",X"00",
		X"04",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"E0",X"70",X"08",
		X"08",X"70",X"E0",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"04",
		X"04",X"00",X"10",X"20",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"60",X"70",X"28",
		X"C0",X"00",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0C",X"3C",X"F8",X"F0",
		X"38",X"70",X"70",X"20",X"00",X"10",X"20",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"18",X"18",
		X"08",X"C0",X"E4",X"88",X"00",X"00",X"00",X"00",X"00",X"10",X"18",X"18",X"0C",X"0C",X"1C",X"18",
		X"20",X"0E",X"1C",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"1C",X"0E",X"20",X"00",
		X"20",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"07",X"0E",X"10",
		X"14",X"0E",X"06",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"04",X"08",X"00",X"00",
		X"20",X"00",X"08",X"04",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"06",X"0E",X"14",
		X"10",X"0E",X"07",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"20",
		X"00",X"04",X"0E",X"0E",X"1C",X"1C",X"38",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"00",X"03",X"07",X"1F",X"7C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"1C",X"0F",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"08",X"1C",X"08",X"00",X"00",X"00",
		X"00",X"10",X"78",X"62",X"46",X"0E",X"1C",X"00",X"00",X"04",X"10",X"80",X"00",X"08",X"02",X"00",
		X"03",X"03",X"06",X"0E",X"3C",X"FC",X"F8",X"E0",X"00",X"08",X"00",X"01",X"00",X"01",X"01",X"01",
		X"01",X"01",X"01",X"00",X"01",X"00",X"08",X"00",X"E0",X"F8",X"FC",X"3C",X"0E",X"06",X"03",X"03",
		X"0C",X"80",X"40",X"20",X"10",X"08",X"00",X"42",X"C4",X"80",X"E0",X"FA",X"C0",X"80",X"60",X"10",
		X"00",X"08",X"10",X"22",X"C0",X"80",X"88",X"20",X"00",X"00",X"00",X"0C",X"0C",X"00",X"00",X"00",
		X"E0",X"E0",X"C0",X"80",X"C3",X"E0",X"E0",X"C0",X"00",X"0C",X"00",X"00",X"00",X"80",X"80",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"C0",X"60",X"70",X"3C",X"3F",X"1F",X"07",X"00",X"10",X"00",X"80",X"00",X"80",X"80",X"80",
		X"80",X"80",X"80",X"00",X"80",X"00",X"10",X"00",X"07",X"1F",X"3F",X"3C",X"70",X"60",X"C0",X"C0",
		X"1B",X"19",X"20",X"24",X"00",X"42",X"10",X"00",X"1F",X"1F",X"3F",X"FF",X"3F",X"3F",X"5F",X"0E",
		X"00",X"00",X"24",X"80",X"44",X"45",X"2B",X"2F",X"03",X"00",X"00",X"20",X"00",X"00",X"08",X"00",
		X"3F",X"3F",X"1F",X"1F",X"1F",X"3F",X"3F",X"03",X"00",X"40",X"04",X"00",X"00",X"19",X"1F",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"60",X"78",X"3C",X"1E",X"0E",X"06",X"00",X"00",X"38",X"38",X"38",X"18",X"18",X"38",X"38",
		X"00",X"00",X"07",X"7F",X"FE",X"E0",X"00",X"00",X"03",X"07",X"77",X"DD",X"FF",X"F6",X"3C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"70",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"0C",X"0C",X"0C",X"1C",X"18",X"18",X"38",X"30",
		X"30",X"38",X"18",X"18",X"1C",X"0C",X"0C",X"0C",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"70",
		X"0C",X"1C",X"38",X"70",X"E0",X"C0",X"00",X"00",X"03",X"03",X"03",X"03",X"07",X"06",X"06",X"0E",
		X"0E",X"06",X"06",X"07",X"03",X"03",X"03",X"03",X"00",X"00",X"C0",X"E0",X"70",X"38",X"1C",X"0C",
		X"0E",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"30",X"30",X"30",X"38",X"18",X"18",X"1C",X"0C",
		X"0C",X"1C",X"18",X"18",X"38",X"30",X"30",X"30",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"0E",
		X"30",X"38",X"1C",X"0E",X"07",X"03",X"00",X"00",X"C0",X"C0",X"C0",X"C0",X"E0",X"60",X"60",X"70",
		X"70",X"60",X"60",X"E0",X"C0",X"C0",X"C0",X"C0",X"00",X"00",X"03",X"07",X"0E",X"1C",X"38",X"30",
		X"00",X"00",X"03",X"1F",X"FE",X"F0",X"00",X"00",X"00",X"00",X"C0",X"F8",X"7F",X"0F",X"00",X"00",
		X"00",X"00",X"0F",X"7F",X"F8",X"C0",X"00",X"00",X"00",X"00",X"F0",X"FE",X"1F",X"03",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"0F",X"FF",X"F8",X"00",X"00",X"00",X"00",X"80",X"F0",X"7F",X"1F",
		X"1F",X"FF",X"F0",X"80",X"00",X"00",X"00",X"00",X"F8",X"FF",X"0F",X"01",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
