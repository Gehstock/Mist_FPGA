library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity MOONCR_ROM_PGM_0 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of MOONCR_ROM_PGM_0 is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"AF",X"32",X"01",X"70",X"C3",X"AD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F5",X"3A",X"00",X"78",X"AF",X"32",X"01",X"70",X"F1",X"C3",
		X"DE",X"00",X"3A",X"00",X"78",X"3E",X"01",X"32",X"04",X"70",X"AF",X"32",X"01",X"70",X"21",X"FF",
		X"00",X"22",X"00",X"40",X"31",X"00",X"44",X"CD",X"2B",X"01",X"AF",X"32",X"04",X"40",X"CD",X"CF",
		X"00",X"C3",X"29",X"02",X"AF",X"32",X"01",X"70",X"AF",X"32",X"04",X"40",X"21",X"1D",X"40",X"3E",
		X"04",X"36",X"00",X"23",X"3D",X"C2",X"A1",X"00",X"36",X"20",X"C3",X"29",X"02",X"21",X"00",X"40",
		X"11",X"00",X"04",X"36",X"00",X"23",X"1B",X"7A",X"B3",X"C2",X"B3",X"00",X"31",X"00",X"44",X"3E",
		X"0E",X"CD",X"92",X"08",X"3E",X"02",X"CD",X"32",X"09",X"CD",X"38",X"2F",X"C3",X"72",X"00",X"21",
		X"1D",X"40",X"3E",X"04",X"36",X"20",X"23",X"3D",X"C2",X"D4",X"00",X"36",X"40",X"C9",X"F5",X"C5",
		X"D5",X"E5",X"DD",X"E5",X"FD",X"E5",X"CD",X"32",X"01",X"3A",X"00",X"78",X"31",X"00",X"44",X"3A",
		X"3A",X"40",X"FE",X"04",X"C2",X"FA",X"00",X"32",X"32",X"40",X"00",X"21",X"05",X"40",X"34",X"7E",
		X"B7",X"C2",X"06",X"01",X"23",X"34",X"CD",X"9F",X"03",X"3A",X"05",X"40",X"E6",X"03",X"C2",X"14",
		X"01",X"CD",X"7A",X"04",X"CD",X"4D",X"01",X"CD",X"D6",X"01",X"3A",X"33",X"40",X"E6",X"01",X"C2",
		X"8A",X"00",X"CD",X"F2",X"01",X"CD",X"F2",X"01",X"C3",X"29",X"02",X"21",X"8B",X"03",X"22",X"02",
		X"40",X"C9",X"32",X"07",X"40",X"2A",X"00",X"40",X"7D",X"FE",X"FF",X"C8",X"11",X"09",X"40",X"29",
		X"19",X"EB",X"21",X"00",X"00",X"39",X"23",X"23",X"EB",X"73",X"23",X"72",X"C9",X"3A",X"00",X"60",
		X"E6",X"01",X"C2",X"C0",X"01",X"3A",X"00",X"60",X"E6",X"02",X"C2",X"40",X"03",X"3A",X"31",X"40",
		X"B7",X"C8",X"CD",X"30",X"03",X"B7",X"CA",X"8D",X"01",X"3A",X"32",X"40",X"FE",X"50",X"D2",X"7A",
		X"01",X"47",X"3A",X"3A",X"40",X"80",X"27",X"32",X"32",X"40",X"AF",X"32",X"31",X"40",X"CD",X"61",
		X"0E",X"3A",X"35",X"40",X"B7",X"C0",X"AF",X"32",X"04",X"40",X"C3",X"72",X"00",X"3A",X"39",X"40",
		X"3C",X"32",X"39",X"40",X"47",X"AF",X"32",X"31",X"40",X"3A",X"38",X"40",X"B8",X"C0",X"3E",X"00",
		X"32",X"39",X"40",X"3A",X"32",X"40",X"FE",X"50",X"D2",X"B1",X"01",X"C6",X"01",X"27",X"32",X"32",
		X"40",X"CD",X"61",X"0E",X"3A",X"35",X"40",X"B7",X"C0",X"AF",X"32",X"04",X"40",X"C3",X"72",X"00",
		X"3E",X"00",X"32",X"37",X"40",X"3C",X"32",X"31",X"40",X"32",X"03",X"60",X"C9",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"0A",X"21",X"27",X"40",X"11",X"1D",X"40",X"AF",X"BE",
		X"CA",X"E7",X"01",X"35",X"C2",X"EB",X"01",X"1A",X"E6",X"EF",X"12",X"23",X"13",X"05",X"C2",X"DE",
		X"01",X"C9",X"21",X"1D",X"40",X"3A",X"05",X"40",X"E6",X"00",X"C2",X"01",X"02",X"7E",X"F6",X"40",
		X"77",X"23",X"3A",X"05",X"40",X"E6",X"00",X"C2",X"0E",X"02",X"7E",X"F6",X"40",X"77",X"23",X"3A",
		X"05",X"40",X"E6",X"00",X"C2",X"1B",X"02",X"7E",X"F6",X"40",X"77",X"23",X"3A",X"05",X"40",X"E6",
		X"01",X"C2",X"28",X"02",X"7E",X"F6",X"40",X"77",X"C9",X"3A",X"00",X"78",X"3A",X"04",X"40",X"B7",
		X"C2",X"6C",X"02",X"3E",X"FF",X"32",X"00",X"40",X"00",X"AF",X"32",X"01",X"70",X"3E",X"01",X"32",
		X"01",X"70",X"00",X"01",X"00",X"0F",X"21",X"1D",X"40",X"7E",X"E6",X"30",X"C2",X"55",X"02",X"7E",
		X"E6",X"C0",X"C2",X"5E",X"02",X"23",X"0C",X"05",X"C2",X"49",X"02",X"C3",X"38",X"02",X"AF",X"32",
		X"01",X"70",X"79",X"32",X"00",X"40",X"7E",X"E6",X"80",X"CA",X"8C",X"02",X"2A",X"00",X"40",X"11",
		X"09",X"40",X"29",X"19",X"5E",X"23",X"56",X"EB",X"F9",X"FD",X"E1",X"DD",X"E1",X"E1",X"D1",X"C1",
		X"AF",X"32",X"01",X"70",X"3E",X"01",X"32",X"01",X"70",X"F1",X"ED",X"45",X"36",X"80",X"2A",X"00",
		X"40",X"11",X"95",X"03",X"29",X"19",X"5E",X"23",X"56",X"EB",X"F9",X"2A",X"00",X"40",X"EB",X"2A",
		X"02",X"40",X"19",X"19",X"5E",X"23",X"56",X"EB",X"AF",X"32",X"01",X"70",X"3E",X"01",X"32",X"01",
		X"70",X"E9",X"F5",X"AF",X"32",X"01",X"70",X"F1",X"F5",X"C5",X"D5",X"E5",X"DD",X"E5",X"FD",X"E5",
		X"F5",X"3A",X"04",X"40",X"B7",X"C3",X"E8",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AF",X"32",X"01",X"70",X"3E",X"01",X"32",X"01",
		X"70",X"F1",X"D6",X"01",X"DA",X"07",X"03",X"F5",X"21",X"00",X"01",X"E5",X"E1",X"2B",X"7C",X"B5",
		X"C2",X"FB",X"02",X"F1",X"C3",X"F2",X"02",X"FD",X"E1",X"DD",X"E1",X"E1",X"D1",X"C1",X"F1",X"C9",
		X"AF",X"32",X"01",X"70",X"2A",X"00",X"40",X"11",X"1D",X"40",X"19",X"7E",X"E6",X"7F",X"77",X"C3",
		X"29",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AF",X"32",X"03",X"60",X"32",X"04",X"68",X"3A",X"37",X"40",X"C9",X"00",X"00",X"00",X"00",X"00",
		X"3E",X"01",X"32",X"37",X"40",X"32",X"31",X"40",X"32",X"04",X"68",X"C9",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"00",X"10",X"00",
		X"30",X"00",X"20",X"7C",X"0A",X"E0",X"43",X"A8",X"43",X"70",X"43",X"38",X"43",X"E0",X"43",X"00",
		X"2A",X"EF",X"40",X"7E",X"E6",X"F8",X"FE",X"F8",X"C2",X"39",X"04",X"7E",X"FE",X"FF",X"CA",X"39",
		X"04",X"FE",X"F8",X"C2",X"CA",X"03",X"23",X"7E",X"32",X"06",X"68",X"0F",X"32",X"07",X"68",X"0F",
		X"32",X"FA",X"40",X"23",X"22",X"EF",X"40",X"C3",X"79",X"04",X"FE",X"FA",X"C2",X"DB",X"03",X"23",
		X"7E",X"32",X"F3",X"40",X"23",X"22",X"F5",X"40",X"C3",X"F8",X"03",X"FE",X"FB",X"C2",X"03",X"04",
		X"3A",X"F3",X"40",X"FE",X"00",X"CA",X"F8",X"03",X"2A",X"F5",X"40",X"22",X"EF",X"40",X"3A",X"F3",
		X"40",X"3D",X"32",X"F3",X"40",X"C3",X"79",X"04",X"2A",X"EF",X"40",X"23",X"23",X"22",X"EF",X"40",
		X"C3",X"79",X"04",X"FE",X"FC",X"C2",X"14",X"04",X"23",X"7E",X"32",X"F4",X"40",X"23",X"22",X"F7",
		X"40",X"C3",X"F8",X"03",X"FE",X"FD",X"C2",X"31",X"04",X"3A",X"F4",X"40",X"FE",X"00",X"CA",X"F8",
		X"03",X"2A",X"F7",X"40",X"22",X"EF",X"40",X"3A",X"F4",X"40",X"3D",X"32",X"F4",X"40",X"C3",X"79",
		X"04",X"FE",X"FE",X"C2",X"F8",X"03",X"C3",X"79",X"04",X"7E",X"32",X"00",X"78",X"3A",X"F9",X"40",
		X"47",X"3A",X"F1",X"40",X"3C",X"32",X"F1",X"40",X"B8",X"DA",X"79",X"04",X"AF",X"32",X"F1",X"40",
		X"3A",X"FA",X"40",X"E6",X"01",X"C2",X"62",X"04",X"2A",X"EF",X"40",X"23",X"22",X"EF",X"40",X"C3",
		X"79",X"04",X"3A",X"F2",X"40",X"3C",X"32",X"F2",X"40",X"23",X"46",X"3A",X"F2",X"40",X"B8",X"DA",
		X"79",X"04",X"AF",X"32",X"F2",X"40",X"C3",X"F8",X"03",X"C9",X"00",X"2A",X"FB",X"40",X"7E",X"E6",
		X"F0",X"FE",X"F0",X"C2",X"11",X"05",X"7E",X"FE",X"FA",X"C2",X"99",X"04",X"23",X"7E",X"32",X"FE",
		X"40",X"23",X"22",X"00",X"41",X"22",X"FB",X"40",X"C9",X"FE",X"FB",X"C2",X"B4",X"04",X"3A",X"FE",
		X"40",X"FE",X"00",X"CA",X"E7",X"04",X"2A",X"00",X"41",X"22",X"FB",X"40",X"3A",X"FE",X"40",X"3D",
		X"32",X"FE",X"40",X"C9",X"FE",X"FC",X"C2",X"C6",X"04",X"23",X"7E",X"32",X"FF",X"40",X"23",X"22",
		X"00",X"41",X"22",X"FB",X"40",X"C9",X"FE",X"FD",X"C2",X"E1",X"04",X"3A",X"FF",X"40",X"FE",X"00",
		X"CA",X"E7",X"04",X"2A",X"02",X"41",X"22",X"FB",X"40",X"3A",X"FF",X"40",X"3D",X"32",X"FF",X"40",
		X"C9",X"FE",X"FE",X"C2",X"E7",X"04",X"C9",X"2A",X"FB",X"40",X"23",X"22",X"FB",X"40",X"C9",X"2A",
		X"FB",X"40",X"7E",X"32",X"04",X"60",X"0F",X"32",X"05",X"60",X"0F",X"32",X"06",X"60",X"0F",X"32",
		X"07",X"60",X"0F",X"32",X"00",X"68",X"0F",X"32",X"01",X"68",X"0F",X"32",X"02",X"68",X"C3",X"2C",
		X"05",X"7E",X"E6",X"90",X"FE",X"80",X"C2",X"20",X"05",X"7E",X"32",X"05",X"68",X"C3",X"2C",X"05",
		X"7E",X"E6",X"90",X"FE",X"90",X"C2",X"EF",X"04",X"7E",X"32",X"03",X"68",X"3A",X"04",X"41",X"47",
		X"3A",X"FD",X"40",X"3C",X"32",X"FD",X"40",X"B8",X"D8",X"AF",X"32",X"FD",X"40",X"C3",X"E7",X"04",
		X"F8",X"02",X"FA",X"02",X"1F",X"3F",X"5F",X"3F",X"5F",X"3F",X"5F",X"3F",X"7F",X"E0",X"F0",X"F7",
		X"F7",X"7C",X"BC",X"DC",X"EC",X"F4",X"F7",X"F0",X"E0",X"C0",X"80",X"00",X"00",X"3F",X"5F",X"3F",
		X"5F",X"3F",X"5F",X"3F",X"7F",X"E0",X"F0",X"F7",X"F7",X"7C",X"BC",X"DC",X"EC",X"F4",X"F7",X"F0",
		X"E0",X"C0",X"80",X"00",X"55",X"AA",X"A8",X"A0",X"80",X"00",X"FB",X"00",X"FF",X"FE",X"F8",X"02",
		X"00",X"00",X"01",X"00",X"03",X"00",X"06",X"00",X"0A",X"00",X"0F",X"00",X"15",X"00",X"1C",X"00",
		X"24",X"00",X"2D",X"00",X"37",X"00",X"42",X"00",X"FA",X"02",X"F8",X"01",X"D5",X"D3",X"CD",X"C7",
		X"F8",X"02",X"FC",X"02",X"D5",X"D3",X"CD",X"C7",X"FD",X"00",X"FF",X"FF",X"FF",X"FF",X"FB",X"00",
		X"FF",X"FE",X"F8",X"01",X"FA",X"02",X"D1",X"C9",X"C3",X"B8",X"AF",X"A0",X"94",X"87",X"6F",X"5E",
		X"3F",X"28",X"0D",X"FA",X"05",X"3F",X"0D",X"5E",X"28",X"6F",X"3F",X"87",X"5E",X"3F",X"6F",X"A0",
		X"87",X"AF",X"94",X"B8",X"A0",X"C3",X"AF",X"C9",X"B8",X"D1",X"C3",X"FB",X"00",X"FF",X"FE",X"F8",
		X"02",X"B8",X"B0",X"A8",X"A0",X"98",X"90",X"88",X"80",X"70",X"60",X"50",X"40",X"3C",X"34",X"2C",
		X"24",X"1B",X"17",X"13",X"0F",X"0B",X"07",X"03",X"13",X"FA",X"03",X"1F",X"23",X"27",X"2B",X"2F",
		X"33",X"37",X"3B",X"3B",X"37",X"33",X"2F",X"2B",X"27",X"23",X"1F",X"FB",X"00",X"FF",X"FE",X"F8",
		X"01",X"80",X"81",X"82",X"83",X"84",X"85",X"86",X"87",X"86",X"85",X"84",X"85",X"86",X"87",X"88",
		X"89",X"8A",X"8B",X"8C",X"8D",X"8E",X"8F",X"8E",X"8D",X"8C",X"8D",X"8E",X"8F",X"90",X"91",X"92",
		X"93",X"FA",X"05",X"A0",X"B0",X"C0",X"D0",X"E0",X"C0",X"80",X"7E",X"7C",X"78",X"70",X"68",X"60",
		X"58",X"50",X"48",X"40",X"18",X"10",X"08",X"FB",X"00",X"FF",X"FE",X"F8",X"0B",X"0D",X"D0",X"28",
		X"CA",X"3F",X"C4",X"5E",X"B8",X"6F",X"AF",X"87",X"A0",X"94",X"94",X"87",X"A0",X"6F",X"AF",X"5E",
		X"B8",X"3F",X"C4",X"28",X"CA",X"0D",X"D0",X"D0",X"D0",X"CA",X"28",X"C4",X"3F",X"B8",X"5E",X"AF",
		X"6E",X"A0",X"87",X"94",X"94",X"6B",X"FF",X"F8",X"00",X"FE",X"F8",X"0B",X"80",X"9A",X"AA",X"9A",
		X"80",X"9A",X"AA",X"9A",X"A5",X"8E",X"A5",X"8E",X"A5",X"8E",X"A5",X"8E",X"FF",X"F8",X"00",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"0B",X"13",X"65",X"63",X"51",X"91",X"C3",X"AA",X"A9",X"A5",X"BB",X"D5",X"6A",X"40",X"D5",
		X"80",X"C9",X"12",X"D3",X"D9",X"C9",X"33",X"12",X"C0",X"00",X"FF",X"F8",X"00",X"FE",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"09",X"B8",X"AF",X"A0",X"94",X"AF",X"A0",X"94",X"87",
		X"A0",X"94",X"87",X"6F",X"94",X"87",X"6F",X"5E",X"87",X"6F",X"54",X"3F",X"6F",X"5E",X"3F",X"28",
		X"5E",X"3F",X"28",X"0D",X"FF",X"F8",X"00",X"FE",X"F8",X"0B",X"E0",X"C0",X"80",X"BF",X"9F",X"8F",
		X"87",X"83",X"7B",X"3B",X"1B",X"0B",X"03",X"01",X"00",X"00",X"FF",X"F8",X"00",X"FE",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"07",
		X"FA",X"01",X"00",X"00",X"28",X"00",X"54",X"00",X"FF",X"02",X"54",X"01",X"80",X"10",X"94",X"01",
		X"80",X"02",X"94",X"01",X"AA",X"10",X"FF",X"04",X"FB",X"00",X"F8",X"0F",X"C0",X"00",X"FF",X"06",
		X"C0",X"00",X"FF",X"05",X"C0",X"00",X"FF",X"04",X"C0",X"00",X"FF",X"03",X"C0",X"00",X"FF",X"02",
		X"C0",X"00",X"FF",X"01",X"C0",X"00",X"FF",X"01",X"F8",X"07",X"F8",X"01",X"FA",X"07",X"C0",X"FF",
		X"C0",X"FF",X"E0",X"DF",X"DE",X"DD",X"DC",X"DB",X"DA",X"DC",X"DA",X"DB",X"DC",X"DD",X"DE",X"DF",
		X"E0",X"E1",X"E2",X"E3",X"E4",X"E5",X"E6",X"E7",X"E8",X"E9",X"FB",X"00",X"FF",X"FE",X"F8",X"03",
		X"54",X"67",X"77",X"C7",X"D7",X"E7",X"F7",X"FF",X"F8",X"07",X"FF",X"10",X"54",X"04",X"FF",X"04",
		X"54",X"04",X"77",X"04",X"8E",X"04",X"77",X"04",X"8E",X"04",X"77",X"04",X"67",X"04",X"FF",X"04",
		X"67",X"04",X"80",X"04",X"9A",X"0C",X"A5",X"04",X"8E",X"04",X"77",X"04",X"A5",X"04",X"8E",X"04",
		X"77",X"04",X"A5",X"04",X"8E",X"04",X"AA",X"04",X"FF",X"04",X"A5",X"04",X"AA",X"10",X"FF",X"00",
		X"FE",X"00",X"F8",X"03",X"C7",X"FF",X"D5",X"C7",X"BC",X"FF",X"C7",X"BC",X"AA",X"FF",X"BC",X"AA",
		X"8E",X"8E",X"FF",X"FF",X"8E",X"87",X"8E",X"94",X"9A",X"94",X"9A",X"A5",X"AA",X"AA",X"FF",X"FF",
		X"8E",X"FF",X"8E",X"F8",X"07",X"94",X"03",X"8E",X"05",X"FF",X"02",X"A5",X"00",X"FF",X"03",X"AA",
		X"00",X"FF",X"00",X"FE",X"00",X"F8",X"03",X"FC",X"01",X"1B",X"34",X"44",X"FA",X"07",X"54",X"FB",
		X"00",X"FF",X"54",X"FF",X"54",X"FF",X"54",X"FF",X"FA",X"07",X"54",X"FB",X"00",X"44",X"54",X"67",
		X"FA",X"07",X"77",X"FB",X"00",X"FF",X"77",X"FF",X"77",X"FF",X"77",X"FF",X"FA",X"07",X"77",X"FB",
		X"00",X"54",X"77",X"80",X"FA",X"07",X"8E",X"FB",X"00",X"FF",X"8E",X"FF",X"8E",X"FF",X"8E",X"FF",
		X"FA",X"07",X"8E",X"FB",X"00",X"77",X"8E",X"A5",X"FA",X"07",X"AB",X"FB",X"00",X"FF",X"AB",X"FF",
		X"AB",X"FF",X"AB",X"FF",X"FA",X"07",X"AB",X"FB",X"00",X"FD",X"00",X"FF",X"FE",X"F8",X"00",X"FF",
		X"FE",X"F8",X"17",X"FA",X"0E",X"AA",X"04",X"D5",X"01",X"FF",X"00",X"FB",X"00",X"F8",X"07",X"FE",
		X"00",X"30",X"31",X"32",X"33",X"34",X"35",X"36",X"37",X"38",X"39",X"3A",X"3B",X"3C",X"3D",X"3E",
		X"3F",X"00",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"81",X"80",X"FE",X"80",X"FA",X"08",X"91",X"FB",X"00",X"90",X"FE",X"80",X"90",
		X"00",X"FE",X"00",X"E5",X"D5",X"57",X"FE",X"0E",X"CA",X"C9",X"08",X"3A",X"35",X"40",X"B7",X"CA",
		X"EB",X"08",X"3A",X"FA",X"40",X"E6",X"04",X"C2",X"EB",X"08",X"7A",X"FE",X"10",X"CA",X"D1",X"08",
		X"FE",X"05",X"CA",X"D1",X"08",X"FE",X"06",X"CA",X"D1",X"08",X"FE",X"07",X"CA",X"D1",X"08",X"FE",
		X"08",X"CA",X"D1",X"08",X"FE",X"09",X"CA",X"D1",X"08",X"3A",X"FA",X"40",X"E6",X"02",X"C2",X"EB",
		X"08",X"21",X"EE",X"08",X"7A",X"07",X"07",X"E6",X"FC",X"5F",X"16",X"00",X"19",X"7E",X"32",X"F9",
		X"40",X"23",X"7E",X"32",X"EF",X"40",X"23",X"7E",X"32",X"F0",X"40",X"D1",X"E1",X"C9",X"02",X"40",
		X"05",X"00",X"01",X"7E",X"05",X"00",X"01",X"B2",X"05",X"00",X"01",X"DF",X"05",X"00",X"01",X"0F",
		X"06",X"00",X"01",X"4B",X"06",X"00",X"02",X"7A",X"06",X"00",X"02",X"A0",X"06",X"00",X"02",X"C6",
		X"06",X"00",X"02",X"E8",X"06",X"00",X"03",X"0E",X"07",X"00",X"02",X"6E",X"07",X"00",X"04",X"B2",
		X"07",X"00",X"01",X"E5",X"07",X"00",X"01",X"3D",X"08",X"00",X"03",X"2A",X"07",X"00",X"02",X"41",
		X"08",X"00",X"00",X"E5",X"D5",X"57",X"FE",X"02",X"CA",X"42",X"09",X"3A",X"35",X"40",X"B7",X"CA",
		X"62",X"09",X"00",X"21",X"65",X"09",X"7A",X"07",X"07",X"E6",X"FC",X"5F",X"16",X"00",X"19",X"7E",
		X"32",X"04",X"41",X"23",X"7E",X"32",X"FB",X"40",X"23",X"7E",X"32",X"FC",X"40",X"23",X"7E",X"32",
		X"FD",X"40",X"D1",X"E1",X"C9",X"01",X"83",X"08",X"00",X"01",X"86",X"08",X"00",X"01",X"8E",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"F5",X"C5",X"D5",X"E5",X"D5",X"DD",X"E1",X"DD",X"7E",X"01",X"87",X"06",X"00",X"4F",X"FD",
		X"21",X"00",X"58",X"FD",X"09",X"FD",X"36",X"00",X"00",X"DD",X"7E",X"00",X"FD",X"77",X"01",X"DD",
		X"46",X"02",X"3E",X"1B",X"90",X"B7",X"CA",X"B4",X"09",X"21",X"40",X"50",X"01",X"20",X"00",X"09",
		X"3D",X"C2",X"AF",X"09",X"DD",X"4E",X"01",X"06",X"00",X"09",X"01",X"E0",X"FF",X"DD",X"23",X"DD",
		X"23",X"DD",X"23",X"DD",X"7E",X"00",X"FE",X"FF",X"CA",X"D8",X"09",X"77",X"09",X"7C",X"FE",X"50",
		X"DA",X"D8",X"09",X"DD",X"23",X"C3",X"C3",X"09",X"E1",X"D1",X"C1",X"F1",X"C9",X"00",X"F5",X"C5",
		X"D5",X"E5",X"D5",X"DD",X"E1",X"DD",X"7E",X"01",X"87",X"06",X"00",X"4F",X"FD",X"21",X"00",X"58",
		X"FD",X"09",X"FD",X"36",X"00",X"00",X"DD",X"7E",X"00",X"FD",X"77",X"01",X"DD",X"46",X"02",X"3E",
		X"1B",X"90",X"B7",X"CA",X"13",X"0A",X"FD",X"21",X"40",X"50",X"01",X"20",X"00",X"FD",X"09",X"3D",
		X"C2",X"0D",X"0A",X"DD",X"4E",X"01",X"06",X"00",X"FD",X"09",X"01",X"E0",X"FF",X"DD",X"56",X"05",
		X"DD",X"66",X"04",X"DD",X"6E",X"03",X"CB",X"42",X"CA",X"35",X"0A",X"7E",X"E6",X"0F",X"FD",X"77",
		X"00",X"23",X"C3",X"3F",X"0A",X"7E",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"FD",X"77",X"00",X"FD",
		X"09",X"15",X"C2",X"26",X"0A",X"E1",X"D1",X"C1",X"F1",X"C9",X"00",X"21",X"00",X"50",X"01",X"00",
		X"04",X"36",X"24",X"23",X"0B",X"78",X"B1",X"C2",X"51",X"0A",X"00",X"21",X"40",X"58",X"01",X"40",
		X"00",X"36",X"00",X"23",X"0B",X"78",X"B1",X"C2",X"61",X"0A",X"C9",X"00",X"21",X"40",X"41",X"01",
		X"80",X"01",X"36",X"00",X"23",X"0B",X"78",X"B1",X"C2",X"72",X"0A",X"C9",X"00",X"3A",X"33",X"40",
		X"B7",X"C2",X"3D",X"0B",X"06",X"00",X"3A",X"32",X"40",X"B7",X"CA",X"8E",X"0A",X"04",X"78",X"32",
		X"35",X"40",X"CD",X"A2",X"0A",X"3E",X"01",X"32",X"34",X"40",X"3E",X"01",X"32",X"04",X"40",X"C3",
		X"94",X"00",X"00",X"3E",X"01",X"32",X"3F",X"40",X"CD",X"4A",X"0A",X"CD",X"FC",X"0C",X"CD",X"61",
		X"0E",X"3A",X"35",X"40",X"B7",X"C2",X"CF",X"0A",X"CD",X"A4",X"0D",X"CD",X"6F",X"2D",X"3E",X"FF",
		X"CD",X"B2",X"02",X"3E",X"FF",X"CD",X"B2",X"02",X"AF",X"32",X"3F",X"40",X"C3",X"21",X"0B",X"CD",
		X"6F",X"2D",X"3A",X"32",X"40",X"FE",X"01",X"C2",X"E0",X"0A",X"CD",X"9B",X"0E",X"C3",X"E3",X"0A",
		X"CD",X"D2",X"0E",X"00",X"3A",X"00",X"68",X"E6",X"02",X"FE",X"02",X"CA",X"FB",X"0A",X"3A",X"00",
		X"68",X"E6",X"01",X"FE",X"01",X"CA",X"14",X"0B",X"C3",X"D2",X"0A",X"3A",X"32",X"40",X"FE",X"02",
		X"DA",X"D2",X"0A",X"3E",X"01",X"32",X"3F",X"40",X"3A",X"32",X"40",X"C6",X"98",X"27",X"32",X"32",
		X"40",X"C3",X"21",X"0B",X"AF",X"32",X"3F",X"40",X"3A",X"32",X"40",X"C6",X"99",X"27",X"32",X"32",
		X"40",X"CD",X"61",X"0E",X"CD",X"6B",X"0A",X"CD",X"A1",X"0C",X"AF",X"CD",X"1E",X"0C",X"3E",X"01",
		X"CD",X"1E",X"0C",X"3A",X"BE",X"40",X"32",X"41",X"40",X"CD",X"FC",X"0C",X"C9",X"00",X"AF",X"32",
		X"33",X"40",X"CD",X"5A",X"0A",X"3A",X"97",X"40",X"3D",X"32",X"97",X"40",X"3A",X"40",X"40",X"CD",
		X"1E",X"0C",X"3A",X"97",X"40",X"B7",X"CA",X"A1",X"0B",X"3A",X"3F",X"40",X"B7",X"CA",X"90",X"0B",
		X"3A",X"41",X"40",X"B7",X"CA",X"90",X"0B",X"3A",X"40",X"40",X"3C",X"E6",X"01",X"32",X"40",X"40",
		X"3A",X"3C",X"40",X"B7",X"CA",X"90",X"0B",X"3A",X"40",X"40",X"B7",X"C2",X"89",X"0B",X"3E",X"01",
		X"32",X"06",X"70",X"32",X"07",X"70",X"C3",X"90",X"0B",X"AF",X"32",X"06",X"70",X"32",X"07",X"70",
		X"CD",X"6B",X"0A",X"3A",X"40",X"40",X"CD",X"56",X"0C",X"3E",X"01",X"32",X"04",X"40",X"C3",X"94",
		X"00",X"3A",X"35",X"40",X"B7",X"CA",X"72",X"00",X"CD",X"0C",X"0F",X"3A",X"9E",X"40",X"B7",X"C2",
		X"E8",X"0B",X"3A",X"9D",X"40",X"B7",X"CA",X"E8",X"0B",X"CD",X"A1",X"0C",X"3A",X"9B",X"40",X"C6",
		X"10",X"F6",X"01",X"E6",X"F1",X"32",X"9B",X"40",X"3C",X"32",X"9C",X"40",X"3E",X"01",X"32",X"9E",
		X"40",X"3A",X"40",X"40",X"CD",X"1E",X"0C",X"3A",X"3F",X"40",X"B7",X"CA",X"90",X"0B",X"3A",X"41",
		X"40",X"B7",X"C2",X"67",X"0B",X"C3",X"90",X"0B",X"AF",X"32",X"9D",X"40",X"CD",X"00",X"2A",X"3A",
		X"3F",X"40",X"B7",X"CA",X"FD",X"0B",X"3A",X"41",X"40",X"B7",X"C2",X"67",X"0B",X"CD",X"78",X"0F",
		X"AF",X"32",X"33",X"40",X"32",X"34",X"40",X"32",X"35",X"40",X"32",X"3F",X"40",X"32",X"40",X"40",
		X"3E",X"01",X"32",X"06",X"70",X"32",X"07",X"70",X"32",X"04",X"40",X"C3",X"72",X"00",X"00",X"B7",
		X"C2",X"2A",X"0C",X"FD",X"21",X"9F",X"40",X"C3",X"2E",X"0C",X"FD",X"21",X"BE",X"40",X"DD",X"21",
		X"97",X"40",X"01",X"01",X"00",X"11",X"01",X"00",X"26",X"08",X"CD",X"EC",X"0C",X"DD",X"21",X"40",
		X"41",X"01",X"01",X"00",X"26",X"0F",X"CD",X"EC",X"0C",X"DD",X"21",X"82",X"41",X"01",X"14",X"00",
		X"26",X"08",X"CD",X"EC",X"0C",X"C9",X"00",X"B7",X"C2",X"68",X"0C",X"3A",X"BE",X"40",X"32",X"41",
		X"40",X"DD",X"21",X"9F",X"40",X"C3",X"72",X"0C",X"3A",X"9F",X"40",X"32",X"41",X"40",X"DD",X"21",
		X"BE",X"40",X"FD",X"21",X"97",X"40",X"01",X"01",X"00",X"11",X"01",X"00",X"26",X"08",X"CD",X"EC",
		X"0C",X"FD",X"21",X"40",X"41",X"11",X"01",X"00",X"26",X"0F",X"CD",X"EC",X"0C",X"FD",X"21",X"82",
		X"41",X"11",X"14",X"00",X"26",X"08",X"CD",X"EC",X"0C",X"AF",X"32",X"26",X"42",X"32",X"27",X"42",
		X"C9",X"00",X"3E",X"03",X"32",X"97",X"40",X"3A",X"9D",X"40",X"B7",X"C2",X"C2",X"0C",X"AF",X"32",
		X"98",X"40",X"32",X"99",X"40",X"32",X"9A",X"40",X"3E",X"01",X"32",X"9B",X"40",X"3E",X"02",X"32",
		X"9C",X"40",X"AF",X"32",X"9D",X"40",X"32",X"9E",X"40",X"AF",X"32",X"26",X"42",X"32",X"27",X"42",
		X"3E",X"03",X"32",X"40",X"41",X"32",X"45",X"41",X"32",X"4A",X"41",X"3E",X"01",X"21",X"82",X"41",
		X"11",X"14",X"00",X"06",X"08",X"77",X"19",X"05",X"C2",X"E5",X"0C",X"C9",X"00",X"DD",X"7E",X"00",
		X"FD",X"77",X"00",X"DD",X"09",X"FD",X"19",X"25",X"C2",X"ED",X"0C",X"C9",X"00",X"11",X"5F",X"0D",
		X"CD",X"80",X"09",X"11",X"7E",X"0D",X"CD",X"DD",X"09",X"11",X"84",X"0D",X"CD",X"DD",X"09",X"11",
		X"8A",X"0D",X"CD",X"DD",X"09",X"21",X"54",X"40",X"06",X"0A",X"0E",X"00",X"7E",X"FE",X"24",X"C2",
		X"23",X"0D",X"0C",X"23",X"05",X"C2",X"1C",X"0D",X"79",X"0F",X"E6",X"0F",X"C6",X"09",X"4F",X"DD",
		X"21",X"51",X"40",X"DD",X"36",X"00",X"03",X"DD",X"36",X"01",X"02",X"DD",X"71",X"02",X"DD",X"36",
		X"0D",X"FF",X"11",X"51",X"40",X"CD",X"80",X"09",X"3A",X"3F",X"40",X"B7",X"C0",X"3A",X"35",X"40",
		X"B7",X"C8",X"11",X"90",X"0D",X"CD",X"80",X"09",X"11",X"9A",X"0D",X"CD",X"80",X"09",X"C9",X"04",
		X"00",X"00",X"24",X"01",X"29",X"1C",X"1D",X"24",X"24",X"24",X"24",X"24",X"11",X"12",X"2B",X"1C",
		X"0C",X"18",X"1B",X"0E",X"24",X"24",X"24",X"24",X"24",X"02",X"29",X"17",X"0D",X"FF",X"07",X"01",
		X"00",X"A0",X"40",X"06",X"07",X"01",X"0B",X"42",X"40",X"06",X"07",X"01",X"16",X"BF",X"40",X"06",
		X"04",X"00",X"16",X"24",X"24",X"24",X"24",X"24",X"24",X"FF",X"07",X"01",X"16",X"24",X"24",X"24",
		X"24",X"24",X"24",X"FF",X"00",X"3E",X"01",X"32",X"04",X"40",X"3E",X"40",X"CD",X"B2",X"02",X"11",
		X"F2",X"0D",X"CD",X"48",X"2A",X"3E",X"40",X"CD",X"B2",X"02",X"11",X"0B",X"0E",X"CD",X"48",X"2A",
		X"3E",X"40",X"CD",X"B2",X"02",X"11",X"1A",X"0E",X"CD",X"48",X"2A",X"3E",X"40",X"CD",X"B2",X"02",
		X"11",X"2B",X"0E",X"CD",X"80",X"09",X"3E",X"40",X"CD",X"B2",X"02",X"11",X"40",X"0E",X"CD",X"80",
		X"09",X"3E",X"80",X"CD",X"B2",X"02",X"11",X"55",X"0E",X"CD",X"80",X"09",X"3E",X"FF",X"CD",X"B2",
		X"02",X"C9",X"03",X"06",X"05",X"1D",X"1B",X"12",X"19",X"24",X"1D",X"18",X"24",X"1D",X"11",X"0E",
		X"24",X"1C",X"19",X"0A",X"0C",X"0E",X"24",X"20",X"0A",X"1B",X"FF",X"02",X"09",X"09",X"16",X"18",
		X"18",X"17",X"24",X"0C",X"1B",X"0E",X"1C",X"1D",X"0A",X"FF",X"0E",X"0E",X"09",X"1D",X"1B",X"22",
		X"24",X"12",X"1D",X"24",X"17",X"18",X"20",X"24",X"28",X"28",X"FF",X"04",X"11",X"06",X"22",X"18",
		X"1E",X"24",X"0C",X"0A",X"17",X"24",X"10",X"0E",X"1D",X"24",X"0A",X"24",X"15",X"18",X"1D",X"FF",
		X"04",X"13",X"06",X"18",X"0F",X"24",X"0F",X"1E",X"17",X"24",X"0A",X"17",X"0D",X"24",X"1D",X"11",
		X"1B",X"12",X"15",X"15",X"FF",X"07",X"1B",X"0A",X"3E",X"3C",X"3A",X"38",X"36",X"34",X"32",X"30",
		X"FF",X"00",X"3A",X"3A",X"40",X"FE",X"04",X"CA",X"77",X"0E",X"11",X"8B",X"0E",X"CD",X"80",X"09",
		X"11",X"95",X"0E",X"CD",X"DD",X"09",X"C9",X"11",X"7E",X"0E",X"CD",X"80",X"09",X"C9",X"05",X"1F",
		X"00",X"0F",X"1B",X"0E",X"0E",X"24",X"19",X"15",X"0A",X"22",X"FF",X"05",X"1F",X"00",X"0C",X"1B",
		X"0E",X"0D",X"12",X"1D",X"FF",X"05",X"1F",X"07",X"32",X"40",X"02",X"00",X"11",X"AF",X"0E",X"CD",
		X"80",X"09",X"11",X"B7",X"0E",X"CD",X"80",X"09",X"11",X"CA",X"0E",X"CD",X"80",X"09",X"C9",X"04",
		X"10",X"0C",X"19",X"1E",X"1C",X"11",X"FF",X"04",X"12",X"07",X"01",X"24",X"19",X"15",X"0A",X"22",
		X"0E",X"1B",X"24",X"0B",X"1E",X"1D",X"1D",X"18",X"17",X"FF",X"04",X"14",X"0C",X"18",X"17",X"15",
		X"22",X"FF",X"00",X"11",X"E6",X"0E",X"CD",X"80",X"09",X"11",X"EE",X"0E",X"CD",X"80",X"09",X"11",
		X"02",X"0F",X"CD",X"80",X"09",X"C9",X"04",X"10",X"0C",X"19",X"1E",X"1C",X"11",X"FF",X"04",X"12",
		X"07",X"01",X"24",X"18",X"1B",X"24",X"02",X"24",X"19",X"15",X"0A",X"22",X"0E",X"1B",X"1C",X"24",
		X"24",X"FF",X"04",X"14",X"0B",X"0B",X"1E",X"1D",X"1D",X"18",X"17",X"FF",X"00",X"3A",X"9E",X"40",
		X"B7",X"C2",X"1B",X"0F",X"3A",X"9D",X"40",X"B7",X"C2",X"34",X"0F",X"3A",X"40",X"40",X"B7",X"C2",
		X"28",X"0F",X"11",X"40",X"0F",X"C3",X"2B",X"0F",X"11",X"51",X"0F",X"CD",X"80",X"09",X"3E",X"80",
		X"CD",X"B2",X"02",X"C9",X"11",X"62",X"0F",X"CD",X"80",X"09",X"3E",X"80",X"CD",X"B2",X"02",X"C9",
		X"00",X"0D",X"07",X"19",X"15",X"0A",X"22",X"0E",X"1B",X"24",X"01",X"24",X"18",X"1F",X"0E",X"1B",
		X"FF",X"00",X"0D",X"07",X"19",X"15",X"0A",X"22",X"0E",X"1B",X"24",X"02",X"24",X"18",X"1F",X"0E",
		X"1B",X"FF",X"00",X"0D",X"04",X"0E",X"17",X"13",X"18",X"22",X"24",X"0A",X"17",X"18",X"1D",X"11",
		X"0E",X"1B",X"24",X"10",X"0A",X"16",X"0E",X"FF",X"00",X"11",X"8E",X"0F",X"CD",X"80",X"09",X"3E",
		X"01",X"32",X"04",X"40",X"3E",X"80",X"CD",X"B2",X"02",X"AF",X"32",X"04",X"40",X"C9",X"00",X"11",
		X"09",X"10",X"0A",X"16",X"0E",X"24",X"18",X"1F",X"0E",X"1B",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"3A",X"3A",X"42",X"FE",X"04",X"CA",X"23",X"10",X"3A",X"9B",X"40",X"E6",X"F0",X"FE",X"50",
		X"DA",X"1B",X"10",X"3A",X"3C",X"42",X"FE",X"01",X"CA",X"23",X"10",X"3A",X"05",X"40",X"E6",X"01",
		X"C2",X"7F",X"10",X"3A",X"3B",X"42",X"FE",X"04",X"DA",X"7F",X"10",X"3A",X"3C",X"42",X"B7",X"CA",
		X"7F",X"10",X"3A",X"26",X"42",X"B7",X"C2",X"41",X"10",X"3A",X"27",X"42",X"FE",X"20",X"DA",X"7F",
		X"10",X"3A",X"3A",X"42",X"FE",X"03",X"CA",X"67",X"10",X"06",X"08",X"AF",X"32",X"39",X"42",X"00",
		X"CD",X"6B",X"11",X"3A",X"39",X"42",X"3C",X"32",X"39",X"42",X"05",X"C2",X"4F",X"10",X"CD",X"E7",
		X"10",X"CD",X"82",X"10",X"C3",X"7F",X"10",X"3A",X"3C",X"42",X"3D",X"0F",X"E6",X"03",X"32",X"39",
		X"42",X"CD",X"6B",X"11",X"3A",X"39",X"42",X"C6",X"04",X"32",X"39",X"42",X"CD",X"6B",X"11",X"CD",
		X"10",X"03",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DD",X"21",X"73",X"41",X"DD",X"7E",X"00",X"B7",
		X"C8",X"3A",X"4B",X"42",X"DD",X"86",X"04",X"DD",X"77",X"04",X"DD",X"7E",X"03",X"C6",X"08",X"DD",
		X"77",X"03",X"CD",X"42",X"11",X"DD",X"7E",X"03",X"FE",X"F7",X"D8",X"21",X"E0",X"53",X"06",X"20",
		X"36",X"24",X"23",X"05",X"C2",X"10",X"11",X"DD",X"36",X"00",X"00",X"AF",X"32",X"4D",X"42",X"FD",
		X"21",X"82",X"41",X"11",X"14",X"00",X"06",X"04",X"FD",X"7E",X"13",X"FE",X"FF",X"C2",X"39",X"11",
		X"FD",X"36",X"13",X"00",X"FD",X"36",X"27",X"00",X"C9",X"FD",X"19",X"FD",X"19",X"05",X"C2",X"28",
		X"11",X"C9",X"00",X"DD",X"7E",X"04",X"C6",X"04",X"47",X"DD",X"7E",X"03",X"0F",X"0F",X"E6",X"3E",
		X"21",X"00",X"58",X"5F",X"16",X"00",X"19",X"70",X"23",X"36",X"07",X"FD",X"21",X"E0",X"53",X"7B",
		X"0F",X"E6",X"1F",X"5F",X"FD",X"19",X"FD",X"36",X"00",X"81",X"C9",X"00",X"C5",X"DD",X"21",X"82",
		X"41",X"11",X"14",X"00",X"3A",X"39",X"42",X"B7",X"CA",X"81",X"11",X"DD",X"19",X"3D",X"C2",X"7B",
		X"11",X"DD",X"7E",X"00",X"B7",X"CA",X"E3",X"11",X"3A",X"4E",X"42",X"B7",X"CA",X"97",X"11",X"DD",
		X"36",X"05",X"05",X"DD",X"36",X"07",X"00",X"DD",X"7E",X"05",X"B7",X"CA",X"B6",X"11",X"3D",X"CA",
		X"BC",X"11",X"3D",X"CA",X"C2",X"11",X"3D",X"CA",X"C8",X"11",X"3D",X"CA",X"CE",X"11",X"3D",X"CA",
		X"D4",X"11",X"3D",X"CA",X"DA",X"11",X"CD",X"0E",X"12",X"C3",X"E0",X"11",X"CD",X"89",X"13",X"C3",
		X"E0",X"11",X"CD",X"C7",X"13",X"C3",X"E0",X"11",X"CD",X"A2",X"14",X"C3",X"E0",X"11",X"CD",X"14",
		X"16",X"C3",X"E0",X"11",X"CD",X"DC",X"16",X"C3",X"E0",X"11",X"CD",X"CD",X"17",X"C3",X"E0",X"11",
		X"CD",X"88",X"18",X"C1",X"C9",X"00",X"DD",X"7E",X"03",X"FE",X"08",X"DA",X"F7",X"11",X"DD",X"7E",
		X"04",X"FE",X"F4",X"D8",X"FE",X"FC",X"D0",X"DD",X"36",X"05",X"04",X"DD",X"36",X"07",X"00",X"DD",
		X"36",X"02",X"00",X"3A",X"3A",X"42",X"FE",X"03",X"C0",X"DD",X"36",X"03",X"00",X"C9",X"00",X"3A",
		X"3A",X"42",X"B7",X"CA",X"28",X"12",X"FE",X"01",X"CA",X"41",X"12",X"FE",X"02",X"CA",X"66",X"12",
		X"FE",X"03",X"CA",X"8B",X"12",X"C3",X"A4",X"12",X"DD",X"7E",X"07",X"B7",X"C2",X"3D",X"12",X"3A",
		X"3A",X"42",X"CD",X"92",X"08",X"FD",X"21",X"29",X"13",X"CD",X"BD",X"12",X"C9",X"CD",X"EF",X"12",
		X"C9",X"DD",X"7E",X"07",X"B7",X"C2",X"62",X"12",X"3A",X"3A",X"42",X"CD",X"92",X"08",X"3A",X"39",
		X"42",X"C6",X"08",X"CD",X"20",X"18",X"DD",X"36",X"04",X"78",X"DD",X"36",X"03",X"80",X"DD",X"36",
		X"01",X"24",X"CD",X"20",X"1A",X"C9",X"DD",X"7E",X"07",X"B7",X"C2",X"87",X"12",X"3A",X"3A",X"42",
		X"CD",X"92",X"08",X"3A",X"39",X"42",X"C6",X"10",X"CD",X"20",X"18",X"DD",X"36",X"04",X"78",X"DD",
		X"36",X"03",X"80",X"DD",X"36",X"01",X"24",X"CD",X"20",X"1A",X"C9",X"DD",X"7E",X"07",X"B7",X"C2",
		X"A0",X"12",X"3A",X"3A",X"42",X"CD",X"92",X"08",X"FD",X"21",X"49",X"13",X"CD",X"BD",X"12",X"C9",
		X"CD",X"EF",X"12",X"C9",X"DD",X"7E",X"07",X"B7",X"C2",X"B9",X"12",X"3A",X"3A",X"42",X"CD",X"92",
		X"08",X"FD",X"21",X"69",X"13",X"CD",X"BD",X"12",X"C9",X"CD",X"EF",X"12",X"C9",X"00",X"3A",X"39",
		X"42",X"07",X"07",X"E6",X"1C",X"5F",X"16",X"00",X"FD",X"19",X"FD",X"7E",X"00",X"DD",X"77",X"03",
		X"FD",X"7E",X"01",X"DD",X"77",X"04",X"FD",X"7E",X"02",X"DD",X"77",X"0A",X"FD",X"7E",X"03",X"DD",
		X"77",X"0B",X"DD",X"36",X"01",X"24",X"DD",X"36",X"06",X"10",X"DD",X"36",X"07",X"01",X"C9",X"DD",
		X"7E",X"06",X"E6",X"01",X"CA",X"FA",X"12",X"DD",X"35",X"01",X"DD",X"7E",X"03",X"DD",X"86",X"0A",
		X"DD",X"77",X"03",X"DD",X"7E",X"04",X"DD",X"86",X"0B",X"DD",X"77",X"04",X"DD",X"35",X"06",X"C0",
		X"3A",X"3A",X"42",X"B7",X"CA",X"20",X"13",X"DD",X"36",X"05",X"01",X"DD",X"36",X"07",X"00",X"C9",
		X"DD",X"36",X"05",X"02",X"DD",X"36",X"07",X"00",X"C9",X"60",X"70",X"FE",X"FE",X"60",X"70",X"FE",
		X"FE",X"60",X"78",X"FF",X"00",X"60",X"78",X"FF",X"00",X"60",X"80",X"FE",X"02",X"60",X"80",X"FE",
		X"02",X"58",X"78",X"FE",X"00",X"58",X"78",X"FE",X"00",X"30",X"20",X"06",X"04",X"20",X"B0",X"06",
		X"FD",X"20",X"40",X"06",X"03",X"50",X"90",X"06",X"FC",X"60",X"A0",X"06",X"FD",X"40",X"50",X"04",
		X"02",X"70",X"C0",X"05",X"FC",X"80",X"50",X"06",X"04",X"00",X"20",X"02",X"00",X"00",X"38",X"03",
		X"00",X"00",X"50",X"02",X"00",X"00",X"68",X"03",X"00",X"00",X"88",X"03",X"00",X"00",X"A0",X"02",
		X"00",X"00",X"B8",X"03",X"00",X"00",X"D0",X"02",X"00",X"00",X"3A",X"3A",X"42",X"FE",X"03",X"CA",
		X"BE",X"13",X"FE",X"04",X"CA",X"BE",X"13",X"DD",X"7E",X"07",X"B7",X"C2",X"B7",X"13",X"21",X"41",
		X"42",X"06",X"01",X"0E",X"00",X"3A",X"3A",X"42",X"FE",X"01",X"C2",X"AF",X"13",X"0E",X"50",X"CD",
		X"08",X"18",X"EE",X"01",X"CD",X"20",X"18",X"CD",X"20",X"1A",X"CD",X"E5",X"11",X"C9",X"DD",X"36",
		X"05",X"02",X"DD",X"36",X"07",X"00",X"C9",X"00",X"3A",X"3A",X"42",X"B7",X"CA",X"E1",X"13",X"FE",
		X"01",X"CA",X"2E",X"14",X"FE",X"02",X"CA",X"2E",X"14",X"FE",X"03",X"CA",X"66",X"14",X"C3",X"7C",
		X"14",X"DD",X"7E",X"07",X"B7",X"C2",X"F3",X"13",X"3A",X"27",X"42",X"0F",X"E6",X"01",X"C6",X"02",
		X"CD",X"20",X"18",X"DD",X"7E",X"13",X"FE",X"FF",X"C8",X"CD",X"20",X"1A",X"CD",X"E5",X"11",X"3A",
		X"39",X"42",X"E6",X"01",X"CA",X"1F",X"14",X"3A",X"9B",X"40",X"E6",X"F0",X"CA",X"1F",X"14",X"DD",
		X"E5",X"FD",X"E1",X"11",X"EC",X"FF",X"FD",X"19",X"FD",X"7E",X"00",X"B7",X"CA",X"25",X"14",X"3A",
		X"3C",X"42",X"FE",X"05",X"D0",X"DD",X"36",X"05",X"03",X"DD",X"36",X"07",X"00",X"C9",X"DD",X"7E",
		X"07",X"B7",X"C2",X"4F",X"14",X"3A",X"3D",X"42",X"47",X"3A",X"3E",X"42",X"B8",X"DA",X"56",X"14",
		X"21",X"42",X"42",X"06",X"07",X"0E",X"30",X"CD",X"08",X"18",X"EE",X"01",X"CD",X"20",X"18",X"CD",
		X"20",X"1A",X"CD",X"E5",X"11",X"C9",X"3A",X"3E",X"42",X"3C",X"32",X"3E",X"42",X"DD",X"36",X"05",
		X"03",X"DD",X"36",X"07",X"00",X"C9",X"DD",X"7E",X"03",X"DD",X"86",X"0A",X"DD",X"77",X"03",X"DD",
		X"7E",X"04",X"DD",X"86",X"0B",X"DD",X"77",X"04",X"CD",X"E5",X"11",X"C9",X"DD",X"7E",X"07",X"B7",
		X"C2",X"90",X"14",X"21",X"42",X"42",X"06",X"01",X"0E",X"52",X"CD",X"08",X"18",X"CD",X"20",X"18",
		X"CD",X"20",X"1A",X"CD",X"E5",X"11",X"3A",X"3D",X"42",X"47",X"3A",X"3E",X"42",X"B8",X"DA",X"56",
		X"14",X"C9",X"00",X"3A",X"3A",X"42",X"B7",X"CA",X"BA",X"14",X"FE",X"01",X"CA",X"BA",X"14",X"FE",
		X"02",X"CA",X"BA",X"14",X"FE",X"03",X"C8",X"C3",X"59",X"15",X"3A",X"9B",X"40",X"E6",X"F0",X"FE",
		X"C0",X"DA",X"CC",X"14",X"3A",X"3C",X"42",X"FE",X"01",X"CA",X"9B",X"15",X"DD",X"7E",X"07",X"B7",
		X"C2",X"45",X"15",X"3A",X"2B",X"42",X"D6",X"20",X"47",X"3A",X"2B",X"42",X"C6",X"20",X"4F",X"DD",
		X"7E",X"04",X"B8",X"DA",X"07",X"15",X"B9",X"D2",X"07",X"15",X"DD",X"7E",X"03",X"FE",X"80",X"DA",
		X"FA",X"14",X"FE",X"A0",X"D2",X"FA",X"14",X"C3",X"25",X"15",X"FE",X"60",X"DA",X"11",X"15",X"FE",
		X"80",X"D2",X"11",X"15",X"C3",X"1B",X"15",X"21",X"43",X"42",X"06",X"0F",X"0E",X"40",X"C3",X"2F",
		X"15",X"21",X"44",X"42",X"06",X"0F",X"0E",X"20",X"C3",X"2F",X"15",X"21",X"45",X"42",X"06",X"03",
		X"0E",X"20",X"C3",X"2F",X"15",X"21",X"46",X"42",X"06",X"03",X"0E",X"1C",X"C3",X"2F",X"15",X"CD",
		X"08",X"18",X"47",X"DD",X"7E",X"05",X"FE",X"02",X"C2",X"41",X"15",X"78",X"EE",X"01",X"C3",X"42",
		X"15",X"78",X"CD",X"20",X"18",X"CD",X"20",X"1A",X"CD",X"E5",X"11",X"DD",X"7E",X"05",X"FE",X"04",
		X"C0",X"3A",X"3E",X"42",X"3D",X"32",X"3E",X"42",X"C9",X"DD",X"7E",X"07",X"B7",X"C2",X"78",X"15",
		X"DD",X"36",X"0B",X"00",X"3A",X"9B",X"40",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"E6",X"03",X"C6",
		X"04",X"DD",X"77",X"0A",X"DD",X"36",X"07",X"01",X"DD",X"7E",X"04",X"DD",X"86",X"0B",X"DD",X"77",
		X"04",X"DD",X"7E",X"03",X"DD",X"86",X"0A",X"DD",X"77",X"03",X"CD",X"E5",X"11",X"DD",X"7E",X"05",
		X"FE",X"04",X"C0",X"3A",X"3E",X"42",X"3D",X"32",X"3E",X"42",X"C9",X"3A",X"3A",X"42",X"FE",X"01",
		X"CA",X"F9",X"15",X"DD",X"7E",X"07",X"B7",X"C2",X"F6",X"15",X"3A",X"46",X"42",X"3C",X"32",X"46",
		X"42",X"3A",X"2B",X"42",X"47",X"DD",X"7E",X"04",X"90",X"DA",X"CA",X"15",X"47",X"3A",X"46",X"42",
		X"F6",X"54",X"E6",X"55",X"32",X"46",X"42",X"C3",X"D7",X"15",X"2F",X"3C",X"47",X"3A",X"46",X"42",
		X"F6",X"56",X"E6",X"57",X"32",X"46",X"42",X"CD",X"20",X"18",X"3A",X"46",X"42",X"E6",X"01",X"C2",
		X"F6",X"15",X"78",X"0F",X"0F",X"0F",X"0F",X"0F",X"E6",X"07",X"C6",X"00",X"FE",X"02",X"D2",X"F3",
		X"15",X"3E",X"01",X"DD",X"77",X"11",X"C3",X"45",X"15",X"DD",X"7E",X"07",X"B7",X"C2",X"0D",X"16",
		X"21",X"46",X"42",X"06",X"07",X"0E",X"58",X"CD",X"08",X"18",X"CD",X"20",X"18",X"C3",X"45",X"15",
		X"00",X"00",X"00",X"00",X"00",X"3A",X"3A",X"42",X"B7",X"CA",X"2E",X"16",X"FE",X"01",X"CA",X"58",
		X"16",X"FE",X"02",X"CA",X"2E",X"16",X"FE",X"03",X"CA",X"6D",X"16",X"C3",X"81",X"16",X"DD",X"7E",
		X"07",X"B7",X"C2",X"54",X"16",X"3A",X"3A",X"42",X"CD",X"92",X"08",X"21",X"47",X"42",X"06",X"03",
		X"0E",X"18",X"CD",X"08",X"18",X"DD",X"36",X"04",X"78",X"DD",X"36",X"03",X"50",X"DD",X"36",X"01",
		X"24",X"CD",X"20",X"18",X"CD",X"20",X"1A",X"C9",X"DD",X"7E",X"07",X"B7",X"C2",X"69",X"16",X"3A",
		X"3A",X"42",X"CD",X"92",X"08",X"CD",X"A3",X"16",X"C9",X"CD",X"EF",X"12",X"C9",X"DD",X"36",X"05",
		X"00",X"DD",X"36",X"07",X"00",X"3A",X"3C",X"42",X"3D",X"32",X"3C",X"42",X"DD",X"36",X"00",X"00",
		X"C9",X"3A",X"3A",X"42",X"CD",X"92",X"08",X"DD",X"36",X"05",X"02",X"DD",X"36",X"07",X"00",X"FD",
		X"21",X"69",X"13",X"3A",X"2B",X"42",X"47",X"3A",X"27",X"42",X"E6",X"3F",X"D6",X"20",X"80",X"DD",
		X"77",X"04",X"C9",X"00",X"DD",X"7E",X"03",X"E6",X"3F",X"C6",X"40",X"DD",X"77",X"03",X"3A",X"3C",
		X"42",X"FE",X"01",X"C2",X"BD",X"16",X"DD",X"7E",X"03",X"E6",X"3F",X"C6",X"10",X"DD",X"7E",X"04",
		X"E6",X"3F",X"C6",X"50",X"DD",X"77",X"04",X"DD",X"36",X"0A",X"00",X"DD",X"36",X"0B",X"00",X"DD",
		X"36",X"01",X"24",X"DD",X"36",X"06",X"10",X"DD",X"36",X"07",X"01",X"C9",X"00",X"3A",X"3A",X"42",
		X"FE",X"03",X"CA",X"36",X"17",X"FE",X"04",X"CA",X"4C",X"17",X"DD",X"7E",X"07",X"B7",X"C2",X"00",
		X"17",X"DD",X"36",X"06",X"40",X"DD",X"36",X"07",X"01",X"3A",X"4E",X"42",X"3D",X"32",X"4E",X"42",
		X"DD",X"7E",X"01",X"FE",X"24",X"CA",X"0B",X"17",X"DD",X"34",X"01",X"DD",X"7E",X"04",X"2F",X"0F",
		X"0F",X"0F",X"0F",X"E6",X"0F",X"D6",X"08",X"DD",X"86",X"04",X"DD",X"77",X"04",X"DD",X"7E",X"03",
		X"2F",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"D6",X"08",X"DD",X"86",X"03",X"DD",X"77",X"03",X"DD",
		X"35",X"06",X"CA",X"8A",X"17",X"C9",X"DD",X"7E",X"07",X"B7",X"C2",X"6E",X"17",X"DD",X"36",X"06",
		X"80",X"DD",X"36",X"07",X"01",X"AF",X"32",X"4E",X"42",X"C3",X"6E",X"17",X"DD",X"7E",X"07",X"B7",
		X"C2",X"6E",X"17",X"DD",X"36",X"07",X"01",X"3A",X"4E",X"42",X"3D",X"32",X"4E",X"42",X"DD",X"36",
		X"06",X"80",X"DD",X"36",X"0A",X"02",X"DD",X"36",X"0B",X"00",X"DD",X"36",X"07",X"01",X"DD",X"7E",
		X"04",X"DD",X"86",X"0B",X"DD",X"77",X"04",X"DD",X"7E",X"03",X"DD",X"86",X"0A",X"DD",X"77",X"03",
		X"CD",X"B2",X"17",X"DD",X"35",X"06",X"CA",X"8A",X"17",X"C9",X"3E",X"01",X"32",X"04",X"40",X"3A",
		X"9B",X"40",X"32",X"9C",X"40",X"E6",X"F0",X"F6",X"01",X"32",X"9B",X"40",X"AF",X"32",X"26",X"42",
		X"32",X"27",X"42",X"3E",X"01",X"32",X"33",X"40",X"3E",X"40",X"CD",X"B2",X"02",X"AF",X"32",X"04",
		X"40",X"C9",X"00",X"DD",X"7E",X"03",X"FE",X"02",X"DA",X"C4",X"17",X"DD",X"7E",X"04",X"FE",X"F4",
		X"D8",X"FE",X"FC",X"D0",X"DD",X"36",X"05",X"06",X"DD",X"36",X"07",X"00",X"C9",X"00",X"DD",X"7E",
		X"07",X"B7",X"C2",X"DD",X"17",X"DD",X"36",X"06",X"80",X"DD",X"36",X"07",X"01",X"DD",X"35",X"06",
		X"CA",X"E4",X"17",X"C9",X"3E",X"01",X"32",X"04",X"40",X"3A",X"9B",X"40",X"32",X"9C",X"40",X"E6",
		X"F0",X"F6",X"01",X"32",X"9B",X"40",X"AF",X"32",X"26",X"42",X"32",X"27",X"42",X"3E",X"01",X"32",
		X"33",X"40",X"3E",X"40",X"CD",X"B2",X"02",X"C9",X"00",X"7E",X"C6",X"06",X"A0",X"77",X"E6",X"FE",
		X"81",X"4F",X"DD",X"7E",X"0F",X"FE",X"01",X"CA",X"1C",X"18",X"79",X"C9",X"79",X"F6",X"01",X"C9",
		X"00",X"FD",X"21",X"00",X"1C",X"57",X"07",X"07",X"07",X"E6",X"F8",X"5F",X"7A",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"E6",X"03",X"57",X"FD",X"19",X"FD",X"7E",X"00",X"DD",X"77",X"08",X"3A",X"3A",X"42",
		X"FE",X"01",X"CA",X"63",X"18",X"FE",X"03",X"CA",X"63",X"18",X"FE",X"04",X"CA",X"63",X"18",X"3A",
		X"40",X"41",X"FE",X"01",X"CA",X"63",X"18",X"3A",X"9B",X"40",X"E6",X"F0",X"C2",X"63",X"18",X"DD",
		X"36",X"08",X"02",X"FD",X"7E",X"01",X"DD",X"77",X"0D",X"FD",X"7E",X"02",X"DD",X"77",X"0E",X"FD",
		X"7E",X"03",X"DD",X"77",X"0F",X"FD",X"7E",X"04",X"DD",X"77",X"10",X"FD",X"7E",X"05",X"DD",X"77",
		X"11",X"FD",X"7E",X"06",X"DD",X"77",X"02",X"C9",X"00",X"21",X"A8",X"19",X"DD",X"7E",X"01",X"57",
		X"3A",X"3A",X"42",X"FE",X"04",X"C2",X"A2",X"18",X"DD",X"7E",X"05",X"FE",X"02",X"DA",X"A2",X"18",
		X"16",X"01",X"3A",X"3A",X"42",X"FE",X"03",X"C2",X"B2",X"18",X"7A",X"FE",X"1D",X"D2",X"B2",X"18",
		X"16",X"1D",X"7A",X"5F",X"16",X"00",X"19",X"FD",X"21",X"40",X"58",X"3A",X"3A",X"42",X"FE",X"03",
		X"CA",X"D2",X"18",X"3A",X"39",X"42",X"07",X"07",X"E6",X"FC",X"5F",X"16",X"00",X"FD",X"19",X"C3",
		X"DE",X"18",X"3A",X"39",X"42",X"E6",X"FC",X"CA",X"DE",X"18",X"FD",X"21",X"50",X"58",X"DD",X"7E",
		X"04",X"FD",X"77",X"00",X"7E",X"57",X"3A",X"3A",X"42",X"FE",X"01",X"C2",X"0F",X"19",X"DD",X"7E",
		X"02",X"E6",X"F0",X"FE",X"50",X"C2",X"0F",X"19",X"7A",X"C6",X"08",X"EE",X"07",X"57",X"DD",X"7E",
		X"0E",X"E6",X"18",X"FE",X"00",X"CA",X"0F",X"19",X"FE",X"18",X"CA",X"0F",X"19",X"16",X"E9",X"3A",
		X"3A",X"42",X"B7",X"C2",X"24",X"19",X"3A",X"39",X"42",X"E6",X"01",X"CA",X"24",X"19",X"7A",X"EE",
		X"40",X"EE",X"80",X"57",X"3A",X"3A",X"42",X"FE",X"04",X"C2",X"34",X"19",X"7A",X"F6",X"40",X"E6",
		X"F7",X"C6",X"08",X"57",X"7A",X"C6",X"20",X"FD",X"77",X"01",X"3A",X"3F",X"42",X"FD",X"77",X"02",
		X"DD",X"7E",X"05",X"FE",X"03",X"C2",X"4E",X"19",X"3A",X"40",X"42",X"FD",X"77",X"02",X"DD",X"7E",
		X"03",X"FD",X"77",X"03",X"3A",X"3A",X"42",X"FE",X"04",X"C0",X"DD",X"7E",X"13",X"B7",X"C8",X"2F",
		X"DD",X"E5",X"DD",X"21",X"40",X"58",X"07",X"07",X"E6",X"FC",X"5F",X"16",X"00",X"DD",X"19",X"DD",
		X"36",X"02",X"01",X"FD",X"7E",X"02",X"FE",X"02",X"C2",X"7F",X"19",X"DD",X"36",X"02",X"03",X"FD",
		X"7E",X"01",X"D6",X"08",X"DD",X"77",X"01",X"FD",X"7E",X"00",X"DD",X"77",X"00",X"FD",X"7E",X"03",
		X"C6",X"10",X"DD",X"77",X"03",X"FD",X"E1",X"FD",X"E5",X"FD",X"7E",X"05",X"FE",X"03",X"CA",X"A5",
		X"19",X"DD",X"36",X"01",X"09",X"DD",X"E1",X"C9",X"00",X"C1",X"C2",X"C3",X"C4",X"C5",X"C6",X"C7",
		X"87",X"86",X"85",X"84",X"83",X"82",X"81",X"01",X"02",X"03",X"04",X"05",X"06",X"07",X"47",X"46",
		X"45",X"44",X"43",X"42",X"41",X"08",X"09",X"0A",X"0B",X"0C",X"0D",X"0E",X"0F",X"00",X"FD",X"21",
		X"E8",X"19",X"3D",X"87",X"5F",X"16",X"00",X"FD",X"19",X"FD",X"7E",X"01",X"2F",X"3C",X"DD",X"77",
		X"0A",X"FD",X"7E",X"00",X"DD",X"77",X"0B",X"C9",X"00",X"FD",X"FF",X"FC",X"FD",X"FB",X"FC",X"FC",
		X"FB",X"FD",X"FC",X"FF",X"FD",X"00",X"FD",X"00",X"FC",X"01",X"FB",X"03",X"FC",X"04",X"FD",X"05",
		X"FF",X"04",X"00",X"03",X"00",X"03",X"01",X"04",X"03",X"05",X"04",X"04",X"05",X"03",X"04",X"01",
		X"03",X"00",X"03",X"00",X"04",X"FF",X"05",X"FD",X"04",X"FC",X"03",X"FB",X"01",X"FC",X"00",X"FD",
		X"00",X"DD",X"7E",X"07",X"B7",X"C2",X"35",X"1A",X"DD",X"7E",X"08",X"DD",X"77",X"09",X"DD",X"36",
		X"07",X"01",X"C3",X"38",X"1B",X"DD",X"7E",X"09",X"3D",X"DD",X"77",X"09",X"C0",X"DD",X"7E",X"08",
		X"DD",X"77",X"09",X"DD",X"7E",X"12",X"3D",X"DD",X"77",X"12",X"C2",X"64",X"1B",X"DD",X"35",X"0E",
		X"C2",X"71",X"1A",X"DD",X"36",X"07",X"00",X"DD",X"7E",X"05",X"FE",X"00",X"CA",X"6C",X"1A",X"FE",
		X"01",X"CA",X"6C",X"1A",X"FE",X"04",X"C0",X"DD",X"36",X"05",X"01",X"C9",X"3C",X"DD",X"77",X"05",
		X"C9",X"DD",X"7E",X"0E",X"E6",X"07",X"FE",X"02",X"C2",X"8B",X"1A",X"DD",X"7E",X"02",X"E6",X"0F",
		X"CA",X"8B",X"1A",X"FE",X"05",X"D2",X"8B",X"1A",X"DD",X"35",X"0E",X"DD",X"7E",X"0D",X"DD",X"86",
		X"0F",X"C2",X"96",X"1A",X"3E",X"1C",X"FE",X"1D",X"C2",X"9D",X"1A",X"3E",X"01",X"DD",X"77",X"0D",
		X"DD",X"7E",X"0E",X"E6",X"03",X"C2",X"1D",X"1B",X"DD",X"7E",X"0E",X"E6",X"07",X"C2",X"10",X"1B",
		X"DD",X"7E",X"0E",X"E6",X"0F",X"C2",X"EC",X"1A",X"DD",X"7E",X"02",X"E6",X"0F",X"FE",X"02",X"CA",
		X"CF",X"1A",X"FE",X"03",X"CA",X"D8",X"1A",X"FE",X"04",X"CA",X"E1",X"1A",X"C3",X"EC",X"1A",X"DD",
		X"34",X"10",X"DD",X"34",X"11",X"C3",X"EC",X"1A",X"DD",X"35",X"10",X"DD",X"35",X"11",X"C3",X"EC",
		X"1A",X"DD",X"7E",X"0F",X"2F",X"3C",X"DD",X"77",X"0F",X"C3",X"EC",X"1A",X"DD",X"7E",X"02",X"E6",
		X"0F",X"FE",X"06",X"CA",X"FE",X"1A",X"FE",X"07",X"CA",X"07",X"1B",X"C3",X"10",X"1B",X"DD",X"34",
		X"10",X"DD",X"34",X"11",X"C3",X"10",X"1B",X"DD",X"35",X"10",X"DD",X"35",X"11",X"C3",X"10",X"1B",
		X"DD",X"7E",X"02",X"E6",X"F0",X"FE",X"20",X"C2",X"1D",X"1B",X"DD",X"35",X"01",X"DD",X"7E",X"02",
		X"E6",X"F0",X"FE",X"10",X"CA",X"35",X"1B",X"FE",X"20",X"CA",X"38",X"1B",X"DD",X"7E",X"0D",X"DD",
		X"77",X"01",X"C3",X"38",X"1B",X"DD",X"35",X"01",X"DD",X"7E",X"0D",X"CD",X"CD",X"19",X"DD",X"7E",
		X"0D",X"D6",X"04",X"DA",X"55",X"1B",X"D6",X"07",X"DA",X"5E",X"1B",X"D6",X"07",X"DA",X"55",X"1B",
		X"D6",X"07",X"DA",X"5E",X"1B",X"DD",X"7E",X"10",X"DD",X"77",X"12",X"C3",X"64",X"1B",X"DD",X"7E",
		X"11",X"DD",X"77",X"12",X"DD",X"7E",X"03",X"DD",X"86",X"0A",X"DD",X"77",X"03",X"DD",X"7E",X"04",
		X"DD",X"86",X"0B",X"DD",X"77",X"04",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"0F",X"09",X"01",X"03",X"03",X"00",X"00",X"01",X"0F",X"09",X"FF",X"03",X"03",X"00",X"00",
		X"01",X"01",X"1E",X"01",X"01",X"02",X"00",X"00",X"01",X"01",X"1E",X"FF",X"01",X"02",X"00",X"00",
		X"02",X"08",X"09",X"01",X"01",X"01",X"10",X"00",X"02",X"16",X"09",X"FF",X"01",X"01",X"10",X"00",
		X"01",X"08",X"09",X"01",X"02",X"02",X"10",X"00",X"01",X"16",X"09",X"FF",X"02",X"02",X"10",X"00",
		X"04",X"08",X"09",X"01",X"01",X"01",X"10",X"00",X"04",X"16",X"09",X"FF",X"01",X"01",X"10",X"00",
		X"02",X"08",X"09",X"01",X"02",X"02",X"10",X"00",X"02",X"16",X"09",X"FF",X"02",X"02",X"10",X"00",
		X"01",X"08",X"09",X"01",X"03",X"03",X"10",X"00",X"01",X"16",X"09",X"FF",X"03",X"03",X"10",X"00",
		X"01",X"08",X"09",X"01",X"04",X"04",X"10",X"00",X"01",X"16",X"09",X"FF",X"04",X"04",X"10",X"00",
		X"04",X"08",X"09",X"01",X"01",X"01",X"10",X"00",X"04",X"16",X"09",X"FF",X"01",X"01",X"10",X"00",
		X"02",X"08",X"09",X"01",X"02",X"02",X"10",X"00",X"02",X"16",X"09",X"FF",X"02",X"02",X"10",X"00",
		X"02",X"08",X"09",X"01",X"01",X"03",X"10",X"00",X"02",X"16",X"09",X"FF",X"01",X"03",X"10",X"00",
		X"02",X"08",X"09",X"01",X"02",X"04",X"10",X"00",X"02",X"16",X"09",X"FF",X"02",X"04",X"10",X"00",
		X"01",X"0F",X"1F",X"01",X"01",X"01",X"22",X"00",X"01",X"0F",X"1F",X"FF",X"01",X"01",X"22",X"00",
		X"01",X"01",X"2F",X"01",X"01",X"01",X"22",X"00",X"01",X"01",X"2F",X"FF",X"01",X"01",X"22",X"00",
		X"01",X"16",X"3F",X"01",X"04",X"04",X"03",X"00",X"01",X"08",X"3F",X"FF",X"04",X"04",X"03",X"00",
		X"01",X"16",X"3F",X"01",X"04",X"04",X"03",X"00",X"01",X"08",X"3F",X"FF",X"04",X"04",X"03",X"00",
		X"01",X"16",X"1F",X"01",X"04",X"04",X"07",X"00",X"01",X"08",X"1F",X"FF",X"04",X"04",X"07",X"00",
		X"01",X"16",X"1F",X"01",X"04",X"04",X"07",X"00",X"01",X"08",X"1F",X"FF",X"04",X"04",X"07",X"00",
		X"01",X"16",X"7F",X"01",X"01",X"01",X"04",X"00",X"01",X"08",X"7F",X"FF",X"01",X"01",X"04",X"00",
		X"01",X"16",X"7F",X"01",X"01",X"01",X"04",X"00",X"01",X"08",X"7F",X"FF",X"01",X"01",X"04",X"00",
		X"01",X"16",X"7F",X"01",X"02",X"01",X"04",X"00",X"01",X"08",X"7F",X"FF",X"02",X"01",X"04",X"00",
		X"01",X"16",X"7F",X"01",X"02",X"01",X"04",X"00",X"01",X"08",X"7F",X"FF",X"02",X"01",X"04",X"00",
		X"01",X"16",X"7F",X"01",X"03",X"01",X"04",X"00",X"01",X"08",X"7F",X"FF",X"03",X"01",X"04",X"00",
		X"01",X"16",X"7F",X"01",X"03",X"01",X"04",X"00",X"01",X"08",X"7F",X"FF",X"03",X"01",X"04",X"00",
		X"01",X"08",X"1D",X"01",X"02",X"02",X"00",X"00",X"01",X"08",X"1D",X"FF",X"02",X"02",X"00",X"00",
		X"01",X"16",X"1D",X"01",X"02",X"02",X"00",X"00",X"01",X"08",X"1D",X"FF",X"02",X"02",X"00",X"00",
		X"01",X"16",X"1D",X"01",X"03",X"02",X"00",X"00",X"01",X"08",X"1D",X"FF",X"03",X"02",X"00",X"00",
		X"01",X"16",X"1D",X"01",X"03",X"02",X"00",X"00",X"01",X"08",X"1D",X"FF",X"03",X"02",X"00",X"00",
		X"01",X"16",X"1D",X"01",X"04",X"03",X"00",X"00",X"01",X"08",X"1D",X"FF",X"04",X"03",X"00",X"00",
		X"01",X"16",X"1D",X"01",X"04",X"03",X"00",X"00",X"01",X"08",X"1D",X"FF",X"04",X"03",X"00",X"00",
		X"01",X"16",X"1D",X"01",X"05",X"03",X"00",X"00",X"01",X"08",X"1D",X"FF",X"05",X"03",X"00",X"00",
		X"01",X"16",X"1D",X"01",X"05",X"03",X"00",X"00",X"01",X"08",X"1D",X"FF",X"05",X"03",X"00",X"00",
		X"01",X"16",X"0F",X"01",X"01",X"01",X"06",X"00",X"01",X"08",X"0F",X"FF",X"01",X"01",X"06",X"00",
		X"01",X"16",X"0F",X"01",X"02",X"01",X"06",X"00",X"01",X"08",X"0F",X"FF",X"02",X"01",X"06",X"00",
		X"01",X"16",X"0F",X"01",X"02",X"02",X"07",X"00",X"01",X"08",X"0F",X"FF",X"02",X"02",X"07",X"00",
		X"01",X"16",X"0F",X"01",X"04",X"02",X"07",X"00",X"01",X"08",X"0F",X"FF",X"04",X"02",X"07",X"00",
		X"01",X"16",X"0F",X"01",X"01",X"02",X"06",X"00",X"01",X"08",X"0F",X"FF",X"01",X"02",X"06",X"00",
		X"01",X"16",X"0F",X"01",X"01",X"03",X"06",X"00",X"01",X"08",X"0F",X"FF",X"01",X"03",X"06",X"00",
		X"01",X"16",X"0F",X"01",X"02",X"04",X"07",X"00",X"01",X"08",X"0F",X"FF",X"02",X"04",X"07",X"00",
		X"01",X"16",X"0F",X"01",X"02",X"06",X"07",X"00",X"01",X"08",X"0F",X"FF",X"02",X"06",X"07",X"00",
		X"01",X"0F",X"09",X"01",X"01",X"01",X"00",X"00",X"01",X"0F",X"09",X"01",X"01",X"01",X"00",X"00",
		X"02",X"04",X"08",X"01",X"02",X"02",X"60",X"00",X"02",X"1A",X"08",X"FF",X"02",X"02",X"60",X"00",
		X"01",X"19",X"11",X"01",X"03",X"03",X"00",X"00",X"01",X"0F",X"07",X"01",X"01",X"01",X"00",X"00",
		X"01",X"08",X"15",X"FF",X"03",X"03",X"00",X"00",X"01",X"01",X"07",X"FF",X"01",X"01",X"00",X"00",
		X"01",X"16",X"1F",X"01",X"02",X"03",X"54",X"00",X"01",X"16",X"1F",X"01",X"01",X"03",X"54",X"00",
		X"01",X"16",X"1F",X"01",X"01",X"01",X"54",X"00",X"01",X"16",X"1F",X"01",X"02",X"03",X"54",X"00",
		X"01",X"16",X"1F",X"01",X"02",X"04",X"54",X"00",X"01",X"16",X"1F",X"01",X"01",X"04",X"54",X"00",
		X"01",X"16",X"1F",X"01",X"02",X"02",X"54",X"00",X"01",X"16",X"1F",X"01",X"01",X"02",X"54",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"3A",X"3B",X"42",X"FE",X"04",X"DA",X"12",X"20",X"CD",X"DD",X"23",X"CD",X"20",X"20",X"CD",
		X"6B",X"21",X"3A",X"3B",X"42",X"FE",X"03",X"C2",X"1D",X"20",X"CD",X"50",X"22",X"CD",X"10",X"03",
		X"00",X"11",X"14",X"00",X"01",X"04",X"04",X"DD",X"21",X"40",X"41",X"DD",X"7E",X"00",X"FE",X"01",
		X"C2",X"7B",X"20",X"FD",X"21",X"82",X"41",X"26",X"08",X"2E",X"01",X"FD",X"7E",X"00",X"B7",X"CA",
		X"75",X"20",X"DD",X"7E",X"04",X"D6",X"0E",X"80",X"FD",X"BE",X"04",X"D2",X"75",X"20",X"DD",X"7E",
		X"04",X"C6",X"0F",X"90",X"FD",X"BE",X"04",X"DA",X"75",X"20",X"DD",X"7E",X"03",X"D6",X"08",X"81",
		X"FD",X"BE",X"03",X"D2",X"75",X"20",X"DD",X"7E",X"03",X"C6",X"10",X"91",X"FD",X"BE",X"03",X"DA",
		X"75",X"20",X"C3",X"24",X"21",X"FD",X"19",X"25",X"C2",X"3B",X"20",X"DD",X"21",X"45",X"41",X"DD",
		X"7E",X"00",X"FE",X"01",X"C2",X"CF",X"20",X"FD",X"21",X"82",X"41",X"26",X"08",X"2E",X"02",X"FD",
		X"7E",X"00",X"B7",X"CA",X"C9",X"20",X"DD",X"7E",X"04",X"D6",X"0A",X"80",X"FD",X"BE",X"04",X"D2",
		X"C9",X"20",X"DD",X"7E",X"04",X"C6",X"1B",X"90",X"FD",X"BE",X"04",X"DA",X"C9",X"20",X"DD",X"7E",
		X"03",X"D6",X"08",X"81",X"FD",X"BE",X"03",X"D2",X"C9",X"20",X"DD",X"7E",X"03",X"C6",X"10",X"91",
		X"FD",X"BE",X"03",X"DA",X"C9",X"20",X"C3",X"24",X"21",X"FD",X"19",X"25",X"C2",X"8F",X"20",X"DD",
		X"21",X"4A",X"41",X"DD",X"7E",X"00",X"FE",X"01",X"C2",X"23",X"21",X"FD",X"21",X"82",X"41",X"26",
		X"08",X"2E",X"03",X"FD",X"7E",X"00",X"B7",X"CA",X"1D",X"21",X"DD",X"7E",X"04",X"D6",X"0F",X"80",
		X"FD",X"BE",X"04",X"D2",X"1D",X"21",X"DD",X"7E",X"04",X"C6",X"20",X"90",X"FD",X"BE",X"04",X"DA",
		X"1D",X"21",X"DD",X"7E",X"03",X"D6",X"10",X"81",X"FD",X"BE",X"03",X"D2",X"1D",X"21",X"DD",X"7E",
		X"03",X"C6",X"10",X"91",X"FD",X"BE",X"03",X"DA",X"1D",X"21",X"C3",X"24",X"21",X"FD",X"19",X"25",
		X"C2",X"E3",X"20",X"C9",X"3E",X"01",X"32",X"04",X"40",X"FD",X"36",X"02",X"00",X"7D",X"CD",X"0A",
		X"27",X"3A",X"40",X"41",X"FE",X"01",X"C2",X"3E",X"21",X"3E",X"03",X"32",X"40",X"41",X"3A",X"45",
		X"41",X"FE",X"01",X"C2",X"4B",X"21",X"3E",X"03",X"32",X"45",X"41",X"3A",X"4A",X"41",X"FE",X"01",
		X"C2",X"58",X"21",X"3E",X"03",X"32",X"4A",X"41",X"00",X"AF",X"32",X"28",X"42",X"32",X"29",X"42",
		X"3A",X"3C",X"42",X"32",X"4E",X"42",X"AF",X"32",X"04",X"40",X"C9",X"C9",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DD",X"21",X"45",X"41",X"DD",X"7E",X"00",
		X"FE",X"01",X"C2",X"FF",X"21",X"FD",X"7E",X"00",X"B7",X"CA",X"FF",X"21",X"DD",X"7E",X"04",X"C6",
		X"06",X"80",X"FD",X"BE",X"04",X"D2",X"FF",X"21",X"DD",X"7E",X"04",X"C6",X"1B",X"90",X"FD",X"BE",
		X"04",X"DA",X"FF",X"21",X"DD",X"7E",X"03",X"C6",X"04",X"81",X"FD",X"BE",X"03",X"D2",X"FF",X"21",
		X"DD",X"7E",X"03",X"C6",X"10",X"91",X"FD",X"BE",X"03",X"DA",X"FF",X"21",X"C3",X"46",X"22",X"DD",
		X"21",X"4A",X"41",X"DD",X"7E",X"00",X"FE",X"01",X"C2",X"45",X"22",X"FD",X"7E",X"00",X"B7",X"CA",
		X"45",X"22",X"DD",X"7E",X"04",X"C6",X"01",X"80",X"FD",X"BE",X"04",X"D2",X"45",X"22",X"DD",X"7E",
		X"04",X"C6",X"20",X"90",X"FD",X"BE",X"04",X"DA",X"45",X"22",X"DD",X"7E",X"03",X"D6",X"04",X"81",
		X"FD",X"BE",X"03",X"D2",X"45",X"22",X"DD",X"7E",X"03",X"C6",X"10",X"91",X"FD",X"BE",X"03",X"DA",
		X"45",X"22",X"C3",X"46",X"22",X"C9",X"AF",X"32",X"4D",X"42",X"3E",X"FF",X"32",X"2D",X"42",X"C9",
		X"3A",X"4A",X"41",X"FE",X"01",X"CA",X"DC",X"23",X"3A",X"45",X"41",X"FE",X"01",X"CA",X"6B",X"22",
		X"3A",X"40",X"41",X"FE",X"01",X"CA",X"76",X"22",X"C3",X"DC",X"23",X"3A",X"4A",X"41",X"FE",X"02",
		X"CA",X"EF",X"22",X"C3",X"DC",X"23",X"3A",X"45",X"41",X"FE",X"02",X"CA",X"89",X"22",X"3A",X"4A",
		X"41",X"FE",X"02",X"CA",X"7C",X"23",X"C3",X"DC",X"23",X"06",X"06",X"0E",X"1B",X"16",X"02",X"1E",
		X"0F",X"26",X"0A",X"2E",X"0A",X"DD",X"21",X"45",X"41",X"FD",X"21",X"40",X"41",X"CD",X"40",X"25",
		X"B7",X"C2",X"BA",X"22",X"06",X"0D",X"0E",X"13",X"16",X"05",X"1E",X"0B",X"26",X"08",X"2E",X"10",
		X"CD",X"FC",X"24",X"B7",X"C2",X"D2",X"22",X"C3",X"DC",X"23",X"AF",X"32",X"40",X"41",X"3A",X"97",
		X"40",X"3D",X"32",X"97",X"40",X"3E",X"01",X"CD",X"84",X"25",X"3E",X"01",X"32",X"45",X"41",X"C3",
		X"DC",X"23",X"3E",X"01",X"32",X"45",X"41",X"3A",X"48",X"41",X"D6",X"08",X"32",X"43",X"41",X"3A",
		X"49",X"41",X"C6",X"08",X"32",X"44",X"41",X"3E",X"01",X"CD",X"E5",X"25",X"C3",X"DC",X"23",X"06",
		X"01",X"0E",X"20",X"16",X"06",X"1E",X"1B",X"26",X"02",X"2E",X"0A",X"DD",X"21",X"4A",X"41",X"FD",
		X"21",X"45",X"41",X"CD",X"40",X"25",X"B7",X"C2",X"20",X"23",X"06",X"0D",X"0E",X"13",X"16",X"0D",
		X"1E",X"13",X"26",X"00",X"2E",X"10",X"CD",X"FC",X"24",X"B7",X"C2",X"4A",X"23",X"C3",X"DC",X"23",
		X"3A",X"40",X"41",X"FE",X"01",X"C2",X"2F",X"23",X"3A",X"97",X"40",X"3D",X"32",X"97",X"40",X"AF",
		X"32",X"40",X"41",X"32",X"45",X"41",X"3A",X"97",X"40",X"3D",X"32",X"97",X"40",X"3E",X"02",X"CD",
		X"84",X"25",X"3E",X"01",X"32",X"4A",X"41",X"C3",X"DC",X"23",X"3E",X"01",X"32",X"4A",X"41",X"3A",
		X"4D",X"41",X"D6",X"10",X"32",X"48",X"41",X"D6",X"08",X"32",X"43",X"41",X"3A",X"4E",X"41",X"32",
		X"49",X"41",X"C6",X"08",X"32",X"44",X"41",X"3A",X"40",X"41",X"FE",X"01",X"CA",X"74",X"23",X"3E",
		X"02",X"C3",X"76",X"23",X"3E",X"03",X"CD",X"E5",X"25",X"C3",X"DC",X"23",X"06",X"01",X"0E",X"20",
		X"16",X"02",X"1E",X"0F",X"26",X"02",X"2E",X"0A",X"DD",X"21",X"4A",X"41",X"FD",X"21",X"40",X"41",
		X"CD",X"40",X"25",X"B7",X"C2",X"C7",X"23",X"06",X"0D",X"0E",X"13",X"16",X"05",X"1E",X"0B",X"26",
		X"00",X"2E",X"10",X"CD",X"FC",X"24",X"B7",X"CA",X"DC",X"23",X"3E",X"01",X"32",X"4A",X"41",X"3A",
		X"4D",X"41",X"D6",X"10",X"32",X"43",X"41",X"3A",X"4E",X"41",X"C6",X"08",X"32",X"44",X"41",X"3E",
		X"02",X"CD",X"E5",X"25",X"C3",X"DC",X"23",X"AF",X"32",X"40",X"41",X"3A",X"97",X"40",X"3D",X"32",
		X"97",X"40",X"3E",X"01",X"CD",X"84",X"25",X"3E",X"01",X"32",X"4A",X"41",X"C9",X"00",X"26",X"05",
		X"DD",X"21",X"59",X"41",X"2E",X"08",X"FD",X"21",X"82",X"41",X"11",X"14",X"00",X"DD",X"7E",X"00",
		X"B7",X"CA",X"44",X"24",X"FD",X"7E",X"00",X"B7",X"CA",X"3E",X"24",X"3A",X"3A",X"42",X"FE",X"04",
		X"CA",X"17",X"24",X"DD",X"7E",X"04",X"FD",X"BE",X"04",X"DA",X"3E",X"24",X"D6",X"10",X"FD",X"BE",
		X"04",X"D2",X"3E",X"24",X"C3",X"2A",X"24",X"DD",X"7E",X"04",X"D6",X"04",X"FD",X"BE",X"04",X"DA",
		X"3E",X"24",X"D6",X"08",X"FD",X"BE",X"04",X"D2",X"3E",X"24",X"DD",X"7E",X"03",X"FD",X"BE",X"03",
		X"DA",X"3E",X"24",X"D6",X"0C",X"FD",X"BE",X"03",X"D2",X"3E",X"24",X"C3",X"4E",X"24",X"FD",X"19",
		X"2D",X"C2",X"F4",X"23",X"11",X"05",X"00",X"DD",X"19",X"25",X"C2",X"E4",X"23",X"C9",X"DD",X"36",
		X"04",X"00",X"FD",X"7E",X"05",X"FE",X"03",X"C2",X"61",X"24",X"3A",X"3E",X"42",X"3D",X"32",X"3E",
		X"42",X"3A",X"3A",X"42",X"C6",X"05",X"CD",X"92",X"08",X"3A",X"3A",X"42",X"B7",X"C2",X"7E",X"24",
		X"7D",X"E6",X"01",X"C2",X"7E",X"24",X"FD",X"36",X"19",X"02",X"FD",X"36",X"1B",X"00",X"3A",X"3A",
		X"42",X"FE",X"03",X"CA",X"B9",X"24",X"3E",X"08",X"95",X"CD",X"3A",X"28",X"01",X"00",X"01",X"3A",
		X"3A",X"42",X"FE",X"00",X"CA",X"A7",X"24",X"FE",X"01",X"CA",X"AD",X"24",X"FE",X"02",X"CA",X"B3",
		X"24",X"01",X"00",X"01",X"C3",X"C2",X"24",X"01",X"50",X"00",X"C3",X"C2",X"24",X"01",X"60",X"00",
		X"C3",X"C2",X"24",X"01",X"30",X"00",X"C3",X"C2",X"24",X"3E",X"08",X"95",X"CD",X"BB",X"28",X"01",
		X"00",X"02",X"CD",X"C9",X"24",X"CD",X"E8",X"26",X"C9",X"00",X"3A",X"35",X"40",X"B7",X"C8",X"21",
		X"9A",X"40",X"79",X"86",X"27",X"77",X"2B",X"78",X"8E",X"27",X"77",X"2B",X"3E",X"00",X"8E",X"27",
		X"77",X"47",X"3A",X"3D",X"40",X"B8",X"C0",X"3A",X"9E",X"40",X"B7",X"C0",X"3A",X"9D",X"40",X"B7",
		X"C0",X"3E",X"10",X"CD",X"92",X"08",X"3E",X"01",X"32",X"9D",X"40",X"C9",X"00",X"DD",X"7E",X"00",
		X"FE",X"02",X"C2",X"3E",X"25",X"FD",X"7E",X"00",X"FE",X"01",X"C2",X"3E",X"25",X"DD",X"7E",X"04",
		X"80",X"93",X"FD",X"BE",X"04",X"D2",X"3E",X"25",X"DD",X"7E",X"04",X"81",X"92",X"FD",X"BE",X"04",
		X"DA",X"3E",X"25",X"DD",X"7E",X"03",X"84",X"D6",X"0F",X"FD",X"BE",X"03",X"D2",X"3E",X"25",X"DD",
		X"7E",X"03",X"C6",X"11",X"95",X"FD",X"BE",X"03",X"DA",X"3E",X"25",X"3E",X"01",X"C9",X"AF",X"C9",
		X"00",X"DD",X"7E",X"00",X"FE",X"02",X"C2",X"82",X"25",X"FD",X"7E",X"00",X"FE",X"01",X"C2",X"82",
		X"25",X"DD",X"7E",X"04",X"80",X"93",X"FD",X"BE",X"04",X"D2",X"82",X"25",X"DD",X"7E",X"04",X"81",
		X"92",X"FD",X"BE",X"04",X"DA",X"82",X"25",X"DD",X"7E",X"03",X"84",X"D6",X"0E",X"FD",X"BE",X"03",
		X"D2",X"82",X"25",X"DD",X"7E",X"03",X"C6",X"0E",X"95",X"FD",X"BE",X"03",X"DA",X"82",X"25",X"3E",
		X"01",X"C9",X"AF",X"C9",X"00",X"F5",X"3E",X"01",X"32",X"04",X"40",X"F1",X"CD",X"0A",X"27",X"3E",
		X"0C",X"CD",X"92",X"08",X"11",X"CD",X"25",X"CD",X"80",X"09",X"C3",X"70",X"29",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"3E",X"06",X"CD",X"C3",X"2A",X"3E",X"08",X"CD",X"C3",X"2A",X"3E",X"17",
		X"CD",X"C3",X"2A",X"AF",X"32",X"28",X"42",X"32",X"29",X"42",X"3A",X"9B",X"40",X"3C",X"32",X"9B",
		X"40",X"AF",X"32",X"26",X"42",X"32",X"27",X"42",X"AF",X"32",X"04",X"40",X"C9",X"0C",X"06",X"07",
		X"1C",X"18",X"1B",X"1B",X"22",X"24",X"17",X"18",X"24",X"0B",X"18",X"17",X"1E",X"1C",X"24",X"24",
		X"24",X"24",X"24",X"24",X"FF",X"00",X"32",X"32",X"42",X"3E",X"01",X"32",X"04",X"40",X"3A",X"40",
		X"41",X"FE",X"01",X"C2",X"FB",X"25",X"3E",X"01",X"CD",X"87",X"34",X"3A",X"45",X"41",X"FE",X"01",
		X"C2",X"08",X"26",X"3E",X"02",X"CD",X"87",X"34",X"3A",X"4A",X"41",X"FE",X"01",X"C2",X"15",X"26",
		X"3E",X"03",X"CD",X"87",X"34",X"00",X"3E",X"0B",X"CD",X"92",X"08",X"11",X"AD",X"26",X"CD",X"80",
		X"09",X"11",X"BB",X"26",X"CD",X"80",X"09",X"11",X"CF",X"26",X"CD",X"80",X"09",X"11",X"DB",X"26",
		X"CD",X"DD",X"09",X"3A",X"30",X"42",X"B7",X"CA",X"55",X"26",X"47",X"3A",X"32",X"42",X"4F",X"AF",
		X"32",X"32",X"42",X"3A",X"32",X"42",X"81",X"27",X"32",X"32",X"42",X"78",X"3D",X"27",X"47",X"C2",
		X"43",X"26",X"C3",X"59",X"26",X"AF",X"32",X"32",X"42",X"11",X"E1",X"26",X"CD",X"DD",X"09",X"3E",
		X"FF",X"CD",X"B2",X"02",X"3E",X"FF",X"CD",X"B2",X"02",X"3E",X"FF",X"CD",X"B2",X"02",X"3E",X"FF",
		X"CD",X"B2",X"02",X"3E",X"FF",X"CD",X"B2",X"02",X"3E",X"06",X"CD",X"C3",X"2A",X"3E",X"08",X"CD",
		X"C3",X"2A",X"3E",X"17",X"CD",X"C3",X"2A",X"3A",X"32",X"42",X"47",X"0E",X"00",X"CD",X"C9",X"24",
		X"CD",X"E8",X"26",X"3A",X"9B",X"40",X"3C",X"32",X"9B",X"40",X"AF",X"32",X"26",X"42",X"32",X"27",
		X"42",X"AF",X"32",X"28",X"42",X"32",X"29",X"42",X"AF",X"32",X"04",X"40",X"C9",X"02",X"17",X"09",
		X"1B",X"12",X"10",X"11",X"1D",X"24",X"18",X"17",X"24",X"28",X"FF",X"04",X"06",X"07",X"0D",X"18",
		X"0C",X"14",X"12",X"17",X"10",X"24",X"0B",X"18",X"17",X"1E",X"1C",X"24",X"24",X"24",X"FF",X"04",
		X"08",X"0C",X"24",X"2A",X"24",X"24",X"24",X"24",X"24",X"2E",X"FF",X"04",X"08",X"0F",X"32",X"42",
		X"03",X"04",X"08",X"15",X"32",X"42",X"04",X"C9",X"00",X"3A",X"40",X"40",X"B7",X"C2",X"F7",X"26",
		X"11",X"FE",X"26",X"CD",X"DD",X"09",X"C9",X"11",X"04",X"27",X"CD",X"DD",X"09",X"C9",X"07",X"01",
		X"00",X"98",X"40",X"06",X"07",X"01",X"16",X"98",X"40",X"06",X"00",X"3D",X"CA",X"17",X"27",X"3D",
		X"CA",X"2A",X"27",X"3D",X"CA",X"35",X"27",X"DD",X"21",X"40",X"41",X"DD",X"7E",X"04",X"D6",X"08",
		X"DD",X"77",X"04",X"FD",X"21",X"40",X"58",X"C3",X"3D",X"27",X"DD",X"21",X"45",X"41",X"FD",X"21",
		X"44",X"58",X"C3",X"3D",X"27",X"DD",X"21",X"4A",X"41",X"FD",X"21",X"4C",X"58",X"CD",X"50",X"29",
		X"AF",X"32",X"4F",X"41",X"32",X"59",X"41",X"32",X"5E",X"41",X"32",X"63",X"41",X"32",X"68",X"41",
		X"32",X"6D",X"41",X"CD",X"21",X"28",X"CD",X"10",X"28",X"3E",X"01",X"CD",X"32",X"09",X"3A",X"4D",
		X"42",X"FE",X"01",X"CA",X"6A",X"27",X"FD",X"21",X"50",X"58",X"DD",X"7E",X"03",X"D6",X"08",X"DD",
		X"77",X"03",X"DD",X"36",X"00",X"00",X"21",X"FC",X"27",X"06",X"05",X"00",X"FD",X"21",X"50",X"58",
		X"DD",X"7E",X"04",X"FD",X"77",X"00",X"7E",X"FD",X"77",X"01",X"FD",X"36",X"02",X"0C",X"DD",X"7E",
		X"03",X"FD",X"77",X"03",X"FD",X"21",X"54",X"58",X"DD",X"7E",X"04",X"C6",X"10",X"FD",X"77",X"00",
		X"23",X"7E",X"FD",X"77",X"01",X"FD",X"36",X"02",X"0C",X"DD",X"7E",X"03",X"FD",X"77",X"03",X"FD",
		X"21",X"58",X"58",X"DD",X"7E",X"04",X"FD",X"77",X"00",X"23",X"7E",X"FD",X"77",X"01",X"FD",X"36",
		X"02",X"0C",X"DD",X"7E",X"03",X"C6",X"10",X"FD",X"77",X"03",X"FD",X"21",X"5C",X"58",X"DD",X"7E",
		X"04",X"C6",X"10",X"FD",X"77",X"00",X"23",X"7E",X"FD",X"77",X"01",X"FD",X"36",X"02",X"0C",X"23",
		X"DD",X"7E",X"03",X"C6",X"10",X"FD",X"77",X"03",X"3E",X"20",X"CD",X"B2",X"02",X"05",X"C2",X"7B",
		X"27",X"3E",X"FF",X"CD",X"B2",X"02",X"3E",X"FF",X"CD",X"B2",X"02",X"C9",X"31",X"30",X"39",X"38",
		X"33",X"32",X"3B",X"3A",X"35",X"34",X"3D",X"3C",X"37",X"36",X"3F",X"3E",X"09",X"09",X"09",X"09",
		X"00",X"21",X"40",X"58",X"06",X"08",X"23",X"36",X"09",X"23",X"23",X"23",X"05",X"C2",X"16",X"28",
		X"C9",X"00",X"21",X"00",X"50",X"06",X"20",X"11",X"03",X"00",X"0E",X"1C",X"19",X"36",X"24",X"23",
		X"0D",X"C2",X"2D",X"28",X"23",X"05",X"C2",X"2A",X"28",X"C9",X"00",X"4F",X"DD",X"21",X"40",X"58",
		X"07",X"07",X"E6",X"1C",X"5F",X"16",X"00",X"DD",X"19",X"CD",X"50",X"29",X"FD",X"36",X"00",X"00",
		X"FD",X"7E",X"04",X"DD",X"77",X"00",X"FD",X"7E",X"03",X"DD",X"77",X"03",X"DD",X"36",X"02",X"0C",
		X"DD",X"36",X"01",X"1C",X"06",X"03",X"3E",X"08",X"CD",X"B2",X"02",X"DD",X"34",X"01",X"05",X"C2",
		X"66",X"28",X"3E",X"08",X"CD",X"B2",X"02",X"DD",X"36",X"01",X"09",X"3A",X"3C",X"42",X"3D",X"32",
		X"3C",X"42",X"3A",X"3A",X"42",X"FE",X"04",X"C0",X"21",X"40",X"58",X"06",X"08",X"23",X"36",X"09",
		X"23",X"23",X"23",X"05",X"C2",X"8D",X"28",X"06",X"08",X"DD",X"21",X"82",X"41",X"11",X"14",X"00",
		X"DD",X"7E",X"00",X"B7",X"CA",X"B4",X"28",X"DD",X"7E",X"13",X"B7",X"C2",X"B4",X"28",X"79",X"2F",
		X"DD",X"77",X"13",X"C9",X"DD",X"19",X"05",X"C2",X"A0",X"28",X"C9",X"00",X"DD",X"21",X"40",X"58",
		X"FE",X"04",X"DA",X"C9",X"28",X"DD",X"21",X"50",X"58",X"CD",X"50",X"29",X"DD",X"36",X"02",X"0C",
		X"DD",X"36",X"06",X"0C",X"DD",X"36",X"0A",X"0C",X"DD",X"36",X"0E",X"0C",X"FD",X"36",X"00",X"00",
		X"06",X"08",X"3E",X"08",X"90",X"C6",X"20",X"DD",X"77",X"01",X"F6",X"40",X"DD",X"77",X"05",X"E6",
		X"3F",X"F6",X"80",X"DD",X"77",X"09",X"F6",X"C0",X"DD",X"77",X"0D",X"3E",X"08",X"90",X"4F",X"FD",
		X"7E",X"04",X"C6",X"08",X"81",X"DD",X"77",X"00",X"DD",X"77",X"04",X"FD",X"7E",X"04",X"D6",X"08",
		X"91",X"DD",X"77",X"08",X"DD",X"77",X"0C",X"FD",X"7E",X"03",X"C6",X"08",X"81",X"DD",X"77",X"07",
		X"DD",X"77",X"0F",X"91",X"FD",X"7E",X"03",X"D6",X"08",X"DD",X"77",X"03",X"DD",X"77",X"0B",X"3E",
		X"08",X"CD",X"B2",X"02",X"05",X"C2",X"E2",X"28",X"DD",X"36",X"01",X"09",X"DD",X"36",X"05",X"09",
		X"DD",X"36",X"09",X"09",X"DD",X"36",X"0D",X"09",X"3A",X"3C",X"42",X"3D",X"32",X"3C",X"42",X"C9",
		X"00",X"E5",X"C5",X"06",X"20",X"21",X"60",X"58",X"36",X"00",X"23",X"05",X"C2",X"58",X"29",X"C1",
		X"E1",X"C9",X"E6",X"40",X"28",X"03",X"3E",X"FF",X"C9",X"3A",X"39",X"BC",X"A7",X"C8",X"97",X"37",
		X"3E",X"FF",X"CD",X"B2",X"02",X"3E",X"FF",X"CD",X"B2",X"02",X"3E",X"FF",X"CD",X"B2",X"02",X"00",
		X"3E",X"FF",X"CD",X"B2",X"02",X"3E",X"FF",X"CD",X"B2",X"02",X"C3",X"A4",X"25",X"39",X"BC",X"A7",
		X"20",X"06",X"CD",X"9C",X"BB",X"28",X"04",X"C9",X"2A",X"3A",X"BC",X"3E",X"FF",X"32",X"39",X"BC",
		X"7E",X"F5",X"23",X"22",X"3A",X"BC",X"7E",X"D6",X"FF",X"20",X"03",X"32",X"39",X"BC",X"F1",X"C9",
		X"CD",X"5D",X"BB",X"FE",X"02",X"C0",X"32",X"3C",X"BC",X"32",X"3D",X"BC",X"CD",X"29",X"BC",X"20",
		X"16",X"3E",X"0D",X"32",X"3F",X"BC",X"CD",X"24",X"BC",X"32",X"3E",X"BC",X"3E",X"02",X"20",X"02",
		X"A7",X"C9",X"CD",X"49",X"BC",X"18",X"0F",X"FE",X"02",X"C0",X"CD",X"5D",X"BB",X"32",X"3E",X"BC",
		X"CD",X"5D",X"BB",X"32",X"3F",X"BC",X"21",X"40",X"1F",X"2D",X"20",X"FD",X"25",X"20",X"FA",X"21",
		X"3C",X"BC",X"3A",X"9D",X"BC",X"A7",X"C8",X"3A",X"3E",X"BC",X"47",X"21",X"03",X"BC",X"11",X"0C",
		X"00",X"DD",X"21",X"98",X"40",X"FD",X"21",X"42",X"40",X"26",X"05",X"2E",X"00",X"DD",X"7E",X"00",
		X"FD",X"96",X"00",X"DA",X"34",X"2A",X"C2",X"40",X"2A",X"DD",X"7E",X"01",X"FD",X"96",X"01",X"DA",
		X"34",X"2A",X"C2",X"40",X"2A",X"DD",X"7E",X"02",X"FD",X"96",X"02",X"DA",X"34",X"2A",X"CA",X"34",
		X"2A",X"C3",X"40",X"2A",X"FD",X"23",X"FD",X"23",X"FD",X"23",X"2C",X"25",X"C2",X"0D",X"2A",X"C9",
		X"7D",X"32",X"EE",X"40",X"CD",X"DE",X"2A",X"C9",X"00",X"F5",X"C5",X"D5",X"E5",X"D5",X"DD",X"E1",
		X"DD",X"7E",X"01",X"87",X"06",X"00",X"4F",X"FD",X"21",X"00",X"58",X"FD",X"09",X"DD",X"56",X"02",
		X"3E",X"1C",X"92",X"87",X"87",X"87",X"FD",X"77",X"00",X"DD",X"7E",X"00",X"FD",X"77",X"01",X"DD",
		X"46",X"02",X"3E",X"1B",X"90",X"B7",X"CA",X"84",X"2A",X"21",X"40",X"50",X"01",X"20",X"00",X"09",
		X"3D",X"C2",X"7F",X"2A",X"DD",X"4E",X"01",X"06",X"00",X"09",X"11",X"E0",X"FF",X"DD",X"23",X"DD",
		X"23",X"DD",X"23",X"DD",X"7E",X"00",X"FE",X"FF",X"CA",X"B0",X"2A",X"77",X"19",X"06",X"08",X"FD",
		X"35",X"00",X"3E",X"03",X"CD",X"B2",X"02",X"05",X"C2",X"9F",X"2A",X"DD",X"23",X"C3",X"93",X"2A",
		X"FD",X"35",X"00",X"CA",X"BE",X"2A",X"3E",X"03",X"CD",X"B2",X"02",X"C3",X"B0",X"2A",X"E1",X"D1",
		X"C1",X"F1",X"C9",X"00",X"C5",X"D5",X"E5",X"21",X"00",X"50",X"5F",X"16",X"00",X"19",X"11",X"20",
		X"00",X"06",X"20",X"36",X"24",X"19",X"05",X"C2",X"D3",X"2A",X"E1",X"D1",X"C1",X"C9",X"00",X"CD",
		X"6F",X"2D",X"CD",X"99",X"2E",X"3E",X"60",X"32",X"30",X"42",X"3E",X"10",X"32",X"31",X"42",X"11",
		X"52",X"2D",X"CD",X"80",X"09",X"11",X"5E",X"2D",X"CD",X"80",X"09",X"11",X"63",X"2D",X"CD",X"DD",
		X"09",X"11",X"69",X"2D",X"CD",X"DD",X"09",X"AF",X"32",X"EB",X"40",X"AF",X"32",X"EC",X"40",X"3A",
		X"40",X"40",X"B7",X"C2",X"1C",X"2B",X"3A",X"00",X"60",X"C3",X"1F",X"2B",X"3A",X"00",X"68",X"32",
		X"2E",X"42",X"E6",X"04",X"C2",X"3A",X"2B",X"3A",X"2E",X"42",X"E6",X"08",X"C2",X"48",X"2B",X"3A",
		X"2E",X"42",X"E6",X"10",X"C2",X"C3",X"2B",X"C3",X"57",X"2B",X"3A",X"EB",X"40",X"B7",X"CA",X"40",
		X"2C",X"3D",X"32",X"EB",X"40",X"C3",X"57",X"2B",X"3A",X"EB",X"40",X"FE",X"1C",X"CA",X"40",X"2C",
		X"3C",X"32",X"EB",X"40",X"C3",X"57",X"2B",X"DD",X"21",X"40",X"58",X"21",X"89",X"2B",X"3A",X"EB",
		X"40",X"07",X"E6",X"FE",X"5F",X"16",X"00",X"19",X"7E",X"DD",X"77",X"00",X"23",X"7E",X"DD",X"77",
		X"03",X"DD",X"36",X"01",X"20",X"DD",X"36",X"02",X"02",X"3A",X"40",X"40",X"B7",X"CA",X"40",X"2C",
		X"DD",X"35",X"00",X"DD",X"35",X"00",X"C3",X"40",X"2C",X"35",X"9C",X"45",X"9C",X"55",X"9C",X"65",
		X"9C",X"75",X"9C",X"85",X"9C",X"95",X"9C",X"A5",X"9C",X"B5",X"9C",X"35",X"AC",X"45",X"AC",X"55",
		X"AC",X"65",X"AC",X"75",X"AC",X"85",X"AC",X"95",X"AC",X"A5",X"AC",X"B5",X"AC",X"C9",X"AC",X"35",
		X"BC",X"45",X"BC",X"55",X"BC",X"65",X"BC",X"75",X"BC",X"85",X"BC",X"95",X"BC",X"A5",X"BC",X"B5",
		X"BC",X"C7",X"BC",X"3A",X"EB",X"40",X"FE",X"1C",X"CA",X"84",X"2C",X"FE",X"12",X"CA",X"06",X"2C",
		X"FE",X"12",X"DA",X"DF",X"2B",X"FE",X"1B",X"CA",X"E4",X"2B",X"C6",X"09",X"C3",X"E6",X"2B",X"C6",
		X"0A",X"C3",X"E6",X"2B",X"3E",X"2C",X"32",X"ED",X"40",X"3A",X"EC",X"40",X"FE",X"0B",X"D2",X"40",
		X"2C",X"21",X"E0",X"40",X"5F",X"16",X"00",X"19",X"3A",X"ED",X"40",X"77",X"3A",X"EC",X"40",X"3C",
		X"32",X"EC",X"40",X"C3",X"21",X"2C",X"3E",X"24",X"32",X"ED",X"40",X"3A",X"EC",X"40",X"B7",X"CA",
		X"40",X"2C",X"3D",X"32",X"EC",X"40",X"21",X"E0",X"40",X"5F",X"16",X"00",X"19",X"3A",X"ED",X"40",
		X"77",X"DD",X"21",X"DD",X"40",X"DD",X"36",X"00",X"06",X"DD",X"36",X"01",X"12",X"DD",X"36",X"02",
		X"0B",X"DD",X"36",X"0D",X"FF",X"11",X"DD",X"40",X"CD",X"80",X"09",X"3E",X"50",X"CD",X"B2",X"02",
		X"3E",X"30",X"CD",X"B2",X"02",X"21",X"31",X"42",X"7E",X"D6",X"01",X"27",X"77",X"C2",X"58",X"2C",
		X"36",X"10",X"2B",X"7E",X"D6",X"01",X"27",X"77",X"21",X"30",X"42",X"7E",X"FE",X"00",X"C2",X"75",
		X"2C",X"23",X"7E",X"FE",X"01",X"C2",X"75",X"2C",X"AF",X"32",X"31",X"42",X"11",X"69",X"2D",X"CD",
		X"DD",X"09",X"C3",X"84",X"2C",X"11",X"63",X"2D",X"CD",X"DD",X"09",X"11",X"69",X"2D",X"CD",X"DD",
		X"09",X"C3",X"0F",X"2B",X"3A",X"EE",X"40",X"47",X"3E",X"04",X"90",X"47",X"B7",X"CA",X"DE",X"2C",
		X"DD",X"21",X"4B",X"40",X"FD",X"21",X"4E",X"40",X"11",X"FA",X"FF",X"0E",X"03",X"DD",X"7E",X"00",
		X"FD",X"77",X"00",X"DD",X"23",X"FD",X"23",X"0D",X"C2",X"9D",X"2C",X"DD",X"19",X"FD",X"19",X"05",
		X"C2",X"9B",X"2C",X"3A",X"EE",X"40",X"47",X"3E",X"04",X"90",X"47",X"DD",X"21",X"7E",X"40",X"FD",
		X"21",X"8C",X"40",X"0E",X"0A",X"DD",X"7E",X"00",X"FD",X"77",X"00",X"DD",X"23",X"FD",X"23",X"0D",
		X"C2",X"C5",X"2C",X"11",X"E8",X"FF",X"DD",X"19",X"FD",X"19",X"05",X"C2",X"C3",X"2C",X"3A",X"EE",
		X"40",X"47",X"4F",X"FD",X"21",X"42",X"40",X"B7",X"CA",X"F5",X"2C",X"FD",X"23",X"FD",X"23",X"FD",
		X"23",X"05",X"C2",X"EB",X"2C",X"DD",X"21",X"98",X"40",X"06",X"03",X"DD",X"7E",X"00",X"FD",X"77",
		X"00",X"DD",X"23",X"FD",X"23",X"05",X"C2",X"FB",X"2C",X"FD",X"21",X"54",X"40",X"79",X"B7",X"CA",
		X"1B",X"2D",X"11",X"0E",X"00",X"FD",X"19",X"0D",X"C2",X"15",X"2D",X"DD",X"21",X"E0",X"40",X"0E",
		X"0A",X"DD",X"7E",X"00",X"FD",X"77",X"00",X"DD",X"23",X"FD",X"23",X"0D",X"C2",X"21",X"2D",X"CD",
		X"6F",X"2D",X"AF",X"32",X"40",X"58",X"3E",X"FF",X"CD",X"B2",X"02",X"3E",X"FF",X"CD",X"B2",X"02",
		X"3E",X"FF",X"CD",X"B2",X"02",X"06",X"1C",X"3E",X"02",X"CD",X"C3",X"2A",X"3C",X"05",X"C2",X"49",
		X"2D",X"C9",X"02",X"1A",X"07",X"1B",X"0E",X"10",X"24",X"1D",X"12",X"16",X"0E",X"FF",X"07",X"1C",
		X"0C",X"2D",X"FF",X"07",X"1C",X"0A",X"30",X"42",X"02",X"07",X"1C",X"0D",X"31",X"42",X"01",X"00",
		X"3E",X"02",X"06",X"18",X"CD",X"C3",X"2A",X"3C",X"05",X"C2",X"74",X"2D",X"11",X"41",X"2E",X"CD",
		X"80",X"09",X"11",X"53",X"2E",X"CD",X"80",X"09",X"11",X"7B",X"2E",X"CD",X"DD",X"09",X"DD",X"21",
		X"51",X"40",X"DD",X"36",X"00",X"00",X"DD",X"36",X"01",X"05",X"DD",X"36",X"02",X"11",X"DD",X"36",
		X"0D",X"FF",X"11",X"51",X"40",X"CD",X"80",X"09",X"11",X"5B",X"2E",X"CD",X"80",X"09",X"11",X"81",
		X"2E",X"CD",X"DD",X"09",X"DD",X"21",X"5F",X"40",X"DD",X"36",X"00",X"01",X"DD",X"36",X"01",X"07",
		X"DD",X"36",X"02",X"11",X"DD",X"36",X"0D",X"FF",X"11",X"5F",X"40",X"CD",X"80",X"09",X"11",X"63",
		X"2E",X"CD",X"80",X"09",X"11",X"87",X"2E",X"CD",X"DD",X"09",X"DD",X"21",X"6D",X"40",X"DD",X"36",
		X"00",X"02",X"DD",X"36",X"01",X"09",X"DD",X"36",X"02",X"11",X"DD",X"36",X"0D",X"FF",X"11",X"6D",
		X"40",X"CD",X"80",X"09",X"11",X"6B",X"2E",X"CD",X"80",X"09",X"11",X"8D",X"2E",X"CD",X"DD",X"09",
		X"DD",X"21",X"7B",X"40",X"DD",X"36",X"00",X"03",X"DD",X"36",X"01",X"0B",X"DD",X"36",X"02",X"11",
		X"DD",X"36",X"0D",X"FF",X"11",X"7B",X"40",X"CD",X"80",X"09",X"11",X"73",X"2E",X"CD",X"80",X"09",
		X"11",X"93",X"2E",X"CD",X"DD",X"09",X"DD",X"21",X"89",X"40",X"DD",X"36",X"00",X"04",X"DD",X"36",
		X"01",X"0D",X"DD",X"36",X"02",X"11",X"DD",X"36",X"0D",X"FF",X"11",X"89",X"40",X"CD",X"80",X"09",
		X"C9",X"06",X"03",X"0A",X"1C",X"0C",X"18",X"1B",X"0E",X"24",X"24",X"24",X"24",X"24",X"17",X"0A",
		X"16",X"0E",X"FF",X"0C",X"05",X"04",X"17",X"18",X"01",X"2D",X"FF",X"0C",X"07",X"04",X"17",X"18",
		X"02",X"2D",X"FF",X"0C",X"09",X"04",X"17",X"18",X"03",X"2D",X"FF",X"0C",X"0B",X"04",X"17",X"18",
		X"04",X"2D",X"FF",X"0C",X"0D",X"04",X"17",X"18",X"05",X"2D",X"FF",X"0C",X"05",X"09",X"42",X"40",
		X"06",X"0C",X"07",X"09",X"45",X"40",X"06",X"0C",X"09",X"09",X"48",X"40",X"06",X"0C",X"0B",X"09",
		X"4B",X"40",X"06",X"0C",X"0D",X"09",X"4E",X"40",X"06",X"00",X"11",X"D4",X"2E",X"CD",X"80",X"09",
		X"11",X"E9",X"2E",X"CD",X"80",X"09",X"11",X"F2",X"2E",X"CD",X"80",X"09",X"11",X"08",X"2F",X"CD",
		X"80",X"09",X"11",X"20",X"2F",X"CD",X"80",X"09",X"21",X"E0",X"40",X"06",X"0A",X"36",X"24",X"23",
		X"05",X"C2",X"BD",X"2E",X"3E",X"01",X"32",X"00",X"60",X"3E",X"01",X"32",X"01",X"60",X"3E",X"01",
		X"32",X"02",X"60",X"C9",X"05",X"10",X"06",X"17",X"0A",X"16",X"0E",X"24",X"1B",X"0E",X"10",X"12",
		X"1C",X"1D",X"1B",X"0A",X"1D",X"12",X"18",X"17",X"FF",X"06",X"12",X"05",X"17",X"0A",X"16",X"0E",
		X"2D",X"FF",X"07",X"14",X"05",X"0A",X"24",X"0B",X"24",X"0C",X"24",X"0D",X"24",X"0E",X"24",X"0F",
		X"24",X"10",X"24",X"11",X"24",X"12",X"24",X"FF",X"07",X"16",X"05",X"13",X"24",X"14",X"24",X"15",
		X"24",X"16",X"24",X"17",X"24",X"18",X"24",X"19",X"24",X"1A",X"24",X"1B",X"24",X"A3",X"A1",X"FF",
		X"07",X"18",X"05",X"1C",X"24",X"1D",X"24",X"1E",X"24",X"1F",X"24",X"20",X"24",X"21",X"24",X"22",
		X"24",X"23",X"24",X"2C",X"24",X"A2",X"A0",X"FF",X"3A",X"00",X"70",X"47",X"E6",X"08",X"3E",X"00",
		X"28",X"01",X"3C",X"32",X"3C",X"40",X"78",X"E6",X"04",X"3E",X"00",X"00",X"00",X"3C",X"32",X"36",
		X"40",X"78",X"E6",X"01",X"3E",X"03",X"20",X"02",X"3C",X"3C",X"32",X"3D",X"40",X"3A",X"00",X"68",
		X"47",X"E6",X"40",X"3E",X"01",X"20",X"01",X"3C",X"32",X"38",X"40",X"78",X"E6",X"80",X"3E",X"03",
		X"20",X"02",X"3C",X"3C",X"32",X"3A",X"40",X"3E",X"01",X"00",X"00",X"00",X"32",X"06",X"70",X"32",
		X"07",X"70",X"18",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"21",X"54",
		X"40",X"06",X"05",X"0E",X"0A",X"DD",X"21",X"D3",X"2F",X"3A",X"36",X"40",X"B7",X"CA",X"A4",X"2F",
		X"DD",X"21",X"DD",X"2F",X"DD",X"7E",X"00",X"77",X"23",X"DD",X"23",X"0D",X"C2",X"A4",X"2F",X"23",
		X"23",X"23",X"23",X"05",X"C2",X"93",X"2F",X"21",X"42",X"40",X"06",X"05",X"36",X"00",X"23",X"36",
		X"50",X"23",X"36",X"00",X"23",X"05",X"C2",X"BC",X"2F",X"3A",X"3A",X"40",X"FE",X"04",X"C0",X"32",
		X"32",X"40",X"C9",X"3F",X"3D",X"3B",X"39",X"37",X"35",X"33",X"31",X"2F",X"24",X"3E",X"3C",X"3A",
		X"38",X"36",X"34",X"32",X"30",X"24",X"24",X"00",X"00",X"0E",X"23",X"CD",X"C8",X"B4",X"EB",X"CD",
		X"B6",X"A4",X"D1",X"E1",X"01",X"80",X"00",X"09",X"EB",X"B7",X"28",X"B0",X"11",X"80",X"00",X"73",
		X"00",X"CD",X"FE",X"32",X"3A",X"3B",X"42",X"FE",X"03",X"C2",X"20",X"30",X"3A",X"27",X"42",X"E6",
		X"03",X"C2",X"2B",X"30",X"CD",X"7E",X"30",X"CD",X"EB",X"30",X"CD",X"50",X"31",X"C3",X"2B",X"30",
		X"FE",X"04",X"DA",X"28",X"30",X"CD",X"42",X"30",X"CD",X"50",X"31",X"CD",X"6A",X"33",X"CD",X"D1",
		X"36",X"3A",X"3B",X"42",X"FE",X"04",X"DA",X"3F",X"30",X"CD",X"E7",X"31",X"CD",X"F7",X"33",X"CD",
		X"10",X"03",X"00",X"3A",X"2E",X"42",X"E6",X"04",X"C2",X"58",X"30",X"3A",X"2E",X"42",X"E6",X"08",
		X"C2",X"6B",X"30",X"AF",X"32",X"28",X"42",X"C9",X"3A",X"2D",X"42",X"B7",X"C2",X"65",X"30",X"3E",
		X"FE",X"32",X"28",X"42",X"C9",X"3E",X"FF",X"32",X"28",X"42",X"C9",X"3A",X"2D",X"42",X"B7",X"C2",
		X"78",X"30",X"3E",X"02",X"32",X"28",X"42",X"C9",X"3E",X"01",X"32",X"28",X"42",X"C9",X"00",X"3A",
		X"26",X"42",X"FE",X"02",X"D8",X"AF",X"32",X"28",X"42",X"3A",X"2E",X"42",X"E6",X"04",X"CA",X"A1",
		X"30",X"3A",X"22",X"42",X"FE",X"C0",X"CA",X"B6",X"30",X"C6",X"01",X"32",X"22",X"42",X"C3",X"B6",
		X"30",X"3A",X"2E",X"42",X"E6",X"08",X"CA",X"B6",X"30",X"3A",X"22",X"42",X"FE",X"40",X"CA",X"B6",
		X"30",X"D6",X"01",X"32",X"22",X"42",X"3A",X"24",X"42",X"A7",X"CA",X"C2",X"30",X"3D",X"32",X"24",
		X"42",X"C9",X"3A",X"22",X"42",X"A7",X"F2",X"CB",X"30",X"2F",X"3C",X"D6",X"40",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"E6",X"07",X"32",X"24",X"42",X"3A",X"22",X"42",X"E6",X"80",X"CA",X"E5",X"30",X"3E",
		X"FF",X"32",X"28",X"42",X"C9",X"3E",X"01",X"32",X"28",X"42",X"C9",X"00",X"3A",X"26",X"42",X"FE",
		X"02",X"D8",X"AF",X"32",X"29",X"42",X"3A",X"2E",X"42",X"E6",X"10",X"CA",X"0E",X"31",X"3A",X"23",
		X"42",X"FE",X"C0",X"CA",X"1B",X"31",X"C6",X"01",X"32",X"23",X"42",X"C3",X"1B",X"31",X"3A",X"23",
		X"42",X"FE",X"40",X"CA",X"1B",X"31",X"D6",X"01",X"32",X"23",X"42",X"3A",X"25",X"42",X"A7",X"CA",
		X"27",X"31",X"3D",X"32",X"25",X"42",X"C9",X"3A",X"23",X"42",X"A7",X"F2",X"30",X"31",X"2F",X"3C",
		X"D6",X"40",X"0F",X"0F",X"0F",X"0F",X"0F",X"E6",X"07",X"32",X"25",X"42",X"3A",X"23",X"42",X"E6",
		X"80",X"CA",X"4A",X"31",X"3E",X"FF",X"32",X"29",X"42",X"C9",X"3E",X"01",X"32",X"29",X"42",X"C9",
		X"00",X"06",X"03",X"0E",X"01",X"11",X"FB",X"FF",X"DD",X"21",X"4A",X"41",X"DD",X"7E",X"00",X"FE",
		X"01",X"CA",X"6C",X"31",X"FE",X"02",X"CA",X"D1",X"31",X"C3",X"DF",X"31",X"3A",X"28",X"42",X"FE",
		X"02",X"CA",X"91",X"31",X"FE",X"01",X"CA",X"91",X"31",X"FE",X"FE",X"CA",X"86",X"31",X"FE",X"FF",
		X"CA",X"86",X"31",X"C3",X"A2",X"31",X"3A",X"2B",X"42",X"FE",X"20",X"D2",X"99",X"31",X"C3",X"A2",
		X"31",X"3A",X"2B",X"42",X"FE",X"D8",X"D2",X"A2",X"31",X"3A",X"28",X"42",X"DD",X"86",X"04",X"DD",
		X"77",X"04",X"3A",X"29",X"42",X"FE",X"01",X"CA",X"B2",X"31",X"FE",X"FF",X"CA",X"BD",X"31",X"C3",
		X"DB",X"31",X"3A",X"2C",X"42",X"FE",X"F0",X"DA",X"C5",X"31",X"C3",X"DB",X"31",X"3A",X"2C",X"42",
		X"FE",X"30",X"DA",X"DB",X"31",X"3A",X"29",X"42",X"DD",X"86",X"03",X"DD",X"77",X"03",X"C3",X"DB",
		X"31",X"3A",X"2A",X"42",X"DD",X"66",X"03",X"84",X"DD",X"77",X"03",X"78",X"CD",X"87",X"34",X"DD",
		X"19",X"0C",X"05",X"C2",X"5C",X"31",X"C9",X"00",X"3A",X"2E",X"42",X"E6",X"10",X"C2",X"F5",X"31",
		X"AF",X"32",X"34",X"42",X"C9",X"3A",X"34",X"42",X"B7",X"C0",X"3E",X"01",X"32",X"34",X"42",X"3A",
		X"72",X"41",X"B7",X"CA",X"13",X"32",X"FE",X"01",X"CA",X"23",X"32",X"FE",X"02",X"CA",X"33",X"32",
		X"C3",X"44",X"32",X"3A",X"40",X"41",X"FE",X"01",X"C2",X"44",X"32",X"3A",X"59",X"41",X"A7",X"CA",
		X"54",X"32",X"C9",X"3A",X"45",X"41",X"FE",X"01",X"C2",X"44",X"32",X"3A",X"5E",X"41",X"A7",X"CA",
		X"6A",X"32",X"C9",X"3A",X"4A",X"41",X"FE",X"01",X"C2",X"44",X"32",X"3A",X"68",X"41",X"A7",X"CA",
		X"80",X"32",X"C9",X"B3",X"3A",X"72",X"41",X"3C",X"FE",X"03",X"DA",X"4E",X"32",X"AF",X"32",X"72",
		X"41",X"C3",X"FF",X"31",X"3E",X"01",X"32",X"72",X"41",X"3E",X"00",X"CD",X"32",X"09",X"DD",X"21",
		X"59",X"41",X"FD",X"21",X"59",X"41",X"CD",X"96",X"32",X"C9",X"3E",X"02",X"32",X"72",X"41",X"3E",
		X"00",X"CD",X"32",X"09",X"DD",X"21",X"5E",X"41",X"FD",X"21",X"63",X"41",X"CD",X"AD",X"32",X"C9",
		X"3E",X"00",X"32",X"72",X"41",X"3E",X"00",X"CD",X"32",X"09",X"DD",X"21",X"68",X"41",X"FD",X"21",
		X"6D",X"41",X"CD",X"C6",X"32",X"C9",X"00",X"3A",X"43",X"41",X"D6",X"01",X"32",X"35",X"42",X"3A",
		X"44",X"41",X"C6",X"08",X"32",X"36",X"42",X"32",X"37",X"42",X"C3",X"DF",X"32",X"00",X"3A",X"48",
		X"41",X"C6",X"03",X"32",X"35",X"42",X"3A",X"49",X"41",X"C6",X"08",X"32",X"36",X"42",X"C6",X"10",
		X"32",X"37",X"42",X"C3",X"DF",X"32",X"00",X"3A",X"4D",X"41",X"C6",X"04",X"32",X"35",X"42",X"3A",
		X"4E",X"41",X"C6",X"04",X"32",X"36",X"42",X"C6",X"18",X"32",X"37",X"42",X"C3",X"DF",X"32",X"00",
		X"DD",X"36",X"00",X"01",X"FD",X"36",X"00",X"01",X"3A",X"35",X"42",X"DD",X"77",X"03",X"FD",X"77",
		X"03",X"3A",X"36",X"42",X"DD",X"77",X"04",X"3A",X"37",X"42",X"FD",X"77",X"04",X"C9",X"00",X"3A",
		X"35",X"40",X"A7",X"CA",X"1B",X"33",X"3A",X"40",X"40",X"A7",X"C2",X"13",X"33",X"3A",X"00",X"60",
		X"C3",X"16",X"33",X"3A",X"00",X"68",X"00",X"32",X"2E",X"42",X"C9",X"3A",X"26",X"42",X"FE",X"03",
		X"DA",X"2B",X"33",X"3A",X"3B",X"42",X"FE",X"03",X"CA",X"46",X"33",X"3A",X"27",X"42",X"E6",X"0F",
		X"C0",X"3A",X"2F",X"42",X"3C",X"E6",X"0F",X"32",X"2F",X"42",X"4F",X"06",X"00",X"21",X"5A",X"33",
		X"09",X"7E",X"32",X"2E",X"42",X"C9",X"3A",X"2B",X"42",X"D6",X"81",X"DA",X"54",X"33",X"3E",X"04",
		X"32",X"2E",X"42",X"C9",X"3E",X"08",X"32",X"2E",X"42",X"C9",X"14",X"08",X"14",X"04",X"18",X"08",
		X"14",X"08",X"14",X"04",X"18",X"08",X"14",X"04",X"18",X"08",X"00",X"DD",X"21",X"4F",X"41",X"DD",
		X"7E",X"00",X"B7",X"C8",X"3A",X"27",X"42",X"E6",X"03",X"C2",X"95",X"33",X"DD",X"7E",X"01",X"B7",
		X"C2",X"87",X"33",X"DD",X"36",X"01",X"15",X"DD",X"7E",X"01",X"3C",X"FE",X"18",X"C2",X"92",X"33",
		X"3E",X"15",X"DD",X"77",X"01",X"FD",X"21",X"40",X"41",X"FD",X"7E",X"00",X"B7",X"CA",X"B3",X"33",
		X"FE",X"03",X"CA",X"B3",X"33",X"FD",X"7E",X"04",X"DD",X"77",X"04",X"FD",X"7E",X"03",X"C6",X"10",
		X"DD",X"77",X"03",X"FD",X"21",X"45",X"41",X"FD",X"7E",X"00",X"B7",X"CA",X"D3",X"33",X"FE",X"03",
		X"CA",X"D3",X"33",X"FD",X"7E",X"04",X"C6",X"08",X"DD",X"77",X"04",X"FD",X"7E",X"03",X"C6",X"10",
		X"DD",X"77",X"03",X"FD",X"21",X"4A",X"41",X"FD",X"7E",X"00",X"B7",X"CA",X"F3",X"33",X"FE",X"03",
		X"CA",X"F3",X"33",X"FD",X"7E",X"04",X"C6",X"08",X"DD",X"77",X"04",X"FD",X"7E",X"03",X"C6",X"10",
		X"DD",X"77",X"03",X"CD",X"DE",X"35",X"C9",X"00",X"26",X"05",X"2E",X"01",X"DD",X"21",X"59",X"41",
		X"DD",X"7E",X"00",X"B7",X"CA",X"20",X"34",X"DD",X"7E",X"03",X"D6",X"04",X"DD",X"77",X"03",X"FE",
		X"04",X"D2",X"1C",X"34",X"DD",X"36",X"00",X"00",X"DD",X"36",X"04",X"00",X"7D",X"CD",X"2B",X"34",
		X"11",X"05",X"00",X"DD",X"19",X"2C",X"25",X"C2",X"00",X"34",X"C9",X"00",X"3D",X"47",X"DD",X"21",
		X"59",X"41",X"B7",X"CA",X"3F",X"34",X"11",X"05",X"00",X"DD",X"19",X"3D",X"C2",X"39",X"34",X"78",
		X"FD",X"21",X"60",X"58",X"07",X"07",X"E6",X"FC",X"5F",X"16",X"00",X"FD",X"19",X"DD",X"7E",X"04",
		X"FD",X"77",X"01",X"3A",X"3C",X"40",X"B7",X"CA",X"6B",X"34",X"3A",X"40",X"40",X"B7",X"CA",X"6B",
		X"34",X"DD",X"7E",X"03",X"2F",X"FD",X"77",X"03",X"C3",X"71",X"34",X"DD",X"7E",X"03",X"FD",X"77",
		X"03",X"DD",X"7E",X"04",X"B7",X"C2",X"7C",X"34",X"DD",X"36",X"00",X"00",X"FD",X"7E",X"03",X"FE",
		X"F8",X"D8",X"DD",X"36",X"04",X"00",X"C9",X"00",X"F5",X"3A",X"4D",X"42",X"B7",X"CA",X"41",X"35",
		X"FE",X"FF",X"CA",X"2D",X"35",X"F1",X"3D",X"CA",X"A2",X"34",X"3D",X"CA",X"BF",X"34",X"3D",X"CA",
		X"F6",X"34",X"DD",X"21",X"40",X"41",X"FD",X"21",X"40",X"58",X"DD",X"7E",X"04",X"FD",X"77",X"00",
		X"FD",X"36",X"01",X"10",X"FD",X"36",X"02",X"03",X"DD",X"7E",X"03",X"FD",X"77",X"03",X"C9",X"DD",
		X"21",X"45",X"41",X"FD",X"21",X"44",X"58",X"DD",X"7E",X"04",X"FD",X"77",X"00",X"FD",X"36",X"01",
		X"12",X"FD",X"36",X"02",X"04",X"DD",X"7E",X"03",X"FD",X"77",X"03",X"FD",X"21",X"48",X"58",X"DD",
		X"7E",X"04",X"C6",X"10",X"FD",X"77",X"00",X"FD",X"36",X"01",X"11",X"FD",X"36",X"02",X"04",X"DD",
		X"7E",X"03",X"FD",X"77",X"03",X"C9",X"DD",X"21",X"4A",X"41",X"FD",X"21",X"4C",X"58",X"DD",X"7E",
		X"04",X"FD",X"77",X"00",X"FD",X"36",X"01",X"14",X"FD",X"36",X"02",X"05",X"DD",X"7E",X"03",X"FD",
		X"77",X"03",X"FD",X"21",X"50",X"58",X"DD",X"7E",X"04",X"C6",X"10",X"FD",X"77",X"00",X"FD",X"36",
		X"01",X"13",X"FD",X"36",X"02",X"05",X"DD",X"7E",X"03",X"FD",X"77",X"03",X"C9",X"F1",X"C5",X"D5",
		X"E5",X"DD",X"E5",X"FD",X"E5",X"3D",X"CA",X"98",X"35",X"3D",X"CA",X"A6",X"35",X"3D",X"CA",X"B4",
		X"35",X"C5",X"D5",X"E5",X"DD",X"E5",X"FD",X"E5",X"3A",X"45",X"41",X"FE",X"01",X"C2",X"5E",X"35",
		X"DD",X"21",X"45",X"41",X"21",X"CC",X"35",X"06",X"02",X"0E",X"04",X"CD",X"4A",X"36",X"3A",X"40",
		X"41",X"FE",X"01",X"C2",X"74",X"35",X"DD",X"21",X"40",X"41",X"21",X"C7",X"35",X"06",X"02",X"0E",
		X"02",X"CD",X"4A",X"36",X"3A",X"4A",X"41",X"FE",X"01",X"C2",X"8A",X"35",X"DD",X"21",X"4A",X"41",
		X"21",X"D5",X"35",X"06",X"02",X"0E",X"04",X"CD",X"4A",X"36",X"3E",X"FF",X"32",X"4D",X"42",X"FD",
		X"E1",X"DD",X"E1",X"E1",X"D1",X"C1",X"F1",X"C9",X"DD",X"21",X"40",X"41",X"06",X"01",X"0E",X"02",
		X"CD",X"9D",X"36",X"C3",X"BF",X"35",X"DD",X"21",X"45",X"41",X"06",X"01",X"0E",X"04",X"CD",X"9D",
		X"36",X"C3",X"BF",X"35",X"DD",X"21",X"4A",X"41",X"06",X"02",X"0E",X"04",X"CD",X"9D",X"36",X"FD",
		X"E1",X"DD",X"E1",X"E1",X"D1",X"C1",X"C9",X"03",X"42",X"40",X"43",X"41",X"04",X"4A",X"48",X"46",
		X"44",X"4B",X"49",X"47",X"45",X"05",X"52",X"50",X"4E",X"4C",X"53",X"51",X"4F",X"4D",X"00",X"3A",
		X"4F",X"41",X"B7",X"C8",X"3A",X"4D",X"42",X"FE",X"01",X"C2",X"0B",X"36",X"DD",X"21",X"4F",X"41",
		X"FD",X"21",X"54",X"58",X"DD",X"7E",X"04",X"FD",X"77",X"00",X"DD",X"7E",X"01",X"FD",X"77",X"01",
		X"FD",X"36",X"02",X"06",X"DD",X"7E",X"03",X"FD",X"77",X"03",X"C9",X"3A",X"50",X"41",X"FE",X"15",
		X"CA",X"1D",X"36",X"FE",X"16",X"CA",X"23",X"36",X"FE",X"17",X"CA",X"29",X"36",X"21",X"3B",X"36",
		X"C3",X"2F",X"36",X"21",X"40",X"36",X"C3",X"2F",X"36",X"21",X"45",X"36",X"C3",X"2F",X"36",X"DD",
		X"21",X"4F",X"41",X"06",X"02",X"0E",X"02",X"CD",X"4A",X"36",X"C9",X"06",X"56",X"54",X"57",X"55",
		X"06",X"5A",X"58",X"5B",X"59",X"06",X"5E",X"5C",X"5F",X"5D",X"00",X"DD",X"7E",X"03",X"0F",X"0F",
		X"E6",X"3E",X"5F",X"16",X"00",X"FD",X"21",X"00",X"58",X"FD",X"19",X"DD",X"7E",X"04",X"2F",X"57",
		X"7B",X"0F",X"E6",X"1F",X"5F",X"C5",X"7A",X"2F",X"C6",X"00",X"FD",X"77",X"00",X"7E",X"FD",X"77",
		X"01",X"FD",X"23",X"FD",X"23",X"05",X"C2",X"66",X"36",X"C1",X"FD",X"21",X"E0",X"53",X"16",X"00",
		X"FD",X"19",X"11",X"E0",X"FF",X"FD",X"E5",X"C5",X"23",X"7E",X"FD",X"77",X"00",X"FD",X"19",X"0D",
		X"C2",X"88",X"36",X"C1",X"FD",X"E1",X"FD",X"23",X"05",X"C2",X"85",X"36",X"C9",X"00",X"78",X"FE",
		X"01",X"C2",X"AC",X"36",X"DD",X"7E",X"03",X"C6",X"08",X"C3",X"AF",X"36",X"DD",X"7E",X"03",X"0F",
		X"0F",X"E6",X"3E",X"5F",X"16",X"00",X"FD",X"21",X"00",X"58",X"FD",X"19",X"DD",X"7E",X"04",X"2F",
		X"57",X"7A",X"2F",X"C6",X"00",X"FD",X"77",X"00",X"FD",X"23",X"FD",X"23",X"05",X"C2",X"C1",X"36",
		X"C9",X"00",X"3A",X"3B",X"42",X"FE",X"03",X"C0",X"DD",X"21",X"54",X"41",X"DD",X"7E",X"01",X"B7",
		X"C2",X"E7",X"36",X"DD",X"36",X"01",X"15",X"3A",X"27",X"42",X"E6",X"03",X"C2",X"FD",X"36",X"DD",
		X"7E",X"01",X"3C",X"FE",X"18",X"C2",X"FA",X"36",X"3E",X"15",X"DD",X"77",X"01",X"FD",X"21",X"40",
		X"41",X"FD",X"7E",X"00",X"FE",X"01",X"C2",X"17",X"37",X"FD",X"7E",X"04",X"DD",X"77",X"04",X"FD",
		X"7E",X"03",X"C6",X"10",X"DD",X"77",X"03",X"FD",X"21",X"45",X"41",X"FD",X"7E",X"00",X"FE",X"01",
		X"C2",X"33",X"37",X"FD",X"7E",X"04",X"C6",X"08",X"DD",X"77",X"04",X"FD",X"7E",X"03",X"C6",X"10",
		X"DD",X"77",X"03",X"FD",X"21",X"4A",X"41",X"FD",X"7E",X"00",X"FE",X"01",X"C2",X"4F",X"37",X"FD",
		X"7E",X"04",X"C6",X"08",X"DD",X"77",X"04",X"FD",X"7E",X"03",X"C6",X"10",X"DD",X"77",X"03",X"CD",
		X"53",X"37",X"C9",X"00",X"DD",X"21",X"54",X"41",X"FD",X"21",X"58",X"58",X"FD",X"36",X"01",X"15",
		X"DD",X"7E",X"04",X"FD",X"77",X"00",X"3A",X"2E",X"42",X"E6",X"10",X"C2",X"75",X"37",X"FD",X"36",
		X"01",X"09",X"C3",X"7E",X"37",X"DD",X"7E",X"01",X"FD",X"77",X"01",X"C3",X"7E",X"37",X"FD",X"36",
		X"02",X"0C",X"DD",X"7E",X"03",X"FD",X"77",X"03",X"C9",X"0D",X"0A",X"52",X"65",X"61",X"64",X"2D",
		X"61",X"66",X"74",X"65",X"72",X"2D",X"77",X"72",X"69",X"74",X"65",X"00",X"0D",X"0A",X"4C",X"6F",
		X"67",X"69",X"63",X"61",X"6C",X"20",X"64",X"69",X"73",X"6B",X"20",X"65",X"72",X"72",X"6F",X"72",
		X"20",X"80",X"00",X"00",X"68",X"2C",X"20",X"64",X"72",X"69",X"76",X"65",X"20",X"00",X"2C",X"20",
		X"62",X"6C",X"6F",X"63",X"6B",X"20",X"80",X"00",X"00",X"81",X"00",X"00",X"68",X"0D",X"0A",X"00",
		X"20",X"65",X"72",X"72",X"6F",X"72",X"3A",X"20",X"44",X"72",X"69",X"76",X"65",X"20",X"00",X"00",
		X"0D",X"0A",X"44",X"72",X"69",X"76",X"65",X"20",X"00",X"20",X"6E",X"6F",X"74",X"20",X"72",X"65",
		X"61",X"64",X"79",X"0D",X"0A",X"00",X"0D",X"0A",X"44",X"69",X"73",X"6B",X"65",X"74",X"74",X"65",
		X"00",X"CD",X"27",X"38",X"3A",X"3B",X"42",X"FE",X"04",X"DA",X"24",X"38",X"3A",X"3C",X"42",X"B7",
		X"C2",X"24",X"38",X"3A",X"9B",X"40",X"3C",X"32",X"9B",X"40",X"AF",X"32",X"26",X"42",X"32",X"27",
		X"42",X"CD",X"96",X"39",X"CD",X"10",X"03",X"00",X"CD",X"61",X"3D",X"3A",X"2D",X"42",X"B7",X"CA",
		X"36",X"38",X"3D",X"32",X"2D",X"42",X"00",X"3A",X"26",X"42",X"21",X"27",X"42",X"B6",X"C2",X"9A",
		X"38",X"21",X"FE",X"38",X"3A",X"35",X"40",X"B7",X"C2",X"4E",X"38",X"21",X"1A",X"39",X"3A",X"9B",
		X"40",X"E6",X"0F",X"3D",X"07",X"E6",X"FE",X"4F",X"06",X"00",X"09",X"7E",X"32",X"3B",X"42",X"D6",
		X"04",X"32",X"3A",X"42",X"23",X"7E",X"32",X"3F",X"42",X"32",X"40",X"42",X"AF",X"32",X"3E",X"42",
		X"3A",X"9B",X"40",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"C6",X"01",X"32",X"3D",X"42",X"21",X"2E",
		X"39",X"3A",X"3A",X"42",X"07",X"07",X"E6",X"FC",X"4F",X"06",X"00",X"09",X"7E",X"32",X"00",X"60",
		X"23",X"7E",X"32",X"01",X"60",X"23",X"7E",X"32",X"02",X"60",X"3A",X"3B",X"42",X"3D",X"CA",X"AD",
		X"38",X"3D",X"CA",X"B3",X"38",X"3D",X"CA",X"B9",X"38",X"00",X"C3",X"BF",X"38",X"CD",X"00",X"3A",
		X"C3",X"F2",X"38",X"CD",X"11",X"3B",X"C3",X"F2",X"38",X"CD",X"E0",X"3B",X"C3",X"F2",X"38",X"00",
		X"3A",X"27",X"42",X"21",X"26",X"42",X"B6",X"C2",X"F2",X"38",X"3E",X"01",X"32",X"4F",X"41",X"0E",
		X"00",X"21",X"82",X"41",X"06",X"08",X"11",X"14",X"00",X"7E",X"B7",X"CA",X"DF",X"38",X"0C",X"19",
		X"05",X"C2",X"D9",X"38",X"79",X"32",X"3C",X"42",X"CD",X"81",X"39",X"AF",X"32",X"4D",X"42",X"CD",
		X"5A",X"39",X"21",X"27",X"42",X"34",X"7E",X"B7",X"C2",X"FD",X"38",X"2B",X"34",X"C9",X"01",X"00",
		X"04",X"03",X"04",X"05",X"06",X"00",X"06",X"02",X"03",X"00",X"05",X"00",X"05",X"02",X"07",X"03",
		X"07",X"05",X"03",X"00",X"08",X"00",X"08",X"02",X"02",X"00",X"01",X"00",X"03",X"00",X"06",X"02",
		X"05",X"02",X"03",X"00",X"04",X"05",X"03",X"00",X"08",X"00",X"07",X"03",X"02",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"01",X"01",X"00",X"01",X"01",
		X"01",X"00",X"00",X"21",X"00",X"50",X"06",X"20",X"0E",X"1C",X"23",X"23",X"23",X"36",X"24",X"23",
		X"0D",X"C2",X"4D",X"39",X"23",X"05",X"C2",X"48",X"39",X"C9",X"00",X"21",X"40",X"58",X"06",X"20",
		X"36",X"00",X"23",X"05",X"C2",X"60",X"39",X"C9",X"00",X"21",X"00",X"50",X"06",X"20",X"11",X"19",
		X"00",X"0E",X"06",X"19",X"36",X"24",X"23",X"0D",X"C2",X"74",X"39",X"23",X"05",X"C2",X"71",X"39",
		X"C9",X"00",X"21",X"82",X"41",X"06",X"08",X"0E",X"13",X"23",X"36",X"00",X"23",X"0D",X"C2",X"8A",
		X"39",X"05",X"C2",X"87",X"39",X"C9",X"00",X"21",X"82",X"41",X"06",X"08",X"0E",X"13",X"36",X"01",
		X"23",X"36",X"00",X"23",X"0D",X"C2",X"A1",X"39",X"05",X"C2",X"9C",X"39",X"C9",X"00",X"3A",X"27",
		X"42",X"0F",X"0F",X"0F",X"E6",X"1F",X"47",X"3A",X"26",X"42",X"07",X"07",X"07",X"07",X"07",X"E6",
		X"E0",X"B0",X"C9",X"00",X"3A",X"40",X"41",X"B8",X"C2",X"D0",X"39",X"79",X"32",X"40",X"41",X"C9",
		X"3A",X"45",X"41",X"B8",X"C2",X"DC",X"39",X"79",X"32",X"45",X"41",X"C9",X"3A",X"4A",X"41",X"B8",
		X"C0",X"79",X"32",X"4A",X"41",X"C9",X"00",X"3A",X"4A",X"41",X"B8",X"C2",X"F3",X"39",X"79",X"32",
		X"4A",X"41",X"C9",X"3A",X"45",X"41",X"B8",X"C2",X"FF",X"39",X"79",X"32",X"45",X"41",X"C9",X"C9",
		X"00",X"3A",X"27",X"42",X"E6",X"07",X"C0",X"CD",X"AD",X"39",X"B7",X"CA",X"41",X"3A",X"FE",X"01",
		X"CA",X"6F",X"3A",X"FE",X"03",X"CA",X"82",X"3A",X"FE",X"04",X"CA",X"8F",X"3A",X"FE",X"05",X"CA",
		X"9C",X"3A",X"FE",X"07",X"CA",X"A4",X"3A",X"FE",X"14",X"CA",X"AF",X"3A",X"FE",X"23",X"CA",X"C8",
		X"3A",X"FE",X"24",X"CA",X"DA",X"3A",X"FE",X"25",X"CA",X"E7",X"3A",X"FE",X"2F",X"CA",X"F9",X"3A",
		X"C9",X"CD",X"42",X"39",X"CD",X"5A",X"39",X"3E",X"0A",X"CD",X"92",X"08",X"3E",X"08",X"32",X"43",
		X"41",X"3E",X"00",X"32",X"48",X"41",X"32",X"4D",X"41",X"3E",X"78",X"32",X"44",X"41",X"3E",X"70",
		X"32",X"49",X"41",X"32",X"4E",X"41",X"3E",X"01",X"32",X"4D",X"42",X"CD",X"68",X"39",X"C9",X"3E",
		X"FF",X"32",X"2A",X"42",X"3A",X"40",X"41",X"FE",X"03",X"C0",X"06",X"03",X"0E",X"02",X"CD",X"C3",
		X"39",X"C9",X"3A",X"45",X"41",X"B7",X"C8",X"06",X"03",X"0E",X"02",X"CD",X"C3",X"39",X"C9",X"3A",
		X"45",X"41",X"B7",X"C0",X"06",X"03",X"0E",X"02",X"CD",X"C3",X"39",X"C9",X"06",X"03",X"0E",X"02",
		X"CD",X"C3",X"39",X"C9",X"3E",X"01",X"32",X"4F",X"41",X"3E",X"15",X"32",X"50",X"41",X"C9",X"3E",
		X"00",X"32",X"29",X"42",X"06",X"02",X"0E",X"01",X"CD",X"C3",X"39",X"3E",X"01",X"32",X"2A",X"42",
		X"AF",X"32",X"4F",X"41",X"CD",X"5A",X"39",X"C9",X"3A",X"45",X"41",X"B7",X"C8",X"3A",X"4A",X"41",
		X"B7",X"C8",X"06",X"02",X"0E",X"03",X"CD",X"E6",X"39",X"C9",X"3A",X"45",X"41",X"B7",X"C0",X"06",
		X"02",X"0E",X"03",X"CD",X"E6",X"39",X"C9",X"3E",X"01",X"32",X"29",X"42",X"3E",X"00",X"32",X"2A",
		X"42",X"06",X"02",X"0E",X"03",X"CD",X"C3",X"39",X"C9",X"AF",X"32",X"29",X"42",X"3A",X"9C",X"40",
		X"32",X"9B",X"40",X"21",X"26",X"42",X"36",X"FF",X"23",X"36",X"FF",X"3E",X"01",X"32",X"4F",X"41",
		X"C9",X"00",X"3A",X"27",X"42",X"E6",X"07",X"C0",X"CD",X"AD",X"39",X"B7",X"CA",X"2A",X"3B",X"FE",
		X"01",X"CA",X"4C",X"3B",X"FE",X"14",X"CA",X"53",X"3B",X"C9",X"3E",X"01",X"32",X"4D",X"42",X"AF",
		X"32",X"28",X"42",X"32",X"29",X"42",X"CD",X"50",X"29",X"3E",X"80",X"CD",X"B2",X"02",X"CD",X"68",
		X"39",X"3E",X"0D",X"CD",X"92",X"08",X"3E",X"FF",X"32",X"29",X"42",X"C9",X"11",X"CF",X"3B",X"CD",
		X"80",X"09",X"C9",X"3A",X"40",X"41",X"FE",X"01",X"C2",X"60",X"3B",X"3E",X"03",X"32",X"40",X"41",
		X"3A",X"45",X"41",X"FE",X"01",X"C2",X"6D",X"3B",X"3E",X"03",X"32",X"45",X"41",X"AF",X"32",X"29",
		X"42",X"3E",X"0E",X"CD",X"C3",X"2A",X"3A",X"4A",X"41",X"FE",X"01",X"C2",X"83",X"3B",X"3E",X"03",
		X"32",X"4A",X"41",X"3E",X"01",X"32",X"04",X"40",X"AF",X"32",X"59",X"41",X"32",X"5E",X"41",X"32",
		X"63",X"41",X"32",X"68",X"41",X"32",X"6D",X"41",X"CD",X"50",X"29",X"CD",X"5A",X"39",X"3E",X"FF",
		X"CD",X"B2",X"02",X"3E",X"FF",X"CD",X"B2",X"02",X"AF",X"32",X"28",X"42",X"32",X"29",X"42",X"32",
		X"4F",X"41",X"3A",X"9B",X"40",X"E6",X"F0",X"C6",X"10",X"F6",X"01",X"32",X"9B",X"40",X"3C",X"32",
		X"9C",X"40",X"3E",X"FF",X"32",X"26",X"42",X"32",X"27",X"42",X"AF",X"32",X"04",X"40",X"C9",X"0C",
		X"0E",X"09",X"0F",X"0A",X"1B",X"24",X"18",X"1E",X"1D",X"24",X"28",X"24",X"24",X"24",X"24",X"FF",
		X"00",X"3A",X"26",X"42",X"E6",X"F8",X"FE",X"01",X"D2",X"F3",X"3B",X"CD",X"AD",X"39",X"FE",X"3F",
		X"DA",X"F6",X"3B",X"CD",X"A8",X"3D",X"3A",X"27",X"42",X"E6",X"07",X"C0",X"3A",X"26",X"42",X"E6",
		X"F8",X"FE",X"02",X"D0",X"CD",X"AD",X"39",X"B7",X"CA",X"25",X"3C",X"FE",X"04",X"CA",X"29",X"3C",
		X"FE",X"06",X"CA",X"7D",X"3C",X"FE",X"2C",X"CA",X"8D",X"3C",X"FE",X"32",X"CA",X"C9",X"3C",X"FE",
		X"40",X"CA",X"CF",X"3C",X"C9",X"CD",X"50",X"29",X"C9",X"3A",X"45",X"41",X"FE",X"03",X"CA",X"49",
		X"3C",X"3A",X"4A",X"41",X"FE",X"03",X"CA",X"49",X"3C",X"3A",X"9B",X"40",X"3C",X"32",X"9B",X"40",
		X"3E",X"FF",X"32",X"26",X"42",X"32",X"27",X"42",X"C9",X"3E",X"80",X"32",X"22",X"42",X"32",X"23",
		X"42",X"3E",X"08",X"32",X"24",X"42",X"32",X"25",X"42",X"AF",X"32",X"28",X"42",X"32",X"29",X"42",
		X"3E",X"01",X"32",X"4D",X"42",X"CD",X"68",X"39",X"3A",X"36",X"40",X"B7",X"C2",X"76",X"3C",X"11",
		X"35",X"3D",X"CD",X"80",X"09",X"C9",X"11",X"E5",X"3C",X"CD",X"80",X"09",X"C9",X"3E",X"FF",X"32",
		X"29",X"42",X"3E",X"0F",X"CD",X"92",X"08",X"3E",X"15",X"32",X"55",X"41",X"C9",X"AF",X"32",X"29",
		X"42",X"3E",X"FF",X"32",X"2A",X"42",X"06",X"03",X"0E",X"02",X"CD",X"C3",X"39",X"AF",X"32",X"4F",
		X"41",X"3E",X"0E",X"CD",X"C3",X"2A",X"3E",X"30",X"32",X"30",X"42",X"3E",X"10",X"32",X"31",X"42",
		X"11",X"40",X"3D",X"CD",X"80",X"09",X"11",X"50",X"3D",X"CD",X"80",X"09",X"11",X"55",X"3D",X"CD",
		X"DD",X"09",X"11",X"5B",X"3D",X"CD",X"DD",X"09",X"C9",X"3E",X"01",X"32",X"4F",X"41",X"C9",X"AF",
		X"32",X"2A",X"42",X"3A",X"36",X"40",X"B7",X"C2",X"E1",X"3C",X"11",X"21",X"3D",X"CD",X"80",X"09",
		X"C9",X"11",X"E5",X"3C",X"C9",X"0C",X"0E",X"05",X"16",X"0A",X"14",X"0E",X"24",X"1B",X"18",X"0C",
		X"14",X"0E",X"1D",X"1C",X"24",X"0D",X"18",X"0C",X"14",X"FF",X"0C",X"10",X"07",X"16",X"0E",X"1C",
		X"1C",X"0A",X"10",X"0E",X"24",X"02",X"FF",X"0C",X"12",X"07",X"16",X"0E",X"1C",X"1C",X"0A",X"10",
		X"0E",X"24",X"02",X"FF",X"0C",X"14",X"07",X"16",X"0E",X"1C",X"1C",X"0A",X"10",X"0E",X"24",X"03",
		X"FF",X"0C",X"06",X"07",X"6E",X"6C",X"6A",X"68",X"66",X"64",X"62",X"60",X"24",X"6F",X"6D",X"6B",
		X"69",X"67",X"65",X"63",X"FF",X"0C",X"0E",X"0A",X"6F",X"6D",X"6B",X"69",X"67",X"65",X"63",X"FF",
		X"02",X"06",X"07",X"0D",X"18",X"0C",X"14",X"12",X"17",X"10",X"24",X"1D",X"12",X"16",X"0E",X"FF",
		X"0C",X"08",X"0C",X"2D",X"FF",X"07",X"08",X"0A",X"30",X"42",X"02",X"07",X"08",X"0D",X"31",X"42",
		X"01",X"00",X"3A",X"40",X"41",X"FE",X"01",X"C2",X"7E",X"3D",X"DD",X"21",X"40",X"41",X"DD",X"7E",
		X"04",X"C6",X"08",X"32",X"2B",X"42",X"DD",X"7E",X"03",X"C6",X"08",X"32",X"2C",X"42",X"3A",X"45",
		X"41",X"FE",X"01",X"C2",X"8D",X"3D",X"DD",X"21",X"45",X"41",X"C3",X"97",X"3D",X"3A",X"4A",X"41",
		X"FE",X"01",X"C0",X"DD",X"21",X"4A",X"41",X"DD",X"7E",X"04",X"C6",X"10",X"32",X"2B",X"42",X"DD",
		X"7E",X"03",X"C6",X"10",X"32",X"2C",X"42",X"C9",X"00",X"3A",X"27",X"42",X"E6",X"03",X"C0",X"21",
		X"31",X"42",X"7E",X"D6",X"01",X"27",X"77",X"C2",X"C2",X"3D",X"36",X"10",X"2B",X"7E",X"D6",X"01",
		X"27",X"77",X"21",X"30",X"42",X"7E",X"FE",X"00",X"C2",X"7C",X"3E",X"23",X"7E",X"FE",X"01",X"C2",
		X"7C",X"3E",X"AF",X"32",X"31",X"42",X"11",X"5B",X"3D",X"CD",X"DD",X"09",X"3E",X"0C",X"CD",X"92",
		X"08",X"11",X"89",X"3E",X"CD",X"80",X"09",X"3E",X"01",X"32",X"04",X"40",X"3E",X"FF",X"CD",X"B2",
		X"02",X"3E",X"FF",X"CD",X"B2",X"02",X"3E",X"FF",X"CD",X"B2",X"02",X"3E",X"06",X"CD",X"C3",X"2A",
		X"3E",X"08",X"CD",X"C3",X"2A",X"3A",X"45",X"41",X"FE",X"02",X"C2",X"29",X"3E",X"3E",X"03",X"32",
		X"45",X"41",X"3A",X"49",X"41",X"C6",X"08",X"32",X"44",X"41",X"3A",X"48",X"41",X"D6",X"08",X"32",
		X"43",X"41",X"AF",X"32",X"48",X"41",X"C3",X"61",X"3E",X"3E",X"03",X"32",X"4A",X"41",X"3A",X"4E",
		X"41",X"32",X"49",X"41",X"C6",X"08",X"32",X"44",X"41",X"3A",X"45",X"41",X"FE",X"01",X"C2",X"55",
		X"3E",X"3A",X"4D",X"41",X"D6",X"10",X"32",X"48",X"41",X"D6",X"08",X"32",X"43",X"41",X"AF",X"32",
		X"4D",X"41",X"C3",X"61",X"3E",X"3A",X"4D",X"41",X"D6",X"10",X"32",X"43",X"41",X"AF",X"32",X"4D",
		X"41",X"AF",X"32",X"28",X"42",X"32",X"29",X"42",X"3A",X"9B",X"40",X"3C",X"32",X"9B",X"40",X"3E",
		X"FF",X"32",X"26",X"42",X"32",X"27",X"42",X"AF",X"32",X"04",X"40",X"C9",X"11",X"55",X"3D",X"CD",
		X"DD",X"09",X"11",X"5B",X"3D",X"CD",X"DD",X"09",X"C9",X"0C",X"06",X"07",X"1C",X"18",X"1B",X"1B",
		X"22",X"24",X"17",X"18",X"24",X"0B",X"18",X"17",X"1E",X"1C",X"24",X"24",X"24",X"24",X"24",X"24",
		X"FF",X"00",X"9F",X"D3",X"04",X"21",X"00",X"00",X"CD",X"3C",X"B9",X"CD",X"21",X"B9",X"D3",X"04",
		X"AF",X"C9",X"C5",X"06",X"7F",X"3A",X"5B",X"B9",X"A7",X"28",X"02",X"06",X"7D",X"78",X"C1",X"C9",
		X"21",X"1F",X"00",X"3A",X"58",X"B9",X"E6",X"10",X"20",X"03",X"21",X"4B",X"00",X"2B",X"E3",X"E3",
		X"7D",X"B4",X"20",X"F9",X"C9",X"01",X"06",X"0B",X"10",X"03",X"08",X"0D",X"12",X"05",X"0A",X"0F",
		X"02",X"07",X"0C",X"11",X"04",X"09",X"0E",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"FF",X"FF",X"E4",X"BA",X"EE",X"BA",X"F0",X"BA",X"F6",X"BA",X"FC",X"BA",X"02",X"BB",
		X"7F",X"B9",X"00",X"63",X"B9",X"51",X"B5",X"68",X"93",X"68",X"93",X"00",X"01",X"03",X"AF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"38",X"9A",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
