library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity jng_snd_rom is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of jng_snd_rom is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"21",X"00",X"20",X"06",X"00",X"C3",X"B2",X"01",X"32",X"00",X"50",X"3A",X"00",X"40",X"C9",X"FF",
		X"32",X"00",X"70",X"3A",X"00",X"60",X"C9",X"FF",X"78",X"CF",X"79",X"32",X"00",X"40",X"C9",X"FF",
		X"78",X"D7",X"79",X"32",X"00",X"60",X"C9",X"FF",X"87",X"85",X"6F",X"7C",X"CE",X"00",X"67",X"7E",
		X"23",X"66",X"6F",X"E9",X"FF",X"FF",X"FF",X"FF",X"D9",X"08",X"CD",X"40",X"00",X"08",X"D9",X"C9",
		X"3E",X"0E",X"CF",X"B7",X"28",X"09",X"F2",X"79",X"00",X"CB",X"BF",X"CD",X"6C",X"00",X"C9",X"21",
		X"00",X"20",X"06",X"0C",X"AF",X"77",X"23",X"10",X"FC",X"C9",X"21",X"00",X"20",X"06",X"06",X"0E",
		X"07",X"BE",X"28",X"05",X"23",X"23",X"10",X"F9",X"41",X"79",X"90",X"C9",X"CD",X"5A",X"00",X"C8",
		X"AF",X"77",X"23",X"77",X"C9",X"13",X"23",X"22",X"28",X"32",X"1A",X"20",X"CD",X"5A",X"00",X"28",
		X"04",X"23",X"36",X"00",X"C9",X"3A",X"1A",X"20",X"21",X"75",X"00",X"06",X"02",X"BE",X"28",X"19",
		X"23",X"10",X"FA",X"06",X"02",X"BE",X"28",X"21",X"23",X"10",X"FA",X"AF",X"CD",X"5A",X"00",X"28",
		X"3A",X"3A",X"1A",X"20",X"77",X"23",X"36",X"00",X"C9",X"AF",X"CD",X"5A",X"00",X"28",X"05",X"FE",
		X"04",X"FA",X"C9",X"00",X"CD",X"37",X"01",X"18",X"58",X"AF",X"CD",X"5A",X"00",X"28",X"05",X"FE",
		X"04",X"F2",X"C9",X"00",X"CD",X"62",X"01",X"18",X"40",X"21",X"1A",X"20",X"46",X"0E",X"00",X"21",
		X"00",X"20",X"3D",X"87",X"5F",X"51",X"19",X"70",X"23",X"71",X"C9",X"CD",X"37",X"01",X"CD",X"62",
		X"01",X"B7",X"28",X"2D",X"3A",X"17",X"20",X"B7",X"28",X"1F",X"3A",X"18",X"20",X"21",X"06",X"20",
		X"CD",X"26",X"01",X"CD",X"2E",X"01",X"57",X"3A",X"17",X"20",X"21",X"00",X"20",X"CD",X"26",X"01",
		X"CD",X"2E",X"01",X"BA",X"F2",X"09",X"01",X"18",X"08",X"3A",X"18",X"20",X"21",X"06",X"20",X"18",
		X"06",X"3A",X"17",X"20",X"21",X"00",X"20",X"B7",X"C8",X"3D",X"87",X"4F",X"06",X"00",X"09",X"3A",
		X"1A",X"20",X"77",X"23",X"70",X"C9",X"3D",X"87",X"4F",X"06",X"00",X"09",X"7E",X"C9",X"21",X"87",
		X"07",X"06",X"00",X"4F",X"09",X"7E",X"C9",X"3A",X"00",X"20",X"CD",X"2E",X"01",X"32",X"12",X"20",
		X"3A",X"02",X"20",X"CD",X"2E",X"01",X"32",X"13",X"20",X"3A",X"04",X"20",X"CD",X"2E",X"01",X"32",
		X"14",X"20",X"3A",X"1A",X"20",X"CD",X"2E",X"01",X"32",X"15",X"20",X"CD",X"8D",X"01",X"32",X"17",
		X"20",X"C9",X"3A",X"06",X"20",X"CD",X"2E",X"01",X"32",X"12",X"20",X"3A",X"08",X"20",X"CD",X"2E",
		X"01",X"32",X"13",X"20",X"3A",X"0A",X"20",X"CD",X"2E",X"01",X"32",X"14",X"20",X"3A",X"1A",X"20",
		X"CD",X"2E",X"01",X"32",X"15",X"20",X"CD",X"8D",X"01",X"32",X"18",X"20",X"C9",X"21",X"12",X"20",
		X"3A",X"15",X"20",X"06",X"03",X"4F",X"7E",X"B9",X"F2",X"9C",X"01",X"4F",X"23",X"10",X"F7",X"79",
		X"06",X"03",X"0E",X"01",X"21",X"12",X"20",X"BE",X"28",X"06",X"0C",X"23",X"10",X"F9",X"0E",X"00",
		X"79",X"C9",X"70",X"23",X"7C",X"FE",X"24",X"20",X"F9",X"F9",X"ED",X"56",X"21",X"00",X"30",X"22",
		X"0C",X"20",X"77",X"01",X"3F",X"07",X"DF",X"E7",X"32",X"0E",X"20",X"32",X"0F",X"20",X"CD",X"C8",
		X"02",X"CD",X"CC",X"02",X"CD",X"D0",X"02",X"CD",X"D6",X"02",X"CD",X"DA",X"02",X"CD",X"DE",X"02",
		X"FB",X"3E",X"0F",X"CF",X"E6",X"80",X"20",X"F9",X"3E",X"0F",X"CF",X"E6",X"80",X"28",X"F9",X"F3",
		X"3E",X"01",X"32",X"10",X"20",X"3A",X"01",X"20",X"B7",X"3A",X"00",X"20",X"CA",X"04",X"02",X"CD",
		X"AC",X"02",X"18",X"03",X"CD",X"92",X"02",X"FB",X"00",X"00",X"F3",X"3E",X"02",X"32",X"10",X"20",
		X"3A",X"03",X"20",X"B7",X"3A",X"02",X"20",X"CA",X"1F",X"02",X"CD",X"AC",X"02",X"18",X"03",X"CD",
		X"92",X"02",X"FB",X"00",X"00",X"F3",X"3E",X"03",X"32",X"10",X"20",X"3A",X"05",X"20",X"B7",X"3A",
		X"04",X"20",X"CA",X"3A",X"02",X"CD",X"AC",X"02",X"18",X"03",X"CD",X"92",X"02",X"FB",X"00",X"00",
		X"F3",X"3E",X"04",X"32",X"10",X"20",X"3A",X"07",X"20",X"B7",X"3A",X"06",X"20",X"CA",X"55",X"02",
		X"CD",X"AC",X"02",X"18",X"03",X"CD",X"92",X"02",X"FB",X"00",X"00",X"F3",X"3E",X"05",X"32",X"10",
		X"20",X"3A",X"09",X"20",X"B7",X"3A",X"08",X"20",X"CA",X"70",X"02",X"CD",X"AC",X"02",X"18",X"03",
		X"CD",X"92",X"02",X"FB",X"00",X"00",X"F3",X"3E",X"06",X"32",X"10",X"20",X"3A",X"0B",X"20",X"B7",
		X"3A",X"0A",X"20",X"CA",X"8C",X"02",X"CD",X"AC",X"02",X"C3",X"E0",X"01",X"CD",X"92",X"02",X"C3",
		X"E0",X"01",X"21",X"A1",X"07",X"EF",X"B7",X"20",X"1B",X"E5",X"21",X"01",X"20",X"3A",X"10",X"20",
		X"3D",X"87",X"D5",X"5F",X"16",X"00",X"19",X"D1",X"36",X"01",X"E1",X"C9",X"B7",X"C8",X"21",X"D5",
		X"07",X"EF",X"B7",X"C8",X"57",X"21",X"00",X"20",X"3A",X"10",X"20",X"3D",X"4F",X"06",X"00",X"09",
		X"09",X"15",X"28",X"01",X"70",X"23",X"70",X"C9",X"06",X"08",X"18",X"06",X"06",X"09",X"18",X"02",
		X"06",X"0A",X"0E",X"00",X"DF",X"C9",X"06",X"08",X"18",X"06",X"06",X"09",X"18",X"02",X"06",X"0A",
		X"0E",X"00",X"E7",X"C9",X"3A",X"10",X"20",X"3D",X"21",X"ED",X"02",X"EF",X"C9",X"F9",X"02",X"02",
		X"03",X"0B",X"03",X"14",X"03",X"1D",X"03",X"26",X"03",X"CD",X"C8",X"02",X"0E",X"09",X"CD",X"2F",
		X"03",X"C9",X"CD",X"CC",X"02",X"0E",X"12",X"CD",X"2F",X"03",X"C9",X"CD",X"D0",X"02",X"0E",X"24",
		X"CD",X"2F",X"03",X"C9",X"CD",X"D6",X"02",X"0E",X"09",X"CD",X"3B",X"03",X"C9",X"CD",X"DA",X"02",
		X"0E",X"12",X"CD",X"3B",X"03",X"C9",X"CD",X"DE",X"02",X"0E",X"24",X"CD",X"3B",X"03",X"C9",X"3A",
		X"0E",X"20",X"B1",X"32",X"0E",X"20",X"06",X"07",X"4F",X"DF",X"C9",X"3A",X"0F",X"20",X"B1",X"32",
		X"0F",X"20",X"06",X"07",X"4F",X"E7",X"C9",X"06",X"06",X"3A",X"10",X"20",X"FE",X"04",X"FA",X"53",
		X"03",X"E7",X"C9",X"DF",X"C9",X"06",X"06",X"3A",X"10",X"20",X"FE",X"04",X"FA",X"63",X"03",X"78",
		X"D7",X"4F",X"C9",X"78",X"CF",X"4F",X"C9",X"3A",X"0E",X"20",X"A0",X"B1",X"32",X"0E",X"20",X"4F",
		X"06",X"07",X"DF",X"C9",X"3A",X"0F",X"20",X"A0",X"B1",X"32",X"0F",X"20",X"4F",X"06",X"07",X"E7",
		X"C9",X"3A",X"10",X"20",X"3D",X"21",X"8A",X"03",X"EF",X"C9",X"96",X"03",X"9D",X"03",X"A4",X"03",
		X"AB",X"03",X"B2",X"03",X"B9",X"03",X"01",X"08",X"FE",X"CD",X"67",X"03",X"C9",X"01",X"10",X"FD",
		X"CD",X"67",X"03",X"C9",X"01",X"20",X"FB",X"CD",X"67",X"03",X"C9",X"01",X"08",X"FE",X"CD",X"74",
		X"03",X"C9",X"01",X"10",X"FD",X"CD",X"74",X"03",X"C9",X"01",X"20",X"FB",X"CD",X"74",X"03",X"C9",
		X"3A",X"10",X"20",X"3D",X"21",X"C9",X"03",X"EF",X"C9",X"D5",X"03",X"DC",X"03",X"E3",X"03",X"EA",
		X"03",X"F1",X"03",X"F8",X"03",X"01",X"01",X"F7",X"CD",X"67",X"03",X"C9",X"01",X"02",X"EF",X"CD",
		X"67",X"03",X"C9",X"01",X"04",X"DF",X"CD",X"67",X"03",X"C9",X"01",X"01",X"F7",X"CD",X"74",X"03",
		X"C9",X"01",X"02",X"EF",X"CD",X"74",X"03",X"C9",X"01",X"04",X"DF",X"CD",X"74",X"03",X"C9",X"3A",
		X"10",X"20",X"3D",X"21",X"08",X"04",X"EF",X"C9",X"14",X"04",X"1B",X"04",X"22",X"04",X"29",X"04",
		X"30",X"04",X"37",X"04",X"01",X"00",X"F6",X"CD",X"67",X"03",X"C9",X"01",X"00",X"ED",X"CD",X"67",
		X"03",X"C9",X"01",X"00",X"DB",X"CD",X"67",X"03",X"C9",X"01",X"00",X"F6",X"CD",X"74",X"03",X"C9",
		X"01",X"00",X"ED",X"CD",X"74",X"03",X"C9",X"01",X"00",X"DB",X"CD",X"74",X"03",X"C9",X"3A",X"10",
		X"20",X"FE",X"04",X"30",X"05",X"C6",X"07",X"47",X"DF",X"C9",X"C6",X"04",X"47",X"E7",X"C9",X"3A",
		X"10",X"20",X"FE",X"04",X"30",X"04",X"C6",X"07",X"CF",X"C9",X"C6",X"04",X"D7",X"C9",X"3A",X"10",
		X"20",X"FE",X"04",X"30",X"09",X"3D",X"87",X"47",X"4D",X"DF",X"4C",X"04",X"DF",X"C9",X"D6",X"04",
		X"87",X"47",X"4D",X"E7",X"4C",X"04",X"E7",X"C9",X"3A",X"10",X"20",X"FE",X"04",X"30",X"0A",X"3D",
		X"87",X"67",X"24",X"CF",X"6F",X"7C",X"CF",X"67",X"C9",X"D6",X"04",X"87",X"67",X"24",X"D7",X"6F",
		X"7C",X"D7",X"67",X"C9",X"FE",X"04",X"D0",X"F5",X"CD",X"E4",X"04",X"F1",X"B7",X"20",X"02",X"77",
		X"C9",X"21",X"B4",X"04",X"87",X"87",X"4F",X"87",X"81",X"4F",X"06",X"00",X"09",X"3A",X"10",X"20",
		X"3D",X"EF",X"77",X"C9",X"07",X"05",X"0C",X"05",X"11",X"05",X"16",X"05",X"1B",X"05",X"20",X"05",
		X"25",X"05",X"2A",X"05",X"2F",X"05",X"34",X"05",X"39",X"05",X"3E",X"05",X"43",X"05",X"48",X"05",
		X"4D",X"05",X"52",X"05",X"57",X"05",X"5C",X"05",X"61",X"05",X"66",X"05",X"6B",X"05",X"70",X"05",
		X"75",X"05",X"7A",X"05",X"21",X"B4",X"04",X"3A",X"10",X"20",X"3D",X"EF",X"C9",X"2A",X"0C",X"20",
		X"7B",X"A5",X"6F",X"7A",X"A4",X"67",X"22",X"0C",X"20",X"C9",X"2A",X"0C",X"20",X"7B",X"B5",X"6F",
		X"7A",X"B4",X"67",X"22",X"0C",X"20",X"C9",X"11",X"3F",X"FF",X"18",X"E1",X"11",X"FF",X"FC",X"18",
		X"DC",X"11",X"FF",X"F3",X"18",X"D7",X"11",X"FC",X"FF",X"18",X"D2",X"11",X"F3",X"FF",X"18",X"CD",
		X"11",X"CF",X"FF",X"18",X"C8",X"11",X"80",X"00",X"18",X"D0",X"11",X"00",X"02",X"18",X"CB",X"11",
		X"00",X"08",X"18",X"C6",X"11",X"02",X"00",X"18",X"C1",X"11",X"08",X"00",X"18",X"BC",X"11",X"20",
		X"00",X"18",X"B7",X"11",X"40",X"00",X"18",X"B2",X"11",X"00",X"01",X"18",X"AD",X"11",X"00",X"04",
		X"18",X"A8",X"11",X"01",X"00",X"18",X"A3",X"11",X"04",X"00",X"18",X"9E",X"11",X"10",X"00",X"18",
		X"99",X"11",X"C0",X"00",X"18",X"94",X"11",X"00",X"03",X"18",X"8F",X"11",X"00",X"0C",X"18",X"8A",
		X"11",X"03",X"00",X"18",X"85",X"11",X"0C",X"00",X"18",X"80",X"11",X"30",X"00",X"C3",X"FA",X"04",
		X"DD",X"7E",X"00",X"FE",X"FF",X"C8",X"CD",X"8B",X"05",X"AF",X"C9",X"DD",X"35",X"01",X"C0",X"3A",
		X"42",X"20",X"DD",X"77",X"01",X"DD",X"CB",X"00",X"46",X"C2",X"AB",X"05",X"DD",X"7E",X"07",X"D6",
		X"01",X"FA",X"AB",X"05",X"DD",X"77",X"07",X"4F",X"CD",X"3E",X"04",X"DD",X"35",X"00",X"C0",X"DD",
		X"6E",X"02",X"DD",X"66",X"03",X"7E",X"47",X"E6",X"1F",X"CA",X"46",X"06",X"FE",X"1F",X"C2",X"62",
		X"06",X"23",X"DD",X"75",X"02",X"DD",X"74",X"03",X"78",X"E6",X"E0",X"0F",X"0F",X"0F",X"0F",X"4F",
		X"06",X"00",X"21",X"DB",X"05",X"09",X"5E",X"23",X"56",X"EB",X"E9",X"EB",X"05",X"09",X"06",X"1F",
		X"06",X"3C",X"06",X"3C",X"06",X"3C",X"06",X"3C",X"06",X"3C",X"06",X"DD",X"6E",X"02",X"DD",X"66",
		X"03",X"4E",X"CB",X"21",X"06",X"00",X"21",X"95",X"06",X"09",X"5E",X"23",X"56",X"ED",X"53",X"40",
		X"20",X"DD",X"73",X"04",X"DD",X"72",X"05",X"18",X"23",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"4E",
		X"06",X"00",X"21",X"2D",X"07",X"09",X"7E",X"32",X"42",X"20",X"DD",X"77",X"01",X"18",X"0D",X"DD",
		X"6E",X"02",X"DD",X"66",X"03",X"7E",X"DD",X"77",X"06",X"DD",X"77",X"07",X"DD",X"6E",X"02",X"DD",
		X"66",X"03",X"23",X"DD",X"75",X"02",X"DD",X"74",X"03",X"C3",X"AF",X"05",X"0E",X"00",X"CD",X"3E",
		X"04",X"DD",X"36",X"00",X"FF",X"C9",X"CD",X"50",X"06",X"0E",X"00",X"CD",X"3E",X"04",X"18",X"37",
		X"78",X"E6",X"E0",X"07",X"07",X"07",X"47",X"3E",X"01",X"18",X"01",X"07",X"10",X"FD",X"DD",X"77",
		X"00",X"C9",X"C5",X"CD",X"50",X"06",X"C1",X"78",X"E6",X"1F",X"3D",X"07",X"4F",X"06",X"00",X"DD",
		X"6E",X"04",X"DD",X"66",X"05",X"09",X"5E",X"23",X"56",X"EB",X"CD",X"5E",X"04",X"DD",X"4E",X"06",
		X"79",X"DD",X"77",X"07",X"CD",X"3E",X"04",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"23",X"DD",X"75",
		X"02",X"DD",X"74",X"03",X"C9",X"B5",X"06",X"B9",X"06",X"BD",X"06",X"C1",X"06",X"C5",X"06",X"C9",
		X"06",X"CD",X"06",X"D1",X"06",X"D5",X"06",X"D9",X"06",X"DD",X"06",X"E1",X"06",X"E5",X"06",X"E9",
		X"06",X"ED",X"06",X"F1",X"06",X"6B",X"08",X"F2",X"07",X"80",X"07",X"14",X"07",X"AE",X"06",X"4E",
		X"06",X"F3",X"05",X"9E",X"05",X"4E",X"05",X"01",X"05",X"B9",X"04",X"76",X"04",X"36",X"04",X"F9",
		X"03",X"C0",X"03",X"8A",X"03",X"57",X"03",X"27",X"03",X"FA",X"02",X"CF",X"02",X"A7",X"02",X"81",
		X"02",X"5D",X"02",X"3B",X"02",X"1B",X"02",X"FD",X"01",X"E0",X"01",X"C5",X"01",X"AC",X"01",X"94",
		X"01",X"7D",X"01",X"68",X"01",X"53",X"01",X"40",X"01",X"2E",X"01",X"1D",X"01",X"0D",X"01",X"FE",
		X"00",X"F0",X"00",X"E3",X"00",X"D6",X"00",X"CA",X"00",X"BE",X"00",X"B4",X"00",X"AA",X"00",X"A0",
		X"00",X"97",X"00",X"8F",X"00",X"87",X"00",X"7F",X"00",X"78",X"00",X"71",X"00",X"6B",X"00",X"65",
		X"00",X"5F",X"00",X"5A",X"00",X"55",X"00",X"50",X"00",X"4C",X"00",X"47",X"00",X"57",X"42",X"34",
		X"2C",X"25",X"21",X"1D",X"1A",X"0C",X"0B",X"0A",X"09",X"08",X"07",X"06",X"05",X"21",X"6F",X"07",
		X"11",X"20",X"20",X"01",X"18",X"00",X"ED",X"B0",X"3A",X"43",X"20",X"07",X"4F",X"07",X"81",X"4F",
		X"06",X"00",X"21",X"01",X"0D",X"09",X"11",X"22",X"20",X"CD",X"65",X"07",X"11",X"2A",X"20",X"CD",
		X"65",X"07",X"11",X"32",X"20",X"7E",X"12",X"CD",X"6C",X"07",X"7E",X"12",X"23",X"13",X"C9",X"01",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"0E",X"07",X"06",X"01",X"04",X"03",X"05",
		X"0C",X"02",X"0A",X"09",X"08",X"0D",X"0F",X"11",X"12",X"13",X"14",X"15",X"16",X"17",X"18",X"19",
		X"0B",X"E4",X"02",X"09",X"08",X"43",X"08",X"71",X"08",X"D3",X"08",X"1A",X"09",X"AB",X"09",X"F5",
		X"09",X"57",X"0A",X"BC",X"0A",X"FD",X"0A",X"60",X"0B",X"B0",X"0B",X"F7",X"0B",X"2E",X"0C",X"74",
		X"0C",X"13",X"0D",X"17",X"0D",X"19",X"0D",X"21",X"0D",X"25",X"0D",X"27",X"0D",X"2F",X"0D",X"33",
		X"0D",X"35",X"0D",X"C5",X"0C",X"00",X"00",X"24",X"08",X"64",X"08",X"92",X"08",X"EB",X"08",X"40",
		X"09",X"C3",X"09",X"12",X"0A",X"77",X"0A",X"D5",X"0A",X"1F",X"0B",X"7A",X"0B",X"CA",X"0B",X"11",
		X"0C",X"4B",X"0C",X"8F",X"0C",X"1B",X"0D",X"1D",X"0D",X"1F",X"0D",X"29",X"0D",X"2B",X"0D",X"2D",
		X"0D",X"37",X"0D",X"39",X"0D",X"3B",X"0D",X"E2",X"0C",X"3E",X"03",X"CD",X"94",X"04",X"CD",X"81",
		X"03",X"21",X"00",X"01",X"CD",X"5E",X"04",X"0E",X"0C",X"CD",X"3E",X"04",X"AF",X"32",X"51",X"20",
		X"32",X"50",X"20",X"C9",X"3A",X"50",X"20",X"3D",X"32",X"50",X"20",X"E6",X"03",X"20",X"12",X"CD",
		X"78",X"04",X"3A",X"51",X"20",X"C6",X"DB",X"32",X"51",X"20",X"AD",X"E6",X"7F",X"6F",X"CD",X"5E",
		X"04",X"AF",X"C9",X"3E",X"01",X"CD",X"94",X"04",X"CD",X"81",X"03",X"0E",X"10",X"CD",X"3E",X"04",
		X"21",X"40",X"0D",X"CD",X"5E",X"04",X"CD",X"4F",X"04",X"3D",X"FE",X"04",X"28",X"11",X"4F",X"CD",
		X"3E",X"04",X"AF",X"C9",X"CD",X"78",X"04",X"2D",X"28",X"E6",X"CD",X"5E",X"04",X"AF",X"C9",X"3D",
		X"C9",X"3E",X"01",X"CD",X"94",X"04",X"CD",X"FF",X"03",X"01",X"1F",X"06",X"CD",X"49",X"03",X"21",
		X"00",X"04",X"CD",X"5E",X"04",X"0E",X"0F",X"CD",X"3E",X"04",X"AF",X"32",X"53",X"20",X"32",X"52",
		X"20",X"C9",X"21",X"52",X"20",X"35",X"56",X"CD",X"78",X"04",X"3A",X"53",X"20",X"C6",X"B5",X"32",
		X"53",X"20",X"AD",X"6F",X"7A",X"E6",X"0F",X"20",X"05",X"25",X"20",X"02",X"26",X"01",X"CD",X"5E",
		X"04",X"7A",X"E6",X"3F",X"20",X"19",X"7C",X"FE",X"01",X"20",X"14",X"06",X"06",X"CD",X"57",X"03",
		X"0D",X"0D",X"CD",X"49",X"03",X"CD",X"4F",X"04",X"3D",X"28",X"06",X"4F",X"CD",X"3E",X"04",X"AF",
		X"C9",X"3D",X"C9",X"3E",X"00",X"CD",X"94",X"04",X"CD",X"81",X"03",X"21",X"40",X"00",X"CD",X"5E",
		X"04",X"3E",X"20",X"32",X"55",X"20",X"AF",X"32",X"54",X"20",X"C9",X"3A",X"55",X"20",X"3D",X"32",
		X"55",X"20",X"20",X"02",X"3D",X"C9",X"CB",X"47",X"28",X"07",X"0E",X"0C",X"CD",X"3E",X"04",X"AF",
		X"C9",X"CD",X"78",X"04",X"3A",X"54",X"20",X"3C",X"32",X"54",X"20",X"85",X"6F",X"30",X"01",X"24",
		X"CD",X"5E",X"04",X"0E",X"00",X"CD",X"3E",X"04",X"AF",X"C9",X"AF",X"CD",X"94",X"04",X"CD",X"81",
		X"03",X"21",X"40",X"00",X"CD",X"5E",X"04",X"0E",X"00",X"CD",X"3E",X"04",X"3E",X"08",X"32",X"59",
		X"20",X"32",X"58",X"20",X"3E",X"DB",X"32",X"56",X"20",X"3E",X"AA",X"32",X"57",X"20",X"AF",X"C9",
		X"3A",X"56",X"20",X"3D",X"32",X"56",X"20",X"20",X"02",X"3D",X"C9",X"FE",X"C3",X"38",X"24",X"28",
		X"15",X"FE",X"CF",X"38",X"0A",X"CD",X"4F",X"04",X"3C",X"4F",X"CD",X"3E",X"04",X"AF",X"C9",X"0E",
		X"00",X"CD",X"3E",X"04",X"AF",X"C9",X"0E",X"0C",X"CD",X"3E",X"04",X"21",X"1F",X"00",X"CD",X"5E",
		X"04",X"AF",X"C9",X"3A",X"58",X"20",X"3D",X"32",X"58",X"20",X"28",X"02",X"AF",X"C9",X"3A",X"59",
		X"20",X"32",X"58",X"20",X"21",X"57",X"20",X"CB",X"0E",X"38",X"0C",X"CD",X"78",X"04",X"3E",X"20",
		X"85",X"6F",X"CD",X"5E",X"04",X"AF",X"C9",X"CD",X"78",X"04",X"3E",X"E0",X"85",X"6F",X"CD",X"5E",
		X"04",X"CD",X"4F",X"04",X"3D",X"4F",X"CD",X"3E",X"04",X"AF",X"C9",X"3E",X"00",X"CD",X"94",X"04",
		X"CD",X"81",X"03",X"21",X"30",X"00",X"CD",X"5E",X"04",X"0E",X"08",X"CD",X"3E",X"04",X"AF",X"32",
		X"5A",X"20",X"C9",X"21",X"5A",X"20",X"35",X"7E",X"28",X"29",X"57",X"FE",X"E8",X"28",X"0C",X"38",
		X"11",X"CD",X"4F",X"04",X"3D",X"4F",X"CD",X"3E",X"04",X"AF",X"C9",X"0E",X"0F",X"CD",X"3E",X"04",
		X"AF",X"C9",X"CD",X"78",X"04",X"01",X"02",X"00",X"09",X"CD",X"5E",X"04",X"7A",X"E6",X"0F",X"28",
		X"E0",X"AF",X"C9",X"3D",X"C9",X"AF",X"CD",X"94",X"04",X"CD",X"81",X"03",X"0E",X"0C",X"CD",X"3E",
		X"04",X"21",X"90",X"00",X"CD",X"5E",X"04",X"AF",X"32",X"5B",X"20",X"3E",X"AA",X"32",X"5C",X"20",
		X"AF",X"C9",X"21",X"5C",X"20",X"CB",X"0E",X"30",X"02",X"AF",X"C9",X"3A",X"5B",X"20",X"3D",X"32",
		X"5B",X"20",X"FE",X"EC",X"38",X"18",X"FE",X"F6",X"28",X"0C",X"CD",X"78",X"04",X"3E",X"F0",X"85",
		X"6F",X"CD",X"5E",X"04",X"AF",X"C9",X"21",X"90",X"00",X"CD",X"5E",X"04",X"AF",X"C9",X"CD",X"78",
		X"04",X"3E",X"10",X"85",X"6F",X"CD",X"5E",X"04",X"CD",X"4F",X"04",X"D6",X"02",X"20",X"02",X"3D",
		X"C9",X"4F",X"CD",X"3E",X"04",X"AF",X"C9",X"3E",X"01",X"CD",X"94",X"04",X"CD",X"81",X"03",X"21",
		X"00",X"05",X"CD",X"5E",X"04",X"0E",X"0E",X"CD",X"3E",X"04",X"3E",X"02",X"32",X"5E",X"20",X"AF",
		X"32",X"5F",X"20",X"32",X"5D",X"20",X"C9",X"3A",X"5E",X"20",X"3D",X"32",X"5E",X"20",X"20",X"28",
		X"3E",X"02",X"32",X"5E",X"20",X"21",X"5D",X"20",X"35",X"28",X"1F",X"7E",X"57",X"CD",X"78",X"04",
		X"7A",X"FE",X"E0",X"38",X"18",X"E6",X"07",X"20",X"01",X"25",X"3A",X"5F",X"20",X"C6",X"C3",X"32",
		X"5F",X"20",X"AA",X"AD",X"6F",X"CD",X"5E",X"04",X"AF",X"C9",X"3E",X"FF",X"C9",X"E6",X"0F",X"20",
		X"E9",X"CD",X"4F",X"04",X"3D",X"4F",X"CD",X"3E",X"04",X"C3",X"9A",X"0A",X"AF",X"CD",X"94",X"04",
		X"CD",X"81",X"03",X"21",X"C0",X"01",X"CD",X"5E",X"04",X"0E",X"0F",X"CD",X"3E",X"04",X"3E",X"48",
		X"32",X"60",X"20",X"AF",X"C9",X"3A",X"60",X"20",X"3D",X"32",X"60",X"20",X"20",X"02",X"3D",X"C9",
		X"FE",X"02",X"38",X"12",X"E6",X"07",X"28",X"02",X"AF",X"C9",X"CD",X"78",X"04",X"01",X"D4",X"FF",
		X"09",X"CD",X"5E",X"04",X"AF",X"C9",X"0E",X"0F",X"CD",X"3E",X"04",X"AF",X"C9",X"3E",X"01",X"CD",
		X"94",X"04",X"CD",X"81",X"03",X"21",X"40",X"00",X"CD",X"5E",X"04",X"0E",X"03",X"CD",X"3E",X"04",
		X"3E",X"20",X"32",X"61",X"20",X"32",X"62",X"20",X"3E",X"08",X"32",X"63",X"20",X"AF",X"C9",X"3A",
		X"62",X"20",X"3D",X"32",X"62",X"20",X"28",X"25",X"FE",X"1A",X"28",X"0C",X"38",X"11",X"CD",X"4F",
		X"04",X"C6",X"02",X"CD",X"3E",X"04",X"AF",X"C9",X"0E",X"0F",X"CD",X"3E",X"04",X"AF",X"C9",X"E6",
		X"01",X"28",X"08",X"CD",X"4F",X"04",X"3D",X"4F",X"CD",X"3E",X"04",X"AF",X"C9",X"3A",X"63",X"20",
		X"3D",X"32",X"63",X"20",X"20",X"02",X"3D",X"C9",X"3A",X"61",X"20",X"32",X"62",X"20",X"AF",X"C9",
		X"3E",X"01",X"CD",X"94",X"04",X"CD",X"81",X"03",X"0E",X"0E",X"CD",X"3E",X"04",X"21",X"FF",X"00",
		X"CD",X"5E",X"04",X"3E",X"40",X"32",X"64",X"20",X"AF",X"C9",X"3A",X"64",X"20",X"3D",X"32",X"64",
		X"20",X"20",X"02",X"3D",X"C9",X"E6",X"07",X"20",X"08",X"CD",X"4F",X"04",X"3D",X"4F",X"CD",X"3E",
		X"04",X"3A",X"64",X"20",X"E6",X"08",X"28",X"0C",X"CD",X"78",X"04",X"3E",X"F0",X"85",X"6F",X"CD",
		X"5E",X"04",X"AF",X"C9",X"CD",X"78",X"04",X"3E",X"10",X"85",X"6F",X"CD",X"5E",X"04",X"AF",X"C9",
		X"3E",X"00",X"CD",X"94",X"04",X"CD",X"81",X"03",X"21",X"7C",X"00",X"CD",X"5E",X"04",X"0E",X"0F",
		X"CD",X"3E",X"04",X"3E",X"3F",X"32",X"65",X"20",X"AF",X"C9",X"21",X"65",X"20",X"35",X"7E",X"28",
		X"24",X"FE",X"11",X"38",X"15",X"FE",X"30",X"38",X"08",X"CD",X"4F",X"04",X"3D",X"4F",X"CD",X"3E",
		X"04",X"CD",X"78",X"04",X"2D",X"CD",X"5E",X"04",X"AF",X"C9",X"E6",X"02",X"0E",X"07",X"28",X"EE",
		X"0E",X"0F",X"C3",X"DE",X"0B",X"3D",X"C9",X"3E",X"00",X"CD",X"94",X"04",X"CD",X"81",X"03",X"0E",
		X"0D",X"CD",X"3E",X"04",X"21",X"FF",X"00",X"CD",X"5E",X"04",X"3E",X"0F",X"32",X"66",X"20",X"AF",
		X"C9",X"3A",X"66",X"20",X"3D",X"32",X"66",X"20",X"28",X"02",X"AF",X"C9",X"3E",X"0F",X"32",X"66",
		X"20",X"CD",X"78",X"04",X"3E",X"F0",X"85",X"D0",X"6F",X"CD",X"5E",X"04",X"AF",X"C9",X"3E",X"00",
		X"CD",X"94",X"04",X"CD",X"81",X"03",X"21",X"90",X"00",X"CD",X"5E",X"04",X"0E",X"09",X"CD",X"3E",
		X"04",X"3E",X"F4",X"32",X"68",X"20",X"AF",X"32",X"67",X"20",X"C9",X"21",X"67",X"20",X"35",X"7E",
		X"E6",X"07",X"20",X"11",X"CD",X"78",X"04",X"3A",X"68",X"20",X"3C",X"28",X"15",X"32",X"68",X"20",
		X"85",X"6F",X"CD",X"5E",X"04",X"7E",X"E6",X"08",X"0E",X"09",X"20",X"01",X"4F",X"CD",X"3E",X"04",
		X"AF",X"C9",X"3D",X"C9",X"3E",X"01",X"CD",X"94",X"04",X"CD",X"81",X"03",X"21",X"D0",X"00",X"CD",
		X"5E",X"04",X"3E",X"08",X"32",X"69",X"20",X"32",X"6A",X"20",X"AF",X"32",X"6B",X"20",X"C9",X"3A",
		X"6A",X"20",X"3D",X"57",X"32",X"6A",X"20",X"20",X"1E",X"3A",X"69",X"20",X"32",X"6A",X"20",X"CD",
		X"78",X"04",X"3A",X"6B",X"20",X"3C",X"32",X"6B",X"20",X"FE",X"4E",X"20",X"03",X"3E",X"FF",X"C9",
		X"4F",X"06",X"00",X"09",X"CD",X"5E",X"04",X"7A",X"E6",X"02",X"0E",X"03",X"28",X"02",X"0E",X"0C",
		X"CD",X"3E",X"04",X"AF",X"C9",X"3E",X"01",X"CD",X"94",X"04",X"CD",X"81",X"03",X"0E",X"0E",X"CD",
		X"3E",X"04",X"3E",X"05",X"32",X"6D",X"20",X"21",X"04",X"00",X"CD",X"5E",X"04",X"AF",X"32",X"6C",
		X"20",X"C9",X"21",X"6C",X"20",X"35",X"7E",X"28",X"16",X"FE",X"DA",X"20",X"06",X"21",X"6D",X"20",
		X"35",X"20",X"E4",X"CD",X"78",X"04",X"01",X"0C",X"00",X"09",X"CD",X"5E",X"04",X"AF",X"C9",X"3D",
		X"C9",X"6A",X"0D",X"91",X"0D",X"B6",X"0D",X"D7",X"0D",X"17",X"0E",X"37",X"0E",X"49",X"0E",X"5E",
		X"0E",X"71",X"0E",X"3E",X"00",X"18",X"26",X"18",X"33",X"18",X"31",X"18",X"38",X"18",X"3D",X"18",
		X"42",X"3E",X"01",X"18",X"18",X"18",X"25",X"18",X"23",X"18",X"2A",X"18",X"2F",X"18",X"34",X"3E",
		X"02",X"18",X"0A",X"18",X"17",X"18",X"15",X"18",X"1C",X"18",X"21",X"18",X"26",X"32",X"43",X"20",
		X"CD",X"3D",X"07",X"AF",X"CD",X"94",X"04",X"CD",X"81",X"03",X"AF",X"C9",X"AF",X"CD",X"94",X"04",
		X"CD",X"81",X"03",X"AF",X"C9",X"DD",X"21",X"20",X"20",X"C3",X"80",X"05",X"DD",X"21",X"28",X"20",
		X"C3",X"80",X"05",X"DD",X"21",X"30",X"20",X"C3",X"80",X"05",X"1F",X"0E",X"3F",X"0B",X"5F",X"09",
		X"6D",X"6F",X"72",X"6D",X"6F",X"72",X"6D",X"6F",X"6F",X"71",X"74",X"6F",X"71",X"74",X"6F",X"74",
		X"72",X"72",X"72",X"74",X"74",X"74",X"36",X"36",X"36",X"36",X"36",X"36",X"36",X"36",X"B6",X"A0",
		X"FF",X"1F",X"0E",X"5F",X"09",X"6A",X"6B",X"6F",X"6A",X"6B",X"6F",X"6A",X"6B",X"6C",X"6D",X"71",
		X"6C",X"6D",X"71",X"6C",X"6D",X"6F",X"6F",X"6F",X"70",X"70",X"70",X"32",X"32",X"32",X"32",X"32",
		X"32",X"32",X"32",X"B2",X"A0",X"FF",X"1F",X"05",X"5F",X"09",X"8C",X"60",X"8C",X"60",X"6C",X"6C",
		X"8E",X"60",X"8E",X"60",X"6E",X"6E",X"69",X"69",X"69",X"6A",X"6A",X"6A",X"2C",X"2C",X"2C",X"2C",
		X"2C",X"2C",X"2C",X"2C",X"AC",X"A0",X"FF",X"1F",X"0E",X"3F",X"0C",X"5F",X"09",X"70",X"70",X"60",
		X"70",X"90",X"71",X"71",X"60",X"71",X"91",X"93",X"91",X"70",X"71",X"70",X"71",X"90",X"71",X"73",
		X"71",X"73",X"91",X"93",X"91",X"2E",X"2F",X"30",X"31",X"2F",X"30",X"31",X"32",X"30",X"31",X"32",
		X"33",X"31",X"32",X"33",X"34",X"32",X"33",X"34",X"35",X"33",X"34",X"35",X"36",X"34",X"35",X"36",
		X"37",X"35",X"36",X"37",X"38",X"A0",X"FF",X"1F",X"0E",X"5F",X"09",X"6C",X"6C",X"60",X"6C",X"8C",
		X"6E",X"6E",X"60",X"6E",X"8E",X"90",X"8E",X"6C",X"6E",X"6C",X"6E",X"8C",X"6E",X"70",X"6E",X"70",
		X"8E",X"90",X"8E",X"A0",X"A0",X"A0",X"FF",X"1F",X"08",X"5F",X"09",X"AC",X"A0",X"A0",X"80",X"87",
		X"AC",X"A0",X"A0",X"80",X"87",X"A0",X"A0",X"A0",X"FF",X"1F",X"0E",X"3F",X"0B",X"5F",X"09",X"69",
		X"69",X"60",X"6C",X"60",X"69",X"60",X"67",X"89",X"8C",X"6E",X"70",X"73",X"B5",X"FF",X"1F",X"08",
		X"5F",X"09",X"69",X"69",X"60",X"6C",X"60",X"69",X"60",X"67",X"89",X"8C",X"6E",X"70",X"73",X"B5",
		X"FF",X"1F",X"02",X"5F",X"08",X"69",X"69",X"60",X"6C",X"60",X"69",X"60",X"67",X"89",X"8C",X"6E",
		X"70",X"73",X"B5",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
