library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity cclimber_tile_bit0 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of cclimber_tile_bit0 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1C",X"36",X"63",X"63",X"7F",X"63",X"63",X"00",X"7E",X"63",X"63",X"7E",X"63",X"63",X"7E",X"00",
		X"1E",X"33",X"60",X"60",X"60",X"33",X"1E",X"00",X"7C",X"66",X"63",X"63",X"63",X"66",X"7C",X"00",
		X"3F",X"30",X"30",X"3E",X"30",X"30",X"3F",X"00",X"7F",X"60",X"60",X"7E",X"60",X"60",X"60",X"00",
		X"1F",X"30",X"60",X"67",X"63",X"33",X"1F",X"00",X"63",X"63",X"63",X"7F",X"63",X"63",X"63",X"00",
		X"3F",X"0C",X"0C",X"0C",X"0C",X"0C",X"3F",X"00",X"03",X"03",X"03",X"03",X"03",X"63",X"3E",X"00",
		X"63",X"66",X"6C",X"78",X"7C",X"6E",X"67",X"00",X"30",X"30",X"30",X"30",X"30",X"30",X"3F",X"00",
		X"63",X"77",X"7F",X"7F",X"6B",X"63",X"63",X"00",X"63",X"73",X"7B",X"7F",X"6F",X"67",X"63",X"00",
		X"3E",X"63",X"63",X"63",X"63",X"63",X"3E",X"00",X"7E",X"63",X"63",X"63",X"7E",X"60",X"60",X"00",
		X"3E",X"63",X"63",X"63",X"6F",X"66",X"3D",X"00",X"7E",X"63",X"63",X"67",X"7C",X"6E",X"67",X"00",
		X"3C",X"66",X"60",X"3E",X"03",X"63",X"3E",X"00",X"3F",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"00",
		X"63",X"63",X"63",X"63",X"63",X"63",X"3E",X"00",X"63",X"63",X"63",X"77",X"3E",X"1C",X"08",X"00",
		X"63",X"63",X"6B",X"7F",X"7F",X"36",X"22",X"00",X"63",X"77",X"3E",X"1C",X"3E",X"77",X"63",X"00",
		X"33",X"33",X"12",X"1E",X"0C",X"0C",X"0C",X"00",X"7F",X"07",X"0E",X"1C",X"38",X"70",X"7F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"06",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",
		X"00",X"00",X"00",X"18",X"1C",X"04",X"08",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"40",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"10",X"02",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"41",X"46",X"18",X"01",X"0E",X"18",X"2B",X"14",X"80",X"20",X"C0",X"00",X"68",X"88",X"34",X"04",
		X"03",X"04",X"03",X"05",X"03",X"00",X"00",X"00",X"C8",X"02",X"E4",X"40",X"E0",X"80",X"00",X"00",
		X"00",X"00",X"08",X"04",X"28",X"24",X"0B",X"04",X"00",X"00",X"00",X"00",X"20",X"90",X"44",X"28",
		X"23",X"24",X"03",X"04",X"23",X"24",X"03",X"0C",X"84",X"68",X"80",X"40",X"80",X"40",X"80",X"40",
		X"22",X"01",X"02",X"40",X"41",X"04",X"00",X"01",X"E0",X"10",X"60",X"88",X"3C",X"44",X"9A",X"21",
		X"00",X"02",X"02",X"04",X"02",X"04",X"00",X"00",X"48",X"88",X"94",X"74",X"48",X"30",X"00",X"00",
		X"00",X"00",X"00",X"00",X"40",X"22",X"4D",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"A6",X"08",X"13",X"44",X"48",X"02",X"04",X"21",X"A0",X"20",X"90",X"00",X"C0",X"00",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",
		X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"28",X"00",X"10",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"10",X"00",X"00",X"00",
		X"00",X"18",X"38",X"30",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"07",X"07",X"1F",X"1C",X"1C",
		X"70",X"F0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"07",X"07",X"1F",X"1C",X"7C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"02",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"10",X"00",X"00",X"00",
		X"00",X"18",X"38",X"30",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"07",X"07",X"1F",X"1C",X"1C",
		X"70",X"F0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"07",X"07",X"1F",X"1C",X"7C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"02",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"10",X"00",X"00",X"00",
		X"00",X"18",X"38",X"30",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"07",X"07",X"1F",X"1C",X"1C",
		X"70",X"F0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"07",X"07",X"1F",X"1C",X"7C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"02",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"10",X"00",X"00",X"00",
		X"00",X"18",X"38",X"30",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"07",X"07",X"1F",X"1C",X"1C",
		X"70",X"F0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"07",X"07",X"1F",X"1C",X"7C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"02",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"10",X"0E",X"08",X"00",X"30",X"78",X"70",X"04",X"04",X"30",X"18",X"08",X"00",X"06",X"06",
		X"61",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"4E",X"66",X"06",X"86",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"30",X"39",X"3D",X"1F",X"1C",X"00",X"00",X"40",X"80",X"8C",X"DC",X"FE",X"1E",
		X"08",X"04",X"04",X"08",X"08",X"10",X"10",X"10",X"0C",X"08",X"04",X"04",X"02",X"02",X"02",X"02",
		X"0E",X"02",X"00",X"02",X"03",X"03",X"01",X"00",X"00",X"00",X"06",X"02",X"10",X"18",X"C1",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"38",X"3C",X"9E",X"CE",X"7D",X"38",X"30",X"60",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"40",
		X"E0",X"E0",X"D0",X"D0",X"20",X"20",X"10",X"11",X"40",X"20",X"10",X"08",X"3E",X"5F",X"07",X"00",
		X"20",X"20",X"0C",X"18",X"10",X"00",X"60",X"60",X"08",X"08",X"70",X"10",X"00",X"0C",X"1E",X"0E",
		X"72",X"66",X"60",X"61",X"00",X"00",X"00",X"00",X"86",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"01",X"31",X"3B",X"7F",X"78",X"00",X"00",X"00",X"0C",X"9C",X"BC",X"FC",X"38",
		X"30",X"10",X"20",X"20",X"40",X"40",X"40",X"40",X"10",X"20",X"20",X"10",X"10",X"08",X"08",X"08",
		X"00",X"00",X"60",X"40",X"08",X"19",X"83",X"03",X"70",X"40",X"00",X"40",X"C0",X"C0",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"02",X"1C",X"8C",X"79",X"73",X"BE",X"1C",X"0C",X"06",
		X"02",X"04",X"08",X"10",X"7C",X"FA",X"E0",X"00",X"07",X"07",X"0B",X"0B",X"04",X"04",X"08",X"08",
		X"8C",X"08",X"DD",X"CB",X"0A",X"76",X"28",X"05",X"CD",X"E7",X"31",X"28",X"0F",X"01",X"04",X"00",
		X"21",X"11",X"39",X"11",X"15",X"39",X"ED",X"B0",X"DD",X"CB",X"09",X"C6",X"DD",X"CB",X"0E",X"5E",
		X"20",X"C7",X"CD",X"F9",X"18",X"28",X"C5",X"18",X"62",X"DD",X"CB",X"0E",X"E6",X"CD",X"49",X"1F",
		X"DA",X"F6",X"11",X"EF",X"3A",X"CA",X"DD",X"11",X"CD",X"0D",X"19",X"0E",X"01",X"CD",X"C0",X"2D",
		X"0E",X"13",X"DD",X"CB",X"0F",X"56",X"20",X"1E",X"21",X"FB",X"0C",X"CD",X"30",X"00",X"38",X"14",
		X"DD",X"CB",X"09",X"D6",X"CD",X"0D",X"19",X"0E",X"00",X"CD",X"D8",X"18",X"0E",X"82",X"CD",X"C0",
		X"2D",X"C3",X"8C",X"08",X"0E",X"07",X"CD",X"73",X"24",X"2E",X"2D",X"41",X"2B",X"DD",X"CB",X"0F",
		X"56",X"28",X"08",X"21",X"FB",X"0C",X"CD",X"30",X"00",X"28",X"D5",X"0E",X"11",X"CD",X"73",X"19",
		X"18",X"15",X"DD",X"CB",X"0E",X"66",X"20",X"0F",X"CD",X"F9",X"18",X"16",X"E1",X"CD",X"83",X"1C",
		X"DD",X"CB",X"09",X"D6",X"C3",X"1D",X"12",X"0E",X"01",X"CD",X"C0",X"2D",X"16",X"E2",X"CD",X"83",
		X"1C",X"DD",X"CB",X"09",X"F6",X"DD",X"CB",X"09",X"D6",X"C3",X"1C",X"10",X"2A",X"37",X"39",X"DD",
		X"CB",X"76",X"66",X"C2",X"2C",X"12",X"E5",X"CD",X"E5",X"04",X"E1",X"22",X"37",X"39",X"DD",X"CB",
		X"0A",X"6E",X"20",X"E1",X"DD",X"36",X"0C",X"07",X"DD",X"CB",X"0A",X"76",X"28",X"05",X"0E",X"6B",
		X"CD",X"56",X"2B",X"0E",X"6D",X"CD",X"56",X"2B",X"0E",X"02",X"CD",X"59",X"1A",X"CD",X"B8",X"34",
		X"CD",X"E3",X"18",X"28",X"C0",X"EF",X"2C",X"28",X"14",X"CD",X"F1",X"34",X"CD",X"9E",X"33",X"CD",
		X"E3",X"18",X"28",X"B1",X"EF",X"2C",X"38",X"F1",X"CD",X"E3",X"18",X"38",X"E8",X"CD",X"8F",X"31",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7C",X"7C",X"00",X"00",X"00",X"00",X"00",X"00",X"7C",X"7C",X"7C",X"00",X"00",X"00",X"00",X"00",
		X"7C",X"7C",X"7C",X"7C",X"00",X"00",X"00",X"00",X"7C",X"7C",X"7C",X"7C",X"7C",X"00",X"00",X"00",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"00",X"00",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"00",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"CB",X"0A",X"5E",X"20",X"05",X"16",X"49",X"CD",
		X"83",X"1C",X"DD",X"7E",X"07",X"CD",X"21",X"00",X"18",X"1F",X"26",X"48",X"4B",X"B3",X"9D",X"CB",
		X"77",X"28",X"3C",X"DD",X"CB",X"08",X"F6",X"DD",X"CB",X"09",X"EE",X"CD",X"49",X"1F",X"28",X"48",
		X"21",X"8F",X"14",X"CD",X"61",X"14",X"28",X"C2",X"21",X"9A",X"14",X"CD",X"61",X"14",X"28",X"BA",
		X"CD",X"49",X"1F",X"28",X"33",X"EF",X"24",X"28",X"25",X"CD",X"22",X"1E",X"28",X"25",X"EF",X"28",
		X"28",X"02",X"37",X"DF",X"CD",X"46",X"13",X"EF",X"29",X"DF",X"CD",X"5E",X"14",X"28",X"9B",X"AF",
		X"C3",X"31",X"22",X"1E",X"08",X"18",X"02",X"1E",X"FF",X"CD",X"15",X"20",X"18",X"EC",X"CD",X"BA",
		X"1F",X"18",X"E7",X"CD",X"0D",X"20",X"18",X"E2",X"DD",X"CB",X"08",X"FE",X"0E",X"02",X"CD",X"73",
		X"24",X"30",X"2F",X"33",X"0B",X"0E",X"11",X"CD",X"73",X"19",X"CD",X"04",X"20",X"18",X"CB",X"DD",
		X"CB",X"08",X"56",X"20",X"1C",X"DD",X"CB",X"08",X"C6",X"DD",X"CB",X"0A",X"5E",X"20",X"12",X"DD",
		X"7E",X"03",X"E6",X"0F",X"20",X"06",X"DD",X"CB",X"09",X"6E",X"28",X"05",X"16",X"29",X"CD",X"83",
		X"1C",X"CD",X"F3",X"1F",X"18",X"A4",X"CD",X"15",X"25",X"18",X"CF",X"CD",X"46",X"13",X"CD",X"3F",
		X"20",X"EF",X"2C",X"38",X"06",X"CD",X"46",X"13",X"CD",X"5C",X"20",X"EF",X"5D",X"DF",X"18",X"8A",
		X"CD",X"49",X"1F",X"DF",X"DD",X"CB",X"08",X"FE",X"0E",X"0A",X"CD",X"73",X"24",X"0A",X"09",X"08",
		X"00",X"07",X"05",X"02",X"07",X"00",X"03",X"0E",X"40",X"B0",X"C8",X"60",X"B0",X"F8",X"0C",X"24",
		X"39",X"05",X"06",X"18",X"63",X"01",X"01",X"01",X"B0",X"F8",X"2E",X"E2",X"30",X"9E",X"80",X"80",
		X"00",X"07",X"05",X"02",X"07",X"00",X"03",X"0E",X"40",X"B0",X"C8",X"60",X"B0",X"F8",X"0C",X"24",
		X"39",X"05",X"06",X"18",X"63",X"01",X"01",X"01",X"B0",X"F8",X"2E",X"E2",X"30",X"9E",X"80",X"80",
		X"00",X"07",X"05",X"02",X"07",X"00",X"03",X"0E",X"40",X"B0",X"C8",X"60",X"B0",X"F8",X"0C",X"24",
		X"39",X"05",X"06",X"18",X"63",X"01",X"01",X"01",X"B0",X"F8",X"2E",X"E2",X"30",X"9E",X"80",X"80",
		X"00",X"00",X"01",X"06",X"3C",X"7C",X"7E",X"7F",X"00",X"38",X"F0",X"00",X"00",X"00",X"F0",X"FC",
		X"1F",X"0F",X"0F",X"0F",X"0C",X"04",X"04",X"00",X"FE",X"FE",X"FE",X"FE",X"3C",X"1E",X"3E",X"00",
		X"00",X"18",X"05",X"3F",X"7E",X"7E",X"7E",X"3D",X"00",X"78",X"F8",X"80",X"00",X"00",X"00",X"F0",
		X"03",X"0F",X"0F",X"0F",X"0C",X"04",X"04",X"00",X"FC",X"FE",X"FE",X"FE",X"3C",X"1E",X"3E",X"00",
		X"00",X"73",X"0F",X"07",X"07",X"0B",X"7C",X"07",X"00",X"CE",X"F0",X"E0",X"E0",X"D0",X"3E",X"E0",
		X"03",X"03",X"07",X"0F",X"3F",X"61",X"01",X"00",X"C0",X"C0",X"E0",X"F0",X"FC",X"86",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"84",X"14",X"48",X"08",X"28",X"88",X"10",X"50",X"8C",X"24",X"08",X"50",X"90",X"08",X"58",X"04",
		X"89",X"22",X"04",X"54",X"4A",X"82",X"26",X"04",X"15",X"22",X"82",X"0A",X"05",X"A1",X"45",X"01",
		X"2C",X"84",X"08",X"28",X"88",X"06",X"2A",X"01",X"90",X"50",X"28",X"08",X"28",X"C8",X"14",X"84",
		X"50",X"10",X"B0",X"10",X"20",X"60",X"A0",X"10",X"4A",X"06",X"94",X"04",X"58",X"28",X"10",X"90",
		X"84",X"20",X"02",X"90",X"4A",X"04",X"91",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DD",X"CB",X"09",X"46",X"CD",X"BF",X"26",X"CD",X"09",X"27",X"DD",X"CB",X"09",X"66",X"CD",X"BF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"40",X"40",X"40",X"40",X"80",X"80",X"80",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"20",X"20",X"20",X"20",
		X"04",X"04",X"04",X"04",X"08",X"08",X"08",X"08",X"20",X"20",X"40",X"40",X"40",X"80",X"80",X"80",
		X"04",X"08",X"08",X"08",X"10",X"10",X"10",X"20",X"00",X"00",X"00",X"00",X"00",X"C0",X"38",X"07",
		X"00",X"00",X"80",X"70",X"0E",X"01",X"00",X"00",X"E0",X"1C",X"03",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"38",X"07",X"00",X"00",X"80",X"70",X"0E",X"01",X"00",X"00",
		X"E0",X"1C",X"03",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"80",X"40",X"20",X"10",X"08",X"04",X"02",X"01",X"80",X"40",X"20",X"10",X"08",X"04",X"02",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"C0",X"30",X"0C",X"03",
		X"C0",X"30",X"0C",X"03",X"00",X"00",X"00",X"00",X"FF",X"FE",X"FC",X"F8",X"F0",X"F8",X"FC",X"FF",
		X"80",X"C0",X"E0",X"F0",X"F8",X"FC",X"FE",X"FF",X"01",X"01",X"01",X"02",X"02",X"02",X"04",X"04",
		X"E0",X"1C",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"70",X"0E",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"38",X"07",X"4F",X"41",X"79",X"A7",X"28",X"EF",X"3E",X"20",
		X"77",X"23",X"10",X"FC",X"C9",X"3A",X"06",X"00",X"5F",X"C6",X"10",X"CD",X"D0",X"26",X"3A",X"07",
		X"00",X"93",X"4F",X"11",X"18",X"39",X"E5",X"21",X"13",X"39",X"CD",X"EA",X"27",X"E1",X"A7",X"C8",
		X"4F",X"06",X"00",X"EB",X"ED",X"B0",X"EB",X"C9",X"11",X"17",X"39",X"E5",X"0E",X"04",X"21",X"15",
		X"39",X"CD",X"EA",X"27",X"E1",X"18",X"02",X"3E",X"22",X"4F",X"E6",X"1F",X"C3",X"07",X"01",X"2A",
		X"47",X"39",X"3E",X"84",X"5E",X"BB",X"C8",X"23",X"56",X"ED",X"53",X"11",X"39",X"23",X"22",X"47",
		X"39",X"21",X"7F",X"39",X"3E",X"09",X"11",X"01",X"28",X"CD",X"FF",X"26",X"3A",X"11",X"39",X"57",
		X"3E",X"E1",X"CD",X"1A",X"27",X"36",X"20",X"23",X"E5",X"11",X"0E",X"00",X"21",X"0A",X"28",X"3A",
		X"11",X"39",X"D6",X"3F",X"28",X"15",X"47",X"19",X"7E",X"FE",X"04",X"28",X"07",X"A7",X"20",X"09",
		X"05",X"23",X"18",X"F4",X"21",X"43",X"29",X"18",X"02",X"10",X"EC",X"7B",X"EB",X"E1",X"CD",X"FF",
		X"26",X"E5",X"21",X"07",X"00",X"7E",X"2B",X"96",X"4F",X"2B",X"2B",X"11",X"40",X"39",X"3A",X"12",
		X"39",X"A7",X"ED",X"52",X"EB",X"06",X"04",X"BE",X"28",X"14",X"38",X"11",X"23",X"10",X"F8",X"2B",
		X"96",X"19",X"2B",X"91",X"28",X"03",X"30",X"FB",X"81",X"1E",X"23",X"18",X"05",X"2B",X"96",X"19",
		X"1E",X"2A",X"86",X"E1",X"CD",X"D7",X"26",X"01",X"0A",X"00",X"B7",X"ED",X"42",X"73",X"23",X"C3",
		X"AE",X"26",X"3A",X"07",X"39",X"A1",X"28",X"0C",X"79",X"FE",X"08",X"0E",X"72",X"28",X"02",X"0E",
		X"44",X"CD",X"56",X"2B",X"3C",X"C9",X"2A",X"17",X"39",X"BF",X"DD",X"CB",X"08",X"56",X"C8",X"AF",
		X"BD",X"20",X"05",X"BC",X"C8",X"3C",X"BC",X"C8",X"21",X"7F",X"39",X"0E",X"05",X"CD",X"DA",X"26",
		X"CD",X"09",X"27",X"CD",X"E6",X"26",X"C3",X"AE",X"26",X"1A",X"B9",X"30",X"01",X"4F",X"91",X"12",
		X"5E",X"23",X"56",X"79",X"E5",X"69",X"26",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"3C",X"18",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"03",X"4C",X"30",X"20",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"20",X"20",X"70",X"CB",X"84",X"88",X"50",X"60",X"10",X"20",
		X"7E",X"81",X"00",X"00",X"00",X"42",X"C3",X"E7",X"0E",X"D3",X"21",X"11",X"0A",X"06",X"08",X"C7",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"20",X"20",X"E0",X"10",X"08",X"07",X"00",X"10",X"18",X"1D",X"1F",X"1F",X"1F",X"FF",X"7F",
		X"27",X"4F",X"CF",X"EF",X"F7",X"F0",X"FC",X"FF",X"E7",X"E7",X"C3",X"C3",X"99",X"3C",X"3C",X"18",
		X"E7",X"F3",X"F3",X"F7",X"EF",X"0F",X"3F",X"FF",X"F0",X"F8",X"F8",X"FC",X"FE",X"FE",X"FE",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"2C",X"7E",X"4F",X"3C",X"C8",X"E5",X"CD",X"56",X"2B",X"E1",X"23",X"18",X"F4",X"CD",X"4E",X"1A",
		X"2A",X"6F",X"39",X"EB",X"CD",X"AE",X"2D",X"C4",X"60",X"2D",X"3E",X"C0",X"CD",X"E5",X"33",X"11",
		X"AF",X"3B",X"18",X"63",X"CD",X"7C",X"2D",X"2A",X"73",X"39",X"73",X"23",X"72",X"C9",X"2A",X"9C",
		X"37",X"3E",X"67",X"CD",X"E0",X"33",X"2A",X"C0",X"37",X"3E",X"69",X"CD",X"E0",X"33",X"2A",X"61",
		X"39",X"3E",X"6D",X"CD",X"E0",X"33",X"CD",X"7C",X"2D",X"ED",X"53",X"61",X"39",X"C9",X"ED",X"5B",
		X"6F",X"39",X"2A",X"61",X"39",X"CD",X"60",X"2D",X"3E",X"CD",X"CD",X"E5",X"33",X"22",X"61",X"39",
		X"3E",X"C7",X"CD",X"E5",X"33",X"EB",X"3E",X"C9",X"CD",X"E5",X"33",X"18",X"1A",X"18",X"48",X"FD",
		X"6E",X"02",X"FD",X"66",X"03",X"2B",X"22",X"5F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
