library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity pooyan_char_grphx2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of pooyan_char_grphx2 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"30",X"70",X"C0",X"80",X"80",X"70",X"30",X"00",X"80",X"C0",X"20",X"20",X"60",X"C0",X"80",X"00",
		X"00",X"00",X"F0",X"F0",X"40",X"00",X"00",X"00",X"20",X"20",X"E0",X"E0",X"20",X"20",X"00",X"00",
		X"60",X"F0",X"B0",X"90",X"90",X"C0",X"40",X"00",X"20",X"20",X"A0",X"A0",X"E0",X"E0",X"60",X"00",
		X"80",X"D0",X"F0",X"B0",X"90",X"80",X"00",X"00",X"C0",X"E0",X"20",X"20",X"20",X"60",X"40",X"00",
		X"00",X"F0",X"F0",X"C0",X"60",X"30",X"10",X"00",X"80",X"E0",X"E0",X"80",X"80",X"80",X"80",X"00",
		X"10",X"B0",X"A0",X"A0",X"A0",X"E0",X"E0",X"00",X"C0",X"E0",X"20",X"20",X"20",X"60",X"40",X"00",
		X"00",X"90",X"90",X"90",X"D0",X"70",X"30",X"00",X"C0",X"E0",X"20",X"20",X"20",X"E0",X"C0",X"00",
		X"C0",X"E0",X"B0",X"90",X"80",X"C0",X"C0",X"00",X"00",X"00",X"00",X"E0",X"E0",X"00",X"00",X"00",
		X"00",X"60",X"90",X"90",X"B0",X"F0",X"60",X"00",X"C0",X"E0",X"A0",X"20",X"20",X"20",X"C0",X"00",
		X"70",X"F0",X"90",X"90",X"90",X"F0",X"60",X"00",X"80",X"C0",X"60",X"20",X"20",X"20",X"00",X"00",
		X"30",X"40",X"80",X"A0",X"A0",X"90",X"40",X"30",X"C0",X"20",X"10",X"50",X"50",X"90",X"20",X"C0",
		X"00",X"00",X"C0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"30",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"30",X"30",X"10",X"00",X"00",X"10",X"10",X"70",X"F0",X"E0",X"C0",X"00",
		X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"70",X"C0",X"80",X"C0",X"70",X"30",X"00",X"E0",X"E0",X"80",X"80",X"80",X"E0",X"E0",X"00",
		X"60",X"F0",X"90",X"90",X"90",X"F0",X"F0",X"00",X"C0",X"E0",X"20",X"20",X"20",X"E0",X"E0",X"00",
		X"40",X"C0",X"80",X"80",X"C0",X"70",X"30",X"00",X"40",X"60",X"20",X"20",X"60",X"C0",X"80",X"00",
		X"30",X"70",X"C0",X"80",X"80",X"F0",X"F0",X"00",X"80",X"C0",X"60",X"20",X"20",X"E0",X"E0",X"00",
		X"80",X"90",X"90",X"90",X"F0",X"F0",X"00",X"00",X"20",X"20",X"20",X"20",X"E0",X"E0",X"00",X"00",
		X"80",X"90",X"90",X"90",X"90",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"00",
		X"90",X"90",X"90",X"90",X"C0",X"70",X"30",X"00",X"E0",X"E0",X"20",X"20",X"60",X"C0",X"80",X"00",
		X"F0",X"F0",X"10",X"10",X"10",X"F0",X"F0",X"00",X"E0",X"E0",X"00",X"00",X"00",X"E0",X"E0",X"00",
		X"80",X"80",X"F0",X"F0",X"80",X"80",X"00",X"00",X"20",X"20",X"E0",X"E0",X"20",X"20",X"00",X"00",
		X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",X"20",X"20",X"20",X"60",X"40",X"00",
		X"80",X"C0",X"60",X"30",X"10",X"F0",X"F0",X"00",X"20",X"60",X"E0",X"C0",X"80",X"E0",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"20",X"20",X"20",X"20",X"E0",X"E0",X"00",X"00",
		X"F0",X"F0",X"70",X"30",X"70",X"F0",X"F0",X"00",X"E0",X"E0",X"00",X"80",X"00",X"E0",X"E0",X"00",
		X"F0",X"F0",X"10",X"30",X"70",X"F0",X"F0",X"00",X"E0",X"E0",X"C0",X"80",X"00",X"E0",X"E0",X"00",
		X"70",X"F0",X"80",X"80",X"80",X"F0",X"70",X"00",X"C0",X"E0",X"20",X"20",X"20",X"E0",X"C0",X"00",
		X"70",X"F0",X"80",X"80",X"80",X"F0",X"F0",X"00",X"00",X"80",X"80",X"80",X"80",X"E0",X"E0",X"00",
		X"70",X"F0",X"80",X"80",X"80",X"F0",X"70",X"00",X"A0",X"C0",X"E0",X"A0",X"60",X"E0",X"C0",X"00",
		X"70",X"F0",X"90",X"80",X"80",X"F0",X"F0",X"00",X"20",X"60",X"E0",X"C0",X"80",X"E0",X"E0",X"00",
		X"00",X"50",X"D0",X"90",X"90",X"F0",X"60",X"00",X"C0",X"E0",X"20",X"20",X"20",X"60",X"40",X"00",
		X"80",X"80",X"F0",X"F0",X"80",X"80",X"00",X"00",X"00",X"00",X"E0",X"E0",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"00",X"00",X"00",X"F0",X"F0",X"00",X"C0",X"E0",X"20",X"20",X"20",X"E0",X"C0",X"00",
		X"F0",X"F0",X"10",X"00",X"10",X"F0",X"F0",X"00",X"00",X"80",X"C0",X"E0",X"C0",X"80",X"00",X"00",
		X"F0",X"F0",X"10",X"30",X"10",X"F0",X"F0",X"00",X"E0",X"E0",X"C0",X"80",X"C0",X"E0",X"E0",X"00",
		X"C0",X"E0",X"70",X"30",X"70",X"E0",X"C0",X"00",X"60",X"E0",X"C0",X"80",X"C0",X"E0",X"60",X"00",
		X"E0",X"F0",X"10",X"10",X"F0",X"E0",X"00",X"00",X"00",X"00",X"E0",X"E0",X"00",X"00",X"00",X"00",
		X"C0",X"E0",X"F0",X"B0",X"90",X"80",X"80",X"00",X"20",X"20",X"20",X"A0",X"E0",X"E0",X"60",X"00",
		X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"60",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"30",X"34",X"C3",X"96",
		X"07",X"87",X"4A",X"06",X"06",X"5A",X"2D",X"07",X"00",X"33",X"00",X"00",X"33",X"00",X"00",X"11",
		X"12",X"12",X"12",X"03",X"00",X"00",X"00",X"00",X"0F",X"0F",X"09",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"FF",X"00",X"00",X"FF",X"00",X"FF",X"33",X"33",X"FF",X"33",X"33",X"FF",X"33",
		X"F0",X"E1",X"B4",X"2D",X"2C",X"59",X"08",X"00",X"87",X"1E",X"0E",X"00",X"00",X"CC",X"33",X"33",
		X"00",X"FF",X"00",X"10",X"BA",X"33",X"11",X"FF",X"33",X"33",X"BB",X"FF",X"F7",X"F3",X"FB",X"FF",
		X"00",X"88",X"F9",X"FF",X"F9",X"F9",X"F9",X"88",X"00",X"33",X"E2",X"E2",X"E2",X"EE",X"E2",X"00",
		X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"F0",X"20",X"20",X"20",X"20",X"20",X"20",X"00",X"F0",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"F0",X"00",X"20",X"20",X"20",X"20",X"20",X"20",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"51",X"11",X"20",X"55",X"00",X"00",X"33",X"FF",X"FF",X"FF",X"FB",X"FE",
		X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"74",X"F7",X"00",X"11",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"50",X"00",X"00",X"00",X"10",X"00",X"10",X"00",X"00",
		X"00",X"60",X"F0",X"F0",X"70",X"F0",X"F0",X"60",X"00",X"00",X"00",X"80",X"C0",X"80",X"00",X"00",
		X"C3",X"0F",X"0F",X"87",X"87",X"87",X"87",X"0F",X"0F",X"0F",X"1E",X"3C",X"1E",X"0F",X"0F",X"0F",
		X"77",X"77",X"77",X"33",X"51",X"00",X"00",X"00",X"FE",X"FE",X"FB",X"FF",X"FF",X"FF",X"33",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"D0",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"5A",X"1E",X"0F",X"2D",X"0F",X"0F",X"0F",X"87",X"E1",X"F0",
		X"0F",X"F0",X"1E",X"C3",X"F0",X"0F",X"1E",X"C3",X"78",X"F0",X"F0",X"78",X"F0",X"0F",X"E1",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"20",X"00",X"00",X"00",X"10",X"00",X"10",X"00",X"00",
		X"00",X"20",X"20",X"20",X"20",X"20",X"20",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"00",
		X"33",X"66",X"33",X"00",X"00",X"10",X"B0",X"E1",X"98",X"DC",X"98",X"00",X"C0",X"D0",X"F0",X"1E",
		X"0E",X"78",X"1E",X"0F",X"0F",X"87",X"87",X"4B",X"00",X"08",X"80",X"4A",X"2C",X"0F",X"0F",X"4B",
		X"1E",X"2D",X"C3",X"3C",X"0F",X"C3",X"F0",X"78",X"87",X"4B",X"0F",X"0F",X"0F",X"78",X"F0",X"87",
		X"0F",X"1E",X"69",X"87",X"0F",X"3C",X"78",X"87",X"69",X"96",X"0F",X"0F",X"0F",X"87",X"0F",X"0F",
		X"3C",X"2D",X"C3",X"0F",X"0F",X"1E",X"E1",X"0F",X"87",X"0F",X"0F",X"3C",X"4B",X"87",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"F0",X"F0",X"87",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"87",X"0F",X"0F",X"0F",
		X"00",X"A5",X"2D",X"1E",X"0F",X"0F",X"87",X"0F",X"00",X"00",X"C0",X"68",X"1E",X"E1",X"69",X"1E",
		X"69",X"69",X"3C",X"03",X"00",X"00",X"FB",X"FB",X"C3",X"0F",X"03",X"00",X"00",X"00",X"FB",X"FB",
		X"00",X"00",X"00",X"00",X"30",X"C3",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"C0",X"2C",X"1E",
		X"00",X"00",X"00",X"00",X"E0",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C3",X"96",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"87",
		X"00",X"10",X"10",X"70",X"70",X"10",X"10",X"00",X"00",X"80",X"80",X"E0",X"E0",X"80",X"80",X"00",
		X"F1",X"FB",X"EE",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"00",X"00",X"00",
		X"0F",X"1E",X"3C",X"78",X"C3",X"1E",X"3C",X"0F",X"3C",X"F0",X"C3",X"0F",X"0F",X"E1",X"F0",X"3C",
		X"3C",X"69",X"C3",X"0F",X"0F",X"1E",X"3C",X"3C",X"0F",X"0F",X"0F",X"0F",X"3C",X"F0",X"E1",X"87",
		X"30",X"30",X"30",X"10",X"10",X"30",X"30",X"30",X"C3",X"E1",X"F0",X"F0",X"E1",X"E1",X"C3",X"C3",
		X"FB",X"FB",X"00",X"00",X"00",X"00",X"00",X"00",X"FB",X"FB",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C3",X"69",X"78",X"3C",X"3C",X"3C",X"1E",X"0F",X"00",X"08",X"84",X"86",X"C2",X"C3",X"E1",X"E1",
		X"C0",X"C0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"80",X"80",X"C0",X"E0",X"E0",
		X"69",X"69",X"3C",X"1E",X"0F",X"1E",X"3C",X"78",X"1E",X"2D",X"96",X"E1",X"B4",X"A5",X"F0",X"96",
		X"00",X"00",X"00",X"11",X"B3",X"32",X"51",X"33",X"00",X"00",X"77",X"FF",X"FF",X"FF",X"FE",X"FD",
		X"0F",X"1E",X"3C",X"78",X"3C",X"3C",X"0F",X"0F",X"87",X"87",X"0F",X"0F",X"87",X"C3",X"C3",X"0F",
		X"0F",X"0F",X"0F",X"3C",X"3C",X"1E",X"0F",X"0F",X"0F",X"0F",X"2D",X"0F",X"87",X"C3",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"1E",X"3C",X"69",X"C3",X"0F",X"0F",X"0F",X"0F",X"87",X"0F",X"0F",X"0F",
		X"3C",X"3C",X"1E",X"1E",X"1E",X"0F",X"0F",X"0F",X"E0",X"E0",X"E0",X"F0",X"E0",X"E0",X"E0",X"F0",
		X"F0",X"78",X"78",X"78",X"78",X"78",X"3C",X"3C",X"C0",X"C0",X"C0",X"E0",X"C0",X"C0",X"C0",X"C0",
		X"0F",X"3C",X"2D",X"2D",X"2D",X"1E",X"1E",X"0F",X"68",X"68",X"C0",X"C0",X"C0",X"68",X"68",X"68",
		X"C3",X"0F",X"0F",X"2D",X"C3",X"1E",X"0F",X"1E",X"4B",X"0F",X"D2",X"D2",X"B4",X"3C",X"69",X"C3",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"78",X"3C",X"68",X"80",X"00",X"3C",X"F0",X"E1",X"C3",X"E1",X"61",X"30",X"00",
		X"43",X"43",X"87",X"96",X"96",X"D2",X"30",X"00",X"78",X"F0",X"F0",X"F0",X"E1",X"96",X"2C",X"C0",
		X"0F",X"0F",X"0F",X"0F",X"87",X"C3",X"F0",X"F0",X"78",X"78",X"87",X"87",X"0F",X"0F",X"3C",X"F0",
		X"0F",X"0F",X"0F",X"87",X"C3",X"78",X"3C",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"4B",X"F0",X"B4",
		X"C3",X"96",X"3C",X"B4",X"69",X"0F",X"B4",X"50",X"96",X"A4",X"A4",X"B4",X"B4",X"E0",X"C0",X"80",
		X"F0",X"F0",X"D2",X"1E",X"3C",X"69",X"87",X"C3",X"96",X"D2",X"D2",X"B4",X"B4",X"3C",X"1E",X"1E",
		X"4B",X"4B",X"4B",X"4B",X"87",X"0F",X"0F",X"87",X"0F",X"0F",X"0F",X"0F",X"0F",X"C3",X"E1",X"3C",
		X"48",X"3C",X"B4",X"0E",X"4A",X"1F",X"1E",X"3C",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"33",X"33",X"CC",X"00",X"00",X"00",X"00",X"00",
		X"B4",X"0E",X"4A",X"78",X"3C",X"3C",X"2C",X"1E",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"10",X"30",X"70",X"90",X"10",X"10",X"10",X"10",X"80",X"C0",X"E0",X"90",X"80",X"80",X"80",X"80",
		X"E0",X"7B",X"B4",X"3C",X"1E",X"1E",X"2D",X"1E",X"00",X"FF",X"00",X"00",X"00",X"F7",X"80",X"C0",
		X"00",X"00",X"22",X"55",X"20",X"55",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"3C",X"C3",
		X"0F",X"96",X"60",X"00",X"00",X"00",X"00",X"00",X"E1",X"0F",X"E1",X"21",X"10",X"00",X"00",X"00",
		X"50",X"11",X"31",X"00",X"00",X"00",X"22",X"66",X"F0",X"F8",X"77",X"22",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"F0",X"F0",X"F0",X"F0",X"3C",X"3C",X"0F",X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"69",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"87",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"03",X"03",X"03",X"03",X"03",X"03",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"11",X"11",X"99",X"DD",X"DD",X"FF",X"F3",X"FF",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"00",X"07",X"0F",X"1E",X"78",X"F0",X"F0",X"F0",X"00",X"0E",X"0F",X"C3",X"F0",X"F0",X"F0",X"F0",
		X"70",X"00",X"00",X"08",X"0F",X"E1",X"F0",X"F0",X"CF",X"09",X"01",X"5C",X"CD",X"FE",X"6F",X"96",
		X"0F",X"0F",X"07",X"03",X"07",X"0F",X"0F",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"08",X"0E",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0C",
		X"0E",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"0C",X"0C",X"08",X"0C",X"0E",X"0E",
		X"08",X"0C",X"0C",X"08",X"0E",X"0F",X"0F",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"01",X"21",X"00",X"00",X"0C",X"0F",X"0F",X"0F",X"0F",X"6F",
		X"00",X"01",X"01",X"07",X"0F",X"3C",X"3C",X"78",X"3C",X"3C",X"78",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"03",X"12",X"16",X"34",X"34",
		X"08",X"0C",X"0C",X"0E",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"06",X"0E",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0E",X"0F",X"0F",X"0F",X"0F",X"0E",X"0D",X"04",X"00",X"08",X"0E",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0E",X"0F",X"0F",X"0F",X"0F",X"0F",X"3C",X"F0",X"00",X"0C",X"0F",X"0F",X"0F",X"78",X"F0",X"F0",
		X"00",X"00",X"08",X"0F",X"0F",X"E1",X"F0",X"F0",X"00",X"00",X"0F",X"0F",X"0F",X"78",X"F0",X"F0",
		X"3C",X"1E",X"0F",X"0F",X"1E",X"0F",X"0F",X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"78",X"78",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"69",X"0F",X"0F",X"0F",X"F0",X"F0",X"F0",X"87",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"C3",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"0F",X"87",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"0F",X"0F",X"1E",X"F0",X"F0",X"F0",X"F0",X"0F",X"0F",X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"87",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"3C",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"C3",X"F0",X"F0",X"F0",X"0F",X"0F",X"0F",X"3C",X"F0",X"F0",X"F0",X"F0",
		X"E1",X"C3",X"87",X"87",X"0F",X"0F",X"0F",X"1E",X"78",X"3C",X"F0",X"78",X"78",X"F0",X"E1",X"C3",
		X"00",X"01",X"0D",X"0F",X"0F",X"E1",X"E1",X"96",X"0E",X"0F",X"0F",X"3C",X"1E",X"3C",X"78",X"F0",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0E",X"0F",X"0F",X"0F",X"0E",X"0F",X"0F",X"0E",
		X"0F",X"0F",X"07",X"03",X"07",X"07",X"0F",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"C3",X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"1E",X"1E",X"3C",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"E1",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"78",X"0F",X"0F",X"0F",X"87",X"F0",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0C",X"0E",X"0E",X"0E",X"0E",X"0C",X"08",X"00",X"00",
		X"25",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"E1",X"E1",X"2D",X"16",X"03",X"07",X"12",X"01",
		X"61",X"43",X"06",X"06",X"02",X"04",X"08",X"08",X"68",X"0C",X"08",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"20",X"20",X"20",X"20",X"20",X"F0",X"00",X"20",X"20",X"22",X"20",X"20",X"00",X"00",X"00",
		X"20",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"A8",X"A8",X"AA",X"22",X"64",X"A8",X"F1",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"D0",X"00",
		X"10",X"10",X"98",X"88",X"66",X"EE",X"D8",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"F7",X"55",
		X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"10",X"60",X"00",X"44",X"77",X"BB",X"44",X"44",
		X"80",X"11",X"22",X"CC",X"00",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"11",X"00",X"11",X"D0",X"00",
		X"10",X"10",X"10",X"44",X"00",X"66",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"F7",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"60",X"00",X"00",X"BB",X"00",X"AA",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"33",X"77",X"54",X"76",X"54",X"77",X"33",X"00",X"88",X"C4",X"C8",X"C0",X"C8",X"C4",X"88",
		X"00",X"72",X"31",X"10",X"10",X"10",X"31",X"72",X"00",X"80",X"80",X"60",X"E0",X"60",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"22",X"75",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"FF",X"FF",X"FF",X"76",X"B3",X"11",X"00",X"00",X"FC",X"FD",X"FE",X"FF",X"FF",X"FF",X"77",X"00",
		X"FF",X"AA",X"FF",X"AA",X"AA",X"FF",X"AA",X"FF",X"FF",X"AA",X"FF",X"AA",X"AA",X"FF",X"AA",X"FF",
		X"F3",X"FF",X"F3",X"FF",X"DD",X"DD",X"99",X"11",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",
		X"F5",X"FD",X"F5",X"DD",X"99",X"B9",X"51",X"11",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",
		X"11",X"11",X"51",X"B9",X"99",X"DD",X"F5",X"FD",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0E",X"0C",X"00",
		X"00",X"00",X"00",X"00",X"01",X"12",X"16",X"16",X"00",X"00",X"00",X"07",X"F0",X"F0",X"C3",X"87",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"30",X"70",X"78",X"78",X"1E",
		X"03",X"07",X"87",X"87",X"C3",X"C3",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"E1",
		X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"07",X"00",X"00",X"00",
		X"1E",X"0F",X"0F",X"0F",X"0F",X"0F",X"03",X"00",X"E1",X"0F",X"0F",X"69",X"3C",X"0F",X"0F",X"03",
		X"87",X"87",X"87",X"2D",X"0F",X"1E",X"0F",X"0F",X"A4",X"48",X"08",X"3B",X"08",X"08",X"33",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"30",X"00",X"22",X"CC",X"CC",X"88",X"00",X"00",X"44",X"00",X"11",X"11",X"11",X"44",X"44",X"00",
		X"00",X"00",X"00",X"03",X"16",X"16",X"12",X"07",X"00",X"00",X"0B",X"F0",X"F0",X"C3",X"87",X"4B",
		X"00",X"01",X"07",X"0F",X"0F",X"0F",X"0F",X"07",X"16",X"78",X"F0",X"F0",X"78",X"78",X"0F",X"0F",
		X"0F",X"0F",X"87",X"87",X"C3",X"C3",X"69",X"1E",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"87",
		X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"07",X"01",X"00",X"00",X"00",
		X"0F",X"0F",X"3C",X"1E",X"0F",X"07",X"03",X"00",X"0F",X"0F",X"0F",X"3C",X"A5",X"0F",X"0F",X"07",
		X"00",X"0B",X"B4",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"08",X"84",X"C2",X"68",X"2C",X"2C",X"3C",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"1E",X"1E",X"0F",X"0F",X"0F",X"0F",X"0E",X"0E",
		X"00",X"FF",X"00",X"00",X"51",X"FF",X"20",X"55",X"00",X"FF",X"33",X"FF",X"FF",X"FF",X"FB",X"FE",
		X"00",X"FF",X"98",X"DC",X"CC",X"FF",X"F2",X"FE",X"00",X"FF",X"00",X"60",X"F1",X"FF",X"F1",X"E0",
		X"77",X"FF",X"77",X"33",X"51",X"FF",X"00",X"00",X"FE",X"FF",X"FB",X"FF",X"FF",X"FF",X"33",X"00",
		X"F2",X"FF",X"F2",X"EE",X"CC",X"FF",X"98",X"00",X"E0",X"FF",X"F1",X"F1",X"F1",X"FF",X"00",X"00",
		X"00",X"FF",X"00",X"11",X"B3",X"FF",X"50",X"BB",X"00",X"FF",X"77",X"FF",X"FF",X"FF",X"FC",X"FB",
		X"00",X"FF",X"40",X"A8",X"98",X"FF",X"FC",X"FC",X"00",X"FF",X"22",X"E2",X"E2",X"FF",X"C0",X"C0",
		X"FF",X"FF",X"FF",X"76",X"B3",X"FF",X"00",X"00",X"F8",X"FF",X"FC",X"FF",X"FF",X"FF",X"77",X"00",
		X"FC",X"FF",X"FC",X"DC",X"98",X"FF",X"40",X"00",X"C0",X"FF",X"C0",X"C0",X"E2",X"FF",X"22",X"00",
		X"00",X"D1",X"C0",X"91",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",
		X"00",X"00",X"CC",X"66",X"EE",X"44",X"EE",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"11",X"00",X"33",X"00",X"00",X"00",X"33",X"F3",X"EE",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"EE",X"CC",X"11",X"00",X"00",X"00",X"00",X"00",X"11",X"DD",X"99",X"11",X"40",X"60",X"C0",
		X"00",X"00",X"51",X"C0",X"D1",X"00",X"00",X"00",X"00",X"00",X"44",X"FF",X"77",X"66",X"AA",X"77",
		X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"11",X"11",X"00",X"00",X"00",X"00",X"33",X"33",X"F3",X"EE",X"00",X"00",X"00",X"00",
		X"33",X"BB",X"88",X"88",X"00",X"10",X"30",X"60",X"88",X"CC",X"CC",X"11",X"11",X"00",X"11",X"77",
		X"00",X"90",X"CC",X"22",X"00",X"00",X"00",X"00",X"00",X"F1",X"11",X"31",X"20",X"20",X"20",X"33",
		X"00",X"F0",X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"F8",X"A8",X"31",X"11",X"31",X"20",X"20",
		X"00",X"00",X"00",X"00",X"22",X"EC",X"F0",X"00",X"00",X"00",X"00",X"20",X"20",X"22",X"F2",X"00",
		X"00",X"00",X"00",X"00",X"88",X"20",X"70",X"00",X"EE",X"33",X"31",X"22",X"64",X"64",X"F4",X"00",
		X"00",X"00",X"00",X"11",X"33",X"33",X"FF",X"FF",X"00",X"00",X"00",X"EE",X"FF",X"FF",X"FF",X"FF",
		X"10",X"10",X"10",X"11",X"33",X"BB",X"FF",X"FF",X"00",X"00",X"00",X"88",X"EF",X"EF",X"CC",X"EF",
		X"FF",X"FF",X"77",X"76",X"33",X"11",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"EE",X"FF",X"E0",X"00",
		X"FF",X"FF",X"FF",X"FE",X"98",X"10",X"10",X"10",X"EF",X"CD",X"88",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"11",X"33",X"33",X"FF",X"FF",X"FF",X"00",X"00",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"10",X"10",X"10",X"11",X"33",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"88",X"CC",X"EF",X"EF",X"CC",
		X"FF",X"76",X"77",X"33",X"11",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"70",X"00",X"00",
		X"FF",X"FE",X"77",X"89",X"10",X"10",X"10",X"10",X"EF",X"EF",X"CD",X"88",X"00",X"00",X"00",X"00",
		X"11",X"33",X"33",X"FF",X"FF",X"FF",X"FF",X"77",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"10",X"10",X"BB",X"FF",X"FF",X"FF",X"FF",X"FE",X"00",X"00",X"00",X"88",X"CC",X"EE",X"EF",X"CD",
		X"76",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"70",X"00",X"00",X"00",X"00",
		X"BB",X"33",X"99",X"01",X"10",X"10",X"10",X"10",X"CC",X"EF",X"AB",X"01",X"00",X"00",X"00",X"00",
		X"61",X"43",X"06",X"06",X"02",X"04",X"08",X"08",X"68",X"1D",X"3B",X"11",X"00",X"00",X"00",X"00",
		X"25",X"89",X"CC",X"88",X"00",X"00",X"00",X"00",X"E1",X"E1",X"2D",X"16",X"03",X"07",X"12",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"11",
		X"00",X"00",X"00",X"00",X"00",X"88",X"CC",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"F0",X"20",X"20",X"20",X"20",X"20",X"20",X"00",X"F0",X"20",X"20",X"20",X"00",X"20",X"20",
		X"00",X"F0",X"20",X"20",X"20",X"20",X"20",X"20",X"00",X"F0",X"20",X"20",X"00",X"00",X"00",X"00",
		X"20",X"20",X"20",X"20",X"20",X"20",X"F0",X"00",X"20",X"20",X"00",X"20",X"20",X"20",X"F0",X"00",
		X"20",X"20",X"20",X"20",X"20",X"20",X"F0",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"F1",X"33",
		X"00",X"F0",X"20",X"20",X"20",X"00",X"20",X"20",X"CC",X"74",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"F0",X"20",X"20",X"00",X"00",X"00",X"20",X"00",X"F0",X"33",X"00",X"00",X"00",X"00",X"00",
		X"20",X"20",X"00",X"20",X"20",X"20",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"F0",X"00",
		X"20",X"00",X"00",X"00",X"20",X"20",X"F1",X"33",X"00",X"00",X"00",X"00",X"00",X"33",X"E0",X"00",
		X"44",X"FC",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"CC",X"22",X"00",X"00",X"00",X"00",
		X"00",X"F0",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"88",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"20",X"F0",X"00",X"00",X"00",X"00",X"00",X"22",X"EC",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"33",X"C0",X"00",X"00",X"00",X"00",X"00",X"A8",X"20",X"70",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
