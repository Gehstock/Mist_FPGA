library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_SND_0 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_SND_0 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"F3",X"31",X"00",X"81",X"C3",X"00",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C3",X"F3",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0E",X"10",X"CD",X"EB",X"03",X"0E",X"40",X"CD",X"EB",X"03",X"32",X"FF",X"9F",X"21",X"00",X"80",
		X"01",X"00",X"04",X"36",X"00",X"23",X"0D",X"20",X"FA",X"10",X"F8",X"CD",X"C9",X"01",X"CD",X"F2",
		X"01",X"ED",X"56",X"DD",X"21",X"62",X"02",X"DD",X"21",X"20",X"81",X"CD",X"97",X"01",X"CD",X"A9",
		X"01",X"DD",X"21",X"46",X"81",X"CD",X"97",X"01",X"CD",X"A9",X"01",X"DD",X"21",X"6C",X"81",X"CD",
		X"97",X"01",X"CD",X"A9",X"01",X"DD",X"21",X"92",X"81",X"CD",X"97",X"01",X"CD",X"A9",X"01",X"11",
		X"B8",X"81",X"0E",X"10",X"CD",X"7E",X"01",X"11",X"C7",X"81",X"0E",X"40",X"CD",X"7E",X"01",X"FB",
		X"3A",X"C6",X"81",X"6F",X"3A",X"D5",X"81",X"0F",X"0F",X"47",X"E6",X"0F",X"67",X"78",X"E6",X"C0",
		X"B5",X"6F",X"11",X"00",X"90",X"19",X"77",X"F3",X"CD",X"F2",X"01",X"C3",X"23",X"01",X"2E",X"00",
		X"06",X"0E",X"7D",X"FE",X"0B",X"1A",X"13",X"38",X"06",X"CD",X"19",X"04",X"BC",X"28",X"04",X"67",
		X"CD",X"0A",X"04",X"2C",X"10",X"EC",X"C9",X"DD",X"4E",X"03",X"DD",X"46",X"04",X"DD",X"6E",X"00",
		X"DD",X"66",X"01",X"E5",X"FD",X"E1",X"C3",X"62",X"02",X"DD",X"71",X"03",X"DD",X"70",X"04",X"0A",
		X"B7",X"20",X"0C",X"DD",X"36",X"02",X"00",X"DD",X"36",X"05",X"00",X"DD",X"E5",X"FD",X"E1",X"FD",
		X"E5",X"E1",X"DD",X"75",X"00",X"DD",X"74",X"01",X"C9",X"3E",X"3F",X"32",X"BF",X"81",X"32",X"CE",
		X"81",X"21",X"20",X"81",X"22",X"20",X"81",X"21",X"46",X"81",X"22",X"46",X"81",X"21",X"6C",X"81",
		X"22",X"6C",X"81",X"21",X"92",X"81",X"22",X"92",X"81",X"C9",X"3E",X"0E",X"D3",X"40",X"DB",X"80",
		X"67",X"C9",X"C9",X"F5",X"C5",X"D5",X"E5",X"CD",X"EA",X"01",X"6C",X"7D",X"32",X"D6",X"81",X"FE",
		X"1F",X"38",X"02",X"2E",X"00",X"26",X"00",X"54",X"5D",X"29",X"29",X"19",X"11",X"22",X"04",X"19",
		X"EB",X"1A",X"F5",X"13",X"21",X"22",X"81",X"01",X"26",X"00",X"B7",X"28",X"04",X"09",X"3D",X"20",
		X"FC",X"F1",X"4F",X"1A",X"13",X"47",X"CB",X"BF",X"BE",X"30",X"03",X"C3",X"5A",X"02",X"2B",X"2B",
		X"44",X"75",X"23",X"70",X"23",X"77",X"23",X"1A",X"13",X"47",X"79",X"FE",X"00",X"20",X"06",X"78",
		X"32",X"25",X"81",X"18",X"0D",X"FE",X"01",X"C2",X"52",X"02",X"3A",X"25",X"81",X"A8",X"A0",X"B8",
		X"20",X"08",X"1A",X"13",X"77",X"23",X"1A",X"13",X"77",X"23",X"E1",X"D1",X"C1",X"F1",X"ED",X"56",
		X"FB",X"C9",X"0A",X"03",X"26",X"00",X"87",X"6F",X"11",X"71",X"02",X"19",X"7E",X"23",X"66",X"6F",
		X"E9",X"9F",X"02",X"A3",X"02",X"A4",X"02",X"B0",X"02",X"BD",X"02",X"C7",X"02",X"D3",X"02",X"E0",
		X"02",X"F2",X"02",X"FC",X"02",X"08",X"03",X"17",X"03",X"31",X"03",X"42",X"03",X"58",X"03",X"6C",
		X"03",X"72",X"03",X"8A",X"03",X"9D",X"03",X"AC",X"03",X"C2",X"03",X"D7",X"03",X"E4",X"03",X"01",
		X"00",X"00",X"C9",X"C9",X"0A",X"03",X"6F",X"87",X"9F",X"67",X"09",X"44",X"4D",X"C3",X"62",X"02",
		X"0A",X"03",X"6F",X"0A",X"03",X"67",X"35",X"20",X"EB",X"03",X"C3",X"62",X"02",X"0A",X"03",X"6F",
		X"0A",X"03",X"67",X"5E",X"C3",X"D6",X"02",X"0A",X"03",X"6F",X"0A",X"03",X"67",X"5E",X"23",X"56",
		X"C3",X"E6",X"02",X"0A",X"03",X"5F",X"0A",X"03",X"6F",X"0A",X"03",X"67",X"73",X"C3",X"62",X"02",
		X"0A",X"03",X"5F",X"0A",X"03",X"57",X"0A",X"03",X"6F",X"0A",X"03",X"67",X"73",X"23",X"72",X"C3",
		X"62",X"02",X"0A",X"03",X"6F",X"0A",X"03",X"67",X"5E",X"C3",X"0B",X"03",X"0A",X"03",X"6F",X"0A",
		X"03",X"67",X"5E",X"23",X"56",X"C3",X"1D",X"03",X"0A",X"03",X"5F",X"0A",X"03",X"6F",X"0A",X"03",
		X"67",X"7E",X"83",X"77",X"C3",X"62",X"02",X"0A",X"03",X"5F",X"0A",X"03",X"57",X"0A",X"03",X"6F",
		X"0A",X"03",X"67",X"E5",X"7E",X"23",X"66",X"6F",X"19",X"EB",X"E1",X"73",X"23",X"72",X"C3",X"62",
		X"02",X"0A",X"03",X"5F",X"0A",X"03",X"6F",X"0A",X"03",X"67",X"CB",X"2E",X"1D",X"20",X"FB",X"C3",
		X"62",X"02",X"0A",X"03",X"5F",X"0A",X"03",X"6F",X"0A",X"03",X"67",X"23",X"CB",X"2E",X"2B",X"CB",
		X"1E",X"23",X"1D",X"20",X"F7",X"C3",X"62",X"02",X"0A",X"03",X"5F",X"0A",X"03",X"6F",X"0A",X"03",
		X"67",X"0A",X"77",X"23",X"03",X"1D",X"C2",X"61",X"03",X"C3",X"62",X"02",X"0A",X"03",X"87",X"C3",
		X"5A",X"03",X"CD",X"EB",X"03",X"01",X"B4",X"01",X"21",X"22",X"81",X"AF",X"77",X"23",X"0D",X"20",
		X"FB",X"10",X"F9",X"CD",X"C9",X"01",X"01",X"00",X"00",X"C9",X"0A",X"03",X"57",X"0A",X"03",X"5F",
		X"0A",X"03",X"6F",X"0A",X"03",X"67",X"7E",X"B2",X"A3",X"77",X"C3",X"62",X"02",X"0A",X"03",X"5F",
		X"0A",X"03",X"6F",X"0A",X"03",X"67",X"7E",X"B3",X"77",X"C3",X"62",X"02",X"0A",X"03",X"6F",X"0A",
		X"03",X"67",X"35",X"20",X"09",X"23",X"7E",X"B7",X"20",X"03",X"C3",X"62",X"02",X"35",X"0B",X"0B",
		X"0B",X"C9",X"0A",X"03",X"6F",X"0A",X"03",X"67",X"FD",X"2B",X"FD",X"2B",X"FD",X"71",X"00",X"FD",
		X"70",X"01",X"44",X"4D",X"C3",X"62",X"02",X"FD",X"4E",X"00",X"FD",X"46",X"01",X"FD",X"23",X"FD",
		X"23",X"C3",X"62",X"02",X"DD",X"36",X"02",X"00",X"C3",X"62",X"02",X"CD",X"F2",X"03",X"0E",X"10",
		X"18",X"02",X"0E",X"40",X"06",X"07",X"ED",X"41",X"CB",X"21",X"16",X"00",X"78",X"FE",X"07",X"20",
		X"02",X"16",X"FF",X"ED",X"51",X"CB",X"39",X"10",X"ED",X"C9",X"ED",X"69",X"CB",X"21",X"ED",X"61",
		X"CB",X"39",X"C9",X"0E",X"10",X"18",X"02",X"0E",X"40",X"ED",X"69",X"CB",X"21",X"ED",X"60",X"CB",
		X"39",X"C9",X"00",X"7F",X"00",X"9A",X"04",X"00",X"7E",X"FF",X"ED",X"07",X"00",X"7D",X"FF",X"6B",
		X"0B",X"02",X"7C",X"F0",X"24",X"0C",X"00",X"7B",X"FF",X"88",X"07",X"00",X"78",X"0F",X"EE",X"0B",
		X"00",X"03",X"03",X"DB",X"0C",X"00",X"04",X"0F",X"01",X"05",X"00",X"05",X"0F",X"59",X"06",X"01",
		X"03",X"04",X"9B",X"04",X"01",X"01",X"04",X"C1",X"06",X"00",X"02",X"0F",X"E1",X"06",X"00",X"01",
		X"03",X"47",X"07",X"02",X"40",X"F0",X"06",X"0E",X"00",X"00",X"03",X"97",X"0C",X"00",X"00",X"03",
		X"7C",X"0C",X"00",X"04",X"04",X"CA",X"04",X"02",X"00",X"F0",X"C9",X"05",X"02",X"02",X"30",X"84",
		X"05",X"02",X"02",X"F0",X"A9",X"0D",X"02",X"03",X"F0",X"F5",X"05",X"00",X"06",X"04",X"6F",X"0D",
		X"01",X"1F",X"04",X"73",X"07",X"00",X"1F",X"07",X"7C",X"07",X"10",X"06",X"0F",X"A2",X"81",X"07",
		X"00",X"05",X"BC",X"81",X"06",X"0D",X"C2",X"81",X"06",X"80",X"A0",X"81",X"11",X"24",X"FB",X"BF",
		X"81",X"11",X"30",X"2F",X"C6",X"81",X"01",X"0B",X"F7",X"FF",X"BC",X"81",X"03",X"A0",X"81",X"F6",
		X"16",X"03",X"A2",X"81",X"DA",X"12",X"24",X"BF",X"81",X"00",X"11",X"00",X"3D",X"C6",X"81",X"06",
		X"03",X"A4",X"81",X"11",X"09",X"FE",X"BF",X"81",X"07",X"00",X"02",X"B8",X"81",X"06",X"0F",X"C0",
		X"81",X"06",X"40",X"A6",X"81",X"01",X"03",X"A6",X"81",X"FB",X"16",X"06",X"00",X"C0",X"81",X"06",
		X"80",X"A6",X"81",X"01",X"03",X"A6",X"81",X"FB",X"03",X"A4",X"81",X"D7",X"12",X"09",X"BF",X"81",
		X"00",X"07",X"00",X"00",X"49",X"81",X"11",X"3F",X"FF",X"BF",X"81",X"0E",X"03",X"C3",X"81",X"00",
		X"00",X"00",X"01",X"06",X"00",X"BE",X"81",X"0E",X"03",X"C0",X"81",X"10",X"10",X"10",X"0F",X"03",
		X"B8",X"81",X"E8",X"03",X"DC",X"05",X"D0",X"07",X"07",X"00",X"C0",X"C3",X"81",X"06",X"03",X"C5",
		X"81",X"11",X"3F",X"C0",X"BF",X"81",X"11",X"3F",X"2A",X"C6",X"81",X"06",X"1E",X"9A",X"81",X"06",
		X"10",X"98",X"81",X"01",X"0B",X"03",X"00",X"B8",X"81",X"0B",X"02",X"00",X"BA",X"81",X"0B",X"01",
		X"00",X"BC",X"81",X"03",X"98",X"81",X"EC",X"0A",X"01",X"BE",X"81",X"03",X"9A",X"81",X"E0",X"06",
		X"20",X"98",X"81",X"06",X"08",X"9A",X"81",X"01",X"0B",X"01",X"00",X"B8",X"81",X"0B",X"01",X"00",
		X"BA",X"81",X"03",X"9A",X"81",X"F1",X"0B",X"01",X"00",X"BC",X"81",X"03",X"98",X"81",X"E4",X"12",
		X"3F",X"BF",X"81",X"00",X"11",X"1B",X"FC",X"CE",X"81",X"11",X"0F",X"30",X"D5",X"81",X"0E",X"02",
		X"CF",X"81",X"0F",X"0F",X"0F",X"02",X"C7",X"81",X"80",X"00",X"90",X"00",X"06",X"0F",X"AA",X"81",
		X"06",X"14",X"A8",X"81",X"14",X"B1",X"05",X"16",X"03",X"AA",X"81",X"F4",X"12",X"1B",X"CE",X"81",
		X"00",X"01",X"0B",X"10",X"00",X"C7",X"81",X"0B",X"12",X"00",X"C9",X"81",X"03",X"A8",X"81",X"F1",
		X"0A",X"FF",X"CF",X"81",X"0A",X"FF",X"D0",X"81",X"15",X"0E",X"02",X"D0",X"81",X"0A",X"09",X"11",
		X"3F",X"F9",X"CE",X"81",X"11",X"2F",X"3F",X"D5",X"81",X"0F",X"02",X"C9",X"81",X"80",X"0C",X"00",
		X"0C",X"0A",X"02",X"C9",X"81",X"0A",X"03",X"CB",X"81",X"06",X"06",X"AE",X"81",X"01",X"03",X"AE",
		X"81",X"FB",X"16",X"02",X"EC",X"11",X"3F",X"FF",X"CE",X"81",X"0E",X"03",X"D2",X"81",X"00",X"00",
		X"00",X"01",X"06",X"00",X"CD",X"81",X"0F",X"03",X"C7",X"81",X"44",X"08",X"D0",X"05",X"D0",X"07",
		X"11",X"3F",X"C0",X"CE",X"81",X"11",X"3F",X"15",X"D5",X"81",X"07",X"00",X"40",X"D2",X"81",X"06",
		X"03",X"D4",X"81",X"0E",X"03",X"CF",X"81",X"10",X"10",X"10",X"06",X"40",X"B0",X"81",X"06",X"10",
		X"B2",X"81",X"01",X"0B",X"01",X"00",X"C7",X"81",X"0B",X"03",X"00",X"C9",X"81",X"0A",X"05",X"CD",
		X"81",X"11",X"10",X"1F",X"CD",X"81",X"03",X"B2",X"81",X"E8",X"0B",X"01",X"00",X"CB",X"81",X"16",
		X"03",X"B0",X"81",X"DA",X"12",X"3F",X"CE",X"81",X"00",X"07",X"00",X"00",X"49",X"81",X"11",X"3F",
		X"FF",X"BF",X"81",X"0E",X"03",X"C3",X"81",X"00",X"00",X"00",X"01",X"06",X"08",X"BE",X"81",X"0F",
		X"03",X"B8",X"81",X"44",X"03",X"D0",X"04",X"D0",X"05",X"11",X"3F",X"D8",X"BF",X"81",X"11",X"3F",
		X"2A",X"C6",X"81",X"07",X"00",X"54",X"C3",X"81",X"06",X"03",X"C5",X"81",X"0E",X"03",X"C0",X"81",
		X"10",X"10",X"10",X"06",X"14",X"98",X"81",X"06",X"20",X"9A",X"81",X"01",X"0B",X"21",X"02",X"B8",
		X"81",X"0B",X"37",X"02",X"BA",X"81",X"03",X"9A",X"81",X"F1",X"0A",X"13",X"BE",X"81",X"11",X"0C",
		X"1F",X"BE",X"81",X"0B",X"06",X"00",X"BC",X"81",X"03",X"98",X"81",X"DB",X"12",X"3F",X"BF",X"81",
		X"00",X"11",X"24",X"FB",X"BF",X"81",X"11",X"30",X"1F",X"C6",X"81",X"06",X"0F",X"C2",X"81",X"07",
		X"E0",X"00",X"BC",X"81",X"07",X"30",X"00",X"A2",X"81",X"13",X"A2",X"81",X"12",X"24",X"BF",X"81",
		X"00",X"07",X"00",X"00",X"49",X"81",X"11",X"3F",X"FF",X"BF",X"81",X"0E",X"03",X"C3",X"81",X"00",
		X"00",X"00",X"01",X"06",X"06",X"BE",X"81",X"0F",X"03",X"B8",X"81",X"45",X"04",X"D1",X"04",X"93",
		X"04",X"11",X"3F",X"C0",X"BF",X"81",X"11",X"3F",X"15",X"C6",X"81",X"07",X"00",X"24",X"C3",X"81",
		X"06",X"03",X"C5",X"81",X"0E",X"03",X"C0",X"81",X"10",X"10",X"10",X"06",X"14",X"9A",X"81",X"06",
		X"04",X"98",X"81",X"01",X"01",X"0A",X"01",X"BE",X"81",X"0A",X"37",X"B8",X"81",X"0A",X"5F",X"BA",
		X"81",X"0A",X"23",X"BC",X"81",X"03",X"98",X"81",X"EA",X"0A",X"FD",X"BE",X"81",X"16",X"03",X"9A",
		X"81",X"DD",X"12",X"FF",X"BF",X"81",X"00",X"0F",X"02",X"B8",X"81",X"D0",X"03",X"43",X"04",X"11",
		X"1B",X"FC",X"BF",X"81",X"11",X"0F",X"30",X"C6",X"81",X"0E",X"02",X"C0",X"81",X"09",X"09",X"06",
		X"18",X"98",X"81",X"01",X"0A",X"34",X"B8",X"81",X"0A",X"35",X"BA",X"81",X"03",X"98",X"81",X"F3",
		X"16",X"02",X"D4",X"12",X"24",X"BF",X"81",X"06",X"00",X"C2",X"81",X"00",X"12",X"3F",X"BF",X"81",
		X"0E",X"03",X"C0",X"81",X"00",X"00",X"00",X"00",X"07",X"00",X"00",X"49",X"81",X"07",X"00",X"00",
		X"6F",X"81",X"07",X"00",X"00",X"95",X"81",X"06",X"01",X"BE",X"81",X"11",X"3F",X"EE",X"BF",X"81",
		X"11",X"3F",X"2A",X"C6",X"81",X"0E",X"02",X"C0",X"81",X"0F",X"06",X"07",X"1D",X"01",X"B8",X"81",
		X"06",X"14",X"98",X"81",X"01",X"03",X"98",X"81",X"FB",X"06",X"8F",X"98",X"81",X"01",X"0B",X"01",
		X"00",X"B8",X"81",X"03",X"98",X"81",X"F6",X"07",X"AC",X"01",X"B8",X"81",X"06",X"32",X"98",X"81",
		X"01",X"03",X"98",X"81",X"FB",X"07",X"FE",X"00",X"B8",X"81",X"06",X"40",X"98",X"81",X"01",X"0B",
		X"FE",X"FF",X"B8",X"81",X"03",X"98",X"81",X"F6",X"12",X"1B",X"BF",X"81",X"00",X"07",X"00",X"00",
		X"49",X"81",X"07",X"00",X"00",X"6F",X"81",X"07",X"00",X"00",X"95",X"81",X"12",X"3F",X"CE",X"81");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
