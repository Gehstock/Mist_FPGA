library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity swimmer_big_sprite_tile_bit0 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of swimmer_big_sprite_tile_bit0 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"70",X"FA",X"CF",X"CF",X"CF",X"EF",X"EE",X"00",X"3C",X"7E",X"EE",X"E2",X"E6",X"C6",X"00",
		X"00",X"00",X"00",X"00",X"00",X"38",X"38",X"21",X"00",X"00",X"00",X"00",X"00",X"40",X"A0",X"B0",
		X"30",X"33",X"3F",X"3D",X"31",X"01",X"01",X"03",X"E0",X"E8",X"8F",X"BF",X"FC",X"F8",X"C0",X"F6",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"3A",X"3F",X"37",X"37",X"37",X"3F",X"7F",X"38",X"7C",X"EC",X"CC",X"1C",X"BF",X"FF",X"FB",
		X"00",X"00",X"01",X"02",X"02",X"02",X"04",X"05",X"00",X"C1",X"20",X"10",X"10",X"08",X"C8",X"29",
		X"05",X"05",X"05",X"01",X"00",X"00",X"00",X"00",X"29",X"24",X"14",X"14",X"14",X"14",X"04",X"04",
		X"00",X"FC",X"00",X"00",X"3F",X"00",X"0C",X"CE",X"27",X"5F",X"1D",X"39",X"C2",X"3C",X"00",X"66",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F8",X"FC",X"80",X"00",X"3F",X"00",X"0C",X"CE",X"00",X"C0",X"00",X"00",X"FB",X"00",X"22",X"2F",
		X"00",X"7F",X"00",X"00",X"00",X"00",X"0C",X"CE",X"00",X"8E",X"4E",X"40",X"3F",X"00",X"23",X"EF",
		X"00",X"00",X"01",X"03",X"02",X"07",X"0C",X"06",X"00",X"00",X"80",X"00",X"03",X"04",X"08",X"08",
		X"8E",X"F8",X"00",X"81",X"00",X"23",X"20",X"33",X"08",X"18",X"70",X"F0",X"C0",X"F0",X"00",X"1F",
		X"00",X"00",X"00",X"30",X"30",X"38",X"30",X"30",X"00",X"00",X"00",X"0C",X"0C",X"1C",X"0C",X"0C",
		X"30",X"30",X"30",X"30",X"30",X"1A",X"1F",X"0F",X"0C",X"0C",X"0C",X"0C",X"3C",X"78",X"F8",X"F0",
		X"1F",X"1F",X"3F",X"3F",X"7F",X"73",X"62",X"70",X"B8",X"FC",X"FC",X"FC",X"F8",X"F0",X"70",X"78",
		X"7C",X"1C",X"10",X"18",X"1C",X"00",X"00",X"00",X"38",X"30",X"38",X"38",X"38",X"70",X"60",X"00",
		X"1F",X"3F",X"3F",X"33",X"39",X"39",X"38",X"38",X"FF",X"FF",X"FF",X"77",X"66",X"67",X"67",X"6E",
		X"78",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"78",X"70",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"3F",X"7F",X"7F",X"7E",X"7E",X"60",X"70",X"FB",X"FB",X"F3",X"03",X"00",X"00",X"00",X"00",
		X"3C",X"1C",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"08",X"2C",X"16",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",
		X"F6",X"F0",X"B8",X"C0",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"C0",X"F0",X"FF",
		X"00",X"00",X"00",X"02",X"06",X"16",X"2E",X"2E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"07",X"0F",X"7F",X"FF",X"DD",X"F9",X"FF",X"F0",X"00",X"80",X"CC",X"FC",X"FC",X"DC",X"98",
		X"3F",X"07",X"0F",X"00",X"00",X"00",X"00",X"00",X"9C",X"1C",X"08",X"1C",X"1C",X"1C",X"1C",X"1C",
		X"1F",X"3F",X"3F",X"3F",X"3F",X"3E",X"3C",X"38",X"D8",X"F8",X"FC",X"FC",X"FC",X"CC",X"5C",X"18",
		X"38",X"38",X"38",X"38",X"18",X"3E",X"3E",X"00",X"20",X"38",X"38",X"38",X"38",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"40",
		X"40",X"40",X"C0",X"C0",X"00",X"00",X"00",X"00",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"07",X"0F",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"07",X"03",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"F8",X"FC",X"FC",X"FE",X"FE",X"C6",X"83",X"00",X"00",X"00",X"0F",X"3C",X"00",X"00",X"00",
		X"81",X"81",X"C1",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",
		X"00",X"00",X"7F",X"FF",X"00",X"00",X"00",X"00",X"00",X"7C",X"FF",X"FF",X"03",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"FF",X"00",X"00",X"00",X"03",X"0F",X"7F",X"FE",X"80",X"00",X"00",
		X"00",X"00",X"C0",X"F0",X"F8",X"7C",X"1C",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"E0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"00",X"07",X"0F",X"00",X"1F",X"00",X"00",X"E0",X"00",X"F0",X"F8",X"00",X"F8",
		X"3F",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"BC",X"BC",X"9E",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"1F",X"7F",X"7F",X"FF",X"FE",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"FF",X"7F",X"7F",X"1F",X"07",X"00",X"80",X"C0",X"FC",X"FF",X"FF",X"FF",X"FF",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"07",X"07",X"0F",X"0F",X"0C",X"08",X"E0",X"F8",X"FC",X"FC",X"FE",X"FE",X"7E",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"1F",X"3F",X"80",X"9F",X"00",X"00",X"00",X"00",X"F8",X"FC",X"01",X"F9",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"1F",X"3F",X"3F",X"7F",X"7F",X"63",X"C1",X"00",X"C0",X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"1F",X"00",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"1F",X"1F",X"1F",X"1F",X"DF",X"DF",X"FF",X"FF",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"00",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"1F",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"1F",X"00",X"F1",X"FB",X"FB",X"FF",X"FF",X"FF",X"FF",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"FF",X"7F",X"7F",X"7F",X"20",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3D",X"3D",X"79",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FC",X"FF",X"FF",X"FF",X"80",X"00",X"00",X"00",X"00",X"E0",X"FC",X"FE",X"0F",
		X"87",X"D0",X"DC",X"CE",X"6E",X"06",X"00",X"00",X"E1",X"0B",X"3B",X"73",X"76",X"60",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"1F",X"38",
		X"81",X"81",X"83",X"07",X"00",X"00",X"00",X"00",X"E0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"09",X"7F",X"FF",X"C0",X"00",X"00",X"00",X"00",X"C0",X"F0",X"F8",X"38",X"18",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"F1",X"FB",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"DF",X"DF",X"DF",X"9F",X"9F",X"1F",X"1F",X"FF",X"FF",X"FF",X"FF",X"E0",X"E1",X"C0",X"40",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"0F",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"0F",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"80",X"80",X"00",X"E0",X"F8",X"FE",X"FE",X"FF",X"7F",X"FF",
		X"81",X"83",X"FF",X"FF",X"FF",X"FF",X"FF",X"83",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FC",X"F8",
		X"E1",X"0B",X"3B",X"73",X"76",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"F8",X"FF",X"7F",X"00",X"00",X"00",X"00",X"01",X"00",X"80",X"FC",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"81",X"41",X"02",X"04",X"09",X"00",X"00",X"00",X"E0",X"80",X"00",X"07",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"1F",X"FF",X"F8",X"00",X"00",X"00",X"E0",X"F0",X"E0",X"C0",X"00",X"00",X"00",X"00",
		X"07",X"1F",X"3F",X"3F",X"7F",X"7F",X"7E",X"FC",X"00",X"C0",X"E0",X"E0",X"F0",X"F0",X"30",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"FF",X"DF",X"DF",X"9F",X"9F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"0F",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"83",X"83",X"83",X"83",X"81",X"81",X"80",X"80",X"F0",X"F0",X"F8",X"FF",X"FF",X"FF",X"FF",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"07",X"07",X"0F",X"FF",X"FF",X"FF",X"FF",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"CF",X"CF",X"07",X"03",X"1F",X"BF",X"FF",X"FF",X"FF",X"FF",X"FB",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"BF",X"FF",X"FF",X"FE",X"FE",X"FC",X"F8",X"1F",X"1F",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"1F",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"70",X"FA",X"CF",X"CF",X"CF",X"EF",X"EE",X"00",X"3C",X"7E",X"EE",X"E2",X"E6",X"C6",X"00",
		X"00",X"00",X"00",X"00",X"00",X"38",X"38",X"21",X"00",X"00",X"00",X"00",X"00",X"40",X"A0",X"B0",
		X"30",X"33",X"3F",X"3D",X"31",X"01",X"01",X"03",X"E0",X"E8",X"8F",X"BF",X"FC",X"F8",X"C0",X"F6",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"3A",X"3F",X"37",X"37",X"37",X"3F",X"7F",X"38",X"7C",X"EC",X"CC",X"1C",X"BF",X"FF",X"FB",
		X"00",X"00",X"01",X"02",X"02",X"02",X"04",X"05",X"00",X"C1",X"20",X"10",X"10",X"08",X"C8",X"29",
		X"05",X"05",X"05",X"01",X"00",X"00",X"00",X"00",X"29",X"24",X"14",X"14",X"14",X"14",X"04",X"04",
		X"00",X"FC",X"00",X"00",X"3F",X"00",X"0C",X"CE",X"27",X"5F",X"1D",X"39",X"C2",X"3C",X"00",X"66",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F8",X"FC",X"80",X"00",X"3F",X"00",X"0C",X"CE",X"00",X"C0",X"00",X"00",X"FB",X"00",X"22",X"2F",
		X"00",X"7F",X"00",X"00",X"00",X"00",X"0C",X"CE",X"00",X"8E",X"4E",X"40",X"3F",X"00",X"23",X"EF",
		X"00",X"00",X"01",X"03",X"02",X"07",X"0C",X"06",X"00",X"00",X"80",X"00",X"03",X"04",X"08",X"08",
		X"8E",X"F8",X"00",X"81",X"00",X"23",X"20",X"33",X"08",X"18",X"70",X"F0",X"C0",X"F0",X"00",X"1F",
		X"00",X"00",X"00",X"30",X"30",X"38",X"30",X"30",X"00",X"00",X"00",X"0C",X"0C",X"1C",X"0C",X"0C",
		X"30",X"30",X"30",X"30",X"30",X"1A",X"1F",X"0F",X"0C",X"0C",X"0C",X"0C",X"3C",X"78",X"F8",X"F0",
		X"1F",X"1F",X"3F",X"3F",X"7F",X"73",X"62",X"70",X"B8",X"FC",X"FC",X"FC",X"F8",X"F0",X"70",X"78",
		X"7C",X"1C",X"10",X"18",X"1C",X"00",X"00",X"00",X"38",X"30",X"38",X"38",X"38",X"70",X"60",X"00",
		X"1F",X"3F",X"3F",X"33",X"39",X"39",X"38",X"38",X"FF",X"FF",X"FF",X"77",X"66",X"67",X"67",X"6E",
		X"78",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"78",X"70",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"3F",X"7F",X"7F",X"7E",X"7E",X"60",X"70",X"FB",X"FB",X"F3",X"03",X"00",X"00",X"00",X"00",
		X"3C",X"1C",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"08",X"2C",X"16",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",
		X"F6",X"F0",X"B8",X"C0",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"C0",X"F0",X"FF",
		X"00",X"00",X"00",X"02",X"06",X"16",X"2E",X"2E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"07",X"0F",X"7F",X"FF",X"DD",X"F9",X"FF",X"F0",X"00",X"80",X"CC",X"FC",X"FC",X"DC",X"98",
		X"3F",X"07",X"0F",X"00",X"00",X"00",X"00",X"00",X"9C",X"1C",X"08",X"1C",X"1C",X"1C",X"1C",X"1C",
		X"1F",X"3F",X"3F",X"3F",X"3F",X"3E",X"3C",X"38",X"D8",X"F8",X"FC",X"FC",X"FC",X"CC",X"5C",X"18",
		X"38",X"38",X"38",X"38",X"18",X"3E",X"3E",X"00",X"20",X"38",X"38",X"38",X"38",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"40",
		X"40",X"40",X"C0",X"C0",X"00",X"00",X"00",X"00",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"07",X"0F",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"07",X"03",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"F8",X"FC",X"FC",X"FE",X"FE",X"C6",X"83",X"00",X"00",X"00",X"0F",X"3C",X"00",X"00",X"00",
		X"81",X"81",X"C1",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",
		X"00",X"00",X"7F",X"FF",X"00",X"00",X"00",X"00",X"00",X"7C",X"FF",X"FF",X"03",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"FF",X"00",X"00",X"00",X"03",X"0F",X"7F",X"FE",X"80",X"00",X"00",
		X"00",X"00",X"C0",X"F0",X"F8",X"7C",X"1C",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"E0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"00",X"07",X"0F",X"00",X"1F",X"00",X"00",X"E0",X"00",X"F0",X"F8",X"00",X"F8",
		X"3F",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"BC",X"BC",X"9E",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"1F",X"7F",X"7F",X"FF",X"FE",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"FF",X"7F",X"7F",X"1F",X"07",X"00",X"80",X"C0",X"FC",X"FF",X"FF",X"FF",X"FF",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"07",X"07",X"0F",X"0F",X"0C",X"08",X"E0",X"F8",X"FC",X"FC",X"FE",X"FE",X"7E",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"1F",X"3F",X"80",X"9F",X"00",X"00",X"00",X"00",X"F8",X"FC",X"01",X"F9",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"1F",X"3F",X"3F",X"7F",X"7F",X"63",X"C1",X"00",X"C0",X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"1F",X"00",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"1F",X"1F",X"1F",X"1F",X"DF",X"DF",X"FF",X"FF",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"00",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"1F",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"1F",X"00",X"F1",X"FB",X"FB",X"FF",X"FF",X"FF",X"FF",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"FF",X"7F",X"7F",X"7F",X"20",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3D",X"3D",X"79",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FC",X"FF",X"FF",X"FF",X"80",X"00",X"00",X"00",X"00",X"E0",X"FC",X"FE",X"0F",
		X"87",X"D0",X"DC",X"CE",X"6E",X"06",X"00",X"00",X"E1",X"0B",X"3B",X"73",X"76",X"60",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"1F",X"38",
		X"81",X"81",X"83",X"07",X"00",X"00",X"00",X"00",X"E0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"09",X"7F",X"FF",X"C0",X"00",X"00",X"00",X"00",X"C0",X"F0",X"F8",X"38",X"18",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"F1",X"FB",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"DF",X"DF",X"DF",X"9F",X"9F",X"1F",X"1F",X"FF",X"FF",X"FF",X"FF",X"E0",X"E1",X"C0",X"40",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"0F",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"0F",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"80",X"80",X"00",X"E0",X"F8",X"FE",X"FE",X"FF",X"7F",X"FF",
		X"81",X"83",X"FF",X"FF",X"FF",X"FF",X"FF",X"83",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FC",X"F8",
		X"E1",X"0B",X"3B",X"73",X"76",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"F8",X"FF",X"7F",X"00",X"00",X"00",X"00",X"01",X"00",X"80",X"FC",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"81",X"41",X"02",X"04",X"09",X"00",X"00",X"00",X"E0",X"80",X"00",X"07",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"1F",X"FF",X"F8",X"00",X"00",X"00",X"E0",X"F0",X"E0",X"C0",X"00",X"00",X"00",X"00",
		X"07",X"1F",X"3F",X"3F",X"7F",X"7F",X"7E",X"FC",X"00",X"C0",X"E0",X"E0",X"F0",X"F0",X"30",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"FF",X"DF",X"DF",X"9F",X"9F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"0F",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"83",X"83",X"83",X"83",X"81",X"81",X"80",X"80",X"F0",X"F0",X"F8",X"FF",X"FF",X"FF",X"FF",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"07",X"07",X"0F",X"FF",X"FF",X"FF",X"FF",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"CF",X"CF",X"07",X"03",X"1F",X"BF",X"FF",X"FF",X"FF",X"FF",X"FB",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"BF",X"FF",X"FF",X"FE",X"FE",X"FC",X"F8",X"1F",X"1F",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"1F",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
