library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_OBJ_0 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_OBJ_0 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"38",X"7C",X"C2",X"82",X"86",X"7C",X"38",X"00",X"02",X"02",X"FE",X"FE",X"42",X"02",X"00",X"00",
		X"62",X"F2",X"BA",X"9A",X"9E",X"CE",X"46",X"00",X"8C",X"DE",X"F2",X"B2",X"92",X"86",X"04",X"00",
		X"08",X"FE",X"FE",X"C8",X"68",X"38",X"18",X"00",X"1C",X"BE",X"A2",X"A2",X"A2",X"E6",X"E4",X"00",
		X"0C",X"9E",X"92",X"92",X"D2",X"7E",X"3C",X"00",X"C0",X"E0",X"B0",X"9E",X"8E",X"C0",X"C0",X"00",
		X"0C",X"6E",X"9A",X"92",X"B2",X"F2",X"6C",X"00",X"78",X"FC",X"96",X"92",X"92",X"F2",X"60",X"00",
		X"3C",X"42",X"81",X"A5",X"A5",X"99",X"42",X"3C",X"00",X"00",X"C0",X"F0",X"FB",X"03",X"00",X"00",
		X"0C",X"1E",X"1E",X"1E",X"3C",X"3C",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"06",X"06",X"00",X"00",X"00",X"00",X"00",X"30",X"78",X"7C",X"3E",X"7C",X"78",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"7E",X"C8",X"88",X"C8",X"7E",X"3E",X"00",
		X"6C",X"FE",X"92",X"92",X"92",X"FE",X"FE",X"00",X"44",X"C6",X"82",X"82",X"C6",X"7C",X"38",X"00",
		X"38",X"7C",X"C6",X"82",X"82",X"FE",X"FE",X"00",X"82",X"92",X"92",X"92",X"FE",X"FE",X"00",X"00",
		X"80",X"90",X"90",X"90",X"90",X"FE",X"FE",X"00",X"9E",X"9E",X"92",X"92",X"C6",X"7C",X"38",X"00",
		X"FE",X"FE",X"10",X"10",X"10",X"FE",X"FE",X"00",X"82",X"82",X"FE",X"FE",X"82",X"82",X"00",X"00",
		X"FC",X"FE",X"02",X"02",X"02",X"06",X"04",X"00",X"82",X"C6",X"6E",X"3C",X"18",X"FE",X"FE",X"00",
		X"02",X"02",X"02",X"02",X"FE",X"FE",X"00",X"00",X"FE",X"FE",X"70",X"38",X"70",X"FE",X"FE",X"00",
		X"FE",X"FE",X"1C",X"38",X"70",X"FE",X"FE",X"00",X"7C",X"FE",X"82",X"82",X"82",X"FE",X"7C",X"00",
		X"70",X"F8",X"88",X"88",X"88",X"FE",X"FE",X"00",X"00",X"00",X"81",X"C3",X"7E",X"3C",X"00",X"00",
		X"72",X"F6",X"9E",X"8C",X"88",X"FE",X"FE",X"00",X"0C",X"5E",X"D2",X"92",X"92",X"F6",X"64",X"00",
		X"80",X"80",X"FE",X"FE",X"80",X"80",X"00",X"00",X"FC",X"FE",X"02",X"02",X"02",X"FE",X"FC",X"00",
		X"F0",X"F8",X"1C",X"0E",X"1C",X"F8",X"F0",X"00",X"FE",X"FE",X"1C",X"38",X"1C",X"FE",X"FE",X"00",
		X"C6",X"EE",X"7C",X"38",X"7C",X"EE",X"C6",X"00",X"E0",X"F0",X"1E",X"1E",X"F0",X"E0",X"00",X"00",
		X"10",X"12",X"1C",X"78",X"1C",X"12",X"10",X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"00",
		X"00",X"1D",X"3F",X"7B",X"71",X"73",X"63",X"37",X"00",X"0C",X"08",X"00",X"32",X"7D",X"FD",X"FC",
		X"7D",X"39",X"01",X"31",X"10",X"00",X"00",X"00",X"F8",X"F8",X"F0",X"F4",X"E8",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"03",X"03",X"03",X"03",X"03",X"03",X"FF",X"FF",X"03",X"03",X"03",X"03",X"03",X"03",X"FF",X"FF",
		X"03",X"03",X"03",X"03",X"03",X"03",X"FF",X"FF",X"03",X"03",X"03",X"03",X"03",X"03",X"FF",X"FF",
		X"03",X"03",X"03",X"03",X"03",X"03",X"FF",X"FF",X"03",X"03",X"03",X"03",X"03",X"03",X"FF",X"FF",
		X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"03",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"07",
		X"03",X"00",X"00",X"00",X"00",X"03",X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"03",X"87",X"87",
		X"03",X"00",X"00",X"00",X"00",X"03",X"87",X"87",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"03",X"03",X"03",X"03",X"03",X"03",X"83",X"83",X"03",X"03",X"03",X"03",X"03",X"03",X"83",X"83",
		X"03",X"03",X"03",X"03",X"03",X"03",X"07",X"07",X"03",X"03",X"03",X"03",X"03",X"03",X"07",X"07",
		X"03",X"03",X"03",X"03",X"03",X"03",X"87",X"87",X"03",X"03",X"03",X"03",X"03",X"03",X"87",X"87",
		X"03",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"03",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"03",X"FF",X"FF",
		X"03",X"00",X"00",X"00",X"00",X"03",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"03",X"FF",X"FF",
		X"03",X"00",X"00",X"00",X"00",X"03",X"FF",X"FF",X"03",X"03",X"03",X"03",X"03",X"03",X"FF",X"FF",
		X"03",X"03",X"03",X"03",X"03",X"03",X"FF",X"FF",X"03",X"03",X"03",X"03",X"03",X"03",X"FF",X"FF",
		X"03",X"03",X"03",X"03",X"03",X"03",X"FF",X"FF",X"03",X"03",X"03",X"03",X"03",X"03",X"FF",X"FF",
		X"03",X"03",X"03",X"03",X"03",X"03",X"FF",X"FF",X"03",X"03",X"03",X"03",X"03",X"03",X"FF",X"FF",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"03",X"03",X"03",X"03",X"03",X"03",X"FF",X"FF",X"1C",X"7E",X"DA",X"FA",X"DA",X"7E",X"1C",X"00",
		X"00",X"0F",X"08",X"08",X"0F",X"00",X"0F",X"08",X"00",X"E0",X"20",X"20",X"E0",X"00",X"E0",X"20",
		X"08",X"0F",X"00",X"0F",X"09",X"08",X"0C",X"00",X"20",X"E0",X"00",X"20",X"A0",X"A0",X"E0",X"00",
		X"00",X"0F",X"08",X"08",X"0F",X"00",X"0F",X"08",X"00",X"E0",X"20",X"20",X"E0",X"00",X"E0",X"20",
		X"08",X"0F",X"00",X"00",X"03",X"00",X"0F",X"00",X"20",X"E0",X"00",X"80",X"E0",X"80",X"80",X"00",
		X"00",X"0F",X"08",X"08",X"0F",X"00",X"0F",X"08",X"00",X"E0",X"20",X"20",X"E0",X"00",X"E0",X"20",
		X"08",X"0F",X"00",X"0F",X"09",X"09",X"0F",X"00",X"20",X"E0",X"00",X"E0",X"20",X"20",X"E0",X"00",
		X"0F",X"08",X"08",X"0F",X"00",X"0F",X"08",X"08",X"E0",X"20",X"20",X"E0",X"00",X"E0",X"20",X"20",
		X"0F",X"00",X"09",X"09",X"09",X"0F",X"00",X"0F",X"E0",X"00",X"E0",X"20",X"20",X"E0",X"00",X"E0",
		X"00",X"0F",X"08",X"0F",X"00",X"0F",X"08",X"0F",X"00",X"E0",X"60",X"E0",X"00",X"E0",X"60",X"E0",
		X"00",X"0F",X"0C",X"0C",X"00",X"0F",X"0D",X"0C",X"00",X"20",X"A0",X"E0",X"00",X"E0",X"20",X"20",
		X"00",X"03",X"1F",X"31",X"20",X"23",X"66",X"74",X"00",X"80",X"D0",X"F0",X"80",X"80",X"B8",X"FC",
		X"7F",X"31",X"03",X"33",X"13",X"01",X"00",X"00",X"FC",X"FD",X"FD",X"F2",X"F0",X"E0",X"00",X"E0",
		X"00",X"00",X"04",X"18",X"1C",X"3E",X"77",X"E3",X"00",X"00",X"38",X"08",X"78",X"F8",X"F8",X"F8",
		X"E3",X"E3",X"77",X"3E",X"1C",X"18",X"04",X"00",X"E8",X"F8",X"F8",X"F8",X"78",X"08",X"38",X"00",
		X"00",X"00",X"18",X"34",X"7E",X"7F",X"7F",X"7F",X"00",X"00",X"00",X"00",X"80",X"40",X"80",X"B8",
		X"3C",X"1F",X"01",X"01",X"01",X"00",X"00",X"00",X"FC",X"7D",X"FD",X"F9",X"F8",X"E0",X"00",X"1C",
		X"03",X"09",X"1F",X"1F",X"1F",X"1F",X"0F",X"1D",X"80",X"C0",X"40",X"C0",X"C0",X"E0",X"80",X"40",
		X"6D",X"5D",X"9F",X"9F",X"5F",X"4F",X"60",X"03",X"80",X"C0",X"C0",X"C0",X"C0",X"80",X"00",X"80",
		X"00",X"11",X"27",X"00",X"16",X"0F",X"03",X"03",X"00",X"C0",X"F0",X"F8",X"3C",X"9C",X"CC",X"CC",
		X"01",X"01",X"01",X"03",X"03",X"00",X"00",X"00",X"C8",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0C",X"1E",X"1E",X"3B",X"71",X"00",X"00",X"20",X"00",X"38",X"7E",X"7E",X"FE",
		X"71",X"71",X"3B",X"3E",X"1E",X"0C",X"00",X"00",X"F4",X"FF",X"7F",X"7D",X"38",X"00",X"80",X"00",
		X"00",X"00",X"00",X"0C",X"1E",X"3E",X"39",X"70",X"00",X"00",X"80",X"00",X"38",X"7D",X"7F",X"FF",
		X"70",X"70",X"39",X"3E",X"1E",X"0C",X"00",X"00",X"F4",X"FE",X"7E",X"7E",X"38",X"00",X"20",X"00",
		X"00",X"0F",X"09",X"01",X"11",X"11",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",
		X"10",X"10",X"10",X"10",X"10",X"00",X"00",X"00",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"09",X"0D",X"0D",X"0D",X"0D",X"0D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",
		X"0C",X"0C",X"0C",X"0C",X"0C",X"00",X"00",X"00",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"78",X"78",X"78",X"01",X"00",X"06",X"3E",X"76",X"00",X"00",X"1C",X"1C",X"8C",X"04",X"A4",X"B4",
		X"7E",X"76",X"3E",X"06",X"00",X"03",X"F0",X"00",X"B0",X"B4",X"A4",X"04",X"8C",X"1C",X"00",X"00",
		X"06",X"07",X"07",X"01",X"00",X"0C",X"7C",X"EC",X"00",X"80",X"80",X"80",X"2C",X"46",X"4E",X"D8",
		X"FC",X"EC",X"7C",X"0C",X"00",X"3C",X"00",X"00",X"C0",X"D8",X"4E",X"46",X"2C",X"00",X"00",X"00",
		X"00",X"00",X"38",X"7C",X"7B",X"7F",X"2E",X"1D",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"7C",
		X"1B",X"F4",X"01",X"00",X"0D",X"0F",X"06",X"00",X"40",X"80",X"20",X"B6",X"9E",X"0C",X"00",X"00",
		X"00",X"00",X"38",X"7C",X"7B",X"7F",X"2E",X"1C",X"00",X"00",X"00",X"40",X"60",X"40",X"58",X"5C",
		X"18",X"F9",X"01",X"00",X"00",X"00",X"00",X"00",X"8C",X"98",X"B0",X"40",X"40",X"60",X"E0",X"E0",
		X"00",X"0F",X"0F",X"0F",X"00",X"06",X"3E",X"76",X"00",X"00",X"00",X"00",X"40",X"26",X"2E",X"6A",
		X"7E",X"76",X"3E",X"06",X"00",X"3C",X"00",X"00",X"60",X"6D",X"27",X"23",X"20",X"20",X"00",X"00",
		X"03",X"03",X"03",X"00",X"00",X"06",X"3E",X"76",X"00",X"C0",X"C0",X"C0",X"10",X"13",X"27",X"6D",
		X"7E",X"76",X"3E",X"06",X"00",X"F0",X"00",X"00",X"60",X"6A",X"2E",X"26",X"40",X"80",X"00",X"00",
		X"00",X"0F",X"0F",X"0F",X"00",X"0C",X"7D",X"ED",X"00",X"00",X"00",X"00",X"40",X"26",X"2E",X"6A",
		X"FD",X"ED",X"7D",X"0C",X"00",X"3C",X"00",X"00",X"60",X"6D",X"27",X"23",X"20",X"20",X"00",X"00",
		X"03",X"03",X"03",X"00",X"00",X"0C",X"7D",X"ED",X"00",X"C0",X"C0",X"C0",X"10",X"13",X"27",X"6D",
		X"FD",X"ED",X"7D",X"0C",X"00",X"F0",X"00",X"00",X"60",X"6A",X"2E",X"26",X"40",X"80",X"00",X"00",
		X"00",X"00",X"01",X"03",X"03",X"1F",X"7E",X"D6",X"00",X"C0",X"E0",X"F0",X"30",X"34",X"9C",X"1C",
		X"FE",X"D6",X"7E",X"1F",X"03",X"01",X"00",X"00",X"00",X"18",X"98",X"28",X"C0",X"EC",X"FC",X"30",
		X"00",X"00",X"00",X"03",X"03",X"1F",X"7A",X"DA",X"00",X"30",X"FC",X"EC",X"C0",X"28",X"98",X"18",
		X"FA",X"DA",X"7A",X"1F",X"03",X"03",X"01",X"00",X"00",X"1C",X"9C",X"34",X"30",X"F0",X"E0",X"C0",
		X"00",X"00",X"01",X"03",X"03",X"07",X"07",X"0F",X"00",X"00",X"E0",X"FC",X"FC",X"94",X"10",X"00",
		X"1F",X"7F",X"FF",X"F7",X"DE",X"46",X"02",X"00",X"18",X"FC",X"F0",X"DC",X"0C",X"04",X"00",X"00",
		X"00",X"00",X"01",X"03",X"03",X"07",X"07",X"0F",X"00",X"38",X"F8",X"E8",X"F0",X"FC",X"1C",X"04",
		X"1F",X"7F",X"FF",X"FF",X"DB",X"4A",X"02",X"00",X"00",X"3C",X"BC",X"84",X"C0",X"E0",X"70",X"18",
		X"00",X"00",X"01",X"03",X"03",X"07",X"07",X"0F",X"00",X"00",X"E0",X"FC",X"FC",X"F4",X"90",X"00",
		X"1F",X"7F",X"FF",X"F6",X"DE",X"46",X"02",X"00",X"D8",X"FC",X"F0",X"7C",X"0C",X"04",X"00",X"00",
		X"00",X"00",X"01",X"03",X"03",X"07",X"07",X"0F",X"00",X"38",X"F8",X"E8",X"F0",X"FC",X"9C",X"04",
		X"1F",X"7F",X"FF",X"FF",X"DB",X"4A",X"02",X"00",X"C0",X"FC",X"FC",X"04",X"C0",X"E0",X"70",X"18",
		X"00",X"00",X"00",X"3F",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"F0",X"0C",X"04",X"04",X"FC",
		X"03",X"03",X"03",X"03",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"3F",X"3F",X"00",X"01",X"00",X"00",X"00",X"00",X"FC",X"F4",X"04",X"FC",
		X"03",X"03",X"03",X"03",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"01",X"00",X"39",X"3F",X"47",X"C6",X"8C",X"AF",X"AD",
		X"00",X"01",X"03",X"01",X"00",X"00",X"00",X"00",X"2F",X"AD",X"AF",X"8C",X"C0",X"40",X"01",X"38",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"07",X"06",X"10",X"16",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"1F",X"16",X"10",X"02",X"0E",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"CC",X"10",X"3B",X"3F",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"3F",X"3F",X"3B",X"10",X"CC",X"C0",X"80",
		X"00",X"00",X"00",X"00",X"39",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"C0",X"F0",X"F8",X"FC",
		X"5B",X"0B",X"03",X"01",X"03",X"03",X"01",X"00",X"FE",X"FF",X"BF",X"BC",X"1F",X"1F",X"0D",X"00",
		X"00",X"70",X"78",X"FC",X"BE",X"3F",X"3F",X"2F",X"00",X"00",X"00",X"00",X"00",X"C0",X"F0",X"F8",
		X"0F",X"1B",X"2E",X"1C",X"18",X"30",X"00",X"00",X"FC",X"FC",X"7C",X"1E",X"0F",X"6F",X"61",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"1C",X"3E",X"0E",X"1F",X"3F",X"7F",X"3F",X"FF",
		X"0B",X"00",X"00",X"00",X"03",X"03",X"03",X"00",X"FF",X"1F",X"0F",X"0F",X"9E",X"FE",X"FE",X"3C",
		X"00",X"0F",X"08",X"0F",X"00",X"0F",X"08",X"0F",X"00",X"E0",X"60",X"E0",X"00",X"E0",X"60",X"E0",
		X"00",X"0F",X"08",X"0F",X"00",X"0D",X"0D",X"0F",X"00",X"E0",X"60",X"E0",X"00",X"E0",X"20",X"20",
		X"00",X"1C",X"14",X"22",X"21",X"10",X"10",X"08",X"00",X"00",X"00",X"00",X"00",X"8C",X"5F",X"33",
		X"08",X"10",X"10",X"20",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"14",X"24",X"45",X"82",X"40",X"20",X"00",X"00",X"00",X"80",X"40",X"20",X"18",X"18",
		X"20",X"40",X"80",X"40",X"20",X"00",X"00",X"00",X"30",X"18",X"0C",X"00",X"00",X"00",X"00",X"00",
		X"04",X"0A",X"11",X"00",X"00",X"00",X"00",X"00",X"20",X"50",X"88",X"04",X"02",X"1C",X"20",X"10",
		X"00",X"00",X"01",X"03",X"06",X"04",X"00",X"00",X"08",X"10",X"20",X"C0",X"C0",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
