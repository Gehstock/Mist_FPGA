library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity cpu1_rom is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of cpu1_rom is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"F3",X"ED",X"56",X"C3",X"68",X"00",X"00",X"00",X"87",X"30",X"05",X"24",X"C3",X"10",X"00",X"00",
		X"85",X"6F",X"D0",X"24",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E5",X"D5",X"C5",X"F5",X"CD",X"80",X"00",X"F1",
		X"C1",X"D1",X"E1",X"FB",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"ED",X"45",X"AF",X"32",X"21",X"68",X"31",X"80",X"9A",X"CD",
		X"07",X"1F",X"3E",X"01",X"32",X"21",X"68",X"FB",X"31",X"80",X"9A",X"CD",X"DC",X"1D",X"18",X"F8",
		X"AF",X"32",X"21",X"68",X"32",X"02",X"A0",X"3A",X"9A",X"87",X"A7",X"C2",X"DF",X"02",X"CD",X"4C",
		X"0E",X"CD",X"9F",X"1B",X"3A",X"CF",X"87",X"CB",X"6F",X"CA",X"D0",X"02",X"3A",X"8C",X"89",X"A7",
		X"20",X"02",X"3E",X"05",X"32",X"09",X"84",X"21",X"E5",X"89",X"11",X"EF",X"89",X"06",X"04",X"C5",
		X"CD",X"6F",X"04",X"C1",X"10",X"F9",X"3A",X"E2",X"89",X"E6",X"0F",X"32",X"E2",X"89",X"3A",X"F3",
		X"89",X"FE",X"3C",X"20",X"12",X"AF",X"32",X"F3",X"89",X"21",X"E8",X"89",X"06",X"03",X"37",X"7E",
		X"CE",X"00",X"27",X"77",X"2B",X"10",X"F8",X"21",X"CC",X"87",X"CB",X"4E",X"28",X"05",X"CB",X"56",
		X"CA",X"D0",X"02",X"00",X"3A",X"57",X"86",X"E6",X"03",X"C2",X"9B",X"04",X"21",X"85",X"87",X"11",
		X"00",X"84",X"1A",X"CB",X"4F",X"20",X"06",X"CB",X"56",X"20",X"33",X"18",X"10",X"CB",X"5E",X"20",
		X"33",X"3A",X"81",X"9A",X"FE",X"00",X"CA",X"D0",X"02",X"CB",X"DE",X"18",X"0A",X"3A",X"81",X"9A",
		X"FE",X"00",X"CA",X"D0",X"02",X"CB",X"D6",X"21",X"87",X"04",X"22",X"5A",X"86",X"3E",X"0A",X"32",
		X"5C",X"86",X"21",X"00",X"00",X"22",X"5E",X"86",X"CD",X"51",X"03",X"C3",X"D0",X"02",X"CB",X"46",
		X"20",X"0A",X"18",X"04",X"CB",X"4E",X"20",X"04",X"CB",X"FE",X"18",X"23",X"CB",X"BE",X"3A",X"D5",
		X"85",X"A7",X"C2",X"E5",X"02",X"21",X"00",X"84",X"CB",X"6E",X"CA",X"E5",X"02",X"23",X"CB",X"7E",
		X"28",X"03",X"C3",X"E5",X"02",X"CB",X"6E",X"20",X"06",X"CD",X"51",X"03",X"C3",X"E5",X"02",X"CD",
		X"51",X"12",X"3A",X"01",X"84",X"CB",X"7F",X"C2",X"D0",X"02",X"3A",X"85",X"87",X"CB",X"7F",X"20",
		X"0F",X"3A",X"6F",X"89",X"CB",X"47",X"CA",X"D0",X"02",X"3A",X"57",X"86",X"CB",X"4F",X"28",X"40",
		X"3A",X"5C",X"86",X"A7",X"CA",X"DF",X"02",X"2A",X"5E",X"86",X"7D",X"B4",X"20",X"25",X"2A",X"5A",
		X"86",X"7E",X"32",X"77",X"86",X"23",X"56",X"23",X"5E",X"ED",X"53",X"5E",X"86",X"23",X"22",X"5A",
		X"86",X"3A",X"5C",X"86",X"3D",X"32",X"5C",X"86",X"7B",X"B2",X"20",X"07",X"AF",X"32",X"5C",X"86",
		X"C3",X"DF",X"02",X"2A",X"5E",X"86",X"2B",X"22",X"5E",X"86",X"3A",X"77",X"86",X"32",X"70",X"89",
		X"3A",X"01",X"84",X"CB",X"5F",X"F5",X"C4",X"4E",X"10",X"F1",X"C2",X"9D",X"02",X"3A",X"46",X"86",
		X"CB",X"47",X"C2",X"35",X"02",X"21",X"03",X"84",X"CB",X"56",X"28",X"4F",X"3A",X"85",X"87",X"CB",
		X"7F",X"20",X"07",X"3A",X"57",X"86",X"CB",X"4F",X"28",X"05",X"3A",X"70",X"89",X"18",X"03",X"3A",
		X"B0",X"85",X"4F",X"E6",X"0F",X"FE",X"08",X"CA",X"4E",X"02",X"79",X"CB",X"6F",X"28",X"4F",X"21",
		X"9F",X"87",X"7E",X"E6",X"0F",X"FE",X"00",X"28",X"03",X"35",X"18",X"47",X"21",X"03",X"84",X"CB",
		X"96",X"23",X"CB",X"96",X"AF",X"32",X"41",X"86",X"32",X"A0",X"98",X"32",X"A1",X"98",X"21",X"82",
		X"98",X"06",X"08",X"36",X"00",X"23",X"32",X"30",X"68",X"10",X"F8",X"CD",X"C7",X"10",X"21",X"04",
		X"84",X"CB",X"96",X"18",X"68",X"AF",X"32",X"A0",X"98",X"32",X"A1",X"98",X"3A",X"AE",X"85",X"CB",
		X"4F",X"28",X"04",X"3E",X"1D",X"18",X"02",X"3E",X"1C",X"32",X"22",X"98",X"18",X"4F",X"3E",X"01",
		X"32",X"9F",X"87",X"3A",X"A2",X"98",X"32",X"A0",X"98",X"3A",X"A3",X"98",X"32",X"A1",X"98",X"3A",
		X"22",X"99",X"32",X"20",X"99",X"3E",X"07",X"32",X"21",X"98",X"3A",X"03",X"84",X"CB",X"5F",X"20",
		X"17",X"3A",X"E4",X"87",X"CB",X"4F",X"28",X"08",X"11",X"0E",X"0C",X"CD",X"0E",X"04",X"18",X"1D",
		X"11",X"0A",X"08",X"CD",X"0E",X"04",X"18",X"15",X"3A",X"AE",X"85",X"CB",X"4F",X"28",X"08",X"11",
		X"0F",X"0D",X"CD",X"0E",X"04",X"18",X"06",X"11",X"0B",X"09",X"CD",X"0E",X"04",X"CD",X"0E",X"13",
		X"CD",X"67",X"19",X"3A",X"46",X"86",X"CB",X"47",X"20",X"1C",X"CB",X"4F",X"20",X"18",X"21",X"01",
		X"84",X"CB",X"66",X"20",X"11",X"CD",X"15",X"03",X"3A",X"A2",X"98",X"32",X"80",X"98",X"3A",X"A3",
		X"98",X"32",X"81",X"98",X"18",X"0A",X"AF",X"32",X"80",X"98",X"32",X"81",X"98",X"CD",X"15",X"03",
		X"32",X"30",X"68",X"21",X"56",X"86",X"CB",X"5E",X"28",X"05",X"CB",X"9E",X"CD",X"EA",X"02",X"3E",
		X"01",X"32",X"21",X"68",X"C9",X"CD",X"67",X"19",X"18",X"E6",X"2A",X"DC",X"85",X"E5",X"FD",X"E1",
		X"2A",X"DA",X"85",X"E5",X"DD",X"E1",X"2A",X"D6",X"85",X"ED",X"5B",X"D8",X"85",X"3A",X"AE",X"85",
		X"E6",X"0F",X"CA",X"4D",X"15",X"FE",X"02",X"CA",X"62",X"15",X"FE",X"04",X"CA",X"19",X"15",X"FE",
		X"06",X"CA",X"35",X"15",X"C9",X"3A",X"46",X"86",X"E6",X"03",X"20",X"30",X"3A",X"01",X"84",X"CB",
		X"7F",X"20",X"29",X"3A",X"03",X"84",X"CB",X"57",X"20",X"22",X"3A",X"85",X"87",X"CB",X"7F",X"20",
		X"0C",X"3A",X"57",X"86",X"CB",X"4F",X"20",X"05",X"3A",X"B0",X"85",X"18",X"03",X"3A",X"70",X"89",
		X"E6",X"0F",X"FE",X"08",X"28",X"06",X"3E",X"01",X"32",X"91",X"9A",X"C9",X"AF",X"32",X"91",X"9A",
		X"C9",X"3A",X"00",X"84",X"CB",X"4F",X"20",X"05",X"3A",X"0D",X"84",X"18",X"03",X"3A",X"0E",X"84",
		X"11",X"01",X"00",X"A7",X"28",X"0F",X"1F",X"47",X"30",X"04",X"7A",X"83",X"27",X"57",X"7B",X"87",
		X"27",X"5F",X"78",X"18",X"EE",X"21",X"D5",X"98",X"DD",X"21",X"55",X"98",X"FD",X"21",X"28",X"04",
		X"CD",X"58",X"04",X"DD",X"21",X"54",X"98",X"21",X"D4",X"98",X"7A",X"E6",X"0F",X"5F",X"7A",X"E6",
		X"F0",X"4F",X"16",X"00",X"FE",X"70",X"38",X"04",X"1E",X"08",X"0E",X"60",X"79",X"FD",X"21",X"3A",
		X"04",X"FE",X"00",X"28",X"2C",X"FD",X"21",X"52",X"04",X"FE",X"10",X"28",X"24",X"FD",X"21",X"4C",
		X"04",X"FE",X"20",X"28",X"1C",X"FD",X"21",X"46",X"04",X"FE",X"30",X"28",X"14",X"FD",X"21",X"40",
		X"04",X"FE",X"40",X"28",X"0C",X"FD",X"21",X"34",X"04",X"FE",X"50",X"28",X"04",X"FD",X"21",X"2E",
		X"04",X"CD",X"58",X"04",X"21",X"8A",X"98",X"06",X"09",X"3E",X"61",X"91",X"77",X"23",X"36",X"08",
		X"23",X"C6",X"10",X"10",X"F7",X"21",X"16",X"04",X"19",X"11",X"0A",X"98",X"06",X"09",X"7E",X"12",
		X"23",X"13",X"3E",X"19",X"12",X"13",X"10",X"F6",X"3A",X"00",X"84",X"CB",X"4F",X"C8",X"CB",X"57",
		X"C8",X"21",X"D4",X"98",X"06",X"06",X"3E",X"10",X"86",X"77",X"23",X"10",X"F9",X"C9",X"21",X"20",
		X"98",X"73",X"23",X"23",X"72",X"C9",X"32",X"32",X"32",X"32",X"32",X"32",X"32",X"32",X"32",X"69",
		X"69",X"69",X"69",X"69",X"69",X"69",X"69",X"69",X"00",X"00",X"00",X"18",X"18",X"18",X"D1",X"B1",
		X"91",X"CE",X"CE",X"CE",X"E1",X"C1",X"A1",X"CE",X"CE",X"CE",X"00",X"00",X"00",X"32",X"32",X"32",
		X"00",X"D1",X"B1",X"32",X"CE",X"CE",X"00",X"E1",X"C1",X"32",X"CE",X"CE",X"00",X"00",X"D1",X"32",
		X"32",X"CE",X"00",X"00",X"E1",X"32",X"32",X"CE",X"06",X"03",X"FD",X"7E",X"03",X"DD",X"77",X"00",
		X"FD",X"7E",X"00",X"77",X"23",X"23",X"FD",X"23",X"DD",X"23",X"DD",X"23",X"10",X"EC",X"C9",X"1A",
		X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"47",X"13",X"1A",X"CB",X"27",X"CB",X"27",X"CB",
		X"27",X"CB",X"27",X"B0",X"77",X"2B",X"C9",X"36",X"00",X"01",X"38",X"00",X"1E",X"36",X"00",X"64",
		X"34",X"00",X"E4",X"32",X"00",X"08",X"38",X"01",X"00",X"FF",X"FF",X"21",X"87",X"87",X"36",X"FF",
		X"21",X"57",X"86",X"CB",X"46",X"CA",X"17",X"05",X"CB",X"CE",X"CB",X"76",X"20",X"0A",X"CB",X"F6",
		X"21",X"58",X"86",X"36",X"00",X"C3",X"17",X"05",X"21",X"58",X"86",X"7E",X"E6",X"0F",X"47",X"CB",
		X"66",X"20",X"2B",X"78",X"A7",X"CA",X"26",X"05",X"3D",X"CA",X"A2",X"06",X"3D",X"CA",X"0D",X"07",
		X"3D",X"CA",X"48",X"07",X"3D",X"3D",X"3D",X"CA",X"5D",X"07",X"3D",X"CA",X"85",X"07",X"3D",X"CA",
		X"C0",X"07",X"3D",X"CA",X"5E",X"08",X"3D",X"CA",X"7D",X"08",X"36",X"00",X"18",X"29",X"78",X"A7",
		X"CA",X"82",X"08",X"3D",X"CA",X"B5",X"09",X"3D",X"CA",X"18",X"0A",X"3D",X"CA",X"BC",X"0B",X"3D",
		X"3D",X"3D",X"CA",X"BF",X"0B",X"3D",X"CA",X"C7",X"0B",X"3D",X"CA",X"DC",X"0B",X"3D",X"CA",X"EB",
		X"0B",X"3D",X"CA",X"F3",X"0B",X"36",X"00",X"21",X"57",X"86",X"CB",X"46",X"20",X"02",X"36",X"00",
		X"3E",X"01",X"32",X"21",X"68",X"C9",X"CB",X"E6",X"21",X"80",X"98",X"06",X"80",X"36",X"00",X"23",
		X"10",X"FB",X"21",X"00",X"A0",X"36",X"01",X"23",X"36",X"01",X"23",X"23",X"36",X"00",X"21",X"10",
		X"80",X"11",X"30",X"80",X"06",X"10",X"3E",X"7F",X"77",X"12",X"23",X"13",X"10",X"F8",X"11",X"1B",
		X"80",X"21",X"9C",X"05",X"06",X"06",X"7E",X"12",X"23",X"1B",X"10",X"FA",X"21",X"13",X"80",X"36",
		X"10",X"21",X"40",X"80",X"01",X"80",X"03",X"36",X"7F",X"23",X"0B",X"32",X"30",X"68",X"79",X"B0",
		X"20",X"F5",X"21",X"68",X"86",X"06",X"07",X"36",X"00",X"23",X"10",X"FB",X"21",X"59",X"86",X"36",
		X"01",X"21",X"40",X"98",X"06",X"0A",X"0E",X"86",X"71",X"0C",X"23",X"36",X"0B",X"23",X"10",X"F8",
		X"21",X"40",X"99",X"06",X"14",X"36",X"00",X"23",X"10",X"FB",X"18",X"1A",X"1C",X"2B",X"1E",X"1D",
		X"22",X"2D",X"31",X"10",X"51",X"10",X"71",X"10",X"91",X"10",X"B1",X"10",X"31",X"30",X"51",X"30",
		X"71",X"30",X"91",X"30",X"B1",X"30",X"21",X"A2",X"05",X"11",X"C0",X"98",X"01",X"14",X"00",X"ED",
		X"B0",X"3E",X"F1",X"32",X"80",X"98",X"32",X"A2",X"98",X"32",X"E4",X"98",X"32",X"EC",X"98",X"21",
		X"D4",X"98",X"CD",X"9A",X"06",X"3E",X"10",X"32",X"81",X"98",X"32",X"A3",X"98",X"32",X"E5",X"98",
		X"32",X"ED",X"98",X"21",X"D5",X"98",X"CD",X"9A",X"06",X"3E",X"02",X"32",X"22",X"98",X"21",X"22",
		X"99",X"CD",X"9A",X"06",X"32",X"64",X"99",X"32",X"6C",X"99",X"32",X"6D",X"98",X"AF",X"32",X"23",
		X"98",X"21",X"54",X"99",X"CD",X"9A",X"06",X"3E",X"20",X"32",X"64",X"98",X"3E",X"01",X"32",X"65",
		X"98",X"3E",X"24",X"32",X"6C",X"98",X"3E",X"05",X"32",X"25",X"98",X"32",X"27",X"98",X"32",X"29",
		X"98",X"3E",X"09",X"21",X"55",X"98",X"CD",X"9A",X"06",X"21",X"DD",X"06",X"11",X"8A",X"98",X"01",
		X"18",X"00",X"C5",X"ED",X"B0",X"C1",X"21",X"F5",X"06",X"11",X"0A",X"98",X"ED",X"B0",X"21",X"0A",
		X"99",X"06",X"0C",X"36",X"00",X"23",X"23",X"10",X"FA",X"21",X"54",X"98",X"06",X"04",X"3E",X"48",
		X"77",X"3C",X"23",X"23",X"10",X"FA",X"21",X"F6",X"0B",X"22",X"5A",X"86",X"21",X"48",X"0C",X"22",
		X"5C",X"86",X"21",X"2C",X"0C",X"22",X"5E",X"86",X"21",X"04",X"0C",X"22",X"60",X"86",X"21",X"0E",
		X"0C",X"22",X"62",X"86",X"21",X"18",X"0C",X"22",X"64",X"86",X"21",X"22",X"0C",X"22",X"66",X"86",
		X"21",X"C0",X"83",X"06",X"3F",X"7E",X"FE",X"8C",X"20",X"02",X"36",X"0C",X"23",X"10",X"F6",X"3E",
		X"00",X"32",X"04",X"A0",X"32",X"05",X"A0",X"C3",X"17",X"05",X"06",X"04",X"77",X"23",X"23",X"10",
		X"FB",X"C9",X"CB",X"E6",X"21",X"03",X"A0",X"36",X"01",X"21",X"40",X"80",X"01",X"80",X"03",X"36",
		X"7D",X"7D",X"E6",X"1F",X"FE",X"04",X"30",X"02",X"36",X"8C",X"23",X"0B",X"79",X"B0",X"20",X"EF",
		X"21",X"84",X"80",X"11",X"20",X"00",X"0E",X"08",X"06",X"18",X"E5",X"36",X"7F",X"19",X"10",X"FB",
		X"E1",X"23",X"0D",X"20",X"F3",X"21",X"76",X"86",X"36",X"00",X"C3",X"17",X"05",X"21",X"90",X"41",
		X"90",X"A9",X"90",X"C9",X"90",X"21",X"B0",X"41",X"B0",X"A9",X"B0",X"C9",X"B0",X"21",X"B0",X"89",
		X"B0",X"B9",X"90",X"31",X"90",X"C0",X"1A",X"C1",X"1A",X"C2",X"1B",X"C3",X"1B",X"C4",X"1A",X"C5",
		X"1A",X"C6",X"1B",X"C7",X"1B",X"C8",X"1C",X"CB",X"1A",X"CC",X"1C",X"CD",X"1C",X"CB",X"E6",X"21",
		X"76",X"86",X"36",X"00",X"AF",X"32",X"E4",X"98",X"32",X"E5",X"98",X"32",X"EC",X"98",X"32",X"ED",
		X"98",X"32",X"A2",X"98",X"32",X"A3",X"98",X"32",X"80",X"98",X"32",X"81",X"98",X"21",X"0A",X"98",
		X"11",X"8A",X"98",X"06",X"18",X"3E",X"00",X"0E",X"32",X"71",X"12",X"23",X"13",X"10",X"FA",X"21",
		X"5F",X"80",X"22",X"5A",X"86",X"C3",X"17",X"05",X"CB",X"E6",X"21",X"00",X"99",X"06",X"80",X"36",
		X"00",X"23",X"10",X"FB",X"21",X"00",X"00",X"22",X"5A",X"86",X"C3",X"17",X"05",X"CB",X"E6",X"06",
		X"80",X"21",X"00",X"98",X"11",X"80",X"98",X"DD",X"21",X"00",X"99",X"AF",X"77",X"12",X"DD",X"77",
		X"00",X"23",X"13",X"DD",X"23",X"10",X"F4",X"21",X"00",X"A0",X"AF",X"77",X"23",X"77",X"23",X"77",
		X"23",X"77",X"C3",X"17",X"05",X"CB",X"E6",X"21",X"0D",X"84",X"11",X"A9",X"87",X"7E",X"12",X"4F",
		X"23",X"13",X"7E",X"12",X"79",X"13",X"12",X"21",X"76",X"86",X"36",X"10",X"23",X"36",X"00",X"21",
		X"80",X"87",X"34",X"CB",X"46",X"20",X"05",X"21",X"E3",X"15",X"18",X"03",X"21",X"6D",X"16",X"22",
		X"5A",X"86",X"3E",X"7E",X"32",X"5C",X"86",X"21",X"00",X"00",X"22",X"5E",X"86",X"C3",X"17",X"05",
		X"CB",X"E6",X"21",X"0D",X"84",X"11",X"A9",X"87",X"1A",X"77",X"23",X"13",X"1A",X"77",X"21",X"40",
		X"80",X"01",X"80",X"03",X"36",X"0C",X"23",X"0B",X"79",X"B0",X"20",X"F8",X"21",X"80",X"98",X"06",
		X"80",X"36",X"00",X"23",X"10",X"FB",X"21",X"00",X"98",X"06",X"40",X"36",X"32",X"23",X"36",X"00",
		X"23",X"10",X"F8",X"21",X"C0",X"83",X"06",X"3F",X"7E",X"FE",X"8C",X"20",X"02",X"36",X"0C",X"32",
		X"30",X"68",X"23",X"10",X"F3",X"21",X"A2",X"05",X"11",X"C0",X"98",X"01",X"14",X"00",X"ED",X"B0",
		X"21",X"40",X"98",X"06",X"0A",X"0E",X"86",X"71",X"0C",X"23",X"36",X"0B",X"23",X"10",X"F8",X"21",
		X"40",X"99",X"06",X"14",X"36",X"00",X"23",X"10",X"FB",X"21",X"2B",X"81",X"11",X"20",X"00",X"06",
		X"0E",X"DD",X"21",X"50",X"08",X"DD",X"7E",X"00",X"77",X"DD",X"23",X"19",X"10",X"F7",X"21",X"03",
		X"A0",X"36",X"01",X"21",X"5E",X"86",X"36",X"FF",X"21",X"CC",X"87",X"CB",X"C6",X"C3",X"17",X"05",
		X"7F",X"7F",X"7F",X"7F",X"15",X"7F",X"2D",X"2C",X"1E",X"1B",X"7F",X"7F",X"7F",X"7F",X"CB",X"E6",
		X"3E",X"01",X"2A",X"00",X"A0",X"77",X"23",X"77",X"23",X"23",X"36",X"00",X"21",X"40",X"80",X"01",
		X"80",X"03",X"36",X"7F",X"23",X"0B",X"79",X"B0",X"20",X"F8",X"C3",X"17",X"05",X"CB",X"E6",X"C3",
		X"17",X"05",X"21",X"4E",X"0C",X"3A",X"59",X"86",X"96",X"32",X"59",X"86",X"D2",X"17",X"05",X"3A",
		X"68",X"86",X"A7",X"20",X"27",X"2A",X"5A",X"86",X"7E",X"32",X"6F",X"86",X"23",X"7E",X"23",X"22",
		X"5A",X"86",X"FE",X"09",X"20",X"13",X"32",X"68",X"86",X"3E",X"8C",X"32",X"82",X"80",X"32",X"A2",
		X"80",X"32",X"83",X"80",X"32",X"A3",X"80",X"18",X"03",X"32",X"68",X"86",X"3A",X"68",X"86",X"3D",
		X"32",X"68",X"86",X"CD",X"4F",X"0C",X"3A",X"A2",X"98",X"32",X"80",X"98",X"3A",X"A3",X"98",X"32",
		X"81",X"98",X"FE",X"10",X"20",X"08",X"21",X"80",X"98",X"36",X"00",X"23",X"36",X"00",X"3E",X"38",
		X"32",X"00",X"98",X"3E",X"06",X"32",X"01",X"98",X"3A",X"A3",X"98",X"FE",X"10",X"28",X"03",X"CD",
		X"0E",X"13",X"3A",X"69",X"86",X"A7",X"20",X"10",X"2A",X"5C",X"86",X"7E",X"32",X"70",X"86",X"23",
		X"7E",X"23",X"22",X"5C",X"86",X"32",X"69",X"86",X"3A",X"69",X"86",X"3D",X"32",X"69",X"86",X"CD",
		X"EE",X"0C",X"3A",X"6A",X"86",X"A7",X"20",X"10",X"2A",X"5E",X"86",X"7E",X"32",X"71",X"86",X"23",
		X"7E",X"23",X"22",X"5E",X"86",X"32",X"6A",X"86",X"3A",X"6A",X"86",X"3D",X"32",X"6A",X"86",X"CD",
		X"4D",X"0D",X"3A",X"6B",X"86",X"A7",X"20",X"10",X"2A",X"60",X"86",X"7E",X"32",X"72",X"86",X"23",
		X"7E",X"23",X"22",X"60",X"86",X"32",X"6B",X"86",X"3A",X"6B",X"86",X"3D",X"32",X"6B",X"86",X"CD",
		X"FB",X"0C",X"3A",X"6C",X"86",X"A7",X"20",X"10",X"2A",X"62",X"86",X"7E",X"32",X"73",X"86",X"23",
		X"7E",X"23",X"22",X"62",X"86",X"32",X"6C",X"86",X"3A",X"6C",X"86",X"3D",X"32",X"6C",X"86",X"CD",
		X"08",X"0D",X"3A",X"6D",X"86",X"A7",X"20",X"10",X"2A",X"64",X"86",X"7E",X"32",X"74",X"86",X"23",
		X"7E",X"23",X"22",X"64",X"86",X"32",X"6D",X"86",X"3A",X"6D",X"86",X"3D",X"32",X"6D",X"86",X"CD",
		X"15",X"0D",X"3A",X"6E",X"86",X"A7",X"20",X"10",X"2A",X"66",X"86",X"7E",X"32",X"75",X"86",X"23",
		X"7E",X"23",X"22",X"66",X"86",X"32",X"6E",X"86",X"3A",X"6E",X"86",X"3D",X"32",X"6E",X"86",X"CD",
		X"22",X"0D",X"C3",X"17",X"05",X"21",X"76",X"86",X"34",X"7E",X"FE",X"05",X"30",X"0F",X"F5",X"21",
		X"C1",X"98",X"06",X"0A",X"34",X"34",X"34",X"34",X"23",X"23",X"10",X"F8",X"F1",X"FE",X"05",X"38",
		X"15",X"FE",X"09",X"30",X"11",X"F5",X"21",X"E5",X"98",X"11",X"ED",X"98",X"34",X"34",X"34",X"34",
		X"EB",X"34",X"34",X"34",X"34",X"F1",X"FE",X"09",X"20",X"0A",X"21",X"64",X"98",X"36",X"23",X"21",
		X"6C",X"98",X"36",X"27",X"FE",X"05",X"38",X"13",X"FE",X"37",X"30",X"0F",X"F5",X"21",X"D5",X"98",
		X"06",X"04",X"34",X"34",X"34",X"34",X"23",X"23",X"10",X"F8",X"F1",X"FE",X"72",X"C2",X"FB",X"0D",
		X"21",X"58",X"86",X"36",X"02",X"C3",X"FB",X"0D",X"21",X"76",X"86",X"34",X"CB",X"46",X"CA",X"17",
		X"05",X"2A",X"5A",X"86",X"11",X"3F",X"80",X"A7",X"ED",X"52",X"20",X"02",X"18",X"1B",X"2A",X"5A",
		X"86",X"11",X"F0",X"87",X"1A",X"CB",X"DF",X"12",X"11",X"20",X"00",X"06",X"1C",X"36",X"7F",X"19",
		X"10",X"FB",X"2A",X"5A",X"86",X"2B",X"22",X"5A",X"86",X"21",X"76",X"86",X"7E",X"FE",X"07",X"20",
		X"28",X"AF",X"21",X"D4",X"98",X"06",X"08",X"77",X"23",X"10",X"FC",X"21",X"D4",X"93",X"06",X"08",
		X"77",X"23",X"10",X"FC",X"21",X"72",X"0A",X"11",X"9C",X"81",X"06",X"07",X"CD",X"3B",X"0E",X"C3",
		X"17",X"05",X"BF",X"BE",X"BD",X"BC",X"BB",X"BA",X"B9",X"FE",X"0B",X"20",X"1F",X"21",X"8B",X"0A",
		X"11",X"FA",X"80",X"06",X"11",X"CD",X"3B",X"0E",X"C3",X"17",X"05",X"35",X"1D",X"2D",X"25",X"7F",
		X"28",X"1C",X"26",X"1A",X"27",X"7F",X"12",X"18",X"19",X"11",X"7F",X"38",X"FE",X"15",X"20",X"20",
		X"21",X"AE",X"0A",X"11",X"D5",X"80",X"06",X"12",X"CD",X"3B",X"0E",X"C3",X"17",X"05",X"6B",X"5A",
		X"60",X"72",X"5F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"5A",X"64",X"68",X"68",X"69",
		X"FE",X"23",X"20",X"17",X"21",X"D2",X"0A",X"11",X"6E",X"81",X"06",X"09",X"CD",X"3B",X"0E",X"C3",
		X"17",X"05",X"6B",X"5E",X"6D",X"5C",X"5A",X"6B",X"5A",X"61",X"5C",X"FE",X"61",X"20",X"33",X"21",
		X"F0",X"87",X"CB",X"9E",X"AF",X"32",X"64",X"99",X"3C",X"32",X"65",X"98",X"3C",X"32",X"6D",X"98",
		X"32",X"6C",X"99",X"3E",X"90",X"32",X"E5",X"98",X"32",X"ED",X"98",X"3E",X"B2",X"32",X"EC",X"98",
		X"3E",X"52",X"32",X"E4",X"98",X"3E",X"20",X"32",X"64",X"98",X"3E",X"24",X"32",X"6C",X"98",X"C3",
		X"17",X"05",X"21",X"6D",X"98",X"FE",X"77",X"20",X"05",X"36",X"0C",X"C3",X"17",X"05",X"FE",X"7F",
		X"20",X"05",X"36",X"02",X"C3",X"17",X"05",X"FE",X"87",X"20",X"02",X"18",X"EC",X"FE",X"8F",X"20",
		X"02",X"18",X"EF",X"FE",X"B3",X"20",X"13",X"36",X"02",X"DD",X"21",X"A4",X"98",X"06",X"06",X"DD",
		X"36",X"00",X"00",X"DD",X"23",X"10",X"F8",X"C3",X"17",X"05",X"DD",X"21",X"24",X"98",X"FD",X"21",
		X"A4",X"98",X"11",X"EC",X"98",X"FE",X"97",X"20",X"2D",X"36",X"0C",X"1A",X"D6",X"10",X"FD",X"77",
		X"00",X"D6",X"10",X"FD",X"77",X"02",X"D6",X"10",X"FD",X"77",X"04",X"13",X"1A",X"FD",X"77",X"01",
		X"FD",X"77",X"03",X"FD",X"77",X"05",X"3E",X"2C",X"DD",X"77",X"00",X"3E",X"32",X"DD",X"77",X"02",
		X"DD",X"77",X"04",X"C3",X"17",X"05",X"FE",X"9D",X"20",X"11",X"3E",X"2D",X"DD",X"77",X"00",X"3C",
		X"DD",X"77",X"02",X"3E",X"32",X"DD",X"77",X"04",X"C3",X"17",X"05",X"FE",X"A3",X"20",X"10",X"3E",
		X"2F",X"DD",X"77",X"00",X"3C",X"DD",X"77",X"02",X"3C",X"DD",X"77",X"04",X"C3",X"17",X"05",X"FE",
		X"FF",X"C2",X"17",X"05",X"21",X"58",X"86",X"36",X"03",X"C3",X"17",X"05",X"C3",X"00",X"17",X"21",
		X"58",X"86",X"36",X"07",X"C3",X"17",X"05",X"3A",X"76",X"86",X"FE",X"80",X"CA",X"5F",X"01",X"FE",
		X"90",X"C2",X"17",X"05",X"21",X"58",X"86",X"36",X"08",X"C3",X"5F",X"07",X"21",X"5E",X"86",X"35",
		X"C2",X"17",X"05",X"21",X"58",X"86",X"36",X"09",X"C3",X"17",X"05",X"21",X"58",X"86",X"36",X"00",
		X"C3",X"17",X"05",X"C3",X"17",X"05",X"13",X"68",X"12",X"20",X"11",X"58",X"10",X"20",X"11",X"09",
		X"13",X"01",X"20",X"00",X"00",X"78",X"10",X"28",X"00",X"10",X"10",X"20",X"00",X"FA",X"00",X"80",
		X"10",X"20",X"00",X"10",X"10",X"20",X"00",X"FA",X"00",X"88",X"10",X"18",X"00",X"10",X"10",X"20",
		X"00",X"FA",X"00",X"90",X"10",X"10",X"00",X"10",X"10",X"20",X"00",X"FA",X"00",X"68",X"10",X"38",
		X"31",X"02",X"30",X"02",X"31",X"02",X"30",X"02",X"31",X"02",X"21",X"01",X"22",X"01",X"23",X"03",
		X"20",X"01",X"30",X"01",X"10",X"1F",X"00",X"FA",X"00",X"B0",X"10",X"20",X"00",X"FA",X"40",X"3A",
		X"6F",X"86",X"E6",X"F0",X"FE",X"20",X"20",X"06",X"21",X"58",X"86",X"36",X"01",X"C9",X"FE",X"10",
		X"C0",X"3A",X"AE",X"85",X"32",X"AF",X"85",X"21",X"22",X"98",X"11",X"22",X"99",X"3A",X"6F",X"86",
		X"E6",X"03",X"20",X"15",X"36",X"00",X"AF",X"12",X"21",X"A3",X"98",X"35",X"35",X"AF",X"32",X"AE",
		X"85",X"3E",X"04",X"32",X"8B",X"80",X"C3",X"D4",X"0C",X"FE",X"01",X"20",X"15",X"36",X"02",X"AF",
		X"12",X"21",X"A2",X"98",X"34",X"34",X"3E",X"02",X"32",X"AE",X"85",X"3E",X"05",X"32",X"6B",X"83",
		X"18",X"32",X"FE",X"02",X"20",X"1F",X"36",X"00",X"3E",X"01",X"12",X"21",X"A3",X"98",X"34",X"34",
		X"3E",X"04",X"32",X"AE",X"85",X"3E",X"8C",X"32",X"63",X"83",X"32",X"43",X"83",X"32",X"62",X"83",
		X"32",X"42",X"83",X"18",X"0F",X"36",X"02",X"3E",X"02",X"12",X"21",X"A2",X"98",X"35",X"35",X"3E",
		X"06",X"32",X"AE",X"85",X"3A",X"A3",X"98",X"FE",X"10",X"20",X"07",X"21",X"22",X"98",X"34",X"34",
		X"34",X"34",X"21",X"76",X"86",X"34",X"CB",X"46",X"C0",X"21",X"22",X"98",X"34",X"C9",X"3A",X"70",
		X"86",X"21",X"E4",X"98",X"11",X"64",X"98",X"CD",X"2F",X"0D",X"C9",X"3A",X"72",X"86",X"21",X"D4",
		X"98",X"11",X"54",X"98",X"CD",X"47",X"0D",X"C9",X"3A",X"73",X"86",X"21",X"D6",X"98",X"11",X"56",
		X"98",X"CD",X"47",X"0D",X"C9",X"3A",X"74",X"86",X"21",X"D8",X"98",X"11",X"58",X"98",X"CD",X"47",
		X"0D",X"C9",X"3A",X"75",X"86",X"21",X"DA",X"98",X"11",X"5A",X"98",X"CD",X"47",X"0D",X"C9",X"F5",
		X"3E",X"21",X"12",X"01",X"77",X"86",X"0A",X"3C",X"02",X"E6",X"07",X"FE",X"02",X"30",X"03",X"1A",
		X"3D",X"12",X"F1",X"CD",X"47",X"0D",X"C9",X"E6",X"F0",X"C8",X"35",X"35",X"C9",X"21",X"6C",X"98",
		X"36",X"24",X"11",X"78",X"86",X"1A",X"3C",X"12",X"CB",X"57",X"20",X"01",X"34",X"3A",X"71",X"86",
		X"E6",X"F0",X"C8",X"FE",X"10",X"20",X"06",X"21",X"EC",X"98",X"35",X"35",X"C9",X"FE",X"30",X"20",
		X"10",X"3A",X"71",X"86",X"21",X"6D",X"98",X"CB",X"47",X"20",X"03",X"36",X"02",X"C9",X"36",X"0C",
		X"C9",X"DD",X"21",X"A4",X"98",X"3A",X"EC",X"98",X"D6",X"10",X"DD",X"77",X"00",X"D6",X"10",X"DD",
		X"77",X"02",X"D6",X"10",X"DD",X"77",X"04",X"3A",X"ED",X"98",X"DD",X"77",X"01",X"DD",X"77",X"03",
		X"DD",X"77",X"05",X"DD",X"21",X"24",X"98",X"3A",X"71",X"86",X"E6",X"0F",X"20",X"1A",X"3E",X"32",
		X"DD",X"77",X"00",X"DD",X"77",X"02",X"DD",X"77",X"04",X"DD",X"21",X"A4",X"98",X"06",X"06",X"DD",
		X"36",X"00",X"00",X"DD",X"23",X"10",X"F8",X"C9",X"FE",X"01",X"20",X"0E",X"3E",X"2C",X"DD",X"77",
		X"00",X"3E",X"32",X"DD",X"77",X"02",X"DD",X"77",X"04",X"C9",X"FE",X"02",X"20",X"0F",X"3E",X"2D",
		X"DD",X"77",X"00",X"3C",X"DD",X"77",X"02",X"3E",X"32",X"DD",X"77",X"04",X"C9",X"3E",X"2F",X"DD",
		X"77",X"00",X"3C",X"DD",X"77",X"02",X"3C",X"DD",X"77",X"04",X"C9",X"FE",X"06",X"DA",X"17",X"05",
		X"FE",X"17",X"30",X"10",X"3A",X"76",X"86",X"CB",X"47",X"CA",X"17",X"05",X"0E",X"FF",X"CD",X"2E",
		X"0E",X"C3",X"17",X"05",X"FE",X"1A",X"DA",X"17",X"05",X"FE",X"29",X"D2",X"17",X"05",X"3A",X"76",
		X"86",X"CB",X"47",X"CA",X"17",X"05",X"0E",X"01",X"CD",X"2E",X"0E",X"C3",X"17",X"05",X"21",X"C1",
		X"98",X"06",X"0A",X"7E",X"81",X"77",X"23",X"23",X"10",X"F9",X"C9",X"EB",X"D5",X"DD",X"E1",X"11",
		X"20",X"00",X"DD",X"7E",X"00",X"DD",X"23",X"77",X"19",X"10",X"F7",X"C9",X"21",X"80",X"98",X"11",
		X"80",X"93",X"06",X"40",X"3A",X"F0",X"87",X"CB",X"5F",X"C0",X"3A",X"00",X"84",X"CB",X"4F",X"28",
		X"06",X"CB",X"57",X"28",X"02",X"18",X"0D",X"7E",X"12",X"23",X"13",X"7E",X"C6",X"37",X"12",X"23",
		X"13",X"10",X"F4",X"C9",X"3E",X"F2",X"96",X"12",X"13",X"23",X"3E",X"27",X"96",X"12",X"23",X"13",
		X"10",X"F2",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3A",X"85",X"87",X"CB",X"7F",X"20",X"07",X"3A",X"57",X"86",X"CB",X"4F",X"28",X"05",X"21",X"70",
		X"89",X"18",X"03",X"21",X"B0",X"85",X"7E",X"E6",X"0E",X"E5",X"7E",X"E6",X"0F",X"FE",X"08",X"20",
		X"07",X"21",X"AE",X"85",X"CB",X"F6",X"E1",X"C9",X"21",X"AE",X"85",X"7E",X"23",X"E6",X"3F",X"77",
		X"E1",X"7E",X"E6",X"3F",X"32",X"AE",X"85",X"E6",X"0F",X"6F",X"3A",X"AF",X"85",X"E6",X"0F",X"BD",
		X"20",X"06",X"21",X"AE",X"85",X"CB",X"BE",X"C9",X"21",X"AE",X"85",X"CB",X"FE",X"C9",X"21",X"01",
		X"84",X"CB",X"5E",X"28",X"30",X"21",X"AE",X"85",X"7E",X"21",X"22",X"98",X"11",X"22",X"99",X"E6",
		X"0F",X"28",X"0D",X"FE",X"04",X"28",X"0E",X"FE",X"02",X"28",X"10",X"FE",X"06",X"28",X"10",X"C9",
		X"36",X"10",X"AF",X"12",X"C9",X"36",X"10",X"3E",X"01",X"12",X"C9",X"36",X"11",X"18",X"F3",X"36",
		X"11",X"3E",X"02",X"12",X"C9",X"21",X"AE",X"85",X"7E",X"21",X"22",X"98",X"11",X"22",X"99",X"01",
		X"00",X"00",X"E6",X"0F",X"28",X"13",X"03",X"FE",X"04",X"28",X"0E",X"01",X"00",X"02",X"FE",X"02",
		X"28",X"07",X"03",X"03",X"FE",X"06",X"28",X"01",X"C9",X"70",X"79",X"12",X"3A",X"01",X"84",X"CB",
		X"67",X"C8",X"34",X"34",X"34",X"34",X"C9",X"3A",X"AE",X"85",X"E6",X"0F",X"20",X"1A",X"3E",X"02",
		X"32",X"AE",X"85",X"CD",X"4E",X"10",X"C9",X"CD",X"00",X"10",X"AF",X"32",X"A0",X"98",X"32",X"A1",
		X"98",X"3A",X"A3",X"98",X"FE",X"08",X"28",X"DF",X"CD",X"1F",X"11",X"CD",X"8F",X"11",X"CD",X"EA",
		X"11",X"21",X"AE",X"85",X"7E",X"E6",X"0F",X"FE",X"08",X"28",X"47",X"7E",X"CB",X"76",X"20",X"42",
		X"3A",X"B3",X"85",X"21",X"B1",X"85",X"96",X"32",X"B3",X"85",X"D0",X"3A",X"AE",X"85",X"CB",X"7F",
		X"28",X"04",X"CD",X"4E",X"10",X"C9",X"CD",X"4E",X"10",X"21",X"B2",X"85",X"34",X"CB",X"46",X"28",
		X"04",X"21",X"22",X"98",X"34",X"3A",X"01",X"84",X"CB",X"57",X"C0",X"CD",X"36",X"11",X"C9",X"3A",
		X"01",X"84",X"CB",X"67",X"20",X"06",X"3E",X"40",X"32",X"B1",X"85",X"C9",X"3E",X"50",X"32",X"B1",
		X"85",X"C9",X"CD",X"4E",X"10",X"C9",X"21",X"AE",X"85",X"7E",X"21",X"A3",X"98",X"E6",X"0F",X"28",
		X"25",X"FE",X"04",X"28",X"13",X"2B",X"FE",X"02",X"28",X"0E",X"FE",X"06",X"28",X"18",X"C9",X"3A",
		X"A3",X"98",X"5F",X"3A",X"A2",X"98",X"57",X"C9",X"34",X"34",X"CD",X"4F",X"11",X"CD",X"74",X"11",
		X"CB",X"49",X"C8",X"35",X"35",X"C9",X"35",X"35",X"CD",X"4F",X"11",X"CD",X"74",X"11",X"CB",X"49",
		X"C8",X"34",X"34",X"C9",X"F5",X"CB",X"89",X"7A",X"FE",X"11",X"38",X"0F",X"FE",X"E2",X"30",X"0B",
		X"7B",X"FE",X"08",X"38",X"06",X"FE",X"F1",X"30",X"02",X"F1",X"C9",X"CB",X"C9",X"F1",X"C9",X"E5",
		X"C5",X"21",X"AE",X"85",X"7E",X"E6",X"0F",X"28",X"04",X"FE",X"04",X"20",X"0B",X"3A",X"A2",X"98",
		X"E6",X"0F",X"FE",X"01",X"28",X"26",X"18",X"19",X"FE",X"02",X"28",X"04",X"FE",X"06",X"20",X"1C",
		X"3A",X"A3",X"98",X"FE",X"20",X"30",X"06",X"FE",X"08",X"28",X"11",X"18",X"04",X"E6",X"0F",X"28",
		X"0B",X"23",X"7E",X"E6",X"0F",X"2B",X"77",X"CB",X"87",X"C1",X"E1",X"C9",X"3A",X"57",X"86",X"CB",
		X"4F",X"20",X"13",X"3A",X"AE",X"85",X"E6",X"0F",X"4F",X"3A",X"AF",X"85",X"E6",X"0F",X"B9",X"28",
		X"05",X"21",X"B3",X"85",X"36",X"02",X"CB",X"C7",X"18",X"DF",X"3A",X"AE",X"85",X"21",X"A2",X"98",
		X"11",X"E1",X"85",X"E6",X"0F",X"28",X"0D",X"FE",X"04",X"28",X"13",X"FE",X"02",X"28",X"19",X"FE",
		X"06",X"28",X"1F",X"C9",X"7E",X"12",X"23",X"1B",X"7E",X"D6",X"10",X"12",X"18",X"1C",X"7E",X"12",
		X"23",X"1B",X"7E",X"C6",X"10",X"12",X"18",X"12",X"7E",X"C6",X"10",X"12",X"23",X"1B",X"7E",X"12",
		X"18",X"08",X"7E",X"D6",X"10",X"12",X"23",X"1B",X"7E",X"12",X"21",X"65",X"84",X"06",X"08",X"11",
		X"08",X"00",X"E5",X"3A",X"E1",X"85",X"BE",X"20",X"0E",X"3A",X"E0",X"85",X"23",X"BE",X"20",X"07",
		X"E1",X"21",X"01",X"84",X"CB",X"D6",X"C9",X"21",X"01",X"84",X"CB",X"96",X"E1",X"19",X"10",X"E2",
		X"C9",X"3A",X"57",X"86",X"CB",X"4F",X"28",X"1C",X"21",X"28",X"85",X"11",X"10",X"00",X"06",X"08",
		X"0E",X"08",X"CB",X"7E",X"28",X"01",X"0D",X"19",X"10",X"F8",X"79",X"FE",X"01",X"20",X"05",X"21",
		X"76",X"86",X"36",X"90",X"2A",X"25",X"86",X"11",X"60",X"09",X"A7",X"ED",X"52",X"20",X"05",X"21",
		X"53",X"86",X"CB",X"CE",X"2A",X"25",X"86",X"7C",X"A7",X"20",X"27",X"7D",X"FE",X"96",X"28",X"0A",
		X"A7",X"20",X"1F",X"21",X"46",X"86",X"CB",X"DE",X"18",X"1C",X"3A",X"4A",X"86",X"CB",X"6F",X"20",
		X"11",X"CB",X"EF",X"32",X"4A",X"86",X"3A",X"F0",X"87",X"CB",X"47",X"20",X"05",X"3E",X"01",X"32",
		X"89",X"9A",X"2B",X"22",X"25",X"86",X"21",X"4A",X"86",X"CB",X"66",X"C0",X"21",X"28",X"85",X"06",
		X"08",X"0E",X"08",X"11",X"10",X"00",X"CB",X"7E",X"28",X"01",X"0D",X"19",X"10",X"F8",X"79",X"A7",
		X"C8",X"21",X"00",X"84",X"3A",X"0D",X"84",X"CB",X"4E",X"28",X"03",X"3A",X"0E",X"84",X"06",X"02",
		X"FE",X"04",X"38",X"1B",X"04",X"FE",X"08",X"38",X"16",X"04",X"FE",X"0C",X"38",X"11",X"04",X"FE",
		X"10",X"38",X"0C",X"04",X"FE",X"14",X"38",X"07",X"04",X"FE",X"18",X"38",X"02",X"18",X"03",X"79",
		X"B8",X"D0",X"21",X"04",X"01",X"22",X"25",X"86",X"21",X"4A",X"86",X"CB",X"E6",X"C9",X"2A",X"D6",
		X"85",X"22",X"DE",X"85",X"3A",X"A2",X"98",X"57",X"3A",X"A3",X"98",X"5F",X"CD",X"93",X"13",X"CD",
		X"53",X"13",X"2A",X"D6",X"85",X"3A",X"DE",X"85",X"BD",X"20",X"06",X"3A",X"DF",X"85",X"BC",X"28",
		X"0C",X"3A",X"46",X"86",X"CB",X"47",X"C0",X"CD",X"0A",X"14",X"CD",X"0A",X"14",X"3A",X"46",X"86",
		X"CB",X"47",X"C0",X"3A",X"AE",X"85",X"E6",X"07",X"47",X"3A",X"AF",X"85",X"E6",X"07",X"B8",X"C4",
		X"EF",X"14",X"C9",X"06",X"00",X"2A",X"D6",X"85",X"CD",X"04",X"14",X"2A",X"D8",X"85",X"CD",X"04",
		X"14",X"2A",X"DA",X"85",X"CD",X"04",X"14",X"2A",X"DC",X"85",X"CD",X"04",X"14",X"78",X"21",X"01",
		X"84",X"CB",X"A6",X"A7",X"C0",X"CB",X"E6",X"C9",X"CD",X"CB",X"13",X"DD",X"21",X"FA",X"85",X"18",
		X"2C",X"CD",X"CB",X"13",X"DD",X"21",X"02",X"86",X"18",X"23",X"CD",X"CB",X"13",X"DD",X"21",X"0A",
		X"86",X"18",X"1A",X"3A",X"AE",X"85",X"E6",X"0F",X"28",X"0C",X"FE",X"06",X"28",X"08",X"3E",X"06",
		X"82",X"57",X"3E",X"06",X"83",X"5F",X"CD",X"CB",X"13",X"DD",X"21",X"D6",X"85",X"DD",X"75",X"00",
		X"DD",X"74",X"01",X"CD",X"FD",X"13",X"DD",X"73",X"02",X"DD",X"72",X"03",X"23",X"DD",X"75",X"04",
		X"DD",X"74",X"05",X"13",X"DD",X"73",X"06",X"DD",X"72",X"07",X"C9",X"7A",X"D6",X"11",X"CB",X"3F",
		X"CB",X"3F",X"57",X"CB",X"3F",X"CB",X"27",X"CB",X"27",X"CB",X"27",X"CB",X"27",X"CB",X"27",X"6F",
		X"7A",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"67",X"16",X"00",X"CB",X"3B",X"CB",X"3B",
		X"CB",X"3B",X"A7",X"ED",X"52",X"EB",X"21",X"A0",X"83",X"A7",X"ED",X"52",X"C9",X"11",X"E0",X"FF",
		X"EB",X"19",X"EB",X"C9",X"7E",X"FE",X"7F",X"C0",X"04",X"C9",X"2A",X"D6",X"85",X"E5",X"DD",X"E1",
		X"ED",X"4B",X"D8",X"85",X"2A",X"DA",X"85",X"ED",X"5B",X"DC",X"85",X"3A",X"AE",X"85",X"E6",X"0F",
		X"28",X"10",X"FE",X"04",X"CA",X"DC",X"14",X"FE",X"02",X"CA",X"D4",X"14",X"FE",X"06",X"CA",X"85",
		X"14",X"C9",X"7E",X"FE",X"08",X"CA",X"E4",X"14",X"FE",X"09",X"CA",X"E4",X"14",X"FE",X"0C",X"28",
		X"1B",X"FE",X"8D",X"38",X"04",X"FE",X"90",X"38",X"13",X"FE",X"8C",X"28",X"0F",X"FE",X"7F",X"CC",
		X"CB",X"15",X"FE",X"7E",X"20",X"04",X"36",X"8C",X"18",X"02",X"36",X"03",X"1A",X"FE",X"08",X"CA",
		X"E7",X"14",X"FE",X"09",X"CA",X"E7",X"14",X"FE",X"0C",X"C8",X"FE",X"8D",X"38",X"03",X"FE",X"90",
		X"D8",X"FE",X"8C",X"C8",X"FE",X"7F",X"CC",X"CB",X"15",X"FE",X"7E",X"20",X"04",X"3E",X"8C",X"12",
		X"C9",X"3E",X"02",X"12",X"C9",X"0A",X"FE",X"02",X"28",X"61",X"FE",X"03",X"28",X"5D",X"FE",X"7F",
		X"28",X"16",X"FE",X"0C",X"28",X"18",X"FE",X"8C",X"28",X"14",X"FE",X"7E",X"28",X"10",X"FE",X"8D",
		X"38",X"04",X"FE",X"90",X"38",X"08",X"FE",X"7F",X"CC",X"CB",X"15",X"3E",X"08",X"02",X"1A",X"FE",
		X"02",X"28",X"34",X"FE",X"03",X"28",X"30",X"FE",X"7F",X"28",X"12",X"FE",X"0C",X"C8",X"FE",X"8C",
		X"C8",X"FE",X"7E",X"C8",X"FE",X"8D",X"38",X"03",X"FE",X"90",X"D8",X"FE",X"7F",X"CC",X"CB",X"15",
		X"3E",X"09",X"12",X"C9",X"DD",X"E5",X"C1",X"E5",X"D1",X"C3",X"85",X"14",X"DD",X"E5",X"E1",X"C5",
		X"D1",X"C3",X"32",X"14",X"36",X"0C",X"C9",X"3E",X"0C",X"12",X"C9",X"3E",X"0C",X"02",X"C9",X"CD",
		X"D3",X"15",X"2A",X"DC",X"85",X"E5",X"FD",X"E1",X"2A",X"DA",X"85",X"E5",X"DD",X"E1",X"2A",X"D6",
		X"85",X"ED",X"5B",X"D8",X"85",X"3A",X"AE",X"85",X"E6",X"0F",X"28",X"0D",X"FE",X"02",X"28",X"25",
		X"FE",X"04",X"28",X"39",X"FE",X"06",X"28",X"4A",X"C9",X"DD",X"7E",X"00",X"CD",X"7B",X"15",X"CB",
		X"47",X"28",X"04",X"DD",X"36",X"00",X"05",X"FD",X"7E",X"00",X"CD",X"7B",X"15",X"CB",X"47",X"C8",
		X"FD",X"36",X"00",X"04",X"C9",X"7E",X"CD",X"7B",X"15",X"CB",X"47",X"28",X"02",X"36",X"06",X"DD",
		X"7E",X"00",X"CD",X"7B",X"15",X"CB",X"47",X"C8",X"DD",X"36",X"00",X"07",X"C9",X"7E",X"CD",X"7B",
		X"15",X"CB",X"47",X"28",X"02",X"36",X"01",X"1A",X"CD",X"7B",X"15",X"CB",X"47",X"C8",X"3E",X"00",
		X"12",X"C9",X"1A",X"CD",X"7B",X"15",X"CB",X"47",X"28",X"03",X"3E",X"0A",X"12",X"FD",X"7E",X"00",
		X"CD",X"7B",X"15",X"CB",X"47",X"C8",X"FD",X"36",X"00",X"0B",X"C9",X"F5",X"3A",X"01",X"84",X"CB",
		X"7F",X"20",X"10",X"3A",X"AE",X"85",X"C6",X"04",X"E6",X"07",X"47",X"3A",X"AF",X"85",X"E6",X"07",
		X"B8",X"20",X"0B",X"F1",X"FE",X"7F",X"CC",X"CB",X"15",X"28",X"2D",X"CB",X"87",X"C9",X"F1",X"FE",
		X"7F",X"CC",X"CB",X"15",X"28",X"22",X"A7",X"28",X"1F",X"FE",X"01",X"28",X"1B",X"FE",X"04",X"28",
		X"17",X"FE",X"05",X"28",X"13",X"FE",X"06",X"28",X"0F",X"FE",X"07",X"28",X"0B",X"FE",X"0A",X"28",
		X"07",X"FE",X"0B",X"28",X"03",X"CB",X"87",X"C9",X"CB",X"C7",X"C9",X"E5",X"21",X"56",X"86",X"CB",
		X"D6",X"E1",X"C9",X"3A",X"A2",X"98",X"57",X"3A",X"A3",X"98",X"5F",X"3A",X"AF",X"85",X"C3",X"96",
		X"13",X"38",X"00",X"38",X"00",X"25",X"32",X"00",X"13",X"38",X"00",X"02",X"30",X"00",X"3B",X"10",
		X"00",X"01",X"00",X"00",X"01",X"10",X"00",X"69",X"30",X"00",X"3F",X"38",X"00",X"01",X"32",X"00",
		X"77",X"12",X"00",X"01",X"02",X"00",X"01",X"12",X"00",X"75",X"32",X"00",X"35",X"38",X"00",X"01",
		X"34",X"01",X"5E",X"38",X"00",X"01",X"36",X"00",X"4B",X"30",X"00",X"28",X"38",X"00",X"01",X"36",
		X"00",X"8C",X"38",X"00",X"01",X"30",X"00",X"3E",X"38",X"00",X"01",X"36",X"00",X"7B",X"38",X"00",
		X"02",X"30",X"00",X"05",X"38",X"00",X"01",X"36",X"00",X"27",X"38",X"00",X"02",X"34",X"00",X"73",
		X"38",X"00",X"01",X"32",X"01",X"7E",X"32",X"00",X"02",X"30",X"00",X"42",X"38",X"00",X"01",X"36",
		X"00",X"9A",X"30",X"00",X"89",X"38",X"00",X"07",X"30",X"00",X"7B",X"38",X"00",X"02",X"34",X"00",
		X"02",X"14",X"00",X"01",X"04",X"00",X"01",X"14",X"00",X"03",X"18",X"00",X"79",X"38",X"00",X"2D",
		X"36",X"00",X"6D",X"38",X"00",X"01",X"34",X"00",X"EE",X"38",X"00",X"04",X"30",X"00",X"3C",X"38",
		X"00",X"02",X"18",X"00",X"01",X"08",X"00",X"01",X"18",X"00",X"2E",X"14",X"00",X"04",X"34",X"00",
		X"0C",X"38",X"00",X"01",X"30",X"00",X"02",X"10",X"00",X"01",X"00",X"00",X"01",X"10",X"00",X"13",
		X"30",X"00",X"9D",X"38",X"00",X"02",X"34",X"00",X"03",X"14",X"00",X"01",X"04",X"00",X"01",X"14",
		X"00",X"04",X"18",X"00",X"33",X"10",X"00",X"03",X"30",X"00",X"60",X"38",X"00",X"01",X"36",X"00",
		X"10",X"38",X"00",X"01",X"30",X"00",X"24",X"32",X"00",X"85",X"38",X"00",X"01",X"34",X"01",X"71",
		X"38",X"00",X"03",X"36",X"00",X"5B",X"38",X"00",X"03",X"32",X"00",X"0F",X"38",X"00",X"01",X"30",
		X"00",X"CF",X"38",X"00",X"01",X"32",X"00",X"76",X"38",X"00",X"01",X"30",X"00",X"47",X"38",X"00",
		X"1F",X"30",X"00",X"11",X"38",X"00",X"01",X"36",X"00",X"26",X"38",X"00",X"01",X"32",X"00",X"B1",
		X"2A",X"5A",X"86",X"23",X"22",X"5A",X"86",X"7C",X"FE",X"03",X"20",X"0E",X"7D",X"FE",X"1A",X"C2",
		X"17",X"05",X"21",X"58",X"86",X"36",X"06",X"C3",X"17",X"05",X"FE",X"02",X"20",X"1D",X"7D",X"FE",
		X"DE",X"CA",X"81",X"18",X"FE",X"32",X"CA",X"21",X"19",X"FE",X"22",X"CA",X"17",X"19",X"FE",X"12",
		X"CA",X"2D",X"18",X"FE",X"02",X"CA",X"FB",X"18",X"C3",X"17",X"05",X"FE",X"01",X"20",X"2F",X"7D",
		X"FE",X"F2",X"CA",X"2D",X"18",X"FE",X"E2",X"CA",X"09",X"19",X"FE",X"BE",X"CA",X"F0",X"18",X"D2",
		X"17",X"05",X"FE",X"BA",X"D2",X"E7",X"17",X"FE",X"B2",X"D2",X"EC",X"17",X"FE",X"AA",X"D2",X"F1",
		X"17",X"FE",X"A9",X"CA",X"A3",X"18",X"FE",X"6D",X"CA",X"81",X"18",X"C3",X"17",X"05",X"7D",X"FE",
		X"C2",X"CA",X"47",X"18",X"FE",X"B2",X"CA",X"33",X"18",X"FE",X"A2",X"CA",X"2D",X"18",X"FE",X"92",
		X"CA",X"04",X"18",X"FE",X"82",X"CA",X"2D",X"18",X"FE",X"72",X"CA",X"16",X"18",X"FE",X"52",X"CA",
		X"F9",X"17",X"D2",X"17",X"05",X"FE",X"4F",X"30",X"3C",X"FE",X"47",X"30",X"3D",X"FE",X"3F",X"30",
		X"3E",X"FE",X"3E",X"CA",X"9F",X"18",X"FE",X"02",X"28",X"03",X"C3",X"17",X"05",X"21",X"A2",X"98",
		X"36",X"82",X"23",X"36",X"90",X"21",X"22",X"98",X"36",X"06",X"23",X"36",X"00",X"21",X"22",X"99",
		X"36",X"02",X"21",X"88",X"98",X"36",X"82",X"23",X"36",X"90",X"21",X"08",X"98",X"36",X"13",X"23",
		X"36",X"06",X"C3",X"17",X"05",X"21",X"82",X"98",X"35",X"35",X"21",X"84",X"98",X"35",X"35",X"21",
		X"86",X"98",X"35",X"35",X"C3",X"17",X"05",X"21",X"82",X"98",X"34",X"34",X"21",X"84",X"98",X"34",
		X"34",X"21",X"86",X"98",X"34",X"34",X"C3",X"17",X"05",X"CD",X"61",X"19",X"21",X"64",X"98",X"36",
		X"23",X"C3",X"17",X"05",X"CD",X"5B",X"19",X"21",X"64",X"98",X"36",X"81",X"21",X"E5",X"98",X"7E",
		X"D6",X"03",X"77",X"C3",X"17",X"05",X"CD",X"5B",X"19",X"21",X"64",X"98",X"36",X"80",X"21",X"E4",
		X"98",X"7E",X"D6",X"08",X"77",X"23",X"7E",X"D6",X"04",X"77",X"C3",X"17",X"05",X"CD",X"61",X"19",
		X"C3",X"17",X"05",X"CD",X"5B",X"19",X"21",X"64",X"98",X"34",X"21",X"82",X"98",X"06",X"06",X"36",
		X"00",X"23",X"10",X"FB",X"C3",X"17",X"05",X"21",X"F4",X"98",X"06",X"04",X"0E",X"90",X"3E",X"37",
		X"77",X"C6",X"10",X"23",X"71",X"23",X"10",X"F8",X"36",X"51",X"23",X"71",X"21",X"64",X"98",X"36",
		X"32",X"21",X"E4",X"98",X"36",X"00",X"23",X"36",X"00",X"21",X"77",X"18",X"11",X"74",X"98",X"01",
		X"0A",X"00",X"ED",X"B0",X"C3",X"8E",X"18",X"39",X"0A",X"47",X"0A",X"3C",X"0A",X"47",X"0A",X"65",
		X"00",X"21",X"F4",X"98",X"06",X"0A",X"36",X"00",X"23",X"10",X"FB",X"C3",X"17",X"05",X"21",X"22",
		X"98",X"36",X"06",X"21",X"22",X"99",X"36",X"00",X"2B",X"2B",X"36",X"00",X"C3",X"17",X"05",X"06",
		X"02",X"18",X"02",X"06",X"00",X"21",X"22",X"98",X"36",X"11",X"DD",X"21",X"82",X"98",X"FD",X"21",
		X"02",X"98",X"3E",X"82",X"0E",X"90",X"DD",X"77",X"00",X"DD",X"77",X"02",X"DD",X"77",X"04",X"DD",
		X"71",X"01",X"DD",X"71",X"03",X"DD",X"71",X"05",X"FD",X"36",X"00",X"37",X"FD",X"36",X"02",X"37",
		X"FD",X"36",X"04",X"36",X"FD",X"36",X"01",X"08",X"FD",X"36",X"03",X"08",X"FD",X"36",X"05",X"08",
		X"DD",X"21",X"02",X"99",X"DD",X"70",X"00",X"DD",X"70",X"02",X"DD",X"70",X"04",X"C3",X"17",X"05",
		X"CD",X"61",X"19",X"21",X"6C",X"98",X"36",X"27",X"C3",X"17",X"05",X"CD",X"5B",X"19",X"21",X"6C",
		X"98",X"36",X"84",X"21",X"ED",X"98",X"C3",X"0F",X"18",X"CD",X"5B",X"19",X"21",X"6C",X"98",X"36",
		X"83",X"21",X"EC",X"98",X"C3",X"21",X"18",X"CD",X"5B",X"19",X"21",X"6C",X"98",X"34",X"C3",X"3A",
		X"18",X"21",X"6C",X"98",X"36",X"32",X"21",X"EC",X"98",X"36",X"00",X"23",X"36",X"00",X"21",X"F4",
		X"98",X"06",X"04",X"0E",X"90",X"3E",X"97",X"77",X"C6",X"10",X"23",X"71",X"23",X"10",X"F8",X"36",
		X"B1",X"23",X"71",X"21",X"51",X"19",X"11",X"74",X"98",X"01",X"0A",X"00",X"ED",X"B0",X"C3",X"8E",
		X"18",X"39",X"0A",X"47",X"0A",X"3F",X"0A",X"47",X"0A",X"65",X"00",X"21",X"22",X"98",X"36",X"0D",
		X"C9",X"21",X"22",X"98",X"36",X"0C",X"C9",X"21",X"6C",X"89",X"CB",X"4E",X"C2",X"E3",X"19",X"CB",
		X"46",X"20",X"30",X"21",X"F0",X"87",X"CB",X"46",X"20",X"51",X"21",X"6D",X"89",X"36",X"00",X"21",
		X"28",X"85",X"0E",X"00",X"06",X"08",X"32",X"30",X"68",X"11",X"10",X"00",X"CB",X"7E",X"28",X"01",
		X"0C",X"19",X"32",X"30",X"68",X"10",X"F5",X"79",X"FE",X"07",X"20",X"2F",X"21",X"F0",X"87",X"CB",
		X"C6",X"18",X"40",X"21",X"A1",X"83",X"36",X"7E",X"23",X"7E",X"FE",X"0E",X"28",X"04",X"FE",X"0F",
		X"20",X"02",X"36",X"7E",X"11",X"20",X"00",X"19",X"3E",X"7E",X"77",X"2B",X"77",X"19",X"77",X"23",
		X"77",X"21",X"86",X"9A",X"36",X"01",X"21",X"6C",X"89",X"CB",X"CE",X"00",X"3A",X"F0",X"87",X"CB",
		X"47",X"28",X"10",X"21",X"6D",X"89",X"7E",X"FE",X"1E",X"20",X"07",X"21",X"6C",X"89",X"CB",X"C6",
		X"18",X"01",X"34",X"00",X"3A",X"00",X"84",X"CB",X"4F",X"20",X"0E",X"2A",X"D4",X"87",X"22",X"ED",
		X"87",X"3A",X"DA",X"87",X"32",X"EB",X"87",X"18",X"0C",X"3A",X"D8",X"87",X"32",X"EB",X"87",X"2A",
		X"D2",X"87",X"22",X"ED",X"87",X"3A",X"99",X"87",X"21",X"EB",X"87",X"CB",X"47",X"28",X"06",X"CB",
		X"87",X"32",X"99",X"87",X"34",X"00",X"3A",X"EB",X"87",X"FE",X"02",X"20",X"21",X"21",X"F0",X"87",
		X"CB",X"EE",X"CD",X"1E",X"1B",X"21",X"EF",X"87",X"36",X"46",X"21",X"F0",X"87",X"CB",X"B6",X"21",
		X"9E",X"98",X"36",X"71",X"23",X"36",X"80",X"21",X"EB",X"87",X"34",X"C3",X"02",X"1B",X"3A",X"F0",
		X"87",X"CB",X"6F",X"28",X"1F",X"2A",X"ED",X"87",X"23",X"22",X"ED",X"87",X"11",X"58",X"02",X"A7",
		X"ED",X"52",X"20",X"10",X"21",X"9E",X"98",X"36",X"00",X"23",X"36",X"E0",X"21",X"F0",X"87",X"CB",
		X"AE",X"C3",X"02",X"1B",X"3A",X"01",X"84",X"CB",X"7F",X"C0",X"3A",X"00",X"84",X"CB",X"6F",X"20",
		X"06",X"3A",X"57",X"86",X"CB",X"4F",X"C8",X"21",X"9E",X"98",X"11",X"A2",X"98",X"1A",X"BE",X"20",
		X"0E",X"23",X"13",X"1A",X"BE",X"20",X"08",X"3A",X"F0",X"87",X"CB",X"F7",X"32",X"F0",X"87",X"3A",
		X"F0",X"87",X"CB",X"77",X"CA",X"02",X"1B",X"21",X"EF",X"87",X"7E",X"A7",X"CA",X"02",X"1B",X"35",
		X"7E",X"FE",X"44",X"20",X"3C",X"21",X"93",X"9A",X"36",X"01",X"21",X"A7",X"87",X"CB",X"C6",X"3A",
		X"E6",X"87",X"32",X"76",X"98",X"AF",X"32",X"77",X"98",X"21",X"7E",X"98",X"36",X"64",X"23",X"36",
		X"00",X"3A",X"9E",X"98",X"D6",X"08",X"32",X"F6",X"98",X"C6",X"10",X"32",X"FE",X"98",X"3A",X"9F",
		X"98",X"32",X"F7",X"98",X"32",X"FF",X"98",X"21",X"9E",X"98",X"36",X"00",X"23",X"36",X"E0",X"18",
		X"21",X"FE",X"02",X"20",X"12",X"21",X"F6",X"98",X"36",X"00",X"23",X"36",X"00",X"21",X"FE",X"98",
		X"36",X"00",X"23",X"36",X"00",X"18",X"0B",X"FE",X"01",X"20",X"07",X"36",X"00",X"21",X"F0",X"87",
		X"CB",X"B6",X"3A",X"00",X"84",X"CB",X"4F",X"2A",X"ED",X"87",X"3A",X"EB",X"87",X"20",X"08",X"32",
		X"DA",X"87",X"22",X"D4",X"87",X"18",X"06",X"32",X"D8",X"87",X"22",X"D2",X"87",X"C9",X"3A",X"00",
		X"84",X"CB",X"4F",X"20",X"05",X"21",X"0D",X"84",X"18",X"03",X"21",X"0E",X"84",X"7E",X"21",X"E8",
		X"87",X"FE",X"12",X"38",X"02",X"3E",X"12",X"77",X"D6",X"01",X"87",X"87",X"5F",X"16",X"00",X"21",
		X"57",X"1B",X"19",X"7E",X"32",X"1E",X"98",X"23",X"7E",X"32",X"1F",X"98",X"23",X"7E",X"32",X"E7",
		X"87",X"23",X"7E",X"32",X"E6",X"87",X"C9",X"53",X"0E",X"04",X"5D",X"55",X"10",X"06",X"5E",X"58",
		X"12",X"08",X"5F",X"54",X"0F",X"10",X"60",X"54",X"0F",X"10",X"60",X"57",X"11",X"20",X"4E",X"57",
		X"11",X"20",X"4E",X"56",X"10",X"30",X"4F",X"56",X"10",X"30",X"4F",X"59",X"13",X"40",X"61",X"59",
		X"13",X"40",X"61",X"5A",X"14",X"50",X"50",X"5A",X"14",X"50",X"50",X"52",X"0D",X"60",X"62",X"52",
		X"0D",X"60",X"62",X"5B",X"15",X"70",X"51",X"5B",X"15",X"70",X"51",X"5C",X"16",X"80",X"63",X"3A",
		X"57",X"86",X"CB",X"4F",X"28",X"04",X"3E",X"02",X"18",X"05",X"3A",X"8D",X"89",X"E6",X"03",X"87",
		X"87",X"87",X"87",X"6F",X"26",X"00",X"3A",X"10",X"84",X"3D",X"5F",X"16",X"00",X"19",X"EB",X"21",
		X"FE",X"1B",X"19",X"7E",X"32",X"BD",X"87",X"3A",X"00",X"84",X"CB",X"4F",X"20",X"05",X"3A",X"0D",
		X"84",X"18",X"03",X"3A",X"0E",X"84",X"21",X"BD",X"87",X"D6",X"1E",X"38",X"06",X"86",X"77",X"30",
		X"02",X"36",X"FF",X"21",X"3E",X"1C",X"06",X"06",X"DD",X"21",X"A0",X"87",X"E5",X"19",X"7E",X"E1",
		X"DD",X"77",X"00",X"D5",X"11",X"40",X"00",X"19",X"D1",X"DD",X"23",X"10",X"EF",X"C9",X"73",X"73",
		X"78",X"78",X"78",X"80",X"80",X"80",X"84",X"84",X"84",X"84",X"87",X"8C",X"96",X"80",X"78",X"78",
		X"78",X"78",X"78",X"80",X"80",X"84",X"84",X"84",X"84",X"84",X"87",X"8C",X"96",X"80",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"80",X"80",X"84",X"84",X"84",X"84",X"84",X"87",X"8C",X"96",X"80",X"7E",X"7E",
		X"7E",X"7E",X"7E",X"87",X"87",X"87",X"87",X"87",X"87",X"8A",X"8C",X"90",X"96",X"80",X"7C",X"80",
		X"80",X"85",X"89",X"92",X"96",X"9A",X"9F",X"9F",X"A3",X"A3",X"A3",X"A3",X"A8",X"80",X"80",X"85",
		X"89",X"89",X"8D",X"96",X"96",X"9A",X"9F",X"9F",X"A3",X"A3",X"A3",X"A3",X"A8",X"80",X"89",X"8D",
		X"91",X"92",X"92",X"9A",X"9A",X"9F",X"9F",X"A3",X"A3",X"A3",X"A3",X"A3",X"A8",X"80",X"92",X"92",
		X"96",X"96",X"9A",X"9F",X"9F",X"A3",X"A3",X"A8",X"A8",X"A8",X"AC",X"AC",X"B4",X"80",X"80",X"89",
		X"8D",X"92",X"9A",X"A3",X"A8",X"AC",X"AC",X"AC",X"B0",X"B4",X"B4",X"B8",X"BC",X"80",X"85",X"8D",
		X"96",X"9A",X"9F",X"A8",X"A8",X"AC",X"AC",X"B0",X"B0",X"B4",X"B4",X"B8",X"BC",X"80",X"92",X"96",
		X"9A",X"9F",X"A3",X"A8",X"A8",X"AC",X"AC",X"B0",X"B0",X"B4",X"B4",X"B8",X"BC",X"80",X"9A",X"9F",
		X"A3",X"A3",X"A8",X"AC",X"B0",X"B4",X"B4",X"B4",X"B8",X"B8",X"BC",X"C1",X"C5",X"80",X"AC",X"B0",
		X"B4",X"B4",X"BC",X"C1",X"C5",X"CA",X"CE",X"D2",X"D2",X"DB",X"DB",X"DF",X"DF",X"80",X"B0",X"B4",
		X"B8",X"BC",X"C1",X"CA",X"CA",X"CE",X"CE",X"D2",X"D7",X"DB",X"DB",X"DF",X"DF",X"80",X"B8",X"BC",
		X"C1",X"C5",X"CA",X"CE",X"CE",X"D2",X"D2",X"D7",X"D7",X"D2",X"D2",X"DF",X"DF",X"80",X"C1",X"C5",
		X"CA",X"CA",X"CE",X"D2",X"D7",X"DB",X"DB",X"DB",X"DF",X"DF",X"DF",X"DF",X"DF",X"80",X"85",X"89",
		X"89",X"8D",X"8D",X"9A",X"9F",X"A3",X"A8",X"A8",X"AC",X"AC",X"AC",X"AC",X"B0",X"80",X"89",X"8D",
		X"92",X"92",X"96",X"9F",X"9F",X"A3",X"A8",X"A8",X"AC",X"AC",X"AC",X"AC",X"B0",X"80",X"92",X"96",
		X"9A",X"9A",X"A4",X"A3",X"A3",X"A8",X"A8",X"AC",X"AC",X"AC",X"AC",X"AC",X"B0",X"80",X"9F",X"9F",
		X"A3",X"A3",X"A8",X"AC",X"B0",X"B0",X"B0",X"B4",X"B4",X"B4",X"B8",X"B8",X"C1",X"80",X"8D",X"96",
		X"9A",X"9F",X"A8",X"B0",X"B4",X"B4",X"B8",X"B8",X"BC",X"C1",X"C1",X"C5",X"CA",X"80",X"92",X"9A",
		X"A3",X"A8",X"AC",X"B4",X"B4",X"B8",X"B8",X"BC",X"BC",X"C1",X"C1",X"C5",X"CA",X"80",X"9F",X"A3",
		X"A8",X"AC",X"B0",X"B4",X"B4",X"B8",X"B8",X"BC",X"BC",X"C1",X"C1",X"C5",X"CA",X"80",X"A8",X"AC",
		X"B0",X"B0",X"B4",X"B8",X"BC",X"C1",X"C1",X"C1",X"C5",X"C5",X"CA",X"CE",X"D2",X"80",X"B7",X"BB",
		X"BF",X"BF",X"C7",X"CC",X"D0",X"D5",X"D9",X"DD",X"DD",X"E2",X"E6",X"EA",X"EA",X"80",X"BB",X"BF",
		X"C3",X"C7",X"CC",X"D5",X"D5",X"D9",X"D9",X"DD",X"E2",X"E6",X"E6",X"EA",X"EA",X"80",X"C3",X"C7",
		X"CF",X"D1",X"D5",X"D9",X"D9",X"DD",X"DD",X"E2",X"E2",X"E6",X"E6",X"EA",X"EA",X"80",X"CC",X"D0",
		X"D5",X"D5",X"D9",X"DD",X"E2",X"E6",X"E6",X"E6",X"EA",X"EA",X"EA",X"EA",X"EA",X"80",X"40",X"40",
		X"40",X"40",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"46",X"48",X"51",X"51",X"51",
		X"51",X"51",X"53",X"53",X"53",X"53",X"53",X"53",X"53",X"53",X"53",X"55",X"3A",X"CF",X"89",X"A7",
		X"20",X"0F",X"3A",X"3D",X"9B",X"FE",X"05",X"D0",X"21",X"F6",X"1D",X"CF",X"7E",X"23",X"66",X"6F",
		X"E9",X"AF",X"32",X"3D",X"9B",X"C9",X"00",X"1E",X"3A",X"1E",X"34",X"1F",X"0B",X"1E",X"01",X"1E",
		X"C9",X"CD",X"AB",X"1E",X"20",X"05",X"AF",X"32",X"3D",X"9B",X"C9",X"21",X"DE",X"1E",X"CD",X"7A",
		X"1E",X"11",X"30",X"B8",X"06",X"04",X"CD",X"7F",X"1E",X"11",X"DE",X"1E",X"21",X"00",X"B8",X"06",
		X"25",X"CD",X"B3",X"1E",X"CC",X"AB",X"1E",X"32",X"CF",X"89",X"21",X"DE",X"1E",X"11",X"A0",X"89",
		X"01",X"25",X"00",X"ED",X"B0",X"AF",X"32",X"3D",X"9B",X"C9",X"21",X"00",X"B8",X"11",X"A0",X"89",
		X"06",X"25",X"36",X"00",X"3E",X"08",X"32",X"40",X"B8",X"3C",X"32",X"40",X"B8",X"00",X"3E",X"08",
		X"32",X"40",X"B8",X"3E",X"0C",X"00",X"32",X"40",X"B8",X"3E",X"0D",X"32",X"40",X"B8",X"00",X"0E",
		X"01",X"ED",X"A0",X"3E",X"04",X"32",X"40",X"B8",X"10",X"D8",X"AF",X"32",X"3D",X"9B",X"C9",X"CD",
		X"77",X"1E",X"AF",X"32",X"3D",X"9B",X"C9",X"21",X"A0",X"89",X"11",X"00",X"B8",X"06",X"25",X"0E",
		X"01",X"ED",X"A0",X"3E",X"0E",X"32",X"40",X"B8",X"CD",X"A0",X"1E",X"3E",X"04",X"32",X"40",X"B8",
		X"3E",X"0A",X"32",X"40",X"B8",X"CD",X"A0",X"1E",X"3E",X"04",X"32",X"40",X"B8",X"10",X"E0",X"C9",
		X"C5",X"01",X"DB",X"24",X"0D",X"20",X"FD",X"10",X"FB",X"C1",X"C9",X"21",X"30",X"B8",X"11",X"03",
		X"1F",X"06",X"04",X"36",X"00",X"3E",X"08",X"32",X"40",X"B8",X"3C",X"32",X"40",X"B8",X"00",X"3E",
		X"08",X"32",X"40",X"B8",X"3E",X"0C",X"00",X"32",X"40",X"B8",X"3E",X"0D",X"32",X"40",X"B8",X"00",
		X"1A",X"AE",X"C0",X"23",X"13",X"3E",X"04",X"32",X"40",X"B8",X"10",X"D7",X"AF",X"C9",X"01",X"00",
		X"00",X"01",X"00",X"00",X"01",X"00",X"00",X"01",X"00",X"00",X"01",X"00",X"00",X"00",X"28",X"35",
		X"28",X"1C",X"35",X"1C",X"26",X"35",X"26",X"1A",X"35",X"1A",X"27",X"35",X"27",X"00",X"01",X"01",
		X"01",X"01",X"01",X"A5",X"C3",X"EE",X"18",X"21",X"00",X"00",X"F3",X"11",X"FE",X"1F",X"06",X"10",
		X"AF",X"86",X"2C",X"20",X"FC",X"24",X"10",X"F9",X"EB",X"BE",X"20",X"10",X"EB",X"1C",X"20",X"EE",
		X"3E",X"FF",X"32",X"00",X"8A",X"3A",X"00",X"8A",X"A7",X"20",X"FA",X"C9",X"3E",X"06",X"85",X"32",
		X"00",X"8A",X"18",X"F8",X"CD",X"77",X"1E",X"11",X"A0",X"89",X"21",X"00",X"B8",X"06",X"25",X"CD",
		X"B3",X"1E",X"3A",X"CF",X"89",X"A7",X"28",X"0B",X"21",X"57",X"1F",X"11",X"30",X"B8",X"06",X"04",
		X"CD",X"7F",X"1E",X"32",X"3D",X"9B",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"D9",X"11",X"BB");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
