library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_D8 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(8 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_D8 is
	type rom is array(0 to  511) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"0C",X"0C",X"0E",X"0E",X"0E",X"0E",X"0E",X"06",X"06",X"06",X"0E",X"0C",X"0C",X"08",X"0C",
		X"00",X"00",X"00",X"08",X"08",X"0C",X"0C",X"0C",X"0E",X"06",X"02",X"0A",X"0E",X"0E",X"07",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"0C",X"0C",X"04",X"06",X"0E",X"0E",X"87",X"03",X"02",
		X"00",X"00",X"00",X"00",X"00",X"08",X"0C",X"0E",X"06",X"0B",X"0D",X"87",X"E1",X"C0",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"0E",X"03",X"89",X"CF",X"F3",X"60",X"40",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"8F",X"D9",X"FC",X"FF",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"DF",X"F1",X"DF",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"20",X"FF",X"FC",X"D9",X"8F",X"0E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"40",X"60",X"F3",X"CF",X"89",X"03",X"0E",X"0C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"C0",X"E1",X"87",X"0D",X"0B",X"06",X"0E",X"0C",X"08",X"00",X"00",X"00",X"00",
		X"00",X"02",X"03",X"87",X"0E",X"0E",X"06",X"04",X"0C",X"0C",X"08",X"08",X"00",X"00",X"00",X"00",
		X"00",X"0E",X"07",X"0E",X"0E",X"0A",X"02",X"06",X"0E",X"0C",X"0C",X"0C",X"08",X"08",X"00",X"00",
		X"00",X"0C",X"08",X"0C",X"0C",X"0E",X"06",X"06",X"06",X"0E",X"0E",X"0E",X"0E",X"0E",X"0C",X"0C",
		X"00",X"08",X"00",X"08",X"0C",X"0C",X"06",X"06",X"0E",X"0F",X"0F",X"8F",X"8F",X"8F",X"87",X"03",
		X"00",X"00",X"00",X"00",X"08",X"0C",X"06",X"03",X"0B",X"8F",X"8F",X"CF",X"C7",X"C3",X"81",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0E",X"07",X"8F",X"8F",X"CF",X"C7",X"81",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0F",X"87",X"CF",X"EF",X"E7",X"C1",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"0F",X"CF",X"EF",X"FF",X"F7",X"E1",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"CF",X"FF",X"F7",X"FF",X"CF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"E1",X"F7",X"FF",X"EF",X"CF",X"0F",X"08",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"C1",X"E7",X"EF",X"CF",X"87",X"0F",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"81",X"C7",X"CF",X"8F",X"8F",X"07",X"0E",X"0C",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"81",X"C3",X"C7",X"CF",X"8F",X"8F",X"0B",X"03",X"06",X"0C",X"08",X"00",X"00",X"00",
		X"00",X"03",X"87",X"8F",X"8F",X"8F",X"0F",X"0F",X"0E",X"06",X"06",X"0C",X"0C",X"08",X"00",X"08",
		X"00",X"0A",X"00",X"80",X"01",X"48",X"28",X"02",X"00",X"22",X"08",X"21",X"08",X"82",X"00",X"04",
		X"04",X"00",X"80",X"02",X"20",X"04",X"00",X"94",X"00",X"48",X"00",X"84",X"01",X"02",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
