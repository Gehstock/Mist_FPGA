library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity char_rom1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of char_rom1 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"0F",X"0C",X"00",X"3F",X"00",X"0C",X"0F",X"0F",X"07",X"03",X"23",X"07",X"23",X"03",X"07",X"0F",
		X"06",X"00",X"00",X"00",X"08",X"0C",X"0E",X"0F",X"3F",X"1F",X"07",X"03",X"00",X"01",X"01",X"00",
		X"9F",X"FF",X"FF",X"FF",X"7F",X"3F",X"1F",X"0F",X"0C",X"0E",X"8F",X"CF",X"FF",X"EF",X"EF",X"FF",
		X"06",X"00",X"00",X"00",X"08",X"0C",X"0E",X"0F",X"0C",X"0E",X"07",X"03",X"00",X"01",X"01",X"00",
		X"9F",X"FF",X"FF",X"FF",X"7F",X"3F",X"1F",X"0F",X"3F",X"1F",X"8F",X"CF",X"FF",X"EF",X"EF",X"FF",
		X"00",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",
		X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"8F",X"CF",X"7F",X"4F",X"4F",X"0F",X"0F",X"0F",X"0F",X"0F",X"EF",X"EF",X"6F",X"0F",X"0F",X"0F",
		X"6F",X"FF",X"BF",X"9F",X"9F",X"4F",X"0F",X"0F",X"0F",X"2F",X"2F",X"2F",X"EF",X"EF",X"6F",X"0F",
		X"0F",X"1F",X"1F",X"1F",X"1F",X"1F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"6F",X"8F",X"8F",X"CF",X"7F",X"3F",X"1F",X"0F",X"4F",X"6F",X"2F",X"2F",X"2F",X"EF",X"CF",X"0F",
		X"7F",X"7F",X"CF",X"8F",X"FF",X"9F",X"0F",X"0F",X"8F",X"CF",X"6F",X"2F",X"2F",X"EF",X"6F",X"0F",
		X"8F",X"9F",X"9F",X"FF",X"FF",X"9F",X"0F",X"0F",X"0F",X"2F",X"2F",X"2F",X"EF",X"EF",X"6F",X"0F",
		X"CF",X"FF",X"3F",X"1F",X"DF",X"3F",X"0F",X"0F",X"0F",X"8F",X"EF",X"6F",X"0F",X"8F",X"6F",X"0F",
		X"8F",X"8F",X"EF",X"FF",X"8F",X"0F",X"0F",X"0F",X"0F",X"0F",X"2F",X"EF",X"EF",X"2F",X"2F",X"0F",
		X"7F",X"FF",X"8F",X"8F",X"CF",X"7F",X"1F",X"0F",X"0F",X"CF",X"6F",X"2F",X"2F",X"EF",X"CF",X"0F",
		X"7F",X"DF",X"8F",X"CF",X"FF",X"9F",X"0F",X"0F",X"0F",X"8F",X"8F",X"8F",X"8F",X"EF",X"6F",X"0F",
		X"6F",X"FF",X"9F",X"9F",X"FF",X"9F",X"0F",X"0F",X"0F",X"6F",X"EF",X"8F",X"0F",X"EF",X"6F",X"0F",
		X"8F",X"5F",X"9F",X"BF",X"FF",X"6F",X"0F",X"0F",X"CF",X"EF",X"AF",X"2F",X"2F",X"4F",X"2F",X"0F",
		X"8F",X"8F",X"CF",X"FF",X"BF",X"8F",X"0F",X"0F",X"0F",X"0F",X"0F",X"8F",X"EF",X"6F",X"0F",X"0F",
		X"CF",X"3F",X"0F",X"CF",X"FF",X"BF",X"8F",X"0F",X"0F",X"0F",X"CF",X"2F",X"AF",X"EF",X"CF",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"FF",X"FF",X"CF",X"AF",X"1F",X"0F",X"0F",X"2F",X"EF",X"EF",X"8F",X"8F",X"8F",X"EF",X"0F",
		X"6F",X"FF",X"9F",X"9F",X"FF",X"9F",X"0F",X"0F",X"CF",X"EF",X"2F",X"2F",X"2F",X"EF",X"6F",X"0F",
		X"5F",X"9F",X"9F",X"8F",X"4F",X"3F",X"1F",X"0F",X"8F",X"EF",X"4F",X"2F",X"2F",X"EF",X"CF",X"0F",
		X"8F",X"4F",X"3F",X"DF",X"FF",X"3F",X"0F",X"0F",X"2F",X"6F",X"CF",X"8F",X"0F",X"EF",X"EF",X"0F",
		X"0F",X"0F",X"0F",X"CF",X"FF",X"9F",X"0F",X"0F",X"0F",X"6F",X"2F",X"2F",X"2F",X"EF",X"6F",X"0F",
		X"0F",X"FF",X"3F",X"1F",X"FF",X"3F",X"0F",X"0F",X"6F",X"EF",X"0F",X"EF",X"0F",X"8F",X"6F",X"0F",
		X"CF",X"3F",X"0F",X"3F",X"FF",X"3F",X"0F",X"0F",X"0F",X"8F",X"EF",X"EF",X"8F",X"0F",X"EF",X"0F",
		X"CF",X"3F",X"1F",X"FF",X"1F",X"FF",X"CF",X"0F",X"0F",X"8F",X"EF",X"0F",X"8F",X"EF",X"0F",X"0F",
		X"CF",X"2F",X"1F",X"7F",X"EF",X"CF",X"0F",X"0F",X"0F",X"0F",X"8F",X"EF",X"6F",X"0F",X"0F",X"0F",
		X"8F",X"6F",X"1F",X"0F",X"FF",X"FF",X"8F",X"0F",X"0F",X"0F",X"8F",X"4F",X"EF",X"EF",X"0F",X"0F",
		X"0F",X"0E",X"0E",X"0E",X"0E",X"0E",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"09",X"09",X"0F",X"0F",X"0F",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"08",X"00",X"07",X"07",X"03",X"08",X"0E",X"0F",X"0F",X"03",X"09",X"0D",X"0D",X"01",X"03",X"0F",
		X"07",X"03",X"08",X"0B",X"0B",X"0F",X"0F",X"0F",X"0F",X"0F",X"01",X"01",X"09",X"0F",X"0F",X"0F",
		X"09",X"00",X"04",X"06",X"06",X"0B",X"0F",X"0F",X"0F",X"0D",X"0D",X"0D",X"01",X"01",X"09",X"0F",
		X"09",X"01",X"06",X"06",X"06",X"0B",X"0F",X"0F",X"0F",X"03",X"01",X"0D",X"0D",X"0D",X"0B",X"0F",
		X"0F",X"03",X"00",X"06",X"0B",X"0D",X"0E",X"0F",X"07",X"07",X"07",X"01",X"01",X"07",X"07",X"0F",
		X"07",X"02",X"02",X"02",X"02",X"08",X"0F",X"0F",X"03",X"01",X"0D",X"0D",X"0D",X"09",X"0B",X"0F",
		X"07",X"06",X"06",X"0A",X"08",X"0C",X"0E",X"0F",X"03",X"01",X"0D",X"0D",X"0D",X"01",X"03",X"0F",
		X"07",X"03",X"01",X"02",X"03",X"0B",X"0D",X"0F",X"0F",X"0F",X"0F",X"0F",X"01",X"09",X"0F",X"0F",
		X"09",X"01",X"06",X"04",X"00",X"09",X"0F",X"0F",X"0F",X"03",X"05",X"05",X"0D",X"05",X"03",X"0F",
		X"08",X"00",X"06",X"06",X"02",X"08",X"0D",X"0F",X"0F",X"07",X"03",X"0B",X"0D",X"0D",X"0D",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"00",X"00",X"03",X"05",X"0E",X"0F",X"0F",X"0D",X"01",X"01",X"07",X"07",X"07",X"01",X"0F",
		X"09",X"00",X"06",X"06",X"00",X"06",X"0F",X"0F",X"03",X"01",X"0D",X"0D",X"0D",X"01",X"09",X"0F",
		X"09",X"07",X"07",X"03",X"08",X"0C",X"0E",X"0F",X"0B",X"09",X"0D",X"0D",X"0D",X"01",X"03",X"0F",
		X"08",X"08",X"03",X"07",X"00",X"06",X"0F",X"0F",X"07",X"03",X"09",X"0D",X"0D",X"01",X"09",X"0F",
		X"07",X"06",X"06",X"00",X"00",X"06",X"0F",X"0F",X"0F",X"0D",X"0D",X"0D",X"01",X"01",X"09",X"0F",
		X"07",X"06",X"06",X"00",X"00",X"06",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"03",X"01",X"09",X"0F",
		X"0A",X"06",X"06",X"07",X"0B",X"0C",X"0E",X"0F",X"07",X"01",X"0B",X"0D",X"0D",X"01",X"03",X"0F",
		X"03",X"00",X"0C",X"0E",X"02",X"0C",X"0F",X"0F",X"0F",X"07",X"01",X"09",X"0F",X"07",X"09",X"0F",
		X"07",X"07",X"01",X"00",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"0D",X"01",X"01",X"0D",X"0D",X"0F",
		X"07",X"03",X"00",X"06",X"07",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"03",X"09",X"0D",X"09",X"0F",
		X"07",X"0B",X"0C",X"02",X"00",X"0C",X"0F",X"0F",X"0D",X"09",X"03",X"07",X"0F",X"01",X"01",X"0F",
		X"0F",X"0F",X"0F",X"03",X"00",X"06",X"0F",X"0F",X"0F",X"09",X"0D",X"0D",X"0D",X"01",X"09",X"0F",
		X"0F",X"00",X"0C",X"0E",X"00",X"0C",X"0F",X"0F",X"09",X"01",X"0F",X"01",X"0F",X"07",X"09",X"0F",
		X"03",X"0C",X"0F",X"0C",X"00",X"0C",X"0F",X"0F",X"0F",X"07",X"01",X"01",X"07",X"0F",X"01",X"0F",
		X"08",X"00",X"07",X"07",X"03",X"08",X"0E",X"0F",X"0F",X"03",X"09",X"0D",X"0D",X"01",X"03",X"0F",
		X"08",X"02",X"07",X"03",X"00",X"06",X"0F",X"0F",X"0F",X"07",X"07",X"07",X"07",X"01",X"09",X"0F",
		X"08",X"00",X"07",X"07",X"03",X"08",X"0E",X"0F",X"0D",X"01",X"03",X"05",X"0D",X"01",X"03",X"0F",
		X"09",X"00",X"06",X"06",X"00",X"06",X"0F",X"0F",X"0F",X"09",X"01",X"07",X"0F",X"01",X"09",X"0F",
		X"07",X"0A",X"06",X"04",X"00",X"09",X"0F",X"0F",X"03",X"01",X"05",X"0D",X"0D",X"0B",X"0D",X"0F",
		X"07",X"07",X"03",X"00",X"04",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"01",X"09",X"0F",X"0F",
		X"03",X"0C",X"0F",X"03",X"00",X"04",X"07",X"0F",X"0F",X"0F",X"03",X"0D",X"05",X"01",X"03",X"0F",
		X"07",X"09",X"0E",X"0F",X"00",X"00",X"07",X"0F",X"0F",X"0F",X"07",X"0B",X"01",X"01",X"0F",X"0F",
		X"03",X"0C",X"0E",X"00",X"0E",X"00",X"03",X"0F",X"0F",X"07",X"01",X"0F",X"07",X"01",X"0F",X"0F",
		X"07",X"0B",X"0D",X"08",X"01",X"07",X"0F",X"0F",X"0F",X"0D",X"01",X"03",X"07",X"0B",X"0D",X"0F",
		X"03",X"0D",X"0E",X"08",X"01",X"03",X"0F",X"0F",X"0F",X"0F",X"07",X"01",X"09",X"0F",X"0F",X"0F",
		X"07",X"03",X"01",X"04",X"06",X"03",X"0F",X"0F",X"0F",X"09",X"0D",X"0D",X"05",X"01",X"09",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"09",X"09",X"0F",X"0F",X"0F",
		X"0F",X"0C",X"0B",X"05",X"05",X"06",X"0B",X"0C",X"0F",X"07",X"0B",X"05",X"05",X"0D",X"0B",X"07",
		X"0F",X"0F",X"0F",X"0F",X"08",X"09",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"0F",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"1F",X"0F",X"0F",X"0F",X"3F",X"3F",X"3F",X"3F",X"EF",X"FF",X"7F",X"3F",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"0F",X"8F",X"CF",X"EF",X"FF",X"7F",X"3F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"8F",X"CF",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"3F",X"2F",X"3F",X"3F",X"1F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"3F",X"3F",X"3F",X"0F",X"0F",X"0F",X"1F",X"3F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"1F",X"3F",X"3F",X"3F",X"1F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"1F",X"3F",X"3F",X"3F",X"3F",X"3F",X"1F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"1F",X"3F",X"3F",X"3F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"3F",X"3F",X"1F",X"1F",X"3F",X"3F",X"3F",X"3F",
		X"1F",X"1F",X"1F",X"0F",X"0F",X"0F",X"0F",X"0F",X"BF",X"BF",X"BF",X"0F",X"0F",X"0F",X"1F",X"3F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"2F",X"2F",X"2F",X"2F",X"1F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"1F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"7F",X"FF",X"EF",X"EF",X"FF",X"FF",X"FF",X"FF",X"0F",X"0F",X"0F",X"0F",X"CF",X"CF",X"CF",X"CF",
		X"FF",X"FF",X"FF",X"1F",X"0F",X"1F",X"1F",X"3F",X"0F",X"8F",X"CF",X"CF",X"CF",X"CF",X"8F",X"8F",
		X"0F",X"0F",X"0F",X"FF",X"FF",X"FF",X"0F",X"0F",X"CF",X"4F",X"CF",X"CF",X"8F",X"0F",X"0F",X"0F",
		X"FF",X"FF",X"FF",X"0F",X"0F",X"FF",X"FF",X"FF",X"CF",X"CF",X"CF",X"0F",X"0F",X"0F",X"8F",X"CF",
		X"0F",X"0F",X"FF",X"FF",X"FF",X"0F",X"0F",X"8F",X"0F",X"0F",X"CF",X"CF",X"CF",X"0F",X"0F",X"0F",
		X"FF",X"FF",X"6F",X"2F",X"2F",X"BF",X"9F",X"9F",X"CF",X"8F",X"CF",X"4F",X"4F",X"4F",X"CF",X"8F",
		X"8F",X"FF",X"FF",X"FF",X"0F",X"0F",X"0F",X"FF",X"0F",X"CF",X"CF",X"CF",X"0F",X"0F",X"4F",X"CF",
		X"0F",X"0F",X"8F",X"FF",X"FF",X"FF",X"0F",X"0F",X"0F",X"0F",X"0F",X"CF",X"CF",X"CF",X"0F",X"0F",
		X"FF",X"FF",X"FF",X"0F",X"0F",X"FF",X"FF",X"FF",X"CF",X"CF",X"CF",X"0F",X"0F",X"CF",X"CF",X"CF",
		X"5F",X"AF",X"AF",X"FF",X"0F",X"FF",X"0F",X"0F",X"4F",X"4F",X"4F",X"4F",X"8F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"FF",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"8F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"1F",X"0F",X"0F",X"0F",X"3F",X"3F",X"3F",X"3F",X"EF",X"FF",X"7F",X"3F",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"0F",X"8F",X"CF",X"EF",X"FF",X"7F",X"3F",X"1F",X"1F",X"1F",X"0F",X"0F",X"0F",X"8F",X"CF",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"08",X"0C",X"0E",X"0F",X"0F",X"0F",X"0F",
		X"30",X"00",X"00",X"00",X"00",X"00",X"0C",X"0E",X"F7",X"F3",X"71",X"30",X"10",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"13",X"81",X"0F",X"CF",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"8F",X"EF",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"FF",X"7F",X"1F",X"07",X"07",X"07",X"0F",X"0F",X"8F",X"CF",X"CF",X"4F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"CF",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"8F",X"8F",
		X"0F",X"8F",X"8F",X"8F",X"CF",X"CF",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"CF",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"8F",X"8F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"1E",X"0F",X"3C",X"3C",X"1E",X"1E",X"0F",X"0F",
		X"3C",X"1E",X"1E",X"1E",X"0F",X"0F",X"0F",X"0F",X"B2",X"D0",X"D1",X"E0",X"E0",X"F0",X"F0",X"78",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"3F",X"3E",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"1E",X"1E",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"F3",X"7B",X"79",X"79",X"3C",X"3C",X"2C",X"0F",
		X"3F",X"2E",X"2E",X"0F",X"1E",X"1E",X"0F",X"0F",X"77",X"7F",X"FF",X"EE",X"FF",X"FF",X"F7",X"F7",
		X"7F",X"FF",X"EF",X"EF",X"FF",X"FF",X"FF",X"FF",X"0F",X"0F",X"0F",X"0F",X"CF",X"CF",X"CF",X"CF",
		X"FF",X"FF",X"FF",X"1F",X"0F",X"1F",X"1F",X"3F",X"0F",X"8F",X"CF",X"CF",X"CF",X"CF",X"8F",X"8F",
		X"43",X"43",X"61",X"21",X"21",X"29",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"FF",X"FF",X"FF",X"7F",X"37",X"07",X"07",X"03",X"8F",X"CF",X"CF",X"CF",X"EF",X"EF",X"6F",X"3F",
		X"0F",X"0F",X"0F",X"0F",X"CF",X"FF",X"FF",X"FF",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"8F",X"8F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"3F",X"2F",X"3F",X"3F",X"1F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"3F",X"3F",X"3F",X"0F",X"0F",X"0F",X"1F",X"3F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"1E",X"1E",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"00",X"08",X"08",X"08",X"0C",X"0E",
		X"0C",X"0E",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"01",X"08",X"0C",X"0E",X"0E",X"0F",
		X"5A",X"FC",X"11",X"E0",X"F0",X"2D",X"1E",X"0F",X"E1",X"78",X"CB",X"33",X"C0",X"F0",X"5A",X"1E",
		X"D1",X"E0",X"E0",X"E0",X"F8",X"F0",X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",X"74",X"74",X"F0",X"F0",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"1F",X"FF",X"D1",X"0F",X"0F",X"0F",X"0F",X"0F",X"FF",X"F0",X"F0",
		X"00",X"10",X"21",X"43",X"0F",X"0F",X"0F",X"0F",X"E7",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"00",X"00",X"10",X"21",X"42",X"84",X"18",X"00",X"73",X"E7",X"CF",X"FF",X"31",X"C3",X"CF",X"C7",
		X"73",X"73",X"E6",X"4C",X"4C",X"80",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"10",X"31",
		X"0F",X"0F",X"0F",X"FF",X"FF",X"FF",X"0F",X"0F",X"CF",X"4F",X"CF",X"CF",X"8F",X"0F",X"0F",X"0F",
		X"FF",X"FF",X"FF",X"0F",X"0F",X"FF",X"FF",X"FF",X"CF",X"CF",X"CF",X"0F",X"0F",X"0F",X"8F",X"CF",
		X"0F",X"0F",X"FF",X"FF",X"FF",X"0F",X"0F",X"8F",X"0F",X"0F",X"CF",X"CF",X"CF",X"0F",X"0F",X"0F",
		X"FF",X"FF",X"6F",X"2F",X"2F",X"BF",X"9F",X"9F",X"CF",X"8F",X"CF",X"4F",X"4F",X"4F",X"CF",X"8F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"3C",X"1E",X"1E",X"1E",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"32",X"32",X"32",X"19",X"19",X"08",X"0C",X"0C",
		X"0C",X"0E",X"0F",X"1C",X"0C",X"0E",X"0E",X"0E",X"31",X"31",X"10",X"08",X"80",X"84",X"62",X"73",
		X"00",X"08",X"84",X"42",X"31",X"10",X"08",X"0C",X"E6",X"71",X"10",X"00",X"00",X"88",X"C4",X"62",
		X"08",X"0C",X"0E",X"00",X"00",X"00",X"24",X"10",X"B7",X"53",X"21",X"10",X"00",X"00",X"00",X"08",
		X"00",X"00",X"00",X"84",X"42",X"21",X"10",X"10",X"21",X"21",X"10",X"10",X"10",X"88",X"6E",X"3F",
		X"E0",X"F0",X"F0",X"F0",X"FE",X"00",X"F0",X"F0",X"FF",X"07",X"07",X"77",X"B3",X"FF",X"33",X"D1",
		X"77",X"B3",X"B3",X"B3",X"D1",X"D1",X"D1",X"E0",X"8F",X"CF",X"CF",X"CF",X"EF",X"EF",X"EF",X"FF",
		X"0E",X"0E",X"0E",X"0E",X"1F",X"7F",X"F7",X"F7",X"10",X"10",X"00",X"07",X"0C",X"00",X"88",X"88",
		X"00",X"00",X"08",X"08",X"08",X"0C",X"0C",X"0C",X"42",X"00",X"00",X"00",X"00",X"00",X"10",X"10",
		X"0F",X"0F",X"0F",X"CF",X"0F",X"0E",X"08",X"00",X"0F",X"0F",X"3F",X"7F",X"7F",X"F7",X"B7",X"B7",
		X"00",X"00",X"70",X"73",X"73",X"E7",X"CF",X"8F",X"73",X"87",X"8F",X"8F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"1F",X"3F",X"3F",X"3F",X"3F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"1F",X"3F",X"3F",X"3F",X"3F",X"3F",X"1F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"1F",X"3F",X"3F",X"3F",X"0F",X"0F",X"0F",X"0F",
		X"1D",X"1D",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"11",X"08",X"0C",X"0C",X"0E",X"0E",X"0F",X"0F",
		X"32",X"11",X"11",X"00",X"00",X"00",X"2A",X"2B",X"86",X"C3",X"E1",X"F8",X"74",X"74",X"32",X"11",
		X"88",X"8C",X"8C",X"CE",X"CF",X"E7",X"77",X"73",X"62",X"31",X"10",X"10",X"00",X"08",X"08",X"8C",
		X"00",X"88",X"CC",X"E6",X"73",X"31",X"10",X"00",X"73",X"31",X"10",X"10",X"10",X"00",X"88",X"C4",
		X"00",X"88",X"CE",X"E7",X"73",X"31",X"10",X"00",X"87",X"87",X"43",X"0F",X"0F",X"CF",X"EF",X"F7",
		X"FF",X"FF",X"FF",X"FF",X"77",X"3B",X"1D",X"0E",X"FC",X"FC",X"FC",X"FE",X"FF",X"FF",X"FE",X"FF",
		X"E0",X"2C",X"0E",X"0F",X"0F",X"8F",X"CB",X"E1",X"33",X"00",X"00",X"00",X"0C",X"4F",X"3B",X"08",
		X"00",X"FF",X"0F",X"CF",X"FF",X"FF",X"FC",X"CC",X"00",X"8C",X"0F",X"0F",X"CF",X"CF",X"EF",X"E1",
		X"00",X"31",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"F1",X"10",X"00",X"00",X"00",
		X"7F",X"0F",X"B7",X"6E",X"00",X"00",X"00",X"00",X"0F",X"7F",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"30",X"F7",X"7F",X"00",X"00",X"00",X"10",X"43",X"0F",X"8F",X"8F",
		X"0F",X"8F",X"8F",X"8F",X"8F",X"CF",X"CE",X"88",X"0F",X"0F",X"0F",X"0F",X"0E",X"08",X"00",X"00",
		X"8F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"8F",X"FF",X"FF",X"FF",X"0F",X"0F",X"0F",X"FF",X"0F",X"CF",X"CF",X"CF",X"0F",X"0F",X"4F",X"CF",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0C",X"0E",X"0E",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"08",X"0C",X"0E",X"0E",X"0F",X"0F",X"0F",X"0F",X"74",X"32",X"32",X"11",X"00",X"00",X"08",X"0C",
		X"F0",X"F8",X"74",X"32",X"32",X"11",X"00",X"08",X"1D",X"1D",X"87",X"C3",X"E1",X"E1",X"F8",X"F8",
		X"00",X"00",X"08",X"08",X"8C",X"8E",X"CF",X"EF",X"F7",X"F7",X"73",X"73",X"53",X"31",X"21",X"29",
		X"43",X"43",X"A9",X"EF",X"F7",X"73",X"31",X"10",X"FF",X"7F",X"3F",X"1F",X"0F",X"8F",X"CF",X"EF",
		X"86",X"C2",X"E0",X"F0",X"78",X"F8",X"BC",X"9E",X"11",X"11",X"00",X"00",X"00",X"80",X"C0",X"E0",
		X"00",X"00",X"08",X"08",X"08",X"0C",X"0C",X"0C",X"FC",X"32",X"11",X"00",X"00",X"00",X"22",X"11",
		X"33",X"00",X"00",X"00",X"08",X"8E",X"47",X"23",X"F8",X"76",X"11",X"00",X"00",X"00",X"00",X"0C",
		X"F7",X"70",X"00",X"00",X"00",X"08",X"0E",X"D3",X"FF",X"F7",X"71",X"10",X"00",X"00",X"00",X"88",
		X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"FF",X"FF",X"00",X"00",X"0C",X"0F",X"0F",X"0F",X"8F",X"FF",
		X"00",X"FF",X"FF",X"FF",X"F0",X"00",X"00",X"00",X"00",X"EE",X"FF",X"FF",X"F0",X"00",X"00",X"00",
		X"FF",X"FF",X"1E",X"1E",X"0F",X"0F",X"0F",X"0F",X"FF",X"BC",X"B4",X"B4",X"D2",X"D2",X"69",X"69",
		X"FD",X"FD",X"EF",X"0F",X"0F",X"0F",X"0F",X"0F",X"F8",X"CB",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"1E",X"7C",X"F6",X"F6",X"FB",X"FB",X"1F",X"7F",X"F3",X"F3",X"F1",X"F1",X"F0",X"F0",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0E",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"11",X"11",X"19",X"08",X"0C",X"0E",X"0F",X"0F",
		X"11",X"11",X"00",X"00",X"08",X"0C",X"0C",X"0E",X"F0",X"F0",X"F8",X"74",X"56",X"23",X"23",X"23",
		X"C3",X"E1",X"E1",X"F0",X"F8",X"74",X"74",X"32",X"0F",X"0F",X"0F",X"0F",X"87",X"87",X"C3",X"E1",
		X"3C",X"1E",X"0F",X"0F",X"0F",X"0F",X"0F",X"87",X"87",X"87",X"C3",X"4B",X"2D",X"0F",X"0F",X"0F",
		X"0F",X"87",X"C3",X"E1",X"F0",X"F0",X"F0",X"78",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"87",
		X"00",X"0C",X"86",X"87",X"87",X"4B",X"0F",X"0F",X"00",X"00",X"00",X"00",X"08",X"0C",X"0E",X"0F",
		X"80",X"68",X"E8",X"BC",X"56",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"00",
		X"0F",X"CF",X"67",X"3B",X"0C",X"0F",X"E1",X"E1",X"0F",X"0F",X"0F",X"8F",X"EF",X"33",X"1D",X"4A",
		X"0F",X"CF",X"77",X"08",X"0E",X"87",X"D2",X"E1",X"0F",X"0F",X"0F",X"EF",X"33",X"08",X"0E",X"0F",
		X"FF",X"FF",X"FF",X"11",X"0E",X"0F",X"0F",X"0F",X"2D",X"2D",X"9E",X"9E",X"07",X"0B",X"0F",X"0F",
		X"FC",X"FC",X"FE",X"0F",X"0F",X"0E",X"1E",X"0F",X"F8",X"F8",X"F4",X"F4",X"0F",X"01",X"C4",X"F4",
		X"F8",X"F8",X"F4",X"F4",X"F2",X"F2",X"F9",X"F9",X"F3",X"F1",X"F1",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"CF",X"E1",X"E1",X"F0",X"F0",X"F0",X"F0",X"F0",X"19",X"1D",X"1D",X"0C",X"0E",X"86",X"86",X"C3",
		X"83",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"FF",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"3F",X"FF",
		X"F7",X"F7",X"F3",X"73",X"73",X"71",X"21",X"21",X"FF",X"FF",X"FF",X"FF",X"FF",X"CF",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"1F",X"7F",X"FF",X"0F",X"0F",X"0F",X"2F",X"6F",X"FF",X"FF",X"FF",
		X"3C",X"3C",X"1E",X"0F",X"8F",X"8F",X"47",X"07",X"87",X"87",X"87",X"C3",X"C3",X"4B",X"2D",X"2D",
		X"0F",X"87",X"C3",X"C3",X"E1",X"F0",X"F0",X"78",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0C",X"0E",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"08",X"0C",X"0E",X"0F",X"0F",
		X"4B",X"87",X"E1",X"D2",X"F0",X"F0",X"B4",X"B4",X"77",X"77",X"77",X"3B",X"3B",X"3B",X"95",X"4A",
		X"3B",X"3B",X"1D",X"1D",X"95",X"86",X"86",X"C2",X"8F",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0E",X"0F",X"0F",X"0F",X"0F",X"8F",X"CF",X"77",X"33",X"08",X"0E",X"1E",X"0F",X"0F",X"0F",X"0F",
		X"2D",X"2D",X"1E",X"1E",X"8F",X"EF",X"33",X"08",X"78",X"78",X"3C",X"3C",X"96",X"96",X"8F",X"EF",
		X"78",X"78",X"3C",X"3C",X"96",X"96",X"4B",X"4B",X"D1",X"C0",X"C0",X"E0",X"E0",X"E0",X"F0",X"F0",
		X"E0",X"E0",X"E0",X"F0",X"3C",X"1F",X"00",X"E0",X"0F",X"0F",X"07",X"07",X"77",X"FF",X"FF",X"11",
		X"77",X"33",X"3B",X"3B",X"19",X"95",X"D1",X"D1",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"77",X"77",X"CF",X"CF",X"CF",X"EF",X"EF",X"EF",X"FF",X"FF",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"3F",X"FF",X"FF",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"8F",X"8F",
		X"0F",X"8F",X"8F",X"CF",X"8F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"5F",X"AF",X"AF",X"FF",X"0F",X"FF",X"0F",X"0F",X"4F",X"4F",X"4F",X"4F",X"8F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"3F",X"3F",X"1F",X"1F",X"3F",X"3F",X"3F",X"3F",
		X"0F",X"0F",X"8F",X"FF",X"FF",X"FF",X"0F",X"0F",X"0F",X"0F",X"0F",X"CF",X"CF",X"CF",X"0F",X"0F",
		X"1F",X"1F",X"1F",X"0F",X"0F",X"0F",X"0F",X"0F",X"BF",X"BF",X"BF",X"0F",X"0F",X"0F",X"1F",X"3F",
		X"0E",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"08",X"0C",X"0E",X"0F",X"0F",X"0F",
		X"73",X"31",X"10",X"00",X"00",X"00",X"08",X"0C",X"FF",X"FF",X"FF",X"F3",X"31",X"10",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"CF",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"88",X"EE",X"EF",X"EF",X"FF",X"FF",X"30",X"10",X"10",X"10",X"08",X"0C",X"0F",X"0F",
		X"8E",X"FF",X"33",X"0C",X"86",X"87",X"4B",X"0F",X"77",X"FF",X"FF",X"FF",X"33",X"91",X"59",X"59",
		X"33",X"91",X"91",X"91",X"C0",X"C0",X"C0",X"E0",X"FF",X"FF",X"FF",X"FF",X"7F",X"0F",X"0F",X"07",
		X"FF",X"FF",X"FF",X"FF",X"77",X"77",X"77",X"33",X"CF",X"CF",X"CF",X"EF",X"EF",X"EF",X"FF",X"FF",
		X"6F",X"0F",X"0F",X"0F",X"FF",X"FF",X"FF",X"FF",X"0F",X"0F",X"0F",X"0F",X"0F",X"8F",X"8F",X"8F",
		X"0F",X"8F",X"8F",X"8F",X"CF",X"CF",X"CF",X"EF",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"FF",X"FF",X"FF",X"0F",X"0F",X"FF",X"FF",X"FF",X"CF",X"CF",X"CF",X"0F",X"0F",X"CF",X"CF",X"CF",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"2F",X"2F",X"2F",X"2F",X"1F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"1F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"FF",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"8F",
		X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",
		X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"0F",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"0F",X"70",X"70",X"70",X"70",X"70",X"70",X"00",X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"0F",X"0F",X"B3",X"B3",X"B3",X"B3",X"B3",X"B3",X"0F",X"0F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"B3",X"B3",X"B3",X"B3",X"B3",X"B3",X"B3",X"B3",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"08",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",
		X"0F",X"87",X"C2",X"D3",X"D3",X"C3",X"80",X"00",X"0F",X"1E",X"30",X"B8",X"B8",X"3C",X"10",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"70",X"70",X"70",X"07",X"03",X"30",X"30",X"30",
		X"F0",X"F0",X"F0",X"E0",X"E1",X"E1",X"E1",X"E1",X"F0",X"F0",X"F0",X"00",X"00",X"78",X"3C",X"1E",
		X"F0",X"F0",X"F0",X"30",X"10",X"C0",X"E0",X"F0",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"61",X"01",
		X"E1",X"D3",X"3F",X"7E",X"FC",X"F0",X"F0",X"F0",X"ED",X"E9",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"30",X"30",X"00",X"70",X"70",X"70",X"07",X"B7",
		X"CE",X"CE",X"CE",X"CE",X"CC",X"88",X"11",X"33",X"70",X"74",X"33",X"00",X"00",X"0F",X"FF",X"FF",
		X"30",X"11",X"88",X"CC",X"CE",X"CE",X"CE",X"CE",X"F0",X"FF",X"0F",X"00",X"00",X"33",X"74",X"70",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"01",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",
		X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",
		X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",
		X"B3",X"B3",X"B3",X"B3",X"B3",X"B3",X"0F",X"0F",X"B3",X"B3",X"B3",X"B3",X"B3",X"B3",X"0F",X"0F",
		X"B3",X"B3",X"B3",X"B3",X"B3",X"B3",X"B3",X"B3",X"B3",X"B3",X"B3",X"B3",X"B3",X"B3",X"B3",X"B3",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",
		X"F0",X"F0",X"F0",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"F0",X"F0",X"F0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"D0",X"B0",X"F0",X"70",X"70",X"70",X"00",X"00",X"F0",X"F0",X"F0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",
		X"F0",X"F0",X"F0",X"00",X"10",X"E0",X"E0",X"E8",X"F0",X"F0",X"F0",X"70",X"70",X"70",X"70",X"70",
		X"F0",X"F0",X"F0",X"0F",X"0F",X"E1",X"E1",X"E1",X"3F",X"3F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"70",X"70",X"70",X"70",X"00",X"00",X"70",X"FF",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"F0",X"FF",
		X"8F",X"F7",X"77",X"70",X"70",X"70",X"70",X"70",X"0F",X"FF",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"E2",X"C6",X"8C",X"00",X"00",X"0F",X"FF",X"FF",X"36",X"36",X"36",X"36",X"32",X"10",X"88",X"CC",
		X"F0",X"FF",X"0F",X"00",X"00",X"8C",X"C6",X"E2",X"C0",X"88",X"10",X"32",X"36",X"36",X"36",X"36",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E1",X"F1",X"F1",X"E1",X"E1",X"F1",X"F1",X"E1",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E1",X"E1",X"F1",X"F1",X"F1",X"F1",X"E1",X"E1",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E1",X"E1",X"E1",X"E0",X"E0",X"E1",X"E1",X"E1",
		X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"0F",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"01",
		X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"38",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"30",X"30",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"E1",X"E1",X"E1",X"10",X"00",X"F0",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"87",X"C3",X"E1",X"F0",
		X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"F0",X"FF",X"E1",X"E1",X"E1",X"E1",X"01",X"10",X"F0",X"FF",
		X"0F",X"FF",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"EF",X"EF",X"E1",X"E1",X"E1",X"E1",X"E1",
		X"C3",X"C3",X"C3",X"C3",X"C3",X"C3",X"C3",X"C3",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",
		X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"78",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",
		X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"07",X"0F",X"0F",X"00",X"00",X"0F",X"0F",X"07",
		X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"3F",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"CF",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"9E",X"9E",X"9E",X"9E",X"9E",X"8F",X"8F",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"0F",X"FF",
		X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"00",X"E1",X"E1",X"F1",X"F1",X"F1",X"E1",X"E1",X"01",
		X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"E1",X"E1",X"F1",X"F1",X"F1",X"F1",X"E1",X"E1",
		X"0F",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"0F",X"E1",X"E1",X"F1",X"F1",X"F1",X"E1",X"E1",
		X"D0",X"D0",X"D0",X"C1",X"E0",X"E0",X"E0",X"E0",X"F0",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"F0",
		X"70",X"70",X"70",X"60",X"50",X"21",X"D2",X"C0",X"D0",X"A1",X"52",X"B4",X"78",X"F0",X"F0",X"00",
		X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"E1",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",
		X"C3",X"D0",X"24",X"52",X"61",X"70",X"70",X"70",X"0F",X"F0",X"F0",X"70",X"B0",X"58",X"A4",X"D2",
		X"B0",X"B0",X"B0",X"B0",X"D0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"F0",
		X"F0",X"F0",X"F1",X"F2",X"B0",X"B0",X"B0",X"B0",X"F0",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"00",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"01",
		X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",
		X"0F",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"0F",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",
		X"0E",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"07",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"0F",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"0F",X"FF",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"08",X"08",X"0B",X"0F",
		X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"1F",X"70",X"70",X"70",X"70",X"70",X"70",X"00",X"CF",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",
		X"08",X"00",X"05",X"06",X"02",X"0B",X"0F",X"0F",X"03",X"07",X"0B",X"0B",X"03",X"07",X"0F",X"0B",
		X"E0",X"F1",X"F1",X"F0",X"E0",X"F1",X"F1",X"F0",X"70",X"70",X"70",X"F0",X"70",X"70",X"70",X"F0",
		X"E0",X"E0",X"68",X"58",X"58",X"1C",X"2D",X"FF",X"F0",X"F0",X"00",X"F0",X"F0",X"F0",X"0F",X"FF",
		X"78",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"E1",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",
		X"B0",X"58",X"A4",X"D2",X"D0",X"A1",X"52",X"B4",X"D0",X"A1",X"52",X"B4",X"B0",X"58",X"A4",X"D2",
		X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"70",X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"F0",X"F2",X"F2",X"F2",X"F2",X"F4",X"F8",X"F0",X"F0",
		X"F0",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F8",X"F4",X"F2",X"F2",X"F2",X"F2",
		X"F0",X"C3",X"B4",X"B1",X"91",X"80",X"C0",X"F0",X"F0",X"3C",X"1E",X"9E",X"DA",X"D2",X"34",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"0F",X"0F",X"0F",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0B",X"03",X"03",X"0B",X"0F",X"0F",
		X"6F",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"6F",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"0F",X"FF",X"E0",X"E0",X"E0",X"E0",X"E0",X"0E",X"0E",X"EE",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"3F",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"CF",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",
		X"05",X"0E",X"00",X"00",X"0F",X"0F",X"0F",X"08",X"0F",X"0B",X"03",X"03",X"0B",X"0F",X"0B",X"03",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"07",X"02",X"0F",X"0F",X"0F",X"0F",X"0F",X"0B",X"03",X"07",
		X"D3",X"D3",X"D3",X"1F",X"1F",X"97",X"97",X"97",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",
		X"B0",X"58",X"A4",X"D2",X"E1",X"F0",X"F0",X"00",X"E1",X"E1",X"E1",X"61",X"A1",X"49",X"B4",X"30",
		X"78",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"70",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",
		X"0F",X"F0",X"F0",X"E0",X"D0",X"A1",X"52",X"B4",X"3C",X"B0",X"43",X"A5",X"69",X"E1",X"E1",X"E1",
		X"70",X"70",X"70",X"70",X"70",X"70",X"60",X"11",X"F0",X"F0",X"F0",X"C0",X"80",X"30",X"34",X"3C",
		X"73",X"71",X"70",X"70",X"70",X"70",X"70",X"70",X"3C",X"9E",X"CF",X"E7",X"F3",X"F0",X"F0",X"F0",
		X"30",X"30",X"30",X"30",X"30",X"30",X"00",X"00",X"E3",X"E3",X"E3",X"E3",X"E3",X"E3",X"01",X"01",
		X"0F",X"73",X"30",X"30",X"30",X"30",X"30",X"30",X"0F",X"EF",X"E3",X"E3",X"E3",X"E3",X"E3",X"E3",
		X"0F",X"33",X"30",X"30",X"30",X"30",X"00",X"00",X"0F",X"FF",X"F0",X"F0",X"F0",X"F0",X"00",X"00",
		X"C7",X"73",X"31",X"10",X"10",X"00",X"00",X"70",X"0F",X"FF",X"FF",X"F0",X"F0",X"00",X"00",X"F0",
		X"0F",X"FF",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"0F",X"FF",X"F0",X"F0",X"F0",X"F0",X"00",X"00",
		X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"E3",X"E3",X"E3",X"E3",X"E3",X"E3",X"E3",X"E3",
		X"97",X"97",X"97",X"D3",X"D3",X"D3",X"1F",X"FF",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",
		X"3F",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"8F",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"01",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F3",X"F3",X"30",X"B0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"C7",X"CF",
		X"30",X"30",X"30",X"30",X"30",X"30",X"00",X"00",X"E1",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",
		X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",
		X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E1",
		X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",
		X"78",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",
		X"07",X"03",X"04",X"0F",X"04",X"01",X"07",X"0F",X"0F",X"0F",X"0F",X"03",X"05",X"0E",X"0D",X"0F",
		X"90",X"90",X"90",X"90",X"90",X"80",X"80",X"00",X"E7",X"E7",X"E7",X"E7",X"E7",X"63",X"31",X"10",
		X"0F",X"87",X"C3",X"B1",X"90",X"90",X"90",X"90",X"0F",X"0F",X"2F",X"EF",X"E7",X"E7",X"E7",X"E7",
		X"0F",X"FF",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"0F",X"EF",X"E3",X"E3",X"E3",X"E3",X"21",X"01",
		X"0F",X"FF",X"FF",X"F0",X"F0",X"00",X"00",X"F0",X"0F",X"CF",X"8F",X"8F",X"8F",X"C7",X"63",X"F1",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",
		X"E1",X"E1",X"01",X"E1",X"E1",X"E1",X"0F",X"FF",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"FF",
		X"08",X"00",X"07",X"0B",X"00",X"00",X"0F",X"0F",X"03",X"03",X"0F",X"0B",X"03",X"03",X"0B",X"0F",
		X"00",X"07",X"0B",X"00",X"00",X"07",X"0F",X"0F",X"03",X"0F",X"0B",X"03",X"03",X"0B",X"0F",X"0B",
		X"3C",X"3C",X"FC",X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F8",X"FC",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"78",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E1",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"E1",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E1",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"70",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",
		X"78",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"70",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"0F",X"08",X"00",X"07",X"07",X"00",X"08",X"0F",X"0F",X"07",X"03",X"0B",X"0B",X"03",X"07",X"0F",
		X"0F",X"00",X"00",X"07",X"0F",X"00",X"00",X"07",X"0B",X"03",X"07",X"03",X"0B",X"03",X"07",X"0F",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"F0",X"F0",X"F0",X"70",X"70",X"70",X"00",X"00",X"F0",X"F0",X"F0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"D4",X"D4",X"D4",X"D4",X"D4",X"D4",X"1A",X"3C",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"30",X"30",X"90",X"D4",X"D4",X"D4",X"D4",X"D4",
		X"6F",X"6F",X"6F",X"6F",X"6F",X"6F",X"6F",X"6F",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"F0",X"F0",X"0F",X"07",X"37",X"70",X"70",X"70",
		X"F0",X"F0",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"F0",X"F0",X"F0",X"F0",
		X"FF",X"FF",X"FF",X"0F",X"0F",X"F0",X"F0",X"F0",X"FF",X"FF",X"FF",X"0F",X"0F",X"F0",X"F0",X"F0",
		X"C4",X"6A",X"62",X"62",X"62",X"62",X"62",X"66",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"CC",
		X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"33",X"62",X"66",X"D3",X"44",X"D3",X"62",X"62",X"66",
		X"31",X"31",X"31",X"33",X"61",X"33",X"61",X"31",X"EA",X"FB",X"7A",X"62",X"EA",X"62",X"EA",X"62",
		X"31",X"31",X"31",X"31",X"33",X"69",X"31",X"31",X"C2",X"C2",X"C2",X"62",X"62",X"6E",X"D3",X"D3",
		X"62",X"62",X"62",X"62",X"62",X"73",X"70",X"31",X"62",X"62",X"66",X"E2",X"C2",X"EE",X"F0",X"0E",
		X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"33",X"62",X"66",X"D3",X"66",X"D3",X"62",X"62",X"66",
		X"31",X"31",X"31",X"33",X"61",X"33",X"61",X"31",X"62",X"FB",X"7A",X"62",X"EA",X"62",X"EA",X"62",
		X"07",X"07",X"43",X"61",X"77",X"F0",X"31",X"31",X"8F",X"8F",X"43",X"61",X"66",X"7F",X"F0",X"62",
		X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"33",X"62",X"62",X"62",X"62",X"62",X"62",X"62",X"66",
		X"6F",X"6F",X"6F",X"6F",X"5E",X"3C",X"78",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F1",X"F1",X"F1",X"F1",X"F1",X"F0",X"F0",X"F0",X"3C",X"3C",X"0F",X"0F",X"FF",X"F0",X"F0",X"F0",
		X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",
		X"F0",X"F0",X"F0",X"E0",X"F1",X"F1",X"F1",X"F1",X"F0",X"F0",X"F0",X"00",X"00",X"3C",X"3C",X"3C",
		X"F0",X"F0",X"0F",X"0F",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"0F",X"FF",X"F0",X"F0",X"F0",
		X"FF",X"FF",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"FF",X"FF",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"E0",X"E8",X"EC",X"0E",X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"FF",X"F7",X"F3",X"E1",X"E0",X"E0",X"E0",X"E0",X"FF",X"FF",X"FF",X"0F",X"0F",X"F0",X"F0",X"F0",
		X"11",X"EF",X"4C",X"D5",X"E7",X"C4",X"C4",X"C4",X"C4",X"A6",X"C4",X"C4",X"A6",X"C4",X"C4",X"C4",
		X"C4",X"C4",X"C4",X"F7",X"78",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"4C",X"C4",X"C4",X"C4",
		X"62",X"62",X"A6",X"C4",X"92",X"B9",X"C2",X"C4",X"C4",X"C4",X"C4",X"C4",X"4C",X"00",X"00",X"00",
		X"07",X"43",X"70",X"57",X"31",X"31",X"31",X"33",X"EA",X"EA",X"EA",X"EA",X"62",X"62",X"62",X"66",
		X"31",X"31",X"31",X"31",X"77",X"47",X"07",X"07",X"62",X"62",X"62",X"62",X"EA",X"EA",X"EA",X"EA",
		X"FB",X"FE",X"9F",X"9F",X"1F",X"97",X"D3",X"33",X"77",X"F0",X"FF",X"1F",X"1F",X"97",X"D3",X"62",
		X"C4",X"C4",X"D5",X"E7",X"15",X"0E",X"0F",X"97",X"62",X"CC",X"2E",X"0E",X"0C",X"CC",X"62",X"62",
		X"F0",X"F0",X"F0",X"00",X"00",X"E0",X"E0",X"E0",X"F0",X"F0",X"F0",X"70",X"70",X"70",X"70",X"70",
		X"F0",X"F0",X"0F",X"0C",X"34",X"13",X"80",X"F0",X"F0",X"F0",X"0F",X"00",X"F0",X"FF",X"00",X"F0",
		X"87",X"C3",X"E1",X"F0",X"F0",X"E0",X"C0",X"80",X"1E",X"3D",X"7B",X"F7",X"77",X"73",X"31",X"10",
		X"F0",X"84",X"3B",X"3C",X"00",X"F0",X"F0",X"F0",X"F0",X"00",X"FF",X"F0",X"00",X"F0",X"F0",X"F0",
		X"E0",X"E0",X"0E",X"0E",X"FF",X"F0",X"F0",X"F0",X"70",X"70",X"70",X"70",X"70",X"F0",X"F0",X"F0",
		X"97",X"97",X"17",X"30",X"F0",X"F0",X"F0",X"F0",X"3C",X"78",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"97",X"97",X"97",X"97",X"97",X"97",X"97",X"97",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",
		X"F0",X"F0",X"84",X"97",X"97",X"97",X"97",X"97",X"F0",X"F0",X"00",X"00",X"3C",X"3C",X"3C",X"3C",
		X"A1",X"A1",X"A1",X"A1",X"A1",X"B0",X"80",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"00",X"F0",
		X"A1",X"A1",X"A1",X"A1",X"A1",X"A1",X"A1",X"A1",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"FF",X"F7",X"83",X"A1",X"A1",X"A1",X"A1",X"A1",X"FF",X"FF",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"00",X"F0",X"3F",X"3F",X"3F",X"3F",X"3F",X"F3",X"11",X"F0",
		X"31",X"33",X"34",X"31",X"31",X"31",X"31",X"33",X"62",X"62",X"6A",X"66",X"69",X"62",X"62",X"66",
		X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"33",X"69",X"69",X"35",X"42",X"62",X"62",
		X"FF",X"69",X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"31",X"33",X"69",X"69",X"31",
		X"00",X"00",X"00",X"11",X"12",X"31",X"31",X"31",X"31",X"31",X"31",X"FD",X"B5",X"31",X"31",X"31",
		X"F0",X"F0",X"F0",X"F0",X"0F",X"EF",X"EF",X"6F",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"0F",X"00",X"F0",X"FF",X"00",X"F0",X"F0",X"F0",X"0F",X"01",X"E1",X"DA",X"34",X"F0",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"08",X"08",X"0B",X"0F",X"0F",X"0F",
		X"F0",X"00",X"FF",X"F0",X"00",X"F0",X"F0",X"F0",X"F0",X"30",X"88",X"C0",X"00",X"F0",X"F0",X"F0",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"30",X"30",X"00",X"00",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",
		X"F0",X"F0",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"30",X"30",X"30",X"30",X"30",X"30",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"00",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"00",X"F0",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"FF",X"FF",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"FF",X"FF",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"09",X"00",X"06",X"00",X"09",X"0F",X"0F",X"08",X"08",X"0A",X"0A",X"00",X"01",X"0F",X"0B",X"03",
		X"72",X"72",X"72",X"72",X"72",X"72",X"72",X"77",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"FF",
		X"EE",X"A6",X"62",X"62",X"73",X"61",X"72",X"72",X"62",X"62",X"66",X"D3",X"62",X"EA",X"EA",X"EA",
		X"62",X"62",X"26",X"61",X"61",X"62",X"62",X"62",X"62",X"62",X"62",X"62",X"62",X"62",X"62",X"62",
		X"62",X"62",X"62",X"FB",X"E3",X"62",X"62",X"62",X"00",X"00",X"00",X"EE",X"A6",X"62",X"62",X"62",
		X"07",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0B",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"F0",X"F0",X"0F",X"0F",X"FF",X"F1",X"F1",X"F1",X"F0",X"F0",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0B",X"07",X"08",X"0C",
		X"F1",X"F1",X"E1",X"00",X"00",X"F0",X"F0",X"F0",X"3C",X"3C",X"3C",X"34",X"30",X"F0",X"F0",X"F0",
		X"B2",X"B2",X"B2",X"B2",X"B2",X"92",X"81",X"C0",X"34",X"34",X"34",X"34",X"34",X"34",X"3C",X"3C",
		X"E1",X"D2",X"B4",X"B2",X"B2",X"B2",X"B2",X"B2",X"3C",X"34",X"34",X"34",X"34",X"34",X"34",X"34",
		X"E1",X"E1",X"E1",X"E1",X"E1",X"F0",X"F0",X"F0",X"7F",X"7F",X"7F",X"0F",X"0F",X"F0",X"F0",X"F0",
		X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"FF",X"FF",X"FF",X"0F",X"0F",X"E1",X"E1",X"E1",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"30",X"30",X"30",X"30",X"30",X"30",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",
		X"00",X"07",X"0B",X"00",X"00",X"07",X"0F",X"0F",X"03",X"0F",X"0B",X"03",X"03",X"0B",X"0F",X"0B",
		X"87",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",
		X"F7",X"73",X"30",X"30",X"30",X"30",X"30",X"30",X"FF",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"E1",X"D3",X"87",X"F0",X"F0",X"F0",X"F0",X"0F",X"FF",X"FF",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"0F",X"0F",X"09",X"09",X"0F",X"0F",X"0F",X"0D",
		X"07",X"00",X"08",X"0F",X"07",X"07",X"00",X"00",X"0B",X"03",X"07",X"0F",X"0F",X"0B",X"03",X"03",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"00",X"00",X"C0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"E0",X"E0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"70",X"00",
		X"70",X"70",X"70",X"30",X"30",X"10",X"00",X"00",X"E0",X"E0",X"E0",X"C0",X"C0",X"80",X"00",X"00",
		X"04",X"01",X"07",X"0F",X"0F",X"08",X"00",X"05",X"05",X"0E",X"0D",X"0F",X"0B",X"03",X"07",X"0B",
		X"E6",X"E6",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"E6",X"E6",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",
		X"0F",X"F0",X"F0",X"F0",X"F0",X"80",X"E6",X"E6",X"0F",X"F0",X"F0",X"F0",X"F0",X"80",X"E6",X"E6",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"F3",X"F3",X"F3",X"F3",X"F3",X"F3",X"31",X"10",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F3",X"F3",X"F3",X"F3",X"F3",X"F3",X"F3",X"F3",
		X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"1E",X"F3",X"F3",X"F3",X"F3",X"F3",X"F3",X"F3",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"F3",X"F3",X"F3",X"F3",X"F3",X"F3",X"F3",X"10",
		X"FF",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"FF",X"FF",X"F3",X"F3",X"F3",X"F3",X"F3",X"F3",
		X"F0",X"F0",X"F0",X"F0",X"0F",X"FF",X"FF",X"0F",X"F0",X"F0",X"F0",X"F0",X"0F",X"FF",X"FF",X"0F",
		X"FF",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"FF",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"70",X"70",X"70",X"30",X"30",X"30",X"30",X"30",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"30",X"30",X"10",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"70",X"30",X"00",X"00",
		X"0D",X"00",X"00",X"07",X"0F",X"08",X"00",X"07",X"0B",X"03",X"03",X"0B",X"0F",X"07",X"03",X"0B",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"00",X"00",X"E0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"08",X"08",X"0B",
		X"00",X"00",X"07",X"0F",X"07",X"01",X"04",X"0F",X"03",X"03",X"0B",X"0F",X"0F",X"0F",X"0F",X"03",
		X"F1",X"F1",X"F1",X"F1",X"F1",X"F0",X"F0",X"00",X"78",X"78",X"78",X"0F",X"FF",X"F0",X"F0",X"00",
		X"0F",X"F0",X"F0",X"E0",X"F1",X"F1",X"F1",X"F1",X"0F",X"F0",X"F0",X"00",X"78",X"78",X"78",X"78",
		X"6F",X"6F",X"6F",X"6F",X"5E",X"3C",X"78",X"F0",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",
		X"6F",X"6F",X"6F",X"6F",X"6F",X"6F",X"6F",X"6F",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",
		X"F0",X"F0",X"F0",X"F0",X"0F",X"EF",X"EF",X"6F",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",
		X"F0",X"F0",X"90",X"D4",X"D4",X"D4",X"F0",X"F0",X"F0",X"F0",X"90",X"D4",X"D4",X"D4",X"F0",X"F0",
		X"3F",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"CF",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E1",X"E1",X"F1",X"F1",X"F1",X"F1",X"E1",X"E1",
		X"78",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",
		X"70",X"70",X"30",X"10",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"70",X"00",X"00",
		X"30",X"30",X"30",X"10",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"70",X"30",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"C0",X"00",X"C0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"09",X"01",X"0B",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"08",X"00",X"03",X"0B",X"00",X"00",X"07",X"0F",X"07",X"03",X"03",X"06",X"00",X"00",X"0E",
		X"06",X"02",X"0B",X"0F",X"0F",X"00",X"00",X"0F",X"0B",X"03",X"07",X"0F",X"0B",X"03",X"03",X"0B",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"09",X"09",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"F0",X"F0",X"F0",X"0F",X"FF",X"F0",X"F0",X"00",X"70",X"70",X"70",X"70",X"70",X"F0",X"F0",X"00",
		X"0F",X"F0",X"F0",X"00",X"F0",X"F0",X"F0",X"F0",X"0F",X"F0",X"F0",X"70",X"70",X"70",X"70",X"70",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"E1",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E1",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"78",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E1",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"70",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E1",
		X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"70",X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
