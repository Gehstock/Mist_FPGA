library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity spr_rom2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of spr_rom2 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"30",X"70",X"00",X"89",X"66",X"00",X"30",X"F0",X"C0",X"22",X"57",X"0F",X"A3",
		X"60",X"C0",X"80",X"00",X"4C",X"C8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"B0",X"32",X"56",X"21",X"22",X"00",X"00",X"D1",X"F1",X"F1",X"E2",X"5C",X"B8",X"F8",X"00",
		X"55",X"2C",X"CC",X"44",X"F0",X"E1",X"0E",X"00",X"00",X"00",X"00",X"00",X"86",X"08",X"00",X"00",
		X"00",X"00",X"10",X"30",X"30",X"70",X"E0",X"D1",X"60",X"C0",X"C0",X"80",X"80",X"10",X"AE",X"4E",
		X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C3",X"94",X"38",X"D8",X"20",X"22",X"10",X"00",X"23",X"D1",X"E0",X"F1",X"F1",X"F1",X"3E",X"98",
		X"30",X"4C",X"0C",X"F8",X"F0",X"F0",X"C3",X"80",X"00",X"00",X"70",X"E0",X"84",X"08",X"00",X"00",
		X"00",X"00",X"10",X"10",X"30",X"74",X"30",X"70",X"00",X"00",X"00",X"00",X"22",X"10",X"77",X"AE",
		X"00",X"00",X"00",X"00",X"00",X"08",X"11",X"31",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"30",
		X"70",X"71",X"61",X"02",X"10",X"23",X"00",X"00",X"EF",X"08",X"70",X"F0",X"F0",X"30",X"89",X"74",
		X"2A",X"2E",X"54",X"F4",X"B0",X"B0",X"38",X"04",X"60",X"C2",X"C2",X"84",X"08",X"80",X"00",X"00",
		X"00",X"00",X"40",X"62",X"40",X"60",X"60",X"70",X"00",X"00",X"00",X"00",X"20",X"00",X"66",X"07",
		X"00",X"00",X"00",X"00",X"40",X"00",X"66",X"0E",X"00",X"00",X"20",X"64",X"20",X"60",X"60",X"E0",
		X"30",X"30",X"30",X"30",X"10",X"00",X"00",X"00",X"37",X"14",X"38",X"78",X"34",X"CA",X"11",X"00",
		X"CE",X"82",X"C1",X"E1",X"C2",X"35",X"88",X"00",X"C0",X"C0",X"C0",X"C0",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"00",X"22",X"45",X"B9",X"35",X"47",X"52",X"52",
		X"00",X"44",X"2A",X"D9",X"CA",X"2E",X"A4",X"A4",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"40",
		X"20",X"20",X"02",X"02",X"02",X"20",X"00",X"00",X"50",X"50",X"41",X"23",X"03",X"10",X"00",X"00",
		X"60",X"60",X"E8",X"C8",X"0C",X"08",X"00",X"00",X"40",X"40",X"04",X"04",X"04",X"40",X"00",X"00",
		X"00",X"00",X"00",X"02",X"32",X"32",X"12",X"11",X"00",X"00",X"86",X"1E",X"C3",X"1E",X"F8",X"D0",
		X"00",X"CC",X"CE",X"6E",X"6E",X"80",X"49",X"19",X"00",X"00",X"00",X"80",X"80",X"80",X"40",X"40",
		X"60",X"20",X"02",X"01",X"01",X"11",X"00",X"00",X"E3",X"F9",X"64",X"DC",X"80",X"48",X"C0",X"00",
		X"9D",X"1D",X"0C",X"62",X"CA",X"00",X"00",X"00",X"60",X"02",X"65",X"00",X"00",X"00",X"00",X"00",
		X"00",X"10",X"00",X"41",X"43",X"43",X"71",X"30",X"00",X"00",X"84",X"6A",X"2C",X"69",X"3D",X"E3",
		X"00",X"40",X"20",X"10",X"00",X"11",X"08",X"8C",X"00",X"00",X"00",X"00",X"80",X"C8",X"24",X"52",
		X"10",X"40",X"20",X"01",X"00",X"00",X"00",X"00",X"F1",X"70",X"54",X"44",X"4C",X"04",X"02",X"10",
		X"4E",X"AF",X"D7",X"26",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"70",X"03",X"C3",X"43",X"00",X"00",X"0C",X"11",X"26",X"E0",X"2D",X"3C",
		X"00",X"80",X"E0",X"10",X"CD",X"67",X"2A",X"87",X"00",X"00",X"00",X"00",X"E0",X"20",X"00",X"00",
		X"61",X"30",X"00",X"00",X"10",X"00",X"00",X"00",X"F2",X"F9",X"F0",X"00",X"80",X"43",X"00",X"00",
		X"1D",X"CF",X"F3",X"88",X"08",X"C0",X"68",X"20",X"08",X"08",X"88",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"11",X"33",X"30",X"03",X"00",X"00",X"30",X"00",X"FF",X"BF",X"C0",X"3C",
		X"00",X"00",X"00",X"02",X"CE",X"EE",X"FF",X"0F",X"00",X"00",X"00",X"88",X"00",X"00",X"88",X"0C",
		X"03",X"21",X"10",X"00",X"00",X"00",X"00",X"00",X"3C",X"3C",X"7C",X"F0",X"00",X"30",X"00",X"00",
		X"0F",X"F7",X"C0",X"82",X"22",X"0F",X"00",X"00",X"48",X"88",X"00",X"00",X"40",X"48",X"00",X"00",
		X"00",X"00",X"00",X"10",X"00",X"00",X"44",X"01",X"00",X"00",X"30",X"80",X"22",X"00",X"E9",X"96",
		X"20",X"E0",X"80",X"08",X"8C",X"CF",X"2D",X"96",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"88",
		X"B8",X"03",X"03",X"43",X"30",X"00",X"00",X"00",X"78",X"2C",X"78",X"B6",X"E0",X"80",X"00",X"00",
		X"5D",X"71",X"E3",X"81",X"01",X"C2",X"80",X"00",X"00",X"00",X"20",X"84",X"C4",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"20",X"40",X"00",X"10",X"30",X"71",X"C4",X"06",X"55",X"23",X"57",
		X"00",X"00",X"00",X"00",X"26",X"5F",X"BF",X"4C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"31",X"03",X"43",X"41",X"00",X"10",X"00",X"A7",X"79",X"7A",X"1E",X"3E",X"3C",X"E0",X"00",
		X"A8",X"60",X"C0",X"C0",X"81",X"20",X"40",X"00",X"10",X"20",X"40",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"10",X"01",X"02",X"20",X"60",X"00",X"80",X"80",X"00",X"0D",X"45",X"89",X"32",
		X"00",X"00",X"00",X"4A",X"06",X"C2",X"2E",X"5D",X"00",X"00",X"00",X"00",X"00",X"64",X"64",X"68",
		X"11",X"00",X"22",X"10",X"10",X"10",X"00",X"00",X"32",X"F8",X"5A",X"C3",X"0F",X"0F",X"92",X"00",
		X"D5",X"D9",X"E0",X"C4",X"6A",X"80",X"44",X"00",X"04",X"04",X"00",X"80",X"80",X"00",X"00",X"00",
		X"00",X"00",X"20",X"31",X"20",X"31",X"20",X"20",X"00",X"00",X"00",X"32",X"23",X"AB",X"63",X"50",
		X"00",X"00",X"08",X"4C",X"08",X"19",X"68",X"68",X"00",X"00",X"40",X"C8",X"40",X"C8",X"40",X"40",
		X"20",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"C7",X"87",X"43",X"03",X"00",X"00",
		X"78",X"78",X"3E",X"1E",X"2C",X"0C",X"00",X"00",X"40",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"11",X"00",X"10",X"90",X"90",X"90",X"98",
		X"00",X"88",X"00",X"80",X"90",X"90",X"90",X"91",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",
		X"40",X"42",X"36",X"27",X"40",X"00",X"00",X"00",X"2A",X"F2",X"F2",X"5C",X"45",X"45",X"11",X"01",
		X"C5",X"74",X"74",X"A3",X"A2",X"A2",X"88",X"80",X"20",X"24",X"C6",X"4E",X"20",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"20",X"10",X"01",X"11",X"44",X"62",X"62",X"61",X"31",X"30",X"10",X"10",
		X"00",X"00",X"40",X"62",X"20",X"03",X"08",X"34",X"00",X"00",X"00",X"04",X"40",X"20",X"AC",X"24",
		X"04",X"00",X"53",X"03",X"03",X"00",X"00",X"00",X"3A",X"72",X"F2",X"FA",X"88",X"00",X"00",X"00",
		X"94",X"92",X"6B",X"49",X"86",X"24",X"04",X"00",X"D6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"22",X"55",X"30",X"01",X"00",X"40",X"02",X"00",X"20",X"10",X"88",X"C4",X"6A",X"71",X"30",
		X"00",X"02",X"00",X"00",X"25",X"70",X"1C",X"CE",X"00",X"00",X"00",X"80",X"40",X"6E",X"80",X"00",
		X"10",X"00",X"26",X"31",X"01",X"00",X"00",X"00",X"23",X"6A",X"F1",X"78",X"AC",X"4C",X"40",X"00",
		X"A3",X"59",X"A5",X"FB",X"89",X"00",X"00",X"00",X"08",X"00",X"04",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"44",X"E8",X"30",X"11",X"00",X"00",X"00",X"71",X"10",X"88",X"49",X"43",
		X"00",X"28",X"10",X"33",X"28",X"B8",X"1F",X"67",X"00",X"00",X"80",X"48",X"88",X"00",X"00",X"08",
		X"00",X"31",X"00",X"00",X"00",X"01",X"00",X"00",X"32",X"00",X"94",X"04",X"33",X"43",X"03",X"00",
		X"A4",X"43",X"74",X"F3",X"00",X"88",X"08",X"80",X"22",X"8C",X"48",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"74",X"00",X"01",X"00",X"00",X"D1",X"00",X"00",X"F0",
		X"00",X"34",X"37",X"00",X"48",X"81",X"17",X"66",X"00",X"00",X"00",X"00",X"00",X"0C",X"CD",X"33",
		X"47",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"E0",X"00",X"00",X"01",X"00",
		X"E1",X"81",X"D1",X"F8",X"20",X"17",X"16",X"00",X"2E",X"1D",X"CC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"30",X"00",X"00",X"70",X"87",X"22",X"34",X"A4",X"11",X"13",
		X"80",X"08",X"08",X"00",X"C7",X"AE",X"18",X"43",X"00",X"00",X"00",X"08",X"44",X"08",X"2C",X"A2",
		X"11",X"30",X"A8",X"66",X"00",X"00",X"00",X"00",X"70",X"F3",X"88",X"11",X"42",X"80",X"00",X"00",
		X"1D",X"FC",X"F0",X"79",X"23",X"03",X"28",X"00",X"88",X"00",X"00",X"08",X"4C",X"08",X"00",X"00",
		X"00",X"00",X"00",X"10",X"11",X"04",X"00",X"00",X"00",X"44",X"84",X"8C",X"28",X"41",X"59",X"02",
		X"00",X"00",X"22",X"08",X"CF",X"A9",X"52",X"B5",X"00",X"00",X"00",X"00",X"08",X"44",X"00",X"88",
		X"20",X"40",X"00",X"11",X"32",X"45",X"22",X"00",X"10",X"65",X"CA",X"84",X"08",X"01",X"20",X"00",
		X"6A",X"54",X"70",X"05",X"11",X"10",X"02",X"00",X"00",X"80",X"4C",X"8C",X"08",X"00",X"00",X"00",
		X"00",X"00",X"11",X"21",X"21",X"53",X"00",X"04",X"00",X"00",X"00",X"8D",X"33",X"E2",X"62",X"18",
		X"00",X"40",X"06",X"06",X"71",X"B5",X"6A",X"7C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D7",
		X"11",X"01",X"10",X"00",X"00",X"00",X"00",X"00",X"81",X"21",X"16",X"46",X"2D",X"8C",X"62",X"44",
		X"F4",X"C8",X"03",X"20",X"26",X"04",X"00",X"00",X"AC",X"8E",X"04",X"00",X"04",X"00",X"00",X"00",
		X"00",X"00",X"00",X"44",X"52",X"36",X"26",X"40",X"23",X"01",X"45",X"45",X"C5",X"F2",X"F2",X"58",
		X"C4",X"08",X"A2",X"A2",X"32",X"74",X"F4",X"E5",X"00",X"00",X"00",X"22",X"A4",X"C6",X"46",X"20",
		X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"98",X"90",X"18",X"81",X"01",X"01",X"00",X"00",
		X"91",X"90",X"81",X"90",X"80",X"08",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"13",X"00",X"00",X"10",X"03",X"77",X"88",X"88",X"04",
		X"00",X"00",X"80",X"48",X"2C",X"90",X"CD",X"65",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",
		X"13",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"34",X"30",X"98",X"00",X"33",X"01",X"00",X"00",
		X"31",X"11",X"81",X"46",X"8C",X"08",X"00",X"00",X"48",X"08",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"26",X"00",X"10",X"03",X"77",X"10",X"10",X"00",X"C0",
		X"00",X"80",X"48",X"2C",X"80",X"80",X"CC",X"74",X"00",X"00",X"00",X"00",X"00",X"80",X"48",X"68",
		X"26",X"22",X"11",X"00",X"00",X"00",X"00",X"00",X"F0",X"30",X"10",X"10",X"00",X"33",X"01",X"00",
		X"30",X"00",X"80",X"80",X"46",X"8C",X"08",X"00",X"AC",X"8C",X"08",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"22",X"66",X"5C",X"10",X"03",X"77",X"10",X"11",X"10",X"00",X"C8",
		X"80",X"48",X"2C",X"80",X"88",X"80",X"CC",X"75",X"00",X"00",X"00",X"00",X"00",X"40",X"24",X"B4",
		X"5C",X"44",X"22",X"00",X"00",X"00",X"00",X"00",X"F8",X"30",X"10",X"11",X"10",X"00",X"33",X"01",
		X"31",X"00",X"80",X"88",X"80",X"46",X"8C",X"08",X"D6",X"46",X"04",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"31",X"22",X"00",X"00",X"00",X"07",X"08",X"CC",X"00",X"00",X"30",X"11",
		X"00",X"00",X"09",X"04",X"0E",X"0E",X"87",X"40",X"04",X"02",X"03",X"8B",X"06",X"04",X"88",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"30",X"20",X"20",X"00",X"22",X"11",X"00",
		X"C8",X"80",X"08",X"0C",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"13",X"22",X"00",X"00",X"00",X"07",X"0F",X"0C",X"00",X"00",X"30",X"11",
		X"00",X"00",X"09",X"04",X"0E",X"0E",X"87",X"40",X"04",X"02",X"03",X"0B",X"8E",X"8C",X"88",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"30",X"20",X"20",X"00",X"22",X"11",X"00",
		X"C8",X"80",X"08",X"0E",X"06",X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"13",X"22",X"26",X"00",X"00",X"07",X"0F",X"4B",X"EE",X"33",X"30",X"11",
		X"00",X"00",X"38",X"0D",X"1F",X"1F",X"97",X"42",X"0C",X"06",X"07",X"87",X"4A",X"4A",X"08",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"30",X"31",X"30",X"00",X"22",X"11",X"00",
		X"C8",X"84",X"0E",X"0F",X"07",X"56",X"8C",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"03",X"13",X"26",X"44",X"00",X"07",X"0F",X"0F",X"EF",X"FF",X"23",X"20",
		X"00",X"60",X"38",X"2F",X"1F",X"17",X"97",X"73",X"0C",X"0E",X"07",X"87",X"4A",X"4A",X"0C",X"08",
		X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"31",X"21",X"30",X"30",X"00",X"22",X"11",X"00",
		X"EB",X"86",X"0F",X"07",X"23",X"56",X"8C",X"00",X"00",X"00",X"0E",X"0C",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"03",X"13",X"26",X"44",X"00",X"07",X"0F",X"0F",X"EF",X"FF",X"23",X"20",
		X"01",X"41",X"3C",X"0F",X"0F",X"2F",X"B7",X"73",X"0C",X"0E",X"0F",X"87",X"4B",X"4B",X"0E",X"0C",
		X"44",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"31",X"21",X"30",X"30",X"00",X"22",X"11",X"00",
		X"EB",X"87",X"8F",X"33",X"23",X"56",X"8C",X"00",X"08",X"0F",X"0E",X"48",X"80",X"00",X"00",X"00",
		X"00",X"00",X"01",X"12",X"25",X"17",X"26",X"04",X"01",X"1C",X"0E",X"0F",X"EF",X"FF",X"23",X"02",
		X"0F",X"C3",X"3C",X"0F",X"4F",X"2B",X"7F",X"B7",X"00",X"08",X"0C",X"84",X"4A",X"4A",X"0C",X"0E",
		X"44",X"44",X"22",X"22",X"11",X"00",X"00",X"00",X"97",X"29",X"38",X"38",X"00",X"00",X"11",X"00",
		X"27",X"0F",X"33",X"33",X"33",X"67",X"CC",X"00",X"0E",X"4E",X"8E",X"8E",X"0C",X"08",X"00",X"00",
		X"00",X"00",X"01",X"13",X"21",X"17",X"26",X"44",X"03",X"3C",X"C3",X"11",X"EE",X"FF",X"23",X"02",
		X"0F",X"C3",X"3C",X"0F",X"47",X"AB",X"3B",X"B7",X"00",X"0C",X"0E",X"86",X"4B",X"4B",X"2D",X"2D",
		X"44",X"44",X"22",X"22",X"11",X"00",X"00",X"00",X"D7",X"A5",X"B4",X"34",X"02",X"CE",X"33",X"00",
		X"27",X"1F",X"33",X"33",X"23",X"56",X"8E",X"00",X"AD",X"AD",X"4A",X"4A",X"84",X"08",X"00",X"00",
		X"00",X"00",X"01",X"13",X"21",X"17",X"26",X"44",X"03",X"3C",X"C3",X"88",X"FF",X"EF",X"02",X"15",
		X"0F",X"C3",X"3C",X"0F",X"47",X"2B",X"B7",X"53",X"00",X"0C",X"0E",X"86",X"4B",X"4B",X"2D",X"AD",
		X"44",X"44",X"22",X"22",X"11",X"00",X"00",X"00",X"9D",X"4A",X"69",X"24",X"04",X"CE",X"33",X"00",
		X"9B",X"37",X"4F",X"33",X"23",X"56",X"8E",X"00",X"AD",X"2D",X"4A",X"4A",X"84",X"08",X"00",X"00",
		X"F1",X"F1",X"00",X"00",X"00",X"30",X"F3",X"44",X"CF",X"CF",X"03",X"61",X"E0",X"FC",X"30",X"10",
		X"80",X"80",X"18",X"30",X"50",X"80",X"80",X"C0",X"1F",X"C3",X"E1",X"E1",X"C0",X"80",X"80",X"F4",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"70",X"32",X"32",X"64",X"64",X"40",X"00",X"87",X"87",X"B3",X"33",X"33",X"30",X"30",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"00",X"00",X"11",X"33",X"77",X"FF",X"FF",X"FF",
		X"47",X"CD",X"EF",X"EE",X"FF",X"CC",X"8B",X"16",X"3C",X"3C",X"3C",X"3F",X"3F",X"00",X"00",X"09",
		X"77",X"F3",X"30",X"00",X"00",X"1E",X"F1",X"F1",X"EE",X"CD",X"8F",X"C2",X"60",X"87",X"CF",X"CF",
		X"2C",X"18",X"12",X"01",X"43",X"81",X"80",X"80",X"8F",X"F0",X"78",X"3C",X"4C",X"CC",X"0F",X"0E",
		X"8C",X"0C",X"2F",X"2F",X"03",X"01",X"10",X"E0",X"E1",X"E1",X"69",X"2D",X"08",X"80",X"C1",X"C7",
		X"99",X"11",X"01",X"DD",X"17",X"3F",X"7F",X"FF",X"F8",X"F8",X"0F",X"0F",X"47",X"DD",X"EF",X"EE",
		X"1E",X"1E",X"DF",X"FD",X"FD",X"F1",X"F1",X"D3",X"97",X"B7",X"F7",X"F3",X"73",X"71",X"31",X"20",
		X"FF",X"FF",X"FF",X"EE",X"CC",X"88",X"00",X"00",X"CC",X"88",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C3",X"C3",X"C3",X"CF",X"CF",X"01",X"07",X"0F",X"0E",X"1E",X"3C",X"3C",X"78",X"78",X"B0",X"50",
		X"00",X"00",X"80",X"C0",X"E0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",
		X"1F",X"E1",X"E1",X"C3",X"03",X"21",X"3C",X"04",X"20",X"10",X"08",X"0E",X"0F",X"69",X"E1",X"E1",
		X"F0",X"70",X"B0",X"07",X"4B",X"0D",X"1D",X"19",X"E0",X"C3",X"0F",X"0F",X"0F",X"0F",X"F8",X"F8",
		X"F1",X"F1",X"00",X"00",X"00",X"30",X"F3",X"44",X"CF",X"CF",X"03",X"70",X"F0",X"FC",X"30",X"10",
		X"80",X"80",X"90",X"BC",X"10",X"11",X"80",X"C2",X"1F",X"C3",X"E1",X"E1",X"C0",X"80",X"88",X"3C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"70",X"32",X"32",X"64",X"64",X"40",X"00",X"87",X"87",X"B3",X"33",X"33",X"30",X"30",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"00",X"00",X"11",X"33",X"77",X"FF",X"FF",X"FF",
		X"47",X"CD",X"EF",X"EE",X"FF",X"CC",X"8B",X"06",X"3C",X"3C",X"3C",X"3F",X"3F",X"00",X"00",X"89",
		X"77",X"F3",X"30",X"00",X"00",X"1E",X"F1",X"F1",X"EE",X"CD",X"8F",X"C3",X"70",X"87",X"CF",X"CF",
		X"0C",X"08",X"04",X"A9",X"4F",X"81",X"80",X"80",X"07",X"70",X"78",X"3C",X"4C",X"CC",X"0F",X"0E",
		X"8C",X"0C",X"2F",X"2F",X"03",X"01",X"10",X"F0",X"E1",X"E1",X"69",X"1F",X"0C",X"02",X"01",X"03",
		X"99",X"11",X"01",X"D1",X"9F",X"3F",X"7F",X"FF",X"F8",X"F8",X"0F",X"0F",X"47",X"DD",X"EF",X"EE",
		X"1E",X"1E",X"DF",X"FD",X"FD",X"F1",X"F1",X"D3",X"17",X"B7",X"F7",X"F3",X"73",X"71",X"31",X"20",
		X"FF",X"FF",X"FF",X"EE",X"CC",X"88",X"00",X"00",X"CC",X"88",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C3",X"C3",X"C3",X"CF",X"CF",X"01",X"07",X"0F",X"0E",X"1E",X"3C",X"3C",X"78",X"78",X"B0",X"50",
		X"00",X"00",X"80",X"C0",X"E0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",
		X"1F",X"E1",X"E1",X"C3",X"03",X"21",X"3C",X"04",X"E0",X"14",X"08",X"0C",X"1F",X"69",X"E1",X"E1",
		X"F0",X"70",X"B0",X"43",X"0F",X"0D",X"1D",X"19",X"E0",X"C3",X"0F",X"0F",X"0F",X"0F",X"F8",X"F8",
		X"F1",X"F1",X"00",X"00",X"00",X"30",X"F3",X"44",X"CF",X"CF",X"03",X"60",X"E0",X"FC",X"30",X"10",
		X"80",X"80",X"10",X"30",X"52",X"E9",X"F5",X"E2",X"1F",X"C3",X"E1",X"E1",X"C0",X"80",X"00",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"70",X"32",X"32",X"64",X"64",X"40",X"00",X"07",X"87",X"B3",X"33",X"33",X"30",X"30",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"00",X"00",X"11",X"33",X"77",X"FF",X"FF",X"FF",
		X"47",X"CD",X"EF",X"EE",X"FF",X"CC",X"8B",X"06",X"3C",X"3C",X"3C",X"3F",X"3F",X"00",X"00",X"09",
		X"77",X"F3",X"30",X"00",X"00",X"1E",X"F1",X"F1",X"EE",X"CD",X"8F",X"C2",X"70",X"87",X"CF",X"CF",
		X"2E",X"19",X"41",X"43",X"03",X"81",X"80",X"80",X"07",X"70",X"78",X"3C",X"4C",X"CC",X"0F",X"0E",
		X"8C",X"0C",X"2F",X"2F",X"03",X"01",X"00",X"E0",X"E1",X"E1",X"69",X"0C",X"6A",X"D5",X"09",X"03",
		X"99",X"11",X"01",X"D1",X"97",X"3F",X"7F",X"FF",X"F8",X"F8",X"0F",X"0F",X"47",X"DD",X"EF",X"EE",
		X"1E",X"1E",X"DF",X"FD",X"FD",X"F1",X"F1",X"D3",X"17",X"B7",X"F7",X"F3",X"73",X"71",X"31",X"20",
		X"FF",X"FF",X"FF",X"EE",X"CC",X"88",X"00",X"00",X"CC",X"88",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C3",X"C3",X"C3",X"CF",X"CF",X"01",X"07",X"0F",X"0E",X"1E",X"3C",X"3C",X"78",X"78",X"30",X"10",
		X"00",X"00",X"80",X"C0",X"E0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",
		X"0E",X"E1",X"E1",X"C3",X"03",X"21",X"3C",X"04",X"64",X"5C",X"3F",X"2C",X"0E",X"69",X"E1",X"E1",
		X"F0",X"70",X"30",X"03",X"0F",X"0D",X"1D",X"19",X"E0",X"C3",X"0F",X"0F",X"0F",X"0F",X"F8",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"C0",
		X"70",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"F3",X"F0",X"30",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"50",X"80",X"00",X"10",X"30",X"00",X"00",X"C0",X"C0",X"80",X"80",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"30",X"30",X"30",X"71",X"71",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"20",X"30",X"10",X"00",X"00",X"00",X"51",X"31",X"10",X"30",X"F0",X"30",X"00",X"00",
		X"00",X"00",X"00",X"00",X"B0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"00",X"00",X"00",X"20",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"03",X"B0",X"F0",X"43",
		X"00",X"50",X"42",X"4A",X"86",X"96",X"2D",X"2D",X"00",X"00",X"00",X"40",X"08",X"08",X"00",X"00",
		X"20",X"00",X"00",X"00",X"40",X"10",X"00",X"00",X"60",X"16",X"04",X"97",X"86",X"03",X"02",X"04",
		X"42",X"E1",X"68",X"16",X"18",X"00",X"80",X"02",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"60",X"30",X"08",X"00",X"10",X"05",X"03",X"02",X"00",X"10",X"87",X"A5",X"4B",X"69",X"24",
		X"00",X"0C",X"0F",X"69",X"C3",X"C0",X"59",X"AE",X"20",X"40",X"04",X"C0",X"08",X"C2",X"05",X"04",
		X"02",X"03",X"01",X"05",X"01",X"90",X"10",X"20",X"8A",X"89",X"CF",X"11",X"3B",X"0C",X"03",X"00",
		X"09",X"4F",X"0F",X"CF",X"02",X"06",X"09",X"00",X"68",X"A4",X"A4",X"0C",X"42",X"20",X"10",X"00",
		X"00",X"20",X"16",X"91",X"81",X"12",X"00",X"2A",X"43",X"D2",X"69",X"3C",X"86",X"0C",X"3B",X"2A",
		X"B0",X"4B",X"A4",X"0B",X"4D",X"45",X"03",X"2A",X"08",X"84",X"4A",X"86",X"C3",X"43",X"C3",X"06",
		X"2A",X"1D",X"04",X"57",X"05",X"04",X"03",X"00",X"66",X"01",X"0B",X"CC",X"99",X"15",X"02",X"02",
		X"5D",X"3B",X"18",X"47",X"9B",X"8B",X"00",X"00",X"0E",X"0C",X"84",X"88",X"88",X"00",X"00",X"00",
		X"00",X"01",X"04",X"00",X"10",X"10",X"03",X"00",X"58",X"34",X"1C",X"E0",X"2D",X"1A",X"45",X"9F",
		X"0C",X"C0",X"C2",X"21",X"1A",X"5E",X"5E",X"8F",X"00",X"08",X"00",X"0A",X"84",X"0C",X"08",X"08",
		X"01",X"01",X"00",X"01",X"01",X"00",X"00",X"00",X"11",X"08",X"3B",X"0A",X"0D",X"0B",X"01",X"80",
		X"2F",X"45",X"DC",X"9A",X"25",X"0E",X"08",X"0A",X"80",X"82",X"00",X"00",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"16",X"78",X"96",X"07",X"02",
		X"00",X"00",X"11",X"08",X"87",X"69",X"2D",X"9E",X"00",X"00",X"00",X"04",X"08",X"00",X"00",X"11",
		X"08",X"00",X"00",X"00",X"02",X"04",X"00",X"00",X"33",X"02",X"40",X"2D",X"05",X"17",X"02",X"01",
		X"02",X"24",X"0F",X"2F",X"4D",X"8B",X"04",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"10",X"2D",X"4B",X"13",
		X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"37",X"13",X"11",X"00",X"00",X"00",X"00",X"00",
		X"AC",X"0E",X"4E",X"88",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"0C",X"0F",X"03",X"00",X"00",X"00",X"00",
		X"31",X"80",X"2E",X"79",X"49",X"06",X"1D",X"0F",X"04",X"06",X"28",X"0B",X"12",X"76",X"08",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"4B",X"07",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"12",X"78",X"00",X"00",X"00",X"00",X"00",X"00",X"C2",X"87",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"21",X"03",X"43",X"17",X"E6",X"2A",X"08",
		X"C3",X"0F",X"1F",X"7F",X"ED",X"32",X"67",X"77",X"0F",X"0F",X"FB",X"33",X"00",X"F1",X"B3",X"04",
		X"60",X"EE",X"55",X"11",X"01",X"67",X"0E",X"BB",X"70",X"23",X"08",X"2A",X"77",X"88",X"34",X"43",
		X"80",X"48",X"48",X"04",X"04",X"40",X"80",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"3C",X"87",X"0C",X"00",X"00",X"00",X"00",X"86",X"86",X"08",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"0E",X"E1",X"3C",X"00",X"00",X"00",X"00",X"00",X"04",X"0E",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"5A",X"25",X"C3",X"C3",X"97",X"08",X"6A",X"58",X"96",X"0F",X"0F",X"89",X"1C",X"0F",X"0F",X"1E",
		X"80",X"C0",X"48",X"48",X"48",X"84",X"80",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2E",X"1F",X"07",X"03",X"01",X"00",X"00",X"00",
		X"88",X"CC",X"4C",X"7F",X"7F",X"3F",X"3F",X"0F",X"66",X"CC",X"DD",X"FF",X"7F",X"BF",X"EE",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"0F",X"0F",X"07",X"01",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"C3",X"00",X"00",X"00",X"30",X"61",X"87",X"0F",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"21",X"21",X"21",X"21",X"53",X"97",
		X"87",X"1D",X"6E",X"6E",X"CC",X"BB",X"77",X"77",X"7F",X"CC",X"FF",X"FF",X"01",X"AB",X"89",X"EF",
		X"CD",X"EE",X"44",X"01",X"0F",X"16",X"07",X"8A",X"4B",X"4A",X"0E",X"D1",X"2A",X"95",X"1F",X"05",
		X"69",X"5E",X"8D",X"0E",X"02",X"99",X"EF",X"0F",X"80",X"E0",X"68",X"2C",X"68",X"0E",X"2C",X"0C",
		X"13",X"15",X"0E",X"0F",X"0F",X"12",X"00",X"00",X"0B",X"9E",X"0E",X"48",X"80",X"00",X"00",X"00",
		X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"3C",X"0F",X"2F",X"9D",X"CC",X"00",X"00",X"00",X"40",X"C1",X"4B",X"3C",X"8F",
		X"00",X"00",X"00",X"07",X"69",X"96",X"1E",X"5E",X"00",X"00",X"00",X"00",X"0C",X"08",X"08",X"80",
		X"EF",X"47",X"AF",X"6E",X"4C",X"DD",X"CC",X"FF",X"3F",X"2E",X"0E",X"17",X"DF",X"DF",X"47",X"47",
		X"AB",X"23",X"47",X"CF",X"8F",X"8F",X"0F",X"0F",X"C0",X"0E",X"0E",X"C0",X"80",X"80",X"80",X"80",
		X"03",X"03",X"01",X"01",X"01",X"00",X"00",X"00",X"33",X"77",X"19",X"0E",X"0C",X"5F",X"77",X"19",
		X"AB",X"15",X"15",X"DB",X"3B",X"32",X"EC",X"70",X"BB",X"11",X"99",X"4C",X"B7",X"FB",X"AE",X"E6",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"06",X"07",X"03",X"01",X"00",X"00",X"00",
		X"B1",X"FC",X"88",X"3F",X"0F",X"00",X"00",X"00",X"80",X"12",X"AD",X"5A",X"07",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"00",X"00",X"00",X"00",X"70",X"7C",X"3B",X"3F",
		X"02",X"01",X"21",X"71",X"D3",X"C2",X"0E",X"DF",X"00",X"C0",X"F0",X"3C",X"01",X"ED",X"DA",X"83",
		X"10",X"00",X"00",X"00",X"00",X"10",X"30",X"71",X"0C",X"B7",X"84",X"97",X"C7",X"C9",X"89",X"08",
		X"33",X"99",X"EF",X"CF",X"9F",X"2E",X"66",X"0C",X"0F",X"7F",X"2E",X"88",X"00",X"44",X"FF",X"F7",
		X"FF",X"99",X"66",X"67",X"03",X"56",X"DF",X"AA",X"43",X"42",X"0E",X"D1",X"2A",X"95",X"EF",X"05",
		X"08",X"09",X"17",X"0E",X"02",X"99",X"6E",X"48",X"0C",X"E0",X"2C",X"8E",X"AC",X"8E",X"2C",X"8C",
		X"22",X"55",X"66",X"08",X"0F",X"12",X"03",X"02",X"08",X"98",X"03",X"52",X"A4",X"84",X"00",X"00",
		X"B7",X"0F",X"1E",X"08",X"00",X"00",X"00",X"00",X"48",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0C",X"C3",X"F0",X"E1",X"C3",X"4B",X"3F",X"00",X"01",X"5A",X"F0",X"0F",X"AB",X"A9",X"5B",
		X"00",X"0C",X"C3",X"78",X"1E",X"EF",X"AB",X"99",X"00",X"00",X"00",X"0C",X"C2",X"4A",X"4A",X"4A",
		X"BF",X"FF",X"11",X"00",X"66",X"77",X"77",X"33",X"1E",X"1F",X"AD",X"56",X"22",X"AB",X"AB",X"AB",
		X"11",X"23",X"CF",X"B4",X"03",X"01",X"44",X"66",X"86",X"4A",X"E1",X"87",X"E1",X"78",X"78",X"3C",
		X"06",X"06",X"03",X"01",X"01",X"00",X"00",X"00",X"33",X"77",X"11",X"0C",X"0C",X"1F",X"47",X"1D",
		X"8A",X"05",X"05",X"CB",X"2B",X"12",X"EC",X"70",X"F7",X"F7",X"73",X"38",X"94",X"48",X"2E",X"E6",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0C",X"0F",X"07",X"03",X"03",X"44",X"00",
		X"F7",X"CC",X"05",X"0F",X"0F",X"0E",X"00",X"00",X"C5",X"88",X"2C",X"5A",X"0F",X"03",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"10",X"61",X"C3",X"97",X"95",X"08",
		X"00",X"10",X"E1",X"C3",X"5B",X"CA",X"1F",X"8F",X"00",X"C0",X"0D",X"0F",X"0E",X"8F",X"8D",X"0F",
		X"10",X"10",X"10",X"10",X"00",X"01",X"10",X"21",X"6E",X"3B",X"01",X"2B",X"A7",X"85",X"09",X"08",
		X"47",X"8F",X"1F",X"7F",X"08",X"4C",X"55",X"0C",X"0F",X"0F",X"EF",X"33",X"DD",X"CC",X"EE",X"F6",
		X"CF",X"EF",X"99",X"55",X"23",X"03",X"33",X"67",X"17",X"9F",X"AE",X"59",X"AA",X"9D",X"77",X"F7",
		X"CC",X"88",X"00",X"07",X"FF",X"FF",X"77",X"77",X"74",X"60",X"68",X"2C",X"78",X"1E",X"34",X"B8",
		X"4E",X"BF",X"00",X"00",X"01",X"1E",X"0F",X"0E",X"3B",X"9A",X"03",X"5A",X"A4",X"84",X"00",X"00",
		X"B3",X"19",X"0F",X"0F",X"00",X"00",X"00",X"00",X"0E",X"0E",X"0C",X"08",X"00",X"00",X"00",X"00",
		X"00",X"0E",X"87",X"0F",X"08",X"00",X"00",X"00",X"00",X"00",X"70",X"F0",X"5A",X"25",X"21",X"43",
		X"00",X"F0",X"F0",X"0F",X"0F",X"09",X"00",X"22",X"00",X"80",X"C0",X"E0",X"78",X"3C",X"3C",X"2C",
		X"8B",X"34",X"69",X"C3",X"C3",X"06",X"11",X"33",X"F0",X"F0",X"07",X"13",X"03",X"01",X"8B",X"8B",
		X"2F",X"B4",X"0F",X"8B",X"01",X"00",X"08",X"CC",X"2C",X"A4",X"E0",X"F0",X"78",X"3C",X"34",X"34",
		X"84",X"86",X"43",X"0F",X"12",X"01",X"00",X"10",X"66",X"66",X"33",X"3B",X"08",X"0E",X"05",X"49",
		X"4A",X"60",X"16",X"01",X"40",X"07",X"0F",X"00",X"FF",X"33",X"00",X"C0",X"3C",X"07",X"06",X"00",
		X"21",X"41",X"01",X"30",X"20",X"60",X"40",X"80",X"0E",X"87",X"C3",X"43",X"21",X"01",X"20",X"40",
		X"33",X"77",X"22",X"0E",X"1E",X"C3",X"04",X"00",X"66",X"FF",X"00",X"0C",X"4A",X"2D",X"07",X"03",
		X"00",X"00",X"01",X"01",X"03",X"12",X"30",X"52",X"00",X"C3",X"2D",X"E1",X"B0",X"81",X"08",X"45",
		X"00",X"03",X"1E",X"1E",X"96",X"F0",X"07",X"0F",X"0F",X"78",X"87",X"0C",X"3B",X"08",X"0B",X"1A",
		X"42",X"03",X"21",X"21",X"03",X"42",X"42",X"C0",X"03",X"45",X"01",X"07",X"07",X"34",X"03",X"45",
		X"1E",X"78",X"87",X"87",X"07",X"87",X"87",X"0E",X"96",X"78",X"87",X"0F",X"0F",X"09",X"00",X"EE",
		X"00",X"99",X"FF",X"CC",X"89",X"12",X"0F",X"00",X"07",X"05",X"00",X"05",X"4A",X"84",X"1A",X"3D",
		X"66",X"01",X"1E",X"2D",X"6B",X"7B",X"91",X"44",X"69",X"C3",X"C2",X"48",X"48",X"0E",X"2C",X"07",
		X"EE",X"FF",X"FF",X"01",X"12",X"69",X"0F",X"0A",X"06",X"06",X"4B",X"0F",X"1E",X"38",X"38",X"20",
		X"FF",X"77",X"00",X"0F",X"87",X"3C",X"00",X"00",X"07",X"24",X"2C",X"48",X"80",X"00",X"00",X"00",
		X"11",X"D1",X"F1",X"F0",X"3C",X"0F",X"0F",X"0F",X"00",X"07",X"1E",X"69",X"87",X"0F",X"0C",X"0F",
		X"00",X"0E",X"E1",X"78",X"78",X"30",X"0F",X"F0",X"00",X"00",X"08",X"0C",X"86",X"C2",X"4A",X"0E",
		X"96",X"F0",X"E1",X"E1",X"2D",X"03",X"01",X"00",X"5A",X"1E",X"1E",X"0B",X"0B",X"1A",X"12",X"01",
		X"78",X"F0",X"0F",X"09",X"86",X"C2",X"0E",X"0C",X"84",X"86",X"87",X"78",X"3C",X"16",X"07",X"16",
		X"06",X"06",X"03",X"01",X"01",X"00",X"00",X"00",X"33",X"77",X"11",X"0C",X"0C",X"1F",X"47",X"1D",
		X"8A",X"05",X"05",X"CB",X"2B",X"12",X"EC",X"70",X"F7",X"F7",X"73",X"38",X"94",X"48",X"2E",X"E6",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2E",X"1F",X"1F",X"0F",X"03",X"01",X"00",X"00",
		X"F7",X"DD",X"AF",X"0F",X"0F",X"0C",X"00",X"00",X"E7",X"EE",X"3D",X"5A",X"0F",X"03",X"01",X"00",
		X"00",X"00",X"80",X"0E",X"23",X"00",X"00",X"10",X"00",X"00",X"10",X"70",X"C3",X"97",X"95",X"08",
		X"02",X"10",X"F0",X"E1",X"C3",X"E8",X"2D",X"BC",X"10",X"D0",X"C1",X"0F",X"0E",X"8F",X"0D",X"0F",
		X"10",X"10",X"10",X"10",X"00",X"07",X"98",X"61",X"6E",X"3B",X"01",X"2B",X"A7",X"85",X"09",X"08",
		X"47",X"9E",X"3C",X"78",X"E1",X"C2",X"06",X"0C",X"C3",X"E1",X"F0",X"1E",X"01",X"44",X"EE",X"F6",
		X"8F",X"CF",X"01",X"01",X"03",X"12",X"03",X"07",X"52",X"5A",X"0E",X"D1",X"2A",X"85",X"0F",X"07",
		X"C0",X"08",X"00",X"07",X"0F",X"1F",X"77",X"77",X"06",X"60",X"68",X"2C",X"78",X"1E",X"34",X"30",
		X"0E",X"3F",X"00",X"00",X"01",X"1E",X"0F",X"0E",X"0B",X"9A",X"03",X"5A",X"A4",X"84",X"00",X"00",
		X"B3",X"08",X"1E",X"09",X"00",X"00",X"00",X"00",X"9A",X"56",X"A4",X"48",X"08",X"00",X"00",X"00",
		X"00",X"0E",X"87",X"0F",X"08",X"00",X"00",X"00",X"00",X"00",X"70",X"F0",X"5A",X"25",X"21",X"43",
		X"00",X"E0",X"F0",X"1E",X"0F",X"0F",X"01",X"22",X"00",X"00",X"80",X"80",X"C0",X"68",X"3C",X"2C",
		X"8B",X"34",X"69",X"C3",X"C3",X"06",X"11",X"33",X"F0",X"F0",X"07",X"13",X"03",X"10",X"9A",X"9A",
		X"2F",X"B4",X"0F",X"8B",X"01",X"00",X"88",X"84",X"2C",X"A4",X"E0",X"F0",X"78",X"3C",X"34",X"34",
		X"03",X"03",X"01",X"01",X"01",X"00",X"00",X"00",X"33",X"77",X"19",X"0E",X"0C",X"5F",X"77",X"19",
		X"8B",X"05",X"05",X"CB",X"2B",X"12",X"EC",X"70",X"3B",X"19",X"08",X"0C",X"87",X"4B",X"2E",X"E6",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0E",X"07",X"07",X"03",X"01",X"44",X"00",
		X"B1",X"70",X"00",X"0F",X"0F",X"0C",X"00",X"00",X"87",X"16",X"25",X"5A",X"01",X"01",X"00",X"00",
		X"00",X"00",X"80",X"1E",X"23",X"10",X"10",X"10",X"00",X"00",X"00",X"C0",X"F0",X"7C",X"3B",X"3F",
		X"02",X"10",X"30",X"61",X"C3",X"E0",X"2C",X"BC",X"00",X"C0",X"F0",X"3C",X"01",X"ED",X"DA",X"83",
		X"10",X"00",X"00",X"00",X"00",X"07",X"98",X"30",X"0C",X"B7",X"84",X"B4",X"E1",X"C1",X"81",X"08",
		X"03",X"89",X"CF",X"0F",X"87",X"0E",X"06",X"0C",X"0F",X"0F",X"0E",X"88",X"00",X"44",X"FF",X"F7",
		X"FF",X"99",X"66",X"67",X"03",X"16",X"0F",X"8A",X"43",X"42",X"0E",X"D1",X"2A",X"85",X"0F",X"05",
		X"08",X"09",X"07",X"0E",X"02",X"19",X"A6",X"C0",X"0C",X"E0",X"68",X"2C",X"68",X"0E",X"2C",X"48",
		X"02",X"15",X"06",X"08",X"0F",X"12",X"03",X"02",X"08",X"98",X"03",X"52",X"A4",X"84",X"00",X"00",
		X"A7",X"3C",X"1E",X"09",X"00",X"00",X"00",X"00",X"C0",X"80",X"80",X"08",X"08",X"00",X"00",X"00",
		X"00",X"00",X"80",X"F0",X"F0",X"C3",X"49",X"0F",X"00",X"00",X"40",X"F0",X"D2",X"78",X"2D",X"4B",
		X"00",X"01",X"F0",X"78",X"F0",X"B4",X"1E",X"2B",X"00",X"00",X"00",X"80",X"C0",X"C2",X"C2",X"86",
		X"0F",X"0F",X"01",X"00",X"66",X"77",X"77",X"33",X"F0",X"4B",X"2D",X"16",X"02",X"9A",X"8B",X"9A",
		X"23",X"03",X"0F",X"B4",X"03",X"01",X"44",X"66",X"84",X"68",X"E0",X"86",X"E0",X"78",X"78",X"3C",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"19",X"3B",X"2A",X"0C",X"0F",X"07",X"03",X"03",
		X"8B",X"05",X"0D",X"4B",X"AB",X"1C",X"2C",X"78",X"3B",X"19",X"0C",X"0E",X"87",X"4B",X"2E",X"E6",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"03",X"01",X"00",X"00",X"01",X"44",X"88",
		X"B1",X"70",X"0C",X"0F",X"0F",X"08",X"00",X"00",X"87",X"16",X"25",X"5A",X"01",X"01",X"00",X"00",
		X"00",X"00",X"80",X"1E",X"23",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"0F",X"03",X"27",
		X"02",X"00",X"00",X"00",X"14",X"3C",X"2C",X"F0",X"00",X"08",X"1E",X"F0",X"01",X"ED",X"DA",X"83",
		X"00",X"00",X"01",X"00",X"00",X"07",X"88",X"30",X"0C",X"3B",X"00",X"38",X"05",X"29",X"61",X"84",
		X"16",X"8B",X"CD",X"08",X"86",X"0B",X"47",X"67",X"C3",X"84",X"4B",X"16",X"1E",X"0C",X"00",X"80",
		X"CC",X"22",X"08",X"0D",X"0F",X"16",X"07",X"8A",X"43",X"42",X"0E",X"D1",X"2A",X"85",X"0F",X"05",
		X"08",X"09",X"07",X"0E",X"02",X"19",X"86",X"E1",X"0C",X"E0",X"68",X"2C",X"78",X"1E",X"34",X"2C",
		X"02",X"15",X"06",X"08",X"0F",X"12",X"03",X"02",X"08",X"98",X"03",X"52",X"A4",X"84",X"00",X"00",
		X"B4",X"0E",X"0D",X"01",X"00",X"00",X"00",X"00",X"E0",X"40",X"00",X"00",X"08",X"00",X"00",X"00",
		X"00",X"00",X"80",X"F0",X"F0",X"C3",X"59",X"0C",X"00",X"00",X"00",X"43",X"C3",X"4B",X"3C",X"CB",
		X"00",X"01",X"0F",X"0F",X"69",X"F0",X"B4",X"1E",X"00",X"00",X"00",X"00",X"0C",X"0A",X"0A",X"86",
		X"8F",X"34",X"69",X"C2",X"C0",X"19",X"33",X"77",X"F0",X"C3",X"2D",X"16",X"02",X"9A",X"8B",X"9A",
		X"0B",X"03",X"0F",X"B4",X"12",X"01",X"44",X"66",X"C0",X"0E",X"0E",X"C2",X"C0",X"C0",X"68",X"2C",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"06",X"03",X"00",X"00",X"00",X"00",X"00",
		X"88",X"04",X"0C",X"4B",X"2B",X"15",X"04",X"1E",X"66",X"CC",X"4D",X"0F",X"93",X"5B",X"2E",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",
		X"4B",X"30",X"00",X"06",X"08",X"08",X"00",X"00",X"0F",X"1E",X"A5",X"52",X"01",X"01",X"00",X"00",
		X"00",X"00",X"00",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"0F",X"03",X"01",
		X"00",X"00",X"00",X"00",X"04",X"1E",X"3C",X"F0",X"10",X"18",X"1E",X"30",X"61",X"E1",X"D2",X"83",
		X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"30",X"14",X"10",X"30",X"30",X"25",X"29",X"61",X"E1",
		X"96",X"85",X"C2",X"86",X"84",X"3B",X"77",X"77",X"C3",X"84",X"4B",X"1E",X"10",X"9A",X"98",X"9E",
		X"CD",X"EE",X"44",X"01",X"0F",X"16",X"07",X"8A",X"4B",X"4A",X"0E",X"D1",X"2A",X"85",X"0F",X"05",
		X"69",X"5E",X"8D",X"0E",X"02",X"19",X"86",X"E1",X"80",X"E0",X"68",X"2C",X"78",X"1E",X"34",X"2C",
		X"02",X"15",X"06",X"08",X"0F",X"12",X"03",X"02",X"09",X"9A",X"06",X"40",X"84",X"80",X"00",X"00",
		X"B4",X"06",X"01",X"01",X"00",X"00",X"00",X"00",X"E0",X"40",X"00",X"00",X"08",X"00",X"00",X"00",
		X"84",X"84",X"C0",X"F0",X"F0",X"C3",X"59",X"0C",X"00",X"00",X"00",X"43",X"C3",X"4B",X"3C",X"CB",
		X"00",X"01",X"0F",X"0F",X"69",X"F0",X"B4",X"1E",X"00",X"00",X"00",X"00",X"0C",X"0A",X"0A",X"86",
		X"8F",X"34",X"4B",X"86",X"84",X"1D",X"0C",X"0F",X"F0",X"87",X"2D",X"16",X"DE",X"DE",X"47",X"47",
		X"0B",X"03",X"0F",X"A5",X"1E",X"B4",X"A5",X"A5",X"C0",X"0E",X"0E",X"C2",X"0E",X"0A",X"02",X"08",
		X"00",X"01",X"11",X"00",X"00",X"00",X"00",X"00",X"18",X"0C",X"0F",X"8B",X"08",X"00",X"00",X"00",
		X"31",X"80",X"2E",X"79",X"49",X"06",X"1D",X"0F",X"04",X"06",X"28",X"0B",X"12",X"76",X"08",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"4B",X"07",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"12",X"78",X"00",X"00",X"10",X"00",X"00",X"00",X"C2",X"E1",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"21",X"30",X"70",X"43",X"C6",X"82",X"80",
		X"F0",X"C3",X"C3",X"1F",X"6D",X"32",X"67",X"77",X"D2",X"96",X"5A",X"16",X"12",X"F0",X"92",X"16",
		X"60",X"EE",X"45",X"01",X"01",X"16",X"0E",X"BB",X"70",X"23",X"80",X"A2",X"77",X"80",X"34",X"43",
		X"C0",X"68",X"68",X"60",X"60",X"60",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"3C",X"87",X"0C",X"00",X"00",X"00",X"00",X"86",X"86",X"08",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0E",X"0E",X"E1",X"3C",X"00",X"00",X"00",X"00",X"00",X"04",X"0E",X"E1",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"5A",X"25",X"C3",X"C3",X"97",X"08",X"6A",X"58",X"96",X"0F",X"0F",X"89",X"1C",X"0F",X"0F",X"1E",
		X"4C",X"C0",X"6A",X"48",X"48",X"84",X"80",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"00",X"10",X"10",X"20",X"03",X"03",X"01",X"84",X"86",X"28",X"08",X"33",X"77",X"00",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"43",X"07",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"1E",X"00",X"00",X"10",X"00",X"00",X"00",X"0E",X"E1",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"10",X"10",X"00",X"00",X"00",X"00",
		X"1E",X"87",X"C2",X"86",X"84",X"84",X"61",X"A5",X"D2",X"96",X"5A",X"1E",X"12",X"9A",X"12",X"16",
		X"CD",X"EE",X"44",X"01",X"0F",X"16",X"40",X"BB",X"68",X"78",X"0F",X"C1",X"0A",X"82",X"24",X"43",
		X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"3C",X"87",X"0C",X"00",X"00",X"00",X"00",X"86",X"86",X"08",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0E",X"0E",X"E1",X"3C",X"00",X"00",X"00",X"00",X"00",X"04",X"0E",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"4B",X"16",X"4B",X"87",X"84",X"0C",X"0C",X"0F",X"96",X"C2",X"68",X"2D",X"1E",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"08",X"00",X"08",X"80",X"08",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C2",X"2E",X"26",X"9F",X"17",X"13",X"23",X"44",X"46",X"67",X"44",X"00",X"88",X"55",X"6F",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"70",X"34",X"5B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"12",X"12",X"21",X"21",X"21",X"10",X"10",
		X"F0",X"87",X"6F",X"4C",X"4C",X"08",X"0C",X"0E",X"F3",X"C3",X"E9",X"BC",X"3C",X"2D",X"5B",X"87",
		X"EF",X"DF",X"AF",X"03",X"03",X"8F",X"0D",X"00",X"48",X"48",X"2C",X"48",X"0C",X"8C",X"CC",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"70",X"D1",X"7E",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7E",X"78",X"F6",X"3B",X"1D",X"87",X"03",X"12",X"80",X"C0",X"E0",X"E0",X"C0",X"C0",X"E0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"0F",X"0F",X"0F",X"3C",X"F0",X"43",X"C0",X"C0",X"0C",X"6B",X"E3",X"F3",X"3D",X"1E",
		X"8D",X"8D",X"0E",X"0E",X"08",X"91",X"8B",X"44",X"00",X"08",X"01",X"0E",X"07",X"09",X"8F",X"F3",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"07",X"03",X"01",X"00",X"00",
		X"E6",X"7B",X"3C",X"3C",X"69",X"69",X"4B",X"07",X"80",X"88",X"B4",X"3C",X"3C",X"3C",X"3C",X"3C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"00",X"00",X"10",X"30",X"70",X"F0",X"F0",X"F0",
		X"40",X"C2",X"E0",X"E1",X"F0",X"C3",X"84",X"19",X"33",X"33",X"33",X"30",X"30",X"0F",X"0F",X"06",
		X"70",X"FC",X"3F",X"0F",X"0F",X"11",X"F0",X"F0",X"E1",X"C2",X"80",X"CC",X"6B",X"88",X"C0",X"C0",
		X"21",X"12",X"11",X"31",X"6E",X"AE",X"8F",X"8E",X"07",X"AE",X"ED",X"8F",X"1F",X"4C",X"19",X"BB",
		X"66",X"47",X"EE",X"4C",X"37",X"0F",X"1E",X"EF",X"2F",X"2F",X"AF",X"8E",X"06",X"8E",X"0C",X"C0",
		X"96",X"1E",X"0E",X"D2",X"10",X"30",X"70",X"F0",X"F7",X"F7",X"00",X"00",X"48",X"D2",X"E0",X"E0",
		X"11",X"11",X"D0",X"F2",X"F2",X"F2",X"F2",X"D0",X"98",X"B8",X"F8",X"FC",X"7C",X"7E",X"3E",X"2E",
		X"F0",X"F0",X"F0",X"E0",X"C0",X"80",X"00",X"00",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CE",X"CE",X"CE",X"C2",X"C2",X"0E",X"09",X"0E",X"02",X"13",X"37",X"37",X"7F",X"7F",X"BF",X"57",
		X"00",X"00",X"88",X"CC",X"EE",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"CC",
		X"CF",X"23",X"CD",X"02",X"04",X"15",X"04",X"02",X"03",X"16",X"9E",X"57",X"23",X"8B",X"CD",X"03",
		X"FF",X"7F",X"BF",X"0B",X"44",X"03",X"12",X"16",X"EE",X"CF",X"0C",X"00",X"00",X"0F",X"F7",X"F7",
		X"F0",X"F0",X"0F",X"0F",X"0F",X"3C",X"F0",X"43",X"C0",X"C0",X"0C",X"6B",X"E3",X"F3",X"3D",X"1E",
		X"98",X"8C",X"2E",X"7E",X"4C",X"91",X"AA",X"4C",X"33",X"33",X"44",X"88",X"80",X"FF",X"AF",X"F3",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"07",X"03",X"01",X"00",X"00",
		X"E6",X"7B",X"3C",X"3C",X"69",X"69",X"4B",X"07",X"80",X"88",X"B4",X"3C",X"3C",X"3C",X"3C",X"3C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"00",X"00",X"10",X"30",X"70",X"F0",X"F0",X"F0",
		X"40",X"C2",X"E0",X"E1",X"F0",X"C3",X"84",X"19",X"33",X"33",X"33",X"30",X"30",X"0F",X"0F",X"06",
		X"70",X"FC",X"3F",X"0F",X"0F",X"11",X"F0",X"F0",X"E1",X"C2",X"80",X"CC",X"6B",X"88",X"C0",X"C0",
		X"21",X"12",X"11",X"00",X"4C",X"8E",X"8C",X"8E",X"87",X"DD",X"44",X"00",X"40",X"C0",X"00",X"11",
		X"88",X"00",X"00",X"00",X"08",X"0E",X"1F",X"EF",X"EF",X"EF",X"67",X"22",X"00",X"88",X"C0",X"C0",
		X"96",X"1E",X"0E",X"D2",X"10",X"30",X"70",X"F0",X"F7",X"F7",X"00",X"00",X"48",X"D2",X"E0",X"E0",
		X"11",X"11",X"D0",X"F2",X"F2",X"F2",X"F2",X"D0",X"98",X"B8",X"F8",X"FC",X"7C",X"7E",X"3E",X"2E",
		X"F0",X"F0",X"F0",X"E0",X"C0",X"80",X"00",X"00",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CE",X"CE",X"CE",X"C2",X"C2",X"0E",X"09",X"00",X"02",X"13",X"37",X"37",X"7F",X"7F",X"BF",X"56",
		X"00",X"00",X"88",X"CC",X"EE",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"CC",
		X"1E",X"BA",X"8B",X"C0",X"18",X"22",X"DC",X"CC",X"02",X"11",X"00",X"83",X"02",X"67",X"67",X"AB",
		X"FF",X"7F",X"BF",X"0B",X"44",X"03",X"12",X"16",X"EE",X"CF",X"0C",X"00",X"00",X"0F",X"F7",X"F7",
		X"10",X"30",X"31",X"87",X"87",X"43",X"43",X"21",X"F0",X"F0",X"FF",X"78",X"0F",X"2F",X"A7",X"B6",
		X"D0",X"E4",X"E9",X"C2",X"0C",X"0C",X"1B",X"17",X"B9",X"F2",X"60",X"81",X"07",X"69",X"2D",X"0F",
		X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"B6",X"43",X"10",X"00",X"00",X"00",X"00",
		X"D3",X"D3",X"D3",X"97",X"13",X"01",X"00",X"00",X"0F",X"87",X"C3",X"87",X"0F",X"C3",X"21",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"01",X"16",X"3E",X"B6",
		X"00",X"00",X"01",X"17",X"5B",X"D3",X"D3",X"D3",X"00",X"03",X"0D",X"01",X"01",X"C1",X"E1",X"E1",
		X"32",X"30",X"43",X"87",X"87",X"30",X"30",X"10",X"B6",X"B6",X"3E",X"2F",X"0F",X"F0",X"F0",X"F0",
		X"D3",X"D3",X"D3",X"1F",X"0F",X"97",X"D0",X"E1",X"E1",X"E1",X"F3",X"C3",X"A9",X"10",X"14",X"28",
		X"F0",X"90",X"83",X"52",X"4D",X"E9",X"F8",X"F8",X"0F",X"C3",X"0F",X"D3",X"1E",X"5E",X"4F",X"4F",
		X"44",X"80",X"80",X"FF",X"E0",X"F0",X"78",X"78",X"00",X"00",X"00",X"EF",X"11",X"11",X"A2",X"A2",
		X"F8",X"BC",X"BC",X"9E",X"9E",X"F8",X"88",X"08",X"4F",X"4F",X"4F",X"4F",X"5E",X"4C",X"0C",X"00",
		X"3C",X"3C",X"2C",X"C0",X"00",X"00",X"00",X"00",X"C4",X"C4",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"88",X"88",X"88",X"88",X"88",X"88",X"00",X"0C",X"4C",X"5F",X"4E",X"4E",X"5E",X"5E",
		X"00",X"00",X"00",X"00",X"EE",X"11",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"88",X"44",X"44",
		X"C8",X"48",X"AE",X"04",X"D5",X"90",X"44",X"88",X"4E",X"09",X"01",X"8B",X"03",X"07",X"43",X"0F",
		X"E0",X"F0",X"78",X"78",X"FF",X"80",X"80",X"00",X"22",X"22",X"91",X"91",X"EF",X"00",X"00",X"00",
		X"00",X"33",X"70",X"77",X"F0",X"78",X"78",X"78",X"00",X"FF",X"F1",X"FF",X"01",X"FC",X"FC",X"FC",
		X"11",X"FF",X"85",X"97",X"1D",X"A2",X"DC",X"5E",X"FD",X"FE",X"FB",X"F7",X"DC",X"60",X"CF",X"E0",
		X"78",X"78",X"78",X"0F",X"34",X"34",X"03",X"00",X"FC",X"FC",X"FF",X"00",X"F0",X"F0",X"0F",X"00",
		X"96",X"B6",X"B4",X"96",X"96",X"A5",X"0F",X"00",X"E0",X"C3",X"F0",X"E0",X"E1",X"0F",X"0F",X"00",
		X"00",X"33",X"70",X"77",X"F0",X"78",X"78",X"78",X"00",X"FF",X"F0",X"FF",X"00",X"FC",X"FC",X"FC",
		X"00",X"FF",X"95",X"96",X"B6",X"B4",X"96",X"96",X"00",X"FF",X"FF",X"E1",X"F0",X"E0",X"C3",X"E0",
		X"78",X"78",X"78",X"0F",X"34",X"07",X"00",X"00",X"FC",X"FC",X"FF",X"00",X"F0",X"0F",X"00",X"00",
		X"96",X"B6",X"B4",X"96",X"97",X"0F",X"04",X"00",X"E0",X"C3",X"F0",X"AC",X"47",X"EE",X"B9",X"FF",
		X"80",X"DC",X"01",X"0B",X"56",X"8E",X"0F",X"9E",X"66",X"90",X"0F",X"78",X"F0",X"F0",X"78",X"F0",
		X"F3",X"F3",X"3F",X"F3",X"E0",X"83",X"83",X"83",X"88",X"88",X"88",X"FF",X"F1",X"F1",X"F1",X"F1",
		X"8E",X"0F",X"9E",X"46",X"0F",X"0F",X"0C",X"00",X"F0",X"78",X"F0",X"F0",X"C3",X"0C",X"00",X"00",
		X"83",X"83",X"83",X"E0",X"0F",X"00",X"00",X"00",X"F1",X"F1",X"F1",X"79",X"1F",X"00",X"00",X"00",
		X"00",X"CC",X"FF",X"0F",X"D6",X"8E",X"0F",X"9E",X"00",X"00",X"CC",X"F3",X"F0",X"F0",X"78",X"F1",
		X"00",X"00",X"00",X"FF",X"E0",X"83",X"83",X"8B",X"00",X"00",X"00",X"FF",X"79",X"F1",X"F1",X"F1",
		X"8E",X"0F",X"DF",X"F7",X"33",X"FF",X"F7",X"EA",X"CE",X"EF",X"FE",X"EE",X"CC",X"FF",X"0A",X"17",
		X"8B",X"83",X"83",X"33",X"00",X"FF",X"F3",X"73",X"F1",X"F1",X"31",X"19",X"11",X"88",X"88",X"88",
		X"11",X"31",X"30",X"88",X"8B",X"44",X"44",X"22",X"FF",X"FF",X"F0",X"77",X"0F",X"24",X"A4",X"B4",
		X"EE",X"EA",X"E7",X"FF",X"0F",X"12",X"12",X"92",X"95",X"86",X"8B",X"7F",X"0F",X"67",X"23",X"01",
		X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"34",X"BC",X"46",X"11",X"00",X"00",X"00",X"00",
		X"D2",X"D2",X"D2",X"9A",X"12",X"01",X"00",X"00",X"01",X"81",X"C1",X"81",X"01",X"CD",X"23",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"01",X"17",X"3D",X"BD",
		X"00",X"00",X"01",X"16",X"5E",X"DE",X"DE",X"DE",X"00",X"03",X"0F",X"0F",X"0F",X"CF",X"EF",X"EF",
		X"31",X"37",X"44",X"88",X"88",X"31",X"31",X"11",X"BD",X"BD",X"35",X"24",X"00",X"FF",X"FF",X"FF",
		X"DE",X"DE",X"DE",X"12",X"00",X"98",X"DF",X"EE",X"EF",X"EF",X"FC",X"8F",X"87",X"0F",X"16",X"14",
		X"C2",X"16",X"0C",X"FF",X"0F",X"F7",X"F7",X"F7",X"03",X"C3",X"03",X"DE",X"1F",X"5B",X"4A",X"4A",
		X"44",X"80",X"80",X"F0",X"EF",X"FF",X"77",X"77",X"00",X"00",X"00",X"E1",X"1E",X"1E",X"AC",X"AC",
		X"F7",X"B3",X"B3",X"91",X"91",X"F7",X"87",X"08",X"4A",X"4A",X"4A",X"4A",X"5B",X"48",X"0C",X"00",
		X"33",X"33",X"23",X"CE",X"00",X"00",X"00",X"00",X"C8",X"C8",X"08",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"87",X"87",X"87",X"87",X"87",X"87",X"00",X"0C",X"48",X"5A",X"4B",X"4B",X"5B",X"5B",
		X"00",X"00",X"00",X"00",X"E0",X"1E",X"0F",X"CF",X"00",X"00",X"00",X"00",X"00",X"80",X"48",X"48",
		X"C7",X"C7",X"F0",X"0F",X"0F",X"3F",X"97",X"C2",X"5B",X"4A",X"C2",X"0E",X"1E",X"CF",X"CF",X"03",
		X"EF",X"FF",X"77",X"77",X"F0",X"80",X"80",X"00",X"2C",X"2C",X"9E",X"9E",X"E1",X"00",X"00",X"00",
		X"00",X"30",X"00",X"70",X"00",X"80",X"80",X"80",X"00",X"F0",X"00",X"F0",X"0F",X"C0",X"C0",X"C0",
		X"00",X"F0",X"52",X"60",X"60",X"40",X"60",X"60",X"00",X"F0",X"F0",X"00",X"00",X"01",X"10",X"01",
		X"80",X"80",X"80",X"F0",X"40",X"40",X"30",X"00",X"C0",X"C0",X"F0",X"0F",X"00",X"00",X"F0",X"00",
		X"60",X"60",X"40",X"60",X"60",X"70",X"F0",X"00",X"01",X"10",X"00",X"01",X"10",X"F0",X"F0",X"00",
		X"00",X"30",X"00",X"70",X"00",X"80",X"80",X"80",X"00",X"F0",X"00",X"F0",X"0F",X"C0",X"C0",X"C0",
		X"00",X"F0",X"52",X"60",X"60",X"40",X"60",X"60",X"00",X"F0",X"F0",X"00",X"00",X"01",X"10",X"01",
		X"80",X"80",X"80",X"F0",X"40",X"70",X"03",X"00",X"C0",X"C0",X"F0",X"0F",X"00",X"F0",X"0F",X"00",
		X"60",X"60",X"40",X"60",X"60",X"F0",X"4F",X"00",X"01",X"10",X"00",X"01",X"10",X"F0",X"0F",X"00",
		X"4B",X"E4",X"4A",X"F0",X"4A",X"87",X"F0",X"86",X"66",X"00",X"F0",X"00",X"00",X"00",X"80",X"00",
		X"30",X"30",X"F0",X"30",X"01",X"07",X"07",X"07",X"80",X"80",X"80",X"F0",X"10",X"98",X"98",X"98",
		X"87",X"F0",X"86",X"4B",X"F0",X"F0",X"C0",X"00",X"00",X"80",X"00",X"00",X"30",X"C0",X"00",X"00",
		X"07",X"07",X"07",X"01",X"F0",X"00",X"00",X"00",X"98",X"DC",X"DC",X"5C",X"90",X"00",X"00",X"00",
		X"00",X"C0",X"F0",X"F0",X"5B",X"87",X"F0",X"97",X"00",X"00",X"C0",X"30",X"00",X"88",X"80",X"00",
		X"00",X"00",X"00",X"F0",X"01",X"07",X"07",X"07",X"00",X"00",X"00",X"F0",X"18",X"98",X"98",X"98",
		X"87",X"F0",X"97",X"C3",X"F0",X"5B",X"F5",X"5B",X"88",X"80",X"00",X"8B",X"87",X"F0",X"CF",X"78",
		X"07",X"07",X"07",X"3C",X"0F",X"F0",X"FC",X"7C",X"DC",X"DC",X"3E",X"1E",X"1E",X"80",X"80",X"80",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F0",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"10",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
