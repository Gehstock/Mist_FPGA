library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity prom_ic39 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of prom_ic39 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7C",X"12",X"12",X"12",X"7E",X"7C",X"00",
		X"00",X"34",X"4A",X"4A",X"4A",X"7E",X"7E",X"00",X"00",X"24",X"42",X"42",X"42",X"7E",X"3C",X"00",
		X"00",X"3C",X"42",X"42",X"42",X"7E",X"7E",X"00",X"00",X"42",X"4A",X"4A",X"4A",X"7E",X"7E",X"00",
		X"00",X"02",X"0A",X"0A",X"0A",X"7E",X"7E",X"00",X"00",X"34",X"52",X"52",X"42",X"7E",X"3C",X"00",
		X"00",X"7E",X"08",X"08",X"08",X"7E",X"7E",X"00",X"00",X"42",X"42",X"7E",X"7E",X"42",X"42",X"00",
		X"00",X"7E",X"7E",X"7E",X"40",X"40",X"30",X"00",X"00",X"42",X"24",X"18",X"08",X"7E",X"7E",X"00",
		X"00",X"40",X"40",X"40",X"40",X"7E",X"7E",X"00",X"00",X"7E",X"02",X"7C",X"02",X"7E",X"7E",X"00",
		X"00",X"7E",X"20",X"18",X"04",X"7E",X"7E",X"00",X"00",X"3C",X"42",X"42",X"42",X"7E",X"3C",X"00",
		X"00",X"0C",X"12",X"12",X"12",X"7E",X"7E",X"00",X"00",X"40",X"3C",X"62",X"42",X"7E",X"3C",X"00",
		X"00",X"44",X"2A",X"1A",X"0A",X"7E",X"7E",X"00",X"00",X"34",X"72",X"4A",X"4A",X"4E",X"2C",X"00",
		X"00",X"02",X"02",X"7E",X"7E",X"02",X"02",X"00",X"00",X"3E",X"40",X"40",X"40",X"7E",X"7E",X"00",
		X"00",X"1E",X"20",X"40",X"20",X"3E",X"1E",X"00",X"00",X"3E",X"40",X"38",X"40",X"7E",X"3E",X"00",
		X"00",X"42",X"26",X"1C",X"38",X"74",X"62",X"00",X"00",X"06",X"08",X"70",X"08",X"0E",X"06",X"00",
		X"00",X"42",X"46",X"4E",X"5A",X"72",X"62",X"00",X"00",X"00",X"00",X"42",X"42",X"7E",X"00",X"00",
		X"00",X"00",X"00",X"7E",X"42",X"42",X"00",X"00",X"00",X"00",X"42",X"66",X"3C",X"18",X"00",X"00",
		X"00",X"00",X"00",X"18",X"3C",X"66",X"42",X"00",X"00",X"00",X"24",X"18",X"7E",X"18",X"24",X"00",
		X"00",X"00",X"3C",X"46",X"4A",X"52",X"3C",X"00",X"00",X"00",X"40",X"40",X"7E",X"42",X"44",X"00",
		X"00",X"00",X"64",X"4A",X"52",X"62",X"44",X"00",X"00",X"00",X"34",X"4A",X"4A",X"4A",X"42",X"00",
		X"00",X"00",X"08",X"7E",X"08",X"08",X"0E",X"00",X"00",X"00",X"30",X"4A",X"4A",X"4A",X"4E",X"00",
		X"00",X"00",X"30",X"4A",X"4A",X"4A",X"3C",X"00",X"00",X"00",X"06",X"1A",X"32",X"62",X"06",X"00",
		X"00",X"00",X"34",X"4A",X"4A",X"4A",X"34",X"00",X"00",X"00",X"3C",X"52",X"52",X"52",X"0C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"00",X"00",X"08",X"08",X"08",X"08",X"08",X"00",
		X"3C",X"42",X"81",X"81",X"81",X"81",X"42",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"09",X"51",X"01",X"02",X"00",
		X"FC",X"E0",X"70",X"38",X"1C",X"3E",X"00",X"00",X"00",X"3E",X"1C",X"38",X"70",X"E0",X"FC",X"9F",
		X"E0",X"70",X"38",X"7C",X"00",X"00",X"00",X"00",X"00",X"7C",X"38",X"70",X"E0",X"FC",X"9F",X"FC",
		X"70",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"70",X"E0",X"FC",X"9F",X"FC",X"E0",
		X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"70",X"E0",X"FC",X"9F",X"FC",X"E0",X"70",
		X"70",X"E0",X"FC",X"9F",X"FC",X"E0",X"70",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",
		X"E0",X"FC",X"9F",X"FC",X"E0",X"70",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"70",
		X"FC",X"9F",X"FC",X"E0",X"70",X"38",X"7C",X"00",X"00",X"00",X"00",X"00",X"7C",X"38",X"70",X"E0",
		X"9F",X"FC",X"E0",X"70",X"38",X"1C",X"3E",X"00",X"00",X"00",X"3E",X"1C",X"38",X"70",X"E0",X"FC",
		X"7F",X"C7",X"0E",X"1C",X"38",X"70",X"FC",X"00",X"FC",X"70",X"38",X"1C",X"0E",X"C7",X"7F",X"E3",
		X"CE",X"1C",X"38",X"70",X"FC",X"00",X"00",X"00",X"FC",X"70",X"38",X"1C",X"CE",X"7F",X"E3",X"7F",
		X"3C",X"78",X"FC",X"00",X"00",X"00",X"00",X"00",X"FC",X"78",X"3C",X"DE",X"7F",X"E3",X"7F",X"DE",
		X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"78",X"FC",X"7F",X"E3",X"7F",X"FC",X"78",
		X"78",X"FC",X"7F",X"E3",X"7F",X"FC",X"78",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",
		X"DE",X"7F",X"E3",X"7F",X"DE",X"3C",X"78",X"FC",X"00",X"00",X"00",X"00",X"00",X"FC",X"78",X"3C",
		X"7F",X"E3",X"7F",X"CE",X"1C",X"38",X"70",X"FC",X"00",X"00",X"00",X"FC",X"70",X"38",X"1C",X"CE",
		X"E3",X"7F",X"C7",X"0E",X"1C",X"38",X"70",X"FC",X"00",X"FC",X"70",X"38",X"1C",X"0E",X"C7",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"00",X"00",X"00",
		X"00",X"00",X"00",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"00",X"00",X"00",X"00",X"0F",X"0F",X"00",X"00",
		X"00",X"00",X"0F",X"0F",X"00",X"00",X"00",X"00",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",
		X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7E",X"CC",X"38",X"FE",X"38",X"CC",X"7E",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",
		X"78",X"3E",X"78",X"9C",X"0E",X"FF",X"3E",X"00",X"00",X"00",X"00",X"00",X"3E",X"FF",X"0E",X"9C",
		X"38",X"5C",X"4E",X"87",X"0F",X"3E",X"FC",X"00",X"FC",X"3E",X"0F",X"87",X"4E",X"5C",X"38",X"3E",
		X"0E",X"FF",X"3E",X"00",X"00",X"00",X"00",X"00",X"3E",X"FF",X"0E",X"9C",X"78",X"3E",X"78",X"9C",
		X"FF",X"1C",X"38",X"FE",X"38",X"1C",X"FF",X"00",X"82",X"92",X"D6",X"FE",X"FE",X"BA",X"92",X"92",
		X"FF",X"38",X"1C",X"7F",X"1C",X"38",X"FF",X"00",X"92",X"92",X"BA",X"FE",X"FE",X"D6",X"92",X"82",
		X"00",X"00",X"10",X"38",X"10",X"00",X"00",X"00",X"00",X"08",X"30",X"7C",X"30",X"08",X"00",X"00",
		X"00",X"0C",X"38",X"FE",X"38",X"0C",X"00",X"00",X"1E",X"0C",X"38",X"FE",X"38",X"0C",X"1E",X"00",
		X"3D",X"3E",X"5C",X"18",X"10",X"20",X"00",X"00",X"00",X"00",X"04",X"08",X"18",X"3A",X"74",X"B8",
		X"7C",X"3A",X"18",X"08",X"04",X"00",X"00",X"00",X"00",X"20",X"10",X"18",X"5C",X"2E",X"1D",X"BC",
		X"BC",X"1D",X"2E",X"5C",X"18",X"10",X"20",X"00",X"00",X"00",X"00",X"04",X"08",X"18",X"3A",X"7C",
		X"74",X"3A",X"18",X"08",X"04",X"00",X"00",X"00",X"00",X"20",X"10",X"18",X"5C",X"3E",X"3D",X"B8",
		X"18",X"F8",X"F0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"38",X"38",X"18",
		X"FE",X"BA",X"92",X"92",X"00",X"10",X"28",X"10",X"00",X"00",X"00",X"00",X"82",X"92",X"D6",X"FE",
		X"18",X"1F",X"0F",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"1C",X"1C",X"18",
		X"00",X"00",X"00",X"00",X"00",X"0A",X"0E",X"00",X"00",X"C3",X"66",X"BC",X"E7",X"BC",X"66",X"C3",
		X"F0",X"F8",X"3C",X"0C",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"C0",
		X"A0",X"C0",X"E0",X"F0",X"70",X"38",X"18",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"DC",X"0C",X"0C",X"1C",X"18",X"10",X"00",X"00",X"00",X"00",X"00",X"80",X"E8",X"F0",X"78",
		X"00",X"40",X"88",X"70",X"E0",X"C0",X"80",X"00",X"80",X"40",X"E0",X"F0",X"F8",X"C4",X"20",X"00",
		X"00",X"40",X"88",X"F0",X"E0",X"C0",X"80",X"00",X"80",X"40",X"E0",X"F0",X"B8",X"44",X"20",X"00",
		X"F0",X"C0",X"80",X"E0",X"80",X"C0",X"F0",X"00",X"F0",X"80",X"C2",X"F5",X"C2",X"80",X"F0",X"00",
		X"FE",X"D6",X"92",X"82",X"00",X"00",X"00",X"00",X"10",X"28",X"10",X"00",X"92",X"92",X"BA",X"FE",
		X"7C",X"E0",X"C0",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"C0",X"E0",X"7C",X"F0",
		X"0F",X"0C",X"10",X"00",X"00",X"00",X"00",X"00",X"70",X"38",X"1C",X"1C",X"0E",X"0E",X"07",X"07",
		X"07",X"03",X"01",X"03",X"03",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"1C",X"1F",
		X"00",X"00",X"01",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"0F",X"1C",X"00",
		X"02",X"04",X"0E",X"1F",X"3F",X"47",X"08",X"01",X"00",X"04",X"22",X"1D",X"0F",X"07",X"02",X"01",
		X"02",X"04",X"0F",X"1F",X"3B",X"45",X"08",X"01",X"00",X"04",X"23",X"1F",X"0F",X"07",X"02",X"01",
		X"0F",X"01",X"43",X"AF",X"43",X"01",X"0F",X"00",X"0F",X"03",X"01",X"07",X"01",X"03",X"0F",X"00",
		X"78",X"FA",X"DC",X"9F",X"BF",X"33",X"43",X"1E",X"1E",X"47",X"33",X"BF",X"9F",X"DC",X"FA",X"78",
		X"00",X"00",X"01",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"01",X"00",X"00",X"01",
		X"C0",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"C0",X"00",
		X"E8",X"F0",X"60",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"20",X"C0",X"C4",
		X"C4",X"C0",X"20",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"E0",X"F0",X"C8",
		X"C8",X"F0",X"E0",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"20",X"C0",X"C4",
		X"C4",X"C0",X"20",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"60",X"F0",X"E8",
		X"C0",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0C",X"3C",X"F8",X"F0",
		X"38",X"70",X"F0",X"E0",X"C0",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"18",X"18",
		X"78",X"F0",X"E8",X"80",X"00",X"00",X"00",X"00",X"00",X"10",X"18",X"18",X"0C",X"0C",X"DC",X"F8",
		X"07",X"0E",X"1C",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"1C",X"0E",X"07",X"1F",
		X"23",X"03",X"04",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"07",X"0F",X"13",
		X"17",X"0F",X"06",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"04",X"03",X"23",
		X"23",X"03",X"04",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"06",X"0F",X"17",
		X"13",X"0F",X"07",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"04",X"03",X"23",
		X"07",X"07",X"0E",X"0E",X"1C",X"1C",X"38",X"70",X"00",X"00",X"00",X"00",X"20",X"10",X"0C",X"0F",
		X"04",X"03",X"03",X"01",X"03",X"07",X"1F",X"7C",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"1C",X"0F",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"01",X"00",X"00",
		X"00",X"60",X"60",X"00",X"08",X"00",X"00",X"00",X"40",X"00",X"08",X"1C",X"08",X"00",X"00",X"00",
		X"18",X"7E",X"CF",X"BD",X"BD",X"F3",X"7F",X"3C",X"08",X"24",X"01",X"84",X"50",X"09",X"22",X"08",
		X"FF",X"FF",X"FE",X"FE",X"FC",X"FC",X"F8",X"E0",X"A1",X"29",X"23",X"B3",X"77",X"77",X"FF",X"FF",
		X"FF",X"FF",X"77",X"77",X"B3",X"23",X"A9",X"25",X"E0",X"F8",X"FC",X"FC",X"FE",X"FE",X"FF",X"FF",
		X"8C",X"C2",X"C0",X"F0",X"3A",X"38",X"0C",X"46",X"C4",X"80",X"FC",X"FF",X"F0",X"82",X"F0",X"38",
		X"05",X"1C",X"78",X"F2",X"F0",X"C4",X"98",X"72",X"E2",X"80",X"0C",X"1E",X"1A",X"8C",X"00",X"00",
		X"F8",X"78",X"B0",X"60",X"F3",X"DB",X"D8",X"30",X"0C",X"1E",X"0C",X"80",X"C0",X"C0",X"64",X"B2",
		X"00",X"00",X"08",X"1C",X"3E",X"36",X"22",X"00",X"00",X"00",X"0E",X"1C",X"38",X"1C",X"0E",X"00",
		X"00",X"00",X"3E",X"3E",X"3E",X"3E",X"3E",X"00",X"60",X"70",X"78",X"7C",X"3C",X"1C",X"0C",X"04",
		X"20",X"30",X"38",X"1C",X"0E",X"06",X"02",X"00",X"00",X"10",X"38",X"7C",X"FE",X"7C",X"38",X"10",
		X"FF",X"FF",X"7F",X"7F",X"3F",X"3F",X"1F",X"07",X"A4",X"85",X"D4",X"C6",X"EE",X"EF",X"FF",X"FF",
		X"FF",X"FF",X"EF",X"EE",X"C6",X"D4",X"84",X"A5",X"07",X"1F",X"3F",X"3F",X"7F",X"7F",X"FF",X"FF",
		X"3F",X"3D",X"2D",X"66",X"26",X"43",X"12",X"20",X"3B",X"3B",X"75",X"EE",X"F5",X"3B",X"7B",X"9F",
		X"20",X"09",X"2C",X"84",X"44",X"ED",X"6D",X"7F",X"77",X"27",X"03",X"20",X"00",X"08",X"1C",X"08",
		X"EF",X"F9",X"77",X"37",X"7C",X"DF",X"EB",X"7D",X"20",X"41",X"04",X"31",X"7B",X"7E",X"33",X"6F",
		X"00",X"00",X"22",X"36",X"3E",X"1C",X"08",X"00",X"00",X"38",X"1C",X"0E",X"1C",X"38",X"00",X"00",
		X"00",X"60",X"78",X"3C",X"1E",X"0E",X"06",X"00",X"00",X"38",X"38",X"38",X"18",X"18",X"38",X"38",
		X"00",X"00",X"07",X"7F",X"FE",X"E0",X"00",X"00",X"03",X"07",X"77",X"DD",X"FF",X"F6",X"3C",X"00",
		X"9E",X"F8",X"E0",X"70",X"38",X"7C",X"00",X"00",X"00",X"00",X"00",X"7C",X"38",X"70",X"E0",X"F8",
		X"79",X"3F",X"67",X"0E",X"1C",X"38",X"7C",X"00",X"00",X"00",X"7C",X"38",X"1C",X"0E",X"67",X"3F",
		X"90",X"20",X"40",X"80",X"00",X"00",X"00",X"00",X"34",X"34",X"34",X"64",X"68",X"68",X"C8",X"D0",
		X"D0",X"C8",X"68",X"68",X"64",X"34",X"34",X"34",X"00",X"00",X"00",X"00",X"80",X"40",X"20",X"90",
		X"34",X"64",X"C8",X"90",X"20",X"C0",X"00",X"00",X"0D",X"0D",X"0D",X"0D",X"19",X"1A",X"1A",X"32",
		X"32",X"1A",X"1A",X"19",X"0D",X"0D",X"0D",X"0D",X"00",X"00",X"C0",X"20",X"90",X"C8",X"64",X"34",
		X"09",X"04",X"02",X"01",X"00",X"00",X"00",X"00",X"2C",X"2C",X"2C",X"26",X"16",X"16",X"13",X"0B",
		X"0B",X"03",X"06",X"06",X"26",X"2C",X"2C",X"2C",X"00",X"00",X"00",X"00",X"01",X"02",X"04",X"09",
		X"2C",X"26",X"13",X"09",X"04",X"03",X"00",X"00",X"B0",X"B0",X"B0",X"B0",X"98",X"58",X"58",X"4C",
		X"4C",X"58",X"50",X"98",X"B0",X"B0",X"B0",X"B0",X"00",X"00",X"03",X"04",X"09",X"13",X"26",X"2C",
		X"03",X"1F",X"FC",X"E1",X"0E",X"F0",X"00",X"00",X"C0",X"F8",X"3F",X"87",X"70",X"0F",X"00",X"00",
		X"00",X"00",X"0F",X"70",X"87",X"3F",X"F8",X"C0",X"00",X"00",X"F0",X"0E",X"E1",X"FC",X"1F",X"03",
		X"00",X"00",X"01",X"0F",X"FE",X"F0",X"07",X"F8",X"00",X"00",X"80",X"F0",X"7F",X"0F",X"E0",X"1F",
		X"1F",X"E0",X"0F",X"7F",X"F0",X"80",X"00",X"00",X"F8",X"07",X"F0",X"FE",X"0F",X"01",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
